module basic_750_5000_1000_50_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_146,In_507);
and U1 (N_1,In_522,In_353);
nand U2 (N_2,In_470,In_52);
nand U3 (N_3,In_164,In_580);
xnor U4 (N_4,In_307,In_655);
nand U5 (N_5,In_729,In_492);
xnor U6 (N_6,In_700,In_114);
nor U7 (N_7,In_202,In_546);
nor U8 (N_8,In_160,In_620);
xnor U9 (N_9,In_721,In_211);
or U10 (N_10,In_268,In_531);
or U11 (N_11,In_319,In_683);
nand U12 (N_12,In_446,In_709);
nor U13 (N_13,In_14,In_90);
and U14 (N_14,In_107,In_624);
xnor U15 (N_15,In_565,In_714);
or U16 (N_16,In_13,In_647);
and U17 (N_17,In_725,In_664);
and U18 (N_18,In_255,In_738);
xor U19 (N_19,In_460,In_554);
nand U20 (N_20,In_277,In_48);
xnor U21 (N_21,In_430,In_359);
nand U22 (N_22,In_734,In_465);
or U23 (N_23,In_555,In_458);
or U24 (N_24,In_448,In_409);
or U25 (N_25,In_590,In_665);
nand U26 (N_26,In_656,In_547);
nand U27 (N_27,In_557,In_365);
nor U28 (N_28,In_240,In_605);
nand U29 (N_29,In_380,In_343);
or U30 (N_30,In_421,In_216);
and U31 (N_31,In_227,In_454);
nor U32 (N_32,In_232,In_340);
xnor U33 (N_33,In_49,In_702);
or U34 (N_34,In_313,In_21);
and U35 (N_35,In_170,In_103);
or U36 (N_36,In_196,In_637);
and U37 (N_37,In_198,In_606);
and U38 (N_38,In_719,In_370);
nand U39 (N_39,In_427,In_135);
or U40 (N_40,In_229,In_213);
nor U41 (N_41,In_670,In_635);
nand U42 (N_42,In_748,In_60);
and U43 (N_43,In_397,In_77);
nor U44 (N_44,In_39,In_183);
or U45 (N_45,In_325,In_117);
and U46 (N_46,In_403,In_366);
nor U47 (N_47,In_242,In_607);
or U48 (N_48,In_206,In_243);
and U49 (N_49,In_134,In_511);
nor U50 (N_50,In_379,In_499);
nor U51 (N_51,In_331,In_125);
or U52 (N_52,In_425,In_519);
nand U53 (N_53,In_395,In_578);
or U54 (N_54,In_710,In_233);
or U55 (N_55,In_387,In_603);
and U56 (N_56,In_740,In_471);
nand U57 (N_57,In_323,In_609);
nand U58 (N_58,In_562,In_34);
xnor U59 (N_59,In_496,In_177);
nand U60 (N_60,In_338,In_66);
and U61 (N_61,In_377,In_685);
nand U62 (N_62,In_457,In_686);
and U63 (N_63,In_551,In_78);
and U64 (N_64,In_147,In_116);
nor U65 (N_65,In_80,In_261);
xnor U66 (N_66,In_472,In_598);
or U67 (N_67,In_40,In_391);
and U68 (N_68,In_559,In_661);
nor U69 (N_69,In_102,In_99);
and U70 (N_70,In_20,In_489);
or U71 (N_71,In_724,In_735);
nand U72 (N_72,In_297,In_672);
nor U73 (N_73,In_81,In_180);
and U74 (N_74,In_541,In_212);
or U75 (N_75,In_256,In_178);
and U76 (N_76,In_731,In_596);
or U77 (N_77,In_15,In_636);
and U78 (N_78,In_136,In_628);
nor U79 (N_79,In_3,In_10);
nor U80 (N_80,In_399,In_150);
nor U81 (N_81,In_422,In_384);
nor U82 (N_82,In_376,In_17);
and U83 (N_83,In_101,In_167);
nand U84 (N_84,In_417,In_357);
nand U85 (N_85,In_431,In_210);
or U86 (N_86,In_601,In_44);
and U87 (N_87,In_192,In_548);
or U88 (N_88,In_737,In_704);
nor U89 (N_89,In_528,In_515);
nor U90 (N_90,In_70,In_494);
and U91 (N_91,In_461,In_218);
or U92 (N_92,In_653,In_663);
or U93 (N_93,In_273,In_575);
or U94 (N_94,In_481,In_226);
nor U95 (N_95,In_689,In_296);
nor U96 (N_96,In_254,In_8);
xor U97 (N_97,In_367,In_314);
and U98 (N_98,In_26,In_477);
nand U99 (N_99,In_563,In_643);
nand U100 (N_100,In_361,In_219);
and U101 (N_101,In_287,In_627);
xnor U102 (N_102,In_223,In_251);
nand U103 (N_103,In_746,In_231);
or U104 (N_104,N_19,In_324);
nor U105 (N_105,N_27,In_732);
or U106 (N_106,N_52,In_209);
nand U107 (N_107,In_483,In_67);
or U108 (N_108,In_248,In_728);
nor U109 (N_109,In_317,In_75);
xnor U110 (N_110,In_584,In_388);
and U111 (N_111,In_744,In_514);
or U112 (N_112,In_626,N_6);
xor U113 (N_113,N_99,In_272);
or U114 (N_114,In_513,In_200);
nand U115 (N_115,N_11,In_692);
nor U116 (N_116,In_600,In_708);
nand U117 (N_117,In_623,In_439);
nor U118 (N_118,In_311,In_346);
nor U119 (N_119,In_159,In_139);
nand U120 (N_120,N_15,In_718);
nor U121 (N_121,In_695,N_82);
nor U122 (N_122,In_74,In_257);
and U123 (N_123,In_516,In_303);
and U124 (N_124,N_71,In_312);
and U125 (N_125,In_293,In_382);
nor U126 (N_126,In_173,In_290);
and U127 (N_127,In_260,In_646);
and U128 (N_128,N_79,N_94);
nor U129 (N_129,In_364,N_85);
and U130 (N_130,In_572,In_100);
and U131 (N_131,In_599,In_411);
nor U132 (N_132,In_249,In_749);
nor U133 (N_133,In_535,In_484);
nand U134 (N_134,In_156,In_32);
and U135 (N_135,In_502,N_16);
and U136 (N_136,In_28,N_17);
nor U137 (N_137,N_45,In_330);
nor U138 (N_138,In_383,In_687);
or U139 (N_139,In_269,N_43);
and U140 (N_140,In_539,In_703);
and U141 (N_141,N_24,In_322);
and U142 (N_142,In_487,In_564);
nor U143 (N_143,In_130,In_529);
nand U144 (N_144,In_142,In_321);
nand U145 (N_145,In_360,In_410);
and U146 (N_146,In_190,In_94);
nand U147 (N_147,In_45,In_642);
and U148 (N_148,In_280,In_726);
and U149 (N_149,N_91,N_26);
nand U150 (N_150,In_684,In_730);
and U151 (N_151,N_60,In_12);
xor U152 (N_152,In_381,In_447);
or U153 (N_153,In_118,In_154);
and U154 (N_154,In_553,In_350);
nand U155 (N_155,In_586,In_239);
or U156 (N_156,In_328,In_583);
nor U157 (N_157,In_705,In_406);
nand U158 (N_158,In_292,In_463);
nor U159 (N_159,In_301,In_259);
nor U160 (N_160,In_650,In_124);
nand U161 (N_161,In_358,In_452);
nor U162 (N_162,In_540,N_1);
or U163 (N_163,In_385,N_98);
and U164 (N_164,In_23,In_660);
or U165 (N_165,In_476,In_244);
nand U166 (N_166,In_720,In_413);
and U167 (N_167,In_195,In_404);
nor U168 (N_168,In_674,N_48);
or U169 (N_169,In_374,In_71);
or U170 (N_170,In_83,N_97);
nor U171 (N_171,In_445,In_205);
nand U172 (N_172,N_75,In_733);
and U173 (N_173,In_671,In_85);
or U174 (N_174,N_7,In_144);
nand U175 (N_175,In_594,In_128);
or U176 (N_176,In_393,In_87);
and U177 (N_177,In_434,In_250);
xnor U178 (N_178,In_204,In_175);
nand U179 (N_179,In_129,In_263);
or U180 (N_180,In_176,In_500);
and U181 (N_181,In_161,In_27);
xnor U182 (N_182,In_690,In_741);
or U183 (N_183,In_1,In_420);
nor U184 (N_184,In_711,In_652);
or U185 (N_185,In_334,N_38);
nand U186 (N_186,In_394,In_675);
nor U187 (N_187,In_508,In_274);
nor U188 (N_188,In_0,In_59);
and U189 (N_189,In_181,In_490);
or U190 (N_190,In_629,In_577);
nand U191 (N_191,In_651,N_61);
xnor U192 (N_192,In_220,In_739);
or U193 (N_193,In_625,N_25);
or U194 (N_194,N_46,In_123);
and U195 (N_195,In_315,In_677);
xnor U196 (N_196,N_88,In_299);
or U197 (N_197,N_44,In_649);
and U198 (N_198,N_72,N_41);
or U199 (N_199,In_47,In_571);
nand U200 (N_200,In_437,N_190);
xor U201 (N_201,In_18,In_469);
and U202 (N_202,In_194,In_172);
nand U203 (N_203,In_407,In_478);
nand U204 (N_204,In_532,N_92);
nor U205 (N_205,N_77,N_57);
xor U206 (N_206,N_134,In_716);
nand U207 (N_207,N_117,In_444);
nand U208 (N_208,In_199,N_114);
or U209 (N_209,In_713,N_127);
or U210 (N_210,In_57,N_74);
nor U211 (N_211,N_169,In_168);
or U212 (N_212,N_175,In_441);
nor U213 (N_213,In_275,In_72);
nand U214 (N_214,In_148,N_23);
nor U215 (N_215,N_102,In_561);
nand U216 (N_216,N_161,N_108);
and U217 (N_217,In_111,In_262);
and U218 (N_218,In_602,In_581);
xor U219 (N_219,N_76,In_63);
or U220 (N_220,In_641,In_166);
xnor U221 (N_221,In_568,N_145);
or U222 (N_222,In_402,In_574);
xnor U223 (N_223,In_179,N_18);
and U224 (N_224,N_62,In_668);
and U225 (N_225,In_106,In_222);
nor U226 (N_226,In_294,In_33);
xnor U227 (N_227,In_622,In_6);
or U228 (N_228,In_658,N_35);
nor U229 (N_229,In_22,N_138);
and U230 (N_230,In_187,In_433);
or U231 (N_231,In_46,In_424);
xor U232 (N_232,In_482,In_537);
and U233 (N_233,In_50,In_302);
and U234 (N_234,In_369,In_246);
xor U235 (N_235,In_140,In_579);
nand U236 (N_236,In_373,In_612);
or U237 (N_237,In_38,N_105);
xor U238 (N_238,In_171,N_109);
nand U239 (N_239,In_694,In_284);
or U240 (N_240,In_98,In_197);
and U241 (N_241,In_279,In_525);
or U242 (N_242,In_419,In_504);
or U243 (N_243,N_69,In_610);
nor U244 (N_244,In_89,N_73);
or U245 (N_245,In_132,In_267);
and U246 (N_246,In_65,N_118);
or U247 (N_247,N_187,N_191);
or U248 (N_248,In_722,N_144);
nor U249 (N_249,N_120,In_336);
or U250 (N_250,In_310,N_39);
and U251 (N_251,N_193,In_632);
or U252 (N_252,In_247,N_199);
nand U253 (N_253,In_105,In_621);
and U254 (N_254,N_133,N_0);
nor U255 (N_255,In_108,In_122);
and U256 (N_256,In_618,N_55);
and U257 (N_257,N_198,N_173);
nor U258 (N_258,In_283,In_688);
nand U259 (N_259,In_682,In_186);
and U260 (N_260,In_208,In_435);
or U261 (N_261,In_698,N_122);
or U262 (N_262,In_468,In_432);
xnor U263 (N_263,In_604,In_597);
nand U264 (N_264,In_405,N_21);
and U265 (N_265,N_140,In_556);
or U266 (N_266,N_112,N_93);
nand U267 (N_267,N_22,In_669);
nor U268 (N_268,In_592,In_318);
nor U269 (N_269,N_164,In_582);
xnor U270 (N_270,In_491,In_97);
nor U271 (N_271,N_152,In_423);
xnor U272 (N_272,N_137,N_166);
nand U273 (N_273,In_201,N_151);
xnor U274 (N_274,N_146,In_520);
or U275 (N_275,N_142,In_127);
and U276 (N_276,In_16,In_149);
nand U277 (N_277,In_631,In_230);
nor U278 (N_278,N_186,In_305);
or U279 (N_279,In_113,N_148);
nor U280 (N_280,N_197,In_245);
or U281 (N_281,In_4,In_506);
nand U282 (N_282,In_332,In_30);
nand U283 (N_283,N_188,N_156);
nand U284 (N_284,In_193,N_49);
nand U285 (N_285,In_640,In_400);
nor U286 (N_286,In_86,N_47);
nor U287 (N_287,In_495,N_54);
xor U288 (N_288,In_137,In_480);
nor U289 (N_289,N_2,N_184);
or U290 (N_290,N_100,In_174);
xor U291 (N_291,In_188,In_339);
or U292 (N_292,In_608,In_415);
and U293 (N_293,N_20,In_617);
xnor U294 (N_294,In_466,In_585);
nor U295 (N_295,In_473,In_428);
nor U296 (N_296,In_459,N_14);
nand U297 (N_297,N_119,In_51);
or U298 (N_298,In_566,In_589);
and U299 (N_299,N_107,In_408);
and U300 (N_300,In_191,In_104);
or U301 (N_301,N_128,In_182);
nand U302 (N_302,In_35,In_386);
nor U303 (N_303,N_10,N_64);
nand U304 (N_304,N_8,In_276);
nor U305 (N_305,N_113,N_106);
nor U306 (N_306,In_510,In_228);
nand U307 (N_307,In_550,N_65);
or U308 (N_308,In_54,In_691);
and U309 (N_309,N_215,In_265);
and U310 (N_310,In_56,N_250);
nand U311 (N_311,N_121,In_157);
nor U312 (N_312,In_523,N_204);
and U313 (N_313,In_110,In_630);
nor U314 (N_314,N_202,In_309);
and U315 (N_315,N_183,N_125);
and U316 (N_316,N_78,N_165);
or U317 (N_317,N_168,In_440);
nand U318 (N_318,N_89,In_271);
nor U319 (N_319,In_236,In_153);
and U320 (N_320,In_163,In_569);
and U321 (N_321,N_154,N_241);
or U322 (N_322,N_153,N_271);
nor U323 (N_323,N_70,In_349);
nand U324 (N_324,In_326,In_112);
xor U325 (N_325,N_143,In_368);
and U326 (N_326,N_68,In_9);
nor U327 (N_327,N_298,N_272);
and U328 (N_328,N_253,In_253);
nor U329 (N_329,N_287,In_234);
or U330 (N_330,In_185,N_257);
and U331 (N_331,N_32,N_292);
nand U332 (N_332,In_345,In_717);
nor U333 (N_333,N_248,N_249);
and U334 (N_334,In_462,In_449);
and U335 (N_335,In_25,In_533);
xnor U336 (N_336,In_79,N_232);
nand U337 (N_337,In_662,In_11);
or U338 (N_338,In_371,In_436);
and U339 (N_339,In_37,In_680);
xor U340 (N_340,In_450,N_42);
nor U341 (N_341,In_614,N_149);
nor U342 (N_342,N_295,In_667);
nand U343 (N_343,N_104,N_63);
nand U344 (N_344,In_488,In_362);
nand U345 (N_345,N_34,N_226);
nor U346 (N_346,In_501,In_518);
or U347 (N_347,N_158,In_96);
xor U348 (N_348,N_224,N_284);
nor U349 (N_349,In_645,N_33);
and U350 (N_350,N_227,In_29);
nand U351 (N_351,In_426,In_320);
xnor U352 (N_352,In_88,N_254);
nor U353 (N_353,N_116,In_288);
nor U354 (N_354,In_467,N_277);
nand U355 (N_355,In_289,N_195);
nand U356 (N_356,In_36,N_245);
and U357 (N_357,N_200,N_218);
nand U358 (N_358,N_259,N_196);
nand U359 (N_359,In_92,N_150);
or U360 (N_360,N_251,In_453);
nand U361 (N_361,In_474,In_638);
and U362 (N_362,In_295,N_29);
nand U363 (N_363,In_414,In_576);
nor U364 (N_364,In_155,N_234);
and U365 (N_365,N_192,In_55);
and U366 (N_366,In_352,N_273);
and U367 (N_367,In_126,N_194);
or U368 (N_368,N_110,In_258);
nand U369 (N_369,In_152,In_475);
or U370 (N_370,In_354,N_243);
or U371 (N_371,N_160,In_19);
nor U372 (N_372,N_5,In_389);
or U373 (N_373,N_285,N_67);
and U374 (N_374,N_274,N_291);
nand U375 (N_375,In_316,N_56);
nand U376 (N_376,In_536,N_86);
xnor U377 (N_377,In_464,N_278);
or U378 (N_378,In_31,In_68);
nor U379 (N_379,N_237,In_165);
or U380 (N_380,In_412,N_31);
xor U381 (N_381,In_438,N_66);
and U382 (N_382,N_176,In_567);
or U383 (N_383,In_329,N_281);
nor U384 (N_384,In_286,N_294);
nor U385 (N_385,N_282,N_201);
or U386 (N_386,N_135,In_742);
nand U387 (N_387,N_130,In_455);
and U388 (N_388,N_269,N_189);
and U389 (N_389,In_616,In_43);
and U390 (N_390,In_372,In_418);
xor U391 (N_391,N_174,N_289);
xor U392 (N_392,In_138,In_356);
or U393 (N_393,N_267,In_69);
or U394 (N_394,In_264,N_141);
xnor U395 (N_395,In_207,N_225);
nand U396 (N_396,In_456,N_238);
and U397 (N_397,In_696,In_545);
and U398 (N_398,N_203,In_278);
and U399 (N_399,N_9,N_283);
nand U400 (N_400,N_235,N_335);
or U401 (N_401,N_136,N_332);
or U402 (N_402,In_611,N_129);
nand U403 (N_403,N_181,N_312);
and U404 (N_404,In_347,In_306);
xnor U405 (N_405,In_727,N_209);
nand U406 (N_406,N_301,N_179);
and U407 (N_407,In_429,N_28);
xnor U408 (N_408,N_275,In_723);
and U409 (N_409,In_699,In_238);
or U410 (N_410,In_5,In_648);
xnor U411 (N_411,N_384,N_244);
nor U412 (N_412,N_276,In_91);
or U413 (N_413,N_255,N_307);
and U414 (N_414,In_706,N_381);
or U415 (N_415,N_162,N_385);
or U416 (N_416,In_162,N_124);
xor U417 (N_417,In_497,N_352);
or U418 (N_418,In_390,N_131);
and U419 (N_419,N_354,N_366);
or U420 (N_420,N_84,N_319);
or U421 (N_421,N_239,N_383);
or U422 (N_422,N_330,In_712);
nor U423 (N_423,N_233,N_300);
and U424 (N_424,In_396,In_587);
nand U425 (N_425,N_362,In_521);
or U426 (N_426,N_229,In_308);
nor U427 (N_427,N_348,N_50);
xnor U428 (N_428,N_375,N_103);
nand U429 (N_429,In_378,In_225);
and U430 (N_430,N_167,N_213);
or U431 (N_431,N_388,N_182);
and U432 (N_432,In_486,N_262);
nand U433 (N_433,In_679,N_95);
xor U434 (N_434,N_216,N_115);
nor U435 (N_435,In_543,In_681);
nand U436 (N_436,In_570,In_351);
and U437 (N_437,N_208,N_96);
or U438 (N_438,N_367,In_593);
or U439 (N_439,N_353,N_37);
nand U440 (N_440,N_221,N_155);
nand U441 (N_441,In_534,N_374);
nand U442 (N_442,N_318,N_80);
xor U443 (N_443,N_172,In_659);
nand U444 (N_444,In_634,In_342);
and U445 (N_445,N_240,N_322);
nor U446 (N_446,In_115,N_53);
nand U447 (N_447,N_347,In_184);
and U448 (N_448,In_701,N_314);
nor U449 (N_449,In_524,In_743);
xor U450 (N_450,In_84,In_375);
nor U451 (N_451,N_258,In_573);
nor U452 (N_452,N_217,N_310);
nand U453 (N_453,In_644,N_256);
or U454 (N_454,In_666,N_365);
nor U455 (N_455,N_247,In_591);
or U456 (N_456,In_285,N_293);
xnor U457 (N_457,N_51,In_613);
xor U458 (N_458,N_13,In_2);
nand U459 (N_459,In_619,In_109);
nor U460 (N_460,In_633,N_313);
nand U461 (N_461,In_24,In_560);
nand U462 (N_462,In_451,N_337);
and U463 (N_463,In_41,In_715);
nor U464 (N_464,N_356,In_736);
and U465 (N_465,N_302,N_346);
xor U466 (N_466,N_210,N_333);
or U467 (N_467,N_359,In_657);
nand U468 (N_468,N_123,N_205);
nor U469 (N_469,In_141,N_392);
nor U470 (N_470,In_189,In_214);
and U471 (N_471,N_290,N_327);
nand U472 (N_472,In_266,N_320);
nor U473 (N_473,N_369,N_361);
nand U474 (N_474,N_379,N_296);
nand U475 (N_475,In_203,In_493);
xnor U476 (N_476,In_615,N_126);
and U477 (N_477,In_552,N_315);
or U478 (N_478,In_588,In_530);
xnor U479 (N_479,In_544,In_745);
and U480 (N_480,N_338,In_131);
nand U481 (N_481,N_323,N_393);
nor U482 (N_482,N_36,N_230);
and U483 (N_483,N_372,In_401);
nand U484 (N_484,N_58,In_538);
and U485 (N_485,N_339,N_180);
xnor U486 (N_486,N_101,In_120);
or U487 (N_487,N_340,N_334);
nor U488 (N_488,N_139,N_268);
and U489 (N_489,N_211,In_707);
xnor U490 (N_490,N_336,N_59);
and U491 (N_491,In_398,In_697);
nand U492 (N_492,N_345,N_261);
and U493 (N_493,N_394,N_342);
and U494 (N_494,N_363,N_328);
nor U495 (N_495,N_380,In_639);
nand U496 (N_496,In_344,In_282);
and U497 (N_497,N_266,N_4);
nor U498 (N_498,N_325,N_304);
nor U499 (N_499,In_270,In_158);
nor U500 (N_500,N_371,N_461);
and U501 (N_501,N_483,N_428);
or U502 (N_502,In_224,N_491);
and U503 (N_503,N_324,N_485);
or U504 (N_504,N_264,In_747);
or U505 (N_505,In_151,N_411);
or U506 (N_506,N_458,N_457);
nor U507 (N_507,N_481,N_418);
and U508 (N_508,N_157,N_430);
or U509 (N_509,N_403,N_265);
nor U510 (N_510,N_344,In_512);
nor U511 (N_511,N_443,In_237);
nor U512 (N_512,In_517,N_220);
nand U513 (N_513,N_389,N_357);
and U514 (N_514,In_42,N_465);
or U515 (N_515,N_406,In_64);
and U516 (N_516,N_454,N_462);
nor U517 (N_517,N_398,N_490);
and U518 (N_518,In_93,N_469);
or U519 (N_519,In_416,In_333);
xor U520 (N_520,N_441,N_421);
nor U521 (N_521,N_228,N_309);
nand U522 (N_522,N_178,In_348);
or U523 (N_523,N_431,In_509);
and U524 (N_524,N_409,N_223);
nor U525 (N_525,N_299,N_410);
nor U526 (N_526,N_397,In_95);
and U527 (N_527,N_350,N_378);
and U528 (N_528,N_207,In_82);
nand U529 (N_529,In_281,In_479);
xnor U530 (N_530,N_246,In_335);
xnor U531 (N_531,N_396,N_426);
nand U532 (N_532,N_445,N_434);
nor U533 (N_533,N_163,N_185);
and U534 (N_534,In_76,N_317);
nor U535 (N_535,N_231,In_121);
nor U536 (N_536,N_30,N_370);
and U537 (N_537,In_53,In_300);
nand U538 (N_538,N_437,In_485);
nand U539 (N_539,N_479,N_422);
or U540 (N_540,N_467,In_526);
nand U541 (N_541,N_478,N_413);
or U542 (N_542,In_678,In_503);
nand U543 (N_543,N_159,N_387);
or U544 (N_544,N_405,N_450);
or U545 (N_545,In_133,N_242);
or U546 (N_546,N_331,N_316);
and U547 (N_547,N_382,In_143);
and U548 (N_548,N_476,N_463);
nand U549 (N_549,In_549,N_494);
and U550 (N_550,N_453,N_386);
nor U551 (N_551,N_425,N_308);
nand U552 (N_552,N_390,N_83);
nor U553 (N_553,N_466,N_306);
nand U554 (N_554,In_595,In_298);
and U555 (N_555,N_305,In_235);
and U556 (N_556,N_477,In_693);
or U557 (N_557,In_654,N_493);
nor U558 (N_558,N_402,N_401);
or U559 (N_559,N_489,N_455);
or U560 (N_560,In_241,In_676);
xnor U561 (N_561,N_448,N_472);
xor U562 (N_562,N_373,N_496);
nor U563 (N_563,N_288,N_447);
or U564 (N_564,N_495,In_61);
and U565 (N_565,N_464,N_341);
or U566 (N_566,N_260,N_360);
nor U567 (N_567,N_326,N_475);
xnor U568 (N_568,N_355,N_470);
nand U569 (N_569,In_252,N_270);
and U570 (N_570,N_90,N_480);
and U571 (N_571,In_7,N_415);
and U572 (N_572,In_443,N_280);
or U573 (N_573,N_81,N_456);
nor U574 (N_574,N_399,In_527);
nand U575 (N_575,N_206,N_351);
xnor U576 (N_576,N_343,N_404);
or U577 (N_577,N_460,N_311);
nor U578 (N_578,N_432,N_297);
nand U579 (N_579,N_433,In_291);
and U580 (N_580,N_487,N_358);
or U581 (N_581,N_446,N_279);
nor U582 (N_582,N_468,N_321);
or U583 (N_583,N_364,N_349);
xnor U584 (N_584,N_214,N_132);
and U585 (N_585,N_40,In_58);
or U586 (N_586,N_212,N_424);
and U587 (N_587,N_252,N_170);
and U588 (N_588,N_429,N_482);
and U589 (N_589,N_499,N_459);
and U590 (N_590,N_408,N_376);
nand U591 (N_591,N_451,N_147);
nor U592 (N_592,N_497,N_414);
xnor U593 (N_593,N_87,N_486);
nand U594 (N_594,N_452,In_355);
nand U595 (N_595,N_263,In_145);
or U596 (N_596,N_377,N_303);
nand U597 (N_597,N_412,N_419);
and U598 (N_598,In_392,N_400);
and U599 (N_599,In_341,In_673);
or U600 (N_600,In_498,N_563);
and U601 (N_601,N_420,N_427);
nor U602 (N_602,N_599,N_524);
or U603 (N_603,N_473,N_546);
nand U604 (N_604,N_592,N_587);
or U605 (N_605,N_549,N_545);
nor U606 (N_606,N_575,In_221);
nand U607 (N_607,N_548,N_525);
nand U608 (N_608,In_215,N_579);
nor U609 (N_609,N_568,N_286);
xor U610 (N_610,N_597,N_554);
nand U611 (N_611,N_559,N_488);
and U612 (N_612,N_567,N_566);
and U613 (N_613,N_530,N_177);
xor U614 (N_614,N_581,N_506);
or U615 (N_615,N_236,N_442);
nor U616 (N_616,N_553,N_560);
or U617 (N_617,In_217,N_542);
or U618 (N_618,N_593,In_304);
nand U619 (N_619,N_521,N_502);
and U620 (N_620,N_557,N_595);
nand U621 (N_621,N_529,N_532);
or U622 (N_622,N_551,N_501);
and U623 (N_623,N_12,N_531);
and U624 (N_624,N_583,N_518);
and U625 (N_625,N_515,N_391);
and U626 (N_626,N_570,In_73);
xnor U627 (N_627,N_584,In_505);
or U628 (N_628,N_543,N_588);
and U629 (N_629,N_511,N_423);
or U630 (N_630,N_541,N_517);
nand U631 (N_631,N_561,In_327);
xor U632 (N_632,N_503,N_565);
nand U633 (N_633,N_520,In_442);
or U634 (N_634,N_471,N_513);
or U635 (N_635,N_440,N_578);
nand U636 (N_636,N_585,N_574);
xor U637 (N_637,N_596,N_572);
nand U638 (N_638,N_474,N_582);
and U639 (N_639,N_171,N_500);
nand U640 (N_640,N_510,N_484);
nor U641 (N_641,N_519,N_562);
nor U642 (N_642,N_368,N_407);
or U643 (N_643,N_556,In_62);
or U644 (N_644,N_598,N_555);
or U645 (N_645,N_537,N_527);
xnor U646 (N_646,N_558,N_550);
or U647 (N_647,N_571,N_594);
and U648 (N_648,N_535,N_492);
and U649 (N_649,N_577,N_444);
xnor U650 (N_650,N_534,N_522);
or U651 (N_651,N_449,N_508);
or U652 (N_652,N_222,N_591);
nor U653 (N_653,N_509,N_538);
nand U654 (N_654,N_569,N_528);
xnor U655 (N_655,N_580,N_539);
nor U656 (N_656,N_564,N_435);
or U657 (N_657,In_169,N_552);
nand U658 (N_658,In_119,N_507);
xor U659 (N_659,N_526,N_219);
or U660 (N_660,N_533,N_540);
or U661 (N_661,N_514,N_416);
xor U662 (N_662,N_523,In_558);
and U663 (N_663,N_504,N_417);
xor U664 (N_664,N_536,N_547);
nor U665 (N_665,N_586,N_590);
and U666 (N_666,N_516,N_573);
nor U667 (N_667,N_498,N_329);
and U668 (N_668,In_542,N_505);
and U669 (N_669,In_337,N_544);
nand U670 (N_670,N_512,N_436);
and U671 (N_671,N_439,N_589);
nand U672 (N_672,N_576,N_438);
and U673 (N_673,N_3,N_395);
and U674 (N_674,In_363,N_111);
or U675 (N_675,N_440,N_595);
and U676 (N_676,N_588,N_556);
nor U677 (N_677,In_73,In_119);
and U678 (N_678,N_518,N_570);
nand U679 (N_679,N_519,N_420);
nand U680 (N_680,N_572,N_12);
nand U681 (N_681,N_513,N_395);
and U682 (N_682,N_535,N_588);
nand U683 (N_683,N_511,N_527);
nor U684 (N_684,N_583,N_407);
and U685 (N_685,N_571,N_560);
or U686 (N_686,N_575,N_534);
xnor U687 (N_687,N_473,N_548);
xor U688 (N_688,N_3,N_529);
nand U689 (N_689,N_510,N_556);
and U690 (N_690,N_416,N_492);
and U691 (N_691,N_534,N_514);
or U692 (N_692,N_435,N_498);
or U693 (N_693,N_581,N_515);
and U694 (N_694,N_560,N_577);
or U695 (N_695,N_506,N_552);
and U696 (N_696,N_580,N_588);
and U697 (N_697,N_520,In_327);
or U698 (N_698,N_554,N_524);
xnor U699 (N_699,N_420,N_395);
xnor U700 (N_700,N_693,N_646);
nor U701 (N_701,N_685,N_650);
nand U702 (N_702,N_670,N_689);
nor U703 (N_703,N_618,N_686);
or U704 (N_704,N_633,N_663);
nor U705 (N_705,N_688,N_661);
nor U706 (N_706,N_662,N_674);
or U707 (N_707,N_698,N_660);
or U708 (N_708,N_697,N_630);
or U709 (N_709,N_625,N_647);
or U710 (N_710,N_657,N_610);
xnor U711 (N_711,N_695,N_669);
and U712 (N_712,N_692,N_629);
nand U713 (N_713,N_683,N_602);
or U714 (N_714,N_643,N_601);
and U715 (N_715,N_619,N_664);
or U716 (N_716,N_631,N_611);
nand U717 (N_717,N_627,N_684);
or U718 (N_718,N_673,N_644);
and U719 (N_719,N_656,N_606);
nor U720 (N_720,N_626,N_636);
and U721 (N_721,N_600,N_666);
nand U722 (N_722,N_604,N_690);
xor U723 (N_723,N_675,N_648);
or U724 (N_724,N_655,N_605);
nor U725 (N_725,N_612,N_617);
or U726 (N_726,N_696,N_637);
xnor U727 (N_727,N_624,N_681);
or U728 (N_728,N_623,N_622);
nor U729 (N_729,N_668,N_645);
nand U730 (N_730,N_680,N_608);
nand U731 (N_731,N_658,N_638);
nor U732 (N_732,N_621,N_607);
and U733 (N_733,N_671,N_652);
or U734 (N_734,N_659,N_613);
nand U735 (N_735,N_641,N_609);
nor U736 (N_736,N_614,N_654);
and U737 (N_737,N_667,N_628);
or U738 (N_738,N_634,N_653);
or U739 (N_739,N_651,N_665);
or U740 (N_740,N_603,N_642);
nor U741 (N_741,N_682,N_677);
and U742 (N_742,N_635,N_639);
xor U743 (N_743,N_676,N_694);
and U744 (N_744,N_640,N_679);
nor U745 (N_745,N_649,N_678);
nor U746 (N_746,N_672,N_616);
or U747 (N_747,N_632,N_691);
xnor U748 (N_748,N_615,N_699);
or U749 (N_749,N_687,N_620);
and U750 (N_750,N_624,N_618);
nor U751 (N_751,N_601,N_647);
and U752 (N_752,N_619,N_696);
nor U753 (N_753,N_606,N_649);
and U754 (N_754,N_611,N_668);
nand U755 (N_755,N_695,N_665);
xnor U756 (N_756,N_653,N_676);
or U757 (N_757,N_603,N_688);
and U758 (N_758,N_661,N_663);
nand U759 (N_759,N_666,N_634);
and U760 (N_760,N_608,N_614);
nand U761 (N_761,N_690,N_692);
nand U762 (N_762,N_682,N_608);
nor U763 (N_763,N_681,N_679);
nand U764 (N_764,N_649,N_638);
nand U765 (N_765,N_670,N_676);
nand U766 (N_766,N_654,N_657);
nor U767 (N_767,N_614,N_616);
or U768 (N_768,N_685,N_684);
and U769 (N_769,N_636,N_662);
and U770 (N_770,N_674,N_648);
nor U771 (N_771,N_636,N_652);
nand U772 (N_772,N_639,N_612);
or U773 (N_773,N_619,N_620);
or U774 (N_774,N_692,N_654);
nor U775 (N_775,N_693,N_688);
or U776 (N_776,N_654,N_610);
nand U777 (N_777,N_646,N_613);
nor U778 (N_778,N_625,N_652);
or U779 (N_779,N_627,N_670);
and U780 (N_780,N_692,N_651);
and U781 (N_781,N_669,N_617);
nor U782 (N_782,N_611,N_637);
or U783 (N_783,N_639,N_669);
or U784 (N_784,N_695,N_699);
and U785 (N_785,N_623,N_629);
and U786 (N_786,N_609,N_639);
or U787 (N_787,N_625,N_698);
nand U788 (N_788,N_617,N_633);
nand U789 (N_789,N_673,N_613);
nor U790 (N_790,N_665,N_652);
nor U791 (N_791,N_665,N_630);
or U792 (N_792,N_621,N_633);
or U793 (N_793,N_602,N_609);
nand U794 (N_794,N_605,N_676);
xor U795 (N_795,N_602,N_619);
nor U796 (N_796,N_662,N_675);
or U797 (N_797,N_663,N_697);
nand U798 (N_798,N_684,N_639);
nor U799 (N_799,N_623,N_632);
or U800 (N_800,N_770,N_745);
nand U801 (N_801,N_796,N_712);
xor U802 (N_802,N_797,N_764);
nor U803 (N_803,N_715,N_730);
and U804 (N_804,N_771,N_760);
and U805 (N_805,N_772,N_753);
and U806 (N_806,N_720,N_719);
nand U807 (N_807,N_755,N_711);
and U808 (N_808,N_731,N_710);
and U809 (N_809,N_733,N_776);
and U810 (N_810,N_736,N_757);
nand U811 (N_811,N_748,N_729);
nand U812 (N_812,N_700,N_721);
and U813 (N_813,N_762,N_774);
or U814 (N_814,N_703,N_756);
nand U815 (N_815,N_784,N_775);
and U816 (N_816,N_769,N_763);
nor U817 (N_817,N_702,N_754);
nor U818 (N_818,N_778,N_785);
and U819 (N_819,N_705,N_701);
and U820 (N_820,N_709,N_722);
and U821 (N_821,N_761,N_751);
and U822 (N_822,N_718,N_707);
nor U823 (N_823,N_746,N_791);
or U824 (N_824,N_750,N_765);
nand U825 (N_825,N_792,N_723);
or U826 (N_826,N_766,N_758);
or U827 (N_827,N_768,N_744);
or U828 (N_828,N_706,N_734);
xor U829 (N_829,N_790,N_795);
or U830 (N_830,N_704,N_725);
xor U831 (N_831,N_783,N_743);
nand U832 (N_832,N_798,N_782);
xnor U833 (N_833,N_786,N_794);
nor U834 (N_834,N_727,N_713);
nor U835 (N_835,N_728,N_793);
or U836 (N_836,N_716,N_773);
nor U837 (N_837,N_777,N_781);
nand U838 (N_838,N_740,N_767);
and U839 (N_839,N_788,N_732);
nor U840 (N_840,N_714,N_708);
nand U841 (N_841,N_789,N_735);
nor U842 (N_842,N_717,N_747);
and U843 (N_843,N_787,N_726);
and U844 (N_844,N_741,N_737);
and U845 (N_845,N_738,N_752);
nor U846 (N_846,N_799,N_759);
nor U847 (N_847,N_739,N_780);
or U848 (N_848,N_779,N_742);
or U849 (N_849,N_724,N_749);
xnor U850 (N_850,N_777,N_798);
or U851 (N_851,N_778,N_721);
nor U852 (N_852,N_799,N_746);
or U853 (N_853,N_788,N_761);
nor U854 (N_854,N_754,N_704);
and U855 (N_855,N_767,N_771);
nor U856 (N_856,N_736,N_744);
and U857 (N_857,N_775,N_750);
and U858 (N_858,N_791,N_745);
or U859 (N_859,N_755,N_745);
and U860 (N_860,N_713,N_780);
nor U861 (N_861,N_759,N_727);
nor U862 (N_862,N_701,N_769);
xnor U863 (N_863,N_788,N_736);
xor U864 (N_864,N_717,N_781);
and U865 (N_865,N_741,N_721);
xor U866 (N_866,N_715,N_799);
or U867 (N_867,N_739,N_716);
or U868 (N_868,N_784,N_778);
and U869 (N_869,N_710,N_718);
and U870 (N_870,N_733,N_734);
and U871 (N_871,N_760,N_717);
nand U872 (N_872,N_783,N_753);
or U873 (N_873,N_717,N_722);
nor U874 (N_874,N_738,N_796);
and U875 (N_875,N_714,N_778);
or U876 (N_876,N_785,N_736);
or U877 (N_877,N_747,N_753);
and U878 (N_878,N_773,N_740);
nor U879 (N_879,N_752,N_733);
nor U880 (N_880,N_744,N_702);
nand U881 (N_881,N_763,N_718);
and U882 (N_882,N_749,N_748);
or U883 (N_883,N_702,N_755);
nand U884 (N_884,N_714,N_785);
nor U885 (N_885,N_753,N_765);
and U886 (N_886,N_746,N_764);
xor U887 (N_887,N_725,N_719);
nand U888 (N_888,N_764,N_727);
nor U889 (N_889,N_729,N_762);
or U890 (N_890,N_734,N_759);
nand U891 (N_891,N_773,N_784);
nor U892 (N_892,N_723,N_761);
nor U893 (N_893,N_727,N_709);
or U894 (N_894,N_714,N_706);
and U895 (N_895,N_787,N_751);
xor U896 (N_896,N_729,N_704);
or U897 (N_897,N_797,N_751);
or U898 (N_898,N_721,N_716);
xor U899 (N_899,N_798,N_746);
nand U900 (N_900,N_857,N_838);
and U901 (N_901,N_884,N_872);
and U902 (N_902,N_822,N_865);
or U903 (N_903,N_862,N_811);
nor U904 (N_904,N_889,N_844);
xnor U905 (N_905,N_834,N_882);
and U906 (N_906,N_875,N_810);
nand U907 (N_907,N_895,N_897);
and U908 (N_908,N_877,N_878);
nand U909 (N_909,N_829,N_896);
and U910 (N_910,N_867,N_831);
nand U911 (N_911,N_858,N_814);
nor U912 (N_912,N_854,N_869);
or U913 (N_913,N_821,N_894);
nor U914 (N_914,N_851,N_813);
or U915 (N_915,N_886,N_828);
xor U916 (N_916,N_839,N_888);
nand U917 (N_917,N_866,N_879);
nor U918 (N_918,N_803,N_876);
nor U919 (N_919,N_891,N_804);
xor U920 (N_920,N_848,N_824);
and U921 (N_921,N_812,N_893);
nor U922 (N_922,N_883,N_818);
nor U923 (N_923,N_849,N_807);
or U924 (N_924,N_805,N_840);
nand U925 (N_925,N_808,N_827);
or U926 (N_926,N_890,N_853);
or U927 (N_927,N_837,N_800);
nor U928 (N_928,N_850,N_820);
or U929 (N_929,N_892,N_899);
and U930 (N_930,N_868,N_815);
nand U931 (N_931,N_863,N_873);
xor U932 (N_932,N_806,N_819);
or U933 (N_933,N_836,N_898);
nor U934 (N_934,N_885,N_842);
nand U935 (N_935,N_856,N_847);
or U936 (N_936,N_843,N_835);
nand U937 (N_937,N_833,N_861);
nand U938 (N_938,N_859,N_825);
xor U939 (N_939,N_826,N_845);
nor U940 (N_940,N_855,N_841);
nand U941 (N_941,N_832,N_860);
nand U942 (N_942,N_802,N_874);
or U943 (N_943,N_801,N_881);
xnor U944 (N_944,N_809,N_830);
nand U945 (N_945,N_846,N_852);
nor U946 (N_946,N_823,N_887);
nor U947 (N_947,N_870,N_817);
and U948 (N_948,N_871,N_864);
nor U949 (N_949,N_880,N_816);
nand U950 (N_950,N_883,N_834);
nor U951 (N_951,N_821,N_826);
and U952 (N_952,N_805,N_886);
or U953 (N_953,N_893,N_824);
xnor U954 (N_954,N_807,N_806);
nor U955 (N_955,N_851,N_814);
and U956 (N_956,N_874,N_873);
or U957 (N_957,N_866,N_819);
and U958 (N_958,N_850,N_810);
nor U959 (N_959,N_881,N_809);
and U960 (N_960,N_887,N_821);
or U961 (N_961,N_877,N_863);
and U962 (N_962,N_815,N_871);
nor U963 (N_963,N_870,N_846);
or U964 (N_964,N_823,N_849);
xnor U965 (N_965,N_862,N_895);
or U966 (N_966,N_824,N_801);
xnor U967 (N_967,N_825,N_835);
and U968 (N_968,N_853,N_845);
or U969 (N_969,N_839,N_820);
nand U970 (N_970,N_859,N_801);
and U971 (N_971,N_823,N_859);
and U972 (N_972,N_833,N_885);
or U973 (N_973,N_820,N_844);
xnor U974 (N_974,N_860,N_802);
or U975 (N_975,N_825,N_807);
or U976 (N_976,N_867,N_878);
and U977 (N_977,N_801,N_818);
nand U978 (N_978,N_867,N_896);
and U979 (N_979,N_889,N_836);
nand U980 (N_980,N_841,N_829);
nor U981 (N_981,N_854,N_808);
and U982 (N_982,N_883,N_809);
nand U983 (N_983,N_832,N_827);
or U984 (N_984,N_877,N_872);
nor U985 (N_985,N_844,N_893);
nand U986 (N_986,N_860,N_868);
and U987 (N_987,N_816,N_891);
nor U988 (N_988,N_814,N_832);
nor U989 (N_989,N_864,N_845);
nor U990 (N_990,N_884,N_849);
nand U991 (N_991,N_861,N_835);
or U992 (N_992,N_802,N_867);
nand U993 (N_993,N_834,N_879);
and U994 (N_994,N_895,N_881);
nand U995 (N_995,N_823,N_818);
and U996 (N_996,N_800,N_839);
nor U997 (N_997,N_896,N_894);
or U998 (N_998,N_844,N_873);
or U999 (N_999,N_806,N_850);
or U1000 (N_1000,N_958,N_975);
and U1001 (N_1001,N_929,N_942);
or U1002 (N_1002,N_920,N_985);
and U1003 (N_1003,N_907,N_973);
nor U1004 (N_1004,N_943,N_955);
nand U1005 (N_1005,N_970,N_917);
and U1006 (N_1006,N_911,N_949);
nand U1007 (N_1007,N_914,N_948);
and U1008 (N_1008,N_998,N_924);
or U1009 (N_1009,N_902,N_953);
or U1010 (N_1010,N_964,N_984);
nand U1011 (N_1011,N_963,N_956);
nor U1012 (N_1012,N_972,N_976);
or U1013 (N_1013,N_989,N_968);
and U1014 (N_1014,N_981,N_990);
xor U1015 (N_1015,N_918,N_926);
or U1016 (N_1016,N_901,N_994);
or U1017 (N_1017,N_909,N_978);
nor U1018 (N_1018,N_905,N_969);
nor U1019 (N_1019,N_939,N_959);
nand U1020 (N_1020,N_925,N_977);
or U1021 (N_1021,N_946,N_903);
nor U1022 (N_1022,N_999,N_950);
nand U1023 (N_1023,N_921,N_988);
nor U1024 (N_1024,N_997,N_993);
or U1025 (N_1025,N_991,N_935);
or U1026 (N_1026,N_995,N_915);
and U1027 (N_1027,N_936,N_906);
or U1028 (N_1028,N_933,N_940);
nand U1029 (N_1029,N_938,N_913);
nor U1030 (N_1030,N_982,N_922);
nor U1031 (N_1031,N_937,N_954);
nand U1032 (N_1032,N_992,N_931);
xnor U1033 (N_1033,N_951,N_934);
and U1034 (N_1034,N_961,N_916);
or U1035 (N_1035,N_944,N_912);
xnor U1036 (N_1036,N_923,N_932);
nand U1037 (N_1037,N_910,N_987);
and U1038 (N_1038,N_960,N_908);
or U1039 (N_1039,N_967,N_957);
and U1040 (N_1040,N_996,N_979);
or U1041 (N_1041,N_941,N_919);
xor U1042 (N_1042,N_962,N_965);
xor U1043 (N_1043,N_900,N_928);
nand U1044 (N_1044,N_904,N_974);
and U1045 (N_1045,N_983,N_927);
xnor U1046 (N_1046,N_945,N_980);
nand U1047 (N_1047,N_952,N_986);
nor U1048 (N_1048,N_930,N_971);
or U1049 (N_1049,N_947,N_966);
nor U1050 (N_1050,N_901,N_962);
nand U1051 (N_1051,N_995,N_922);
xnor U1052 (N_1052,N_963,N_908);
xor U1053 (N_1053,N_910,N_939);
or U1054 (N_1054,N_953,N_930);
nor U1055 (N_1055,N_971,N_976);
and U1056 (N_1056,N_901,N_904);
and U1057 (N_1057,N_925,N_902);
nor U1058 (N_1058,N_957,N_945);
nor U1059 (N_1059,N_900,N_974);
nand U1060 (N_1060,N_935,N_934);
or U1061 (N_1061,N_971,N_954);
nor U1062 (N_1062,N_985,N_939);
and U1063 (N_1063,N_962,N_927);
nand U1064 (N_1064,N_901,N_951);
or U1065 (N_1065,N_974,N_966);
or U1066 (N_1066,N_948,N_922);
and U1067 (N_1067,N_919,N_956);
nand U1068 (N_1068,N_975,N_966);
nand U1069 (N_1069,N_986,N_902);
nand U1070 (N_1070,N_970,N_926);
nor U1071 (N_1071,N_983,N_988);
and U1072 (N_1072,N_933,N_908);
nand U1073 (N_1073,N_987,N_936);
nand U1074 (N_1074,N_981,N_979);
or U1075 (N_1075,N_958,N_916);
xor U1076 (N_1076,N_994,N_972);
nand U1077 (N_1077,N_954,N_945);
xor U1078 (N_1078,N_978,N_955);
and U1079 (N_1079,N_921,N_904);
nor U1080 (N_1080,N_940,N_901);
nand U1081 (N_1081,N_916,N_943);
nor U1082 (N_1082,N_911,N_989);
or U1083 (N_1083,N_973,N_956);
nand U1084 (N_1084,N_928,N_910);
and U1085 (N_1085,N_997,N_967);
or U1086 (N_1086,N_938,N_922);
or U1087 (N_1087,N_994,N_949);
and U1088 (N_1088,N_944,N_978);
or U1089 (N_1089,N_907,N_955);
nand U1090 (N_1090,N_958,N_980);
nand U1091 (N_1091,N_914,N_907);
xor U1092 (N_1092,N_949,N_962);
and U1093 (N_1093,N_901,N_902);
and U1094 (N_1094,N_982,N_920);
or U1095 (N_1095,N_952,N_974);
and U1096 (N_1096,N_946,N_963);
or U1097 (N_1097,N_977,N_967);
nand U1098 (N_1098,N_918,N_954);
nand U1099 (N_1099,N_987,N_919);
and U1100 (N_1100,N_1005,N_1031);
or U1101 (N_1101,N_1022,N_1048);
and U1102 (N_1102,N_1019,N_1066);
and U1103 (N_1103,N_1015,N_1032);
and U1104 (N_1104,N_1055,N_1082);
nand U1105 (N_1105,N_1028,N_1021);
nand U1106 (N_1106,N_1008,N_1020);
and U1107 (N_1107,N_1002,N_1069);
xor U1108 (N_1108,N_1051,N_1004);
or U1109 (N_1109,N_1001,N_1018);
or U1110 (N_1110,N_1014,N_1059);
nor U1111 (N_1111,N_1053,N_1009);
nand U1112 (N_1112,N_1090,N_1049);
and U1113 (N_1113,N_1068,N_1075);
xor U1114 (N_1114,N_1098,N_1050);
and U1115 (N_1115,N_1030,N_1029);
and U1116 (N_1116,N_1093,N_1076);
and U1117 (N_1117,N_1074,N_1037);
nand U1118 (N_1118,N_1071,N_1000);
and U1119 (N_1119,N_1025,N_1063);
nor U1120 (N_1120,N_1016,N_1060);
nor U1121 (N_1121,N_1026,N_1058);
and U1122 (N_1122,N_1036,N_1023);
and U1123 (N_1123,N_1043,N_1045);
and U1124 (N_1124,N_1038,N_1027);
nor U1125 (N_1125,N_1094,N_1034);
or U1126 (N_1126,N_1047,N_1086);
or U1127 (N_1127,N_1070,N_1057);
nor U1128 (N_1128,N_1096,N_1092);
or U1129 (N_1129,N_1095,N_1056);
nand U1130 (N_1130,N_1097,N_1083);
and U1131 (N_1131,N_1065,N_1062);
or U1132 (N_1132,N_1041,N_1011);
and U1133 (N_1133,N_1061,N_1072);
or U1134 (N_1134,N_1024,N_1040);
nand U1135 (N_1135,N_1088,N_1064);
nor U1136 (N_1136,N_1044,N_1081);
xnor U1137 (N_1137,N_1042,N_1089);
nor U1138 (N_1138,N_1003,N_1035);
and U1139 (N_1139,N_1087,N_1010);
nor U1140 (N_1140,N_1078,N_1052);
nor U1141 (N_1141,N_1073,N_1007);
or U1142 (N_1142,N_1099,N_1012);
and U1143 (N_1143,N_1085,N_1077);
or U1144 (N_1144,N_1084,N_1006);
and U1145 (N_1145,N_1080,N_1067);
xor U1146 (N_1146,N_1079,N_1013);
nor U1147 (N_1147,N_1046,N_1091);
nor U1148 (N_1148,N_1017,N_1033);
and U1149 (N_1149,N_1039,N_1054);
and U1150 (N_1150,N_1032,N_1010);
xnor U1151 (N_1151,N_1043,N_1089);
nand U1152 (N_1152,N_1068,N_1001);
and U1153 (N_1153,N_1083,N_1041);
nor U1154 (N_1154,N_1017,N_1098);
nor U1155 (N_1155,N_1015,N_1008);
or U1156 (N_1156,N_1017,N_1013);
nor U1157 (N_1157,N_1008,N_1051);
xnor U1158 (N_1158,N_1059,N_1061);
nand U1159 (N_1159,N_1069,N_1043);
and U1160 (N_1160,N_1076,N_1085);
nand U1161 (N_1161,N_1006,N_1081);
nand U1162 (N_1162,N_1041,N_1052);
nand U1163 (N_1163,N_1020,N_1075);
or U1164 (N_1164,N_1077,N_1046);
and U1165 (N_1165,N_1027,N_1026);
and U1166 (N_1166,N_1068,N_1023);
nand U1167 (N_1167,N_1093,N_1033);
nand U1168 (N_1168,N_1013,N_1045);
nand U1169 (N_1169,N_1012,N_1071);
nor U1170 (N_1170,N_1061,N_1087);
nor U1171 (N_1171,N_1032,N_1090);
xnor U1172 (N_1172,N_1055,N_1005);
xor U1173 (N_1173,N_1071,N_1055);
or U1174 (N_1174,N_1041,N_1045);
nor U1175 (N_1175,N_1050,N_1034);
nor U1176 (N_1176,N_1056,N_1034);
nor U1177 (N_1177,N_1008,N_1084);
nand U1178 (N_1178,N_1022,N_1021);
nand U1179 (N_1179,N_1090,N_1095);
or U1180 (N_1180,N_1019,N_1095);
nor U1181 (N_1181,N_1030,N_1072);
or U1182 (N_1182,N_1097,N_1042);
nor U1183 (N_1183,N_1085,N_1009);
or U1184 (N_1184,N_1093,N_1024);
xor U1185 (N_1185,N_1063,N_1030);
nand U1186 (N_1186,N_1058,N_1065);
or U1187 (N_1187,N_1096,N_1059);
or U1188 (N_1188,N_1008,N_1067);
xor U1189 (N_1189,N_1082,N_1044);
and U1190 (N_1190,N_1027,N_1085);
xnor U1191 (N_1191,N_1034,N_1054);
nand U1192 (N_1192,N_1061,N_1000);
nand U1193 (N_1193,N_1060,N_1096);
xor U1194 (N_1194,N_1031,N_1047);
or U1195 (N_1195,N_1025,N_1054);
or U1196 (N_1196,N_1084,N_1011);
or U1197 (N_1197,N_1086,N_1065);
or U1198 (N_1198,N_1004,N_1099);
nor U1199 (N_1199,N_1050,N_1058);
nor U1200 (N_1200,N_1134,N_1160);
and U1201 (N_1201,N_1172,N_1184);
nor U1202 (N_1202,N_1169,N_1143);
or U1203 (N_1203,N_1187,N_1100);
or U1204 (N_1204,N_1135,N_1153);
and U1205 (N_1205,N_1103,N_1101);
and U1206 (N_1206,N_1102,N_1141);
nor U1207 (N_1207,N_1198,N_1195);
and U1208 (N_1208,N_1157,N_1197);
xor U1209 (N_1209,N_1130,N_1183);
and U1210 (N_1210,N_1167,N_1155);
nor U1211 (N_1211,N_1137,N_1148);
nor U1212 (N_1212,N_1173,N_1149);
and U1213 (N_1213,N_1161,N_1193);
xnor U1214 (N_1214,N_1162,N_1132);
nor U1215 (N_1215,N_1185,N_1182);
and U1216 (N_1216,N_1147,N_1179);
and U1217 (N_1217,N_1196,N_1145);
xor U1218 (N_1218,N_1146,N_1163);
or U1219 (N_1219,N_1123,N_1138);
nor U1220 (N_1220,N_1122,N_1117);
and U1221 (N_1221,N_1154,N_1109);
or U1222 (N_1222,N_1125,N_1128);
nor U1223 (N_1223,N_1116,N_1139);
nor U1224 (N_1224,N_1112,N_1181);
or U1225 (N_1225,N_1118,N_1107);
nor U1226 (N_1226,N_1188,N_1140);
or U1227 (N_1227,N_1192,N_1165);
or U1228 (N_1228,N_1175,N_1152);
nor U1229 (N_1229,N_1151,N_1121);
or U1230 (N_1230,N_1120,N_1124);
and U1231 (N_1231,N_1186,N_1199);
or U1232 (N_1232,N_1177,N_1106);
nor U1233 (N_1233,N_1105,N_1190);
nor U1234 (N_1234,N_1166,N_1142);
or U1235 (N_1235,N_1164,N_1129);
nand U1236 (N_1236,N_1191,N_1110);
nor U1237 (N_1237,N_1180,N_1178);
or U1238 (N_1238,N_1108,N_1136);
or U1239 (N_1239,N_1176,N_1104);
nand U1240 (N_1240,N_1114,N_1115);
or U1241 (N_1241,N_1127,N_1194);
and U1242 (N_1242,N_1170,N_1113);
nand U1243 (N_1243,N_1150,N_1168);
and U1244 (N_1244,N_1133,N_1174);
and U1245 (N_1245,N_1111,N_1156);
or U1246 (N_1246,N_1158,N_1189);
xor U1247 (N_1247,N_1131,N_1171);
and U1248 (N_1248,N_1144,N_1126);
nor U1249 (N_1249,N_1119,N_1159);
nand U1250 (N_1250,N_1156,N_1133);
nand U1251 (N_1251,N_1164,N_1189);
nor U1252 (N_1252,N_1132,N_1185);
and U1253 (N_1253,N_1121,N_1179);
or U1254 (N_1254,N_1124,N_1134);
nor U1255 (N_1255,N_1181,N_1115);
xnor U1256 (N_1256,N_1167,N_1129);
nand U1257 (N_1257,N_1172,N_1149);
and U1258 (N_1258,N_1184,N_1159);
xnor U1259 (N_1259,N_1186,N_1151);
or U1260 (N_1260,N_1144,N_1161);
or U1261 (N_1261,N_1107,N_1145);
nand U1262 (N_1262,N_1129,N_1157);
nor U1263 (N_1263,N_1131,N_1152);
or U1264 (N_1264,N_1135,N_1136);
or U1265 (N_1265,N_1189,N_1126);
and U1266 (N_1266,N_1105,N_1108);
or U1267 (N_1267,N_1103,N_1143);
xor U1268 (N_1268,N_1166,N_1177);
nand U1269 (N_1269,N_1178,N_1162);
or U1270 (N_1270,N_1132,N_1126);
nand U1271 (N_1271,N_1101,N_1100);
nand U1272 (N_1272,N_1122,N_1149);
or U1273 (N_1273,N_1162,N_1159);
nand U1274 (N_1274,N_1100,N_1114);
nor U1275 (N_1275,N_1188,N_1131);
or U1276 (N_1276,N_1170,N_1127);
and U1277 (N_1277,N_1117,N_1155);
nor U1278 (N_1278,N_1125,N_1131);
or U1279 (N_1279,N_1128,N_1105);
and U1280 (N_1280,N_1199,N_1111);
or U1281 (N_1281,N_1117,N_1175);
xnor U1282 (N_1282,N_1156,N_1159);
xnor U1283 (N_1283,N_1181,N_1158);
and U1284 (N_1284,N_1106,N_1149);
nand U1285 (N_1285,N_1135,N_1120);
nor U1286 (N_1286,N_1134,N_1149);
or U1287 (N_1287,N_1141,N_1103);
xor U1288 (N_1288,N_1182,N_1125);
and U1289 (N_1289,N_1179,N_1163);
xnor U1290 (N_1290,N_1152,N_1196);
nor U1291 (N_1291,N_1165,N_1171);
or U1292 (N_1292,N_1101,N_1160);
or U1293 (N_1293,N_1165,N_1177);
and U1294 (N_1294,N_1166,N_1192);
or U1295 (N_1295,N_1168,N_1180);
and U1296 (N_1296,N_1120,N_1129);
and U1297 (N_1297,N_1118,N_1173);
nand U1298 (N_1298,N_1124,N_1114);
nand U1299 (N_1299,N_1133,N_1153);
nand U1300 (N_1300,N_1277,N_1270);
xnor U1301 (N_1301,N_1274,N_1212);
and U1302 (N_1302,N_1272,N_1244);
nand U1303 (N_1303,N_1266,N_1287);
or U1304 (N_1304,N_1225,N_1202);
nand U1305 (N_1305,N_1226,N_1201);
nand U1306 (N_1306,N_1298,N_1257);
or U1307 (N_1307,N_1261,N_1262);
and U1308 (N_1308,N_1264,N_1234);
nor U1309 (N_1309,N_1281,N_1250);
and U1310 (N_1310,N_1288,N_1218);
and U1311 (N_1311,N_1236,N_1258);
xnor U1312 (N_1312,N_1299,N_1240);
and U1313 (N_1313,N_1278,N_1271);
nand U1314 (N_1314,N_1200,N_1228);
nand U1315 (N_1315,N_1224,N_1291);
nand U1316 (N_1316,N_1283,N_1233);
and U1317 (N_1317,N_1211,N_1248);
or U1318 (N_1318,N_1210,N_1252);
nor U1319 (N_1319,N_1232,N_1221);
nand U1320 (N_1320,N_1247,N_1245);
nor U1321 (N_1321,N_1259,N_1239);
nand U1322 (N_1322,N_1205,N_1251);
xnor U1323 (N_1323,N_1249,N_1222);
and U1324 (N_1324,N_1294,N_1276);
and U1325 (N_1325,N_1273,N_1297);
or U1326 (N_1326,N_1207,N_1254);
nor U1327 (N_1327,N_1229,N_1296);
or U1328 (N_1328,N_1267,N_1208);
or U1329 (N_1329,N_1204,N_1293);
nand U1330 (N_1330,N_1243,N_1265);
nand U1331 (N_1331,N_1213,N_1255);
nor U1332 (N_1332,N_1206,N_1231);
and U1333 (N_1333,N_1289,N_1295);
and U1334 (N_1334,N_1253,N_1269);
nor U1335 (N_1335,N_1282,N_1219);
and U1336 (N_1336,N_1238,N_1275);
and U1337 (N_1337,N_1214,N_1235);
nor U1338 (N_1338,N_1279,N_1209);
and U1339 (N_1339,N_1227,N_1242);
nand U1340 (N_1340,N_1290,N_1223);
xor U1341 (N_1341,N_1217,N_1260);
xor U1342 (N_1342,N_1263,N_1256);
and U1343 (N_1343,N_1230,N_1215);
nand U1344 (N_1344,N_1285,N_1220);
or U1345 (N_1345,N_1268,N_1216);
and U1346 (N_1346,N_1246,N_1203);
or U1347 (N_1347,N_1286,N_1292);
xnor U1348 (N_1348,N_1280,N_1284);
xnor U1349 (N_1349,N_1237,N_1241);
xnor U1350 (N_1350,N_1228,N_1283);
nand U1351 (N_1351,N_1212,N_1287);
nor U1352 (N_1352,N_1251,N_1226);
or U1353 (N_1353,N_1267,N_1276);
or U1354 (N_1354,N_1282,N_1228);
nor U1355 (N_1355,N_1213,N_1244);
nand U1356 (N_1356,N_1201,N_1250);
nor U1357 (N_1357,N_1262,N_1205);
and U1358 (N_1358,N_1294,N_1219);
or U1359 (N_1359,N_1265,N_1264);
nor U1360 (N_1360,N_1272,N_1241);
or U1361 (N_1361,N_1245,N_1290);
xnor U1362 (N_1362,N_1240,N_1290);
or U1363 (N_1363,N_1266,N_1241);
nand U1364 (N_1364,N_1239,N_1251);
nor U1365 (N_1365,N_1298,N_1223);
or U1366 (N_1366,N_1283,N_1204);
and U1367 (N_1367,N_1287,N_1271);
and U1368 (N_1368,N_1226,N_1210);
nor U1369 (N_1369,N_1276,N_1213);
nand U1370 (N_1370,N_1222,N_1264);
nor U1371 (N_1371,N_1208,N_1237);
nand U1372 (N_1372,N_1296,N_1264);
and U1373 (N_1373,N_1246,N_1217);
xor U1374 (N_1374,N_1258,N_1274);
and U1375 (N_1375,N_1294,N_1207);
and U1376 (N_1376,N_1227,N_1285);
nor U1377 (N_1377,N_1276,N_1272);
or U1378 (N_1378,N_1228,N_1267);
or U1379 (N_1379,N_1252,N_1264);
and U1380 (N_1380,N_1214,N_1239);
nor U1381 (N_1381,N_1272,N_1224);
nor U1382 (N_1382,N_1231,N_1220);
or U1383 (N_1383,N_1226,N_1271);
and U1384 (N_1384,N_1296,N_1249);
nand U1385 (N_1385,N_1258,N_1287);
and U1386 (N_1386,N_1245,N_1269);
nor U1387 (N_1387,N_1273,N_1220);
or U1388 (N_1388,N_1237,N_1265);
nor U1389 (N_1389,N_1201,N_1242);
nor U1390 (N_1390,N_1286,N_1226);
nor U1391 (N_1391,N_1222,N_1286);
nand U1392 (N_1392,N_1264,N_1279);
xnor U1393 (N_1393,N_1280,N_1207);
nor U1394 (N_1394,N_1258,N_1248);
and U1395 (N_1395,N_1252,N_1250);
nand U1396 (N_1396,N_1227,N_1230);
xnor U1397 (N_1397,N_1290,N_1289);
nor U1398 (N_1398,N_1223,N_1240);
nor U1399 (N_1399,N_1242,N_1245);
or U1400 (N_1400,N_1352,N_1356);
or U1401 (N_1401,N_1331,N_1308);
nand U1402 (N_1402,N_1368,N_1305);
nor U1403 (N_1403,N_1391,N_1371);
xor U1404 (N_1404,N_1375,N_1383);
nand U1405 (N_1405,N_1379,N_1323);
xor U1406 (N_1406,N_1392,N_1319);
nor U1407 (N_1407,N_1318,N_1369);
and U1408 (N_1408,N_1328,N_1316);
nand U1409 (N_1409,N_1300,N_1354);
xor U1410 (N_1410,N_1311,N_1387);
nand U1411 (N_1411,N_1361,N_1340);
nor U1412 (N_1412,N_1389,N_1326);
and U1413 (N_1413,N_1343,N_1336);
nand U1414 (N_1414,N_1386,N_1370);
and U1415 (N_1415,N_1362,N_1344);
or U1416 (N_1416,N_1376,N_1381);
or U1417 (N_1417,N_1333,N_1312);
and U1418 (N_1418,N_1398,N_1353);
nand U1419 (N_1419,N_1338,N_1394);
xnor U1420 (N_1420,N_1324,N_1365);
and U1421 (N_1421,N_1395,N_1378);
nor U1422 (N_1422,N_1337,N_1355);
nor U1423 (N_1423,N_1346,N_1329);
nor U1424 (N_1424,N_1306,N_1372);
nand U1425 (N_1425,N_1399,N_1303);
nand U1426 (N_1426,N_1384,N_1350);
and U1427 (N_1427,N_1339,N_1390);
or U1428 (N_1428,N_1304,N_1347);
and U1429 (N_1429,N_1309,N_1320);
nor U1430 (N_1430,N_1366,N_1382);
nor U1431 (N_1431,N_1325,N_1364);
and U1432 (N_1432,N_1385,N_1327);
nand U1433 (N_1433,N_1380,N_1313);
nor U1434 (N_1434,N_1334,N_1393);
nor U1435 (N_1435,N_1335,N_1315);
or U1436 (N_1436,N_1396,N_1307);
and U1437 (N_1437,N_1322,N_1332);
nor U1438 (N_1438,N_1397,N_1317);
nor U1439 (N_1439,N_1349,N_1330);
or U1440 (N_1440,N_1360,N_1348);
or U1441 (N_1441,N_1310,N_1377);
nand U1442 (N_1442,N_1351,N_1321);
nor U1443 (N_1443,N_1302,N_1342);
nand U1444 (N_1444,N_1374,N_1345);
or U1445 (N_1445,N_1363,N_1359);
or U1446 (N_1446,N_1341,N_1388);
nand U1447 (N_1447,N_1367,N_1373);
or U1448 (N_1448,N_1358,N_1301);
nand U1449 (N_1449,N_1314,N_1357);
nor U1450 (N_1450,N_1347,N_1307);
and U1451 (N_1451,N_1352,N_1344);
nor U1452 (N_1452,N_1342,N_1354);
nor U1453 (N_1453,N_1356,N_1362);
nor U1454 (N_1454,N_1337,N_1371);
and U1455 (N_1455,N_1312,N_1346);
and U1456 (N_1456,N_1310,N_1361);
nand U1457 (N_1457,N_1371,N_1396);
and U1458 (N_1458,N_1398,N_1363);
nor U1459 (N_1459,N_1337,N_1303);
and U1460 (N_1460,N_1313,N_1306);
xor U1461 (N_1461,N_1397,N_1307);
nand U1462 (N_1462,N_1373,N_1310);
and U1463 (N_1463,N_1307,N_1301);
nor U1464 (N_1464,N_1364,N_1365);
nor U1465 (N_1465,N_1311,N_1303);
or U1466 (N_1466,N_1334,N_1327);
nand U1467 (N_1467,N_1354,N_1313);
or U1468 (N_1468,N_1356,N_1378);
nand U1469 (N_1469,N_1304,N_1335);
or U1470 (N_1470,N_1334,N_1342);
and U1471 (N_1471,N_1364,N_1328);
or U1472 (N_1472,N_1355,N_1369);
nand U1473 (N_1473,N_1318,N_1357);
xor U1474 (N_1474,N_1320,N_1314);
and U1475 (N_1475,N_1382,N_1307);
nor U1476 (N_1476,N_1375,N_1330);
or U1477 (N_1477,N_1310,N_1336);
xnor U1478 (N_1478,N_1375,N_1390);
xor U1479 (N_1479,N_1337,N_1393);
or U1480 (N_1480,N_1384,N_1348);
xnor U1481 (N_1481,N_1340,N_1335);
nand U1482 (N_1482,N_1332,N_1303);
nor U1483 (N_1483,N_1363,N_1341);
and U1484 (N_1484,N_1315,N_1346);
and U1485 (N_1485,N_1359,N_1376);
xor U1486 (N_1486,N_1317,N_1301);
and U1487 (N_1487,N_1331,N_1309);
nor U1488 (N_1488,N_1394,N_1324);
nor U1489 (N_1489,N_1328,N_1378);
and U1490 (N_1490,N_1355,N_1362);
or U1491 (N_1491,N_1367,N_1304);
nor U1492 (N_1492,N_1374,N_1391);
or U1493 (N_1493,N_1321,N_1381);
and U1494 (N_1494,N_1358,N_1376);
and U1495 (N_1495,N_1365,N_1378);
or U1496 (N_1496,N_1358,N_1371);
nor U1497 (N_1497,N_1303,N_1353);
and U1498 (N_1498,N_1340,N_1382);
nor U1499 (N_1499,N_1346,N_1367);
nand U1500 (N_1500,N_1453,N_1419);
or U1501 (N_1501,N_1424,N_1462);
nor U1502 (N_1502,N_1404,N_1497);
nand U1503 (N_1503,N_1466,N_1484);
and U1504 (N_1504,N_1483,N_1454);
nand U1505 (N_1505,N_1433,N_1486);
nor U1506 (N_1506,N_1494,N_1426);
and U1507 (N_1507,N_1490,N_1458);
and U1508 (N_1508,N_1413,N_1444);
nor U1509 (N_1509,N_1475,N_1415);
and U1510 (N_1510,N_1461,N_1428);
nand U1511 (N_1511,N_1438,N_1498);
or U1512 (N_1512,N_1409,N_1481);
nor U1513 (N_1513,N_1446,N_1429);
or U1514 (N_1514,N_1499,N_1423);
or U1515 (N_1515,N_1439,N_1408);
nor U1516 (N_1516,N_1401,N_1478);
nand U1517 (N_1517,N_1440,N_1487);
nand U1518 (N_1518,N_1434,N_1437);
nor U1519 (N_1519,N_1464,N_1447);
or U1520 (N_1520,N_1435,N_1422);
nor U1521 (N_1521,N_1489,N_1456);
and U1522 (N_1522,N_1493,N_1449);
nor U1523 (N_1523,N_1436,N_1476);
nand U1524 (N_1524,N_1406,N_1425);
nor U1525 (N_1525,N_1414,N_1495);
xnor U1526 (N_1526,N_1431,N_1421);
or U1527 (N_1527,N_1482,N_1488);
or U1528 (N_1528,N_1479,N_1491);
and U1529 (N_1529,N_1410,N_1469);
nand U1530 (N_1530,N_1432,N_1427);
and U1531 (N_1531,N_1448,N_1411);
or U1532 (N_1532,N_1473,N_1430);
or U1533 (N_1533,N_1452,N_1455);
and U1534 (N_1534,N_1471,N_1492);
and U1535 (N_1535,N_1463,N_1460);
or U1536 (N_1536,N_1402,N_1412);
and U1537 (N_1537,N_1467,N_1465);
xor U1538 (N_1538,N_1496,N_1420);
nor U1539 (N_1539,N_1403,N_1445);
nand U1540 (N_1540,N_1441,N_1459);
and U1541 (N_1541,N_1457,N_1418);
and U1542 (N_1542,N_1443,N_1477);
nor U1543 (N_1543,N_1451,N_1405);
nor U1544 (N_1544,N_1407,N_1417);
and U1545 (N_1545,N_1485,N_1474);
nor U1546 (N_1546,N_1442,N_1450);
nor U1547 (N_1547,N_1472,N_1416);
or U1548 (N_1548,N_1480,N_1468);
and U1549 (N_1549,N_1470,N_1400);
or U1550 (N_1550,N_1407,N_1460);
xor U1551 (N_1551,N_1467,N_1438);
or U1552 (N_1552,N_1450,N_1492);
xnor U1553 (N_1553,N_1476,N_1457);
nor U1554 (N_1554,N_1499,N_1409);
xor U1555 (N_1555,N_1479,N_1403);
nor U1556 (N_1556,N_1421,N_1443);
or U1557 (N_1557,N_1462,N_1443);
or U1558 (N_1558,N_1466,N_1435);
xor U1559 (N_1559,N_1489,N_1402);
nand U1560 (N_1560,N_1485,N_1491);
or U1561 (N_1561,N_1454,N_1463);
nand U1562 (N_1562,N_1488,N_1499);
or U1563 (N_1563,N_1404,N_1450);
nor U1564 (N_1564,N_1412,N_1451);
nor U1565 (N_1565,N_1445,N_1434);
nor U1566 (N_1566,N_1462,N_1469);
or U1567 (N_1567,N_1499,N_1492);
nor U1568 (N_1568,N_1458,N_1422);
nor U1569 (N_1569,N_1466,N_1489);
or U1570 (N_1570,N_1473,N_1434);
nor U1571 (N_1571,N_1415,N_1433);
nor U1572 (N_1572,N_1412,N_1490);
nor U1573 (N_1573,N_1482,N_1424);
and U1574 (N_1574,N_1495,N_1488);
or U1575 (N_1575,N_1491,N_1414);
nor U1576 (N_1576,N_1483,N_1477);
nand U1577 (N_1577,N_1454,N_1439);
nand U1578 (N_1578,N_1441,N_1455);
and U1579 (N_1579,N_1442,N_1414);
or U1580 (N_1580,N_1494,N_1428);
and U1581 (N_1581,N_1454,N_1430);
nor U1582 (N_1582,N_1489,N_1457);
or U1583 (N_1583,N_1464,N_1418);
nor U1584 (N_1584,N_1456,N_1414);
or U1585 (N_1585,N_1445,N_1440);
and U1586 (N_1586,N_1411,N_1479);
xor U1587 (N_1587,N_1461,N_1402);
nand U1588 (N_1588,N_1402,N_1436);
nor U1589 (N_1589,N_1486,N_1487);
and U1590 (N_1590,N_1467,N_1433);
nor U1591 (N_1591,N_1414,N_1463);
nand U1592 (N_1592,N_1406,N_1411);
nand U1593 (N_1593,N_1487,N_1416);
nor U1594 (N_1594,N_1435,N_1462);
or U1595 (N_1595,N_1499,N_1438);
or U1596 (N_1596,N_1417,N_1412);
nor U1597 (N_1597,N_1409,N_1432);
or U1598 (N_1598,N_1439,N_1414);
nand U1599 (N_1599,N_1447,N_1448);
and U1600 (N_1600,N_1584,N_1524);
and U1601 (N_1601,N_1592,N_1599);
and U1602 (N_1602,N_1563,N_1559);
nor U1603 (N_1603,N_1539,N_1527);
xnor U1604 (N_1604,N_1582,N_1503);
and U1605 (N_1605,N_1572,N_1530);
nor U1606 (N_1606,N_1511,N_1594);
nand U1607 (N_1607,N_1567,N_1518);
and U1608 (N_1608,N_1564,N_1502);
nand U1609 (N_1609,N_1566,N_1551);
or U1610 (N_1610,N_1583,N_1580);
and U1611 (N_1611,N_1519,N_1522);
or U1612 (N_1612,N_1509,N_1533);
nor U1613 (N_1613,N_1545,N_1595);
nand U1614 (N_1614,N_1571,N_1500);
and U1615 (N_1615,N_1535,N_1516);
nor U1616 (N_1616,N_1529,N_1531);
or U1617 (N_1617,N_1510,N_1525);
and U1618 (N_1618,N_1561,N_1515);
nand U1619 (N_1619,N_1555,N_1578);
nand U1620 (N_1620,N_1590,N_1586);
nand U1621 (N_1621,N_1543,N_1593);
or U1622 (N_1622,N_1556,N_1534);
or U1623 (N_1623,N_1520,N_1577);
nor U1624 (N_1624,N_1540,N_1576);
nand U1625 (N_1625,N_1588,N_1597);
nor U1626 (N_1626,N_1513,N_1512);
xnor U1627 (N_1627,N_1506,N_1547);
nor U1628 (N_1628,N_1565,N_1562);
nand U1629 (N_1629,N_1532,N_1574);
or U1630 (N_1630,N_1526,N_1507);
nor U1631 (N_1631,N_1589,N_1596);
and U1632 (N_1632,N_1560,N_1541);
nor U1633 (N_1633,N_1553,N_1504);
and U1634 (N_1634,N_1517,N_1508);
or U1635 (N_1635,N_1521,N_1536);
and U1636 (N_1636,N_1523,N_1575);
nor U1637 (N_1637,N_1591,N_1514);
and U1638 (N_1638,N_1554,N_1568);
nor U1639 (N_1639,N_1528,N_1550);
nor U1640 (N_1640,N_1573,N_1569);
or U1641 (N_1641,N_1537,N_1585);
or U1642 (N_1642,N_1581,N_1557);
or U1643 (N_1643,N_1542,N_1505);
xor U1644 (N_1644,N_1570,N_1544);
nor U1645 (N_1645,N_1587,N_1546);
or U1646 (N_1646,N_1558,N_1538);
or U1647 (N_1647,N_1598,N_1548);
nand U1648 (N_1648,N_1552,N_1501);
or U1649 (N_1649,N_1549,N_1579);
nand U1650 (N_1650,N_1593,N_1595);
nor U1651 (N_1651,N_1584,N_1543);
and U1652 (N_1652,N_1522,N_1588);
or U1653 (N_1653,N_1521,N_1510);
nand U1654 (N_1654,N_1556,N_1537);
and U1655 (N_1655,N_1576,N_1564);
xnor U1656 (N_1656,N_1526,N_1510);
nand U1657 (N_1657,N_1558,N_1582);
nor U1658 (N_1658,N_1506,N_1598);
nor U1659 (N_1659,N_1573,N_1506);
nor U1660 (N_1660,N_1555,N_1503);
and U1661 (N_1661,N_1577,N_1540);
xor U1662 (N_1662,N_1554,N_1531);
or U1663 (N_1663,N_1513,N_1555);
nand U1664 (N_1664,N_1574,N_1570);
nand U1665 (N_1665,N_1559,N_1525);
or U1666 (N_1666,N_1597,N_1596);
or U1667 (N_1667,N_1537,N_1571);
or U1668 (N_1668,N_1552,N_1532);
or U1669 (N_1669,N_1517,N_1520);
or U1670 (N_1670,N_1539,N_1555);
nor U1671 (N_1671,N_1584,N_1540);
nand U1672 (N_1672,N_1571,N_1596);
nor U1673 (N_1673,N_1528,N_1597);
and U1674 (N_1674,N_1551,N_1529);
or U1675 (N_1675,N_1564,N_1531);
and U1676 (N_1676,N_1554,N_1591);
nor U1677 (N_1677,N_1595,N_1526);
and U1678 (N_1678,N_1573,N_1528);
or U1679 (N_1679,N_1522,N_1550);
and U1680 (N_1680,N_1527,N_1535);
and U1681 (N_1681,N_1531,N_1599);
or U1682 (N_1682,N_1551,N_1508);
nand U1683 (N_1683,N_1592,N_1533);
nor U1684 (N_1684,N_1577,N_1583);
nor U1685 (N_1685,N_1564,N_1563);
nor U1686 (N_1686,N_1548,N_1557);
and U1687 (N_1687,N_1520,N_1533);
and U1688 (N_1688,N_1593,N_1572);
and U1689 (N_1689,N_1541,N_1576);
or U1690 (N_1690,N_1571,N_1577);
or U1691 (N_1691,N_1502,N_1537);
nand U1692 (N_1692,N_1527,N_1521);
xor U1693 (N_1693,N_1591,N_1577);
and U1694 (N_1694,N_1570,N_1550);
nor U1695 (N_1695,N_1537,N_1534);
nand U1696 (N_1696,N_1501,N_1557);
nand U1697 (N_1697,N_1538,N_1593);
and U1698 (N_1698,N_1598,N_1546);
nor U1699 (N_1699,N_1571,N_1563);
xor U1700 (N_1700,N_1648,N_1639);
and U1701 (N_1701,N_1633,N_1617);
or U1702 (N_1702,N_1664,N_1645);
nor U1703 (N_1703,N_1638,N_1632);
or U1704 (N_1704,N_1650,N_1622);
nand U1705 (N_1705,N_1687,N_1663);
and U1706 (N_1706,N_1618,N_1676);
and U1707 (N_1707,N_1651,N_1691);
and U1708 (N_1708,N_1655,N_1681);
and U1709 (N_1709,N_1644,N_1693);
xor U1710 (N_1710,N_1688,N_1669);
or U1711 (N_1711,N_1671,N_1656);
nor U1712 (N_1712,N_1699,N_1609);
nand U1713 (N_1713,N_1659,N_1692);
nand U1714 (N_1714,N_1649,N_1696);
xnor U1715 (N_1715,N_1625,N_1602);
nand U1716 (N_1716,N_1654,N_1642);
or U1717 (N_1717,N_1640,N_1653);
nor U1718 (N_1718,N_1606,N_1662);
or U1719 (N_1719,N_1629,N_1636);
and U1720 (N_1720,N_1667,N_1660);
nand U1721 (N_1721,N_1658,N_1698);
nand U1722 (N_1722,N_1635,N_1601);
nand U1723 (N_1723,N_1685,N_1603);
or U1724 (N_1724,N_1689,N_1674);
nand U1725 (N_1725,N_1621,N_1668);
nand U1726 (N_1726,N_1657,N_1661);
xnor U1727 (N_1727,N_1647,N_1683);
nor U1728 (N_1728,N_1605,N_1612);
or U1729 (N_1729,N_1678,N_1686);
nand U1730 (N_1730,N_1624,N_1611);
or U1731 (N_1731,N_1652,N_1675);
nand U1732 (N_1732,N_1614,N_1680);
or U1733 (N_1733,N_1630,N_1684);
xor U1734 (N_1734,N_1682,N_1608);
or U1735 (N_1735,N_1600,N_1604);
or U1736 (N_1736,N_1670,N_1641);
or U1737 (N_1737,N_1697,N_1677);
and U1738 (N_1738,N_1665,N_1694);
nand U1739 (N_1739,N_1690,N_1620);
or U1740 (N_1740,N_1643,N_1679);
or U1741 (N_1741,N_1673,N_1628);
or U1742 (N_1742,N_1615,N_1607);
and U1743 (N_1743,N_1626,N_1672);
nand U1744 (N_1744,N_1619,N_1627);
nand U1745 (N_1745,N_1637,N_1623);
and U1746 (N_1746,N_1613,N_1610);
and U1747 (N_1747,N_1634,N_1666);
nor U1748 (N_1748,N_1631,N_1695);
xnor U1749 (N_1749,N_1646,N_1616);
nand U1750 (N_1750,N_1676,N_1671);
nor U1751 (N_1751,N_1601,N_1668);
nand U1752 (N_1752,N_1692,N_1600);
or U1753 (N_1753,N_1676,N_1686);
or U1754 (N_1754,N_1684,N_1656);
or U1755 (N_1755,N_1653,N_1667);
nand U1756 (N_1756,N_1600,N_1617);
or U1757 (N_1757,N_1602,N_1662);
nand U1758 (N_1758,N_1610,N_1629);
xnor U1759 (N_1759,N_1660,N_1642);
nor U1760 (N_1760,N_1661,N_1608);
xnor U1761 (N_1761,N_1650,N_1695);
nor U1762 (N_1762,N_1613,N_1603);
and U1763 (N_1763,N_1627,N_1607);
xor U1764 (N_1764,N_1628,N_1603);
or U1765 (N_1765,N_1672,N_1646);
nor U1766 (N_1766,N_1629,N_1622);
xnor U1767 (N_1767,N_1643,N_1621);
or U1768 (N_1768,N_1601,N_1648);
or U1769 (N_1769,N_1618,N_1607);
xor U1770 (N_1770,N_1609,N_1607);
nand U1771 (N_1771,N_1629,N_1685);
xor U1772 (N_1772,N_1614,N_1637);
or U1773 (N_1773,N_1632,N_1619);
or U1774 (N_1774,N_1608,N_1691);
or U1775 (N_1775,N_1656,N_1695);
nor U1776 (N_1776,N_1624,N_1605);
and U1777 (N_1777,N_1677,N_1674);
or U1778 (N_1778,N_1665,N_1653);
or U1779 (N_1779,N_1675,N_1617);
or U1780 (N_1780,N_1601,N_1666);
or U1781 (N_1781,N_1672,N_1664);
and U1782 (N_1782,N_1607,N_1674);
nor U1783 (N_1783,N_1626,N_1637);
nor U1784 (N_1784,N_1634,N_1636);
and U1785 (N_1785,N_1669,N_1684);
and U1786 (N_1786,N_1693,N_1671);
and U1787 (N_1787,N_1628,N_1663);
nand U1788 (N_1788,N_1623,N_1641);
nor U1789 (N_1789,N_1643,N_1605);
nor U1790 (N_1790,N_1665,N_1685);
or U1791 (N_1791,N_1671,N_1605);
nor U1792 (N_1792,N_1653,N_1629);
nand U1793 (N_1793,N_1683,N_1627);
xnor U1794 (N_1794,N_1656,N_1660);
and U1795 (N_1795,N_1637,N_1663);
nand U1796 (N_1796,N_1695,N_1635);
nor U1797 (N_1797,N_1620,N_1637);
xnor U1798 (N_1798,N_1695,N_1605);
nand U1799 (N_1799,N_1630,N_1628);
and U1800 (N_1800,N_1732,N_1739);
or U1801 (N_1801,N_1770,N_1772);
nand U1802 (N_1802,N_1792,N_1786);
nor U1803 (N_1803,N_1765,N_1768);
nand U1804 (N_1804,N_1734,N_1767);
nand U1805 (N_1805,N_1716,N_1711);
nand U1806 (N_1806,N_1777,N_1722);
nand U1807 (N_1807,N_1728,N_1738);
and U1808 (N_1808,N_1727,N_1759);
nor U1809 (N_1809,N_1721,N_1729);
and U1810 (N_1810,N_1785,N_1713);
nand U1811 (N_1811,N_1758,N_1710);
or U1812 (N_1812,N_1782,N_1714);
xor U1813 (N_1813,N_1730,N_1771);
xnor U1814 (N_1814,N_1720,N_1702);
or U1815 (N_1815,N_1784,N_1725);
or U1816 (N_1816,N_1778,N_1715);
or U1817 (N_1817,N_1747,N_1737);
xnor U1818 (N_1818,N_1773,N_1700);
nand U1819 (N_1819,N_1726,N_1744);
nor U1820 (N_1820,N_1752,N_1746);
nor U1821 (N_1821,N_1798,N_1775);
nand U1822 (N_1822,N_1799,N_1751);
nor U1823 (N_1823,N_1709,N_1701);
nor U1824 (N_1824,N_1763,N_1795);
and U1825 (N_1825,N_1733,N_1757);
nand U1826 (N_1826,N_1797,N_1750);
or U1827 (N_1827,N_1736,N_1742);
and U1828 (N_1828,N_1760,N_1735);
or U1829 (N_1829,N_1724,N_1756);
or U1830 (N_1830,N_1703,N_1790);
and U1831 (N_1831,N_1780,N_1755);
nand U1832 (N_1832,N_1761,N_1769);
xor U1833 (N_1833,N_1748,N_1749);
nor U1834 (N_1834,N_1794,N_1740);
and U1835 (N_1835,N_1754,N_1762);
or U1836 (N_1836,N_1788,N_1753);
or U1837 (N_1837,N_1717,N_1705);
nor U1838 (N_1838,N_1707,N_1793);
nand U1839 (N_1839,N_1766,N_1787);
or U1840 (N_1840,N_1791,N_1764);
nor U1841 (N_1841,N_1779,N_1718);
and U1842 (N_1842,N_1776,N_1712);
or U1843 (N_1843,N_1704,N_1731);
and U1844 (N_1844,N_1741,N_1781);
nor U1845 (N_1845,N_1796,N_1783);
and U1846 (N_1846,N_1719,N_1745);
nand U1847 (N_1847,N_1723,N_1774);
xor U1848 (N_1848,N_1708,N_1789);
nand U1849 (N_1849,N_1743,N_1706);
and U1850 (N_1850,N_1745,N_1705);
or U1851 (N_1851,N_1754,N_1791);
and U1852 (N_1852,N_1777,N_1772);
and U1853 (N_1853,N_1794,N_1701);
or U1854 (N_1854,N_1714,N_1710);
nand U1855 (N_1855,N_1744,N_1754);
or U1856 (N_1856,N_1744,N_1715);
nand U1857 (N_1857,N_1713,N_1704);
or U1858 (N_1858,N_1768,N_1735);
or U1859 (N_1859,N_1782,N_1720);
and U1860 (N_1860,N_1787,N_1732);
and U1861 (N_1861,N_1744,N_1708);
or U1862 (N_1862,N_1782,N_1733);
or U1863 (N_1863,N_1732,N_1715);
xnor U1864 (N_1864,N_1766,N_1747);
or U1865 (N_1865,N_1713,N_1765);
and U1866 (N_1866,N_1794,N_1721);
or U1867 (N_1867,N_1750,N_1798);
and U1868 (N_1868,N_1797,N_1730);
or U1869 (N_1869,N_1707,N_1753);
or U1870 (N_1870,N_1766,N_1703);
and U1871 (N_1871,N_1790,N_1723);
nor U1872 (N_1872,N_1748,N_1792);
nand U1873 (N_1873,N_1741,N_1793);
nand U1874 (N_1874,N_1780,N_1754);
and U1875 (N_1875,N_1782,N_1771);
or U1876 (N_1876,N_1729,N_1762);
and U1877 (N_1877,N_1785,N_1776);
xnor U1878 (N_1878,N_1781,N_1709);
nand U1879 (N_1879,N_1749,N_1709);
nor U1880 (N_1880,N_1784,N_1781);
or U1881 (N_1881,N_1792,N_1737);
or U1882 (N_1882,N_1757,N_1775);
nor U1883 (N_1883,N_1747,N_1733);
nor U1884 (N_1884,N_1715,N_1735);
and U1885 (N_1885,N_1721,N_1760);
xnor U1886 (N_1886,N_1737,N_1741);
or U1887 (N_1887,N_1761,N_1793);
and U1888 (N_1888,N_1796,N_1790);
nor U1889 (N_1889,N_1762,N_1796);
xor U1890 (N_1890,N_1741,N_1768);
or U1891 (N_1891,N_1724,N_1703);
or U1892 (N_1892,N_1796,N_1776);
nand U1893 (N_1893,N_1728,N_1722);
or U1894 (N_1894,N_1734,N_1773);
or U1895 (N_1895,N_1715,N_1745);
nand U1896 (N_1896,N_1736,N_1755);
nor U1897 (N_1897,N_1798,N_1726);
or U1898 (N_1898,N_1740,N_1761);
nor U1899 (N_1899,N_1714,N_1744);
nand U1900 (N_1900,N_1846,N_1850);
nand U1901 (N_1901,N_1888,N_1808);
xor U1902 (N_1902,N_1891,N_1882);
nor U1903 (N_1903,N_1852,N_1832);
nor U1904 (N_1904,N_1813,N_1802);
xnor U1905 (N_1905,N_1805,N_1800);
nor U1906 (N_1906,N_1865,N_1856);
nor U1907 (N_1907,N_1874,N_1877);
nor U1908 (N_1908,N_1854,N_1836);
and U1909 (N_1909,N_1851,N_1849);
nand U1910 (N_1910,N_1870,N_1831);
nor U1911 (N_1911,N_1895,N_1830);
and U1912 (N_1912,N_1872,N_1869);
xnor U1913 (N_1913,N_1839,N_1890);
nand U1914 (N_1914,N_1892,N_1811);
or U1915 (N_1915,N_1864,N_1866);
nand U1916 (N_1916,N_1860,N_1819);
xor U1917 (N_1917,N_1889,N_1833);
or U1918 (N_1918,N_1816,N_1894);
or U1919 (N_1919,N_1875,N_1884);
nand U1920 (N_1920,N_1859,N_1809);
and U1921 (N_1921,N_1876,N_1871);
nand U1922 (N_1922,N_1825,N_1806);
nor U1923 (N_1923,N_1883,N_1807);
or U1924 (N_1924,N_1868,N_1834);
or U1925 (N_1925,N_1817,N_1867);
nand U1926 (N_1926,N_1887,N_1861);
nor U1927 (N_1927,N_1842,N_1899);
and U1928 (N_1928,N_1862,N_1801);
or U1929 (N_1929,N_1822,N_1835);
nor U1930 (N_1930,N_1873,N_1820);
nor U1931 (N_1931,N_1885,N_1844);
nand U1932 (N_1932,N_1810,N_1818);
nor U1933 (N_1933,N_1863,N_1898);
xor U1934 (N_1934,N_1853,N_1837);
nand U1935 (N_1935,N_1804,N_1840);
or U1936 (N_1936,N_1845,N_1824);
nand U1937 (N_1937,N_1843,N_1879);
or U1938 (N_1938,N_1803,N_1826);
nand U1939 (N_1939,N_1896,N_1880);
or U1940 (N_1940,N_1857,N_1838);
and U1941 (N_1941,N_1878,N_1841);
nor U1942 (N_1942,N_1855,N_1827);
nor U1943 (N_1943,N_1893,N_1848);
or U1944 (N_1944,N_1858,N_1823);
and U1945 (N_1945,N_1847,N_1821);
nor U1946 (N_1946,N_1829,N_1828);
nand U1947 (N_1947,N_1881,N_1897);
and U1948 (N_1948,N_1815,N_1814);
nor U1949 (N_1949,N_1812,N_1886);
nor U1950 (N_1950,N_1868,N_1899);
nand U1951 (N_1951,N_1849,N_1834);
and U1952 (N_1952,N_1800,N_1886);
nor U1953 (N_1953,N_1845,N_1875);
and U1954 (N_1954,N_1813,N_1862);
nand U1955 (N_1955,N_1829,N_1835);
or U1956 (N_1956,N_1866,N_1837);
and U1957 (N_1957,N_1876,N_1896);
nand U1958 (N_1958,N_1856,N_1839);
nor U1959 (N_1959,N_1809,N_1873);
nand U1960 (N_1960,N_1879,N_1884);
nand U1961 (N_1961,N_1844,N_1817);
nand U1962 (N_1962,N_1885,N_1856);
xor U1963 (N_1963,N_1883,N_1810);
xnor U1964 (N_1964,N_1844,N_1878);
xnor U1965 (N_1965,N_1831,N_1863);
nand U1966 (N_1966,N_1896,N_1858);
nand U1967 (N_1967,N_1881,N_1820);
and U1968 (N_1968,N_1811,N_1838);
nand U1969 (N_1969,N_1882,N_1835);
nor U1970 (N_1970,N_1869,N_1860);
nor U1971 (N_1971,N_1801,N_1876);
nand U1972 (N_1972,N_1847,N_1849);
nand U1973 (N_1973,N_1855,N_1873);
and U1974 (N_1974,N_1899,N_1800);
nor U1975 (N_1975,N_1860,N_1814);
nor U1976 (N_1976,N_1859,N_1880);
and U1977 (N_1977,N_1819,N_1837);
xor U1978 (N_1978,N_1866,N_1851);
nand U1979 (N_1979,N_1818,N_1802);
nor U1980 (N_1980,N_1837,N_1808);
nand U1981 (N_1981,N_1841,N_1837);
and U1982 (N_1982,N_1826,N_1823);
nand U1983 (N_1983,N_1845,N_1867);
and U1984 (N_1984,N_1817,N_1843);
nand U1985 (N_1985,N_1802,N_1810);
nor U1986 (N_1986,N_1866,N_1876);
or U1987 (N_1987,N_1847,N_1800);
nor U1988 (N_1988,N_1837,N_1870);
nor U1989 (N_1989,N_1867,N_1887);
nor U1990 (N_1990,N_1824,N_1876);
and U1991 (N_1991,N_1815,N_1825);
nand U1992 (N_1992,N_1867,N_1878);
or U1993 (N_1993,N_1810,N_1870);
or U1994 (N_1994,N_1827,N_1828);
and U1995 (N_1995,N_1869,N_1854);
or U1996 (N_1996,N_1877,N_1885);
nor U1997 (N_1997,N_1879,N_1822);
and U1998 (N_1998,N_1845,N_1858);
or U1999 (N_1999,N_1887,N_1812);
nor U2000 (N_2000,N_1918,N_1940);
nor U2001 (N_2001,N_1941,N_1960);
nor U2002 (N_2002,N_1905,N_1963);
and U2003 (N_2003,N_1924,N_1906);
and U2004 (N_2004,N_1931,N_1996);
xor U2005 (N_2005,N_1913,N_1966);
or U2006 (N_2006,N_1977,N_1955);
and U2007 (N_2007,N_1987,N_1968);
nor U2008 (N_2008,N_1912,N_1944);
and U2009 (N_2009,N_1970,N_1903);
nand U2010 (N_2010,N_1927,N_1971);
nor U2011 (N_2011,N_1943,N_1911);
and U2012 (N_2012,N_1929,N_1993);
and U2013 (N_2013,N_1997,N_1909);
xor U2014 (N_2014,N_1999,N_1974);
nand U2015 (N_2015,N_1956,N_1928);
nor U2016 (N_2016,N_1915,N_1964);
nor U2017 (N_2017,N_1989,N_1948);
nor U2018 (N_2018,N_1957,N_1933);
nand U2019 (N_2019,N_1979,N_1992);
xor U2020 (N_2020,N_1945,N_1949);
or U2021 (N_2021,N_1990,N_1923);
and U2022 (N_2022,N_1961,N_1901);
nand U2023 (N_2023,N_1969,N_1930);
and U2024 (N_2024,N_1902,N_1975);
nand U2025 (N_2025,N_1939,N_1926);
nor U2026 (N_2026,N_1998,N_1936);
and U2027 (N_2027,N_1934,N_1967);
and U2028 (N_2028,N_1986,N_1937);
nor U2029 (N_2029,N_1922,N_1976);
nand U2030 (N_2030,N_1947,N_1965);
nor U2031 (N_2031,N_1988,N_1921);
nand U2032 (N_2032,N_1958,N_1991);
or U2033 (N_2033,N_1914,N_1972);
or U2034 (N_2034,N_1916,N_1925);
and U2035 (N_2035,N_1982,N_1942);
nor U2036 (N_2036,N_1983,N_1932);
nand U2037 (N_2037,N_1907,N_1951);
nor U2038 (N_2038,N_1900,N_1946);
and U2039 (N_2039,N_1994,N_1953);
xor U2040 (N_2040,N_1910,N_1919);
nor U2041 (N_2041,N_1908,N_1973);
xor U2042 (N_2042,N_1980,N_1920);
nand U2043 (N_2043,N_1959,N_1995);
and U2044 (N_2044,N_1950,N_1917);
nand U2045 (N_2045,N_1952,N_1935);
and U2046 (N_2046,N_1978,N_1938);
nor U2047 (N_2047,N_1962,N_1981);
nor U2048 (N_2048,N_1904,N_1954);
xor U2049 (N_2049,N_1984,N_1985);
or U2050 (N_2050,N_1945,N_1913);
and U2051 (N_2051,N_1905,N_1974);
nand U2052 (N_2052,N_1959,N_1943);
xnor U2053 (N_2053,N_1958,N_1920);
nor U2054 (N_2054,N_1935,N_1951);
nand U2055 (N_2055,N_1960,N_1990);
or U2056 (N_2056,N_1915,N_1975);
or U2057 (N_2057,N_1904,N_1995);
or U2058 (N_2058,N_1987,N_1955);
nand U2059 (N_2059,N_1979,N_1937);
or U2060 (N_2060,N_1938,N_1912);
and U2061 (N_2061,N_1933,N_1912);
nor U2062 (N_2062,N_1939,N_1962);
nand U2063 (N_2063,N_1953,N_1918);
or U2064 (N_2064,N_1943,N_1985);
and U2065 (N_2065,N_1930,N_1912);
xnor U2066 (N_2066,N_1903,N_1976);
or U2067 (N_2067,N_1985,N_1993);
xor U2068 (N_2068,N_1966,N_1983);
or U2069 (N_2069,N_1901,N_1925);
nand U2070 (N_2070,N_1955,N_1953);
xnor U2071 (N_2071,N_1962,N_1989);
or U2072 (N_2072,N_1929,N_1904);
and U2073 (N_2073,N_1999,N_1994);
nor U2074 (N_2074,N_1987,N_1989);
nand U2075 (N_2075,N_1901,N_1971);
and U2076 (N_2076,N_1928,N_1954);
nand U2077 (N_2077,N_1969,N_1911);
nand U2078 (N_2078,N_1976,N_1920);
and U2079 (N_2079,N_1902,N_1990);
or U2080 (N_2080,N_1916,N_1918);
nor U2081 (N_2081,N_1931,N_1997);
nor U2082 (N_2082,N_1905,N_1915);
and U2083 (N_2083,N_1991,N_1972);
nand U2084 (N_2084,N_1919,N_1991);
nand U2085 (N_2085,N_1943,N_1989);
and U2086 (N_2086,N_1944,N_1954);
nor U2087 (N_2087,N_1903,N_1929);
nand U2088 (N_2088,N_1926,N_1961);
or U2089 (N_2089,N_1952,N_1965);
nor U2090 (N_2090,N_1981,N_1977);
or U2091 (N_2091,N_1905,N_1958);
and U2092 (N_2092,N_1923,N_1946);
and U2093 (N_2093,N_1997,N_1967);
nor U2094 (N_2094,N_1974,N_1956);
nand U2095 (N_2095,N_1993,N_1975);
nor U2096 (N_2096,N_1923,N_1962);
nand U2097 (N_2097,N_1918,N_1984);
and U2098 (N_2098,N_1921,N_1983);
nor U2099 (N_2099,N_1973,N_1972);
nand U2100 (N_2100,N_2045,N_2089);
and U2101 (N_2101,N_2014,N_2063);
or U2102 (N_2102,N_2093,N_2020);
nor U2103 (N_2103,N_2037,N_2058);
nand U2104 (N_2104,N_2092,N_2040);
nor U2105 (N_2105,N_2016,N_2090);
nand U2106 (N_2106,N_2022,N_2067);
nor U2107 (N_2107,N_2098,N_2082);
xor U2108 (N_2108,N_2047,N_2094);
nand U2109 (N_2109,N_2003,N_2019);
nor U2110 (N_2110,N_2002,N_2041);
nand U2111 (N_2111,N_2087,N_2055);
or U2112 (N_2112,N_2068,N_2065);
nor U2113 (N_2113,N_2005,N_2064);
xor U2114 (N_2114,N_2027,N_2039);
or U2115 (N_2115,N_2091,N_2008);
nor U2116 (N_2116,N_2096,N_2025);
nand U2117 (N_2117,N_2099,N_2084);
or U2118 (N_2118,N_2072,N_2073);
or U2119 (N_2119,N_2048,N_2053);
and U2120 (N_2120,N_2043,N_2017);
nor U2121 (N_2121,N_2034,N_2015);
and U2122 (N_2122,N_2062,N_2069);
and U2123 (N_2123,N_2028,N_2024);
xnor U2124 (N_2124,N_2086,N_2009);
nor U2125 (N_2125,N_2011,N_2071);
nor U2126 (N_2126,N_2032,N_2013);
and U2127 (N_2127,N_2049,N_2036);
and U2128 (N_2128,N_2054,N_2044);
and U2129 (N_2129,N_2075,N_2052);
or U2130 (N_2130,N_2083,N_2077);
or U2131 (N_2131,N_2095,N_2035);
nor U2132 (N_2132,N_2079,N_2018);
nor U2133 (N_2133,N_2010,N_2000);
and U2134 (N_2134,N_2080,N_2059);
nand U2135 (N_2135,N_2088,N_2031);
nand U2136 (N_2136,N_2076,N_2001);
and U2137 (N_2137,N_2085,N_2012);
or U2138 (N_2138,N_2097,N_2060);
xnor U2139 (N_2139,N_2021,N_2026);
or U2140 (N_2140,N_2050,N_2042);
nand U2141 (N_2141,N_2056,N_2081);
and U2142 (N_2142,N_2051,N_2046);
xnor U2143 (N_2143,N_2033,N_2038);
nor U2144 (N_2144,N_2030,N_2004);
or U2145 (N_2145,N_2061,N_2007);
nand U2146 (N_2146,N_2078,N_2074);
nand U2147 (N_2147,N_2023,N_2029);
nand U2148 (N_2148,N_2070,N_2057);
or U2149 (N_2149,N_2066,N_2006);
nor U2150 (N_2150,N_2027,N_2070);
nor U2151 (N_2151,N_2010,N_2075);
nand U2152 (N_2152,N_2041,N_2036);
nand U2153 (N_2153,N_2068,N_2097);
nand U2154 (N_2154,N_2072,N_2067);
and U2155 (N_2155,N_2075,N_2069);
xor U2156 (N_2156,N_2039,N_2004);
nand U2157 (N_2157,N_2067,N_2095);
and U2158 (N_2158,N_2085,N_2053);
nor U2159 (N_2159,N_2073,N_2063);
nor U2160 (N_2160,N_2069,N_2019);
nor U2161 (N_2161,N_2024,N_2005);
nor U2162 (N_2162,N_2049,N_2041);
or U2163 (N_2163,N_2098,N_2046);
nand U2164 (N_2164,N_2067,N_2017);
nor U2165 (N_2165,N_2068,N_2009);
nor U2166 (N_2166,N_2064,N_2018);
and U2167 (N_2167,N_2057,N_2072);
nor U2168 (N_2168,N_2053,N_2061);
nor U2169 (N_2169,N_2063,N_2018);
and U2170 (N_2170,N_2031,N_2007);
and U2171 (N_2171,N_2011,N_2089);
nand U2172 (N_2172,N_2086,N_2096);
and U2173 (N_2173,N_2005,N_2013);
or U2174 (N_2174,N_2048,N_2086);
nand U2175 (N_2175,N_2026,N_2082);
xor U2176 (N_2176,N_2065,N_2099);
or U2177 (N_2177,N_2077,N_2060);
or U2178 (N_2178,N_2068,N_2022);
and U2179 (N_2179,N_2082,N_2021);
nor U2180 (N_2180,N_2054,N_2052);
nor U2181 (N_2181,N_2024,N_2079);
and U2182 (N_2182,N_2023,N_2000);
nand U2183 (N_2183,N_2083,N_2072);
nand U2184 (N_2184,N_2036,N_2082);
or U2185 (N_2185,N_2075,N_2020);
nor U2186 (N_2186,N_2026,N_2024);
nand U2187 (N_2187,N_2072,N_2080);
nor U2188 (N_2188,N_2022,N_2086);
xnor U2189 (N_2189,N_2045,N_2047);
nor U2190 (N_2190,N_2016,N_2007);
nand U2191 (N_2191,N_2071,N_2016);
nor U2192 (N_2192,N_2025,N_2057);
or U2193 (N_2193,N_2019,N_2086);
nor U2194 (N_2194,N_2020,N_2050);
nor U2195 (N_2195,N_2083,N_2080);
xor U2196 (N_2196,N_2046,N_2031);
nor U2197 (N_2197,N_2008,N_2044);
and U2198 (N_2198,N_2099,N_2096);
and U2199 (N_2199,N_2032,N_2073);
nor U2200 (N_2200,N_2120,N_2124);
nor U2201 (N_2201,N_2110,N_2118);
or U2202 (N_2202,N_2139,N_2113);
nor U2203 (N_2203,N_2138,N_2122);
xnor U2204 (N_2204,N_2179,N_2132);
nor U2205 (N_2205,N_2128,N_2103);
xor U2206 (N_2206,N_2196,N_2147);
or U2207 (N_2207,N_2152,N_2130);
nor U2208 (N_2208,N_2192,N_2116);
and U2209 (N_2209,N_2143,N_2183);
or U2210 (N_2210,N_2127,N_2189);
or U2211 (N_2211,N_2117,N_2195);
and U2212 (N_2212,N_2159,N_2107);
and U2213 (N_2213,N_2169,N_2182);
or U2214 (N_2214,N_2174,N_2186);
nor U2215 (N_2215,N_2170,N_2141);
xnor U2216 (N_2216,N_2176,N_2163);
and U2217 (N_2217,N_2184,N_2115);
nand U2218 (N_2218,N_2160,N_2188);
xor U2219 (N_2219,N_2175,N_2190);
nor U2220 (N_2220,N_2173,N_2158);
and U2221 (N_2221,N_2112,N_2198);
nand U2222 (N_2222,N_2162,N_2166);
nand U2223 (N_2223,N_2149,N_2180);
nor U2224 (N_2224,N_2199,N_2114);
nand U2225 (N_2225,N_2131,N_2136);
or U2226 (N_2226,N_2108,N_2172);
or U2227 (N_2227,N_2171,N_2125);
xor U2228 (N_2228,N_2135,N_2105);
or U2229 (N_2229,N_2150,N_2104);
nor U2230 (N_2230,N_2164,N_2167);
xnor U2231 (N_2231,N_2185,N_2102);
and U2232 (N_2232,N_2161,N_2146);
nor U2233 (N_2233,N_2109,N_2177);
nor U2234 (N_2234,N_2168,N_2134);
and U2235 (N_2235,N_2126,N_2140);
and U2236 (N_2236,N_2151,N_2144);
nor U2237 (N_2237,N_2142,N_2148);
nand U2238 (N_2238,N_2121,N_2123);
and U2239 (N_2239,N_2153,N_2165);
nand U2240 (N_2240,N_2106,N_2157);
nor U2241 (N_2241,N_2181,N_2178);
and U2242 (N_2242,N_2187,N_2119);
xor U2243 (N_2243,N_2155,N_2145);
and U2244 (N_2244,N_2154,N_2193);
and U2245 (N_2245,N_2133,N_2100);
nor U2246 (N_2246,N_2111,N_2197);
nor U2247 (N_2247,N_2194,N_2129);
and U2248 (N_2248,N_2191,N_2156);
nand U2249 (N_2249,N_2101,N_2137);
or U2250 (N_2250,N_2154,N_2171);
or U2251 (N_2251,N_2110,N_2125);
and U2252 (N_2252,N_2199,N_2144);
nand U2253 (N_2253,N_2117,N_2138);
or U2254 (N_2254,N_2108,N_2113);
xor U2255 (N_2255,N_2159,N_2185);
xor U2256 (N_2256,N_2130,N_2199);
nor U2257 (N_2257,N_2138,N_2107);
nor U2258 (N_2258,N_2114,N_2118);
or U2259 (N_2259,N_2111,N_2145);
nor U2260 (N_2260,N_2112,N_2194);
nor U2261 (N_2261,N_2149,N_2165);
nor U2262 (N_2262,N_2160,N_2108);
or U2263 (N_2263,N_2117,N_2153);
nand U2264 (N_2264,N_2174,N_2193);
nand U2265 (N_2265,N_2161,N_2113);
or U2266 (N_2266,N_2111,N_2193);
and U2267 (N_2267,N_2191,N_2189);
or U2268 (N_2268,N_2161,N_2110);
and U2269 (N_2269,N_2181,N_2127);
and U2270 (N_2270,N_2187,N_2174);
nand U2271 (N_2271,N_2146,N_2118);
or U2272 (N_2272,N_2181,N_2123);
nand U2273 (N_2273,N_2157,N_2169);
and U2274 (N_2274,N_2105,N_2129);
xnor U2275 (N_2275,N_2106,N_2142);
or U2276 (N_2276,N_2113,N_2153);
or U2277 (N_2277,N_2110,N_2193);
nor U2278 (N_2278,N_2172,N_2104);
nor U2279 (N_2279,N_2109,N_2190);
nand U2280 (N_2280,N_2113,N_2182);
and U2281 (N_2281,N_2121,N_2118);
and U2282 (N_2282,N_2180,N_2148);
or U2283 (N_2283,N_2183,N_2159);
or U2284 (N_2284,N_2147,N_2117);
xnor U2285 (N_2285,N_2116,N_2174);
nand U2286 (N_2286,N_2103,N_2124);
xor U2287 (N_2287,N_2119,N_2137);
or U2288 (N_2288,N_2141,N_2181);
nand U2289 (N_2289,N_2126,N_2115);
xor U2290 (N_2290,N_2129,N_2158);
or U2291 (N_2291,N_2151,N_2156);
and U2292 (N_2292,N_2192,N_2121);
or U2293 (N_2293,N_2108,N_2158);
nor U2294 (N_2294,N_2157,N_2190);
or U2295 (N_2295,N_2182,N_2135);
or U2296 (N_2296,N_2182,N_2105);
nor U2297 (N_2297,N_2128,N_2150);
nand U2298 (N_2298,N_2130,N_2124);
and U2299 (N_2299,N_2144,N_2129);
nand U2300 (N_2300,N_2207,N_2222);
nand U2301 (N_2301,N_2276,N_2285);
nor U2302 (N_2302,N_2254,N_2288);
nand U2303 (N_2303,N_2266,N_2268);
and U2304 (N_2304,N_2220,N_2265);
or U2305 (N_2305,N_2280,N_2267);
and U2306 (N_2306,N_2241,N_2259);
xor U2307 (N_2307,N_2296,N_2275);
nor U2308 (N_2308,N_2235,N_2295);
nand U2309 (N_2309,N_2200,N_2224);
nor U2310 (N_2310,N_2273,N_2223);
or U2311 (N_2311,N_2233,N_2248);
or U2312 (N_2312,N_2283,N_2219);
nor U2313 (N_2313,N_2299,N_2215);
nor U2314 (N_2314,N_2221,N_2263);
nor U2315 (N_2315,N_2211,N_2246);
nor U2316 (N_2316,N_2230,N_2258);
nor U2317 (N_2317,N_2271,N_2245);
nor U2318 (N_2318,N_2239,N_2226);
and U2319 (N_2319,N_2294,N_2284);
nor U2320 (N_2320,N_2297,N_2286);
and U2321 (N_2321,N_2231,N_2278);
and U2322 (N_2322,N_2261,N_2210);
nand U2323 (N_2323,N_2217,N_2203);
nand U2324 (N_2324,N_2244,N_2234);
or U2325 (N_2325,N_2216,N_2214);
nand U2326 (N_2326,N_2201,N_2298);
nor U2327 (N_2327,N_2277,N_2237);
and U2328 (N_2328,N_2289,N_2243);
or U2329 (N_2329,N_2202,N_2208);
nand U2330 (N_2330,N_2251,N_2229);
or U2331 (N_2331,N_2240,N_2227);
nand U2332 (N_2332,N_2293,N_2290);
nor U2333 (N_2333,N_2272,N_2212);
or U2334 (N_2334,N_2206,N_2232);
xnor U2335 (N_2335,N_2205,N_2292);
nor U2336 (N_2336,N_2242,N_2252);
nor U2337 (N_2337,N_2247,N_2282);
or U2338 (N_2338,N_2253,N_2250);
and U2339 (N_2339,N_2238,N_2255);
nand U2340 (N_2340,N_2209,N_2236);
and U2341 (N_2341,N_2274,N_2225);
nand U2342 (N_2342,N_2287,N_2269);
nor U2343 (N_2343,N_2213,N_2204);
nor U2344 (N_2344,N_2279,N_2256);
and U2345 (N_2345,N_2257,N_2249);
nor U2346 (N_2346,N_2228,N_2218);
nor U2347 (N_2347,N_2270,N_2281);
nor U2348 (N_2348,N_2264,N_2260);
xnor U2349 (N_2349,N_2291,N_2262);
or U2350 (N_2350,N_2228,N_2204);
or U2351 (N_2351,N_2232,N_2259);
nand U2352 (N_2352,N_2263,N_2274);
nor U2353 (N_2353,N_2246,N_2225);
and U2354 (N_2354,N_2281,N_2265);
xor U2355 (N_2355,N_2276,N_2291);
nor U2356 (N_2356,N_2277,N_2204);
and U2357 (N_2357,N_2275,N_2288);
xor U2358 (N_2358,N_2224,N_2261);
or U2359 (N_2359,N_2248,N_2275);
nand U2360 (N_2360,N_2228,N_2268);
xnor U2361 (N_2361,N_2276,N_2219);
nor U2362 (N_2362,N_2201,N_2224);
nor U2363 (N_2363,N_2263,N_2278);
or U2364 (N_2364,N_2226,N_2281);
xnor U2365 (N_2365,N_2285,N_2242);
nor U2366 (N_2366,N_2238,N_2237);
and U2367 (N_2367,N_2250,N_2210);
nor U2368 (N_2368,N_2229,N_2231);
nor U2369 (N_2369,N_2246,N_2250);
or U2370 (N_2370,N_2222,N_2280);
and U2371 (N_2371,N_2289,N_2209);
xor U2372 (N_2372,N_2295,N_2225);
nor U2373 (N_2373,N_2203,N_2285);
nor U2374 (N_2374,N_2251,N_2243);
or U2375 (N_2375,N_2254,N_2236);
and U2376 (N_2376,N_2291,N_2281);
xnor U2377 (N_2377,N_2208,N_2277);
or U2378 (N_2378,N_2278,N_2277);
and U2379 (N_2379,N_2255,N_2230);
nand U2380 (N_2380,N_2277,N_2248);
and U2381 (N_2381,N_2208,N_2299);
or U2382 (N_2382,N_2290,N_2268);
or U2383 (N_2383,N_2286,N_2287);
or U2384 (N_2384,N_2290,N_2236);
nor U2385 (N_2385,N_2204,N_2224);
and U2386 (N_2386,N_2234,N_2205);
nand U2387 (N_2387,N_2207,N_2293);
nor U2388 (N_2388,N_2291,N_2296);
or U2389 (N_2389,N_2238,N_2207);
nor U2390 (N_2390,N_2273,N_2270);
or U2391 (N_2391,N_2280,N_2273);
and U2392 (N_2392,N_2206,N_2267);
and U2393 (N_2393,N_2216,N_2212);
nor U2394 (N_2394,N_2286,N_2255);
and U2395 (N_2395,N_2251,N_2257);
nand U2396 (N_2396,N_2256,N_2209);
or U2397 (N_2397,N_2264,N_2294);
nor U2398 (N_2398,N_2266,N_2258);
nand U2399 (N_2399,N_2262,N_2216);
and U2400 (N_2400,N_2318,N_2314);
nand U2401 (N_2401,N_2335,N_2385);
nand U2402 (N_2402,N_2388,N_2304);
and U2403 (N_2403,N_2396,N_2365);
nand U2404 (N_2404,N_2303,N_2333);
xnor U2405 (N_2405,N_2319,N_2370);
nand U2406 (N_2406,N_2366,N_2343);
nand U2407 (N_2407,N_2308,N_2315);
and U2408 (N_2408,N_2334,N_2306);
and U2409 (N_2409,N_2316,N_2320);
nand U2410 (N_2410,N_2307,N_2349);
nand U2411 (N_2411,N_2384,N_2331);
nor U2412 (N_2412,N_2324,N_2380);
xor U2413 (N_2413,N_2310,N_2311);
nand U2414 (N_2414,N_2375,N_2348);
or U2415 (N_2415,N_2329,N_2374);
or U2416 (N_2416,N_2382,N_2341);
or U2417 (N_2417,N_2389,N_2360);
nor U2418 (N_2418,N_2317,N_2362);
or U2419 (N_2419,N_2336,N_2340);
and U2420 (N_2420,N_2323,N_2359);
or U2421 (N_2421,N_2327,N_2300);
and U2422 (N_2422,N_2352,N_2390);
xor U2423 (N_2423,N_2368,N_2344);
nand U2424 (N_2424,N_2353,N_2332);
and U2425 (N_2425,N_2356,N_2325);
and U2426 (N_2426,N_2381,N_2364);
nand U2427 (N_2427,N_2376,N_2386);
nor U2428 (N_2428,N_2378,N_2337);
nand U2429 (N_2429,N_2342,N_2369);
xor U2430 (N_2430,N_2394,N_2367);
and U2431 (N_2431,N_2339,N_2346);
nand U2432 (N_2432,N_2350,N_2393);
nor U2433 (N_2433,N_2338,N_2379);
nand U2434 (N_2434,N_2395,N_2361);
and U2435 (N_2435,N_2321,N_2387);
and U2436 (N_2436,N_2330,N_2328);
or U2437 (N_2437,N_2312,N_2345);
nand U2438 (N_2438,N_2354,N_2358);
nand U2439 (N_2439,N_2377,N_2302);
nor U2440 (N_2440,N_2309,N_2398);
nor U2441 (N_2441,N_2392,N_2371);
nand U2442 (N_2442,N_2363,N_2397);
nand U2443 (N_2443,N_2383,N_2372);
nand U2444 (N_2444,N_2399,N_2313);
or U2445 (N_2445,N_2373,N_2305);
or U2446 (N_2446,N_2322,N_2347);
or U2447 (N_2447,N_2357,N_2301);
nand U2448 (N_2448,N_2351,N_2326);
or U2449 (N_2449,N_2391,N_2355);
and U2450 (N_2450,N_2380,N_2305);
or U2451 (N_2451,N_2325,N_2388);
nand U2452 (N_2452,N_2372,N_2380);
and U2453 (N_2453,N_2374,N_2354);
xnor U2454 (N_2454,N_2374,N_2305);
or U2455 (N_2455,N_2323,N_2391);
nor U2456 (N_2456,N_2322,N_2342);
and U2457 (N_2457,N_2322,N_2392);
nor U2458 (N_2458,N_2356,N_2387);
or U2459 (N_2459,N_2343,N_2373);
nor U2460 (N_2460,N_2366,N_2327);
and U2461 (N_2461,N_2364,N_2303);
or U2462 (N_2462,N_2302,N_2343);
nor U2463 (N_2463,N_2391,N_2379);
nand U2464 (N_2464,N_2377,N_2382);
nand U2465 (N_2465,N_2325,N_2360);
nand U2466 (N_2466,N_2372,N_2359);
and U2467 (N_2467,N_2329,N_2303);
or U2468 (N_2468,N_2320,N_2389);
or U2469 (N_2469,N_2344,N_2365);
xnor U2470 (N_2470,N_2306,N_2387);
nand U2471 (N_2471,N_2370,N_2389);
nor U2472 (N_2472,N_2329,N_2387);
or U2473 (N_2473,N_2322,N_2329);
nand U2474 (N_2474,N_2390,N_2384);
xor U2475 (N_2475,N_2366,N_2300);
nor U2476 (N_2476,N_2371,N_2386);
or U2477 (N_2477,N_2333,N_2321);
or U2478 (N_2478,N_2300,N_2325);
nor U2479 (N_2479,N_2342,N_2330);
nand U2480 (N_2480,N_2343,N_2321);
or U2481 (N_2481,N_2383,N_2322);
nand U2482 (N_2482,N_2360,N_2398);
nor U2483 (N_2483,N_2374,N_2369);
or U2484 (N_2484,N_2375,N_2327);
and U2485 (N_2485,N_2372,N_2355);
nand U2486 (N_2486,N_2324,N_2323);
or U2487 (N_2487,N_2311,N_2313);
and U2488 (N_2488,N_2369,N_2335);
or U2489 (N_2489,N_2399,N_2359);
nor U2490 (N_2490,N_2337,N_2395);
nand U2491 (N_2491,N_2389,N_2381);
and U2492 (N_2492,N_2311,N_2340);
and U2493 (N_2493,N_2369,N_2306);
and U2494 (N_2494,N_2383,N_2365);
or U2495 (N_2495,N_2381,N_2370);
and U2496 (N_2496,N_2397,N_2337);
or U2497 (N_2497,N_2346,N_2396);
nand U2498 (N_2498,N_2372,N_2367);
or U2499 (N_2499,N_2389,N_2399);
nor U2500 (N_2500,N_2414,N_2463);
or U2501 (N_2501,N_2456,N_2484);
and U2502 (N_2502,N_2477,N_2442);
xnor U2503 (N_2503,N_2438,N_2485);
nand U2504 (N_2504,N_2409,N_2492);
xnor U2505 (N_2505,N_2406,N_2482);
xor U2506 (N_2506,N_2432,N_2473);
or U2507 (N_2507,N_2417,N_2496);
and U2508 (N_2508,N_2451,N_2486);
nor U2509 (N_2509,N_2441,N_2468);
nand U2510 (N_2510,N_2470,N_2457);
nor U2511 (N_2511,N_2421,N_2418);
or U2512 (N_2512,N_2444,N_2412);
nand U2513 (N_2513,N_2474,N_2476);
and U2514 (N_2514,N_2454,N_2404);
xnor U2515 (N_2515,N_2460,N_2448);
nor U2516 (N_2516,N_2475,N_2471);
nand U2517 (N_2517,N_2447,N_2429);
nand U2518 (N_2518,N_2413,N_2439);
nor U2519 (N_2519,N_2462,N_2452);
nand U2520 (N_2520,N_2425,N_2420);
nor U2521 (N_2521,N_2489,N_2498);
and U2522 (N_2522,N_2416,N_2483);
and U2523 (N_2523,N_2400,N_2478);
nand U2524 (N_2524,N_2465,N_2495);
nand U2525 (N_2525,N_2437,N_2401);
or U2526 (N_2526,N_2466,N_2455);
and U2527 (N_2527,N_2459,N_2453);
nor U2528 (N_2528,N_2422,N_2405);
and U2529 (N_2529,N_2407,N_2433);
nand U2530 (N_2530,N_2446,N_2415);
or U2531 (N_2531,N_2411,N_2458);
or U2532 (N_2532,N_2402,N_2480);
nor U2533 (N_2533,N_2435,N_2490);
nand U2534 (N_2534,N_2450,N_2426);
or U2535 (N_2535,N_2461,N_2445);
and U2536 (N_2536,N_2467,N_2449);
and U2537 (N_2537,N_2487,N_2436);
and U2538 (N_2538,N_2464,N_2443);
nor U2539 (N_2539,N_2472,N_2493);
nand U2540 (N_2540,N_2403,N_2494);
and U2541 (N_2541,N_2430,N_2423);
or U2542 (N_2542,N_2427,N_2431);
xnor U2543 (N_2543,N_2499,N_2419);
nor U2544 (N_2544,N_2497,N_2424);
xnor U2545 (N_2545,N_2488,N_2440);
or U2546 (N_2546,N_2408,N_2479);
xor U2547 (N_2547,N_2434,N_2491);
and U2548 (N_2548,N_2481,N_2410);
nor U2549 (N_2549,N_2469,N_2428);
and U2550 (N_2550,N_2484,N_2467);
nor U2551 (N_2551,N_2494,N_2475);
xor U2552 (N_2552,N_2414,N_2458);
nand U2553 (N_2553,N_2490,N_2417);
nor U2554 (N_2554,N_2494,N_2451);
or U2555 (N_2555,N_2416,N_2459);
or U2556 (N_2556,N_2485,N_2427);
xor U2557 (N_2557,N_2435,N_2494);
or U2558 (N_2558,N_2486,N_2413);
or U2559 (N_2559,N_2441,N_2480);
nand U2560 (N_2560,N_2438,N_2431);
nand U2561 (N_2561,N_2454,N_2413);
or U2562 (N_2562,N_2435,N_2474);
nand U2563 (N_2563,N_2456,N_2466);
nor U2564 (N_2564,N_2462,N_2478);
xnor U2565 (N_2565,N_2472,N_2402);
or U2566 (N_2566,N_2484,N_2498);
nand U2567 (N_2567,N_2471,N_2486);
or U2568 (N_2568,N_2464,N_2420);
or U2569 (N_2569,N_2407,N_2430);
nor U2570 (N_2570,N_2447,N_2434);
nor U2571 (N_2571,N_2453,N_2444);
nor U2572 (N_2572,N_2462,N_2416);
nand U2573 (N_2573,N_2419,N_2459);
nand U2574 (N_2574,N_2428,N_2407);
nand U2575 (N_2575,N_2469,N_2466);
or U2576 (N_2576,N_2444,N_2476);
nand U2577 (N_2577,N_2447,N_2425);
nand U2578 (N_2578,N_2462,N_2409);
nor U2579 (N_2579,N_2436,N_2466);
nand U2580 (N_2580,N_2408,N_2456);
and U2581 (N_2581,N_2411,N_2432);
and U2582 (N_2582,N_2426,N_2466);
and U2583 (N_2583,N_2444,N_2446);
and U2584 (N_2584,N_2419,N_2454);
nand U2585 (N_2585,N_2400,N_2426);
and U2586 (N_2586,N_2446,N_2422);
and U2587 (N_2587,N_2489,N_2434);
or U2588 (N_2588,N_2474,N_2475);
nor U2589 (N_2589,N_2458,N_2475);
nor U2590 (N_2590,N_2428,N_2405);
nand U2591 (N_2591,N_2453,N_2475);
or U2592 (N_2592,N_2478,N_2422);
or U2593 (N_2593,N_2408,N_2483);
nor U2594 (N_2594,N_2460,N_2459);
and U2595 (N_2595,N_2414,N_2455);
or U2596 (N_2596,N_2469,N_2403);
and U2597 (N_2597,N_2419,N_2430);
nand U2598 (N_2598,N_2468,N_2499);
nand U2599 (N_2599,N_2459,N_2433);
or U2600 (N_2600,N_2550,N_2510);
or U2601 (N_2601,N_2521,N_2551);
nor U2602 (N_2602,N_2505,N_2508);
and U2603 (N_2603,N_2559,N_2592);
or U2604 (N_2604,N_2527,N_2585);
and U2605 (N_2605,N_2553,N_2542);
nand U2606 (N_2606,N_2504,N_2588);
nand U2607 (N_2607,N_2534,N_2586);
nand U2608 (N_2608,N_2572,N_2537);
nor U2609 (N_2609,N_2528,N_2578);
nand U2610 (N_2610,N_2532,N_2591);
and U2611 (N_2611,N_2566,N_2580);
nor U2612 (N_2612,N_2570,N_2563);
or U2613 (N_2613,N_2520,N_2565);
xor U2614 (N_2614,N_2573,N_2546);
or U2615 (N_2615,N_2576,N_2581);
nor U2616 (N_2616,N_2577,N_2543);
nand U2617 (N_2617,N_2541,N_2547);
or U2618 (N_2618,N_2568,N_2582);
or U2619 (N_2619,N_2552,N_2539);
nor U2620 (N_2620,N_2587,N_2530);
or U2621 (N_2621,N_2522,N_2555);
nand U2622 (N_2622,N_2519,N_2562);
and U2623 (N_2623,N_2569,N_2525);
nor U2624 (N_2624,N_2526,N_2513);
nand U2625 (N_2625,N_2590,N_2560);
and U2626 (N_2626,N_2583,N_2571);
or U2627 (N_2627,N_2558,N_2524);
xor U2628 (N_2628,N_2556,N_2506);
nor U2629 (N_2629,N_2548,N_2517);
xor U2630 (N_2630,N_2595,N_2564);
or U2631 (N_2631,N_2557,N_2575);
xor U2632 (N_2632,N_2502,N_2597);
xor U2633 (N_2633,N_2561,N_2516);
nor U2634 (N_2634,N_2507,N_2523);
and U2635 (N_2635,N_2594,N_2518);
nor U2636 (N_2636,N_2574,N_2598);
nand U2637 (N_2637,N_2540,N_2593);
xor U2638 (N_2638,N_2584,N_2589);
nor U2639 (N_2639,N_2544,N_2531);
nand U2640 (N_2640,N_2533,N_2503);
and U2641 (N_2641,N_2567,N_2500);
nor U2642 (N_2642,N_2596,N_2554);
nor U2643 (N_2643,N_2514,N_2515);
nor U2644 (N_2644,N_2511,N_2529);
and U2645 (N_2645,N_2579,N_2536);
nor U2646 (N_2646,N_2512,N_2509);
or U2647 (N_2647,N_2599,N_2501);
nor U2648 (N_2648,N_2535,N_2538);
nor U2649 (N_2649,N_2549,N_2545);
nand U2650 (N_2650,N_2571,N_2531);
and U2651 (N_2651,N_2571,N_2552);
nand U2652 (N_2652,N_2577,N_2592);
and U2653 (N_2653,N_2527,N_2545);
nand U2654 (N_2654,N_2515,N_2578);
and U2655 (N_2655,N_2503,N_2564);
or U2656 (N_2656,N_2559,N_2546);
or U2657 (N_2657,N_2581,N_2587);
or U2658 (N_2658,N_2525,N_2531);
nand U2659 (N_2659,N_2510,N_2572);
nand U2660 (N_2660,N_2537,N_2529);
nor U2661 (N_2661,N_2522,N_2590);
and U2662 (N_2662,N_2563,N_2584);
or U2663 (N_2663,N_2543,N_2522);
xnor U2664 (N_2664,N_2551,N_2567);
nand U2665 (N_2665,N_2544,N_2557);
or U2666 (N_2666,N_2517,N_2537);
and U2667 (N_2667,N_2559,N_2541);
and U2668 (N_2668,N_2558,N_2505);
or U2669 (N_2669,N_2575,N_2599);
or U2670 (N_2670,N_2534,N_2569);
nor U2671 (N_2671,N_2593,N_2546);
and U2672 (N_2672,N_2562,N_2587);
nand U2673 (N_2673,N_2534,N_2547);
nand U2674 (N_2674,N_2519,N_2553);
nor U2675 (N_2675,N_2536,N_2520);
and U2676 (N_2676,N_2517,N_2561);
nor U2677 (N_2677,N_2579,N_2586);
xor U2678 (N_2678,N_2598,N_2591);
and U2679 (N_2679,N_2513,N_2500);
nand U2680 (N_2680,N_2555,N_2516);
and U2681 (N_2681,N_2512,N_2567);
nor U2682 (N_2682,N_2586,N_2529);
nor U2683 (N_2683,N_2523,N_2542);
and U2684 (N_2684,N_2599,N_2531);
nor U2685 (N_2685,N_2545,N_2565);
or U2686 (N_2686,N_2597,N_2516);
and U2687 (N_2687,N_2591,N_2540);
nor U2688 (N_2688,N_2524,N_2530);
xor U2689 (N_2689,N_2580,N_2570);
and U2690 (N_2690,N_2510,N_2529);
nand U2691 (N_2691,N_2572,N_2511);
nand U2692 (N_2692,N_2594,N_2516);
nor U2693 (N_2693,N_2551,N_2571);
nand U2694 (N_2694,N_2507,N_2563);
nand U2695 (N_2695,N_2584,N_2524);
nor U2696 (N_2696,N_2560,N_2585);
xor U2697 (N_2697,N_2579,N_2521);
nand U2698 (N_2698,N_2514,N_2564);
or U2699 (N_2699,N_2580,N_2527);
or U2700 (N_2700,N_2627,N_2643);
and U2701 (N_2701,N_2667,N_2637);
nor U2702 (N_2702,N_2658,N_2616);
nand U2703 (N_2703,N_2623,N_2673);
nand U2704 (N_2704,N_2654,N_2657);
or U2705 (N_2705,N_2612,N_2625);
nor U2706 (N_2706,N_2691,N_2610);
nor U2707 (N_2707,N_2652,N_2651);
xnor U2708 (N_2708,N_2694,N_2699);
nand U2709 (N_2709,N_2622,N_2642);
xnor U2710 (N_2710,N_2656,N_2671);
nand U2711 (N_2711,N_2698,N_2603);
nor U2712 (N_2712,N_2647,N_2630);
nor U2713 (N_2713,N_2655,N_2607);
nor U2714 (N_2714,N_2693,N_2649);
nor U2715 (N_2715,N_2681,N_2688);
xor U2716 (N_2716,N_2646,N_2665);
or U2717 (N_2717,N_2633,N_2608);
or U2718 (N_2718,N_2660,N_2617);
nor U2719 (N_2719,N_2620,N_2650);
or U2720 (N_2720,N_2605,N_2600);
nor U2721 (N_2721,N_2690,N_2653);
and U2722 (N_2722,N_2614,N_2645);
or U2723 (N_2723,N_2664,N_2663);
nand U2724 (N_2724,N_2641,N_2666);
and U2725 (N_2725,N_2695,N_2661);
xor U2726 (N_2726,N_2634,N_2618);
nor U2727 (N_2727,N_2672,N_2697);
nor U2728 (N_2728,N_2636,N_2674);
nand U2729 (N_2729,N_2684,N_2639);
xor U2730 (N_2730,N_2680,N_2629);
nor U2731 (N_2731,N_2662,N_2683);
nand U2732 (N_2732,N_2602,N_2644);
nor U2733 (N_2733,N_2668,N_2613);
xnor U2734 (N_2734,N_2669,N_2685);
or U2735 (N_2735,N_2621,N_2632);
or U2736 (N_2736,N_2615,N_2659);
and U2737 (N_2737,N_2675,N_2676);
or U2738 (N_2738,N_2611,N_2638);
nand U2739 (N_2739,N_2635,N_2686);
nand U2740 (N_2740,N_2601,N_2640);
nand U2741 (N_2741,N_2609,N_2624);
nor U2742 (N_2742,N_2682,N_2689);
nor U2743 (N_2743,N_2678,N_2679);
nor U2744 (N_2744,N_2619,N_2677);
xnor U2745 (N_2745,N_2670,N_2687);
or U2746 (N_2746,N_2628,N_2696);
nor U2747 (N_2747,N_2692,N_2604);
nand U2748 (N_2748,N_2648,N_2606);
and U2749 (N_2749,N_2626,N_2631);
nor U2750 (N_2750,N_2601,N_2660);
and U2751 (N_2751,N_2666,N_2688);
or U2752 (N_2752,N_2648,N_2686);
nand U2753 (N_2753,N_2675,N_2696);
and U2754 (N_2754,N_2604,N_2685);
or U2755 (N_2755,N_2678,N_2676);
nor U2756 (N_2756,N_2643,N_2635);
nor U2757 (N_2757,N_2670,N_2686);
and U2758 (N_2758,N_2681,N_2651);
and U2759 (N_2759,N_2603,N_2601);
and U2760 (N_2760,N_2658,N_2697);
and U2761 (N_2761,N_2606,N_2619);
nand U2762 (N_2762,N_2619,N_2622);
nor U2763 (N_2763,N_2667,N_2689);
or U2764 (N_2764,N_2696,N_2689);
nand U2765 (N_2765,N_2661,N_2620);
or U2766 (N_2766,N_2657,N_2693);
or U2767 (N_2767,N_2605,N_2649);
xnor U2768 (N_2768,N_2637,N_2604);
nand U2769 (N_2769,N_2620,N_2603);
nor U2770 (N_2770,N_2699,N_2638);
and U2771 (N_2771,N_2679,N_2612);
xnor U2772 (N_2772,N_2676,N_2604);
and U2773 (N_2773,N_2655,N_2603);
or U2774 (N_2774,N_2614,N_2640);
nand U2775 (N_2775,N_2639,N_2655);
or U2776 (N_2776,N_2675,N_2603);
or U2777 (N_2777,N_2641,N_2678);
and U2778 (N_2778,N_2637,N_2646);
xnor U2779 (N_2779,N_2674,N_2668);
nand U2780 (N_2780,N_2646,N_2644);
nand U2781 (N_2781,N_2601,N_2696);
and U2782 (N_2782,N_2602,N_2691);
nand U2783 (N_2783,N_2659,N_2647);
or U2784 (N_2784,N_2684,N_2617);
nor U2785 (N_2785,N_2627,N_2663);
nor U2786 (N_2786,N_2686,N_2697);
or U2787 (N_2787,N_2653,N_2642);
and U2788 (N_2788,N_2639,N_2666);
nand U2789 (N_2789,N_2674,N_2692);
nand U2790 (N_2790,N_2664,N_2693);
or U2791 (N_2791,N_2630,N_2658);
nor U2792 (N_2792,N_2600,N_2662);
or U2793 (N_2793,N_2653,N_2665);
or U2794 (N_2794,N_2669,N_2670);
and U2795 (N_2795,N_2675,N_2664);
nor U2796 (N_2796,N_2604,N_2622);
and U2797 (N_2797,N_2674,N_2603);
nand U2798 (N_2798,N_2665,N_2696);
or U2799 (N_2799,N_2615,N_2688);
and U2800 (N_2800,N_2767,N_2717);
and U2801 (N_2801,N_2758,N_2775);
nor U2802 (N_2802,N_2740,N_2795);
nand U2803 (N_2803,N_2751,N_2777);
nand U2804 (N_2804,N_2716,N_2742);
nor U2805 (N_2805,N_2786,N_2756);
nor U2806 (N_2806,N_2715,N_2711);
and U2807 (N_2807,N_2744,N_2754);
and U2808 (N_2808,N_2797,N_2760);
and U2809 (N_2809,N_2766,N_2738);
nand U2810 (N_2810,N_2737,N_2710);
nand U2811 (N_2811,N_2781,N_2774);
nor U2812 (N_2812,N_2707,N_2743);
or U2813 (N_2813,N_2727,N_2759);
or U2814 (N_2814,N_2761,N_2732);
or U2815 (N_2815,N_2701,N_2793);
xor U2816 (N_2816,N_2763,N_2718);
or U2817 (N_2817,N_2784,N_2752);
and U2818 (N_2818,N_2757,N_2705);
and U2819 (N_2819,N_2798,N_2724);
nor U2820 (N_2820,N_2748,N_2782);
nand U2821 (N_2821,N_2764,N_2787);
nand U2822 (N_2822,N_2791,N_2762);
and U2823 (N_2823,N_2722,N_2792);
nand U2824 (N_2824,N_2729,N_2713);
and U2825 (N_2825,N_2773,N_2772);
or U2826 (N_2826,N_2703,N_2725);
and U2827 (N_2827,N_2736,N_2750);
nor U2828 (N_2828,N_2770,N_2789);
or U2829 (N_2829,N_2768,N_2720);
or U2830 (N_2830,N_2745,N_2790);
or U2831 (N_2831,N_2721,N_2712);
and U2832 (N_2832,N_2753,N_2733);
nand U2833 (N_2833,N_2778,N_2700);
and U2834 (N_2834,N_2785,N_2788);
nand U2835 (N_2835,N_2739,N_2771);
nor U2836 (N_2836,N_2747,N_2765);
nor U2837 (N_2837,N_2796,N_2769);
nand U2838 (N_2838,N_2728,N_2749);
or U2839 (N_2839,N_2799,N_2708);
nand U2840 (N_2840,N_2780,N_2779);
nand U2841 (N_2841,N_2730,N_2702);
or U2842 (N_2842,N_2709,N_2746);
nand U2843 (N_2843,N_2776,N_2723);
and U2844 (N_2844,N_2755,N_2706);
and U2845 (N_2845,N_2734,N_2726);
or U2846 (N_2846,N_2783,N_2719);
and U2847 (N_2847,N_2735,N_2714);
nor U2848 (N_2848,N_2794,N_2731);
xor U2849 (N_2849,N_2741,N_2704);
or U2850 (N_2850,N_2728,N_2784);
or U2851 (N_2851,N_2781,N_2788);
and U2852 (N_2852,N_2754,N_2791);
nor U2853 (N_2853,N_2702,N_2714);
or U2854 (N_2854,N_2792,N_2744);
nor U2855 (N_2855,N_2776,N_2751);
nor U2856 (N_2856,N_2785,N_2740);
nand U2857 (N_2857,N_2738,N_2713);
nand U2858 (N_2858,N_2736,N_2795);
nand U2859 (N_2859,N_2703,N_2795);
nand U2860 (N_2860,N_2706,N_2777);
nand U2861 (N_2861,N_2786,N_2724);
or U2862 (N_2862,N_2759,N_2751);
and U2863 (N_2863,N_2755,N_2736);
or U2864 (N_2864,N_2773,N_2735);
nor U2865 (N_2865,N_2736,N_2788);
or U2866 (N_2866,N_2700,N_2772);
and U2867 (N_2867,N_2718,N_2741);
and U2868 (N_2868,N_2790,N_2775);
or U2869 (N_2869,N_2778,N_2719);
nor U2870 (N_2870,N_2791,N_2720);
nor U2871 (N_2871,N_2761,N_2723);
and U2872 (N_2872,N_2747,N_2746);
or U2873 (N_2873,N_2748,N_2710);
nor U2874 (N_2874,N_2758,N_2721);
nor U2875 (N_2875,N_2774,N_2722);
nor U2876 (N_2876,N_2744,N_2702);
nor U2877 (N_2877,N_2740,N_2762);
and U2878 (N_2878,N_2785,N_2775);
nor U2879 (N_2879,N_2753,N_2736);
xor U2880 (N_2880,N_2750,N_2738);
nand U2881 (N_2881,N_2749,N_2715);
nor U2882 (N_2882,N_2750,N_2708);
nand U2883 (N_2883,N_2736,N_2790);
or U2884 (N_2884,N_2703,N_2704);
nand U2885 (N_2885,N_2708,N_2756);
nor U2886 (N_2886,N_2796,N_2790);
nand U2887 (N_2887,N_2767,N_2727);
or U2888 (N_2888,N_2780,N_2723);
or U2889 (N_2889,N_2713,N_2723);
and U2890 (N_2890,N_2740,N_2708);
nand U2891 (N_2891,N_2714,N_2783);
and U2892 (N_2892,N_2749,N_2706);
or U2893 (N_2893,N_2790,N_2751);
and U2894 (N_2894,N_2796,N_2760);
nor U2895 (N_2895,N_2788,N_2726);
nor U2896 (N_2896,N_2795,N_2793);
nor U2897 (N_2897,N_2736,N_2784);
and U2898 (N_2898,N_2789,N_2711);
or U2899 (N_2899,N_2765,N_2756);
nand U2900 (N_2900,N_2847,N_2887);
or U2901 (N_2901,N_2839,N_2806);
or U2902 (N_2902,N_2859,N_2836);
xor U2903 (N_2903,N_2830,N_2844);
or U2904 (N_2904,N_2814,N_2853);
and U2905 (N_2905,N_2868,N_2898);
nand U2906 (N_2906,N_2819,N_2831);
nor U2907 (N_2907,N_2840,N_2801);
or U2908 (N_2908,N_2871,N_2896);
or U2909 (N_2909,N_2807,N_2870);
nor U2910 (N_2910,N_2826,N_2852);
nand U2911 (N_2911,N_2829,N_2845);
nor U2912 (N_2912,N_2842,N_2862);
nand U2913 (N_2913,N_2854,N_2874);
xnor U2914 (N_2914,N_2849,N_2835);
and U2915 (N_2915,N_2821,N_2841);
xnor U2916 (N_2916,N_2810,N_2805);
or U2917 (N_2917,N_2869,N_2877);
or U2918 (N_2918,N_2891,N_2864);
nor U2919 (N_2919,N_2822,N_2851);
nor U2920 (N_2920,N_2800,N_2817);
nor U2921 (N_2921,N_2856,N_2889);
xor U2922 (N_2922,N_2855,N_2812);
xor U2923 (N_2923,N_2897,N_2813);
and U2924 (N_2924,N_2833,N_2886);
and U2925 (N_2925,N_2825,N_2808);
xnor U2926 (N_2926,N_2828,N_2820);
xnor U2927 (N_2927,N_2878,N_2892);
nor U2928 (N_2928,N_2837,N_2866);
xnor U2929 (N_2929,N_2895,N_2809);
or U2930 (N_2930,N_2843,N_2893);
or U2931 (N_2931,N_2823,N_2883);
nor U2932 (N_2932,N_2899,N_2818);
nand U2933 (N_2933,N_2861,N_2850);
xor U2934 (N_2934,N_2827,N_2882);
and U2935 (N_2935,N_2875,N_2824);
nand U2936 (N_2936,N_2848,N_2888);
and U2937 (N_2937,N_2816,N_2894);
nand U2938 (N_2938,N_2802,N_2857);
nand U2939 (N_2939,N_2846,N_2834);
xnor U2940 (N_2940,N_2884,N_2815);
nor U2941 (N_2941,N_2890,N_2873);
nor U2942 (N_2942,N_2860,N_2858);
nor U2943 (N_2943,N_2880,N_2867);
or U2944 (N_2944,N_2863,N_2832);
and U2945 (N_2945,N_2872,N_2811);
nor U2946 (N_2946,N_2876,N_2804);
or U2947 (N_2947,N_2838,N_2885);
or U2948 (N_2948,N_2881,N_2865);
and U2949 (N_2949,N_2879,N_2803);
nor U2950 (N_2950,N_2880,N_2838);
nor U2951 (N_2951,N_2875,N_2846);
xnor U2952 (N_2952,N_2893,N_2852);
nor U2953 (N_2953,N_2890,N_2819);
nor U2954 (N_2954,N_2827,N_2820);
and U2955 (N_2955,N_2859,N_2806);
and U2956 (N_2956,N_2803,N_2832);
nor U2957 (N_2957,N_2870,N_2820);
nor U2958 (N_2958,N_2801,N_2887);
nor U2959 (N_2959,N_2850,N_2897);
nor U2960 (N_2960,N_2877,N_2862);
nor U2961 (N_2961,N_2884,N_2857);
or U2962 (N_2962,N_2840,N_2855);
and U2963 (N_2963,N_2834,N_2890);
nor U2964 (N_2964,N_2851,N_2860);
or U2965 (N_2965,N_2884,N_2863);
nor U2966 (N_2966,N_2887,N_2820);
and U2967 (N_2967,N_2855,N_2888);
nor U2968 (N_2968,N_2880,N_2858);
nand U2969 (N_2969,N_2843,N_2834);
or U2970 (N_2970,N_2832,N_2805);
and U2971 (N_2971,N_2842,N_2829);
nand U2972 (N_2972,N_2822,N_2843);
or U2973 (N_2973,N_2806,N_2899);
nor U2974 (N_2974,N_2826,N_2810);
nor U2975 (N_2975,N_2897,N_2835);
nor U2976 (N_2976,N_2865,N_2827);
nand U2977 (N_2977,N_2866,N_2803);
nand U2978 (N_2978,N_2895,N_2815);
nor U2979 (N_2979,N_2811,N_2834);
or U2980 (N_2980,N_2892,N_2832);
and U2981 (N_2981,N_2837,N_2812);
or U2982 (N_2982,N_2898,N_2830);
nand U2983 (N_2983,N_2867,N_2801);
and U2984 (N_2984,N_2892,N_2880);
or U2985 (N_2985,N_2888,N_2826);
xnor U2986 (N_2986,N_2812,N_2844);
and U2987 (N_2987,N_2860,N_2875);
and U2988 (N_2988,N_2849,N_2898);
nor U2989 (N_2989,N_2827,N_2840);
nand U2990 (N_2990,N_2858,N_2803);
and U2991 (N_2991,N_2847,N_2836);
nor U2992 (N_2992,N_2854,N_2896);
nor U2993 (N_2993,N_2867,N_2816);
and U2994 (N_2994,N_2857,N_2845);
and U2995 (N_2995,N_2854,N_2837);
and U2996 (N_2996,N_2894,N_2840);
xnor U2997 (N_2997,N_2879,N_2874);
nor U2998 (N_2998,N_2845,N_2869);
or U2999 (N_2999,N_2842,N_2811);
and U3000 (N_3000,N_2954,N_2981);
and U3001 (N_3001,N_2985,N_2995);
nand U3002 (N_3002,N_2941,N_2977);
nor U3003 (N_3003,N_2996,N_2933);
or U3004 (N_3004,N_2936,N_2973);
and U3005 (N_3005,N_2929,N_2901);
and U3006 (N_3006,N_2984,N_2914);
or U3007 (N_3007,N_2945,N_2902);
and U3008 (N_3008,N_2918,N_2969);
nor U3009 (N_3009,N_2956,N_2906);
or U3010 (N_3010,N_2938,N_2932);
and U3011 (N_3011,N_2990,N_2967);
nor U3012 (N_3012,N_2998,N_2907);
nor U3013 (N_3013,N_2993,N_2950);
nor U3014 (N_3014,N_2909,N_2982);
or U3015 (N_3015,N_2952,N_2957);
nand U3016 (N_3016,N_2944,N_2949);
xor U3017 (N_3017,N_2935,N_2904);
or U3018 (N_3018,N_2999,N_2928);
nand U3019 (N_3019,N_2912,N_2910);
nor U3020 (N_3020,N_2961,N_2927);
or U3021 (N_3021,N_2926,N_2921);
or U3022 (N_3022,N_2923,N_2979);
nor U3023 (N_3023,N_2931,N_2917);
and U3024 (N_3024,N_2900,N_2948);
nand U3025 (N_3025,N_2966,N_2964);
nor U3026 (N_3026,N_2937,N_2913);
or U3027 (N_3027,N_2908,N_2953);
nor U3028 (N_3028,N_2991,N_2962);
nor U3029 (N_3029,N_2997,N_2925);
and U3030 (N_3030,N_2986,N_2922);
nor U3031 (N_3031,N_2916,N_2911);
nor U3032 (N_3032,N_2942,N_2974);
or U3033 (N_3033,N_2943,N_2920);
xor U3034 (N_3034,N_2975,N_2980);
nand U3035 (N_3035,N_2946,N_2987);
nand U3036 (N_3036,N_2905,N_2989);
nor U3037 (N_3037,N_2971,N_2992);
nor U3038 (N_3038,N_2958,N_2903);
xnor U3039 (N_3039,N_2919,N_2970);
and U3040 (N_3040,N_2978,N_2960);
xnor U3041 (N_3041,N_2940,N_2968);
nand U3042 (N_3042,N_2947,N_2924);
nand U3043 (N_3043,N_2934,N_2915);
nand U3044 (N_3044,N_2951,N_2983);
nor U3045 (N_3045,N_2994,N_2939);
nand U3046 (N_3046,N_2972,N_2965);
xor U3047 (N_3047,N_2930,N_2959);
nand U3048 (N_3048,N_2963,N_2955);
xnor U3049 (N_3049,N_2988,N_2976);
nand U3050 (N_3050,N_2947,N_2932);
xor U3051 (N_3051,N_2944,N_2931);
xor U3052 (N_3052,N_2961,N_2932);
xor U3053 (N_3053,N_2908,N_2927);
nand U3054 (N_3054,N_2907,N_2914);
xnor U3055 (N_3055,N_2942,N_2984);
or U3056 (N_3056,N_2948,N_2930);
or U3057 (N_3057,N_2983,N_2917);
nand U3058 (N_3058,N_2923,N_2927);
or U3059 (N_3059,N_2901,N_2919);
nor U3060 (N_3060,N_2929,N_2965);
or U3061 (N_3061,N_2978,N_2981);
and U3062 (N_3062,N_2923,N_2921);
or U3063 (N_3063,N_2915,N_2976);
nand U3064 (N_3064,N_2959,N_2975);
nor U3065 (N_3065,N_2926,N_2936);
nand U3066 (N_3066,N_2907,N_2947);
nor U3067 (N_3067,N_2907,N_2979);
nand U3068 (N_3068,N_2979,N_2940);
or U3069 (N_3069,N_2974,N_2931);
or U3070 (N_3070,N_2956,N_2948);
nand U3071 (N_3071,N_2915,N_2952);
or U3072 (N_3072,N_2930,N_2996);
or U3073 (N_3073,N_2916,N_2908);
nor U3074 (N_3074,N_2940,N_2973);
nor U3075 (N_3075,N_2963,N_2931);
and U3076 (N_3076,N_2956,N_2934);
or U3077 (N_3077,N_2903,N_2912);
and U3078 (N_3078,N_2926,N_2990);
nor U3079 (N_3079,N_2900,N_2927);
nand U3080 (N_3080,N_2967,N_2907);
and U3081 (N_3081,N_2965,N_2987);
nand U3082 (N_3082,N_2996,N_2928);
nor U3083 (N_3083,N_2948,N_2963);
or U3084 (N_3084,N_2996,N_2914);
or U3085 (N_3085,N_2938,N_2948);
xor U3086 (N_3086,N_2999,N_2908);
and U3087 (N_3087,N_2963,N_2944);
or U3088 (N_3088,N_2921,N_2912);
nor U3089 (N_3089,N_2917,N_2916);
and U3090 (N_3090,N_2950,N_2926);
nor U3091 (N_3091,N_2917,N_2944);
or U3092 (N_3092,N_2932,N_2935);
nor U3093 (N_3093,N_2934,N_2977);
or U3094 (N_3094,N_2939,N_2980);
nor U3095 (N_3095,N_2902,N_2997);
xor U3096 (N_3096,N_2990,N_2995);
or U3097 (N_3097,N_2907,N_2924);
nor U3098 (N_3098,N_2959,N_2949);
nand U3099 (N_3099,N_2920,N_2945);
and U3100 (N_3100,N_3093,N_3010);
or U3101 (N_3101,N_3038,N_3047);
xnor U3102 (N_3102,N_3067,N_3063);
and U3103 (N_3103,N_3044,N_3088);
nor U3104 (N_3104,N_3004,N_3042);
and U3105 (N_3105,N_3094,N_3021);
xnor U3106 (N_3106,N_3076,N_3008);
or U3107 (N_3107,N_3041,N_3073);
nand U3108 (N_3108,N_3015,N_3046);
and U3109 (N_3109,N_3043,N_3027);
nor U3110 (N_3110,N_3053,N_3003);
or U3111 (N_3111,N_3040,N_3002);
xor U3112 (N_3112,N_3070,N_3035);
xnor U3113 (N_3113,N_3066,N_3024);
nand U3114 (N_3114,N_3095,N_3017);
and U3115 (N_3115,N_3086,N_3006);
nor U3116 (N_3116,N_3092,N_3048);
nand U3117 (N_3117,N_3029,N_3049);
nor U3118 (N_3118,N_3037,N_3036);
and U3119 (N_3119,N_3026,N_3080);
and U3120 (N_3120,N_3075,N_3059);
nor U3121 (N_3121,N_3025,N_3009);
and U3122 (N_3122,N_3085,N_3082);
nand U3123 (N_3123,N_3060,N_3081);
or U3124 (N_3124,N_3089,N_3055);
nor U3125 (N_3125,N_3018,N_3062);
nor U3126 (N_3126,N_3012,N_3030);
nand U3127 (N_3127,N_3083,N_3077);
nor U3128 (N_3128,N_3034,N_3084);
or U3129 (N_3129,N_3098,N_3064);
nor U3130 (N_3130,N_3051,N_3045);
and U3131 (N_3131,N_3031,N_3022);
or U3132 (N_3132,N_3028,N_3005);
nor U3133 (N_3133,N_3078,N_3011);
xnor U3134 (N_3134,N_3019,N_3068);
nor U3135 (N_3135,N_3023,N_3032);
nor U3136 (N_3136,N_3016,N_3061);
xor U3137 (N_3137,N_3013,N_3039);
xor U3138 (N_3138,N_3054,N_3071);
or U3139 (N_3139,N_3079,N_3096);
nand U3140 (N_3140,N_3014,N_3099);
and U3141 (N_3141,N_3097,N_3091);
nor U3142 (N_3142,N_3065,N_3052);
nand U3143 (N_3143,N_3072,N_3057);
xnor U3144 (N_3144,N_3069,N_3020);
and U3145 (N_3145,N_3001,N_3007);
nand U3146 (N_3146,N_3000,N_3058);
nor U3147 (N_3147,N_3050,N_3074);
nand U3148 (N_3148,N_3090,N_3087);
xnor U3149 (N_3149,N_3056,N_3033);
and U3150 (N_3150,N_3088,N_3072);
nand U3151 (N_3151,N_3021,N_3064);
nand U3152 (N_3152,N_3038,N_3084);
nor U3153 (N_3153,N_3065,N_3018);
xnor U3154 (N_3154,N_3074,N_3003);
or U3155 (N_3155,N_3076,N_3051);
nor U3156 (N_3156,N_3089,N_3028);
nand U3157 (N_3157,N_3087,N_3026);
xor U3158 (N_3158,N_3030,N_3078);
nor U3159 (N_3159,N_3090,N_3073);
nor U3160 (N_3160,N_3041,N_3083);
nor U3161 (N_3161,N_3036,N_3083);
nand U3162 (N_3162,N_3002,N_3045);
xor U3163 (N_3163,N_3079,N_3010);
nor U3164 (N_3164,N_3006,N_3018);
nand U3165 (N_3165,N_3005,N_3027);
xnor U3166 (N_3166,N_3001,N_3086);
and U3167 (N_3167,N_3003,N_3031);
nand U3168 (N_3168,N_3007,N_3040);
nand U3169 (N_3169,N_3011,N_3009);
nand U3170 (N_3170,N_3039,N_3054);
or U3171 (N_3171,N_3082,N_3060);
nor U3172 (N_3172,N_3037,N_3073);
nor U3173 (N_3173,N_3095,N_3004);
xor U3174 (N_3174,N_3076,N_3065);
nor U3175 (N_3175,N_3032,N_3062);
xor U3176 (N_3176,N_3022,N_3068);
and U3177 (N_3177,N_3077,N_3053);
nand U3178 (N_3178,N_3031,N_3099);
nor U3179 (N_3179,N_3043,N_3096);
or U3180 (N_3180,N_3081,N_3034);
nor U3181 (N_3181,N_3033,N_3059);
nor U3182 (N_3182,N_3032,N_3016);
or U3183 (N_3183,N_3046,N_3036);
xor U3184 (N_3184,N_3090,N_3049);
and U3185 (N_3185,N_3006,N_3080);
nor U3186 (N_3186,N_3053,N_3009);
nor U3187 (N_3187,N_3079,N_3087);
nor U3188 (N_3188,N_3052,N_3037);
nand U3189 (N_3189,N_3093,N_3054);
or U3190 (N_3190,N_3032,N_3096);
and U3191 (N_3191,N_3047,N_3050);
xor U3192 (N_3192,N_3077,N_3024);
nand U3193 (N_3193,N_3091,N_3067);
and U3194 (N_3194,N_3015,N_3032);
or U3195 (N_3195,N_3091,N_3031);
nand U3196 (N_3196,N_3093,N_3002);
nor U3197 (N_3197,N_3032,N_3034);
nand U3198 (N_3198,N_3012,N_3073);
nand U3199 (N_3199,N_3025,N_3074);
nand U3200 (N_3200,N_3114,N_3104);
or U3201 (N_3201,N_3158,N_3191);
nand U3202 (N_3202,N_3127,N_3129);
nor U3203 (N_3203,N_3109,N_3132);
or U3204 (N_3204,N_3195,N_3184);
nand U3205 (N_3205,N_3121,N_3101);
nor U3206 (N_3206,N_3159,N_3181);
and U3207 (N_3207,N_3128,N_3143);
nand U3208 (N_3208,N_3162,N_3166);
nor U3209 (N_3209,N_3170,N_3113);
or U3210 (N_3210,N_3171,N_3185);
or U3211 (N_3211,N_3173,N_3139);
and U3212 (N_3212,N_3150,N_3163);
nand U3213 (N_3213,N_3177,N_3118);
nor U3214 (N_3214,N_3136,N_3178);
nor U3215 (N_3215,N_3183,N_3146);
and U3216 (N_3216,N_3103,N_3154);
or U3217 (N_3217,N_3110,N_3172);
and U3218 (N_3218,N_3176,N_3182);
nor U3219 (N_3219,N_3165,N_3156);
nand U3220 (N_3220,N_3179,N_3115);
xnor U3221 (N_3221,N_3174,N_3125);
xor U3222 (N_3222,N_3120,N_3100);
nor U3223 (N_3223,N_3168,N_3144);
nor U3224 (N_3224,N_3186,N_3188);
nor U3225 (N_3225,N_3119,N_3108);
or U3226 (N_3226,N_3193,N_3106);
xor U3227 (N_3227,N_3138,N_3187);
or U3228 (N_3228,N_3197,N_3135);
and U3229 (N_3229,N_3142,N_3123);
nand U3230 (N_3230,N_3112,N_3134);
nor U3231 (N_3231,N_3105,N_3133);
and U3232 (N_3232,N_3180,N_3116);
nand U3233 (N_3233,N_3157,N_3199);
nor U3234 (N_3234,N_3155,N_3153);
nand U3235 (N_3235,N_3169,N_3117);
and U3236 (N_3236,N_3152,N_3198);
xnor U3237 (N_3237,N_3122,N_3164);
and U3238 (N_3238,N_3148,N_3145);
nand U3239 (N_3239,N_3111,N_3137);
xor U3240 (N_3240,N_3192,N_3160);
and U3241 (N_3241,N_3107,N_3190);
or U3242 (N_3242,N_3161,N_3149);
nand U3243 (N_3243,N_3140,N_3189);
or U3244 (N_3244,N_3126,N_3130);
nor U3245 (N_3245,N_3141,N_3102);
nor U3246 (N_3246,N_3194,N_3131);
nor U3247 (N_3247,N_3175,N_3147);
nor U3248 (N_3248,N_3167,N_3124);
xor U3249 (N_3249,N_3196,N_3151);
or U3250 (N_3250,N_3122,N_3100);
nand U3251 (N_3251,N_3152,N_3171);
nand U3252 (N_3252,N_3127,N_3113);
nand U3253 (N_3253,N_3122,N_3114);
or U3254 (N_3254,N_3189,N_3196);
or U3255 (N_3255,N_3182,N_3110);
nor U3256 (N_3256,N_3163,N_3164);
nor U3257 (N_3257,N_3182,N_3166);
nor U3258 (N_3258,N_3186,N_3109);
xor U3259 (N_3259,N_3173,N_3181);
nand U3260 (N_3260,N_3104,N_3127);
nor U3261 (N_3261,N_3149,N_3163);
and U3262 (N_3262,N_3139,N_3185);
or U3263 (N_3263,N_3154,N_3158);
nand U3264 (N_3264,N_3145,N_3189);
nor U3265 (N_3265,N_3132,N_3149);
or U3266 (N_3266,N_3198,N_3164);
or U3267 (N_3267,N_3121,N_3132);
or U3268 (N_3268,N_3156,N_3113);
nor U3269 (N_3269,N_3156,N_3119);
and U3270 (N_3270,N_3199,N_3159);
nor U3271 (N_3271,N_3132,N_3193);
and U3272 (N_3272,N_3169,N_3136);
or U3273 (N_3273,N_3133,N_3138);
nor U3274 (N_3274,N_3174,N_3188);
xnor U3275 (N_3275,N_3118,N_3136);
nand U3276 (N_3276,N_3198,N_3184);
and U3277 (N_3277,N_3128,N_3164);
or U3278 (N_3278,N_3184,N_3178);
nor U3279 (N_3279,N_3167,N_3126);
nand U3280 (N_3280,N_3154,N_3155);
nor U3281 (N_3281,N_3114,N_3128);
and U3282 (N_3282,N_3159,N_3152);
nor U3283 (N_3283,N_3194,N_3182);
or U3284 (N_3284,N_3179,N_3103);
or U3285 (N_3285,N_3105,N_3112);
nand U3286 (N_3286,N_3122,N_3101);
nand U3287 (N_3287,N_3133,N_3151);
xor U3288 (N_3288,N_3193,N_3177);
and U3289 (N_3289,N_3109,N_3104);
and U3290 (N_3290,N_3177,N_3147);
nand U3291 (N_3291,N_3126,N_3174);
or U3292 (N_3292,N_3109,N_3144);
nand U3293 (N_3293,N_3131,N_3175);
nor U3294 (N_3294,N_3134,N_3118);
nor U3295 (N_3295,N_3174,N_3132);
xnor U3296 (N_3296,N_3158,N_3159);
nand U3297 (N_3297,N_3111,N_3139);
nand U3298 (N_3298,N_3163,N_3135);
nor U3299 (N_3299,N_3113,N_3102);
xnor U3300 (N_3300,N_3248,N_3262);
nor U3301 (N_3301,N_3232,N_3268);
and U3302 (N_3302,N_3256,N_3225);
and U3303 (N_3303,N_3274,N_3251);
or U3304 (N_3304,N_3255,N_3236);
xor U3305 (N_3305,N_3276,N_3279);
nand U3306 (N_3306,N_3213,N_3241);
nor U3307 (N_3307,N_3209,N_3263);
nor U3308 (N_3308,N_3240,N_3283);
nand U3309 (N_3309,N_3281,N_3222);
and U3310 (N_3310,N_3289,N_3264);
nor U3311 (N_3311,N_3245,N_3260);
nand U3312 (N_3312,N_3219,N_3290);
nand U3313 (N_3313,N_3200,N_3214);
or U3314 (N_3314,N_3216,N_3261);
and U3315 (N_3315,N_3299,N_3297);
or U3316 (N_3316,N_3269,N_3285);
or U3317 (N_3317,N_3202,N_3286);
or U3318 (N_3318,N_3284,N_3293);
nor U3319 (N_3319,N_3266,N_3238);
nand U3320 (N_3320,N_3224,N_3246);
and U3321 (N_3321,N_3250,N_3296);
nor U3322 (N_3322,N_3234,N_3204);
nand U3323 (N_3323,N_3244,N_3207);
nor U3324 (N_3324,N_3217,N_3282);
or U3325 (N_3325,N_3298,N_3231);
or U3326 (N_3326,N_3242,N_3203);
nor U3327 (N_3327,N_3277,N_3257);
and U3328 (N_3328,N_3218,N_3210);
nand U3329 (N_3329,N_3239,N_3223);
and U3330 (N_3330,N_3237,N_3273);
nand U3331 (N_3331,N_3221,N_3278);
xnor U3332 (N_3332,N_3220,N_3292);
nor U3333 (N_3333,N_3212,N_3275);
xnor U3334 (N_3334,N_3253,N_3252);
and U3335 (N_3335,N_3291,N_3267);
nand U3336 (N_3336,N_3249,N_3254);
and U3337 (N_3337,N_3258,N_3227);
nand U3338 (N_3338,N_3265,N_3259);
and U3339 (N_3339,N_3235,N_3271);
and U3340 (N_3340,N_3228,N_3288);
or U3341 (N_3341,N_3233,N_3211);
or U3342 (N_3342,N_3280,N_3295);
or U3343 (N_3343,N_3205,N_3229);
or U3344 (N_3344,N_3226,N_3247);
nand U3345 (N_3345,N_3230,N_3243);
or U3346 (N_3346,N_3294,N_3272);
or U3347 (N_3347,N_3215,N_3206);
and U3348 (N_3348,N_3270,N_3208);
and U3349 (N_3349,N_3201,N_3287);
or U3350 (N_3350,N_3243,N_3285);
and U3351 (N_3351,N_3236,N_3230);
xnor U3352 (N_3352,N_3200,N_3230);
and U3353 (N_3353,N_3293,N_3236);
nand U3354 (N_3354,N_3239,N_3287);
nor U3355 (N_3355,N_3282,N_3219);
or U3356 (N_3356,N_3286,N_3221);
and U3357 (N_3357,N_3288,N_3252);
nor U3358 (N_3358,N_3222,N_3284);
nor U3359 (N_3359,N_3200,N_3298);
nor U3360 (N_3360,N_3202,N_3218);
nor U3361 (N_3361,N_3279,N_3202);
or U3362 (N_3362,N_3279,N_3224);
and U3363 (N_3363,N_3252,N_3243);
or U3364 (N_3364,N_3234,N_3201);
or U3365 (N_3365,N_3226,N_3205);
or U3366 (N_3366,N_3267,N_3251);
nor U3367 (N_3367,N_3213,N_3224);
and U3368 (N_3368,N_3282,N_3290);
and U3369 (N_3369,N_3224,N_3264);
nand U3370 (N_3370,N_3208,N_3274);
and U3371 (N_3371,N_3218,N_3294);
nand U3372 (N_3372,N_3206,N_3258);
and U3373 (N_3373,N_3241,N_3208);
xnor U3374 (N_3374,N_3207,N_3271);
nand U3375 (N_3375,N_3256,N_3251);
and U3376 (N_3376,N_3244,N_3228);
and U3377 (N_3377,N_3213,N_3222);
and U3378 (N_3378,N_3225,N_3240);
or U3379 (N_3379,N_3215,N_3225);
or U3380 (N_3380,N_3223,N_3284);
nand U3381 (N_3381,N_3230,N_3212);
and U3382 (N_3382,N_3249,N_3264);
or U3383 (N_3383,N_3208,N_3255);
or U3384 (N_3384,N_3204,N_3220);
or U3385 (N_3385,N_3228,N_3250);
nor U3386 (N_3386,N_3297,N_3228);
and U3387 (N_3387,N_3265,N_3253);
xor U3388 (N_3388,N_3229,N_3260);
or U3389 (N_3389,N_3272,N_3207);
or U3390 (N_3390,N_3251,N_3284);
nor U3391 (N_3391,N_3256,N_3205);
and U3392 (N_3392,N_3244,N_3290);
nand U3393 (N_3393,N_3279,N_3285);
or U3394 (N_3394,N_3272,N_3236);
and U3395 (N_3395,N_3213,N_3239);
or U3396 (N_3396,N_3276,N_3206);
nor U3397 (N_3397,N_3211,N_3272);
or U3398 (N_3398,N_3229,N_3228);
nand U3399 (N_3399,N_3234,N_3206);
and U3400 (N_3400,N_3310,N_3378);
nand U3401 (N_3401,N_3307,N_3368);
and U3402 (N_3402,N_3332,N_3399);
xor U3403 (N_3403,N_3380,N_3382);
nor U3404 (N_3404,N_3358,N_3355);
nor U3405 (N_3405,N_3329,N_3347);
nor U3406 (N_3406,N_3353,N_3372);
nor U3407 (N_3407,N_3331,N_3344);
nor U3408 (N_3408,N_3324,N_3337);
and U3409 (N_3409,N_3311,N_3320);
nand U3410 (N_3410,N_3393,N_3377);
nand U3411 (N_3411,N_3392,N_3300);
and U3412 (N_3412,N_3376,N_3314);
xnor U3413 (N_3413,N_3370,N_3304);
nor U3414 (N_3414,N_3305,N_3356);
nand U3415 (N_3415,N_3365,N_3342);
nand U3416 (N_3416,N_3387,N_3306);
and U3417 (N_3417,N_3395,N_3374);
nand U3418 (N_3418,N_3317,N_3302);
and U3419 (N_3419,N_3367,N_3398);
or U3420 (N_3420,N_3383,N_3309);
nand U3421 (N_3421,N_3318,N_3352);
nor U3422 (N_3422,N_3321,N_3328);
and U3423 (N_3423,N_3346,N_3364);
xnor U3424 (N_3424,N_3389,N_3359);
nor U3425 (N_3425,N_3322,N_3361);
or U3426 (N_3426,N_3384,N_3351);
nand U3427 (N_3427,N_3391,N_3357);
nand U3428 (N_3428,N_3362,N_3330);
xor U3429 (N_3429,N_3394,N_3336);
xnor U3430 (N_3430,N_3396,N_3375);
and U3431 (N_3431,N_3341,N_3326);
and U3432 (N_3432,N_3363,N_3301);
nand U3433 (N_3433,N_3366,N_3348);
and U3434 (N_3434,N_3315,N_3319);
nor U3435 (N_3435,N_3390,N_3333);
nor U3436 (N_3436,N_3354,N_3312);
or U3437 (N_3437,N_3325,N_3339);
xnor U3438 (N_3438,N_3388,N_3381);
and U3439 (N_3439,N_3316,N_3369);
and U3440 (N_3440,N_3308,N_3340);
nand U3441 (N_3441,N_3385,N_3313);
nor U3442 (N_3442,N_3350,N_3327);
and U3443 (N_3443,N_3360,N_3303);
or U3444 (N_3444,N_3397,N_3349);
nor U3445 (N_3445,N_3334,N_3343);
xor U3446 (N_3446,N_3345,N_3338);
nor U3447 (N_3447,N_3371,N_3373);
xnor U3448 (N_3448,N_3386,N_3323);
xor U3449 (N_3449,N_3335,N_3379);
or U3450 (N_3450,N_3358,N_3369);
nor U3451 (N_3451,N_3324,N_3333);
nand U3452 (N_3452,N_3397,N_3323);
nand U3453 (N_3453,N_3365,N_3331);
nor U3454 (N_3454,N_3360,N_3395);
and U3455 (N_3455,N_3396,N_3319);
nand U3456 (N_3456,N_3335,N_3386);
nand U3457 (N_3457,N_3397,N_3347);
or U3458 (N_3458,N_3357,N_3310);
or U3459 (N_3459,N_3374,N_3385);
nand U3460 (N_3460,N_3359,N_3330);
or U3461 (N_3461,N_3347,N_3353);
or U3462 (N_3462,N_3357,N_3389);
nand U3463 (N_3463,N_3366,N_3379);
nor U3464 (N_3464,N_3359,N_3351);
nand U3465 (N_3465,N_3328,N_3346);
xnor U3466 (N_3466,N_3344,N_3367);
and U3467 (N_3467,N_3317,N_3334);
nand U3468 (N_3468,N_3366,N_3383);
nand U3469 (N_3469,N_3335,N_3307);
and U3470 (N_3470,N_3382,N_3363);
and U3471 (N_3471,N_3338,N_3308);
and U3472 (N_3472,N_3325,N_3347);
and U3473 (N_3473,N_3315,N_3329);
and U3474 (N_3474,N_3322,N_3399);
nand U3475 (N_3475,N_3306,N_3346);
and U3476 (N_3476,N_3368,N_3348);
xnor U3477 (N_3477,N_3397,N_3332);
nor U3478 (N_3478,N_3353,N_3396);
xor U3479 (N_3479,N_3321,N_3304);
nand U3480 (N_3480,N_3304,N_3311);
xor U3481 (N_3481,N_3364,N_3384);
nor U3482 (N_3482,N_3309,N_3384);
and U3483 (N_3483,N_3384,N_3322);
or U3484 (N_3484,N_3371,N_3358);
nor U3485 (N_3485,N_3371,N_3338);
nand U3486 (N_3486,N_3381,N_3393);
or U3487 (N_3487,N_3310,N_3307);
nand U3488 (N_3488,N_3353,N_3316);
and U3489 (N_3489,N_3347,N_3309);
and U3490 (N_3490,N_3369,N_3310);
nand U3491 (N_3491,N_3369,N_3327);
and U3492 (N_3492,N_3303,N_3353);
nor U3493 (N_3493,N_3377,N_3341);
nor U3494 (N_3494,N_3373,N_3368);
or U3495 (N_3495,N_3381,N_3382);
and U3496 (N_3496,N_3331,N_3370);
or U3497 (N_3497,N_3348,N_3372);
nor U3498 (N_3498,N_3338,N_3303);
nand U3499 (N_3499,N_3392,N_3381);
nand U3500 (N_3500,N_3433,N_3477);
or U3501 (N_3501,N_3485,N_3404);
nand U3502 (N_3502,N_3416,N_3479);
nor U3503 (N_3503,N_3467,N_3463);
nor U3504 (N_3504,N_3417,N_3461);
nand U3505 (N_3505,N_3401,N_3465);
or U3506 (N_3506,N_3495,N_3452);
xor U3507 (N_3507,N_3439,N_3437);
nand U3508 (N_3508,N_3444,N_3457);
and U3509 (N_3509,N_3453,N_3454);
and U3510 (N_3510,N_3450,N_3470);
nor U3511 (N_3511,N_3409,N_3432);
nand U3512 (N_3512,N_3425,N_3490);
nand U3513 (N_3513,N_3423,N_3498);
and U3514 (N_3514,N_3446,N_3471);
or U3515 (N_3515,N_3405,N_3411);
or U3516 (N_3516,N_3483,N_3431);
or U3517 (N_3517,N_3484,N_3402);
xnor U3518 (N_3518,N_3419,N_3447);
and U3519 (N_3519,N_3445,N_3403);
or U3520 (N_3520,N_3418,N_3458);
nor U3521 (N_3521,N_3455,N_3487);
xor U3522 (N_3522,N_3436,N_3459);
or U3523 (N_3523,N_3468,N_3469);
and U3524 (N_3524,N_3466,N_3499);
nor U3525 (N_3525,N_3426,N_3497);
nor U3526 (N_3526,N_3456,N_3472);
and U3527 (N_3527,N_3481,N_3413);
and U3528 (N_3528,N_3440,N_3407);
or U3529 (N_3529,N_3427,N_3422);
nand U3530 (N_3530,N_3493,N_3428);
and U3531 (N_3531,N_3434,N_3435);
or U3532 (N_3532,N_3415,N_3489);
or U3533 (N_3533,N_3410,N_3462);
or U3534 (N_3534,N_3443,N_3442);
nor U3535 (N_3535,N_3430,N_3438);
or U3536 (N_3536,N_3414,N_3475);
nor U3537 (N_3537,N_3486,N_3476);
nor U3538 (N_3538,N_3400,N_3491);
and U3539 (N_3539,N_3412,N_3406);
nor U3540 (N_3540,N_3496,N_3488);
nor U3541 (N_3541,N_3429,N_3482);
xnor U3542 (N_3542,N_3421,N_3420);
and U3543 (N_3543,N_3474,N_3464);
nand U3544 (N_3544,N_3460,N_3478);
nand U3545 (N_3545,N_3494,N_3449);
nor U3546 (N_3546,N_3448,N_3424);
or U3547 (N_3547,N_3408,N_3480);
nor U3548 (N_3548,N_3492,N_3441);
nand U3549 (N_3549,N_3473,N_3451);
nand U3550 (N_3550,N_3416,N_3419);
or U3551 (N_3551,N_3468,N_3413);
nand U3552 (N_3552,N_3449,N_3428);
nor U3553 (N_3553,N_3493,N_3469);
and U3554 (N_3554,N_3422,N_3408);
nor U3555 (N_3555,N_3499,N_3416);
xor U3556 (N_3556,N_3470,N_3455);
xor U3557 (N_3557,N_3487,N_3469);
and U3558 (N_3558,N_3494,N_3410);
or U3559 (N_3559,N_3425,N_3486);
or U3560 (N_3560,N_3470,N_3413);
nand U3561 (N_3561,N_3471,N_3461);
nor U3562 (N_3562,N_3467,N_3433);
xnor U3563 (N_3563,N_3487,N_3479);
nor U3564 (N_3564,N_3479,N_3418);
nand U3565 (N_3565,N_3494,N_3477);
or U3566 (N_3566,N_3496,N_3487);
nor U3567 (N_3567,N_3444,N_3492);
or U3568 (N_3568,N_3495,N_3467);
and U3569 (N_3569,N_3470,N_3460);
and U3570 (N_3570,N_3471,N_3449);
xnor U3571 (N_3571,N_3452,N_3469);
xnor U3572 (N_3572,N_3470,N_3420);
nor U3573 (N_3573,N_3432,N_3441);
or U3574 (N_3574,N_3489,N_3476);
xor U3575 (N_3575,N_3475,N_3471);
nand U3576 (N_3576,N_3474,N_3452);
nand U3577 (N_3577,N_3440,N_3461);
and U3578 (N_3578,N_3407,N_3433);
nand U3579 (N_3579,N_3414,N_3401);
nand U3580 (N_3580,N_3433,N_3430);
nor U3581 (N_3581,N_3458,N_3435);
and U3582 (N_3582,N_3467,N_3488);
or U3583 (N_3583,N_3432,N_3423);
or U3584 (N_3584,N_3485,N_3458);
nor U3585 (N_3585,N_3442,N_3456);
or U3586 (N_3586,N_3406,N_3457);
and U3587 (N_3587,N_3485,N_3410);
and U3588 (N_3588,N_3416,N_3441);
nor U3589 (N_3589,N_3415,N_3452);
nand U3590 (N_3590,N_3417,N_3473);
or U3591 (N_3591,N_3438,N_3428);
nand U3592 (N_3592,N_3454,N_3413);
nand U3593 (N_3593,N_3435,N_3467);
nand U3594 (N_3594,N_3493,N_3484);
nand U3595 (N_3595,N_3434,N_3433);
or U3596 (N_3596,N_3400,N_3423);
and U3597 (N_3597,N_3482,N_3497);
or U3598 (N_3598,N_3497,N_3473);
nor U3599 (N_3599,N_3437,N_3409);
and U3600 (N_3600,N_3583,N_3529);
nand U3601 (N_3601,N_3533,N_3582);
nand U3602 (N_3602,N_3563,N_3560);
or U3603 (N_3603,N_3561,N_3573);
nor U3604 (N_3604,N_3523,N_3562);
nand U3605 (N_3605,N_3521,N_3531);
nand U3606 (N_3606,N_3559,N_3537);
and U3607 (N_3607,N_3592,N_3506);
nor U3608 (N_3608,N_3545,N_3536);
or U3609 (N_3609,N_3596,N_3558);
and U3610 (N_3610,N_3519,N_3598);
and U3611 (N_3611,N_3579,N_3593);
nor U3612 (N_3612,N_3597,N_3591);
or U3613 (N_3613,N_3526,N_3547);
or U3614 (N_3614,N_3549,N_3567);
nor U3615 (N_3615,N_3522,N_3511);
xor U3616 (N_3616,N_3564,N_3508);
and U3617 (N_3617,N_3552,N_3502);
nand U3618 (N_3618,N_3530,N_3541);
or U3619 (N_3619,N_3557,N_3574);
nand U3620 (N_3620,N_3590,N_3586);
nor U3621 (N_3621,N_3527,N_3539);
or U3622 (N_3622,N_3551,N_3548);
and U3623 (N_3623,N_3504,N_3515);
xor U3624 (N_3624,N_3575,N_3538);
and U3625 (N_3625,N_3584,N_3507);
or U3626 (N_3626,N_3569,N_3518);
xor U3627 (N_3627,N_3570,N_3503);
or U3628 (N_3628,N_3513,N_3553);
and U3629 (N_3629,N_3525,N_3544);
xnor U3630 (N_3630,N_3524,N_3578);
and U3631 (N_3631,N_3514,N_3568);
and U3632 (N_3632,N_3572,N_3500);
nand U3633 (N_3633,N_3554,N_3516);
nand U3634 (N_3634,N_3520,N_3534);
nand U3635 (N_3635,N_3577,N_3543);
or U3636 (N_3636,N_3599,N_3587);
nand U3637 (N_3637,N_3580,N_3501);
xor U3638 (N_3638,N_3550,N_3546);
nor U3639 (N_3639,N_3576,N_3505);
nor U3640 (N_3640,N_3542,N_3509);
or U3641 (N_3641,N_3566,N_3589);
or U3642 (N_3642,N_3517,N_3571);
xnor U3643 (N_3643,N_3588,N_3512);
nand U3644 (N_3644,N_3532,N_3594);
and U3645 (N_3645,N_3581,N_3595);
and U3646 (N_3646,N_3510,N_3556);
and U3647 (N_3647,N_3528,N_3585);
xnor U3648 (N_3648,N_3555,N_3540);
nand U3649 (N_3649,N_3535,N_3565);
nor U3650 (N_3650,N_3557,N_3561);
xor U3651 (N_3651,N_3535,N_3590);
nand U3652 (N_3652,N_3520,N_3547);
xor U3653 (N_3653,N_3544,N_3505);
and U3654 (N_3654,N_3546,N_3527);
and U3655 (N_3655,N_3548,N_3517);
and U3656 (N_3656,N_3542,N_3558);
xor U3657 (N_3657,N_3531,N_3582);
xor U3658 (N_3658,N_3543,N_3514);
or U3659 (N_3659,N_3587,N_3596);
nand U3660 (N_3660,N_3568,N_3519);
xor U3661 (N_3661,N_3534,N_3559);
and U3662 (N_3662,N_3566,N_3574);
and U3663 (N_3663,N_3550,N_3579);
xor U3664 (N_3664,N_3514,N_3503);
and U3665 (N_3665,N_3551,N_3584);
and U3666 (N_3666,N_3515,N_3513);
nor U3667 (N_3667,N_3538,N_3592);
nor U3668 (N_3668,N_3594,N_3569);
and U3669 (N_3669,N_3506,N_3596);
and U3670 (N_3670,N_3580,N_3575);
nand U3671 (N_3671,N_3505,N_3546);
nor U3672 (N_3672,N_3590,N_3520);
and U3673 (N_3673,N_3536,N_3528);
nor U3674 (N_3674,N_3504,N_3582);
nor U3675 (N_3675,N_3537,N_3501);
and U3676 (N_3676,N_3558,N_3548);
nor U3677 (N_3677,N_3522,N_3559);
nor U3678 (N_3678,N_3599,N_3576);
and U3679 (N_3679,N_3506,N_3572);
nor U3680 (N_3680,N_3503,N_3564);
and U3681 (N_3681,N_3503,N_3532);
or U3682 (N_3682,N_3502,N_3508);
or U3683 (N_3683,N_3567,N_3515);
or U3684 (N_3684,N_3532,N_3558);
nor U3685 (N_3685,N_3575,N_3548);
or U3686 (N_3686,N_3564,N_3565);
nand U3687 (N_3687,N_3507,N_3582);
and U3688 (N_3688,N_3572,N_3586);
or U3689 (N_3689,N_3512,N_3599);
nand U3690 (N_3690,N_3595,N_3524);
or U3691 (N_3691,N_3587,N_3570);
nor U3692 (N_3692,N_3557,N_3502);
xnor U3693 (N_3693,N_3556,N_3595);
or U3694 (N_3694,N_3527,N_3508);
and U3695 (N_3695,N_3569,N_3575);
and U3696 (N_3696,N_3556,N_3554);
nor U3697 (N_3697,N_3593,N_3531);
nor U3698 (N_3698,N_3537,N_3523);
or U3699 (N_3699,N_3589,N_3519);
or U3700 (N_3700,N_3609,N_3645);
xor U3701 (N_3701,N_3642,N_3611);
or U3702 (N_3702,N_3628,N_3615);
and U3703 (N_3703,N_3654,N_3668);
and U3704 (N_3704,N_3632,N_3663);
nor U3705 (N_3705,N_3604,N_3689);
xor U3706 (N_3706,N_3695,N_3636);
or U3707 (N_3707,N_3666,N_3683);
and U3708 (N_3708,N_3682,N_3605);
nor U3709 (N_3709,N_3675,N_3618);
nor U3710 (N_3710,N_3698,N_3655);
nand U3711 (N_3711,N_3662,N_3680);
or U3712 (N_3712,N_3641,N_3684);
and U3713 (N_3713,N_3624,N_3650);
and U3714 (N_3714,N_3620,N_3661);
nor U3715 (N_3715,N_3676,N_3687);
nand U3716 (N_3716,N_3633,N_3603);
or U3717 (N_3717,N_3613,N_3651);
nand U3718 (N_3718,N_3647,N_3610);
and U3719 (N_3719,N_3634,N_3670);
and U3720 (N_3720,N_3619,N_3601);
nand U3721 (N_3721,N_3659,N_3600);
nand U3722 (N_3722,N_3625,N_3699);
or U3723 (N_3723,N_3614,N_3674);
and U3724 (N_3724,N_3665,N_3622);
nor U3725 (N_3725,N_3690,N_3691);
and U3726 (N_3726,N_3686,N_3696);
and U3727 (N_3727,N_3629,N_3671);
nor U3728 (N_3728,N_3631,N_3644);
or U3729 (N_3729,N_3630,N_3688);
xor U3730 (N_3730,N_3653,N_3673);
nand U3731 (N_3731,N_3623,N_3617);
and U3732 (N_3732,N_3692,N_3669);
or U3733 (N_3733,N_3685,N_3627);
or U3734 (N_3734,N_3656,N_3658);
or U3735 (N_3735,N_3602,N_3679);
and U3736 (N_3736,N_3697,N_3621);
or U3737 (N_3737,N_3678,N_3677);
and U3738 (N_3738,N_3664,N_3616);
nor U3739 (N_3739,N_3672,N_3626);
nor U3740 (N_3740,N_3646,N_3635);
nand U3741 (N_3741,N_3667,N_3612);
or U3742 (N_3742,N_3660,N_3607);
nor U3743 (N_3743,N_3640,N_3637);
nand U3744 (N_3744,N_3693,N_3681);
nor U3745 (N_3745,N_3639,N_3606);
nor U3746 (N_3746,N_3643,N_3694);
or U3747 (N_3747,N_3652,N_3657);
nor U3748 (N_3748,N_3649,N_3608);
or U3749 (N_3749,N_3638,N_3648);
and U3750 (N_3750,N_3664,N_3629);
nor U3751 (N_3751,N_3691,N_3631);
and U3752 (N_3752,N_3622,N_3656);
and U3753 (N_3753,N_3680,N_3688);
and U3754 (N_3754,N_3645,N_3692);
nor U3755 (N_3755,N_3697,N_3650);
nand U3756 (N_3756,N_3628,N_3664);
nand U3757 (N_3757,N_3635,N_3684);
nor U3758 (N_3758,N_3619,N_3608);
nor U3759 (N_3759,N_3651,N_3623);
and U3760 (N_3760,N_3688,N_3649);
and U3761 (N_3761,N_3678,N_3675);
or U3762 (N_3762,N_3638,N_3614);
nand U3763 (N_3763,N_3614,N_3611);
xor U3764 (N_3764,N_3609,N_3627);
nand U3765 (N_3765,N_3633,N_3632);
or U3766 (N_3766,N_3617,N_3631);
nand U3767 (N_3767,N_3647,N_3671);
and U3768 (N_3768,N_3627,N_3634);
and U3769 (N_3769,N_3638,N_3693);
nand U3770 (N_3770,N_3603,N_3651);
xor U3771 (N_3771,N_3622,N_3626);
nor U3772 (N_3772,N_3649,N_3616);
xnor U3773 (N_3773,N_3671,N_3641);
or U3774 (N_3774,N_3667,N_3663);
nand U3775 (N_3775,N_3601,N_3692);
and U3776 (N_3776,N_3649,N_3638);
xor U3777 (N_3777,N_3609,N_3602);
nand U3778 (N_3778,N_3658,N_3600);
nand U3779 (N_3779,N_3637,N_3665);
nor U3780 (N_3780,N_3622,N_3604);
nand U3781 (N_3781,N_3632,N_3642);
xnor U3782 (N_3782,N_3698,N_3665);
nor U3783 (N_3783,N_3611,N_3610);
and U3784 (N_3784,N_3663,N_3624);
nor U3785 (N_3785,N_3613,N_3618);
nand U3786 (N_3786,N_3676,N_3659);
nand U3787 (N_3787,N_3642,N_3641);
and U3788 (N_3788,N_3694,N_3609);
nand U3789 (N_3789,N_3601,N_3668);
and U3790 (N_3790,N_3659,N_3635);
and U3791 (N_3791,N_3610,N_3689);
or U3792 (N_3792,N_3698,N_3644);
xor U3793 (N_3793,N_3648,N_3609);
and U3794 (N_3794,N_3674,N_3644);
or U3795 (N_3795,N_3628,N_3614);
nand U3796 (N_3796,N_3693,N_3615);
and U3797 (N_3797,N_3655,N_3607);
and U3798 (N_3798,N_3630,N_3678);
nand U3799 (N_3799,N_3643,N_3612);
nor U3800 (N_3800,N_3772,N_3759);
nor U3801 (N_3801,N_3756,N_3721);
nor U3802 (N_3802,N_3793,N_3717);
nand U3803 (N_3803,N_3727,N_3776);
or U3804 (N_3804,N_3745,N_3760);
or U3805 (N_3805,N_3714,N_3729);
nor U3806 (N_3806,N_3703,N_3779);
and U3807 (N_3807,N_3720,N_3702);
and U3808 (N_3808,N_3722,N_3784);
nand U3809 (N_3809,N_3708,N_3766);
nor U3810 (N_3810,N_3768,N_3731);
nor U3811 (N_3811,N_3777,N_3786);
and U3812 (N_3812,N_3744,N_3797);
nor U3813 (N_3813,N_3757,N_3781);
or U3814 (N_3814,N_3735,N_3719);
and U3815 (N_3815,N_3743,N_3794);
or U3816 (N_3816,N_3733,N_3747);
and U3817 (N_3817,N_3758,N_3737);
and U3818 (N_3818,N_3700,N_3775);
nand U3819 (N_3819,N_3767,N_3763);
nand U3820 (N_3820,N_3723,N_3732);
xor U3821 (N_3821,N_3738,N_3785);
and U3822 (N_3822,N_3780,N_3754);
nand U3823 (N_3823,N_3778,N_3704);
nor U3824 (N_3824,N_3791,N_3782);
nor U3825 (N_3825,N_3787,N_3709);
or U3826 (N_3826,N_3726,N_3746);
or U3827 (N_3827,N_3707,N_3774);
nand U3828 (N_3828,N_3705,N_3799);
xnor U3829 (N_3829,N_3740,N_3715);
nor U3830 (N_3830,N_3750,N_3769);
xor U3831 (N_3831,N_3790,N_3788);
nor U3832 (N_3832,N_3718,N_3713);
and U3833 (N_3833,N_3771,N_3761);
and U3834 (N_3834,N_3789,N_3773);
nand U3835 (N_3835,N_3716,N_3762);
and U3836 (N_3836,N_3795,N_3753);
and U3837 (N_3837,N_3783,N_3765);
and U3838 (N_3838,N_3755,N_3798);
nor U3839 (N_3839,N_3751,N_3770);
or U3840 (N_3840,N_3736,N_3739);
or U3841 (N_3841,N_3749,N_3710);
and U3842 (N_3842,N_3741,N_3701);
or U3843 (N_3843,N_3728,N_3734);
or U3844 (N_3844,N_3712,N_3742);
and U3845 (N_3845,N_3724,N_3764);
nor U3846 (N_3846,N_3730,N_3748);
nor U3847 (N_3847,N_3711,N_3792);
nand U3848 (N_3848,N_3725,N_3796);
or U3849 (N_3849,N_3752,N_3706);
nor U3850 (N_3850,N_3747,N_3727);
and U3851 (N_3851,N_3759,N_3743);
nor U3852 (N_3852,N_3735,N_3709);
and U3853 (N_3853,N_3702,N_3751);
and U3854 (N_3854,N_3726,N_3767);
xor U3855 (N_3855,N_3762,N_3721);
nand U3856 (N_3856,N_3707,N_3755);
or U3857 (N_3857,N_3734,N_3708);
and U3858 (N_3858,N_3786,N_3700);
nand U3859 (N_3859,N_3716,N_3752);
or U3860 (N_3860,N_3787,N_3754);
or U3861 (N_3861,N_3759,N_3721);
nor U3862 (N_3862,N_3716,N_3706);
nand U3863 (N_3863,N_3748,N_3731);
nand U3864 (N_3864,N_3735,N_3799);
or U3865 (N_3865,N_3700,N_3746);
nand U3866 (N_3866,N_3757,N_3766);
nor U3867 (N_3867,N_3782,N_3727);
and U3868 (N_3868,N_3715,N_3750);
nand U3869 (N_3869,N_3731,N_3789);
xor U3870 (N_3870,N_3773,N_3731);
nand U3871 (N_3871,N_3766,N_3753);
or U3872 (N_3872,N_3737,N_3783);
xor U3873 (N_3873,N_3750,N_3757);
nand U3874 (N_3874,N_3754,N_3731);
and U3875 (N_3875,N_3763,N_3701);
or U3876 (N_3876,N_3790,N_3737);
and U3877 (N_3877,N_3794,N_3785);
and U3878 (N_3878,N_3761,N_3742);
nand U3879 (N_3879,N_3764,N_3721);
nor U3880 (N_3880,N_3729,N_3774);
nor U3881 (N_3881,N_3712,N_3720);
nor U3882 (N_3882,N_3718,N_3701);
nand U3883 (N_3883,N_3768,N_3716);
or U3884 (N_3884,N_3722,N_3796);
and U3885 (N_3885,N_3710,N_3735);
or U3886 (N_3886,N_3749,N_3760);
or U3887 (N_3887,N_3774,N_3747);
or U3888 (N_3888,N_3752,N_3700);
nand U3889 (N_3889,N_3752,N_3755);
nand U3890 (N_3890,N_3756,N_3789);
or U3891 (N_3891,N_3787,N_3705);
nor U3892 (N_3892,N_3745,N_3773);
or U3893 (N_3893,N_3745,N_3790);
xnor U3894 (N_3894,N_3726,N_3797);
and U3895 (N_3895,N_3788,N_3711);
nor U3896 (N_3896,N_3786,N_3744);
or U3897 (N_3897,N_3710,N_3750);
xnor U3898 (N_3898,N_3766,N_3703);
and U3899 (N_3899,N_3717,N_3776);
nand U3900 (N_3900,N_3881,N_3803);
nand U3901 (N_3901,N_3842,N_3822);
and U3902 (N_3902,N_3888,N_3839);
or U3903 (N_3903,N_3897,N_3886);
nor U3904 (N_3904,N_3854,N_3808);
and U3905 (N_3905,N_3817,N_3809);
or U3906 (N_3906,N_3806,N_3862);
and U3907 (N_3907,N_3826,N_3813);
or U3908 (N_3908,N_3887,N_3846);
xor U3909 (N_3909,N_3891,N_3857);
nand U3910 (N_3910,N_3878,N_3876);
and U3911 (N_3911,N_3816,N_3855);
nor U3912 (N_3912,N_3820,N_3879);
and U3913 (N_3913,N_3827,N_3858);
or U3914 (N_3914,N_3838,N_3843);
xor U3915 (N_3915,N_3890,N_3895);
xor U3916 (N_3916,N_3883,N_3896);
nor U3917 (N_3917,N_3872,N_3869);
and U3918 (N_3918,N_3829,N_3812);
nor U3919 (N_3919,N_3844,N_3892);
nand U3920 (N_3920,N_3814,N_3823);
nand U3921 (N_3921,N_3852,N_3859);
or U3922 (N_3922,N_3866,N_3899);
nand U3923 (N_3923,N_3882,N_3804);
nor U3924 (N_3924,N_3837,N_3832);
and U3925 (N_3925,N_3853,N_3849);
and U3926 (N_3926,N_3835,N_3867);
nor U3927 (N_3927,N_3871,N_3811);
nand U3928 (N_3928,N_3877,N_3861);
or U3929 (N_3929,N_3893,N_3851);
nor U3930 (N_3930,N_3870,N_3841);
xnor U3931 (N_3931,N_3824,N_3863);
nand U3932 (N_3932,N_3874,N_3856);
nand U3933 (N_3933,N_3830,N_3840);
nand U3934 (N_3934,N_3821,N_3815);
or U3935 (N_3935,N_3873,N_3818);
or U3936 (N_3936,N_3845,N_3885);
nand U3937 (N_3937,N_3898,N_3889);
nand U3938 (N_3938,N_3834,N_3805);
or U3939 (N_3939,N_3875,N_3860);
xnor U3940 (N_3940,N_3864,N_3807);
or U3941 (N_3941,N_3847,N_3880);
and U3942 (N_3942,N_3831,N_3802);
xor U3943 (N_3943,N_3833,N_3819);
nand U3944 (N_3944,N_3828,N_3868);
or U3945 (N_3945,N_3801,N_3894);
nor U3946 (N_3946,N_3850,N_3800);
nor U3947 (N_3947,N_3825,N_3836);
nor U3948 (N_3948,N_3884,N_3848);
nand U3949 (N_3949,N_3865,N_3810);
nor U3950 (N_3950,N_3800,N_3833);
or U3951 (N_3951,N_3812,N_3869);
nor U3952 (N_3952,N_3833,N_3864);
nand U3953 (N_3953,N_3839,N_3833);
nor U3954 (N_3954,N_3878,N_3877);
and U3955 (N_3955,N_3876,N_3825);
nor U3956 (N_3956,N_3898,N_3821);
nor U3957 (N_3957,N_3885,N_3869);
or U3958 (N_3958,N_3877,N_3816);
and U3959 (N_3959,N_3839,N_3827);
nor U3960 (N_3960,N_3812,N_3804);
and U3961 (N_3961,N_3838,N_3812);
nor U3962 (N_3962,N_3847,N_3877);
and U3963 (N_3963,N_3869,N_3802);
nand U3964 (N_3964,N_3831,N_3889);
and U3965 (N_3965,N_3887,N_3873);
and U3966 (N_3966,N_3860,N_3861);
or U3967 (N_3967,N_3857,N_3818);
nor U3968 (N_3968,N_3867,N_3861);
nor U3969 (N_3969,N_3846,N_3802);
nor U3970 (N_3970,N_3874,N_3807);
or U3971 (N_3971,N_3866,N_3801);
and U3972 (N_3972,N_3833,N_3830);
or U3973 (N_3973,N_3822,N_3860);
and U3974 (N_3974,N_3850,N_3890);
or U3975 (N_3975,N_3852,N_3823);
or U3976 (N_3976,N_3866,N_3830);
nand U3977 (N_3977,N_3838,N_3823);
nand U3978 (N_3978,N_3837,N_3860);
nand U3979 (N_3979,N_3837,N_3813);
and U3980 (N_3980,N_3818,N_3885);
nor U3981 (N_3981,N_3825,N_3865);
nand U3982 (N_3982,N_3842,N_3848);
and U3983 (N_3983,N_3819,N_3823);
and U3984 (N_3984,N_3869,N_3894);
nand U3985 (N_3985,N_3855,N_3893);
and U3986 (N_3986,N_3817,N_3848);
and U3987 (N_3987,N_3846,N_3884);
nand U3988 (N_3988,N_3892,N_3831);
and U3989 (N_3989,N_3855,N_3827);
nand U3990 (N_3990,N_3820,N_3862);
xor U3991 (N_3991,N_3800,N_3808);
or U3992 (N_3992,N_3888,N_3872);
or U3993 (N_3993,N_3856,N_3899);
nand U3994 (N_3994,N_3852,N_3809);
or U3995 (N_3995,N_3840,N_3800);
and U3996 (N_3996,N_3819,N_3822);
or U3997 (N_3997,N_3843,N_3868);
nor U3998 (N_3998,N_3839,N_3834);
and U3999 (N_3999,N_3862,N_3853);
and U4000 (N_4000,N_3990,N_3944);
or U4001 (N_4001,N_3933,N_3938);
nor U4002 (N_4002,N_3979,N_3922);
nand U4003 (N_4003,N_3927,N_3984);
nand U4004 (N_4004,N_3951,N_3970);
or U4005 (N_4005,N_3946,N_3965);
or U4006 (N_4006,N_3973,N_3982);
nor U4007 (N_4007,N_3931,N_3959);
or U4008 (N_4008,N_3958,N_3953);
or U4009 (N_4009,N_3978,N_3923);
and U4010 (N_4010,N_3918,N_3957);
and U4011 (N_4011,N_3907,N_3971);
xor U4012 (N_4012,N_3992,N_3967);
nor U4013 (N_4013,N_3915,N_3916);
or U4014 (N_4014,N_3964,N_3932);
nor U4015 (N_4015,N_3924,N_3960);
nor U4016 (N_4016,N_3909,N_3952);
nand U4017 (N_4017,N_3997,N_3980);
and U4018 (N_4018,N_3977,N_3903);
nand U4019 (N_4019,N_3963,N_3904);
xor U4020 (N_4020,N_3940,N_3947);
and U4021 (N_4021,N_3985,N_3987);
and U4022 (N_4022,N_3975,N_3906);
and U4023 (N_4023,N_3939,N_3908);
nor U4024 (N_4024,N_3913,N_3943);
nand U4025 (N_4025,N_3935,N_3945);
or U4026 (N_4026,N_3936,N_3954);
nand U4027 (N_4027,N_3974,N_3994);
nand U4028 (N_4028,N_3949,N_3998);
xnor U4029 (N_4029,N_3996,N_3948);
nand U4030 (N_4030,N_3914,N_3900);
xor U4031 (N_4031,N_3955,N_3966);
nor U4032 (N_4032,N_3919,N_3917);
and U4033 (N_4033,N_3910,N_3911);
nor U4034 (N_4034,N_3930,N_3950);
nand U4035 (N_4035,N_3993,N_3972);
xnor U4036 (N_4036,N_3962,N_3925);
and U4037 (N_4037,N_3905,N_3968);
nand U4038 (N_4038,N_3983,N_3921);
nor U4039 (N_4039,N_3934,N_3902);
and U4040 (N_4040,N_3976,N_3920);
nand U4041 (N_4041,N_3986,N_3999);
xnor U4042 (N_4042,N_3969,N_3901);
and U4043 (N_4043,N_3991,N_3989);
and U4044 (N_4044,N_3956,N_3937);
or U4045 (N_4045,N_3926,N_3942);
and U4046 (N_4046,N_3961,N_3988);
nand U4047 (N_4047,N_3929,N_3995);
nand U4048 (N_4048,N_3928,N_3941);
nand U4049 (N_4049,N_3912,N_3981);
nor U4050 (N_4050,N_3937,N_3938);
nand U4051 (N_4051,N_3941,N_3924);
and U4052 (N_4052,N_3910,N_3966);
and U4053 (N_4053,N_3944,N_3972);
and U4054 (N_4054,N_3989,N_3919);
nor U4055 (N_4055,N_3900,N_3995);
nor U4056 (N_4056,N_3956,N_3978);
and U4057 (N_4057,N_3983,N_3966);
nor U4058 (N_4058,N_3953,N_3931);
nor U4059 (N_4059,N_3979,N_3978);
xor U4060 (N_4060,N_3907,N_3929);
nor U4061 (N_4061,N_3900,N_3908);
nor U4062 (N_4062,N_3972,N_3961);
nor U4063 (N_4063,N_3923,N_3960);
or U4064 (N_4064,N_3978,N_3957);
nor U4065 (N_4065,N_3997,N_3978);
nand U4066 (N_4066,N_3937,N_3968);
or U4067 (N_4067,N_3920,N_3975);
nand U4068 (N_4068,N_3979,N_3934);
and U4069 (N_4069,N_3942,N_3973);
nand U4070 (N_4070,N_3977,N_3993);
nand U4071 (N_4071,N_3901,N_3937);
nand U4072 (N_4072,N_3997,N_3974);
xor U4073 (N_4073,N_3923,N_3965);
and U4074 (N_4074,N_3904,N_3943);
or U4075 (N_4075,N_3991,N_3905);
nor U4076 (N_4076,N_3943,N_3997);
and U4077 (N_4077,N_3918,N_3971);
and U4078 (N_4078,N_3950,N_3977);
or U4079 (N_4079,N_3989,N_3961);
nand U4080 (N_4080,N_3938,N_3936);
or U4081 (N_4081,N_3970,N_3941);
and U4082 (N_4082,N_3950,N_3968);
xor U4083 (N_4083,N_3996,N_3913);
and U4084 (N_4084,N_3997,N_3985);
and U4085 (N_4085,N_3962,N_3938);
or U4086 (N_4086,N_3999,N_3957);
xnor U4087 (N_4087,N_3985,N_3945);
or U4088 (N_4088,N_3953,N_3985);
nor U4089 (N_4089,N_3959,N_3957);
nor U4090 (N_4090,N_3995,N_3984);
nor U4091 (N_4091,N_3929,N_3936);
and U4092 (N_4092,N_3919,N_3918);
nand U4093 (N_4093,N_3990,N_3934);
nor U4094 (N_4094,N_3910,N_3968);
and U4095 (N_4095,N_3925,N_3948);
nand U4096 (N_4096,N_3983,N_3912);
nor U4097 (N_4097,N_3941,N_3976);
xnor U4098 (N_4098,N_3971,N_3914);
and U4099 (N_4099,N_3922,N_3961);
xor U4100 (N_4100,N_4045,N_4094);
nand U4101 (N_4101,N_4082,N_4041);
and U4102 (N_4102,N_4087,N_4026);
nor U4103 (N_4103,N_4077,N_4070);
or U4104 (N_4104,N_4052,N_4043);
or U4105 (N_4105,N_4009,N_4076);
nand U4106 (N_4106,N_4096,N_4097);
nor U4107 (N_4107,N_4039,N_4008);
nand U4108 (N_4108,N_4061,N_4035);
nand U4109 (N_4109,N_4065,N_4000);
and U4110 (N_4110,N_4057,N_4089);
or U4111 (N_4111,N_4085,N_4071);
nand U4112 (N_4112,N_4074,N_4086);
and U4113 (N_4113,N_4038,N_4046);
and U4114 (N_4114,N_4080,N_4064);
nand U4115 (N_4115,N_4090,N_4069);
xor U4116 (N_4116,N_4019,N_4048);
nor U4117 (N_4117,N_4095,N_4088);
or U4118 (N_4118,N_4013,N_4033);
or U4119 (N_4119,N_4053,N_4058);
xor U4120 (N_4120,N_4036,N_4078);
or U4121 (N_4121,N_4011,N_4040);
nor U4122 (N_4122,N_4056,N_4002);
and U4123 (N_4123,N_4005,N_4001);
xor U4124 (N_4124,N_4092,N_4029);
nor U4125 (N_4125,N_4099,N_4066);
xnor U4126 (N_4126,N_4017,N_4044);
and U4127 (N_4127,N_4068,N_4059);
or U4128 (N_4128,N_4030,N_4023);
xnor U4129 (N_4129,N_4047,N_4067);
and U4130 (N_4130,N_4054,N_4072);
nor U4131 (N_4131,N_4021,N_4042);
and U4132 (N_4132,N_4025,N_4050);
nor U4133 (N_4133,N_4028,N_4016);
nand U4134 (N_4134,N_4010,N_4032);
and U4135 (N_4135,N_4020,N_4098);
and U4136 (N_4136,N_4062,N_4073);
nor U4137 (N_4137,N_4049,N_4006);
or U4138 (N_4138,N_4012,N_4083);
or U4139 (N_4139,N_4063,N_4081);
and U4140 (N_4140,N_4075,N_4018);
xnor U4141 (N_4141,N_4055,N_4022);
and U4142 (N_4142,N_4091,N_4079);
nand U4143 (N_4143,N_4037,N_4027);
and U4144 (N_4144,N_4003,N_4024);
nor U4145 (N_4145,N_4031,N_4051);
nor U4146 (N_4146,N_4034,N_4014);
nor U4147 (N_4147,N_4015,N_4004);
and U4148 (N_4148,N_4007,N_4084);
nor U4149 (N_4149,N_4093,N_4060);
and U4150 (N_4150,N_4019,N_4008);
and U4151 (N_4151,N_4089,N_4052);
or U4152 (N_4152,N_4047,N_4049);
nand U4153 (N_4153,N_4094,N_4009);
and U4154 (N_4154,N_4010,N_4023);
or U4155 (N_4155,N_4039,N_4029);
xnor U4156 (N_4156,N_4095,N_4004);
nand U4157 (N_4157,N_4051,N_4020);
or U4158 (N_4158,N_4088,N_4046);
nand U4159 (N_4159,N_4060,N_4064);
and U4160 (N_4160,N_4039,N_4067);
or U4161 (N_4161,N_4081,N_4050);
and U4162 (N_4162,N_4059,N_4069);
and U4163 (N_4163,N_4060,N_4074);
or U4164 (N_4164,N_4081,N_4070);
or U4165 (N_4165,N_4080,N_4069);
and U4166 (N_4166,N_4014,N_4047);
nor U4167 (N_4167,N_4027,N_4026);
nor U4168 (N_4168,N_4093,N_4027);
or U4169 (N_4169,N_4085,N_4066);
and U4170 (N_4170,N_4000,N_4066);
nor U4171 (N_4171,N_4045,N_4059);
and U4172 (N_4172,N_4098,N_4058);
or U4173 (N_4173,N_4096,N_4079);
xor U4174 (N_4174,N_4007,N_4003);
or U4175 (N_4175,N_4020,N_4039);
and U4176 (N_4176,N_4025,N_4024);
xnor U4177 (N_4177,N_4038,N_4092);
nor U4178 (N_4178,N_4033,N_4023);
or U4179 (N_4179,N_4006,N_4009);
xnor U4180 (N_4180,N_4098,N_4060);
nor U4181 (N_4181,N_4032,N_4038);
or U4182 (N_4182,N_4029,N_4026);
and U4183 (N_4183,N_4053,N_4098);
and U4184 (N_4184,N_4003,N_4062);
and U4185 (N_4185,N_4071,N_4019);
nor U4186 (N_4186,N_4081,N_4059);
and U4187 (N_4187,N_4064,N_4012);
nor U4188 (N_4188,N_4088,N_4076);
nand U4189 (N_4189,N_4080,N_4011);
or U4190 (N_4190,N_4009,N_4051);
or U4191 (N_4191,N_4000,N_4015);
nor U4192 (N_4192,N_4016,N_4050);
nor U4193 (N_4193,N_4027,N_4036);
and U4194 (N_4194,N_4047,N_4010);
xnor U4195 (N_4195,N_4018,N_4058);
nand U4196 (N_4196,N_4037,N_4087);
nor U4197 (N_4197,N_4056,N_4063);
and U4198 (N_4198,N_4027,N_4024);
and U4199 (N_4199,N_4054,N_4082);
xor U4200 (N_4200,N_4185,N_4119);
or U4201 (N_4201,N_4145,N_4182);
and U4202 (N_4202,N_4194,N_4136);
and U4203 (N_4203,N_4164,N_4113);
or U4204 (N_4204,N_4124,N_4181);
or U4205 (N_4205,N_4190,N_4165);
and U4206 (N_4206,N_4196,N_4160);
xor U4207 (N_4207,N_4108,N_4118);
and U4208 (N_4208,N_4100,N_4172);
nor U4209 (N_4209,N_4104,N_4174);
nor U4210 (N_4210,N_4173,N_4162);
nand U4211 (N_4211,N_4116,N_4140);
nor U4212 (N_4212,N_4168,N_4142);
nand U4213 (N_4213,N_4139,N_4138);
and U4214 (N_4214,N_4106,N_4122);
nand U4215 (N_4215,N_4131,N_4127);
nor U4216 (N_4216,N_4105,N_4176);
or U4217 (N_4217,N_4149,N_4128);
or U4218 (N_4218,N_4126,N_4110);
or U4219 (N_4219,N_4132,N_4179);
and U4220 (N_4220,N_4159,N_4192);
xor U4221 (N_4221,N_4178,N_4171);
and U4222 (N_4222,N_4198,N_4199);
nor U4223 (N_4223,N_4137,N_4107);
or U4224 (N_4224,N_4195,N_4146);
nor U4225 (N_4225,N_4154,N_4188);
nand U4226 (N_4226,N_4177,N_4129);
nor U4227 (N_4227,N_4161,N_4197);
xnor U4228 (N_4228,N_4155,N_4150);
and U4229 (N_4229,N_4193,N_4166);
and U4230 (N_4230,N_4148,N_4183);
xor U4231 (N_4231,N_4123,N_4187);
nor U4232 (N_4232,N_4111,N_4158);
or U4233 (N_4233,N_4125,N_4121);
and U4234 (N_4234,N_4152,N_4101);
nand U4235 (N_4235,N_4102,N_4115);
nand U4236 (N_4236,N_4163,N_4103);
nor U4237 (N_4237,N_4133,N_4153);
or U4238 (N_4238,N_4114,N_4120);
nor U4239 (N_4239,N_4143,N_4141);
or U4240 (N_4240,N_4109,N_4134);
or U4241 (N_4241,N_4151,N_4130);
or U4242 (N_4242,N_4156,N_4112);
and U4243 (N_4243,N_4180,N_4135);
or U4244 (N_4244,N_4117,N_4170);
xor U4245 (N_4245,N_4144,N_4169);
or U4246 (N_4246,N_4191,N_4189);
or U4247 (N_4247,N_4184,N_4186);
nor U4248 (N_4248,N_4157,N_4175);
nand U4249 (N_4249,N_4167,N_4147);
xor U4250 (N_4250,N_4139,N_4110);
and U4251 (N_4251,N_4131,N_4180);
or U4252 (N_4252,N_4101,N_4120);
nand U4253 (N_4253,N_4175,N_4179);
and U4254 (N_4254,N_4145,N_4151);
and U4255 (N_4255,N_4139,N_4106);
nand U4256 (N_4256,N_4143,N_4152);
or U4257 (N_4257,N_4172,N_4166);
nor U4258 (N_4258,N_4128,N_4121);
and U4259 (N_4259,N_4113,N_4142);
and U4260 (N_4260,N_4177,N_4171);
nand U4261 (N_4261,N_4147,N_4106);
xor U4262 (N_4262,N_4156,N_4171);
nand U4263 (N_4263,N_4113,N_4150);
nor U4264 (N_4264,N_4153,N_4123);
or U4265 (N_4265,N_4114,N_4119);
xnor U4266 (N_4266,N_4176,N_4137);
nand U4267 (N_4267,N_4120,N_4132);
nor U4268 (N_4268,N_4103,N_4146);
or U4269 (N_4269,N_4151,N_4173);
or U4270 (N_4270,N_4101,N_4160);
nand U4271 (N_4271,N_4146,N_4120);
or U4272 (N_4272,N_4181,N_4191);
and U4273 (N_4273,N_4104,N_4124);
nor U4274 (N_4274,N_4137,N_4172);
or U4275 (N_4275,N_4151,N_4198);
nand U4276 (N_4276,N_4174,N_4132);
nand U4277 (N_4277,N_4121,N_4106);
nor U4278 (N_4278,N_4168,N_4195);
and U4279 (N_4279,N_4137,N_4138);
nand U4280 (N_4280,N_4159,N_4170);
and U4281 (N_4281,N_4172,N_4168);
or U4282 (N_4282,N_4172,N_4175);
or U4283 (N_4283,N_4104,N_4113);
or U4284 (N_4284,N_4192,N_4167);
nand U4285 (N_4285,N_4130,N_4165);
nor U4286 (N_4286,N_4109,N_4186);
and U4287 (N_4287,N_4130,N_4180);
and U4288 (N_4288,N_4182,N_4121);
nor U4289 (N_4289,N_4154,N_4139);
nand U4290 (N_4290,N_4147,N_4154);
nand U4291 (N_4291,N_4184,N_4167);
and U4292 (N_4292,N_4122,N_4135);
nor U4293 (N_4293,N_4155,N_4169);
nand U4294 (N_4294,N_4143,N_4134);
nand U4295 (N_4295,N_4111,N_4113);
and U4296 (N_4296,N_4106,N_4136);
or U4297 (N_4297,N_4115,N_4137);
and U4298 (N_4298,N_4132,N_4102);
or U4299 (N_4299,N_4181,N_4197);
and U4300 (N_4300,N_4295,N_4218);
nand U4301 (N_4301,N_4242,N_4281);
or U4302 (N_4302,N_4221,N_4283);
and U4303 (N_4303,N_4217,N_4255);
xor U4304 (N_4304,N_4244,N_4264);
nand U4305 (N_4305,N_4235,N_4253);
xor U4306 (N_4306,N_4233,N_4210);
and U4307 (N_4307,N_4268,N_4241);
nand U4308 (N_4308,N_4260,N_4280);
and U4309 (N_4309,N_4246,N_4216);
and U4310 (N_4310,N_4204,N_4273);
nand U4311 (N_4311,N_4276,N_4223);
nand U4312 (N_4312,N_4293,N_4226);
or U4313 (N_4313,N_4252,N_4256);
nand U4314 (N_4314,N_4278,N_4207);
or U4315 (N_4315,N_4294,N_4229);
nor U4316 (N_4316,N_4288,N_4237);
or U4317 (N_4317,N_4213,N_4239);
or U4318 (N_4318,N_4208,N_4209);
and U4319 (N_4319,N_4271,N_4258);
and U4320 (N_4320,N_4254,N_4206);
xnor U4321 (N_4321,N_4249,N_4257);
or U4322 (N_4322,N_4263,N_4220);
and U4323 (N_4323,N_4215,N_4224);
nand U4324 (N_4324,N_4269,N_4296);
nand U4325 (N_4325,N_4279,N_4265);
or U4326 (N_4326,N_4267,N_4291);
nor U4327 (N_4327,N_4251,N_4274);
nor U4328 (N_4328,N_4234,N_4222);
and U4329 (N_4329,N_4289,N_4275);
nand U4330 (N_4330,N_4250,N_4282);
nand U4331 (N_4331,N_4248,N_4262);
nand U4332 (N_4332,N_4202,N_4214);
or U4333 (N_4333,N_4285,N_4219);
nand U4334 (N_4334,N_4272,N_4290);
and U4335 (N_4335,N_4286,N_4259);
xnor U4336 (N_4336,N_4298,N_4211);
and U4337 (N_4337,N_4240,N_4247);
or U4338 (N_4338,N_4245,N_4225);
xnor U4339 (N_4339,N_4266,N_4201);
nor U4340 (N_4340,N_4238,N_4236);
or U4341 (N_4341,N_4228,N_4227);
nand U4342 (N_4342,N_4299,N_4297);
and U4343 (N_4343,N_4212,N_4270);
xor U4344 (N_4344,N_4205,N_4232);
and U4345 (N_4345,N_4200,N_4292);
or U4346 (N_4346,N_4243,N_4261);
xnor U4347 (N_4347,N_4277,N_4231);
nand U4348 (N_4348,N_4284,N_4230);
and U4349 (N_4349,N_4203,N_4287);
and U4350 (N_4350,N_4233,N_4242);
or U4351 (N_4351,N_4253,N_4297);
xor U4352 (N_4352,N_4297,N_4239);
or U4353 (N_4353,N_4272,N_4251);
xor U4354 (N_4354,N_4237,N_4282);
nor U4355 (N_4355,N_4211,N_4292);
or U4356 (N_4356,N_4242,N_4217);
nand U4357 (N_4357,N_4236,N_4264);
and U4358 (N_4358,N_4233,N_4243);
nand U4359 (N_4359,N_4225,N_4256);
nand U4360 (N_4360,N_4207,N_4275);
nor U4361 (N_4361,N_4253,N_4290);
or U4362 (N_4362,N_4289,N_4230);
or U4363 (N_4363,N_4217,N_4213);
nor U4364 (N_4364,N_4282,N_4253);
or U4365 (N_4365,N_4210,N_4224);
and U4366 (N_4366,N_4224,N_4291);
nand U4367 (N_4367,N_4206,N_4258);
and U4368 (N_4368,N_4289,N_4258);
or U4369 (N_4369,N_4263,N_4287);
or U4370 (N_4370,N_4283,N_4212);
or U4371 (N_4371,N_4243,N_4297);
nor U4372 (N_4372,N_4217,N_4240);
xor U4373 (N_4373,N_4285,N_4207);
nand U4374 (N_4374,N_4243,N_4295);
xor U4375 (N_4375,N_4251,N_4290);
nand U4376 (N_4376,N_4273,N_4252);
nand U4377 (N_4377,N_4201,N_4293);
nor U4378 (N_4378,N_4268,N_4253);
or U4379 (N_4379,N_4240,N_4254);
or U4380 (N_4380,N_4285,N_4261);
nor U4381 (N_4381,N_4222,N_4220);
or U4382 (N_4382,N_4224,N_4213);
and U4383 (N_4383,N_4248,N_4202);
or U4384 (N_4384,N_4261,N_4259);
nor U4385 (N_4385,N_4261,N_4219);
nor U4386 (N_4386,N_4255,N_4230);
nand U4387 (N_4387,N_4260,N_4256);
nor U4388 (N_4388,N_4275,N_4205);
or U4389 (N_4389,N_4296,N_4221);
nor U4390 (N_4390,N_4292,N_4285);
xnor U4391 (N_4391,N_4205,N_4245);
nand U4392 (N_4392,N_4275,N_4282);
nand U4393 (N_4393,N_4221,N_4209);
or U4394 (N_4394,N_4202,N_4254);
and U4395 (N_4395,N_4209,N_4230);
nand U4396 (N_4396,N_4261,N_4280);
xor U4397 (N_4397,N_4253,N_4222);
nor U4398 (N_4398,N_4276,N_4266);
or U4399 (N_4399,N_4239,N_4243);
and U4400 (N_4400,N_4309,N_4321);
and U4401 (N_4401,N_4340,N_4304);
or U4402 (N_4402,N_4348,N_4324);
nand U4403 (N_4403,N_4367,N_4372);
xor U4404 (N_4404,N_4350,N_4381);
xnor U4405 (N_4405,N_4301,N_4362);
nand U4406 (N_4406,N_4308,N_4319);
or U4407 (N_4407,N_4371,N_4384);
nand U4408 (N_4408,N_4368,N_4385);
and U4409 (N_4409,N_4361,N_4311);
nand U4410 (N_4410,N_4347,N_4388);
xnor U4411 (N_4411,N_4394,N_4335);
nand U4412 (N_4412,N_4332,N_4358);
or U4413 (N_4413,N_4320,N_4312);
nor U4414 (N_4414,N_4357,N_4354);
nand U4415 (N_4415,N_4339,N_4387);
or U4416 (N_4416,N_4389,N_4349);
or U4417 (N_4417,N_4378,N_4365);
or U4418 (N_4418,N_4398,N_4379);
and U4419 (N_4419,N_4359,N_4333);
nor U4420 (N_4420,N_4383,N_4346);
nor U4421 (N_4421,N_4344,N_4390);
or U4422 (N_4422,N_4395,N_4314);
and U4423 (N_4423,N_4352,N_4373);
and U4424 (N_4424,N_4399,N_4366);
nor U4425 (N_4425,N_4305,N_4386);
nand U4426 (N_4426,N_4318,N_4336);
xnor U4427 (N_4427,N_4393,N_4343);
nand U4428 (N_4428,N_4353,N_4322);
and U4429 (N_4429,N_4337,N_4341);
or U4430 (N_4430,N_4360,N_4307);
nand U4431 (N_4431,N_4323,N_4310);
nand U4432 (N_4432,N_4316,N_4338);
and U4433 (N_4433,N_4345,N_4326);
nor U4434 (N_4434,N_4396,N_4342);
nand U4435 (N_4435,N_4325,N_4382);
nand U4436 (N_4436,N_4363,N_4351);
nor U4437 (N_4437,N_4331,N_4313);
nand U4438 (N_4438,N_4317,N_4334);
xor U4439 (N_4439,N_4330,N_4369);
xor U4440 (N_4440,N_4356,N_4374);
or U4441 (N_4441,N_4302,N_4370);
and U4442 (N_4442,N_4329,N_4300);
nor U4443 (N_4443,N_4391,N_4315);
or U4444 (N_4444,N_4306,N_4328);
nor U4445 (N_4445,N_4380,N_4392);
nor U4446 (N_4446,N_4303,N_4375);
or U4447 (N_4447,N_4355,N_4376);
nor U4448 (N_4448,N_4327,N_4397);
nor U4449 (N_4449,N_4364,N_4377);
nor U4450 (N_4450,N_4388,N_4389);
or U4451 (N_4451,N_4309,N_4346);
nor U4452 (N_4452,N_4374,N_4355);
nand U4453 (N_4453,N_4398,N_4355);
nand U4454 (N_4454,N_4351,N_4388);
nand U4455 (N_4455,N_4332,N_4361);
or U4456 (N_4456,N_4317,N_4378);
xor U4457 (N_4457,N_4312,N_4399);
xor U4458 (N_4458,N_4394,N_4364);
and U4459 (N_4459,N_4336,N_4376);
and U4460 (N_4460,N_4395,N_4391);
nor U4461 (N_4461,N_4346,N_4313);
or U4462 (N_4462,N_4397,N_4324);
nor U4463 (N_4463,N_4379,N_4331);
xor U4464 (N_4464,N_4329,N_4384);
and U4465 (N_4465,N_4301,N_4397);
and U4466 (N_4466,N_4359,N_4383);
and U4467 (N_4467,N_4311,N_4367);
or U4468 (N_4468,N_4353,N_4366);
and U4469 (N_4469,N_4315,N_4320);
nor U4470 (N_4470,N_4342,N_4354);
nand U4471 (N_4471,N_4377,N_4387);
or U4472 (N_4472,N_4337,N_4345);
nor U4473 (N_4473,N_4335,N_4354);
nor U4474 (N_4474,N_4330,N_4307);
or U4475 (N_4475,N_4309,N_4307);
nor U4476 (N_4476,N_4307,N_4329);
and U4477 (N_4477,N_4318,N_4310);
nor U4478 (N_4478,N_4364,N_4376);
and U4479 (N_4479,N_4340,N_4388);
and U4480 (N_4480,N_4304,N_4317);
nand U4481 (N_4481,N_4337,N_4324);
nand U4482 (N_4482,N_4309,N_4313);
or U4483 (N_4483,N_4313,N_4305);
nor U4484 (N_4484,N_4329,N_4352);
nand U4485 (N_4485,N_4327,N_4392);
xor U4486 (N_4486,N_4355,N_4359);
and U4487 (N_4487,N_4357,N_4345);
nor U4488 (N_4488,N_4388,N_4372);
nand U4489 (N_4489,N_4352,N_4305);
and U4490 (N_4490,N_4342,N_4350);
and U4491 (N_4491,N_4383,N_4378);
nor U4492 (N_4492,N_4399,N_4323);
nor U4493 (N_4493,N_4345,N_4322);
nor U4494 (N_4494,N_4352,N_4377);
or U4495 (N_4495,N_4333,N_4334);
nand U4496 (N_4496,N_4357,N_4395);
and U4497 (N_4497,N_4356,N_4398);
nand U4498 (N_4498,N_4338,N_4357);
nor U4499 (N_4499,N_4335,N_4331);
or U4500 (N_4500,N_4495,N_4457);
or U4501 (N_4501,N_4463,N_4412);
and U4502 (N_4502,N_4436,N_4421);
nor U4503 (N_4503,N_4484,N_4411);
or U4504 (N_4504,N_4474,N_4435);
and U4505 (N_4505,N_4410,N_4427);
nor U4506 (N_4506,N_4478,N_4492);
and U4507 (N_4507,N_4455,N_4475);
xor U4508 (N_4508,N_4400,N_4479);
nor U4509 (N_4509,N_4477,N_4468);
xor U4510 (N_4510,N_4429,N_4403);
nor U4511 (N_4511,N_4426,N_4488);
nor U4512 (N_4512,N_4473,N_4481);
or U4513 (N_4513,N_4489,N_4456);
or U4514 (N_4514,N_4458,N_4425);
nand U4515 (N_4515,N_4487,N_4401);
nor U4516 (N_4516,N_4447,N_4444);
and U4517 (N_4517,N_4493,N_4428);
and U4518 (N_4518,N_4483,N_4482);
nor U4519 (N_4519,N_4496,N_4471);
or U4520 (N_4520,N_4442,N_4424);
nand U4521 (N_4521,N_4454,N_4459);
xnor U4522 (N_4522,N_4407,N_4486);
nand U4523 (N_4523,N_4490,N_4422);
or U4524 (N_4524,N_4430,N_4438);
xnor U4525 (N_4525,N_4434,N_4450);
xnor U4526 (N_4526,N_4497,N_4499);
xnor U4527 (N_4527,N_4409,N_4440);
nor U4528 (N_4528,N_4452,N_4451);
nor U4529 (N_4529,N_4423,N_4462);
nor U4530 (N_4530,N_4446,N_4418);
and U4531 (N_4531,N_4406,N_4443);
nand U4532 (N_4532,N_4439,N_4472);
and U4533 (N_4533,N_4413,N_4431);
or U4534 (N_4534,N_4491,N_4465);
xnor U4535 (N_4535,N_4420,N_4408);
nor U4536 (N_4536,N_4402,N_4464);
nand U4537 (N_4537,N_4485,N_4405);
nand U4538 (N_4538,N_4437,N_4448);
and U4539 (N_4539,N_4466,N_4441);
and U4540 (N_4540,N_4467,N_4470);
and U4541 (N_4541,N_4445,N_4469);
or U4542 (N_4542,N_4419,N_4415);
and U4543 (N_4543,N_4404,N_4417);
xor U4544 (N_4544,N_4416,N_4461);
xnor U4545 (N_4545,N_4432,N_4476);
xor U4546 (N_4546,N_4480,N_4453);
nand U4547 (N_4547,N_4449,N_4433);
nand U4548 (N_4548,N_4498,N_4460);
nand U4549 (N_4549,N_4494,N_4414);
and U4550 (N_4550,N_4457,N_4452);
nand U4551 (N_4551,N_4432,N_4460);
or U4552 (N_4552,N_4427,N_4474);
nand U4553 (N_4553,N_4417,N_4441);
nor U4554 (N_4554,N_4408,N_4425);
or U4555 (N_4555,N_4425,N_4470);
nand U4556 (N_4556,N_4439,N_4481);
or U4557 (N_4557,N_4485,N_4429);
or U4558 (N_4558,N_4451,N_4490);
or U4559 (N_4559,N_4446,N_4486);
or U4560 (N_4560,N_4488,N_4410);
or U4561 (N_4561,N_4426,N_4473);
or U4562 (N_4562,N_4468,N_4471);
nand U4563 (N_4563,N_4416,N_4400);
and U4564 (N_4564,N_4414,N_4426);
nand U4565 (N_4565,N_4406,N_4492);
xor U4566 (N_4566,N_4494,N_4423);
nand U4567 (N_4567,N_4409,N_4496);
xor U4568 (N_4568,N_4416,N_4486);
nor U4569 (N_4569,N_4433,N_4428);
nand U4570 (N_4570,N_4488,N_4450);
or U4571 (N_4571,N_4419,N_4418);
xor U4572 (N_4572,N_4404,N_4418);
nand U4573 (N_4573,N_4430,N_4499);
nand U4574 (N_4574,N_4482,N_4405);
nand U4575 (N_4575,N_4403,N_4435);
nand U4576 (N_4576,N_4424,N_4407);
xnor U4577 (N_4577,N_4491,N_4486);
nor U4578 (N_4578,N_4487,N_4433);
and U4579 (N_4579,N_4489,N_4448);
and U4580 (N_4580,N_4459,N_4442);
nor U4581 (N_4581,N_4494,N_4427);
or U4582 (N_4582,N_4493,N_4461);
and U4583 (N_4583,N_4492,N_4480);
and U4584 (N_4584,N_4436,N_4433);
and U4585 (N_4585,N_4401,N_4446);
nor U4586 (N_4586,N_4404,N_4463);
or U4587 (N_4587,N_4411,N_4436);
nand U4588 (N_4588,N_4405,N_4441);
nand U4589 (N_4589,N_4497,N_4489);
and U4590 (N_4590,N_4429,N_4444);
nand U4591 (N_4591,N_4449,N_4442);
or U4592 (N_4592,N_4421,N_4410);
or U4593 (N_4593,N_4400,N_4440);
nand U4594 (N_4594,N_4401,N_4476);
or U4595 (N_4595,N_4472,N_4422);
and U4596 (N_4596,N_4400,N_4474);
nor U4597 (N_4597,N_4467,N_4488);
nor U4598 (N_4598,N_4486,N_4403);
and U4599 (N_4599,N_4423,N_4406);
nor U4600 (N_4600,N_4551,N_4540);
nor U4601 (N_4601,N_4532,N_4567);
and U4602 (N_4602,N_4543,N_4581);
nand U4603 (N_4603,N_4546,N_4585);
nor U4604 (N_4604,N_4535,N_4515);
and U4605 (N_4605,N_4566,N_4572);
nor U4606 (N_4606,N_4598,N_4571);
or U4607 (N_4607,N_4501,N_4557);
and U4608 (N_4608,N_4514,N_4522);
nand U4609 (N_4609,N_4534,N_4510);
xnor U4610 (N_4610,N_4589,N_4556);
or U4611 (N_4611,N_4517,N_4502);
and U4612 (N_4612,N_4579,N_4563);
nor U4613 (N_4613,N_4539,N_4521);
nor U4614 (N_4614,N_4524,N_4525);
or U4615 (N_4615,N_4548,N_4529);
nand U4616 (N_4616,N_4575,N_4520);
and U4617 (N_4617,N_4594,N_4519);
nor U4618 (N_4618,N_4550,N_4507);
and U4619 (N_4619,N_4564,N_4512);
and U4620 (N_4620,N_4593,N_4537);
nor U4621 (N_4621,N_4583,N_4531);
and U4622 (N_4622,N_4576,N_4569);
and U4623 (N_4623,N_4586,N_4530);
and U4624 (N_4624,N_4560,N_4559);
or U4625 (N_4625,N_4595,N_4568);
and U4626 (N_4626,N_4511,N_4528);
xor U4627 (N_4627,N_4553,N_4500);
or U4628 (N_4628,N_4541,N_4513);
xnor U4629 (N_4629,N_4592,N_4542);
nor U4630 (N_4630,N_4555,N_4518);
nor U4631 (N_4631,N_4545,N_4552);
or U4632 (N_4632,N_4596,N_4526);
nand U4633 (N_4633,N_4580,N_4577);
xor U4634 (N_4634,N_4578,N_4527);
or U4635 (N_4635,N_4584,N_4554);
nor U4636 (N_4636,N_4533,N_4516);
and U4637 (N_4637,N_4523,N_4562);
or U4638 (N_4638,N_4547,N_4549);
nor U4639 (N_4639,N_4544,N_4504);
and U4640 (N_4640,N_4565,N_4588);
nand U4641 (N_4641,N_4590,N_4573);
xnor U4642 (N_4642,N_4508,N_4599);
or U4643 (N_4643,N_4582,N_4538);
or U4644 (N_4644,N_4509,N_4574);
nand U4645 (N_4645,N_4587,N_4597);
or U4646 (N_4646,N_4503,N_4558);
or U4647 (N_4647,N_4506,N_4505);
and U4648 (N_4648,N_4591,N_4570);
and U4649 (N_4649,N_4536,N_4561);
nand U4650 (N_4650,N_4550,N_4591);
nor U4651 (N_4651,N_4592,N_4584);
or U4652 (N_4652,N_4589,N_4568);
and U4653 (N_4653,N_4577,N_4564);
nor U4654 (N_4654,N_4521,N_4597);
nor U4655 (N_4655,N_4526,N_4548);
or U4656 (N_4656,N_4508,N_4569);
and U4657 (N_4657,N_4564,N_4520);
and U4658 (N_4658,N_4516,N_4540);
or U4659 (N_4659,N_4532,N_4597);
nor U4660 (N_4660,N_4599,N_4549);
and U4661 (N_4661,N_4596,N_4530);
nor U4662 (N_4662,N_4557,N_4553);
or U4663 (N_4663,N_4594,N_4563);
or U4664 (N_4664,N_4520,N_4596);
nor U4665 (N_4665,N_4581,N_4527);
nand U4666 (N_4666,N_4541,N_4596);
or U4667 (N_4667,N_4548,N_4567);
nor U4668 (N_4668,N_4554,N_4543);
and U4669 (N_4669,N_4572,N_4501);
nand U4670 (N_4670,N_4577,N_4524);
nor U4671 (N_4671,N_4531,N_4591);
and U4672 (N_4672,N_4599,N_4545);
and U4673 (N_4673,N_4586,N_4590);
xor U4674 (N_4674,N_4524,N_4546);
and U4675 (N_4675,N_4570,N_4507);
nand U4676 (N_4676,N_4558,N_4521);
nor U4677 (N_4677,N_4597,N_4517);
and U4678 (N_4678,N_4513,N_4509);
and U4679 (N_4679,N_4536,N_4543);
and U4680 (N_4680,N_4541,N_4588);
or U4681 (N_4681,N_4536,N_4510);
and U4682 (N_4682,N_4584,N_4536);
or U4683 (N_4683,N_4599,N_4531);
nor U4684 (N_4684,N_4543,N_4507);
or U4685 (N_4685,N_4508,N_4594);
or U4686 (N_4686,N_4537,N_4591);
xnor U4687 (N_4687,N_4577,N_4514);
nand U4688 (N_4688,N_4523,N_4537);
nand U4689 (N_4689,N_4520,N_4526);
nand U4690 (N_4690,N_4562,N_4541);
or U4691 (N_4691,N_4521,N_4541);
xor U4692 (N_4692,N_4558,N_4575);
or U4693 (N_4693,N_4572,N_4550);
nor U4694 (N_4694,N_4595,N_4548);
or U4695 (N_4695,N_4564,N_4543);
nand U4696 (N_4696,N_4517,N_4509);
nor U4697 (N_4697,N_4502,N_4549);
or U4698 (N_4698,N_4549,N_4586);
nor U4699 (N_4699,N_4556,N_4592);
nand U4700 (N_4700,N_4605,N_4679);
or U4701 (N_4701,N_4617,N_4635);
nor U4702 (N_4702,N_4632,N_4607);
or U4703 (N_4703,N_4673,N_4612);
xor U4704 (N_4704,N_4663,N_4629);
or U4705 (N_4705,N_4626,N_4609);
nor U4706 (N_4706,N_4647,N_4681);
and U4707 (N_4707,N_4661,N_4646);
or U4708 (N_4708,N_4641,N_4691);
or U4709 (N_4709,N_4693,N_4639);
nand U4710 (N_4710,N_4624,N_4692);
and U4711 (N_4711,N_4657,N_4633);
or U4712 (N_4712,N_4680,N_4616);
or U4713 (N_4713,N_4655,N_4690);
nor U4714 (N_4714,N_4606,N_4613);
nand U4715 (N_4715,N_4688,N_4615);
nor U4716 (N_4716,N_4667,N_4670);
nor U4717 (N_4717,N_4689,N_4630);
and U4718 (N_4718,N_4602,N_4634);
nand U4719 (N_4719,N_4662,N_4683);
xor U4720 (N_4720,N_4698,N_4653);
and U4721 (N_4721,N_4658,N_4644);
and U4722 (N_4722,N_4620,N_4695);
xnor U4723 (N_4723,N_4672,N_4645);
and U4724 (N_4724,N_4699,N_4614);
nor U4725 (N_4725,N_4654,N_4669);
and U4726 (N_4726,N_4652,N_4600);
or U4727 (N_4727,N_4684,N_4625);
nand U4728 (N_4728,N_4675,N_4619);
nand U4729 (N_4729,N_4697,N_4611);
nand U4730 (N_4730,N_4601,N_4671);
nor U4731 (N_4731,N_4682,N_4668);
and U4732 (N_4732,N_4610,N_4608);
nor U4733 (N_4733,N_4656,N_4678);
or U4734 (N_4734,N_4674,N_4650);
or U4735 (N_4735,N_4622,N_4604);
xnor U4736 (N_4736,N_4685,N_4648);
and U4737 (N_4737,N_4696,N_4666);
nand U4738 (N_4738,N_4618,N_4631);
nor U4739 (N_4739,N_4640,N_4638);
nand U4740 (N_4740,N_4649,N_4659);
nor U4741 (N_4741,N_4621,N_4628);
nor U4742 (N_4742,N_4643,N_4686);
xnor U4743 (N_4743,N_4651,N_4636);
nand U4744 (N_4744,N_4660,N_4677);
xnor U4745 (N_4745,N_4627,N_4694);
xor U4746 (N_4746,N_4676,N_4637);
nor U4747 (N_4747,N_4642,N_4603);
nor U4748 (N_4748,N_4623,N_4665);
or U4749 (N_4749,N_4687,N_4664);
nor U4750 (N_4750,N_4657,N_4629);
nor U4751 (N_4751,N_4685,N_4632);
nor U4752 (N_4752,N_4648,N_4677);
nand U4753 (N_4753,N_4603,N_4627);
and U4754 (N_4754,N_4609,N_4625);
nand U4755 (N_4755,N_4690,N_4625);
or U4756 (N_4756,N_4636,N_4661);
or U4757 (N_4757,N_4652,N_4676);
or U4758 (N_4758,N_4645,N_4610);
nand U4759 (N_4759,N_4638,N_4605);
or U4760 (N_4760,N_4637,N_4625);
nor U4761 (N_4761,N_4669,N_4671);
and U4762 (N_4762,N_4652,N_4648);
xnor U4763 (N_4763,N_4661,N_4634);
and U4764 (N_4764,N_4648,N_4622);
nor U4765 (N_4765,N_4626,N_4683);
nor U4766 (N_4766,N_4665,N_4682);
or U4767 (N_4767,N_4627,N_4666);
nor U4768 (N_4768,N_4611,N_4696);
nand U4769 (N_4769,N_4606,N_4648);
and U4770 (N_4770,N_4627,N_4656);
or U4771 (N_4771,N_4650,N_4686);
nor U4772 (N_4772,N_4646,N_4670);
xor U4773 (N_4773,N_4606,N_4670);
and U4774 (N_4774,N_4684,N_4670);
nand U4775 (N_4775,N_4655,N_4606);
xor U4776 (N_4776,N_4697,N_4662);
nand U4777 (N_4777,N_4698,N_4645);
nor U4778 (N_4778,N_4652,N_4614);
nand U4779 (N_4779,N_4699,N_4622);
nor U4780 (N_4780,N_4618,N_4628);
nor U4781 (N_4781,N_4616,N_4676);
nand U4782 (N_4782,N_4692,N_4614);
nor U4783 (N_4783,N_4639,N_4612);
nor U4784 (N_4784,N_4675,N_4697);
nor U4785 (N_4785,N_4634,N_4695);
or U4786 (N_4786,N_4621,N_4682);
or U4787 (N_4787,N_4664,N_4617);
nand U4788 (N_4788,N_4676,N_4661);
xor U4789 (N_4789,N_4642,N_4619);
nor U4790 (N_4790,N_4682,N_4622);
nand U4791 (N_4791,N_4630,N_4656);
nor U4792 (N_4792,N_4662,N_4692);
or U4793 (N_4793,N_4687,N_4662);
xor U4794 (N_4794,N_4638,N_4633);
nand U4795 (N_4795,N_4652,N_4672);
and U4796 (N_4796,N_4697,N_4608);
nor U4797 (N_4797,N_4624,N_4652);
or U4798 (N_4798,N_4635,N_4687);
xor U4799 (N_4799,N_4607,N_4653);
and U4800 (N_4800,N_4758,N_4791);
nand U4801 (N_4801,N_4724,N_4776);
nor U4802 (N_4802,N_4708,N_4741);
nand U4803 (N_4803,N_4786,N_4705);
nand U4804 (N_4804,N_4721,N_4756);
or U4805 (N_4805,N_4787,N_4729);
nor U4806 (N_4806,N_4757,N_4763);
and U4807 (N_4807,N_4754,N_4709);
nor U4808 (N_4808,N_4767,N_4726);
nand U4809 (N_4809,N_4722,N_4751);
nand U4810 (N_4810,N_4738,N_4771);
and U4811 (N_4811,N_4750,N_4784);
xor U4812 (N_4812,N_4752,N_4711);
nor U4813 (N_4813,N_4760,N_4740);
nor U4814 (N_4814,N_4727,N_4733);
and U4815 (N_4815,N_4725,N_4783);
nor U4816 (N_4816,N_4745,N_4768);
nand U4817 (N_4817,N_4706,N_4743);
nor U4818 (N_4818,N_4710,N_4764);
nand U4819 (N_4819,N_4755,N_4794);
or U4820 (N_4820,N_4735,N_4788);
nor U4821 (N_4821,N_4796,N_4716);
nand U4822 (N_4822,N_4799,N_4700);
nor U4823 (N_4823,N_4737,N_4769);
and U4824 (N_4824,N_4736,N_4703);
nor U4825 (N_4825,N_4747,N_4715);
nand U4826 (N_4826,N_4718,N_4714);
xor U4827 (N_4827,N_4761,N_4781);
nor U4828 (N_4828,N_4789,N_4744);
or U4829 (N_4829,N_4774,N_4739);
nand U4830 (N_4830,N_4773,N_4702);
or U4831 (N_4831,N_4748,N_4730);
nor U4832 (N_4832,N_4704,N_4766);
or U4833 (N_4833,N_4759,N_4795);
nor U4834 (N_4834,N_4792,N_4793);
or U4835 (N_4835,N_4734,N_4778);
or U4836 (N_4836,N_4779,N_4765);
or U4837 (N_4837,N_4775,N_4707);
xor U4838 (N_4838,N_4749,N_4782);
nor U4839 (N_4839,N_4797,N_4777);
or U4840 (N_4840,N_4798,N_4772);
or U4841 (N_4841,N_4720,N_4790);
and U4842 (N_4842,N_4780,N_4742);
and U4843 (N_4843,N_4719,N_4753);
nand U4844 (N_4844,N_4723,N_4712);
nor U4845 (N_4845,N_4728,N_4732);
nor U4846 (N_4846,N_4770,N_4762);
nand U4847 (N_4847,N_4731,N_4717);
nand U4848 (N_4848,N_4701,N_4746);
nand U4849 (N_4849,N_4713,N_4785);
nand U4850 (N_4850,N_4733,N_4706);
or U4851 (N_4851,N_4766,N_4748);
and U4852 (N_4852,N_4720,N_4789);
nand U4853 (N_4853,N_4747,N_4759);
and U4854 (N_4854,N_4771,N_4719);
and U4855 (N_4855,N_4782,N_4707);
nand U4856 (N_4856,N_4735,N_4734);
or U4857 (N_4857,N_4742,N_4712);
or U4858 (N_4858,N_4702,N_4740);
nand U4859 (N_4859,N_4741,N_4732);
nor U4860 (N_4860,N_4794,N_4723);
nor U4861 (N_4861,N_4796,N_4774);
nand U4862 (N_4862,N_4709,N_4738);
nor U4863 (N_4863,N_4777,N_4773);
and U4864 (N_4864,N_4761,N_4726);
or U4865 (N_4865,N_4756,N_4729);
nor U4866 (N_4866,N_4758,N_4778);
nand U4867 (N_4867,N_4742,N_4784);
and U4868 (N_4868,N_4727,N_4766);
and U4869 (N_4869,N_4717,N_4797);
nand U4870 (N_4870,N_4761,N_4791);
nor U4871 (N_4871,N_4737,N_4715);
xnor U4872 (N_4872,N_4783,N_4799);
or U4873 (N_4873,N_4757,N_4786);
nand U4874 (N_4874,N_4749,N_4788);
or U4875 (N_4875,N_4735,N_4727);
and U4876 (N_4876,N_4760,N_4716);
xnor U4877 (N_4877,N_4783,N_4719);
nor U4878 (N_4878,N_4771,N_4708);
and U4879 (N_4879,N_4766,N_4775);
nand U4880 (N_4880,N_4751,N_4787);
or U4881 (N_4881,N_4722,N_4756);
nor U4882 (N_4882,N_4799,N_4762);
and U4883 (N_4883,N_4734,N_4700);
and U4884 (N_4884,N_4769,N_4741);
xor U4885 (N_4885,N_4723,N_4741);
nor U4886 (N_4886,N_4715,N_4709);
or U4887 (N_4887,N_4727,N_4778);
or U4888 (N_4888,N_4743,N_4717);
nor U4889 (N_4889,N_4798,N_4793);
or U4890 (N_4890,N_4736,N_4704);
xnor U4891 (N_4891,N_4716,N_4742);
xnor U4892 (N_4892,N_4725,N_4709);
xnor U4893 (N_4893,N_4785,N_4755);
and U4894 (N_4894,N_4753,N_4778);
xnor U4895 (N_4895,N_4707,N_4717);
xnor U4896 (N_4896,N_4704,N_4712);
or U4897 (N_4897,N_4790,N_4713);
and U4898 (N_4898,N_4743,N_4753);
nor U4899 (N_4899,N_4796,N_4765);
nor U4900 (N_4900,N_4819,N_4870);
xor U4901 (N_4901,N_4863,N_4896);
nand U4902 (N_4902,N_4833,N_4818);
nor U4903 (N_4903,N_4846,N_4851);
nor U4904 (N_4904,N_4869,N_4830);
nor U4905 (N_4905,N_4844,N_4885);
nor U4906 (N_4906,N_4805,N_4838);
nand U4907 (N_4907,N_4865,N_4888);
and U4908 (N_4908,N_4824,N_4867);
and U4909 (N_4909,N_4866,N_4880);
nor U4910 (N_4910,N_4839,N_4868);
or U4911 (N_4911,N_4862,N_4860);
nor U4912 (N_4912,N_4875,N_4893);
xor U4913 (N_4913,N_4823,N_4806);
or U4914 (N_4914,N_4871,N_4822);
nand U4915 (N_4915,N_4841,N_4873);
xor U4916 (N_4916,N_4811,N_4874);
nor U4917 (N_4917,N_4872,N_4879);
nor U4918 (N_4918,N_4881,N_4840);
nand U4919 (N_4919,N_4887,N_4831);
nor U4920 (N_4920,N_4876,N_4899);
and U4921 (N_4921,N_4883,N_4803);
xor U4922 (N_4922,N_4853,N_4878);
or U4923 (N_4923,N_4828,N_4884);
and U4924 (N_4924,N_4837,N_4855);
nor U4925 (N_4925,N_4890,N_4847);
and U4926 (N_4926,N_4820,N_4809);
or U4927 (N_4927,N_4832,N_4882);
nand U4928 (N_4928,N_4815,N_4864);
and U4929 (N_4929,N_4849,N_4816);
and U4930 (N_4930,N_4845,N_4877);
nand U4931 (N_4931,N_4834,N_4895);
nor U4932 (N_4932,N_4817,N_4807);
nand U4933 (N_4933,N_4810,N_4808);
or U4934 (N_4934,N_4836,N_4843);
or U4935 (N_4935,N_4852,N_4858);
or U4936 (N_4936,N_4854,N_4800);
nor U4937 (N_4937,N_4892,N_4897);
or U4938 (N_4938,N_4861,N_4889);
nor U4939 (N_4939,N_4827,N_4814);
nand U4940 (N_4940,N_4857,N_4826);
nand U4941 (N_4941,N_4891,N_4802);
nand U4942 (N_4942,N_4848,N_4859);
nand U4943 (N_4943,N_4842,N_4856);
and U4944 (N_4944,N_4804,N_4821);
and U4945 (N_4945,N_4813,N_4898);
and U4946 (N_4946,N_4829,N_4835);
or U4947 (N_4947,N_4894,N_4886);
nand U4948 (N_4948,N_4801,N_4812);
or U4949 (N_4949,N_4850,N_4825);
or U4950 (N_4950,N_4837,N_4864);
xnor U4951 (N_4951,N_4857,N_4815);
nand U4952 (N_4952,N_4861,N_4893);
nor U4953 (N_4953,N_4843,N_4877);
and U4954 (N_4954,N_4834,N_4822);
and U4955 (N_4955,N_4804,N_4845);
or U4956 (N_4956,N_4846,N_4884);
nor U4957 (N_4957,N_4822,N_4800);
or U4958 (N_4958,N_4892,N_4820);
and U4959 (N_4959,N_4831,N_4826);
nor U4960 (N_4960,N_4820,N_4876);
or U4961 (N_4961,N_4814,N_4832);
or U4962 (N_4962,N_4818,N_4880);
nor U4963 (N_4963,N_4850,N_4833);
and U4964 (N_4964,N_4815,N_4830);
nand U4965 (N_4965,N_4862,N_4827);
xnor U4966 (N_4966,N_4880,N_4838);
xor U4967 (N_4967,N_4870,N_4846);
nor U4968 (N_4968,N_4840,N_4860);
nor U4969 (N_4969,N_4849,N_4874);
or U4970 (N_4970,N_4866,N_4809);
or U4971 (N_4971,N_4853,N_4823);
nor U4972 (N_4972,N_4861,N_4828);
nand U4973 (N_4973,N_4882,N_4875);
and U4974 (N_4974,N_4858,N_4819);
nor U4975 (N_4975,N_4811,N_4807);
and U4976 (N_4976,N_4883,N_4806);
nor U4977 (N_4977,N_4800,N_4891);
nor U4978 (N_4978,N_4897,N_4860);
nand U4979 (N_4979,N_4876,N_4851);
and U4980 (N_4980,N_4805,N_4885);
nor U4981 (N_4981,N_4807,N_4822);
or U4982 (N_4982,N_4802,N_4874);
or U4983 (N_4983,N_4852,N_4817);
xnor U4984 (N_4984,N_4881,N_4801);
or U4985 (N_4985,N_4835,N_4845);
and U4986 (N_4986,N_4802,N_4835);
nor U4987 (N_4987,N_4802,N_4894);
or U4988 (N_4988,N_4886,N_4828);
and U4989 (N_4989,N_4891,N_4855);
or U4990 (N_4990,N_4800,N_4859);
and U4991 (N_4991,N_4895,N_4857);
nand U4992 (N_4992,N_4861,N_4805);
and U4993 (N_4993,N_4853,N_4880);
or U4994 (N_4994,N_4833,N_4885);
or U4995 (N_4995,N_4811,N_4830);
nand U4996 (N_4996,N_4828,N_4863);
nor U4997 (N_4997,N_4827,N_4863);
nor U4998 (N_4998,N_4818,N_4800);
nor U4999 (N_4999,N_4870,N_4801);
and UO_0 (O_0,N_4919,N_4909);
nor UO_1 (O_1,N_4931,N_4949);
nor UO_2 (O_2,N_4924,N_4904);
and UO_3 (O_3,N_4984,N_4925);
nand UO_4 (O_4,N_4950,N_4970);
and UO_5 (O_5,N_4978,N_4911);
nor UO_6 (O_6,N_4997,N_4922);
nor UO_7 (O_7,N_4908,N_4920);
and UO_8 (O_8,N_4985,N_4974);
and UO_9 (O_9,N_4902,N_4957);
or UO_10 (O_10,N_4953,N_4972);
or UO_11 (O_11,N_4951,N_4960);
xor UO_12 (O_12,N_4938,N_4992);
nor UO_13 (O_13,N_4961,N_4993);
and UO_14 (O_14,N_4936,N_4965);
nand UO_15 (O_15,N_4939,N_4959);
xor UO_16 (O_16,N_4918,N_4937);
or UO_17 (O_17,N_4966,N_4947);
nor UO_18 (O_18,N_4975,N_4995);
nand UO_19 (O_19,N_4988,N_4930);
nor UO_20 (O_20,N_4907,N_4981);
xor UO_21 (O_21,N_4929,N_4945);
nor UO_22 (O_22,N_4921,N_4910);
xor UO_23 (O_23,N_4932,N_4944);
or UO_24 (O_24,N_4915,N_4905);
nor UO_25 (O_25,N_4967,N_4917);
and UO_26 (O_26,N_4989,N_4983);
or UO_27 (O_27,N_4994,N_4935);
nand UO_28 (O_28,N_4903,N_4996);
nor UO_29 (O_29,N_4906,N_4948);
xnor UO_30 (O_30,N_4991,N_4912);
nand UO_31 (O_31,N_4913,N_4942);
or UO_32 (O_32,N_4956,N_4963);
nor UO_33 (O_33,N_4926,N_4928);
or UO_34 (O_34,N_4969,N_4979);
and UO_35 (O_35,N_4927,N_4916);
nand UO_36 (O_36,N_4977,N_4941);
and UO_37 (O_37,N_4900,N_4968);
nand UO_38 (O_38,N_4999,N_4976);
and UO_39 (O_39,N_4982,N_4933);
nand UO_40 (O_40,N_4986,N_4958);
nor UO_41 (O_41,N_4923,N_4962);
and UO_42 (O_42,N_4980,N_4940);
xnor UO_43 (O_43,N_4998,N_4901);
nor UO_44 (O_44,N_4973,N_4964);
nand UO_45 (O_45,N_4946,N_4934);
nand UO_46 (O_46,N_4952,N_4943);
nand UO_47 (O_47,N_4914,N_4987);
nand UO_48 (O_48,N_4955,N_4990);
or UO_49 (O_49,N_4954,N_4971);
nand UO_50 (O_50,N_4902,N_4936);
and UO_51 (O_51,N_4988,N_4929);
and UO_52 (O_52,N_4938,N_4933);
nor UO_53 (O_53,N_4957,N_4967);
nor UO_54 (O_54,N_4982,N_4965);
nor UO_55 (O_55,N_4987,N_4967);
and UO_56 (O_56,N_4903,N_4999);
and UO_57 (O_57,N_4954,N_4960);
or UO_58 (O_58,N_4922,N_4957);
xnor UO_59 (O_59,N_4952,N_4993);
or UO_60 (O_60,N_4936,N_4944);
nor UO_61 (O_61,N_4948,N_4912);
or UO_62 (O_62,N_4921,N_4987);
and UO_63 (O_63,N_4954,N_4994);
and UO_64 (O_64,N_4977,N_4996);
nor UO_65 (O_65,N_4943,N_4939);
or UO_66 (O_66,N_4978,N_4916);
and UO_67 (O_67,N_4991,N_4915);
or UO_68 (O_68,N_4996,N_4952);
nor UO_69 (O_69,N_4943,N_4947);
or UO_70 (O_70,N_4965,N_4922);
or UO_71 (O_71,N_4985,N_4920);
xnor UO_72 (O_72,N_4913,N_4914);
or UO_73 (O_73,N_4926,N_4934);
nand UO_74 (O_74,N_4990,N_4991);
xor UO_75 (O_75,N_4965,N_4907);
nor UO_76 (O_76,N_4983,N_4951);
or UO_77 (O_77,N_4994,N_4987);
nand UO_78 (O_78,N_4948,N_4970);
nor UO_79 (O_79,N_4965,N_4917);
xnor UO_80 (O_80,N_4962,N_4957);
xor UO_81 (O_81,N_4929,N_4928);
nor UO_82 (O_82,N_4960,N_4966);
xnor UO_83 (O_83,N_4962,N_4928);
or UO_84 (O_84,N_4946,N_4985);
or UO_85 (O_85,N_4941,N_4963);
nand UO_86 (O_86,N_4931,N_4907);
xnor UO_87 (O_87,N_4947,N_4957);
or UO_88 (O_88,N_4910,N_4950);
or UO_89 (O_89,N_4919,N_4984);
or UO_90 (O_90,N_4996,N_4932);
nor UO_91 (O_91,N_4976,N_4945);
or UO_92 (O_92,N_4972,N_4922);
xnor UO_93 (O_93,N_4904,N_4950);
nor UO_94 (O_94,N_4928,N_4961);
and UO_95 (O_95,N_4956,N_4970);
nand UO_96 (O_96,N_4953,N_4975);
and UO_97 (O_97,N_4907,N_4945);
nand UO_98 (O_98,N_4924,N_4944);
or UO_99 (O_99,N_4959,N_4945);
or UO_100 (O_100,N_4978,N_4930);
nand UO_101 (O_101,N_4910,N_4905);
and UO_102 (O_102,N_4990,N_4919);
nand UO_103 (O_103,N_4939,N_4902);
nor UO_104 (O_104,N_4994,N_4901);
and UO_105 (O_105,N_4942,N_4906);
and UO_106 (O_106,N_4955,N_4965);
nor UO_107 (O_107,N_4958,N_4997);
xor UO_108 (O_108,N_4946,N_4942);
and UO_109 (O_109,N_4926,N_4932);
or UO_110 (O_110,N_4901,N_4953);
nand UO_111 (O_111,N_4926,N_4942);
or UO_112 (O_112,N_4914,N_4998);
nand UO_113 (O_113,N_4916,N_4956);
and UO_114 (O_114,N_4907,N_4989);
nand UO_115 (O_115,N_4995,N_4913);
nor UO_116 (O_116,N_4958,N_4967);
and UO_117 (O_117,N_4975,N_4980);
xor UO_118 (O_118,N_4917,N_4977);
and UO_119 (O_119,N_4989,N_4978);
or UO_120 (O_120,N_4931,N_4948);
and UO_121 (O_121,N_4935,N_4987);
nor UO_122 (O_122,N_4990,N_4962);
and UO_123 (O_123,N_4935,N_4989);
xor UO_124 (O_124,N_4995,N_4961);
nor UO_125 (O_125,N_4981,N_4998);
nor UO_126 (O_126,N_4917,N_4932);
or UO_127 (O_127,N_4905,N_4937);
xor UO_128 (O_128,N_4902,N_4990);
and UO_129 (O_129,N_4952,N_4992);
and UO_130 (O_130,N_4957,N_4945);
or UO_131 (O_131,N_4990,N_4958);
and UO_132 (O_132,N_4950,N_4968);
xor UO_133 (O_133,N_4963,N_4948);
nor UO_134 (O_134,N_4926,N_4981);
nor UO_135 (O_135,N_4927,N_4951);
or UO_136 (O_136,N_4991,N_4905);
nor UO_137 (O_137,N_4936,N_4971);
and UO_138 (O_138,N_4916,N_4913);
xnor UO_139 (O_139,N_4956,N_4945);
or UO_140 (O_140,N_4989,N_4999);
or UO_141 (O_141,N_4948,N_4946);
nor UO_142 (O_142,N_4950,N_4930);
xnor UO_143 (O_143,N_4964,N_4972);
or UO_144 (O_144,N_4941,N_4940);
xnor UO_145 (O_145,N_4919,N_4910);
nor UO_146 (O_146,N_4972,N_4925);
or UO_147 (O_147,N_4991,N_4923);
or UO_148 (O_148,N_4960,N_4990);
or UO_149 (O_149,N_4901,N_4992);
nand UO_150 (O_150,N_4923,N_4976);
nand UO_151 (O_151,N_4999,N_4907);
and UO_152 (O_152,N_4931,N_4994);
or UO_153 (O_153,N_4938,N_4944);
xnor UO_154 (O_154,N_4953,N_4995);
nor UO_155 (O_155,N_4947,N_4998);
and UO_156 (O_156,N_4971,N_4938);
nor UO_157 (O_157,N_4945,N_4927);
nand UO_158 (O_158,N_4958,N_4937);
and UO_159 (O_159,N_4916,N_4905);
and UO_160 (O_160,N_4985,N_4982);
nand UO_161 (O_161,N_4997,N_4945);
or UO_162 (O_162,N_4928,N_4911);
nor UO_163 (O_163,N_4976,N_4905);
or UO_164 (O_164,N_4966,N_4941);
nor UO_165 (O_165,N_4910,N_4971);
nand UO_166 (O_166,N_4927,N_4913);
and UO_167 (O_167,N_4983,N_4990);
nor UO_168 (O_168,N_4992,N_4916);
or UO_169 (O_169,N_4907,N_4921);
or UO_170 (O_170,N_4998,N_4974);
nor UO_171 (O_171,N_4955,N_4918);
and UO_172 (O_172,N_4970,N_4967);
or UO_173 (O_173,N_4987,N_4927);
nand UO_174 (O_174,N_4983,N_4979);
nand UO_175 (O_175,N_4996,N_4944);
xor UO_176 (O_176,N_4957,N_4937);
nor UO_177 (O_177,N_4960,N_4959);
and UO_178 (O_178,N_4904,N_4942);
nor UO_179 (O_179,N_4980,N_4957);
nor UO_180 (O_180,N_4965,N_4908);
xor UO_181 (O_181,N_4927,N_4964);
nand UO_182 (O_182,N_4929,N_4922);
or UO_183 (O_183,N_4973,N_4924);
nand UO_184 (O_184,N_4989,N_4948);
or UO_185 (O_185,N_4920,N_4988);
or UO_186 (O_186,N_4961,N_4934);
and UO_187 (O_187,N_4934,N_4921);
xor UO_188 (O_188,N_4912,N_4945);
or UO_189 (O_189,N_4968,N_4932);
or UO_190 (O_190,N_4908,N_4924);
and UO_191 (O_191,N_4911,N_4902);
xor UO_192 (O_192,N_4902,N_4988);
nand UO_193 (O_193,N_4976,N_4998);
nand UO_194 (O_194,N_4946,N_4945);
nand UO_195 (O_195,N_4923,N_4980);
nand UO_196 (O_196,N_4908,N_4919);
nand UO_197 (O_197,N_4985,N_4999);
or UO_198 (O_198,N_4950,N_4913);
nand UO_199 (O_199,N_4977,N_4961);
and UO_200 (O_200,N_4995,N_4945);
and UO_201 (O_201,N_4958,N_4979);
or UO_202 (O_202,N_4950,N_4933);
and UO_203 (O_203,N_4920,N_4963);
or UO_204 (O_204,N_4917,N_4956);
nor UO_205 (O_205,N_4974,N_4951);
nand UO_206 (O_206,N_4977,N_4978);
nor UO_207 (O_207,N_4913,N_4974);
nor UO_208 (O_208,N_4919,N_4927);
or UO_209 (O_209,N_4922,N_4925);
and UO_210 (O_210,N_4999,N_4919);
and UO_211 (O_211,N_4930,N_4963);
nand UO_212 (O_212,N_4991,N_4937);
or UO_213 (O_213,N_4962,N_4913);
or UO_214 (O_214,N_4998,N_4989);
nand UO_215 (O_215,N_4954,N_4925);
xnor UO_216 (O_216,N_4929,N_4926);
nand UO_217 (O_217,N_4909,N_4960);
and UO_218 (O_218,N_4906,N_4915);
or UO_219 (O_219,N_4924,N_4963);
nand UO_220 (O_220,N_4920,N_4912);
or UO_221 (O_221,N_4937,N_4962);
and UO_222 (O_222,N_4945,N_4934);
or UO_223 (O_223,N_4968,N_4975);
nor UO_224 (O_224,N_4986,N_4950);
and UO_225 (O_225,N_4998,N_4924);
nor UO_226 (O_226,N_4984,N_4945);
nand UO_227 (O_227,N_4909,N_4994);
and UO_228 (O_228,N_4924,N_4984);
or UO_229 (O_229,N_4998,N_4910);
or UO_230 (O_230,N_4915,N_4966);
nand UO_231 (O_231,N_4930,N_4990);
nand UO_232 (O_232,N_4936,N_4927);
and UO_233 (O_233,N_4959,N_4938);
or UO_234 (O_234,N_4923,N_4999);
or UO_235 (O_235,N_4957,N_4925);
nand UO_236 (O_236,N_4901,N_4915);
or UO_237 (O_237,N_4953,N_4915);
nand UO_238 (O_238,N_4912,N_4965);
nand UO_239 (O_239,N_4979,N_4933);
nand UO_240 (O_240,N_4983,N_4932);
nor UO_241 (O_241,N_4984,N_4944);
xor UO_242 (O_242,N_4903,N_4973);
and UO_243 (O_243,N_4968,N_4928);
and UO_244 (O_244,N_4900,N_4987);
nand UO_245 (O_245,N_4988,N_4908);
nand UO_246 (O_246,N_4970,N_4952);
nand UO_247 (O_247,N_4932,N_4924);
or UO_248 (O_248,N_4972,N_4963);
nor UO_249 (O_249,N_4988,N_4970);
and UO_250 (O_250,N_4985,N_4934);
and UO_251 (O_251,N_4963,N_4969);
nor UO_252 (O_252,N_4933,N_4987);
and UO_253 (O_253,N_4971,N_4953);
and UO_254 (O_254,N_4932,N_4908);
xnor UO_255 (O_255,N_4908,N_4981);
nor UO_256 (O_256,N_4937,N_4923);
or UO_257 (O_257,N_4903,N_4933);
xor UO_258 (O_258,N_4908,N_4975);
and UO_259 (O_259,N_4918,N_4920);
or UO_260 (O_260,N_4920,N_4909);
nand UO_261 (O_261,N_4962,N_4916);
xor UO_262 (O_262,N_4970,N_4969);
nand UO_263 (O_263,N_4926,N_4958);
xnor UO_264 (O_264,N_4928,N_4989);
xor UO_265 (O_265,N_4913,N_4957);
nor UO_266 (O_266,N_4902,N_4998);
nand UO_267 (O_267,N_4979,N_4954);
and UO_268 (O_268,N_4946,N_4980);
nand UO_269 (O_269,N_4951,N_4902);
and UO_270 (O_270,N_4998,N_4931);
nand UO_271 (O_271,N_4957,N_4994);
nand UO_272 (O_272,N_4942,N_4979);
and UO_273 (O_273,N_4964,N_4903);
or UO_274 (O_274,N_4932,N_4981);
nand UO_275 (O_275,N_4954,N_4933);
xor UO_276 (O_276,N_4947,N_4976);
and UO_277 (O_277,N_4922,N_4959);
nor UO_278 (O_278,N_4945,N_4935);
xor UO_279 (O_279,N_4901,N_4910);
xor UO_280 (O_280,N_4939,N_4945);
nand UO_281 (O_281,N_4904,N_4994);
nand UO_282 (O_282,N_4930,N_4972);
nor UO_283 (O_283,N_4911,N_4942);
nand UO_284 (O_284,N_4991,N_4954);
and UO_285 (O_285,N_4990,N_4946);
and UO_286 (O_286,N_4967,N_4922);
nand UO_287 (O_287,N_4940,N_4931);
and UO_288 (O_288,N_4934,N_4973);
nor UO_289 (O_289,N_4992,N_4934);
or UO_290 (O_290,N_4989,N_4953);
or UO_291 (O_291,N_4933,N_4912);
and UO_292 (O_292,N_4941,N_4927);
xor UO_293 (O_293,N_4956,N_4926);
or UO_294 (O_294,N_4971,N_4908);
or UO_295 (O_295,N_4931,N_4939);
xor UO_296 (O_296,N_4927,N_4990);
or UO_297 (O_297,N_4930,N_4968);
nand UO_298 (O_298,N_4916,N_4986);
nor UO_299 (O_299,N_4900,N_4975);
and UO_300 (O_300,N_4900,N_4928);
or UO_301 (O_301,N_4937,N_4976);
or UO_302 (O_302,N_4999,N_4939);
and UO_303 (O_303,N_4991,N_4928);
nor UO_304 (O_304,N_4922,N_4995);
xor UO_305 (O_305,N_4930,N_4934);
nand UO_306 (O_306,N_4943,N_4946);
nand UO_307 (O_307,N_4975,N_4954);
nor UO_308 (O_308,N_4946,N_4978);
or UO_309 (O_309,N_4910,N_4981);
and UO_310 (O_310,N_4974,N_4969);
nor UO_311 (O_311,N_4999,N_4932);
and UO_312 (O_312,N_4925,N_4975);
xnor UO_313 (O_313,N_4937,N_4919);
xnor UO_314 (O_314,N_4971,N_4919);
or UO_315 (O_315,N_4960,N_4995);
and UO_316 (O_316,N_4990,N_4965);
and UO_317 (O_317,N_4974,N_4971);
or UO_318 (O_318,N_4943,N_4954);
or UO_319 (O_319,N_4954,N_4903);
xnor UO_320 (O_320,N_4929,N_4932);
nor UO_321 (O_321,N_4959,N_4919);
or UO_322 (O_322,N_4922,N_4906);
or UO_323 (O_323,N_4921,N_4956);
or UO_324 (O_324,N_4939,N_4956);
nand UO_325 (O_325,N_4991,N_4989);
nor UO_326 (O_326,N_4925,N_4993);
and UO_327 (O_327,N_4996,N_4989);
nor UO_328 (O_328,N_4940,N_4989);
and UO_329 (O_329,N_4959,N_4966);
nor UO_330 (O_330,N_4911,N_4982);
nand UO_331 (O_331,N_4989,N_4946);
nand UO_332 (O_332,N_4931,N_4992);
nor UO_333 (O_333,N_4912,N_4988);
and UO_334 (O_334,N_4908,N_4916);
and UO_335 (O_335,N_4986,N_4949);
or UO_336 (O_336,N_4979,N_4902);
and UO_337 (O_337,N_4976,N_4902);
and UO_338 (O_338,N_4982,N_4935);
nand UO_339 (O_339,N_4981,N_4918);
or UO_340 (O_340,N_4906,N_4989);
nor UO_341 (O_341,N_4929,N_4914);
xor UO_342 (O_342,N_4995,N_4958);
nor UO_343 (O_343,N_4907,N_4966);
or UO_344 (O_344,N_4983,N_4984);
or UO_345 (O_345,N_4945,N_4915);
xnor UO_346 (O_346,N_4964,N_4934);
and UO_347 (O_347,N_4919,N_4931);
and UO_348 (O_348,N_4930,N_4949);
or UO_349 (O_349,N_4992,N_4953);
nand UO_350 (O_350,N_4924,N_4958);
and UO_351 (O_351,N_4983,N_4994);
nor UO_352 (O_352,N_4982,N_4943);
or UO_353 (O_353,N_4923,N_4916);
or UO_354 (O_354,N_4974,N_4904);
and UO_355 (O_355,N_4932,N_4967);
and UO_356 (O_356,N_4996,N_4909);
and UO_357 (O_357,N_4900,N_4980);
xnor UO_358 (O_358,N_4970,N_4929);
or UO_359 (O_359,N_4906,N_4997);
or UO_360 (O_360,N_4959,N_4915);
nand UO_361 (O_361,N_4976,N_4914);
or UO_362 (O_362,N_4913,N_4992);
nor UO_363 (O_363,N_4994,N_4999);
nand UO_364 (O_364,N_4925,N_4958);
and UO_365 (O_365,N_4902,N_4904);
and UO_366 (O_366,N_4922,N_4955);
xnor UO_367 (O_367,N_4960,N_4927);
xor UO_368 (O_368,N_4907,N_4912);
or UO_369 (O_369,N_4989,N_4931);
or UO_370 (O_370,N_4919,N_4968);
xnor UO_371 (O_371,N_4955,N_4981);
nor UO_372 (O_372,N_4941,N_4967);
xor UO_373 (O_373,N_4946,N_4905);
or UO_374 (O_374,N_4921,N_4989);
nor UO_375 (O_375,N_4902,N_4986);
nand UO_376 (O_376,N_4991,N_4918);
nand UO_377 (O_377,N_4938,N_4925);
nand UO_378 (O_378,N_4936,N_4979);
and UO_379 (O_379,N_4901,N_4975);
nor UO_380 (O_380,N_4997,N_4990);
or UO_381 (O_381,N_4978,N_4998);
nor UO_382 (O_382,N_4920,N_4955);
nand UO_383 (O_383,N_4983,N_4939);
xor UO_384 (O_384,N_4918,N_4925);
and UO_385 (O_385,N_4905,N_4940);
and UO_386 (O_386,N_4949,N_4984);
nand UO_387 (O_387,N_4913,N_4953);
xor UO_388 (O_388,N_4916,N_4959);
nor UO_389 (O_389,N_4978,N_4909);
or UO_390 (O_390,N_4973,N_4959);
nor UO_391 (O_391,N_4993,N_4900);
nor UO_392 (O_392,N_4962,N_4906);
or UO_393 (O_393,N_4912,N_4925);
and UO_394 (O_394,N_4934,N_4908);
nor UO_395 (O_395,N_4917,N_4946);
nand UO_396 (O_396,N_4950,N_4947);
and UO_397 (O_397,N_4922,N_4982);
or UO_398 (O_398,N_4939,N_4971);
xor UO_399 (O_399,N_4962,N_4944);
and UO_400 (O_400,N_4900,N_4955);
and UO_401 (O_401,N_4937,N_4975);
or UO_402 (O_402,N_4952,N_4962);
nand UO_403 (O_403,N_4915,N_4954);
nor UO_404 (O_404,N_4985,N_4971);
or UO_405 (O_405,N_4939,N_4982);
nand UO_406 (O_406,N_4954,N_4936);
or UO_407 (O_407,N_4935,N_4922);
nor UO_408 (O_408,N_4996,N_4910);
or UO_409 (O_409,N_4977,N_4903);
and UO_410 (O_410,N_4976,N_4978);
nand UO_411 (O_411,N_4980,N_4951);
nor UO_412 (O_412,N_4982,N_4924);
and UO_413 (O_413,N_4977,N_4940);
or UO_414 (O_414,N_4923,N_4961);
or UO_415 (O_415,N_4991,N_4933);
or UO_416 (O_416,N_4949,N_4989);
nor UO_417 (O_417,N_4943,N_4907);
nand UO_418 (O_418,N_4959,N_4902);
and UO_419 (O_419,N_4968,N_4952);
nand UO_420 (O_420,N_4936,N_4900);
and UO_421 (O_421,N_4924,N_4917);
nor UO_422 (O_422,N_4960,N_4904);
and UO_423 (O_423,N_4927,N_4915);
and UO_424 (O_424,N_4957,N_4956);
or UO_425 (O_425,N_4976,N_4931);
nor UO_426 (O_426,N_4912,N_4977);
nor UO_427 (O_427,N_4941,N_4969);
xor UO_428 (O_428,N_4904,N_4935);
nand UO_429 (O_429,N_4980,N_4908);
nor UO_430 (O_430,N_4936,N_4961);
nand UO_431 (O_431,N_4996,N_4966);
and UO_432 (O_432,N_4989,N_4981);
or UO_433 (O_433,N_4913,N_4948);
nor UO_434 (O_434,N_4901,N_4932);
and UO_435 (O_435,N_4919,N_4945);
nor UO_436 (O_436,N_4936,N_4945);
and UO_437 (O_437,N_4907,N_4990);
nand UO_438 (O_438,N_4962,N_4999);
nand UO_439 (O_439,N_4965,N_4958);
nor UO_440 (O_440,N_4927,N_4959);
nand UO_441 (O_441,N_4931,N_4934);
and UO_442 (O_442,N_4939,N_4962);
or UO_443 (O_443,N_4931,N_4957);
xnor UO_444 (O_444,N_4985,N_4954);
or UO_445 (O_445,N_4974,N_4942);
nor UO_446 (O_446,N_4907,N_4947);
and UO_447 (O_447,N_4931,N_4967);
and UO_448 (O_448,N_4965,N_4902);
nor UO_449 (O_449,N_4951,N_4977);
nor UO_450 (O_450,N_4998,N_4943);
nor UO_451 (O_451,N_4945,N_4979);
nand UO_452 (O_452,N_4920,N_4996);
and UO_453 (O_453,N_4993,N_4932);
nor UO_454 (O_454,N_4978,N_4961);
nand UO_455 (O_455,N_4922,N_4940);
xnor UO_456 (O_456,N_4910,N_4992);
nor UO_457 (O_457,N_4975,N_4941);
nor UO_458 (O_458,N_4972,N_4981);
nand UO_459 (O_459,N_4911,N_4946);
nand UO_460 (O_460,N_4964,N_4908);
nand UO_461 (O_461,N_4945,N_4986);
nor UO_462 (O_462,N_4964,N_4920);
or UO_463 (O_463,N_4951,N_4936);
or UO_464 (O_464,N_4904,N_4903);
nor UO_465 (O_465,N_4918,N_4951);
or UO_466 (O_466,N_4911,N_4950);
nor UO_467 (O_467,N_4932,N_4919);
and UO_468 (O_468,N_4915,N_4949);
nand UO_469 (O_469,N_4968,N_4913);
and UO_470 (O_470,N_4945,N_4910);
or UO_471 (O_471,N_4971,N_4993);
nand UO_472 (O_472,N_4953,N_4986);
nand UO_473 (O_473,N_4977,N_4923);
and UO_474 (O_474,N_4961,N_4981);
or UO_475 (O_475,N_4911,N_4941);
and UO_476 (O_476,N_4986,N_4912);
and UO_477 (O_477,N_4965,N_4909);
and UO_478 (O_478,N_4964,N_4978);
and UO_479 (O_479,N_4904,N_4932);
or UO_480 (O_480,N_4973,N_4951);
xor UO_481 (O_481,N_4938,N_4962);
nor UO_482 (O_482,N_4966,N_4904);
nor UO_483 (O_483,N_4969,N_4930);
and UO_484 (O_484,N_4936,N_4933);
nor UO_485 (O_485,N_4980,N_4991);
nor UO_486 (O_486,N_4901,N_4912);
nand UO_487 (O_487,N_4991,N_4960);
and UO_488 (O_488,N_4905,N_4958);
nor UO_489 (O_489,N_4996,N_4949);
nand UO_490 (O_490,N_4978,N_4963);
or UO_491 (O_491,N_4997,N_4928);
nor UO_492 (O_492,N_4988,N_4918);
or UO_493 (O_493,N_4938,N_4951);
and UO_494 (O_494,N_4997,N_4926);
nand UO_495 (O_495,N_4939,N_4926);
and UO_496 (O_496,N_4909,N_4973);
nand UO_497 (O_497,N_4985,N_4901);
nand UO_498 (O_498,N_4921,N_4908);
or UO_499 (O_499,N_4978,N_4917);
and UO_500 (O_500,N_4969,N_4919);
and UO_501 (O_501,N_4970,N_4914);
or UO_502 (O_502,N_4936,N_4904);
nor UO_503 (O_503,N_4924,N_4991);
and UO_504 (O_504,N_4987,N_4948);
xor UO_505 (O_505,N_4935,N_4979);
nor UO_506 (O_506,N_4997,N_4934);
and UO_507 (O_507,N_4932,N_4906);
nand UO_508 (O_508,N_4913,N_4938);
nor UO_509 (O_509,N_4937,N_4992);
or UO_510 (O_510,N_4998,N_4970);
nand UO_511 (O_511,N_4929,N_4935);
or UO_512 (O_512,N_4959,N_4981);
xor UO_513 (O_513,N_4970,N_4999);
nor UO_514 (O_514,N_4930,N_4917);
xnor UO_515 (O_515,N_4969,N_4917);
or UO_516 (O_516,N_4981,N_4976);
nor UO_517 (O_517,N_4964,N_4911);
or UO_518 (O_518,N_4929,N_4910);
nor UO_519 (O_519,N_4996,N_4950);
nand UO_520 (O_520,N_4902,N_4948);
nor UO_521 (O_521,N_4986,N_4952);
nor UO_522 (O_522,N_4987,N_4910);
nand UO_523 (O_523,N_4904,N_4954);
and UO_524 (O_524,N_4942,N_4982);
nor UO_525 (O_525,N_4981,N_4988);
nor UO_526 (O_526,N_4963,N_4954);
nand UO_527 (O_527,N_4900,N_4951);
or UO_528 (O_528,N_4970,N_4930);
or UO_529 (O_529,N_4938,N_4995);
nand UO_530 (O_530,N_4914,N_4936);
nand UO_531 (O_531,N_4970,N_4944);
nand UO_532 (O_532,N_4993,N_4986);
or UO_533 (O_533,N_4916,N_4920);
nand UO_534 (O_534,N_4905,N_4913);
or UO_535 (O_535,N_4977,N_4952);
or UO_536 (O_536,N_4929,N_4918);
or UO_537 (O_537,N_4953,N_4939);
and UO_538 (O_538,N_4986,N_4907);
or UO_539 (O_539,N_4921,N_4969);
nand UO_540 (O_540,N_4995,N_4900);
nor UO_541 (O_541,N_4928,N_4967);
nand UO_542 (O_542,N_4952,N_4951);
and UO_543 (O_543,N_4971,N_4906);
nor UO_544 (O_544,N_4963,N_4903);
nor UO_545 (O_545,N_4986,N_4971);
nor UO_546 (O_546,N_4975,N_4926);
nand UO_547 (O_547,N_4947,N_4914);
nand UO_548 (O_548,N_4906,N_4933);
and UO_549 (O_549,N_4995,N_4924);
or UO_550 (O_550,N_4919,N_4986);
xor UO_551 (O_551,N_4932,N_4928);
nand UO_552 (O_552,N_4997,N_4987);
xnor UO_553 (O_553,N_4939,N_4934);
nand UO_554 (O_554,N_4977,N_4921);
or UO_555 (O_555,N_4936,N_4906);
or UO_556 (O_556,N_4971,N_4967);
and UO_557 (O_557,N_4981,N_4966);
nor UO_558 (O_558,N_4915,N_4922);
nor UO_559 (O_559,N_4941,N_4950);
and UO_560 (O_560,N_4991,N_4995);
or UO_561 (O_561,N_4967,N_4946);
and UO_562 (O_562,N_4988,N_4903);
nor UO_563 (O_563,N_4924,N_4937);
and UO_564 (O_564,N_4957,N_4914);
nand UO_565 (O_565,N_4908,N_4942);
nand UO_566 (O_566,N_4914,N_4918);
and UO_567 (O_567,N_4990,N_4945);
or UO_568 (O_568,N_4927,N_4956);
nand UO_569 (O_569,N_4964,N_4991);
nor UO_570 (O_570,N_4939,N_4913);
nand UO_571 (O_571,N_4902,N_4917);
and UO_572 (O_572,N_4903,N_4934);
nand UO_573 (O_573,N_4927,N_4904);
nand UO_574 (O_574,N_4995,N_4916);
and UO_575 (O_575,N_4989,N_4913);
or UO_576 (O_576,N_4989,N_4958);
xor UO_577 (O_577,N_4941,N_4973);
nor UO_578 (O_578,N_4911,N_4987);
nand UO_579 (O_579,N_4903,N_4925);
or UO_580 (O_580,N_4979,N_4926);
and UO_581 (O_581,N_4922,N_4939);
or UO_582 (O_582,N_4938,N_4978);
and UO_583 (O_583,N_4904,N_4916);
nor UO_584 (O_584,N_4926,N_4925);
and UO_585 (O_585,N_4929,N_4924);
nand UO_586 (O_586,N_4930,N_4903);
nor UO_587 (O_587,N_4963,N_4949);
and UO_588 (O_588,N_4901,N_4960);
nor UO_589 (O_589,N_4978,N_4979);
and UO_590 (O_590,N_4901,N_4926);
xor UO_591 (O_591,N_4926,N_4957);
nand UO_592 (O_592,N_4917,N_4906);
nor UO_593 (O_593,N_4915,N_4956);
or UO_594 (O_594,N_4928,N_4916);
nor UO_595 (O_595,N_4984,N_4961);
or UO_596 (O_596,N_4919,N_4993);
nor UO_597 (O_597,N_4948,N_4971);
nand UO_598 (O_598,N_4935,N_4940);
and UO_599 (O_599,N_4901,N_4951);
nand UO_600 (O_600,N_4978,N_4991);
nand UO_601 (O_601,N_4958,N_4957);
nand UO_602 (O_602,N_4980,N_4910);
or UO_603 (O_603,N_4952,N_4905);
and UO_604 (O_604,N_4919,N_4981);
and UO_605 (O_605,N_4951,N_4997);
and UO_606 (O_606,N_4935,N_4965);
or UO_607 (O_607,N_4932,N_4995);
nor UO_608 (O_608,N_4951,N_4917);
nand UO_609 (O_609,N_4968,N_4944);
or UO_610 (O_610,N_4904,N_4933);
nor UO_611 (O_611,N_4968,N_4961);
or UO_612 (O_612,N_4944,N_4997);
nand UO_613 (O_613,N_4952,N_4922);
and UO_614 (O_614,N_4968,N_4949);
and UO_615 (O_615,N_4963,N_4926);
nor UO_616 (O_616,N_4949,N_4929);
nand UO_617 (O_617,N_4985,N_4994);
or UO_618 (O_618,N_4922,N_4971);
and UO_619 (O_619,N_4932,N_4966);
nand UO_620 (O_620,N_4916,N_4999);
and UO_621 (O_621,N_4986,N_4973);
nor UO_622 (O_622,N_4904,N_4937);
nor UO_623 (O_623,N_4975,N_4916);
nand UO_624 (O_624,N_4967,N_4943);
or UO_625 (O_625,N_4946,N_4914);
nand UO_626 (O_626,N_4926,N_4978);
nor UO_627 (O_627,N_4907,N_4978);
nor UO_628 (O_628,N_4903,N_4924);
xor UO_629 (O_629,N_4977,N_4979);
and UO_630 (O_630,N_4937,N_4954);
nor UO_631 (O_631,N_4998,N_4938);
nand UO_632 (O_632,N_4957,N_4921);
xor UO_633 (O_633,N_4930,N_4946);
or UO_634 (O_634,N_4972,N_4949);
and UO_635 (O_635,N_4951,N_4909);
nor UO_636 (O_636,N_4961,N_4974);
nor UO_637 (O_637,N_4900,N_4957);
xnor UO_638 (O_638,N_4924,N_4911);
nand UO_639 (O_639,N_4943,N_4962);
nor UO_640 (O_640,N_4964,N_4984);
and UO_641 (O_641,N_4940,N_4967);
nor UO_642 (O_642,N_4900,N_4910);
or UO_643 (O_643,N_4977,N_4990);
or UO_644 (O_644,N_4993,N_4907);
and UO_645 (O_645,N_4962,N_4934);
and UO_646 (O_646,N_4968,N_4903);
nand UO_647 (O_647,N_4969,N_4947);
nor UO_648 (O_648,N_4964,N_4912);
nand UO_649 (O_649,N_4939,N_4910);
or UO_650 (O_650,N_4994,N_4988);
nand UO_651 (O_651,N_4996,N_4933);
nand UO_652 (O_652,N_4975,N_4934);
and UO_653 (O_653,N_4978,N_4947);
nor UO_654 (O_654,N_4999,N_4902);
nand UO_655 (O_655,N_4937,N_4927);
or UO_656 (O_656,N_4971,N_4916);
nor UO_657 (O_657,N_4923,N_4945);
or UO_658 (O_658,N_4962,N_4969);
or UO_659 (O_659,N_4966,N_4999);
nand UO_660 (O_660,N_4980,N_4947);
nor UO_661 (O_661,N_4948,N_4990);
nor UO_662 (O_662,N_4941,N_4912);
nor UO_663 (O_663,N_4981,N_4937);
and UO_664 (O_664,N_4968,N_4974);
nand UO_665 (O_665,N_4939,N_4908);
and UO_666 (O_666,N_4905,N_4959);
or UO_667 (O_667,N_4973,N_4953);
or UO_668 (O_668,N_4996,N_4964);
nor UO_669 (O_669,N_4996,N_4901);
nand UO_670 (O_670,N_4945,N_4991);
nand UO_671 (O_671,N_4988,N_4925);
nor UO_672 (O_672,N_4915,N_4967);
nand UO_673 (O_673,N_4961,N_4904);
nand UO_674 (O_674,N_4904,N_4992);
nor UO_675 (O_675,N_4911,N_4914);
nor UO_676 (O_676,N_4962,N_4903);
and UO_677 (O_677,N_4955,N_4902);
and UO_678 (O_678,N_4921,N_4928);
nor UO_679 (O_679,N_4962,N_4951);
nor UO_680 (O_680,N_4906,N_4902);
or UO_681 (O_681,N_4981,N_4923);
or UO_682 (O_682,N_4917,N_4963);
nor UO_683 (O_683,N_4903,N_4947);
nand UO_684 (O_684,N_4963,N_4979);
and UO_685 (O_685,N_4917,N_4971);
nor UO_686 (O_686,N_4952,N_4934);
nor UO_687 (O_687,N_4923,N_4986);
nand UO_688 (O_688,N_4969,N_4909);
nand UO_689 (O_689,N_4980,N_4966);
nor UO_690 (O_690,N_4947,N_4920);
nor UO_691 (O_691,N_4922,N_4948);
or UO_692 (O_692,N_4903,N_4981);
and UO_693 (O_693,N_4923,N_4973);
nand UO_694 (O_694,N_4953,N_4947);
and UO_695 (O_695,N_4988,N_4955);
or UO_696 (O_696,N_4918,N_4923);
nand UO_697 (O_697,N_4982,N_4944);
and UO_698 (O_698,N_4963,N_4915);
nand UO_699 (O_699,N_4936,N_4996);
or UO_700 (O_700,N_4946,N_4962);
nor UO_701 (O_701,N_4977,N_4950);
nand UO_702 (O_702,N_4962,N_4914);
nand UO_703 (O_703,N_4909,N_4933);
and UO_704 (O_704,N_4949,N_4941);
or UO_705 (O_705,N_4972,N_4928);
or UO_706 (O_706,N_4983,N_4998);
nand UO_707 (O_707,N_4942,N_4917);
or UO_708 (O_708,N_4918,N_4902);
and UO_709 (O_709,N_4956,N_4940);
or UO_710 (O_710,N_4996,N_4979);
and UO_711 (O_711,N_4901,N_4903);
and UO_712 (O_712,N_4925,N_4973);
or UO_713 (O_713,N_4920,N_4951);
nand UO_714 (O_714,N_4924,N_4940);
xor UO_715 (O_715,N_4960,N_4920);
or UO_716 (O_716,N_4959,N_4988);
nand UO_717 (O_717,N_4973,N_4904);
nand UO_718 (O_718,N_4930,N_4993);
nand UO_719 (O_719,N_4975,N_4932);
or UO_720 (O_720,N_4995,N_4993);
and UO_721 (O_721,N_4926,N_4922);
or UO_722 (O_722,N_4967,N_4984);
nand UO_723 (O_723,N_4952,N_4982);
or UO_724 (O_724,N_4971,N_4975);
and UO_725 (O_725,N_4995,N_4915);
or UO_726 (O_726,N_4962,N_4909);
nand UO_727 (O_727,N_4947,N_4964);
nor UO_728 (O_728,N_4987,N_4981);
nor UO_729 (O_729,N_4931,N_4956);
nor UO_730 (O_730,N_4992,N_4908);
nand UO_731 (O_731,N_4950,N_4912);
nor UO_732 (O_732,N_4951,N_4972);
nor UO_733 (O_733,N_4989,N_4977);
nand UO_734 (O_734,N_4904,N_4991);
nor UO_735 (O_735,N_4907,N_4940);
nor UO_736 (O_736,N_4997,N_4952);
or UO_737 (O_737,N_4909,N_4970);
xnor UO_738 (O_738,N_4976,N_4989);
nor UO_739 (O_739,N_4948,N_4982);
nor UO_740 (O_740,N_4956,N_4982);
and UO_741 (O_741,N_4979,N_4948);
or UO_742 (O_742,N_4922,N_4999);
and UO_743 (O_743,N_4906,N_4952);
nand UO_744 (O_744,N_4975,N_4935);
xnor UO_745 (O_745,N_4966,N_4954);
and UO_746 (O_746,N_4999,N_4904);
and UO_747 (O_747,N_4991,N_4999);
or UO_748 (O_748,N_4946,N_4974);
nor UO_749 (O_749,N_4935,N_4958);
nor UO_750 (O_750,N_4998,N_4961);
and UO_751 (O_751,N_4951,N_4932);
or UO_752 (O_752,N_4968,N_4934);
nand UO_753 (O_753,N_4978,N_4956);
or UO_754 (O_754,N_4935,N_4933);
xnor UO_755 (O_755,N_4982,N_4928);
and UO_756 (O_756,N_4993,N_4970);
and UO_757 (O_757,N_4909,N_4945);
nor UO_758 (O_758,N_4941,N_4929);
xor UO_759 (O_759,N_4921,N_4961);
nor UO_760 (O_760,N_4955,N_4957);
nand UO_761 (O_761,N_4962,N_4987);
nor UO_762 (O_762,N_4956,N_4935);
and UO_763 (O_763,N_4903,N_4976);
and UO_764 (O_764,N_4969,N_4951);
or UO_765 (O_765,N_4997,N_4921);
and UO_766 (O_766,N_4926,N_4912);
nor UO_767 (O_767,N_4966,N_4963);
and UO_768 (O_768,N_4904,N_4965);
or UO_769 (O_769,N_4903,N_4937);
nor UO_770 (O_770,N_4909,N_4937);
nor UO_771 (O_771,N_4967,N_4960);
xnor UO_772 (O_772,N_4952,N_4973);
and UO_773 (O_773,N_4945,N_4913);
or UO_774 (O_774,N_4980,N_4979);
and UO_775 (O_775,N_4903,N_4912);
nand UO_776 (O_776,N_4917,N_4925);
nor UO_777 (O_777,N_4939,N_4947);
or UO_778 (O_778,N_4928,N_4930);
and UO_779 (O_779,N_4935,N_4937);
nor UO_780 (O_780,N_4900,N_4933);
and UO_781 (O_781,N_4979,N_4971);
or UO_782 (O_782,N_4961,N_4994);
or UO_783 (O_783,N_4956,N_4958);
nand UO_784 (O_784,N_4987,N_4946);
and UO_785 (O_785,N_4927,N_4970);
and UO_786 (O_786,N_4983,N_4910);
nand UO_787 (O_787,N_4911,N_4952);
and UO_788 (O_788,N_4970,N_4901);
nand UO_789 (O_789,N_4955,N_4931);
nand UO_790 (O_790,N_4975,N_4957);
nor UO_791 (O_791,N_4953,N_4958);
nor UO_792 (O_792,N_4904,N_4908);
and UO_793 (O_793,N_4994,N_4943);
and UO_794 (O_794,N_4937,N_4988);
nand UO_795 (O_795,N_4996,N_4904);
nor UO_796 (O_796,N_4943,N_4974);
nor UO_797 (O_797,N_4946,N_4952);
or UO_798 (O_798,N_4960,N_4923);
nand UO_799 (O_799,N_4941,N_4984);
and UO_800 (O_800,N_4979,N_4932);
and UO_801 (O_801,N_4944,N_4986);
nor UO_802 (O_802,N_4935,N_4953);
nand UO_803 (O_803,N_4908,N_4969);
or UO_804 (O_804,N_4994,N_4950);
nor UO_805 (O_805,N_4910,N_4917);
nor UO_806 (O_806,N_4944,N_4955);
xnor UO_807 (O_807,N_4914,N_4968);
nand UO_808 (O_808,N_4948,N_4942);
xor UO_809 (O_809,N_4929,N_4994);
and UO_810 (O_810,N_4979,N_4941);
nor UO_811 (O_811,N_4966,N_4988);
nand UO_812 (O_812,N_4998,N_4951);
and UO_813 (O_813,N_4918,N_4995);
nand UO_814 (O_814,N_4984,N_4954);
or UO_815 (O_815,N_4939,N_4952);
or UO_816 (O_816,N_4922,N_4908);
and UO_817 (O_817,N_4967,N_4948);
nor UO_818 (O_818,N_4987,N_4909);
nand UO_819 (O_819,N_4986,N_4965);
nor UO_820 (O_820,N_4990,N_4909);
nor UO_821 (O_821,N_4935,N_4970);
xnor UO_822 (O_822,N_4900,N_4941);
nor UO_823 (O_823,N_4928,N_4935);
xnor UO_824 (O_824,N_4981,N_4938);
nand UO_825 (O_825,N_4942,N_4934);
nor UO_826 (O_826,N_4997,N_4935);
or UO_827 (O_827,N_4923,N_4904);
nor UO_828 (O_828,N_4961,N_4915);
or UO_829 (O_829,N_4986,N_4946);
and UO_830 (O_830,N_4974,N_4914);
xnor UO_831 (O_831,N_4908,N_4911);
or UO_832 (O_832,N_4968,N_4981);
xor UO_833 (O_833,N_4903,N_4997);
or UO_834 (O_834,N_4989,N_4914);
and UO_835 (O_835,N_4953,N_4993);
or UO_836 (O_836,N_4966,N_4901);
or UO_837 (O_837,N_4906,N_4934);
nor UO_838 (O_838,N_4935,N_4968);
or UO_839 (O_839,N_4916,N_4914);
and UO_840 (O_840,N_4989,N_4994);
nand UO_841 (O_841,N_4914,N_4967);
nor UO_842 (O_842,N_4920,N_4950);
nand UO_843 (O_843,N_4906,N_4981);
nand UO_844 (O_844,N_4989,N_4927);
and UO_845 (O_845,N_4913,N_4921);
or UO_846 (O_846,N_4936,N_4901);
and UO_847 (O_847,N_4946,N_4982);
xor UO_848 (O_848,N_4913,N_4946);
nor UO_849 (O_849,N_4937,N_4946);
nand UO_850 (O_850,N_4917,N_4959);
nor UO_851 (O_851,N_4982,N_4972);
or UO_852 (O_852,N_4953,N_4997);
nor UO_853 (O_853,N_4902,N_4996);
xor UO_854 (O_854,N_4968,N_4993);
nor UO_855 (O_855,N_4954,N_4995);
xnor UO_856 (O_856,N_4934,N_4923);
or UO_857 (O_857,N_4924,N_4933);
and UO_858 (O_858,N_4931,N_4973);
or UO_859 (O_859,N_4965,N_4970);
nor UO_860 (O_860,N_4904,N_4912);
or UO_861 (O_861,N_4922,N_4969);
nand UO_862 (O_862,N_4902,N_4913);
or UO_863 (O_863,N_4909,N_4997);
nand UO_864 (O_864,N_4999,N_4929);
nor UO_865 (O_865,N_4902,N_4975);
and UO_866 (O_866,N_4985,N_4968);
nand UO_867 (O_867,N_4989,N_4934);
and UO_868 (O_868,N_4950,N_4900);
or UO_869 (O_869,N_4965,N_4943);
and UO_870 (O_870,N_4966,N_4951);
nor UO_871 (O_871,N_4938,N_4901);
nand UO_872 (O_872,N_4904,N_4988);
or UO_873 (O_873,N_4964,N_4979);
and UO_874 (O_874,N_4907,N_4918);
nand UO_875 (O_875,N_4975,N_4993);
or UO_876 (O_876,N_4985,N_4988);
nor UO_877 (O_877,N_4941,N_4972);
nor UO_878 (O_878,N_4928,N_4973);
nor UO_879 (O_879,N_4991,N_4982);
or UO_880 (O_880,N_4966,N_4990);
and UO_881 (O_881,N_4925,N_4930);
nand UO_882 (O_882,N_4974,N_4999);
and UO_883 (O_883,N_4920,N_4995);
nand UO_884 (O_884,N_4906,N_4972);
nand UO_885 (O_885,N_4948,N_4911);
or UO_886 (O_886,N_4920,N_4925);
nor UO_887 (O_887,N_4953,N_4912);
or UO_888 (O_888,N_4988,N_4919);
and UO_889 (O_889,N_4978,N_4937);
and UO_890 (O_890,N_4925,N_4937);
or UO_891 (O_891,N_4970,N_4938);
xnor UO_892 (O_892,N_4921,N_4990);
nand UO_893 (O_893,N_4911,N_4919);
and UO_894 (O_894,N_4968,N_4983);
nor UO_895 (O_895,N_4912,N_4918);
or UO_896 (O_896,N_4985,N_4997);
xor UO_897 (O_897,N_4917,N_4981);
and UO_898 (O_898,N_4979,N_4988);
and UO_899 (O_899,N_4983,N_4952);
or UO_900 (O_900,N_4933,N_4947);
and UO_901 (O_901,N_4985,N_4975);
nor UO_902 (O_902,N_4974,N_4903);
and UO_903 (O_903,N_4966,N_4992);
and UO_904 (O_904,N_4951,N_4934);
or UO_905 (O_905,N_4991,N_4900);
nand UO_906 (O_906,N_4997,N_4918);
nand UO_907 (O_907,N_4909,N_4992);
nand UO_908 (O_908,N_4931,N_4968);
nor UO_909 (O_909,N_4960,N_4929);
nand UO_910 (O_910,N_4974,N_4935);
nand UO_911 (O_911,N_4967,N_4993);
and UO_912 (O_912,N_4932,N_4964);
nand UO_913 (O_913,N_4987,N_4912);
nor UO_914 (O_914,N_4930,N_4922);
nand UO_915 (O_915,N_4944,N_4966);
xnor UO_916 (O_916,N_4938,N_4946);
or UO_917 (O_917,N_4905,N_4983);
nand UO_918 (O_918,N_4910,N_4902);
nor UO_919 (O_919,N_4946,N_4912);
nor UO_920 (O_920,N_4986,N_4976);
nor UO_921 (O_921,N_4915,N_4973);
nand UO_922 (O_922,N_4974,N_4917);
nor UO_923 (O_923,N_4993,N_4984);
or UO_924 (O_924,N_4972,N_4921);
nand UO_925 (O_925,N_4975,N_4942);
or UO_926 (O_926,N_4912,N_4959);
and UO_927 (O_927,N_4969,N_4933);
nor UO_928 (O_928,N_4924,N_4975);
or UO_929 (O_929,N_4943,N_4951);
or UO_930 (O_930,N_4996,N_4915);
and UO_931 (O_931,N_4987,N_4922);
xor UO_932 (O_932,N_4931,N_4962);
or UO_933 (O_933,N_4906,N_4926);
and UO_934 (O_934,N_4922,N_4901);
nand UO_935 (O_935,N_4936,N_4903);
nor UO_936 (O_936,N_4950,N_4987);
nand UO_937 (O_937,N_4991,N_4929);
or UO_938 (O_938,N_4904,N_4964);
xor UO_939 (O_939,N_4959,N_4969);
nor UO_940 (O_940,N_4967,N_4959);
nor UO_941 (O_941,N_4994,N_4905);
or UO_942 (O_942,N_4973,N_4966);
and UO_943 (O_943,N_4953,N_4929);
or UO_944 (O_944,N_4977,N_4927);
nand UO_945 (O_945,N_4943,N_4950);
nand UO_946 (O_946,N_4913,N_4910);
nand UO_947 (O_947,N_4973,N_4975);
nand UO_948 (O_948,N_4914,N_4927);
or UO_949 (O_949,N_4900,N_4908);
nor UO_950 (O_950,N_4999,N_4952);
nand UO_951 (O_951,N_4947,N_4923);
and UO_952 (O_952,N_4983,N_4925);
nor UO_953 (O_953,N_4967,N_4989);
or UO_954 (O_954,N_4936,N_4950);
or UO_955 (O_955,N_4915,N_4957);
and UO_956 (O_956,N_4923,N_4925);
or UO_957 (O_957,N_4983,N_4941);
nor UO_958 (O_958,N_4934,N_4941);
nor UO_959 (O_959,N_4937,N_4956);
nand UO_960 (O_960,N_4914,N_4921);
nand UO_961 (O_961,N_4973,N_4974);
and UO_962 (O_962,N_4987,N_4979);
nor UO_963 (O_963,N_4972,N_4944);
and UO_964 (O_964,N_4982,N_4905);
and UO_965 (O_965,N_4910,N_4914);
xnor UO_966 (O_966,N_4933,N_4964);
nor UO_967 (O_967,N_4911,N_4912);
and UO_968 (O_968,N_4981,N_4941);
and UO_969 (O_969,N_4902,N_4926);
nor UO_970 (O_970,N_4915,N_4944);
and UO_971 (O_971,N_4956,N_4946);
nand UO_972 (O_972,N_4936,N_4930);
and UO_973 (O_973,N_4995,N_4987);
or UO_974 (O_974,N_4988,N_4991);
nand UO_975 (O_975,N_4943,N_4985);
and UO_976 (O_976,N_4934,N_4936);
xor UO_977 (O_977,N_4970,N_4937);
nor UO_978 (O_978,N_4900,N_4932);
nor UO_979 (O_979,N_4927,N_4946);
or UO_980 (O_980,N_4908,N_4954);
or UO_981 (O_981,N_4969,N_4965);
xnor UO_982 (O_982,N_4992,N_4915);
and UO_983 (O_983,N_4964,N_4943);
nor UO_984 (O_984,N_4964,N_4937);
or UO_985 (O_985,N_4937,N_4906);
xnor UO_986 (O_986,N_4924,N_4954);
nor UO_987 (O_987,N_4903,N_4919);
xor UO_988 (O_988,N_4993,N_4965);
nand UO_989 (O_989,N_4920,N_4935);
or UO_990 (O_990,N_4926,N_4933);
or UO_991 (O_991,N_4984,N_4987);
or UO_992 (O_992,N_4997,N_4940);
or UO_993 (O_993,N_4933,N_4913);
and UO_994 (O_994,N_4970,N_4987);
or UO_995 (O_995,N_4968,N_4945);
nand UO_996 (O_996,N_4910,N_4968);
and UO_997 (O_997,N_4920,N_4962);
and UO_998 (O_998,N_4967,N_4903);
nand UO_999 (O_999,N_4967,N_4985);
endmodule