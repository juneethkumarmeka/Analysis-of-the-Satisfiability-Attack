module basic_3000_30000_3500_30_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_2820,In_1849);
nand U1 (N_1,In_1584,In_2249);
and U2 (N_2,In_2126,In_2074);
and U3 (N_3,In_959,In_731);
and U4 (N_4,In_304,In_1688);
and U5 (N_5,In_2322,In_2796);
nand U6 (N_6,In_1390,In_675);
nand U7 (N_7,In_2933,In_957);
or U8 (N_8,In_2951,In_1520);
xor U9 (N_9,In_605,In_1691);
or U10 (N_10,In_2399,In_2298);
xnor U11 (N_11,In_499,In_1434);
or U12 (N_12,In_1541,In_1542);
xor U13 (N_13,In_2413,In_1357);
and U14 (N_14,In_1954,In_295);
or U15 (N_15,In_2060,In_1415);
and U16 (N_16,In_589,In_880);
nand U17 (N_17,In_165,In_1306);
xnor U18 (N_18,In_1577,In_2116);
nand U19 (N_19,In_1414,In_1429);
or U20 (N_20,In_2523,In_1168);
nor U21 (N_21,In_1275,In_781);
nor U22 (N_22,In_1606,In_1955);
or U23 (N_23,In_824,In_1373);
and U24 (N_24,In_333,In_2783);
nor U25 (N_25,In_2401,In_2636);
or U26 (N_26,In_2115,In_2036);
nor U27 (N_27,In_2017,In_1165);
nand U28 (N_28,In_2473,In_1328);
xnor U29 (N_29,In_81,In_1486);
nand U30 (N_30,In_2346,In_106);
or U31 (N_31,In_2132,In_197);
xor U32 (N_32,In_2880,In_2078);
or U33 (N_33,In_2888,In_1968);
and U34 (N_34,In_1500,In_2133);
and U35 (N_35,In_2252,In_2700);
and U36 (N_36,In_500,In_621);
nand U37 (N_37,In_1387,In_782);
or U38 (N_38,In_1075,In_249);
xnor U39 (N_39,In_2858,In_2351);
or U40 (N_40,In_2824,In_1634);
xnor U41 (N_41,In_2819,In_1060);
or U42 (N_42,In_2665,In_2785);
nor U43 (N_43,In_554,In_1261);
nor U44 (N_44,In_2661,In_2635);
nand U45 (N_45,In_1527,In_1008);
nor U46 (N_46,In_267,In_1811);
nand U47 (N_47,In_1728,In_1488);
or U48 (N_48,In_209,In_1073);
nor U49 (N_49,In_1480,In_1413);
nor U50 (N_50,In_2216,In_2402);
or U51 (N_51,In_1124,In_1513);
or U52 (N_52,In_1462,In_828);
and U53 (N_53,In_882,In_1103);
or U54 (N_54,In_2678,In_212);
xor U55 (N_55,In_1842,In_1865);
nand U56 (N_56,In_1848,In_1810);
and U57 (N_57,In_737,In_437);
and U58 (N_58,In_2142,In_943);
nand U59 (N_59,In_1149,In_1230);
nor U60 (N_60,In_272,In_2258);
xnor U61 (N_61,In_1422,In_839);
nand U62 (N_62,In_74,In_922);
nor U63 (N_63,In_2039,In_139);
nand U64 (N_64,In_2681,In_2251);
nor U65 (N_65,In_1970,In_1337);
or U66 (N_66,In_1067,In_19);
and U67 (N_67,In_1160,In_2941);
nand U68 (N_68,In_486,In_2471);
nand U69 (N_69,In_1863,In_591);
nor U70 (N_70,In_2618,In_1166);
or U71 (N_71,In_125,In_2566);
or U72 (N_72,In_2580,In_1643);
and U73 (N_73,In_421,In_2000);
and U74 (N_74,In_2680,In_2312);
xor U75 (N_75,In_1719,In_2826);
nand U76 (N_76,In_1656,In_721);
nor U77 (N_77,In_169,In_681);
xor U78 (N_78,In_1635,In_211);
and U79 (N_79,In_1477,In_1494);
xnor U80 (N_80,In_1153,In_1806);
nor U81 (N_81,In_1538,In_1482);
xor U82 (N_82,In_448,In_2730);
xnor U83 (N_83,In_1769,In_301);
xnor U84 (N_84,In_2289,In_88);
and U85 (N_85,In_2877,In_524);
xnor U86 (N_86,In_2285,In_2350);
nor U87 (N_87,In_1670,In_692);
and U88 (N_88,In_963,In_2294);
or U89 (N_89,In_315,In_2179);
or U90 (N_90,In_2774,In_1304);
or U91 (N_91,In_2380,In_2794);
nand U92 (N_92,In_2172,In_729);
and U93 (N_93,In_567,In_1664);
xor U94 (N_94,In_1464,In_698);
and U95 (N_95,In_2588,In_473);
or U96 (N_96,In_1123,In_1498);
and U97 (N_97,In_2599,In_124);
nand U98 (N_98,In_2487,In_2182);
and U99 (N_99,In_1640,In_1547);
nor U100 (N_100,In_2746,In_2428);
nand U101 (N_101,In_2984,In_2845);
and U102 (N_102,In_493,In_2079);
and U103 (N_103,In_2367,In_2689);
xor U104 (N_104,In_2027,In_583);
or U105 (N_105,In_1095,In_2156);
nand U106 (N_106,In_2280,In_2099);
or U107 (N_107,In_735,In_2470);
nand U108 (N_108,In_2003,In_287);
nor U109 (N_109,In_649,In_1566);
xnor U110 (N_110,In_2159,In_1391);
or U111 (N_111,In_2989,In_2543);
or U112 (N_112,In_1199,In_2069);
and U113 (N_113,In_2419,In_1928);
or U114 (N_114,In_1809,In_2833);
or U115 (N_115,In_329,In_453);
or U116 (N_116,In_1181,In_2023);
and U117 (N_117,In_2461,In_1180);
and U118 (N_118,In_321,In_748);
or U119 (N_119,In_747,In_1394);
nand U120 (N_120,In_1545,In_1228);
xor U121 (N_121,In_2967,In_2477);
nor U122 (N_122,In_2277,In_2488);
or U123 (N_123,In_702,In_2331);
nand U124 (N_124,In_677,In_2670);
xnor U125 (N_125,In_2956,In_1476);
xor U126 (N_126,In_1558,In_1343);
xnor U127 (N_127,In_966,In_501);
nor U128 (N_128,In_2032,In_1771);
or U129 (N_129,In_1046,In_925);
nor U130 (N_130,In_1405,In_1033);
xnor U131 (N_131,In_2840,In_2708);
xor U132 (N_132,In_661,In_65);
nor U133 (N_133,In_878,In_98);
nand U134 (N_134,In_11,In_381);
nand U135 (N_135,In_2768,In_777);
nand U136 (N_136,In_162,In_862);
or U137 (N_137,In_1010,In_80);
xor U138 (N_138,In_1621,In_2579);
nor U139 (N_139,In_1729,In_995);
xor U140 (N_140,In_931,In_1854);
and U141 (N_141,In_474,In_1085);
nor U142 (N_142,In_544,In_248);
nor U143 (N_143,In_1447,In_2859);
xor U144 (N_144,In_2450,In_2482);
xor U145 (N_145,In_1556,In_1041);
nor U146 (N_146,In_285,In_2766);
or U147 (N_147,In_2398,In_2392);
nor U148 (N_148,In_2709,In_2609);
xor U149 (N_149,In_2047,In_999);
and U150 (N_150,In_879,In_1943);
nor U151 (N_151,In_2662,In_1052);
xor U152 (N_152,In_1990,In_35);
or U153 (N_153,In_1219,In_2653);
nor U154 (N_154,In_2757,In_1291);
or U155 (N_155,In_576,In_548);
xnor U156 (N_156,In_540,In_771);
and U157 (N_157,In_2717,In_2629);
xor U158 (N_158,In_872,In_160);
xnor U159 (N_159,In_1321,In_1758);
and U160 (N_160,In_1187,In_1690);
or U161 (N_161,In_93,In_2037);
and U162 (N_162,In_1828,In_1743);
xnor U163 (N_163,In_1053,In_2022);
or U164 (N_164,In_1280,In_2619);
and U165 (N_165,In_1175,In_2364);
and U166 (N_166,In_1302,In_2842);
xnor U167 (N_167,In_230,In_233);
nor U168 (N_168,In_1455,In_750);
nand U169 (N_169,In_1309,In_2677);
xor U170 (N_170,In_1750,In_1797);
nor U171 (N_171,In_519,In_2961);
and U172 (N_172,In_51,In_1616);
or U173 (N_173,In_1058,In_2712);
xnor U174 (N_174,In_1259,In_1964);
xnor U175 (N_175,In_316,In_2269);
nand U176 (N_176,In_708,In_306);
nor U177 (N_177,In_1649,In_108);
nor U178 (N_178,In_2065,In_1487);
or U179 (N_179,In_147,In_940);
nand U180 (N_180,In_2169,In_1214);
nand U181 (N_181,In_614,In_2589);
xnor U182 (N_182,In_1678,In_1379);
nand U183 (N_183,In_1277,In_2453);
and U184 (N_184,In_1960,In_1303);
nor U185 (N_185,In_2699,In_2046);
nor U186 (N_186,In_345,In_852);
nor U187 (N_187,In_517,In_2434);
nand U188 (N_188,In_514,In_161);
xnor U189 (N_189,In_525,In_1780);
nor U190 (N_190,In_1647,In_1091);
or U191 (N_191,In_559,In_1439);
and U192 (N_192,In_2034,In_1242);
and U193 (N_193,In_562,In_1665);
and U194 (N_194,In_293,In_1612);
or U195 (N_195,In_1300,In_754);
nand U196 (N_196,In_2658,In_1437);
xnor U197 (N_197,In_2632,In_893);
nand U198 (N_198,In_2863,In_1460);
and U199 (N_199,In_656,In_1114);
nand U200 (N_200,In_1004,In_1510);
nor U201 (N_201,In_1875,In_2535);
nand U202 (N_202,In_2314,In_53);
or U203 (N_203,In_2290,In_874);
nor U204 (N_204,In_2226,In_728);
nand U205 (N_205,In_2627,In_2528);
xnor U206 (N_206,In_810,In_1817);
xor U207 (N_207,In_1580,In_1233);
xnor U208 (N_208,In_898,In_2405);
and U209 (N_209,In_388,In_1697);
xnor U210 (N_210,In_2235,In_2024);
and U211 (N_211,In_2317,In_1217);
nand U212 (N_212,In_1912,In_1125);
nand U213 (N_213,In_842,In_330);
or U214 (N_214,In_217,In_783);
and U215 (N_215,In_1258,In_1006);
and U216 (N_216,In_1490,In_2239);
nand U217 (N_217,In_2253,In_1685);
or U218 (N_218,In_1001,In_14);
or U219 (N_219,In_1325,In_24);
and U220 (N_220,In_942,In_1013);
xor U221 (N_221,In_2009,In_706);
nand U222 (N_222,In_2763,In_1724);
and U223 (N_223,In_1398,In_1416);
xor U224 (N_224,In_2170,In_1804);
nor U225 (N_225,In_214,In_951);
nor U226 (N_226,In_2016,In_2546);
and U227 (N_227,In_1568,In_1938);
xnor U228 (N_228,In_276,In_2713);
xnor U229 (N_229,In_1430,In_1502);
xnor U230 (N_230,In_72,In_266);
xnor U231 (N_231,In_1533,In_1521);
and U232 (N_232,In_823,In_2431);
nor U233 (N_233,In_190,In_2098);
or U234 (N_234,In_1479,In_977);
or U235 (N_235,In_761,In_2687);
or U236 (N_236,In_1138,In_2202);
nand U237 (N_237,In_372,In_1076);
or U238 (N_238,In_699,In_353);
xor U239 (N_239,In_418,In_1549);
nand U240 (N_240,In_2043,In_2724);
or U241 (N_241,In_2640,In_1886);
xnor U242 (N_242,In_305,In_602);
or U243 (N_243,In_30,In_2166);
xnor U244 (N_244,In_2622,In_40);
nand U245 (N_245,In_617,In_2444);
xor U246 (N_246,In_323,In_1999);
or U247 (N_247,In_593,In_2574);
and U248 (N_248,In_2711,In_1497);
nor U249 (N_249,In_1748,In_1747);
and U250 (N_250,In_2534,In_2899);
and U251 (N_251,In_2381,In_2674);
and U252 (N_252,In_947,In_875);
nand U253 (N_253,In_2204,In_2209);
nand U254 (N_254,In_159,In_1056);
nand U255 (N_255,In_1826,In_1572);
nand U256 (N_256,In_1663,In_1680);
nor U257 (N_257,In_742,In_1965);
or U258 (N_258,In_773,In_670);
nor U259 (N_259,In_869,In_1911);
and U260 (N_260,In_447,In_1644);
nor U261 (N_261,In_84,In_806);
nand U262 (N_262,In_1475,In_779);
xnor U263 (N_263,In_521,In_1203);
nor U264 (N_264,In_1564,In_1446);
xor U265 (N_265,In_1902,In_269);
nor U266 (N_266,In_2917,In_983);
xnor U267 (N_267,In_1120,In_480);
nand U268 (N_268,In_1198,In_523);
nor U269 (N_269,In_2263,In_795);
nand U270 (N_270,In_1517,In_374);
nor U271 (N_271,In_686,In_1454);
nor U272 (N_272,In_759,In_90);
nor U273 (N_273,In_1236,In_2988);
xor U274 (N_274,In_1731,In_1352);
and U275 (N_275,In_238,In_2673);
or U276 (N_276,In_1910,In_1725);
nor U277 (N_277,In_461,In_1028);
or U278 (N_278,In_1333,In_2987);
and U279 (N_279,In_876,In_2556);
and U280 (N_280,In_1273,In_929);
xor U281 (N_281,In_2141,In_2348);
xnor U282 (N_282,In_1034,In_2621);
xnor U283 (N_283,In_2052,In_1048);
nor U284 (N_284,In_1319,In_2233);
xor U285 (N_285,In_1628,In_116);
xor U286 (N_286,In_2292,In_2306);
or U287 (N_287,In_899,In_17);
xnor U288 (N_288,In_913,In_1109);
xnor U289 (N_289,In_175,In_1511);
xor U290 (N_290,In_1805,In_1677);
and U291 (N_291,In_2737,In_1272);
nand U292 (N_292,In_1285,In_1332);
nor U293 (N_293,In_192,In_2297);
and U294 (N_294,In_2407,In_714);
or U295 (N_295,In_549,In_428);
or U296 (N_296,In_2059,In_2501);
or U297 (N_297,In_1722,In_1971);
nand U298 (N_298,In_71,In_2245);
nand U299 (N_299,In_2552,In_2756);
nor U300 (N_300,In_1478,In_1134);
or U301 (N_301,In_1355,In_624);
nor U302 (N_302,In_696,In_2811);
or U303 (N_303,In_2479,In_5);
and U304 (N_304,In_1066,In_579);
xor U305 (N_305,In_2890,In_2946);
nor U306 (N_306,In_1986,In_2007);
nand U307 (N_307,In_570,In_1732);
and U308 (N_308,In_142,In_1014);
or U309 (N_309,In_690,In_2642);
and U310 (N_310,In_662,In_666);
nor U311 (N_311,In_31,In_2847);
nor U312 (N_312,In_2011,In_442);
nand U313 (N_313,In_1967,In_2849);
xor U314 (N_314,In_2583,In_1829);
nor U315 (N_315,In_2026,In_1183);
nor U316 (N_316,In_550,In_1808);
nor U317 (N_317,In_2992,In_2830);
and U318 (N_318,In_2900,In_466);
nand U319 (N_319,In_2995,In_1624);
nand U320 (N_320,In_324,In_798);
and U321 (N_321,In_2561,In_200);
nand U322 (N_322,In_1721,In_1297);
nand U323 (N_323,In_2323,In_1078);
xnor U324 (N_324,In_2605,In_151);
xnor U325 (N_325,In_896,In_672);
nand U326 (N_326,In_1738,In_462);
nand U327 (N_327,In_1601,In_1839);
nor U328 (N_328,In_1940,In_1435);
nand U329 (N_329,In_2203,In_551);
xor U330 (N_330,In_755,In_263);
and U331 (N_331,In_604,In_1148);
or U332 (N_332,In_994,In_2360);
nor U333 (N_333,In_1659,In_2966);
xnor U334 (N_334,In_877,In_1914);
xor U335 (N_335,In_337,In_543);
nand U336 (N_336,In_173,In_2544);
or U337 (N_337,In_1254,In_2425);
and U338 (N_338,In_2340,In_1833);
xnor U339 (N_339,In_2057,In_1650);
and U340 (N_340,In_1843,In_497);
xor U341 (N_341,In_243,In_2692);
xor U342 (N_342,In_2146,In_2652);
xor U343 (N_343,In_1752,In_432);
xnor U344 (N_344,In_2827,In_1726);
and U345 (N_345,In_1323,In_825);
xor U346 (N_346,In_2856,In_2963);
nand U347 (N_347,In_629,In_1751);
or U348 (N_348,In_2288,In_2457);
or U349 (N_349,In_1264,In_387);
and U350 (N_350,In_987,In_685);
and U351 (N_351,In_1629,In_1684);
nand U352 (N_352,In_2729,In_1947);
xor U353 (N_353,In_7,In_1862);
xnor U354 (N_354,In_2582,In_1852);
nor U355 (N_355,In_76,In_100);
xor U356 (N_356,In_2326,In_150);
or U357 (N_357,In_2685,In_2525);
nor U358 (N_358,In_620,In_547);
and U359 (N_359,In_156,In_2948);
nand U360 (N_360,In_434,In_713);
nor U361 (N_361,In_894,In_1444);
nor U362 (N_362,In_226,In_1757);
nand U363 (N_363,In_1400,In_2498);
nand U364 (N_364,In_50,In_1583);
and U365 (N_365,In_635,In_841);
xnor U366 (N_366,In_347,In_1164);
nor U367 (N_367,In_1873,In_52);
or U368 (N_368,In_2243,In_77);
or U369 (N_369,In_858,In_94);
or U370 (N_370,In_1978,In_157);
or U371 (N_371,In_2897,In_198);
nor U372 (N_372,In_2114,In_2736);
nand U373 (N_373,In_1891,In_294);
nor U374 (N_374,In_2970,In_2307);
and U375 (N_375,In_2028,In_1158);
and U376 (N_376,In_1461,In_826);
or U377 (N_377,In_1672,In_1074);
xnor U378 (N_378,In_1090,In_367);
xor U379 (N_379,In_1451,In_1869);
or U380 (N_380,In_2389,In_719);
xor U381 (N_381,In_988,In_2332);
xnor U382 (N_382,In_1847,In_2529);
nor U383 (N_383,In_1063,In_2705);
and U384 (N_384,In_1247,In_1162);
xor U385 (N_385,In_2408,In_380);
nand U386 (N_386,In_326,In_1108);
nand U387 (N_387,In_2870,In_133);
or U388 (N_388,In_111,In_2531);
and U389 (N_389,In_155,In_2703);
nand U390 (N_390,In_984,In_1881);
xor U391 (N_391,In_1801,In_1346);
and U392 (N_392,In_1215,In_2452);
xnor U393 (N_393,In_2077,In_358);
nand U394 (N_394,In_1384,In_818);
and U395 (N_395,In_476,In_1858);
nand U396 (N_396,In_1313,In_2519);
and U397 (N_397,In_2167,In_2109);
and U398 (N_398,In_1595,In_505);
and U399 (N_399,In_799,In_1054);
xor U400 (N_400,In_2173,In_1452);
xnor U401 (N_401,In_2754,In_1036);
nand U402 (N_402,In_1171,In_2669);
nor U403 (N_403,In_1121,In_1534);
nor U404 (N_404,In_1737,In_2067);
xnor U405 (N_405,In_2119,In_403);
nor U406 (N_406,In_1474,In_2781);
and U407 (N_407,In_2135,In_419);
and U408 (N_408,In_910,In_2887);
xor U409 (N_409,In_2975,In_2295);
and U410 (N_410,In_1330,In_2440);
xor U411 (N_411,In_2810,In_967);
nand U412 (N_412,In_1683,In_612);
nand U413 (N_413,In_338,In_1154);
and U414 (N_414,In_429,In_33);
nor U415 (N_415,In_1651,In_1167);
xnor U416 (N_416,In_1191,In_496);
or U417 (N_417,In_2019,In_1150);
and U418 (N_418,In_1339,In_1961);
xnor U419 (N_419,In_2853,In_68);
nand U420 (N_420,In_2021,In_784);
and U421 (N_421,In_2671,In_1941);
xnor U422 (N_422,In_1399,In_844);
xnor U423 (N_423,In_1625,In_2752);
and U424 (N_424,In_1239,In_2577);
nand U425 (N_425,In_985,In_2160);
and U426 (N_426,In_2363,In_2791);
or U427 (N_427,In_764,In_980);
and U428 (N_428,In_1314,In_1957);
and U429 (N_429,In_1106,In_2753);
nand U430 (N_430,In_166,In_1364);
or U431 (N_431,In_1906,In_2779);
and U432 (N_432,In_2576,In_2391);
and U433 (N_433,In_1689,In_1021);
nand U434 (N_434,In_1386,In_717);
and U435 (N_435,In_1427,In_1469);
or U436 (N_436,In_889,In_1135);
and U437 (N_437,In_1789,In_239);
nor U438 (N_438,In_2570,In_1156);
and U439 (N_439,In_1987,In_2932);
or U440 (N_440,In_1608,In_2615);
and U441 (N_441,In_1798,In_1874);
xnor U442 (N_442,In_976,In_1115);
or U443 (N_443,In_1423,In_123);
nand U444 (N_444,In_1438,In_273);
or U445 (N_445,In_1544,In_2590);
nand U446 (N_446,In_2320,In_75);
xnor U447 (N_447,In_1371,In_179);
xor U448 (N_448,In_204,In_206);
nor U449 (N_449,In_1426,In_701);
nand U450 (N_450,In_867,In_141);
nand U451 (N_451,In_2982,In_1244);
and U452 (N_452,In_809,In_2508);
xnor U453 (N_453,In_2587,In_2663);
nand U454 (N_454,In_2716,In_2148);
xor U455 (N_455,In_885,In_441);
and U456 (N_456,In_187,In_2496);
or U457 (N_457,In_1753,In_787);
or U458 (N_458,In_767,In_1089);
or U459 (N_459,In_2409,In_350);
xnor U460 (N_460,In_2310,In_586);
xnor U461 (N_461,In_1084,In_1495);
or U462 (N_462,In_786,In_21);
and U463 (N_463,In_97,In_830);
or U464 (N_464,In_254,In_1931);
and U465 (N_465,In_626,In_2008);
and U466 (N_466,In_1739,In_1071);
or U467 (N_467,In_1174,In_1585);
nor U468 (N_468,In_848,In_63);
nand U469 (N_469,In_1765,In_43);
nor U470 (N_470,In_412,In_1715);
nor U471 (N_471,In_274,In_2979);
xnor U472 (N_472,In_2818,In_969);
nor U473 (N_473,In_2936,In_791);
and U474 (N_474,In_1504,In_1139);
and U475 (N_475,In_1768,In_2722);
and U476 (N_476,In_821,In_2053);
xor U477 (N_477,In_1069,In_1574);
and U478 (N_478,In_1509,In_2474);
or U479 (N_479,In_1485,In_2293);
nor U480 (N_480,In_1767,In_244);
or U481 (N_481,In_597,In_2105);
or U482 (N_482,In_1284,In_1742);
or U483 (N_483,In_2287,In_2971);
and U484 (N_484,In_2025,In_2219);
or U485 (N_485,In_152,In_569);
nand U486 (N_486,In_1619,In_1468);
nand U487 (N_487,In_2231,In_2211);
nor U488 (N_488,In_1921,In_2762);
and U489 (N_489,In_296,In_611);
nand U490 (N_490,In_2915,In_1717);
nor U491 (N_491,In_402,In_2242);
xor U492 (N_492,In_178,In_526);
nand U493 (N_493,In_1449,In_2198);
nor U494 (N_494,In_1696,In_250);
nand U495 (N_495,In_2324,In_2189);
nand U496 (N_496,In_373,In_682);
or U497 (N_497,In_1617,In_815);
nor U498 (N_498,In_507,In_2603);
nor U499 (N_499,In_1456,In_2907);
and U500 (N_500,In_3,In_2404);
nand U501 (N_501,In_2229,In_2666);
xor U502 (N_502,In_1370,In_1834);
nor U503 (N_503,In_1813,In_907);
and U504 (N_504,In_430,In_2517);
and U505 (N_505,In_95,In_1039);
nor U506 (N_506,In_1213,In_2883);
and U507 (N_507,In_259,In_27);
and U508 (N_508,In_2083,In_1919);
or U509 (N_509,In_2195,In_399);
nor U510 (N_510,In_1492,In_1668);
nor U511 (N_511,In_1404,In_1410);
xnor U512 (N_512,In_2990,In_1023);
or U513 (N_513,In_194,In_596);
nor U514 (N_514,In_1116,In_386);
xor U515 (N_515,In_427,In_1523);
or U516 (N_516,In_1576,In_609);
nor U517 (N_517,In_1626,In_2103);
or U518 (N_518,In_760,In_153);
or U519 (N_519,In_531,In_411);
or U520 (N_520,In_642,In_1336);
or U521 (N_521,In_2744,In_1);
and U522 (N_522,In_2035,In_284);
nor U523 (N_523,In_986,In_1850);
and U524 (N_524,In_2563,In_325);
nand U525 (N_525,In_2527,In_2719);
nor U526 (N_526,In_2725,In_572);
or U527 (N_527,In_2998,In_1779);
and U528 (N_528,In_1372,In_2186);
nand U529 (N_529,In_888,In_484);
and U530 (N_530,In_1019,In_1741);
nand U531 (N_531,In_2336,In_2539);
or U532 (N_532,In_1251,In_1443);
nand U533 (N_533,In_637,In_2630);
or U534 (N_534,In_938,In_1009);
xnor U535 (N_535,In_2061,In_1989);
or U536 (N_536,In_2094,In_2759);
nand U537 (N_537,In_2977,In_1142);
xor U538 (N_538,In_1918,In_1996);
xnor U539 (N_539,In_1604,In_1223);
xor U540 (N_540,In_2553,In_1086);
or U541 (N_541,In_455,In_566);
or U542 (N_542,In_1559,In_1000);
nand U543 (N_543,In_426,In_2532);
xnor U544 (N_544,In_138,In_1367);
or U545 (N_545,In_2247,In_1793);
and U546 (N_546,In_2437,In_1762);
xor U547 (N_547,In_1596,In_193);
or U548 (N_548,In_2345,In_1383);
nand U549 (N_549,In_2925,In_2728);
and U550 (N_550,In_2633,In_512);
and U551 (N_551,In_234,In_137);
or U552 (N_552,In_481,In_618);
or U553 (N_553,In_1051,In_1255);
and U554 (N_554,In_1005,In_952);
and U555 (N_555,In_1407,In_790);
and U556 (N_556,In_2509,In_112);
and U557 (N_557,In_964,In_15);
nor U558 (N_558,In_59,In_2822);
nand U559 (N_559,In_1481,In_1641);
nand U560 (N_560,In_1360,In_1736);
nor U561 (N_561,In_1676,In_1913);
nand U562 (N_562,In_83,In_2373);
or U563 (N_563,In_1632,In_56);
nand U564 (N_564,In_1418,In_2417);
nor U565 (N_565,In_26,In_694);
xnor U566 (N_566,In_908,In_1127);
nor U567 (N_567,In_1231,In_2163);
xor U568 (N_568,In_2514,In_2910);
xor U569 (N_569,In_417,In_2276);
nor U570 (N_570,In_397,In_2940);
xor U571 (N_571,In_2255,In_2934);
xor U572 (N_572,In_1988,In_1335);
xor U573 (N_573,In_62,In_246);
or U574 (N_574,In_163,In_220);
xor U575 (N_575,In_2751,In_2585);
or U576 (N_576,In_1800,In_280);
or U577 (N_577,In_1526,In_946);
nor U578 (N_578,In_2371,In_2524);
and U579 (N_579,In_2999,In_2050);
xnor U580 (N_580,In_2112,In_2442);
nand U581 (N_581,In_2891,In_749);
or U582 (N_582,In_1563,In_1118);
nor U583 (N_583,In_1899,In_2659);
or U584 (N_584,In_2232,In_2834);
nand U585 (N_585,In_2775,In_34);
nand U586 (N_586,In_2879,In_2241);
xor U587 (N_587,In_1368,In_792);
xor U588 (N_588,In_2928,In_1324);
nor U589 (N_589,In_854,In_1221);
and U590 (N_590,In_1857,In_1018);
and U591 (N_591,In_406,In_423);
or U592 (N_592,In_127,In_744);
nand U593 (N_593,In_136,In_1100);
and U594 (N_594,In_1973,In_57);
or U595 (N_595,In_1985,In_780);
and U596 (N_596,In_2789,In_2439);
and U597 (N_597,In_2504,In_2096);
nor U598 (N_598,In_1754,In_511);
or U599 (N_599,In_1945,In_2330);
or U600 (N_600,In_676,In_29);
nand U601 (N_601,In_2884,In_1701);
nand U602 (N_602,In_1939,In_2578);
or U603 (N_603,In_2191,In_585);
nand U604 (N_604,In_1248,In_1727);
nor U605 (N_605,In_2101,In_1463);
and U606 (N_606,In_2937,In_1827);
or U607 (N_607,In_1375,In_2520);
nand U608 (N_608,In_2997,In_613);
or U609 (N_609,In_1508,In_1860);
xnor U610 (N_610,In_1775,In_667);
xnor U611 (N_611,In_1082,In_2644);
xor U612 (N_612,In_1055,In_2397);
and U613 (N_613,In_130,In_414);
and U614 (N_614,In_645,In_1781);
and U615 (N_615,In_1507,In_2218);
and U616 (N_616,In_66,In_1366);
and U617 (N_617,In_327,In_464);
nor U618 (N_618,In_360,In_492);
xor U619 (N_619,In_565,In_309);
nand U620 (N_620,In_2412,In_965);
nor U621 (N_621,In_730,In_1252);
and U622 (N_622,In_1408,In_834);
and U623 (N_623,In_1238,In_1674);
nor U624 (N_624,In_1679,In_1791);
nand U625 (N_625,In_2926,In_912);
nor U626 (N_626,In_868,In_1772);
nor U627 (N_627,In_313,In_1342);
and U628 (N_628,In_242,In_12);
xnor U629 (N_629,In_1122,In_2207);
nand U630 (N_630,In_687,In_494);
nand U631 (N_631,In_2194,In_1312);
nand U632 (N_632,In_2309,In_1812);
or U633 (N_633,In_807,In_2745);
and U634 (N_634,In_498,In_1975);
nand U635 (N_635,In_1376,In_2127);
xor U636 (N_636,In_2248,In_1043);
nand U637 (N_637,In_1040,In_2088);
or U638 (N_638,In_2908,In_1286);
or U639 (N_639,In_2909,In_2068);
nor U640 (N_640,In_2366,In_2418);
nor U641 (N_641,In_2903,In_2387);
nor U642 (N_642,In_953,In_2770);
nand U643 (N_643,In_2410,In_1334);
nand U644 (N_644,In_2876,In_2575);
nor U645 (N_645,In_1655,In_1287);
nor U646 (N_646,In_289,In_1081);
xor U647 (N_647,In_91,In_2104);
xor U648 (N_648,In_283,In_2986);
nand U649 (N_649,In_1581,In_1718);
or U650 (N_650,In_1240,In_1901);
nand U651 (N_651,In_2765,In_1070);
nor U652 (N_652,In_408,In_126);
and U653 (N_653,In_2267,In_633);
xor U654 (N_654,In_1530,In_707);
and U655 (N_655,In_546,In_2361);
xor U656 (N_656,In_2706,In_281);
nor U657 (N_657,In_1694,In_659);
or U658 (N_658,In_520,In_1803);
and U659 (N_659,In_1570,In_595);
nand U660 (N_660,In_568,In_1934);
nor U661 (N_661,In_2177,In_2942);
nor U662 (N_662,In_334,In_1733);
nand U663 (N_663,In_362,In_2904);
nor U664 (N_664,In_42,In_831);
nand U665 (N_665,In_2931,In_1926);
and U666 (N_666,In_314,In_1582);
xor U667 (N_667,In_2443,In_592);
xor U668 (N_668,In_1666,In_1916);
and U669 (N_669,In_1388,In_188);
nor U670 (N_670,In_712,In_2451);
nand U671 (N_671,In_202,In_1260);
xnor U672 (N_672,In_1631,In_817);
nand U673 (N_673,In_1851,In_2395);
nor U674 (N_674,In_2185,In_1903);
or U675 (N_675,In_1755,In_140);
xor U676 (N_676,In_2793,In_535);
xnor U677 (N_677,In_2382,In_0);
nand U678 (N_678,In_2647,In_709);
nor U679 (N_679,In_1349,In_919);
nand U680 (N_680,In_1807,In_1774);
nor U681 (N_681,In_674,In_78);
or U682 (N_682,In_1401,In_2147);
and U683 (N_683,In_1894,In_1607);
and U684 (N_684,In_2620,In_522);
nand U685 (N_685,In_2256,In_2914);
or U686 (N_686,In_1350,In_2560);
xor U687 (N_687,In_1288,In_1361);
nand U688 (N_688,In_2465,In_558);
nor U689 (N_689,In_1378,In_2192);
nand U690 (N_690,In_1278,In_1271);
nor U691 (N_691,In_2038,In_1569);
or U692 (N_692,In_213,In_1578);
nor U693 (N_693,In_2151,In_2093);
or U694 (N_694,In_225,In_2597);
nand U695 (N_695,In_479,In_2954);
nor U696 (N_696,In_1942,In_1880);
xor U697 (N_697,In_2586,In_796);
xnor U698 (N_698,In_542,In_459);
and U699 (N_699,In_2782,In_515);
and U700 (N_700,In_46,In_1623);
nor U701 (N_701,In_948,In_1611);
or U702 (N_702,In_788,In_1420);
and U703 (N_703,In_1706,In_2237);
and U704 (N_704,In_1528,In_1079);
or U705 (N_705,In_2268,In_2001);
xor U706 (N_706,In_10,In_2056);
or U707 (N_707,In_1925,In_2250);
nand U708 (N_708,In_2042,In_1888);
nand U709 (N_709,In_1904,In_1802);
nand U710 (N_710,In_1982,In_1417);
and U711 (N_711,In_1207,In_1363);
nor U712 (N_712,In_705,In_2851);
or U713 (N_713,In_665,In_2343);
xnor U714 (N_714,In_927,In_1981);
or U715 (N_715,In_376,In_2606);
nor U716 (N_716,In_2739,In_865);
nor U717 (N_717,In_1295,In_1318);
and U718 (N_718,In_2178,In_460);
nand U719 (N_719,In_2800,In_1561);
and U720 (N_720,In_2780,In_2807);
nand U721 (N_721,In_2973,In_700);
and U722 (N_722,In_1347,In_1406);
xnor U723 (N_723,In_2741,In_1094);
and U724 (N_724,In_954,In_361);
and U725 (N_725,In_1035,In_1944);
or U726 (N_726,In_483,In_2273);
or U727 (N_727,In_1799,In_379);
xnor U728 (N_728,In_2436,In_1380);
xnor U729 (N_729,In_2801,In_1782);
nand U730 (N_730,In_1917,In_2639);
and U731 (N_731,In_776,In_2555);
and U732 (N_732,In_2902,In_752);
and U733 (N_733,In_1594,In_634);
nand U734 (N_734,In_557,In_435);
nand U735 (N_735,In_843,In_2214);
and U736 (N_736,In_2125,In_2626);
nor U737 (N_737,In_870,In_191);
or U738 (N_738,In_1362,In_1796);
xnor U739 (N_739,In_574,In_2616);
xnor U740 (N_740,In_1083,In_1951);
nor U741 (N_741,In_390,In_2123);
xnor U742 (N_742,In_2548,In_732);
nor U743 (N_743,In_2161,In_103);
nor U744 (N_744,In_2070,In_652);
or U745 (N_745,In_2549,In_1907);
xnor U746 (N_746,In_2758,In_2564);
nand U747 (N_747,In_1020,In_1660);
nor U748 (N_748,In_529,In_405);
nand U749 (N_749,In_2393,In_718);
and U750 (N_750,In_2611,In_972);
or U751 (N_751,In_450,In_2837);
xnor U752 (N_752,In_2422,In_1948);
xnor U753 (N_753,In_2565,In_475);
nor U754 (N_754,In_2804,In_2102);
and U755 (N_755,In_1794,In_121);
and U756 (N_756,In_2347,In_2188);
xor U757 (N_757,In_1243,In_2893);
or U758 (N_758,In_60,In_1923);
or U759 (N_759,In_1551,In_37);
or U760 (N_760,In_2541,In_1537);
and U761 (N_761,In_2139,In_2943);
and U762 (N_762,In_1645,In_1830);
nand U763 (N_763,In_2117,In_2217);
nand U764 (N_764,In_905,In_36);
nor U765 (N_765,In_1316,In_2878);
nor U766 (N_766,In_2006,In_836);
nor U767 (N_767,In_1740,In_2924);
and U768 (N_768,In_503,In_1276);
nor U769 (N_769,In_1389,In_1627);
nand U770 (N_770,In_2672,In_1905);
nor U771 (N_771,In_1871,In_1823);
or U772 (N_772,In_1516,In_2370);
nor U773 (N_773,In_1015,In_1777);
nor U774 (N_774,In_2062,In_1395);
xnor U775 (N_775,In_2374,In_6);
and U776 (N_776,In_1253,In_1909);
xnor U777 (N_777,In_1031,In_265);
xor U778 (N_778,In_2812,In_2180);
or U779 (N_779,In_1227,In_1692);
nor U780 (N_780,In_1897,In_2985);
xnor U781 (N_781,In_2341,In_1867);
nand U782 (N_782,In_955,In_2212);
nor U783 (N_783,In_2489,In_974);
nor U784 (N_784,In_981,In_2815);
nand U785 (N_785,In_552,In_2911);
nand U786 (N_786,In_222,In_172);
nor U787 (N_787,In_195,In_1671);
and U788 (N_788,In_2976,In_863);
and U789 (N_789,In_344,In_916);
or U790 (N_790,In_1972,In_1200);
nor U791 (N_791,In_2369,In_2784);
xor U792 (N_792,In_866,In_23);
and U793 (N_793,In_903,In_451);
nand U794 (N_794,In_85,In_1695);
and U795 (N_795,In_537,In_189);
nand U796 (N_796,In_339,In_1959);
nand U797 (N_797,In_926,In_2675);
xor U798 (N_798,In_2082,In_2272);
nor U799 (N_799,In_1702,In_1433);
and U800 (N_800,In_258,In_1974);
nor U801 (N_801,In_352,In_887);
nand U802 (N_802,In_1457,In_1937);
nor U803 (N_803,In_820,In_2748);
xor U804 (N_804,In_1064,In_892);
nor U805 (N_805,In_802,In_2657);
or U806 (N_806,In_1704,In_1713);
xnor U807 (N_807,In_2221,In_2650);
nand U808 (N_808,In_2690,In_2448);
or U809 (N_809,In_8,In_989);
xnor U810 (N_810,In_310,In_488);
or U811 (N_811,In_1745,In_660);
xnor U812 (N_812,In_171,In_2190);
nor U813 (N_813,In_264,In_2499);
and U814 (N_814,In_2076,In_2264);
nand U815 (N_815,In_581,In_2483);
xor U816 (N_816,In_1709,In_2278);
and U817 (N_817,In_2168,In_1137);
nand U818 (N_818,In_587,In_561);
nor U819 (N_819,In_2707,In_785);
xnor U820 (N_820,In_9,In_2086);
nor U821 (N_821,In_247,In_765);
and U822 (N_822,In_1535,In_734);
nand U823 (N_823,In_2569,In_2234);
or U824 (N_824,In_375,In_833);
xnor U825 (N_825,In_921,In_1552);
nor U826 (N_826,In_275,In_639);
or U827 (N_827,In_1700,In_2459);
or U828 (N_828,In_1838,In_1146);
xnor U829 (N_829,In_1345,In_1102);
or U830 (N_830,In_131,In_2154);
and U831 (N_831,In_2538,In_1151);
and U832 (N_832,In_2200,In_92);
xnor U833 (N_833,In_1268,In_1760);
xnor U834 (N_834,In_2814,In_2704);
and U835 (N_835,In_623,In_2886);
or U836 (N_836,In_1597,In_884);
nand U837 (N_837,In_58,In_641);
nor U838 (N_838,In_1356,In_1246);
or U839 (N_839,In_2857,In_2648);
nor U840 (N_840,In_2486,In_1825);
nand U841 (N_841,In_1204,In_1450);
or U842 (N_842,In_96,In_1241);
xnor U843 (N_843,In_2149,In_1098);
and U844 (N_844,In_1216,In_1790);
xor U845 (N_845,In_1614,In_2727);
nand U846 (N_846,In_1505,In_536);
nand U847 (N_847,In_506,In_1610);
or U848 (N_848,In_2771,In_2894);
nand U849 (N_849,In_1290,In_643);
nor U850 (N_850,In_2557,In_1557);
nand U851 (N_851,In_2420,In_1846);
or U852 (N_852,In_2484,In_1667);
and U853 (N_853,In_2738,In_1262);
xnor U854 (N_854,In_221,In_1946);
nor U855 (N_855,In_804,In_2472);
nand U856 (N_856,In_1887,In_2638);
nor U857 (N_857,In_838,In_215);
xnor U858 (N_858,In_956,In_2848);
or U859 (N_859,In_2433,In_689);
nand U860 (N_860,In_1962,In_2918);
and U861 (N_861,In_1205,In_1605);
xor U862 (N_862,In_1257,In_2787);
nor U863 (N_863,In_909,In_2279);
nand U864 (N_864,In_331,In_2874);
nor U865 (N_865,In_343,In_603);
and U866 (N_866,In_855,In_1396);
nor U867 (N_867,In_727,In_1459);
and U868 (N_868,In_1267,In_1588);
nor U869 (N_869,In_1855,In_1471);
or U870 (N_870,In_1652,In_1331);
or U871 (N_871,In_2137,In_2175);
nand U872 (N_872,In_2421,In_216);
nand U873 (N_873,In_2805,In_2429);
nor U874 (N_874,In_1820,In_2612);
xor U875 (N_875,In_278,In_145);
xnor U876 (N_876,In_181,In_2664);
xor U877 (N_877,In_813,In_650);
nor U878 (N_878,In_415,In_413);
xor U879 (N_879,In_2764,In_2841);
and U880 (N_880,In_2864,In_2960);
xnor U881 (N_881,In_950,In_638);
or U882 (N_882,In_1311,In_1045);
and U883 (N_883,In_1016,In_2731);
or U884 (N_884,In_691,In_1042);
nor U885 (N_885,In_1885,In_1893);
xnor U886 (N_886,In_2165,In_627);
nor U887 (N_887,In_2396,In_2464);
or U888 (N_888,In_2760,In_859);
or U889 (N_889,In_2584,In_1872);
nor U890 (N_890,In_229,In_203);
nor U891 (N_891,In_2788,In_164);
nor U892 (N_892,In_2604,In_2100);
and U893 (N_893,In_61,In_2379);
nor U894 (N_894,In_392,In_18);
or U895 (N_895,In_739,In_262);
and U896 (N_896,In_2660,In_2686);
xor U897 (N_897,In_1744,In_904);
and U898 (N_898,In_2301,In_647);
xnor U899 (N_899,In_370,In_1030);
xnor U900 (N_900,In_2110,In_1930);
nand U901 (N_901,In_132,In_2072);
nor U902 (N_902,In_2353,In_533);
nor U903 (N_903,In_482,In_1385);
nand U904 (N_904,In_2359,In_2005);
xor U905 (N_905,In_1868,In_741);
xor U906 (N_906,In_2817,In_1963);
nand U907 (N_907,In_454,In_553);
nand U908 (N_908,In_2795,In_1193);
nand U909 (N_909,In_1105,In_2512);
nor U910 (N_910,In_257,In_2831);
or U911 (N_911,In_1653,In_1250);
or U912 (N_912,In_2210,In_122);
nand U913 (N_913,In_2930,In_1062);
xnor U914 (N_914,In_2740,In_935);
or U915 (N_915,In_2403,In_2613);
or U916 (N_916,In_1409,In_346);
nor U917 (N_917,In_2438,In_673);
nor U918 (N_918,In_340,In_1421);
xnor U919 (N_919,In_69,In_1491);
xor U920 (N_920,In_697,In_657);
nor U921 (N_921,In_2617,In_1113);
nand U922 (N_922,In_348,In_720);
xor U923 (N_923,In_359,In_1877);
xor U924 (N_924,In_404,In_117);
and U925 (N_925,In_2225,In_282);
and U926 (N_926,In_1466,In_2174);
nor U927 (N_927,In_1994,In_2854);
nor U928 (N_928,In_2607,In_1099);
nor U929 (N_929,In_1831,In_438);
nor U930 (N_930,In_1993,In_1026);
or U931 (N_931,In_154,In_1821);
and U932 (N_932,In_770,In_1841);
or U933 (N_933,In_2825,In_775);
nand U934 (N_934,In_1506,In_297);
xnor U935 (N_935,In_1197,In_342);
nand U936 (N_936,In_2715,In_1412);
xor U937 (N_937,In_1723,In_2208);
and U938 (N_938,In_2545,In_2071);
or U939 (N_939,In_2228,In_2502);
nor U940 (N_940,In_2938,In_2843);
nor U941 (N_941,In_2138,In_2491);
xnor U942 (N_942,In_2018,In_2896);
xnor U943 (N_943,In_678,In_291);
nand U944 (N_944,In_1599,In_2344);
and U945 (N_945,In_932,In_184);
nor U946 (N_946,In_1017,In_1832);
xnor U947 (N_947,In_1602,In_382);
nor U948 (N_948,In_2205,In_2962);
and U949 (N_949,In_2898,In_487);
nor U950 (N_950,In_2772,In_207);
nor U951 (N_951,In_1567,In_2342);
and U952 (N_952,In_1573,In_575);
xnor U953 (N_953,In_2400,In_1932);
or U954 (N_954,In_582,In_1322);
and U955 (N_955,In_1633,In_2839);
or U956 (N_956,In_2377,In_478);
nand U957 (N_957,In_2511,In_2476);
xor U958 (N_958,In_2862,In_2058);
and U959 (N_959,In_1618,In_328);
nor U960 (N_960,In_1184,In_1170);
nor U961 (N_961,In_2386,In_409);
or U962 (N_962,In_1587,In_1734);
or U963 (N_963,In_307,In_1317);
nand U964 (N_964,In_2447,In_2478);
and U965 (N_965,In_2375,In_1189);
xor U966 (N_966,In_1049,In_119);
nand U967 (N_967,In_2865,In_992);
or U968 (N_968,In_2773,In_1326);
nand U969 (N_969,In_2406,In_2357);
nor U970 (N_970,In_2885,In_900);
nor U971 (N_971,In_1687,In_1029);
xor U972 (N_972,In_616,In_716);
or U973 (N_973,In_1419,In_113);
nand U974 (N_974,In_2124,In_2010);
nand U975 (N_975,In_1470,In_651);
nor U976 (N_976,In_636,In_128);
xnor U977 (N_977,In_1374,In_1525);
xnor U978 (N_978,In_1889,In_107);
nand U979 (N_979,In_208,In_2974);
and U980 (N_980,In_625,In_349);
nand U981 (N_981,In_1025,In_2286);
or U982 (N_982,In_436,In_335);
and U983 (N_983,In_174,In_1920);
and U984 (N_984,In_2048,In_1984);
or U985 (N_985,In_356,In_2384);
or U986 (N_986,In_1710,In_2631);
xor U987 (N_987,In_2334,In_990);
or U988 (N_988,In_663,In_1836);
xnor U989 (N_989,In_644,In_2480);
or U990 (N_990,In_2368,In_1093);
or U991 (N_991,In_937,In_628);
or U992 (N_992,In_471,In_110);
nor U993 (N_993,In_2798,In_489);
nor U994 (N_994,In_1249,In_440);
xnor U995 (N_995,In_2424,In_224);
and U996 (N_996,In_1639,In_2767);
nor U997 (N_997,In_1927,In_564);
and U998 (N_998,In_308,In_851);
and U999 (N_999,In_1002,In_2594);
and U1000 (N_1000,In_443,In_2861);
nor U1001 (N_1001,N_432,In_2128);
xor U1002 (N_1002,N_659,N_708);
and U1003 (N_1003,N_581,In_2291);
xor U1004 (N_1004,N_412,N_725);
nor U1005 (N_1005,N_548,In_2855);
nand U1006 (N_1006,N_223,N_462);
xor U1007 (N_1007,In_1024,In_2390);
or U1008 (N_1008,In_2296,N_726);
or U1009 (N_1009,In_2230,In_182);
and U1010 (N_1010,N_145,In_2628);
and U1011 (N_1011,N_510,In_2844);
or U1012 (N_1012,In_1211,N_718);
and U1013 (N_1013,N_497,In_1613);
nor U1014 (N_1014,In_936,N_621);
nand U1015 (N_1015,N_564,N_655);
or U1016 (N_1016,In_1065,N_943);
nand U1017 (N_1017,N_243,N_39);
and U1018 (N_1018,In_1176,N_63);
nor U1019 (N_1019,N_59,N_942);
nand U1020 (N_1020,In_2547,N_416);
nand U1021 (N_1021,N_123,In_1397);
or U1022 (N_1022,N_194,In_1609);
xnor U1023 (N_1023,N_338,N_880);
and U1024 (N_1024,N_47,N_62);
and U1025 (N_1025,In_1218,N_222);
xnor U1026 (N_1026,In_1088,N_939);
xor U1027 (N_1027,In_772,N_347);
and U1028 (N_1028,N_912,In_538);
and U1029 (N_1029,In_1077,In_2327);
and U1030 (N_1030,N_72,N_436);
xor U1031 (N_1031,N_69,In_1104);
or U1032 (N_1032,N_649,In_2319);
and U1033 (N_1033,N_401,In_1458);
nor U1034 (N_1034,In_1882,In_745);
nand U1035 (N_1035,In_2959,N_56);
nand U1036 (N_1036,In_2432,In_2316);
and U1037 (N_1037,N_310,N_825);
xnor U1038 (N_1038,In_371,N_166);
and U1039 (N_1039,In_850,N_614);
nand U1040 (N_1040,In_2157,N_395);
nand U1041 (N_1041,N_728,In_1864);
nor U1042 (N_1042,N_13,In_1703);
xor U1043 (N_1043,In_726,N_299);
nand U1044 (N_1044,N_16,In_1172);
and U1045 (N_1045,N_787,N_64);
or U1046 (N_1046,In_2991,In_218);
xnor U1047 (N_1047,N_910,In_1966);
or U1048 (N_1048,N_842,In_1003);
nand U1049 (N_1049,N_190,N_859);
and U1050 (N_1050,N_304,N_428);
or U1051 (N_1051,N_712,In_1956);
nor U1052 (N_1052,In_2568,In_2676);
nor U1053 (N_1053,N_135,In_2776);
nor U1054 (N_1054,In_928,N_29);
or U1055 (N_1055,N_719,In_146);
xor U1056 (N_1056,In_1776,N_843);
nand U1057 (N_1057,N_660,N_99);
nor U1058 (N_1058,In_1068,In_924);
and U1059 (N_1059,In_2054,In_1658);
and U1060 (N_1060,In_48,N_425);
xor U1061 (N_1061,In_2792,N_421);
or U1062 (N_1062,N_466,N_79);
or U1063 (N_1063,N_346,In_420);
or U1064 (N_1064,N_814,In_2265);
xnor U1065 (N_1065,In_1424,N_477);
xor U1066 (N_1066,In_1540,N_903);
nand U1067 (N_1067,In_2600,N_526);
or U1068 (N_1068,N_812,In_1870);
nor U1069 (N_1069,N_215,In_2063);
or U1070 (N_1070,In_38,N_856);
nor U1071 (N_1071,In_1908,In_1126);
xnor U1072 (N_1072,In_1220,N_525);
and U1073 (N_1073,N_774,N_717);
or U1074 (N_1074,In_2311,In_1087);
nor U1075 (N_1075,In_1007,N_165);
and U1076 (N_1076,N_748,N_117);
or U1077 (N_1077,In_1636,In_2957);
xor U1078 (N_1078,In_2446,In_2111);
xor U1079 (N_1079,In_2274,In_1590);
xnor U1080 (N_1080,N_980,In_1579);
nor U1081 (N_1081,In_86,In_2958);
or U1082 (N_1082,In_1657,In_1152);
or U1083 (N_1083,In_2732,In_1866);
xor U1084 (N_1084,N_973,N_776);
nor U1085 (N_1085,In_610,N_322);
nor U1086 (N_1086,In_2004,In_2494);
and U1087 (N_1087,N_81,In_2654);
nand U1088 (N_1088,In_2947,N_7);
or U1089 (N_1089,N_957,In_1531);
xnor U1090 (N_1090,In_2254,In_384);
nor U1091 (N_1091,N_505,In_2271);
nor U1092 (N_1092,N_790,In_1178);
and U1093 (N_1093,N_558,In_2313);
xor U1094 (N_1094,N_898,N_492);
xnor U1095 (N_1095,N_121,N_890);
xor U1096 (N_1096,N_955,In_252);
nand U1097 (N_1097,In_365,In_129);
and U1098 (N_1098,In_1050,In_1282);
or U1099 (N_1099,N_661,In_2641);
nor U1100 (N_1100,In_2505,In_1720);
xor U1101 (N_1101,N_31,In_253);
nor U1102 (N_1102,N_783,In_87);
or U1103 (N_1103,In_1936,N_131);
and U1104 (N_1104,In_1952,N_629);
xnor U1105 (N_1105,N_592,In_933);
and U1106 (N_1106,N_560,N_146);
nand U1107 (N_1107,In_2643,In_2015);
nand U1108 (N_1108,In_89,N_94);
xnor U1109 (N_1109,In_2922,In_1256);
nor U1110 (N_1110,In_1785,N_265);
nor U1111 (N_1111,N_666,N_167);
or U1112 (N_1112,N_216,In_1856);
nor U1113 (N_1113,N_95,In_2624);
nor U1114 (N_1114,In_2315,N_444);
and U1115 (N_1115,N_788,In_539);
and U1116 (N_1116,In_1787,N_154);
and U1117 (N_1117,In_835,In_2667);
or U1118 (N_1118,N_187,N_839);
nand U1119 (N_1119,In_2598,In_2236);
or U1120 (N_1120,N_506,N_533);
and U1121 (N_1121,N_619,N_188);
nor U1122 (N_1122,In_864,N_625);
and U1123 (N_1123,In_2455,In_2352);
xnor U1124 (N_1124,In_2113,In_991);
or U1125 (N_1125,N_120,In_2304);
nand U1126 (N_1126,In_849,In_1661);
xnor U1127 (N_1127,In_1591,In_2799);
and U1128 (N_1128,In_2416,N_975);
and U1129 (N_1129,In_2972,In_1953);
nor U1130 (N_1130,In_2227,In_400);
or U1131 (N_1131,N_345,In_1411);
or U1132 (N_1132,N_23,In_998);
and U1133 (N_1133,N_398,N_937);
nand U1134 (N_1134,N_115,N_613);
and U1135 (N_1135,In_2073,In_1274);
or U1136 (N_1136,N_575,N_703);
and U1137 (N_1137,In_2710,N_297);
or U1138 (N_1138,N_272,In_1381);
and U1139 (N_1139,N_899,In_1080);
or U1140 (N_1140,In_336,N_175);
and U1141 (N_1141,N_257,N_796);
nor U1142 (N_1142,In_1714,N_132);
xor U1143 (N_1143,N_904,In_2108);
nand U1144 (N_1144,In_185,In_2097);
or U1145 (N_1145,In_1853,In_1296);
or U1146 (N_1146,N_35,In_2522);
nor U1147 (N_1147,In_368,In_545);
xnor U1148 (N_1148,In_918,N_802);
xor U1149 (N_1149,N_677,N_152);
xnor U1150 (N_1150,In_271,N_931);
nor U1151 (N_1151,N_214,N_978);
and U1152 (N_1152,N_765,In_1206);
nor U1153 (N_1153,N_692,N_645);
nor U1154 (N_1154,N_481,In_654);
xnor U1155 (N_1155,In_2562,In_467);
xor U1156 (N_1156,In_2106,N_104);
xnor U1157 (N_1157,N_539,In_766);
xor U1158 (N_1158,In_2964,In_1950);
nand U1159 (N_1159,In_118,In_1515);
xnor U1160 (N_1160,N_826,N_467);
or U1161 (N_1161,N_908,In_2338);
or U1162 (N_1162,In_1773,In_580);
nand U1163 (N_1163,In_1092,In_210);
nand U1164 (N_1164,N_200,In_2266);
nand U1165 (N_1165,N_231,In_2500);
or U1166 (N_1166,In_1465,In_1369);
nor U1167 (N_1167,In_1554,N_394);
nor U1168 (N_1168,In_753,In_1432);
nand U1169 (N_1169,N_339,In_410);
or U1170 (N_1170,N_693,N_543);
xor U1171 (N_1171,N_189,N_312);
and U1172 (N_1172,N_487,In_2030);
xnor U1173 (N_1173,In_1301,N_112);
or U1174 (N_1174,N_571,In_668);
nor U1175 (N_1175,N_114,N_761);
nor U1176 (N_1176,In_2949,In_1234);
and U1177 (N_1177,N_236,In_1145);
xor U1178 (N_1178,In_2260,N_885);
nor U1179 (N_1179,In_819,In_1589);
nand U1180 (N_1180,N_682,N_144);
or U1181 (N_1181,In_939,N_450);
and U1182 (N_1182,N_287,In_469);
and U1183 (N_1183,N_294,N_4);
and U1184 (N_1184,In_2702,N_595);
and U1185 (N_1185,N_845,In_812);
nor U1186 (N_1186,N_9,N_419);
and U1187 (N_1187,In_2087,N_934);
nand U1188 (N_1188,In_2551,In_2723);
xnor U1189 (N_1189,In_2913,N_782);
and U1190 (N_1190,In_2623,In_1536);
or U1191 (N_1191,In_1281,N_233);
and U1192 (N_1192,N_76,N_639);
nand U1193 (N_1193,N_203,N_58);
or U1194 (N_1194,In_571,N_951);
or U1195 (N_1195,In_2130,In_2697);
and U1196 (N_1196,In_2726,N_511);
nand U1197 (N_1197,N_411,In_1320);
or U1198 (N_1198,N_606,In_2832);
xnor U1199 (N_1199,N_838,In_2356);
and U1200 (N_1200,In_723,N_795);
nor U1201 (N_1201,In_1128,In_1705);
and U1202 (N_1202,N_344,N_565);
or U1203 (N_1203,N_71,N_417);
nand U1204 (N_1204,In_601,In_1995);
nand U1205 (N_1205,N_298,N_562);
and U1206 (N_1206,N_330,N_54);
and U1207 (N_1207,In_177,N_391);
and U1208 (N_1208,In_205,N_605);
or U1209 (N_1209,N_535,In_2475);
and U1210 (N_1210,In_199,In_2107);
nor U1211 (N_1211,In_711,N_291);
nor U1212 (N_1212,In_975,N_50);
or U1213 (N_1213,In_167,In_232);
and U1214 (N_1214,In_934,N_656);
or U1215 (N_1215,N_275,In_228);
and U1216 (N_1216,N_174,N_988);
nor U1217 (N_1217,N_65,N_648);
or U1218 (N_1218,In_508,N_410);
or U1219 (N_1219,N_616,In_2318);
or U1220 (N_1220,N_615,In_1929);
and U1221 (N_1221,N_683,In_312);
and U1222 (N_1222,In_2916,In_1699);
or U1223 (N_1223,In_1129,In_2521);
or U1224 (N_1224,In_2875,N_295);
nand U1225 (N_1225,N_83,N_757);
nor U1226 (N_1226,N_638,In_1133);
nor U1227 (N_1227,N_695,In_774);
xor U1228 (N_1228,In_2460,In_2935);
nand U1229 (N_1229,N_241,In_2095);
nand U1230 (N_1230,In_2415,N_953);
nor U1231 (N_1231,In_2394,N_640);
or U1232 (N_1232,In_1047,N_771);
nor U1233 (N_1233,In_1746,N_164);
or U1234 (N_1234,N_680,N_469);
xor U1235 (N_1235,In_1499,N_855);
or U1236 (N_1236,In_2542,In_2376);
nand U1237 (N_1237,N_976,N_256);
or U1238 (N_1238,In_722,N_124);
nor U1239 (N_1239,In_2953,In_1201);
and U1240 (N_1240,In_2155,N_372);
xnor U1241 (N_1241,In_317,In_2750);
xnor U1242 (N_1242,N_803,N_577);
and U1243 (N_1243,N_538,In_504);
nor U1244 (N_1244,In_1598,In_1190);
xor U1245 (N_1245,N_457,N_303);
xnor U1246 (N_1246,In_2952,In_105);
nand U1247 (N_1247,N_784,N_721);
nand U1248 (N_1248,N_986,In_763);
xnor U1249 (N_1249,In_2558,In_993);
nand U1250 (N_1250,N_552,N_536);
or U1251 (N_1251,N_594,N_905);
nor U1252 (N_1252,In_1603,In_917);
nand U1253 (N_1253,In_363,In_1543);
xor U1254 (N_1254,N_106,N_37);
nor U1255 (N_1255,In_241,N_370);
or U1256 (N_1256,N_631,N_18);
or U1257 (N_1257,In_1761,N_250);
nand U1258 (N_1258,In_332,N_940);
nand U1259 (N_1259,In_873,In_532);
and U1260 (N_1260,N_503,In_510);
or U1261 (N_1261,N_228,In_1279);
and U1262 (N_1262,N_82,N_268);
or U1263 (N_1263,In_1707,In_829);
nand U1264 (N_1264,N_524,N_929);
nor U1265 (N_1265,N_210,In_2968);
or U1266 (N_1266,In_2085,In_2718);
xnor U1267 (N_1267,In_2134,In_845);
nor U1268 (N_1268,N_48,N_530);
xor U1269 (N_1269,In_47,N_772);
nor U1270 (N_1270,In_653,In_1353);
or U1271 (N_1271,In_758,N_149);
xnor U1272 (N_1272,In_1698,In_1195);
and U1273 (N_1273,In_1027,N_292);
nor U1274 (N_1274,In_2786,N_206);
nor U1275 (N_1275,N_641,N_663);
and U1276 (N_1276,N_403,In_490);
xor U1277 (N_1277,N_280,N_507);
or U1278 (N_1278,N_686,In_2162);
and U1279 (N_1279,In_2040,N_522);
nor U1280 (N_1280,N_41,In_1208);
or U1281 (N_1281,N_924,N_642);
and U1282 (N_1282,N_596,In_1392);
nand U1283 (N_1283,In_472,In_1341);
and U1284 (N_1284,N_408,In_1716);
or U1285 (N_1285,N_184,In_2806);
nor U1286 (N_1286,N_851,In_2426);
nor U1287 (N_1287,In_2871,In_1393);
and U1288 (N_1288,In_102,In_930);
nand U1289 (N_1289,N_60,In_2454);
or U1290 (N_1290,In_1210,In_2797);
or U1291 (N_1291,N_999,In_1232);
or U1292 (N_1292,In_949,N_133);
or U1293 (N_1293,In_2223,N_341);
or U1294 (N_1294,In_398,In_2996);
or U1295 (N_1295,N_736,In_2645);
nand U1296 (N_1296,N_17,N_690);
nand U1297 (N_1297,N_367,N_113);
nand U1298 (N_1298,In_1061,In_1562);
nand U1299 (N_1299,In_789,N_25);
xor U1300 (N_1300,In_2492,N_990);
xnor U1301 (N_1301,In_180,N_105);
or U1302 (N_1302,In_1130,In_2889);
nand U1303 (N_1303,In_2838,N_618);
nand U1304 (N_1304,N_87,N_388);
nor U1305 (N_1305,N_836,N_441);
or U1306 (N_1306,In_1266,In_1235);
nor U1307 (N_1307,N_563,N_382);
or U1308 (N_1308,In_2734,In_2259);
and U1309 (N_1309,N_588,N_897);
xnor U1310 (N_1310,In_1141,In_502);
nand U1311 (N_1311,In_168,N_311);
and U1312 (N_1312,N_489,N_608);
and U1313 (N_1313,In_640,In_444);
nor U1314 (N_1314,N_151,In_1299);
nand U1315 (N_1315,In_1949,N_249);
and U1316 (N_1316,In_364,In_2064);
nand U1317 (N_1317,In_1489,In_794);
and U1318 (N_1318,In_1473,N_77);
or U1319 (N_1319,In_2591,N_57);
nand U1320 (N_1320,N_248,N_46);
nand U1321 (N_1321,In_648,N_647);
or U1322 (N_1322,N_604,N_674);
xnor U1323 (N_1323,N_260,N_176);
nand U1324 (N_1324,N_1,N_11);
and U1325 (N_1325,In_563,N_499);
xor U1326 (N_1326,In_1340,N_520);
and U1327 (N_1327,N_309,N_3);
nor U1328 (N_1328,N_935,In_808);
and U1329 (N_1329,N_393,N_381);
and U1330 (N_1330,N_70,N_706);
and U1331 (N_1331,In_598,In_588);
nor U1332 (N_1332,In_378,N_415);
xnor U1333 (N_1333,N_326,N_273);
xnor U1334 (N_1334,In_2507,In_2358);
or U1335 (N_1335,In_573,N_390);
and U1336 (N_1336,N_459,N_247);
nand U1337 (N_1337,N_127,In_1571);
nand U1338 (N_1338,In_302,In_2980);
nor U1339 (N_1339,In_2634,In_2769);
or U1340 (N_1340,In_1819,N_657);
nor U1341 (N_1341,N_463,N_224);
or U1342 (N_1342,In_1514,N_496);
nor U1343 (N_1343,N_61,N_982);
nor U1344 (N_1344,In_646,In_2220);
nor U1345 (N_1345,In_2518,In_1711);
and U1346 (N_1346,In_39,In_223);
nand U1347 (N_1347,In_237,N_865);
xnor U1348 (N_1348,In_279,N_484);
and U1349 (N_1349,In_2872,In_2246);
or U1350 (N_1350,N_40,In_2803);
and U1351 (N_1351,In_1896,In_2122);
and U1352 (N_1352,N_961,In_961);
xnor U1353 (N_1353,In_2920,In_311);
xnor U1354 (N_1354,N_125,N_767);
or U1355 (N_1355,In_1022,N_662);
or U1356 (N_1356,In_846,In_1442);
and U1357 (N_1357,In_2602,In_978);
nor U1358 (N_1358,N_523,N_108);
and U1359 (N_1359,In_1770,In_1548);
nand U1360 (N_1360,In_2906,In_1445);
or U1361 (N_1361,In_740,N_894);
or U1362 (N_1362,N_872,N_110);
nor U1363 (N_1363,In_1163,N_383);
and U1364 (N_1364,N_997,In_704);
xor U1365 (N_1365,N_705,In_170);
and U1366 (N_1366,In_594,N_212);
nand U1367 (N_1367,N_407,In_658);
xnor U1368 (N_1368,N_201,N_835);
nor U1369 (N_1369,N_727,In_2184);
nand U1370 (N_1370,N_447,In_491);
and U1371 (N_1371,In_608,In_2625);
xnor U1372 (N_1372,In_2206,N_610);
or U1373 (N_1373,In_196,N_827);
or U1374 (N_1374,N_340,In_911);
nor U1375 (N_1375,N_483,In_255);
or U1376 (N_1376,In_1403,N_413);
nand U1377 (N_1377,In_1883,N_183);
and U1378 (N_1378,N_239,N_422);
nand U1379 (N_1379,N_913,N_816);
and U1380 (N_1380,In_816,In_1185);
and U1381 (N_1381,In_2742,N_494);
and U1382 (N_1382,N_729,N_198);
and U1383 (N_1383,N_895,N_159);
xor U1384 (N_1384,In_2321,N_373);
nor U1385 (N_1385,N_700,In_577);
and U1386 (N_1386,In_322,N_715);
nor U1387 (N_1387,In_622,In_1915);
and U1388 (N_1388,N_668,In_1560);
or U1389 (N_1389,N_926,In_2495);
or U1390 (N_1390,N_375,In_143);
and U1391 (N_1391,N_831,In_1532);
xor U1392 (N_1392,N_587,In_2944);
and U1393 (N_1393,In_2493,In_1365);
xnor U1394 (N_1394,In_1059,N_864);
nor U1395 (N_1395,N_424,In_2823);
xnor U1396 (N_1396,N_139,In_2646);
and U1397 (N_1397,N_336,In_630);
xnor U1398 (N_1398,In_1226,In_2213);
xor U1399 (N_1399,In_1119,N_977);
and U1400 (N_1400,N_991,N_274);
nand U1401 (N_1401,In_1107,In_2329);
xnor U1402 (N_1402,N_584,In_2222);
nor U1403 (N_1403,In_393,In_997);
and U1404 (N_1404,N_993,In_1329);
and U1405 (N_1405,In_801,N_925);
xnor U1406 (N_1406,N_811,N_586);
xnor U1407 (N_1407,In_1979,In_1289);
and U1408 (N_1408,N_128,N_569);
and U1409 (N_1409,N_626,N_556);
xor U1410 (N_1410,In_1144,In_41);
and U1411 (N_1411,In_1822,In_366);
nor U1412 (N_1412,In_1072,N_271);
nor U1413 (N_1413,In_1117,N_490);
nor U1414 (N_1414,In_2090,N_541);
nand U1415 (N_1415,In_2383,N_623);
xor U1416 (N_1416,N_847,In_1344);
or U1417 (N_1417,N_739,In_2905);
nand U1418 (N_1418,In_886,In_778);
nand U1419 (N_1419,In_2813,In_631);
nor U1420 (N_1420,In_1112,In_1539);
nor U1421 (N_1421,N_364,In_477);
xnor U1422 (N_1422,In_607,N_857);
xor U1423 (N_1423,N_766,N_887);
nor U1424 (N_1424,In_2540,In_465);
xor U1425 (N_1425,N_211,N_443);
and U1426 (N_1426,N_701,In_2921);
nor U1427 (N_1427,N_157,In_1662);
nand U1428 (N_1428,N_470,In_303);
nand U1429 (N_1429,In_516,In_2835);
and U1430 (N_1430,In_751,N_513);
and U1431 (N_1431,In_288,N_305);
and U1432 (N_1432,In_2136,N_315);
nor U1433 (N_1433,In_860,In_456);
nand U1434 (N_1434,In_1892,N_808);
nor U1435 (N_1435,In_827,N_965);
xor U1436 (N_1436,N_871,In_2981);
or U1437 (N_1437,N_191,N_597);
or U1438 (N_1438,In_1980,In_2698);
and U1439 (N_1439,N_846,N_884);
nor U1440 (N_1440,N_532,In_2466);
nor U1441 (N_1441,N_220,In_979);
and U1442 (N_1442,In_134,N_26);
or U1443 (N_1443,In_725,N_775);
nor U1444 (N_1444,N_599,In_300);
nand U1445 (N_1445,In_2537,N_285);
nor U1446 (N_1446,In_2,N_967);
or U1447 (N_1447,N_78,In_768);
nand U1448 (N_1448,N_302,In_2777);
nor U1449 (N_1449,In_2530,N_768);
xnor U1450 (N_1450,In_2302,N_916);
xnor U1451 (N_1451,In_2041,In_1991);
xnor U1452 (N_1452,N_675,N_743);
nand U1453 (N_1453,N_528,In_104);
nor U1454 (N_1454,N_468,N_51);
nand U1455 (N_1455,In_1766,In_2281);
nand U1456 (N_1456,In_1763,N_172);
and U1457 (N_1457,N_854,In_351);
nor U1458 (N_1458,In_2299,In_13);
and U1459 (N_1459,N_229,N_451);
xor U1460 (N_1460,In_1815,In_32);
xor U1461 (N_1461,In_840,N_317);
nor U1462 (N_1462,In_1155,N_759);
xnor U1463 (N_1463,In_996,N_12);
nand U1464 (N_1464,In_1592,N_369);
and U1465 (N_1465,In_2463,N_876);
nor U1466 (N_1466,In_1292,In_1924);
and U1467 (N_1467,N_288,In_1840);
nor U1468 (N_1468,In_2411,In_1898);
nor U1469 (N_1469,In_2693,N_349);
nand U1470 (N_1470,In_445,In_2282);
nand U1471 (N_1471,In_2308,In_534);
nand U1472 (N_1472,N_852,In_357);
xnor U1473 (N_1473,In_292,In_2515);
and U1474 (N_1474,N_933,N_445);
or U1475 (N_1475,N_972,N_380);
or U1476 (N_1476,In_1237,N_752);
or U1477 (N_1477,N_637,In_1132);
and U1478 (N_1478,In_797,In_600);
nand U1479 (N_1479,In_2637,N_435);
or U1480 (N_1480,N_707,N_158);
xor U1481 (N_1481,N_434,In_1269);
xnor U1482 (N_1482,N_745,In_1818);
nor U1483 (N_1483,N_261,N_810);
nor U1484 (N_1484,N_716,In_2430);
and U1485 (N_1485,In_1518,In_2044);
or U1486 (N_1486,In_2355,N_833);
or U1487 (N_1487,N_778,In_235);
nor U1488 (N_1488,In_1824,N_366);
or U1489 (N_1489,N_754,N_515);
or U1490 (N_1490,In_439,N_116);
nand U1491 (N_1491,N_414,In_2860);
nor U1492 (N_1492,N_512,N_733);
and U1493 (N_1493,In_1359,N_891);
nor U1494 (N_1494,N_714,N_103);
or U1495 (N_1495,N_225,In_1327);
nor U1496 (N_1496,In_120,In_2150);
or U1497 (N_1497,In_1136,N_437);
or U1498 (N_1498,In_2197,N_837);
nand U1499 (N_1499,N_892,In_2808);
nor U1500 (N_1500,In_2571,In_1524);
xor U1501 (N_1501,N_186,In_2533);
or U1502 (N_1502,N_724,N_337);
nor U1503 (N_1503,N_74,N_781);
xnor U1504 (N_1504,In_2559,In_1265);
nor U1505 (N_1505,N_567,In_982);
and U1506 (N_1506,N_779,In_2333);
and U1507 (N_1507,In_803,In_1294);
nor U1508 (N_1508,N_801,In_2572);
nor U1509 (N_1509,In_958,N_840);
nor U1510 (N_1510,In_2303,In_1169);
and U1511 (N_1511,In_1212,In_1620);
nand U1512 (N_1512,N_673,N_75);
xnor U1513 (N_1513,N_956,In_1708);
and U1514 (N_1514,In_2581,In_1111);
nor U1515 (N_1515,N_475,N_568);
xnor U1516 (N_1516,In_341,In_655);
and U1517 (N_1517,N_537,N_572);
nand U1518 (N_1518,N_566,In_44);
xnor U1519 (N_1519,In_1101,N_19);
xnor U1520 (N_1520,N_452,N_85);
and U1521 (N_1521,In_354,In_1032);
and U1522 (N_1522,N_34,N_653);
nor U1523 (N_1523,N_49,N_267);
or U1524 (N_1524,N_861,N_352);
or U1525 (N_1525,N_356,N_333);
or U1526 (N_1526,N_88,N_284);
nor U1527 (N_1527,In_231,N_476);
xor U1528 (N_1528,N_207,In_396);
and U1529 (N_1529,N_521,In_2176);
or U1530 (N_1530,N_930,N_495);
nor U1531 (N_1531,N_14,N_163);
xor U1532 (N_1532,In_2051,N_455);
xor U1533 (N_1533,N_963,N_92);
and U1534 (N_1534,N_770,N_258);
nor U1535 (N_1535,In_1935,N_141);
and U1536 (N_1536,N_122,N_777);
nand U1537 (N_1537,In_1861,In_219);
nand U1538 (N_1538,N_148,N_180);
or U1539 (N_1539,N_900,In_2385);
xor U1540 (N_1540,N_244,In_446);
nand U1541 (N_1541,In_2171,In_1263);
nor U1542 (N_1542,In_2802,In_286);
nand U1543 (N_1543,In_757,N_555);
nand U1544 (N_1544,In_318,N_889);
or U1545 (N_1545,N_901,In_915);
nand U1546 (N_1546,N_671,N_281);
nand U1547 (N_1547,N_446,N_794);
nand U1548 (N_1548,In_2497,N_449);
nand U1549 (N_1549,In_2029,In_149);
and U1550 (N_1550,In_1879,N_585);
nand U1551 (N_1551,N_658,In_2089);
and U1552 (N_1552,N_829,N_602);
nor U1553 (N_1553,In_1749,N_710);
nor U1554 (N_1554,N_91,N_235);
nand U1555 (N_1555,In_1895,In_857);
and U1556 (N_1556,N_959,N_817);
or U1557 (N_1557,In_2749,In_703);
or U1558 (N_1558,In_2238,N_205);
nor U1559 (N_1559,N_878,N_400);
nand U1560 (N_1560,In_2201,N_888);
or U1561 (N_1561,In_1519,N_150);
nand U1562 (N_1562,N_97,N_971);
nor U1563 (N_1563,In_733,N_651);
nor U1564 (N_1564,In_2867,In_847);
nor U1565 (N_1565,N_473,N_509);
and U1566 (N_1566,In_724,N_101);
xnor U1567 (N_1567,In_1453,In_2684);
and U1568 (N_1568,N_800,N_300);
nor U1569 (N_1569,In_144,In_688);
or U1570 (N_1570,In_401,N_687);
xnor U1571 (N_1571,In_2596,N_44);
or U1572 (N_1572,In_1565,N_129);
xor U1573 (N_1573,In_2187,In_277);
xnor U1574 (N_1574,N_153,In_1890);
or U1575 (N_1575,N_43,N_709);
nor U1576 (N_1576,N_958,In_1177);
xor U1577 (N_1577,N_177,N_118);
and U1578 (N_1578,N_282,In_2595);
or U1579 (N_1579,In_1878,In_2593);
and U1580 (N_1580,N_15,N_365);
or U1581 (N_1581,In_1586,In_560);
nor U1582 (N_1582,In_555,In_2262);
xor U1583 (N_1583,N_763,N_987);
nand U1584 (N_1584,In_2649,N_731);
and U1585 (N_1585,In_902,N_195);
nor U1586 (N_1586,In_2337,N_983);
and U1587 (N_1587,In_1712,N_278);
xor U1588 (N_1588,N_209,In_227);
nor U1589 (N_1589,In_2012,N_80);
nor U1590 (N_1590,In_527,In_2881);
xnor U1591 (N_1591,In_1673,In_2014);
nand U1592 (N_1592,In_1550,In_2592);
nand U1593 (N_1593,N_33,In_1669);
nor U1594 (N_1594,In_2868,N_160);
nand U1595 (N_1595,N_348,In_2901);
or U1596 (N_1596,In_1159,N_598);
and U1597 (N_1597,In_2733,N_946);
or U1598 (N_1598,N_517,N_137);
and U1599 (N_1599,In_1354,N_868);
or U1600 (N_1600,In_1795,N_199);
xor U1601 (N_1601,N_314,In_54);
xor U1602 (N_1602,N_226,In_822);
nor U1603 (N_1603,In_814,In_2013);
and U1604 (N_1604,In_2467,In_319);
nor U1605 (N_1605,In_1675,N_442);
nand U1606 (N_1606,N_385,N_576);
nand U1607 (N_1607,N_136,N_699);
nand U1608 (N_1608,N_860,In_2055);
and U1609 (N_1609,N_374,N_650);
or U1610 (N_1610,In_800,N_126);
nor U1611 (N_1611,In_1784,N_479);
or U1612 (N_1612,In_1179,In_425);
and U1613 (N_1613,In_2994,In_1788);
xor U1614 (N_1614,In_1575,In_2275);
xnor U1615 (N_1615,N_698,In_2481);
xnor U1616 (N_1616,N_156,In_2164);
or U1617 (N_1617,N_170,N_797);
nor U1618 (N_1618,In_619,N_818);
or U1619 (N_1619,N_968,In_16);
or U1620 (N_1620,In_2919,N_902);
xor U1621 (N_1621,N_603,N_335);
or U1622 (N_1622,N_992,N_676);
nor U1623 (N_1623,N_140,N_546);
xnor U1624 (N_1624,N_877,N_922);
xor U1625 (N_1625,N_917,N_646);
and U1626 (N_1626,N_750,In_1131);
nand U1627 (N_1627,N_669,N_746);
xnor U1628 (N_1628,N_196,N_948);
or U1629 (N_1629,N_96,N_685);
xnor U1630 (N_1630,In_1958,N_107);
nor U1631 (N_1631,In_1245,In_101);
or U1632 (N_1632,N_277,N_764);
and U1633 (N_1633,N_960,In_1778);
nand U1634 (N_1634,N_392,N_301);
xnor U1635 (N_1635,N_93,In_2181);
or U1636 (N_1636,N_438,In_2651);
nand U1637 (N_1637,In_1222,In_1637);
nor U1638 (N_1638,N_732,N_290);
and U1639 (N_1639,In_1496,In_1382);
xor U1640 (N_1640,N_68,N_397);
or U1641 (N_1641,N_351,N_670);
and U1642 (N_1642,N_138,In_895);
nor U1643 (N_1643,N_579,N_542);
nor U1644 (N_1644,In_973,N_448);
or U1645 (N_1645,N_279,N_822);
or U1646 (N_1646,N_423,N_276);
nand U1647 (N_1647,N_84,N_881);
nand U1648 (N_1648,N_762,N_823);
nor U1649 (N_1649,N_478,N_8);
or U1650 (N_1650,In_1735,In_960);
or U1651 (N_1651,In_1298,N_21);
and U1652 (N_1652,In_1270,In_2081);
nor U1653 (N_1653,N_918,N_242);
xnor U1654 (N_1654,N_882,N_289);
nand U1655 (N_1655,N_502,In_832);
nor U1656 (N_1656,In_2193,In_891);
xnor U1657 (N_1657,In_1012,N_234);
nand U1658 (N_1658,In_1348,N_919);
nor U1659 (N_1659,N_702,In_1646);
xor U1660 (N_1660,In_1358,N_863);
nand U1661 (N_1661,N_786,N_474);
nor U1662 (N_1662,N_52,In_148);
nand U1663 (N_1663,In_2378,In_1976);
and U1664 (N_1664,In_1681,N_580);
or U1665 (N_1665,In_693,N_332);
nand U1666 (N_1666,In_2485,N_879);
nand U1667 (N_1667,N_540,In_45);
xor U1668 (N_1668,In_615,In_2335);
xnor U1669 (N_1669,In_1983,N_561);
xnor U1670 (N_1670,N_2,N_353);
or U1671 (N_1671,N_213,In_1764);
or U1672 (N_1672,In_1859,N_6);
nand U1673 (N_1673,N_308,In_2550);
or U1674 (N_1674,N_697,N_873);
or U1675 (N_1675,N_90,N_628);
nor U1676 (N_1676,In_736,N_593);
xor U1677 (N_1677,In_424,N_218);
xor U1678 (N_1678,N_550,In_389);
xor U1679 (N_1679,N_549,In_2721);
nor U1680 (N_1680,N_534,N_545);
or U1681 (N_1681,In_2610,N_984);
and U1682 (N_1682,In_2153,In_1110);
nand U1683 (N_1683,N_426,In_298);
or U1684 (N_1684,In_945,N_964);
xnor U1685 (N_1685,In_2554,In_2199);
nand U1686 (N_1686,In_458,N_909);
or U1687 (N_1687,In_738,In_968);
nand U1688 (N_1688,N_634,In_1483);
or U1689 (N_1689,In_2002,In_1642);
nor U1690 (N_1690,In_431,In_270);
nand U1691 (N_1691,N_283,N_161);
xor U1692 (N_1692,N_760,N_197);
xor U1693 (N_1693,In_2140,In_2469);
nand U1694 (N_1694,N_740,N_439);
nand U1695 (N_1695,N_906,In_1293);
nand U1696 (N_1696,In_251,In_743);
and U1697 (N_1697,N_323,In_377);
xnor U1698 (N_1698,In_906,N_730);
nand U1699 (N_1699,N_969,In_2852);
xnor U1700 (N_1700,N_862,In_669);
and U1701 (N_1701,In_2993,In_793);
or U1702 (N_1702,N_547,N_269);
xor U1703 (N_1703,In_433,N_531);
and U1704 (N_1704,In_1992,In_2846);
and U1705 (N_1705,In_1305,In_2365);
xnor U1706 (N_1706,N_259,N_665);
nor U1707 (N_1707,In_2695,In_901);
nor U1708 (N_1708,N_386,In_2020);
nand U1709 (N_1709,N_574,In_320);
nand U1710 (N_1710,In_1522,N_722);
and U1711 (N_1711,N_418,N_232);
and U1712 (N_1712,In_1786,In_2080);
and U1713 (N_1713,In_2516,In_1192);
nor U1714 (N_1714,In_245,In_73);
and U1715 (N_1715,N_622,N_923);
or U1716 (N_1716,In_1997,In_1783);
nand U1717 (N_1717,In_55,N_735);
nand U1718 (N_1718,In_1173,In_1431);
or U1719 (N_1719,In_201,In_606);
or U1720 (N_1720,N_498,In_2614);
nand U1721 (N_1721,N_807,In_2882);
and U1722 (N_1722,In_2601,N_325);
nand U1723 (N_1723,N_893,In_2513);
nand U1724 (N_1724,N_378,In_541);
xor U1725 (N_1725,In_1844,N_630);
nor U1726 (N_1726,N_491,In_1622);
and U1727 (N_1727,In_2462,In_1436);
nor U1728 (N_1728,N_834,In_355);
or U1729 (N_1729,In_856,In_578);
or U1730 (N_1730,N_320,N_67);
nand U1731 (N_1731,N_849,In_970);
nor U1732 (N_1732,In_256,N_554);
xor U1733 (N_1733,In_290,N_624);
nand U1734 (N_1734,In_2683,N_853);
or U1735 (N_1735,N_430,In_391);
xnor U1736 (N_1736,In_890,N_886);
nand U1737 (N_1737,N_780,In_1338);
nor U1738 (N_1738,N_819,N_472);
nand U1739 (N_1739,In_2836,N_245);
nand U1740 (N_1740,In_2829,In_920);
and U1741 (N_1741,N_617,In_1140);
or U1742 (N_1742,N_501,In_2608);
nor U1743 (N_1743,In_762,In_2328);
or U1744 (N_1744,In_2927,In_2456);
and U1745 (N_1745,N_464,N_809);
nand U1746 (N_1746,N_493,In_2244);
nand U1747 (N_1747,N_440,N_420);
and U1748 (N_1748,N_694,N_578);
xnor U1749 (N_1749,N_178,N_0);
or U1750 (N_1750,N_42,N_805);
nand U1751 (N_1751,N_219,In_2694);
and U1752 (N_1752,In_1630,In_1182);
or U1753 (N_1753,N_664,In_2983);
or U1754 (N_1754,In_2354,N_405);
nor U1755 (N_1755,N_321,In_1402);
and U1756 (N_1756,N_828,In_881);
xor U1757 (N_1757,In_769,N_989);
and U1758 (N_1758,In_67,N_799);
xor U1759 (N_1759,N_848,N_179);
nor U1760 (N_1760,In_1310,In_1157);
nand U1761 (N_1761,N_527,N_519);
nand U1762 (N_1762,N_24,In_2828);
xnor U1763 (N_1763,N_793,N_866);
nor U1764 (N_1764,In_811,N_387);
and U1765 (N_1765,In_2049,N_456);
nor U1766 (N_1766,In_2668,N_319);
nand U1767 (N_1767,N_841,N_264);
or U1768 (N_1768,In_1977,N_824);
and U1769 (N_1769,N_785,N_32);
xor U1770 (N_1770,N_22,In_680);
nand U1771 (N_1771,In_485,N_995);
xnor U1772 (N_1772,N_996,In_1440);
nor U1773 (N_1773,In_1011,In_2892);
or U1774 (N_1774,In_1428,N_947);
and U1775 (N_1775,In_2761,N_559);
nor U1776 (N_1776,N_516,N_30);
or U1777 (N_1777,In_556,N_313);
nor U1778 (N_1778,N_192,In_1308);
and U1779 (N_1779,In_2866,In_1186);
nand U1780 (N_1780,In_1143,In_2809);
nand U1781 (N_1781,N_514,In_1792);
or U1782 (N_1782,In_2372,N_792);
or U1783 (N_1783,N_227,N_954);
or U1784 (N_1784,In_2152,N_230);
and U1785 (N_1785,N_488,In_470);
nor U1786 (N_1786,N_756,N_691);
nor U1787 (N_1787,In_2873,N_98);
xor U1788 (N_1788,In_2696,N_844);
nand U1789 (N_1789,N_907,N_688);
or U1790 (N_1790,In_1377,In_299);
nand U1791 (N_1791,In_837,N_962);
nand U1792 (N_1792,N_36,In_509);
nand U1793 (N_1793,N_20,N_204);
xor U1794 (N_1794,N_589,N_361);
and U1795 (N_1795,N_689,In_2978);
nor U1796 (N_1796,N_266,N_368);
or U1797 (N_1797,N_915,N_202);
nor U1798 (N_1798,In_2441,In_679);
or U1799 (N_1799,In_1096,In_1814);
or U1800 (N_1800,In_1484,In_1307);
xor U1801 (N_1801,N_635,N_737);
nor U1802 (N_1802,N_427,N_329);
and U1803 (N_1803,N_162,In_1224);
or U1804 (N_1804,N_263,N_399);
or U1805 (N_1805,N_684,In_941);
xnor U1806 (N_1806,N_465,N_316);
nor U1807 (N_1807,N_518,N_240);
or U1808 (N_1808,N_359,N_143);
nand U1809 (N_1809,In_369,N_821);
nor U1810 (N_1810,In_416,N_5);
nor U1811 (N_1811,N_55,In_2679);
and U1812 (N_1812,In_1441,N_652);
or U1813 (N_1813,N_38,N_966);
or U1814 (N_1814,N_217,In_463);
nor U1815 (N_1815,In_1876,In_2084);
or U1816 (N_1816,In_2714,N_253);
or U1817 (N_1817,N_874,N_773);
or U1818 (N_1818,In_2120,In_1037);
xor U1819 (N_1819,In_1969,In_2183);
and U1820 (N_1820,In_2145,In_1654);
or U1821 (N_1821,N_102,In_1194);
or U1822 (N_1822,N_791,N_343);
nand U1823 (N_1823,N_358,N_109);
and U1824 (N_1824,In_715,In_528);
xnor U1825 (N_1825,N_741,N_485);
nand U1826 (N_1826,N_927,In_2691);
or U1827 (N_1827,N_557,N_582);
xor U1828 (N_1828,In_2092,N_945);
nor U1829 (N_1829,In_1835,In_2567);
and U1830 (N_1830,In_457,N_142);
nor U1831 (N_1831,In_1196,In_914);
nand U1832 (N_1832,In_394,N_404);
nor U1833 (N_1833,In_2031,In_2121);
nor U1834 (N_1834,N_952,N_979);
nand U1835 (N_1835,In_1693,N_221);
or U1836 (N_1836,N_813,In_176);
or U1837 (N_1837,In_99,In_2257);
nor U1838 (N_1838,In_2895,In_1229);
xnor U1839 (N_1839,In_2778,N_185);
nand U1840 (N_1840,N_181,In_115);
nand U1841 (N_1841,In_385,In_135);
nor U1842 (N_1842,N_704,In_599);
or U1843 (N_1843,N_28,N_609);
or U1844 (N_1844,In_1648,N_858);
xor U1845 (N_1845,In_1315,N_169);
nand U1846 (N_1846,N_402,N_89);
xor U1847 (N_1847,N_193,In_2720);
or U1848 (N_1848,N_832,N_806);
nor U1849 (N_1849,N_920,N_654);
or U1850 (N_1850,In_109,N_850);
nor U1851 (N_1851,N_389,In_2349);
nand U1852 (N_1852,In_1209,In_883);
or U1853 (N_1853,In_1686,N_10);
xnor U1854 (N_1854,In_2735,In_1555);
or U1855 (N_1855,In_2414,N_633);
and U1856 (N_1856,N_471,In_1512);
or U1857 (N_1857,In_2965,N_376);
nor U1858 (N_1858,N_208,N_377);
or U1859 (N_1859,N_681,In_756);
and U1860 (N_1860,In_664,In_2045);
or U1861 (N_1861,In_897,In_2300);
or U1862 (N_1862,In_1493,In_495);
or U1863 (N_1863,N_461,In_2033);
and U1864 (N_1864,In_2945,N_237);
nor U1865 (N_1865,In_1351,In_1845);
nor U1866 (N_1866,N_27,N_985);
or U1867 (N_1867,N_789,N_583);
xor U1868 (N_1868,In_1756,In_695);
xnor U1869 (N_1869,In_1188,In_2656);
xnor U1870 (N_1870,In_268,In_1759);
xnor U1871 (N_1871,In_2912,N_119);
and U1872 (N_1872,In_2969,In_2215);
xor U1873 (N_1873,N_590,N_460);
nand U1874 (N_1874,N_738,N_696);
nor U1875 (N_1875,N_601,N_406);
and U1876 (N_1876,In_805,N_911);
nand U1877 (N_1877,N_147,N_720);
xor U1878 (N_1878,N_111,In_2682);
or U1879 (N_1879,N_296,In_2688);
nand U1880 (N_1880,N_734,N_293);
nor U1881 (N_1881,In_236,In_2129);
or U1882 (N_1882,N_350,N_544);
or U1883 (N_1883,In_1038,N_66);
xnor U1884 (N_1884,N_73,In_2362);
and U1885 (N_1885,In_923,N_431);
xor U1886 (N_1886,In_2458,N_328);
or U1887 (N_1887,In_1593,In_261);
and U1888 (N_1888,N_482,In_2816);
nand U1889 (N_1889,In_2339,In_2143);
nand U1890 (N_1890,In_114,N_591);
xor U1891 (N_1891,N_355,In_2435);
nor U1892 (N_1892,In_2270,In_1057);
and U1893 (N_1893,N_611,In_1283);
xnor U1894 (N_1894,In_710,N_384);
nor U1895 (N_1895,In_1529,In_49);
nor U1896 (N_1896,N_830,N_815);
nor U1897 (N_1897,In_2427,In_2445);
and U1898 (N_1898,N_318,N_936);
nor U1899 (N_1899,In_2261,In_1546);
and U1900 (N_1900,In_2325,N_820);
nor U1901 (N_1901,In_2939,In_383);
nand U1902 (N_1902,N_747,N_551);
nand U1903 (N_1903,N_270,In_1147);
xnor U1904 (N_1904,N_944,In_1638);
xnor U1905 (N_1905,In_962,In_2468);
nand U1906 (N_1906,N_612,N_182);
and U1907 (N_1907,N_678,In_260);
nor U1908 (N_1908,In_64,In_1503);
or U1909 (N_1909,N_429,N_570);
xor U1910 (N_1910,In_1837,In_518);
and U1911 (N_1911,In_240,In_1922);
xor U1912 (N_1912,N_553,N_713);
nand U1913 (N_1913,In_1998,In_861);
or U1914 (N_1914,N_255,In_2747);
and U1915 (N_1915,In_2144,N_306);
or U1916 (N_1916,In_632,In_2284);
nand U1917 (N_1917,N_342,N_500);
xnor U1918 (N_1918,N_928,In_2224);
and U1919 (N_1919,N_914,In_407);
nor U1920 (N_1920,In_2821,N_751);
or U1921 (N_1921,In_395,N_433);
or U1922 (N_1922,In_1816,N_667);
nor U1923 (N_1923,In_1161,N_974);
nor U1924 (N_1924,In_2240,N_480);
or U1925 (N_1925,N_409,N_453);
xor U1926 (N_1926,N_486,In_1225);
nand U1927 (N_1927,In_2573,N_458);
nor U1928 (N_1928,N_173,N_286);
and U1929 (N_1929,N_100,N_331);
nor U1930 (N_1930,In_422,N_883);
or U1931 (N_1931,N_254,In_2075);
or U1932 (N_1932,N_171,In_2755);
or U1933 (N_1933,N_749,N_371);
xnor U1934 (N_1934,In_1682,In_2536);
nor U1935 (N_1935,In_590,N_742);
and U1936 (N_1936,N_357,In_158);
nor U1937 (N_1937,N_938,N_950);
xnor U1938 (N_1938,In_1097,In_2196);
xor U1939 (N_1939,N_758,In_28);
xor U1940 (N_1940,N_53,In_1467);
nand U1941 (N_1941,In_971,N_644);
xor U1942 (N_1942,In_452,N_804);
nor U1943 (N_1943,In_79,N_238);
nand U1944 (N_1944,N_994,In_183);
xor U1945 (N_1945,N_875,In_1615);
and U1946 (N_1946,In_2490,In_2850);
and U1947 (N_1947,In_2423,In_671);
or U1948 (N_1948,In_468,N_354);
xnor U1949 (N_1949,N_679,In_853);
and U1950 (N_1950,N_573,In_1600);
xor U1951 (N_1951,In_1884,N_379);
or U1952 (N_1952,N_643,N_921);
nor U1953 (N_1953,In_449,N_360);
or U1954 (N_1954,N_998,In_2091);
xnor U1955 (N_1955,In_2305,In_2869);
nor U1956 (N_1956,N_636,In_746);
nand U1957 (N_1957,N_168,In_1425);
xor U1958 (N_1958,N_251,N_307);
xnor U1959 (N_1959,N_362,N_327);
xor U1960 (N_1960,In_1501,In_2955);
nand U1961 (N_1961,N_896,N_755);
nor U1962 (N_1962,In_2131,N_798);
nand U1963 (N_1963,N_869,In_2923);
nand U1964 (N_1964,In_2743,N_627);
or U1965 (N_1965,In_683,N_620);
nand U1966 (N_1966,N_252,N_753);
nand U1967 (N_1967,In_4,N_867);
nand U1968 (N_1968,In_2503,N_396);
nand U1969 (N_1969,N_155,N_262);
nand U1970 (N_1970,In_2655,In_1933);
xor U1971 (N_1971,In_1900,In_82);
nand U1972 (N_1972,In_186,N_508);
and U1973 (N_1973,In_2790,In_2283);
xnor U1974 (N_1974,N_600,N_744);
and U1975 (N_1975,In_2388,In_2449);
or U1976 (N_1976,N_632,In_2510);
xnor U1977 (N_1977,In_530,In_70);
xnor U1978 (N_1978,N_672,In_1044);
nor U1979 (N_1979,N_246,In_1553);
xnor U1980 (N_1980,In_2158,In_2066);
and U1981 (N_1981,N_941,In_2929);
nor U1982 (N_1982,In_20,N_723);
or U1983 (N_1983,In_25,In_2118);
and U1984 (N_1984,N_86,N_870);
or U1985 (N_1985,In_584,N_769);
nor U1986 (N_1986,N_324,N_949);
nand U1987 (N_1987,In_2701,In_2526);
or U1988 (N_1988,In_684,N_504);
and U1989 (N_1989,N_529,N_981);
or U1990 (N_1990,N_454,In_1730);
nand U1991 (N_1991,N_134,N_363);
or U1992 (N_1992,N_711,In_1472);
xor U1993 (N_1993,N_607,In_2950);
and U1994 (N_1994,N_334,N_932);
nor U1995 (N_1995,In_944,In_22);
or U1996 (N_1996,In_513,In_871);
and U1997 (N_1997,N_45,N_130);
nand U1998 (N_1998,N_970,In_2506);
xnor U1999 (N_1999,In_1202,In_1448);
nand U2000 (N_2000,N_1839,N_1065);
nor U2001 (N_2001,N_1311,N_1336);
nor U2002 (N_2002,N_1795,N_1805);
or U2003 (N_2003,N_1587,N_1716);
and U2004 (N_2004,N_1622,N_1141);
or U2005 (N_2005,N_1613,N_1176);
nor U2006 (N_2006,N_1219,N_1989);
nand U2007 (N_2007,N_1975,N_1812);
or U2008 (N_2008,N_1309,N_1786);
xnor U2009 (N_2009,N_1612,N_1059);
nor U2010 (N_2010,N_1379,N_1441);
xor U2011 (N_2011,N_1516,N_1746);
xnor U2012 (N_2012,N_1035,N_1632);
nand U2013 (N_2013,N_1569,N_1578);
and U2014 (N_2014,N_1428,N_1177);
nand U2015 (N_2015,N_1470,N_1500);
or U2016 (N_2016,N_1947,N_1251);
nor U2017 (N_2017,N_1664,N_1029);
and U2018 (N_2018,N_1913,N_1356);
nand U2019 (N_2019,N_1970,N_1170);
nor U2020 (N_2020,N_1886,N_1004);
xor U2021 (N_2021,N_1999,N_1079);
nand U2022 (N_2022,N_1486,N_1210);
or U2023 (N_2023,N_1078,N_1686);
or U2024 (N_2024,N_1061,N_1877);
nand U2025 (N_2025,N_1867,N_1100);
or U2026 (N_2026,N_1396,N_1286);
nor U2027 (N_2027,N_1070,N_1995);
nor U2028 (N_2028,N_1199,N_1451);
or U2029 (N_2029,N_1386,N_1952);
or U2030 (N_2030,N_1002,N_1926);
xnor U2031 (N_2031,N_1399,N_1920);
xnor U2032 (N_2032,N_1841,N_1382);
xnor U2033 (N_2033,N_1791,N_1136);
or U2034 (N_2034,N_1579,N_1343);
nand U2035 (N_2035,N_1284,N_1520);
or U2036 (N_2036,N_1456,N_1505);
and U2037 (N_2037,N_1387,N_1442);
and U2038 (N_2038,N_1123,N_1024);
or U2039 (N_2039,N_1719,N_1640);
xnor U2040 (N_2040,N_1459,N_1419);
and U2041 (N_2041,N_1101,N_1776);
nor U2042 (N_2042,N_1488,N_1750);
nor U2043 (N_2043,N_1190,N_1129);
nor U2044 (N_2044,N_1656,N_1014);
and U2045 (N_2045,N_1221,N_1938);
nand U2046 (N_2046,N_1810,N_1852);
nand U2047 (N_2047,N_1756,N_1925);
and U2048 (N_2048,N_1702,N_1005);
and U2049 (N_2049,N_1067,N_1015);
nand U2050 (N_2050,N_1388,N_1230);
nor U2051 (N_2051,N_1714,N_1836);
xor U2052 (N_2052,N_1769,N_1277);
nand U2053 (N_2053,N_1401,N_1196);
or U2054 (N_2054,N_1711,N_1904);
or U2055 (N_2055,N_1527,N_1993);
nand U2056 (N_2056,N_1148,N_1856);
nand U2057 (N_2057,N_1019,N_1740);
and U2058 (N_2058,N_1205,N_1742);
or U2059 (N_2059,N_1784,N_1151);
and U2060 (N_2060,N_1051,N_1003);
or U2061 (N_2061,N_1454,N_1394);
nand U2062 (N_2062,N_1780,N_1536);
nor U2063 (N_2063,N_1127,N_1305);
nand U2064 (N_2064,N_1771,N_1863);
or U2065 (N_2065,N_1820,N_1627);
xor U2066 (N_2066,N_1888,N_1996);
nand U2067 (N_2067,N_1346,N_1942);
and U2068 (N_2068,N_1404,N_1586);
nand U2069 (N_2069,N_1165,N_1572);
or U2070 (N_2070,N_1918,N_1905);
or U2071 (N_2071,N_1435,N_1432);
nor U2072 (N_2072,N_1935,N_1361);
or U2073 (N_2073,N_1808,N_1338);
nor U2074 (N_2074,N_1718,N_1114);
nor U2075 (N_2075,N_1589,N_1036);
xor U2076 (N_2076,N_1874,N_1258);
xnor U2077 (N_2077,N_1255,N_1526);
nand U2078 (N_2078,N_1312,N_1501);
xnor U2079 (N_2079,N_1697,N_1759);
and U2080 (N_2080,N_1477,N_1460);
nor U2081 (N_2081,N_1507,N_1200);
nor U2082 (N_2082,N_1595,N_1720);
nand U2083 (N_2083,N_1417,N_1032);
xnor U2084 (N_2084,N_1917,N_1717);
and U2085 (N_2085,N_1696,N_1424);
and U2086 (N_2086,N_1704,N_1861);
and U2087 (N_2087,N_1760,N_1733);
or U2088 (N_2088,N_1297,N_1462);
xor U2089 (N_2089,N_1261,N_1037);
nand U2090 (N_2090,N_1367,N_1551);
and U2091 (N_2091,N_1583,N_1809);
and U2092 (N_2092,N_1541,N_1027);
xor U2093 (N_2093,N_1273,N_1131);
nand U2094 (N_2094,N_1490,N_1758);
nand U2095 (N_2095,N_1951,N_1453);
or U2096 (N_2096,N_1646,N_1076);
nor U2097 (N_2097,N_1880,N_1414);
nand U2098 (N_2098,N_1152,N_1864);
nand U2099 (N_2099,N_1039,N_1371);
and U2100 (N_2100,N_1434,N_1408);
or U2101 (N_2101,N_1638,N_1814);
nand U2102 (N_2102,N_1103,N_1008);
nor U2103 (N_2103,N_1498,N_1629);
and U2104 (N_2104,N_1548,N_1609);
or U2105 (N_2105,N_1539,N_1155);
xor U2106 (N_2106,N_1703,N_1360);
nand U2107 (N_2107,N_1057,N_1223);
nand U2108 (N_2108,N_1909,N_1535);
nor U2109 (N_2109,N_1707,N_1824);
xor U2110 (N_2110,N_1243,N_1828);
and U2111 (N_2111,N_1514,N_1392);
nor U2112 (N_2112,N_1363,N_1345);
or U2113 (N_2113,N_1184,N_1274);
nor U2114 (N_2114,N_1482,N_1294);
xor U2115 (N_2115,N_1080,N_1098);
or U2116 (N_2116,N_1436,N_1598);
and U2117 (N_2117,N_1159,N_1971);
and U2118 (N_2118,N_1095,N_1049);
nand U2119 (N_2119,N_1359,N_1953);
nor U2120 (N_2120,N_1492,N_1458);
nand U2121 (N_2121,N_1654,N_1902);
nor U2122 (N_2122,N_1307,N_1940);
and U2123 (N_2123,N_1932,N_1257);
and U2124 (N_2124,N_1204,N_1739);
xnor U2125 (N_2125,N_1285,N_1532);
nor U2126 (N_2126,N_1236,N_1988);
nand U2127 (N_2127,N_1172,N_1213);
and U2128 (N_2128,N_1806,N_1400);
nor U2129 (N_2129,N_1254,N_1679);
nor U2130 (N_2130,N_1556,N_1180);
nor U2131 (N_2131,N_1594,N_1317);
and U2132 (N_2132,N_1683,N_1021);
nor U2133 (N_2133,N_1497,N_1570);
nor U2134 (N_2134,N_1960,N_1997);
or U2135 (N_2135,N_1897,N_1416);
nand U2136 (N_2136,N_1026,N_1238);
or U2137 (N_2137,N_1876,N_1044);
or U2138 (N_2138,N_1410,N_1557);
nand U2139 (N_2139,N_1135,N_1233);
nand U2140 (N_2140,N_1693,N_1573);
xor U2141 (N_2141,N_1253,N_1647);
and U2142 (N_2142,N_1891,N_1964);
and U2143 (N_2143,N_1418,N_1147);
nor U2144 (N_2144,N_1171,N_1485);
or U2145 (N_2145,N_1673,N_1590);
xnor U2146 (N_2146,N_1502,N_1724);
xnor U2147 (N_2147,N_1833,N_1503);
nand U2148 (N_2148,N_1803,N_1741);
or U2149 (N_2149,N_1735,N_1216);
and U2150 (N_2150,N_1464,N_1921);
and U2151 (N_2151,N_1549,N_1798);
nor U2152 (N_2152,N_1788,N_1006);
or U2153 (N_2153,N_1766,N_1232);
xor U2154 (N_2154,N_1937,N_1468);
or U2155 (N_2155,N_1529,N_1827);
or U2156 (N_2156,N_1929,N_1375);
xnor U2157 (N_2157,N_1054,N_1674);
xnor U2158 (N_2158,N_1380,N_1553);
or U2159 (N_2159,N_1649,N_1042);
or U2160 (N_2160,N_1366,N_1473);
xnor U2161 (N_2161,N_1045,N_1685);
nor U2162 (N_2162,N_1241,N_1510);
nor U2163 (N_2163,N_1799,N_1467);
and U2164 (N_2164,N_1242,N_1559);
and U2165 (N_2165,N_1985,N_1637);
or U2166 (N_2166,N_1934,N_1466);
and U2167 (N_2167,N_1099,N_1007);
nor U2168 (N_2168,N_1245,N_1757);
and U2169 (N_2169,N_1561,N_1506);
nor U2170 (N_2170,N_1156,N_1455);
nor U2171 (N_2171,N_1580,N_1504);
nor U2172 (N_2172,N_1882,N_1825);
nand U2173 (N_2173,N_1819,N_1624);
nor U2174 (N_2174,N_1593,N_1672);
xnor U2175 (N_2175,N_1600,N_1818);
and U2176 (N_2176,N_1635,N_1228);
xnor U2177 (N_2177,N_1496,N_1318);
or U2178 (N_2178,N_1671,N_1144);
nand U2179 (N_2179,N_1302,N_1053);
and U2180 (N_2180,N_1816,N_1499);
nand U2181 (N_2181,N_1206,N_1090);
or U2182 (N_2182,N_1352,N_1083);
nor U2183 (N_2183,N_1472,N_1900);
or U2184 (N_2184,N_1325,N_1128);
or U2185 (N_2185,N_1108,N_1109);
nor U2186 (N_2186,N_1288,N_1519);
or U2187 (N_2187,N_1916,N_1730);
nor U2188 (N_2188,N_1287,N_1217);
and U2189 (N_2189,N_1813,N_1789);
xor U2190 (N_2190,N_1142,N_1614);
or U2191 (N_2191,N_1430,N_1933);
and U2192 (N_2192,N_1310,N_1092);
xor U2193 (N_2193,N_1064,N_1249);
xor U2194 (N_2194,N_1817,N_1113);
and U2195 (N_2195,N_1826,N_1163);
nand U2196 (N_2196,N_1901,N_1525);
nand U2197 (N_2197,N_1745,N_1331);
or U2198 (N_2198,N_1038,N_1182);
nand U2199 (N_2199,N_1203,N_1438);
nor U2200 (N_2200,N_1087,N_1889);
xnor U2201 (N_2201,N_1787,N_1568);
or U2202 (N_2202,N_1322,N_1211);
nand U2203 (N_2203,N_1981,N_1262);
and U2204 (N_2204,N_1321,N_1815);
or U2205 (N_2205,N_1732,N_1048);
nand U2206 (N_2206,N_1606,N_1752);
or U2207 (N_2207,N_1911,N_1487);
nor U2208 (N_2208,N_1120,N_1617);
nand U2209 (N_2209,N_1393,N_1692);
and U2210 (N_2210,N_1489,N_1009);
nor U2211 (N_2211,N_1362,N_1154);
nand U2212 (N_2212,N_1316,N_1774);
or U2213 (N_2213,N_1948,N_1138);
xor U2214 (N_2214,N_1370,N_1025);
nand U2215 (N_2215,N_1452,N_1611);
and U2216 (N_2216,N_1373,N_1481);
or U2217 (N_2217,N_1413,N_1461);
xnor U2218 (N_2218,N_1189,N_1094);
nor U2219 (N_2219,N_1082,N_1843);
nand U2220 (N_2220,N_1246,N_1722);
nor U2221 (N_2221,N_1091,N_1829);
and U2222 (N_2222,N_1765,N_1073);
and U2223 (N_2223,N_1097,N_1280);
or U2224 (N_2224,N_1052,N_1945);
nand U2225 (N_2225,N_1830,N_1565);
xnor U2226 (N_2226,N_1515,N_1562);
and U2227 (N_2227,N_1773,N_1471);
and U2228 (N_2228,N_1391,N_1599);
nand U2229 (N_2229,N_1275,N_1639);
or U2230 (N_2230,N_1610,N_1222);
nand U2231 (N_2231,N_1224,N_1320);
nor U2232 (N_2232,N_1353,N_1378);
or U2233 (N_2233,N_1174,N_1162);
xnor U2234 (N_2234,N_1838,N_1134);
nand U2235 (N_2235,N_1081,N_1476);
xor U2236 (N_2236,N_1961,N_1050);
and U2237 (N_2237,N_1256,N_1000);
or U2238 (N_2238,N_1326,N_1509);
nor U2239 (N_2239,N_1969,N_1235);
or U2240 (N_2240,N_1706,N_1063);
xnor U2241 (N_2241,N_1749,N_1423);
or U2242 (N_2242,N_1854,N_1870);
nor U2243 (N_2243,N_1688,N_1849);
or U2244 (N_2244,N_1445,N_1066);
and U2245 (N_2245,N_1178,N_1409);
nor U2246 (N_2246,N_1463,N_1859);
nand U2247 (N_2247,N_1075,N_1865);
xnor U2248 (N_2248,N_1289,N_1313);
nor U2249 (N_2249,N_1832,N_1104);
xnor U2250 (N_2250,N_1479,N_1293);
and U2251 (N_2251,N_1700,N_1149);
nand U2252 (N_2252,N_1919,N_1282);
xor U2253 (N_2253,N_1678,N_1851);
nand U2254 (N_2254,N_1234,N_1040);
and U2255 (N_2255,N_1543,N_1102);
or U2256 (N_2256,N_1350,N_1111);
nand U2257 (N_2257,N_1552,N_1212);
nand U2258 (N_2258,N_1755,N_1764);
and U2259 (N_2259,N_1140,N_1955);
xor U2260 (N_2260,N_1978,N_1582);
xor U2261 (N_2261,N_1695,N_1793);
nor U2262 (N_2262,N_1980,N_1449);
nor U2263 (N_2263,N_1831,N_1124);
or U2264 (N_2264,N_1577,N_1112);
nor U2265 (N_2265,N_1121,N_1540);
or U2266 (N_2266,N_1106,N_1547);
nand U2267 (N_2267,N_1374,N_1967);
nand U2268 (N_2268,N_1943,N_1016);
nand U2269 (N_2269,N_1385,N_1270);
nand U2270 (N_2270,N_1469,N_1575);
or U2271 (N_2271,N_1010,N_1558);
and U2272 (N_2272,N_1324,N_1429);
nand U2273 (N_2273,N_1823,N_1291);
nor U2274 (N_2274,N_1797,N_1369);
and U2275 (N_2275,N_1898,N_1875);
nand U2276 (N_2276,N_1554,N_1560);
and U2277 (N_2277,N_1710,N_1443);
or U2278 (N_2278,N_1998,N_1011);
nand U2279 (N_2279,N_1615,N_1368);
or U2280 (N_2280,N_1330,N_1041);
nor U2281 (N_2281,N_1296,N_1872);
xor U2282 (N_2282,N_1768,N_1146);
and U2283 (N_2283,N_1517,N_1986);
nand U2284 (N_2284,N_1907,N_1398);
and U2285 (N_2285,N_1857,N_1652);
xor U2286 (N_2286,N_1604,N_1523);
and U2287 (N_2287,N_1744,N_1936);
nand U2288 (N_2288,N_1644,N_1893);
nor U2289 (N_2289,N_1194,N_1976);
nand U2290 (N_2290,N_1290,N_1915);
or U2291 (N_2291,N_1491,N_1628);
nand U2292 (N_2292,N_1869,N_1181);
or U2293 (N_2293,N_1546,N_1957);
nor U2294 (N_2294,N_1252,N_1655);
nand U2295 (N_2295,N_1892,N_1340);
and U2296 (N_2296,N_1800,N_1166);
nor U2297 (N_2297,N_1439,N_1950);
xor U2298 (N_2298,N_1447,N_1896);
xor U2299 (N_2299,N_1173,N_1093);
and U2300 (N_2300,N_1618,N_1748);
xor U2301 (N_2301,N_1626,N_1761);
and U2302 (N_2302,N_1145,N_1130);
and U2303 (N_2303,N_1348,N_1690);
xor U2304 (N_2304,N_1364,N_1954);
or U2305 (N_2305,N_1792,N_1931);
xor U2306 (N_2306,N_1751,N_1979);
xnor U2307 (N_2307,N_1992,N_1962);
or U2308 (N_2308,N_1132,N_1747);
nor U2309 (N_2309,N_1862,N_1659);
and U2310 (N_2310,N_1840,N_1033);
nor U2311 (N_2311,N_1648,N_1427);
nand U2312 (N_2312,N_1191,N_1924);
xor U2313 (N_2313,N_1705,N_1390);
xor U2314 (N_2314,N_1956,N_1342);
nor U2315 (N_2315,N_1636,N_1666);
xnor U2316 (N_2316,N_1337,N_1781);
xor U2317 (N_2317,N_1267,N_1984);
nor U2318 (N_2318,N_1737,N_1495);
or U2319 (N_2319,N_1023,N_1949);
xor U2320 (N_2320,N_1143,N_1247);
nor U2321 (N_2321,N_1801,N_1185);
and U2322 (N_2322,N_1259,N_1665);
or U2323 (N_2323,N_1887,N_1349);
nand U2324 (N_2324,N_1058,N_1680);
or U2325 (N_2325,N_1726,N_1405);
nand U2326 (N_2326,N_1314,N_1698);
and U2327 (N_2327,N_1794,N_1890);
xor U2328 (N_2328,N_1069,N_1167);
and U2329 (N_2329,N_1281,N_1608);
nor U2330 (N_2330,N_1446,N_1738);
or U2331 (N_2331,N_1597,N_1778);
xnor U2332 (N_2332,N_1264,N_1512);
or U2333 (N_2333,N_1115,N_1433);
nand U2334 (N_2334,N_1939,N_1117);
nand U2335 (N_2335,N_1567,N_1734);
or U2336 (N_2336,N_1621,N_1725);
or U2337 (N_2337,N_1301,N_1581);
and U2338 (N_2338,N_1871,N_1753);
nand U2339 (N_2339,N_1202,N_1511);
nand U2340 (N_2340,N_1796,N_1187);
and U2341 (N_2341,N_1422,N_1974);
nand U2342 (N_2342,N_1043,N_1475);
and U2343 (N_2343,N_1645,N_1347);
xor U2344 (N_2344,N_1855,N_1474);
and U2345 (N_2345,N_1848,N_1545);
nor U2346 (N_2346,N_1585,N_1723);
nand U2347 (N_2347,N_1183,N_1912);
xor U2348 (N_2348,N_1958,N_1304);
or U2349 (N_2349,N_1341,N_1837);
xor U2350 (N_2350,N_1965,N_1675);
nand U2351 (N_2351,N_1767,N_1195);
or U2352 (N_2352,N_1633,N_1372);
or U2353 (N_2353,N_1885,N_1770);
or U2354 (N_2354,N_1110,N_1508);
or U2355 (N_2355,N_1643,N_1625);
or U2356 (N_2356,N_1339,N_1186);
xnor U2357 (N_2357,N_1743,N_1225);
xnor U2358 (N_2358,N_1914,N_1670);
nand U2359 (N_2359,N_1244,N_1315);
xor U2360 (N_2360,N_1480,N_1853);
and U2361 (N_2361,N_1332,N_1908);
and U2362 (N_2362,N_1013,N_1085);
nand U2363 (N_2363,N_1990,N_1521);
nor U2364 (N_2364,N_1240,N_1616);
nor U2365 (N_2365,N_1335,N_1762);
or U2366 (N_2366,N_1959,N_1383);
nand U2367 (N_2367,N_1518,N_1484);
xor U2368 (N_2368,N_1207,N_1208);
xnor U2369 (N_2369,N_1982,N_1906);
xnor U2370 (N_2370,N_1607,N_1513);
or U2371 (N_2371,N_1116,N_1728);
and U2372 (N_2372,N_1620,N_1214);
or U2373 (N_2373,N_1358,N_1158);
or U2374 (N_2374,N_1689,N_1963);
or U2375 (N_2375,N_1197,N_1031);
nor U2376 (N_2376,N_1701,N_1237);
and U2377 (N_2377,N_1164,N_1623);
xor U2378 (N_2378,N_1930,N_1444);
xor U2379 (N_2379,N_1537,N_1550);
and U2380 (N_2380,N_1239,N_1847);
and U2381 (N_2381,N_1105,N_1642);
nor U2382 (N_2382,N_1403,N_1415);
and U2383 (N_2383,N_1844,N_1528);
xnor U2384 (N_2384,N_1055,N_1641);
nor U2385 (N_2385,N_1420,N_1248);
or U2386 (N_2386,N_1785,N_1062);
or U2387 (N_2387,N_1278,N_1431);
nor U2388 (N_2388,N_1283,N_1653);
xnor U2389 (N_2389,N_1250,N_1319);
nand U2390 (N_2390,N_1691,N_1866);
xnor U2391 (N_2391,N_1001,N_1272);
nor U2392 (N_2392,N_1899,N_1198);
and U2393 (N_2393,N_1402,N_1650);
xnor U2394 (N_2394,N_1096,N_1192);
nor U2395 (N_2395,N_1271,N_1107);
nor U2396 (N_2396,N_1669,N_1715);
or U2397 (N_2397,N_1910,N_1603);
xor U2398 (N_2398,N_1946,N_1457);
or U2399 (N_2399,N_1071,N_1161);
and U2400 (N_2400,N_1987,N_1068);
or U2401 (N_2401,N_1658,N_1821);
xnor U2402 (N_2402,N_1983,N_1088);
or U2403 (N_2403,N_1295,N_1591);
or U2404 (N_2404,N_1160,N_1299);
nor U2405 (N_2405,N_1020,N_1175);
and U2406 (N_2406,N_1133,N_1226);
and U2407 (N_2407,N_1030,N_1169);
or U2408 (N_2408,N_1602,N_1328);
or U2409 (N_2409,N_1588,N_1564);
or U2410 (N_2410,N_1811,N_1357);
nor U2411 (N_2411,N_1660,N_1308);
nor U2412 (N_2412,N_1850,N_1682);
or U2413 (N_2413,N_1651,N_1713);
and U2414 (N_2414,N_1426,N_1351);
or U2415 (N_2415,N_1150,N_1524);
nor U2416 (N_2416,N_1822,N_1736);
and U2417 (N_2417,N_1927,N_1972);
or U2418 (N_2418,N_1542,N_1721);
xnor U2419 (N_2419,N_1994,N_1894);
xor U2420 (N_2420,N_1437,N_1531);
or U2421 (N_2421,N_1306,N_1699);
or U2422 (N_2422,N_1072,N_1846);
and U2423 (N_2423,N_1584,N_1193);
xor U2424 (N_2424,N_1574,N_1712);
xnor U2425 (N_2425,N_1266,N_1268);
and U2426 (N_2426,N_1941,N_1333);
xor U2427 (N_2427,N_1046,N_1534);
nand U2428 (N_2428,N_1977,N_1630);
nor U2429 (N_2429,N_1881,N_1265);
nor U2430 (N_2430,N_1478,N_1137);
xor U2431 (N_2431,N_1018,N_1968);
nor U2432 (N_2432,N_1086,N_1125);
nand U2433 (N_2433,N_1168,N_1201);
nand U2434 (N_2434,N_1571,N_1074);
nand U2435 (N_2435,N_1619,N_1601);
nor U2436 (N_2436,N_1754,N_1779);
or U2437 (N_2437,N_1835,N_1406);
nand U2438 (N_2438,N_1209,N_1298);
nor U2439 (N_2439,N_1012,N_1119);
nand U2440 (N_2440,N_1056,N_1303);
or U2441 (N_2441,N_1631,N_1522);
or U2442 (N_2442,N_1260,N_1538);
or U2443 (N_2443,N_1300,N_1220);
or U2444 (N_2444,N_1448,N_1729);
xor U2445 (N_2445,N_1483,N_1231);
nand U2446 (N_2446,N_1411,N_1028);
or U2447 (N_2447,N_1804,N_1139);
and U2448 (N_2448,N_1060,N_1566);
and U2449 (N_2449,N_1218,N_1858);
nand U2450 (N_2450,N_1407,N_1022);
or U2451 (N_2451,N_1263,N_1709);
xnor U2452 (N_2452,N_1397,N_1563);
and U2453 (N_2453,N_1694,N_1395);
xnor U2454 (N_2454,N_1681,N_1802);
and U2455 (N_2455,N_1276,N_1034);
nand U2456 (N_2456,N_1334,N_1533);
nand U2457 (N_2457,N_1329,N_1188);
or U2458 (N_2458,N_1077,N_1596);
or U2459 (N_2459,N_1879,N_1344);
or U2460 (N_2460,N_1576,N_1544);
or U2461 (N_2461,N_1662,N_1772);
nor U2462 (N_2462,N_1687,N_1269);
and U2463 (N_2463,N_1667,N_1381);
nor U2464 (N_2464,N_1790,N_1425);
nand U2465 (N_2465,N_1676,N_1355);
xor U2466 (N_2466,N_1450,N_1883);
or U2467 (N_2467,N_1834,N_1279);
nor U2468 (N_2468,N_1884,N_1783);
nand U2469 (N_2469,N_1122,N_1389);
nand U2470 (N_2470,N_1047,N_1668);
xor U2471 (N_2471,N_1657,N_1663);
nand U2472 (N_2472,N_1292,N_1966);
or U2473 (N_2473,N_1991,N_1777);
or U2474 (N_2474,N_1323,N_1118);
and U2475 (N_2475,N_1089,N_1421);
xor U2476 (N_2476,N_1605,N_1084);
nand U2477 (N_2477,N_1179,N_1807);
and U2478 (N_2478,N_1493,N_1782);
nand U2479 (N_2479,N_1873,N_1860);
nand U2480 (N_2480,N_1878,N_1327);
nor U2481 (N_2481,N_1227,N_1153);
or U2482 (N_2482,N_1684,N_1842);
nor U2483 (N_2483,N_1973,N_1634);
nand U2484 (N_2484,N_1465,N_1868);
and U2485 (N_2485,N_1555,N_1763);
or U2486 (N_2486,N_1677,N_1708);
nand U2487 (N_2487,N_1215,N_1126);
or U2488 (N_2488,N_1494,N_1661);
xor U2489 (N_2489,N_1017,N_1928);
xnor U2490 (N_2490,N_1530,N_1731);
or U2491 (N_2491,N_1727,N_1903);
nand U2492 (N_2492,N_1775,N_1922);
nor U2493 (N_2493,N_1384,N_1923);
nand U2494 (N_2494,N_1376,N_1845);
xnor U2495 (N_2495,N_1157,N_1229);
xor U2496 (N_2496,N_1895,N_1440);
xnor U2497 (N_2497,N_1377,N_1944);
or U2498 (N_2498,N_1412,N_1592);
nand U2499 (N_2499,N_1354,N_1365);
or U2500 (N_2500,N_1222,N_1622);
and U2501 (N_2501,N_1889,N_1707);
xor U2502 (N_2502,N_1591,N_1251);
nand U2503 (N_2503,N_1413,N_1224);
or U2504 (N_2504,N_1375,N_1463);
nand U2505 (N_2505,N_1860,N_1991);
nor U2506 (N_2506,N_1046,N_1177);
xor U2507 (N_2507,N_1266,N_1251);
nand U2508 (N_2508,N_1228,N_1568);
or U2509 (N_2509,N_1006,N_1883);
nand U2510 (N_2510,N_1435,N_1018);
nand U2511 (N_2511,N_1675,N_1497);
xnor U2512 (N_2512,N_1612,N_1715);
xor U2513 (N_2513,N_1494,N_1397);
or U2514 (N_2514,N_1193,N_1685);
xor U2515 (N_2515,N_1863,N_1772);
or U2516 (N_2516,N_1771,N_1557);
xnor U2517 (N_2517,N_1303,N_1114);
xor U2518 (N_2518,N_1516,N_1709);
or U2519 (N_2519,N_1067,N_1874);
nand U2520 (N_2520,N_1405,N_1880);
xnor U2521 (N_2521,N_1132,N_1457);
nand U2522 (N_2522,N_1744,N_1910);
nand U2523 (N_2523,N_1438,N_1962);
nand U2524 (N_2524,N_1976,N_1764);
xor U2525 (N_2525,N_1837,N_1541);
xor U2526 (N_2526,N_1687,N_1416);
nand U2527 (N_2527,N_1673,N_1707);
nor U2528 (N_2528,N_1666,N_1152);
xnor U2529 (N_2529,N_1529,N_1626);
nand U2530 (N_2530,N_1668,N_1486);
or U2531 (N_2531,N_1034,N_1872);
and U2532 (N_2532,N_1330,N_1752);
xor U2533 (N_2533,N_1011,N_1751);
nor U2534 (N_2534,N_1768,N_1318);
or U2535 (N_2535,N_1259,N_1358);
xor U2536 (N_2536,N_1694,N_1065);
nor U2537 (N_2537,N_1103,N_1078);
or U2538 (N_2538,N_1032,N_1921);
nor U2539 (N_2539,N_1853,N_1800);
and U2540 (N_2540,N_1377,N_1343);
or U2541 (N_2541,N_1265,N_1901);
xnor U2542 (N_2542,N_1760,N_1884);
xor U2543 (N_2543,N_1304,N_1378);
or U2544 (N_2544,N_1802,N_1387);
and U2545 (N_2545,N_1337,N_1514);
or U2546 (N_2546,N_1080,N_1116);
and U2547 (N_2547,N_1900,N_1353);
nor U2548 (N_2548,N_1063,N_1604);
or U2549 (N_2549,N_1811,N_1866);
xnor U2550 (N_2550,N_1051,N_1976);
nor U2551 (N_2551,N_1590,N_1923);
and U2552 (N_2552,N_1316,N_1695);
nor U2553 (N_2553,N_1396,N_1753);
xnor U2554 (N_2554,N_1370,N_1497);
xor U2555 (N_2555,N_1415,N_1680);
nor U2556 (N_2556,N_1160,N_1685);
nand U2557 (N_2557,N_1525,N_1911);
and U2558 (N_2558,N_1604,N_1223);
and U2559 (N_2559,N_1678,N_1599);
nand U2560 (N_2560,N_1859,N_1927);
or U2561 (N_2561,N_1935,N_1068);
nand U2562 (N_2562,N_1826,N_1031);
and U2563 (N_2563,N_1134,N_1546);
and U2564 (N_2564,N_1493,N_1157);
nor U2565 (N_2565,N_1218,N_1233);
and U2566 (N_2566,N_1441,N_1568);
and U2567 (N_2567,N_1866,N_1361);
nor U2568 (N_2568,N_1933,N_1044);
or U2569 (N_2569,N_1969,N_1086);
nor U2570 (N_2570,N_1783,N_1217);
nand U2571 (N_2571,N_1758,N_1355);
or U2572 (N_2572,N_1122,N_1856);
xor U2573 (N_2573,N_1120,N_1972);
nand U2574 (N_2574,N_1323,N_1974);
nand U2575 (N_2575,N_1770,N_1166);
and U2576 (N_2576,N_1623,N_1193);
nor U2577 (N_2577,N_1514,N_1568);
or U2578 (N_2578,N_1998,N_1755);
or U2579 (N_2579,N_1923,N_1023);
nand U2580 (N_2580,N_1469,N_1198);
and U2581 (N_2581,N_1746,N_1242);
nand U2582 (N_2582,N_1320,N_1967);
nor U2583 (N_2583,N_1062,N_1121);
or U2584 (N_2584,N_1046,N_1212);
nor U2585 (N_2585,N_1671,N_1750);
xnor U2586 (N_2586,N_1661,N_1512);
nor U2587 (N_2587,N_1992,N_1195);
xnor U2588 (N_2588,N_1031,N_1347);
and U2589 (N_2589,N_1159,N_1991);
nor U2590 (N_2590,N_1362,N_1938);
or U2591 (N_2591,N_1879,N_1586);
nor U2592 (N_2592,N_1202,N_1284);
and U2593 (N_2593,N_1079,N_1036);
nand U2594 (N_2594,N_1272,N_1134);
or U2595 (N_2595,N_1127,N_1648);
xnor U2596 (N_2596,N_1548,N_1021);
nor U2597 (N_2597,N_1700,N_1738);
nor U2598 (N_2598,N_1575,N_1537);
nand U2599 (N_2599,N_1994,N_1927);
nand U2600 (N_2600,N_1251,N_1196);
nor U2601 (N_2601,N_1577,N_1862);
nor U2602 (N_2602,N_1233,N_1056);
nand U2603 (N_2603,N_1098,N_1459);
nand U2604 (N_2604,N_1901,N_1848);
xnor U2605 (N_2605,N_1498,N_1866);
xor U2606 (N_2606,N_1965,N_1054);
and U2607 (N_2607,N_1903,N_1541);
and U2608 (N_2608,N_1156,N_1853);
or U2609 (N_2609,N_1386,N_1046);
nor U2610 (N_2610,N_1420,N_1593);
xnor U2611 (N_2611,N_1618,N_1373);
or U2612 (N_2612,N_1506,N_1592);
xor U2613 (N_2613,N_1214,N_1682);
and U2614 (N_2614,N_1931,N_1892);
or U2615 (N_2615,N_1913,N_1570);
nand U2616 (N_2616,N_1061,N_1576);
xor U2617 (N_2617,N_1484,N_1052);
nand U2618 (N_2618,N_1111,N_1442);
nand U2619 (N_2619,N_1997,N_1452);
and U2620 (N_2620,N_1934,N_1274);
xor U2621 (N_2621,N_1608,N_1624);
or U2622 (N_2622,N_1320,N_1922);
and U2623 (N_2623,N_1240,N_1196);
or U2624 (N_2624,N_1067,N_1275);
xnor U2625 (N_2625,N_1260,N_1416);
and U2626 (N_2626,N_1722,N_1557);
xor U2627 (N_2627,N_1088,N_1097);
nor U2628 (N_2628,N_1087,N_1816);
nand U2629 (N_2629,N_1335,N_1756);
or U2630 (N_2630,N_1586,N_1294);
xor U2631 (N_2631,N_1717,N_1475);
xnor U2632 (N_2632,N_1787,N_1089);
or U2633 (N_2633,N_1676,N_1273);
or U2634 (N_2634,N_1995,N_1121);
nor U2635 (N_2635,N_1771,N_1143);
and U2636 (N_2636,N_1097,N_1196);
or U2637 (N_2637,N_1650,N_1941);
or U2638 (N_2638,N_1929,N_1376);
nand U2639 (N_2639,N_1518,N_1681);
nand U2640 (N_2640,N_1079,N_1294);
and U2641 (N_2641,N_1155,N_1496);
nand U2642 (N_2642,N_1881,N_1664);
or U2643 (N_2643,N_1545,N_1485);
nor U2644 (N_2644,N_1335,N_1233);
xnor U2645 (N_2645,N_1250,N_1473);
and U2646 (N_2646,N_1451,N_1711);
and U2647 (N_2647,N_1481,N_1334);
nor U2648 (N_2648,N_1898,N_1324);
and U2649 (N_2649,N_1435,N_1867);
or U2650 (N_2650,N_1785,N_1121);
xor U2651 (N_2651,N_1660,N_1196);
xnor U2652 (N_2652,N_1956,N_1004);
xnor U2653 (N_2653,N_1488,N_1132);
nand U2654 (N_2654,N_1741,N_1801);
or U2655 (N_2655,N_1791,N_1165);
xnor U2656 (N_2656,N_1254,N_1204);
nand U2657 (N_2657,N_1596,N_1415);
nor U2658 (N_2658,N_1606,N_1632);
and U2659 (N_2659,N_1815,N_1849);
nand U2660 (N_2660,N_1175,N_1388);
xnor U2661 (N_2661,N_1852,N_1539);
and U2662 (N_2662,N_1870,N_1754);
or U2663 (N_2663,N_1575,N_1806);
nor U2664 (N_2664,N_1463,N_1473);
and U2665 (N_2665,N_1125,N_1664);
or U2666 (N_2666,N_1782,N_1375);
or U2667 (N_2667,N_1190,N_1654);
and U2668 (N_2668,N_1342,N_1580);
xnor U2669 (N_2669,N_1366,N_1809);
xor U2670 (N_2670,N_1300,N_1435);
nor U2671 (N_2671,N_1202,N_1804);
nor U2672 (N_2672,N_1366,N_1763);
or U2673 (N_2673,N_1654,N_1266);
nand U2674 (N_2674,N_1733,N_1534);
and U2675 (N_2675,N_1479,N_1366);
or U2676 (N_2676,N_1264,N_1711);
or U2677 (N_2677,N_1107,N_1560);
or U2678 (N_2678,N_1236,N_1390);
and U2679 (N_2679,N_1838,N_1884);
or U2680 (N_2680,N_1451,N_1293);
and U2681 (N_2681,N_1023,N_1873);
and U2682 (N_2682,N_1561,N_1527);
and U2683 (N_2683,N_1080,N_1871);
and U2684 (N_2684,N_1914,N_1716);
and U2685 (N_2685,N_1936,N_1251);
or U2686 (N_2686,N_1640,N_1015);
xor U2687 (N_2687,N_1136,N_1679);
and U2688 (N_2688,N_1335,N_1354);
nor U2689 (N_2689,N_1120,N_1246);
or U2690 (N_2690,N_1579,N_1959);
xnor U2691 (N_2691,N_1403,N_1855);
xor U2692 (N_2692,N_1865,N_1499);
nor U2693 (N_2693,N_1299,N_1966);
nand U2694 (N_2694,N_1282,N_1222);
nor U2695 (N_2695,N_1112,N_1325);
nand U2696 (N_2696,N_1322,N_1194);
nand U2697 (N_2697,N_1591,N_1819);
or U2698 (N_2698,N_1282,N_1414);
and U2699 (N_2699,N_1413,N_1531);
or U2700 (N_2700,N_1566,N_1891);
and U2701 (N_2701,N_1085,N_1702);
nor U2702 (N_2702,N_1657,N_1388);
xor U2703 (N_2703,N_1751,N_1511);
and U2704 (N_2704,N_1285,N_1638);
or U2705 (N_2705,N_1739,N_1707);
or U2706 (N_2706,N_1763,N_1966);
nor U2707 (N_2707,N_1935,N_1011);
xnor U2708 (N_2708,N_1741,N_1330);
nor U2709 (N_2709,N_1746,N_1014);
nand U2710 (N_2710,N_1533,N_1344);
xor U2711 (N_2711,N_1690,N_1142);
or U2712 (N_2712,N_1463,N_1136);
nor U2713 (N_2713,N_1542,N_1900);
nor U2714 (N_2714,N_1796,N_1275);
xor U2715 (N_2715,N_1387,N_1361);
nor U2716 (N_2716,N_1981,N_1880);
nand U2717 (N_2717,N_1980,N_1651);
or U2718 (N_2718,N_1356,N_1974);
or U2719 (N_2719,N_1675,N_1827);
nand U2720 (N_2720,N_1387,N_1001);
or U2721 (N_2721,N_1586,N_1630);
xnor U2722 (N_2722,N_1128,N_1359);
nand U2723 (N_2723,N_1233,N_1536);
or U2724 (N_2724,N_1589,N_1040);
xnor U2725 (N_2725,N_1685,N_1761);
or U2726 (N_2726,N_1138,N_1406);
xnor U2727 (N_2727,N_1121,N_1624);
nand U2728 (N_2728,N_1303,N_1907);
xor U2729 (N_2729,N_1316,N_1159);
or U2730 (N_2730,N_1163,N_1158);
xor U2731 (N_2731,N_1588,N_1411);
or U2732 (N_2732,N_1441,N_1512);
xor U2733 (N_2733,N_1753,N_1251);
and U2734 (N_2734,N_1424,N_1215);
and U2735 (N_2735,N_1860,N_1982);
or U2736 (N_2736,N_1954,N_1488);
nor U2737 (N_2737,N_1656,N_1414);
xor U2738 (N_2738,N_1458,N_1092);
nand U2739 (N_2739,N_1594,N_1580);
xor U2740 (N_2740,N_1683,N_1467);
and U2741 (N_2741,N_1508,N_1196);
and U2742 (N_2742,N_1437,N_1371);
xor U2743 (N_2743,N_1450,N_1772);
nor U2744 (N_2744,N_1861,N_1968);
nor U2745 (N_2745,N_1104,N_1619);
and U2746 (N_2746,N_1768,N_1591);
xnor U2747 (N_2747,N_1643,N_1658);
or U2748 (N_2748,N_1094,N_1907);
nand U2749 (N_2749,N_1517,N_1178);
xor U2750 (N_2750,N_1181,N_1378);
nand U2751 (N_2751,N_1941,N_1889);
xor U2752 (N_2752,N_1335,N_1246);
nand U2753 (N_2753,N_1954,N_1403);
nor U2754 (N_2754,N_1041,N_1335);
nor U2755 (N_2755,N_1129,N_1755);
and U2756 (N_2756,N_1121,N_1469);
nand U2757 (N_2757,N_1927,N_1546);
and U2758 (N_2758,N_1266,N_1713);
and U2759 (N_2759,N_1412,N_1429);
nand U2760 (N_2760,N_1669,N_1995);
xor U2761 (N_2761,N_1944,N_1848);
and U2762 (N_2762,N_1111,N_1130);
xor U2763 (N_2763,N_1030,N_1097);
xnor U2764 (N_2764,N_1014,N_1264);
xnor U2765 (N_2765,N_1312,N_1040);
nor U2766 (N_2766,N_1241,N_1629);
nor U2767 (N_2767,N_1970,N_1172);
xor U2768 (N_2768,N_1256,N_1248);
and U2769 (N_2769,N_1216,N_1151);
xor U2770 (N_2770,N_1600,N_1112);
and U2771 (N_2771,N_1267,N_1974);
and U2772 (N_2772,N_1317,N_1905);
nand U2773 (N_2773,N_1714,N_1683);
xnor U2774 (N_2774,N_1746,N_1072);
or U2775 (N_2775,N_1850,N_1597);
xnor U2776 (N_2776,N_1452,N_1851);
or U2777 (N_2777,N_1925,N_1573);
or U2778 (N_2778,N_1884,N_1038);
nor U2779 (N_2779,N_1725,N_1999);
nand U2780 (N_2780,N_1619,N_1346);
or U2781 (N_2781,N_1365,N_1289);
or U2782 (N_2782,N_1182,N_1758);
or U2783 (N_2783,N_1012,N_1738);
nor U2784 (N_2784,N_1739,N_1915);
nand U2785 (N_2785,N_1786,N_1840);
and U2786 (N_2786,N_1688,N_1262);
and U2787 (N_2787,N_1527,N_1758);
and U2788 (N_2788,N_1880,N_1863);
or U2789 (N_2789,N_1582,N_1004);
or U2790 (N_2790,N_1341,N_1397);
and U2791 (N_2791,N_1498,N_1814);
and U2792 (N_2792,N_1836,N_1205);
or U2793 (N_2793,N_1210,N_1943);
nor U2794 (N_2794,N_1344,N_1451);
and U2795 (N_2795,N_1479,N_1850);
xor U2796 (N_2796,N_1651,N_1734);
and U2797 (N_2797,N_1680,N_1963);
nor U2798 (N_2798,N_1805,N_1672);
nor U2799 (N_2799,N_1109,N_1716);
and U2800 (N_2800,N_1465,N_1044);
or U2801 (N_2801,N_1700,N_1395);
and U2802 (N_2802,N_1162,N_1149);
xor U2803 (N_2803,N_1380,N_1376);
xor U2804 (N_2804,N_1575,N_1542);
and U2805 (N_2805,N_1533,N_1649);
or U2806 (N_2806,N_1622,N_1050);
and U2807 (N_2807,N_1943,N_1581);
nor U2808 (N_2808,N_1149,N_1869);
and U2809 (N_2809,N_1193,N_1315);
nand U2810 (N_2810,N_1222,N_1511);
nor U2811 (N_2811,N_1102,N_1288);
nor U2812 (N_2812,N_1816,N_1971);
xor U2813 (N_2813,N_1528,N_1177);
xnor U2814 (N_2814,N_1247,N_1715);
or U2815 (N_2815,N_1136,N_1586);
nor U2816 (N_2816,N_1156,N_1253);
nand U2817 (N_2817,N_1520,N_1233);
nand U2818 (N_2818,N_1946,N_1458);
nand U2819 (N_2819,N_1119,N_1798);
and U2820 (N_2820,N_1523,N_1995);
nor U2821 (N_2821,N_1778,N_1492);
nor U2822 (N_2822,N_1297,N_1399);
xor U2823 (N_2823,N_1854,N_1849);
or U2824 (N_2824,N_1945,N_1426);
xnor U2825 (N_2825,N_1710,N_1321);
xor U2826 (N_2826,N_1691,N_1886);
xor U2827 (N_2827,N_1963,N_1429);
and U2828 (N_2828,N_1685,N_1974);
or U2829 (N_2829,N_1813,N_1282);
or U2830 (N_2830,N_1531,N_1872);
nor U2831 (N_2831,N_1241,N_1236);
nand U2832 (N_2832,N_1458,N_1213);
nor U2833 (N_2833,N_1769,N_1944);
and U2834 (N_2834,N_1557,N_1889);
xor U2835 (N_2835,N_1864,N_1766);
nor U2836 (N_2836,N_1512,N_1031);
or U2837 (N_2837,N_1498,N_1436);
and U2838 (N_2838,N_1526,N_1187);
or U2839 (N_2839,N_1948,N_1624);
or U2840 (N_2840,N_1335,N_1901);
nor U2841 (N_2841,N_1693,N_1700);
nor U2842 (N_2842,N_1684,N_1202);
or U2843 (N_2843,N_1332,N_1975);
or U2844 (N_2844,N_1548,N_1979);
xnor U2845 (N_2845,N_1057,N_1102);
xor U2846 (N_2846,N_1175,N_1450);
or U2847 (N_2847,N_1027,N_1551);
nand U2848 (N_2848,N_1748,N_1369);
or U2849 (N_2849,N_1373,N_1076);
xor U2850 (N_2850,N_1476,N_1030);
and U2851 (N_2851,N_1526,N_1892);
xor U2852 (N_2852,N_1702,N_1111);
and U2853 (N_2853,N_1023,N_1679);
nand U2854 (N_2854,N_1436,N_1460);
nor U2855 (N_2855,N_1782,N_1759);
or U2856 (N_2856,N_1784,N_1870);
nor U2857 (N_2857,N_1712,N_1344);
nand U2858 (N_2858,N_1264,N_1723);
nand U2859 (N_2859,N_1883,N_1837);
nor U2860 (N_2860,N_1300,N_1655);
nand U2861 (N_2861,N_1605,N_1394);
nor U2862 (N_2862,N_1248,N_1022);
nand U2863 (N_2863,N_1691,N_1228);
or U2864 (N_2864,N_1139,N_1827);
or U2865 (N_2865,N_1081,N_1757);
nand U2866 (N_2866,N_1752,N_1074);
nor U2867 (N_2867,N_1132,N_1418);
nor U2868 (N_2868,N_1997,N_1579);
or U2869 (N_2869,N_1977,N_1102);
or U2870 (N_2870,N_1093,N_1374);
and U2871 (N_2871,N_1970,N_1738);
nor U2872 (N_2872,N_1640,N_1676);
nor U2873 (N_2873,N_1183,N_1645);
nand U2874 (N_2874,N_1629,N_1858);
nor U2875 (N_2875,N_1476,N_1229);
or U2876 (N_2876,N_1925,N_1901);
nand U2877 (N_2877,N_1137,N_1147);
and U2878 (N_2878,N_1180,N_1942);
or U2879 (N_2879,N_1992,N_1196);
xor U2880 (N_2880,N_1374,N_1527);
or U2881 (N_2881,N_1646,N_1998);
xnor U2882 (N_2882,N_1047,N_1874);
nand U2883 (N_2883,N_1688,N_1188);
and U2884 (N_2884,N_1291,N_1442);
xnor U2885 (N_2885,N_1864,N_1792);
or U2886 (N_2886,N_1652,N_1581);
nor U2887 (N_2887,N_1648,N_1036);
xnor U2888 (N_2888,N_1584,N_1210);
and U2889 (N_2889,N_1608,N_1517);
and U2890 (N_2890,N_1779,N_1125);
nand U2891 (N_2891,N_1551,N_1758);
nand U2892 (N_2892,N_1285,N_1526);
and U2893 (N_2893,N_1227,N_1501);
xnor U2894 (N_2894,N_1711,N_1515);
and U2895 (N_2895,N_1640,N_1633);
nand U2896 (N_2896,N_1183,N_1145);
nor U2897 (N_2897,N_1888,N_1167);
xor U2898 (N_2898,N_1445,N_1805);
nand U2899 (N_2899,N_1207,N_1747);
or U2900 (N_2900,N_1691,N_1403);
nor U2901 (N_2901,N_1899,N_1982);
nand U2902 (N_2902,N_1875,N_1100);
xor U2903 (N_2903,N_1041,N_1879);
or U2904 (N_2904,N_1678,N_1476);
or U2905 (N_2905,N_1678,N_1264);
xnor U2906 (N_2906,N_1664,N_1180);
xnor U2907 (N_2907,N_1297,N_1621);
nor U2908 (N_2908,N_1485,N_1219);
xnor U2909 (N_2909,N_1077,N_1452);
nand U2910 (N_2910,N_1896,N_1779);
or U2911 (N_2911,N_1214,N_1506);
or U2912 (N_2912,N_1592,N_1660);
nand U2913 (N_2913,N_1596,N_1238);
or U2914 (N_2914,N_1309,N_1398);
or U2915 (N_2915,N_1833,N_1791);
nand U2916 (N_2916,N_1430,N_1639);
or U2917 (N_2917,N_1985,N_1214);
nand U2918 (N_2918,N_1421,N_1250);
nand U2919 (N_2919,N_1997,N_1896);
and U2920 (N_2920,N_1939,N_1967);
or U2921 (N_2921,N_1989,N_1373);
xor U2922 (N_2922,N_1504,N_1333);
xnor U2923 (N_2923,N_1944,N_1694);
xor U2924 (N_2924,N_1976,N_1787);
and U2925 (N_2925,N_1491,N_1926);
or U2926 (N_2926,N_1707,N_1477);
xnor U2927 (N_2927,N_1149,N_1647);
nand U2928 (N_2928,N_1420,N_1678);
nand U2929 (N_2929,N_1855,N_1779);
and U2930 (N_2930,N_1132,N_1361);
nand U2931 (N_2931,N_1658,N_1583);
and U2932 (N_2932,N_1924,N_1040);
and U2933 (N_2933,N_1302,N_1034);
nand U2934 (N_2934,N_1276,N_1988);
nor U2935 (N_2935,N_1285,N_1659);
xor U2936 (N_2936,N_1135,N_1002);
nor U2937 (N_2937,N_1774,N_1673);
and U2938 (N_2938,N_1877,N_1164);
nor U2939 (N_2939,N_1786,N_1172);
nor U2940 (N_2940,N_1977,N_1200);
nand U2941 (N_2941,N_1119,N_1980);
nand U2942 (N_2942,N_1637,N_1946);
xor U2943 (N_2943,N_1287,N_1500);
or U2944 (N_2944,N_1645,N_1257);
and U2945 (N_2945,N_1956,N_1926);
nand U2946 (N_2946,N_1269,N_1584);
nor U2947 (N_2947,N_1783,N_1985);
xor U2948 (N_2948,N_1187,N_1229);
and U2949 (N_2949,N_1942,N_1370);
xor U2950 (N_2950,N_1483,N_1712);
and U2951 (N_2951,N_1130,N_1216);
xnor U2952 (N_2952,N_1170,N_1829);
nand U2953 (N_2953,N_1650,N_1395);
nand U2954 (N_2954,N_1762,N_1489);
and U2955 (N_2955,N_1046,N_1086);
nor U2956 (N_2956,N_1013,N_1448);
or U2957 (N_2957,N_1459,N_1630);
and U2958 (N_2958,N_1853,N_1058);
or U2959 (N_2959,N_1504,N_1778);
nor U2960 (N_2960,N_1846,N_1748);
nand U2961 (N_2961,N_1014,N_1138);
nand U2962 (N_2962,N_1508,N_1503);
nor U2963 (N_2963,N_1702,N_1584);
and U2964 (N_2964,N_1580,N_1283);
and U2965 (N_2965,N_1913,N_1797);
or U2966 (N_2966,N_1405,N_1979);
nand U2967 (N_2967,N_1523,N_1226);
and U2968 (N_2968,N_1607,N_1820);
and U2969 (N_2969,N_1869,N_1562);
or U2970 (N_2970,N_1819,N_1686);
nor U2971 (N_2971,N_1173,N_1080);
and U2972 (N_2972,N_1947,N_1620);
or U2973 (N_2973,N_1034,N_1170);
xor U2974 (N_2974,N_1698,N_1498);
nand U2975 (N_2975,N_1926,N_1360);
or U2976 (N_2976,N_1017,N_1806);
nor U2977 (N_2977,N_1208,N_1103);
and U2978 (N_2978,N_1627,N_1162);
or U2979 (N_2979,N_1963,N_1848);
nand U2980 (N_2980,N_1016,N_1755);
nor U2981 (N_2981,N_1866,N_1590);
xnor U2982 (N_2982,N_1968,N_1531);
nor U2983 (N_2983,N_1421,N_1898);
and U2984 (N_2984,N_1752,N_1325);
nand U2985 (N_2985,N_1288,N_1642);
nor U2986 (N_2986,N_1131,N_1802);
and U2987 (N_2987,N_1119,N_1294);
and U2988 (N_2988,N_1111,N_1818);
nand U2989 (N_2989,N_1766,N_1973);
nand U2990 (N_2990,N_1293,N_1112);
or U2991 (N_2991,N_1279,N_1994);
nand U2992 (N_2992,N_1411,N_1787);
xnor U2993 (N_2993,N_1307,N_1439);
xnor U2994 (N_2994,N_1914,N_1105);
nand U2995 (N_2995,N_1006,N_1730);
and U2996 (N_2996,N_1341,N_1564);
and U2997 (N_2997,N_1046,N_1411);
nand U2998 (N_2998,N_1077,N_1232);
nor U2999 (N_2999,N_1006,N_1469);
or U3000 (N_3000,N_2575,N_2074);
or U3001 (N_3001,N_2578,N_2925);
and U3002 (N_3002,N_2482,N_2012);
and U3003 (N_3003,N_2121,N_2404);
nor U3004 (N_3004,N_2547,N_2180);
or U3005 (N_3005,N_2518,N_2468);
xor U3006 (N_3006,N_2480,N_2139);
or U3007 (N_3007,N_2185,N_2982);
and U3008 (N_3008,N_2513,N_2496);
nand U3009 (N_3009,N_2977,N_2862);
nor U3010 (N_3010,N_2786,N_2249);
or U3011 (N_3011,N_2576,N_2902);
or U3012 (N_3012,N_2668,N_2370);
and U3013 (N_3013,N_2057,N_2929);
nand U3014 (N_3014,N_2077,N_2069);
xor U3015 (N_3015,N_2564,N_2631);
nand U3016 (N_3016,N_2304,N_2520);
xnor U3017 (N_3017,N_2937,N_2936);
nor U3018 (N_3018,N_2403,N_2204);
nand U3019 (N_3019,N_2873,N_2845);
and U3020 (N_3020,N_2661,N_2365);
nor U3021 (N_3021,N_2466,N_2971);
nor U3022 (N_3022,N_2130,N_2424);
nor U3023 (N_3023,N_2470,N_2625);
xor U3024 (N_3024,N_2312,N_2944);
nand U3025 (N_3025,N_2748,N_2807);
or U3026 (N_3026,N_2267,N_2038);
nor U3027 (N_3027,N_2718,N_2755);
nor U3028 (N_3028,N_2372,N_2660);
and U3029 (N_3029,N_2603,N_2680);
xnor U3030 (N_3030,N_2949,N_2854);
nor U3031 (N_3031,N_2770,N_2635);
and U3032 (N_3032,N_2445,N_2962);
and U3033 (N_3033,N_2135,N_2871);
or U3034 (N_3034,N_2219,N_2539);
nor U3035 (N_3035,N_2504,N_2376);
and U3036 (N_3036,N_2068,N_2650);
xnor U3037 (N_3037,N_2286,N_2632);
nand U3038 (N_3038,N_2691,N_2614);
or U3039 (N_3039,N_2519,N_2450);
and U3040 (N_3040,N_2942,N_2550);
and U3041 (N_3041,N_2938,N_2382);
and U3042 (N_3042,N_2719,N_2455);
or U3043 (N_3043,N_2213,N_2960);
nand U3044 (N_3044,N_2869,N_2613);
xnor U3045 (N_3045,N_2533,N_2830);
xnor U3046 (N_3046,N_2302,N_2123);
or U3047 (N_3047,N_2900,N_2951);
nor U3048 (N_3048,N_2621,N_2574);
xor U3049 (N_3049,N_2825,N_2326);
nand U3050 (N_3050,N_2605,N_2541);
xnor U3051 (N_3051,N_2814,N_2790);
and U3052 (N_3052,N_2456,N_2910);
nor U3053 (N_3053,N_2051,N_2415);
nor U3054 (N_3054,N_2838,N_2627);
and U3055 (N_3055,N_2958,N_2281);
nand U3056 (N_3056,N_2345,N_2427);
nand U3057 (N_3057,N_2759,N_2463);
xnor U3058 (N_3058,N_2922,N_2887);
xor U3059 (N_3059,N_2610,N_2155);
or U3060 (N_3060,N_2913,N_2401);
xor U3061 (N_3061,N_2393,N_2102);
or U3062 (N_3062,N_2319,N_2842);
xor U3063 (N_3063,N_2216,N_2229);
or U3064 (N_3064,N_2484,N_2258);
nand U3065 (N_3065,N_2451,N_2098);
nor U3066 (N_3066,N_2201,N_2804);
nor U3067 (N_3067,N_2105,N_2889);
xnor U3068 (N_3068,N_2633,N_2572);
nand U3069 (N_3069,N_2993,N_2604);
or U3070 (N_3070,N_2757,N_2747);
xor U3071 (N_3071,N_2386,N_2018);
nor U3072 (N_3072,N_2122,N_2324);
or U3073 (N_3073,N_2502,N_2119);
or U3074 (N_3074,N_2964,N_2850);
and U3075 (N_3075,N_2313,N_2815);
and U3076 (N_3076,N_2876,N_2813);
or U3077 (N_3077,N_2367,N_2731);
nand U3078 (N_3078,N_2543,N_2493);
xor U3079 (N_3079,N_2992,N_2290);
nand U3080 (N_3080,N_2449,N_2760);
or U3081 (N_3081,N_2784,N_2301);
and U3082 (N_3082,N_2440,N_2341);
and U3083 (N_3083,N_2439,N_2835);
xnor U3084 (N_3084,N_2252,N_2497);
xor U3085 (N_3085,N_2752,N_2454);
xnor U3086 (N_3086,N_2309,N_2250);
xnor U3087 (N_3087,N_2965,N_2217);
nand U3088 (N_3088,N_2202,N_2526);
nand U3089 (N_3089,N_2148,N_2967);
and U3090 (N_3090,N_2316,N_2989);
or U3091 (N_3091,N_2169,N_2245);
and U3092 (N_3092,N_2344,N_2397);
nor U3093 (N_3093,N_2409,N_2273);
nor U3094 (N_3094,N_2348,N_2761);
or U3095 (N_3095,N_2713,N_2307);
and U3096 (N_3096,N_2940,N_2389);
and U3097 (N_3097,N_2059,N_2590);
or U3098 (N_3098,N_2985,N_2306);
nor U3099 (N_3099,N_2178,N_2003);
nor U3100 (N_3100,N_2154,N_2181);
nor U3101 (N_3101,N_2329,N_2241);
and U3102 (N_3102,N_2548,N_2930);
nor U3103 (N_3103,N_2226,N_2356);
and U3104 (N_3104,N_2189,N_2395);
nand U3105 (N_3105,N_2186,N_2948);
nor U3106 (N_3106,N_2157,N_2618);
or U3107 (N_3107,N_2089,N_2810);
or U3108 (N_3108,N_2460,N_2638);
nand U3109 (N_3109,N_2061,N_2086);
and U3110 (N_3110,N_2336,N_2612);
xor U3111 (N_3111,N_2999,N_2143);
nor U3112 (N_3112,N_2616,N_2005);
nor U3113 (N_3113,N_2198,N_2602);
nor U3114 (N_3114,N_2834,N_2723);
and U3115 (N_3115,N_2560,N_2857);
or U3116 (N_3116,N_2821,N_2779);
or U3117 (N_3117,N_2371,N_2600);
and U3118 (N_3118,N_2729,N_2274);
xnor U3119 (N_3119,N_2224,N_2682);
nand U3120 (N_3120,N_2002,N_2159);
nor U3121 (N_3121,N_2352,N_2311);
nand U3122 (N_3122,N_2990,N_2218);
nand U3123 (N_3123,N_2400,N_2298);
nand U3124 (N_3124,N_2461,N_2407);
nor U3125 (N_3125,N_2953,N_2820);
xor U3126 (N_3126,N_2765,N_2266);
or U3127 (N_3127,N_2565,N_2885);
and U3128 (N_3128,N_2177,N_2007);
or U3129 (N_3129,N_2692,N_2487);
nor U3130 (N_3130,N_2742,N_2055);
xnor U3131 (N_3131,N_2209,N_2881);
and U3132 (N_3132,N_2131,N_2349);
xor U3133 (N_3133,N_2555,N_2724);
or U3134 (N_3134,N_2655,N_2524);
or U3135 (N_3135,N_2399,N_2727);
and U3136 (N_3136,N_2705,N_2529);
xnor U3137 (N_3137,N_2628,N_2561);
nand U3138 (N_3138,N_2874,N_2553);
or U3139 (N_3139,N_2912,N_2084);
and U3140 (N_3140,N_2340,N_2596);
nand U3141 (N_3141,N_2014,N_2787);
xor U3142 (N_3142,N_2983,N_2859);
xnor U3143 (N_3143,N_2571,N_2443);
xor U3144 (N_3144,N_2355,N_2556);
or U3145 (N_3145,N_2935,N_2646);
or U3146 (N_3146,N_2745,N_2898);
and U3147 (N_3147,N_2617,N_2630);
nor U3148 (N_3148,N_2715,N_2535);
xnor U3149 (N_3149,N_2684,N_2398);
and U3150 (N_3150,N_2255,N_2280);
or U3151 (N_3151,N_2583,N_2128);
nor U3152 (N_3152,N_2537,N_2926);
or U3153 (N_3153,N_2994,N_2700);
and U3154 (N_3154,N_2001,N_2021);
nand U3155 (N_3155,N_2829,N_2338);
xnor U3156 (N_3156,N_2697,N_2961);
and U3157 (N_3157,N_2441,N_2896);
and U3158 (N_3158,N_2040,N_2864);
nor U3159 (N_3159,N_2525,N_2422);
or U3160 (N_3160,N_2416,N_2284);
and U3161 (N_3161,N_2943,N_2923);
xnor U3162 (N_3162,N_2256,N_2762);
and U3163 (N_3163,N_2557,N_2952);
xor U3164 (N_3164,N_2781,N_2243);
xor U3165 (N_3165,N_2136,N_2322);
nor U3166 (N_3166,N_2037,N_2152);
or U3167 (N_3167,N_2380,N_2421);
nor U3168 (N_3168,N_2698,N_2467);
or U3169 (N_3169,N_2819,N_2702);
nand U3170 (N_3170,N_2963,N_2891);
or U3171 (N_3171,N_2469,N_2447);
nor U3172 (N_3172,N_2199,N_2282);
nor U3173 (N_3173,N_2088,N_2031);
nor U3174 (N_3174,N_2688,N_2339);
and U3175 (N_3175,N_2689,N_2150);
nor U3176 (N_3176,N_2653,N_2183);
and U3177 (N_3177,N_2234,N_2894);
or U3178 (N_3178,N_2453,N_2151);
nor U3179 (N_3179,N_2945,N_2333);
nor U3180 (N_3180,N_2300,N_2235);
nand U3181 (N_3181,N_2562,N_2364);
nand U3182 (N_3182,N_2052,N_2078);
nand U3183 (N_3183,N_2939,N_2946);
nor U3184 (N_3184,N_2405,N_2414);
xnor U3185 (N_3185,N_2207,N_2381);
and U3186 (N_3186,N_2335,N_2764);
xor U3187 (N_3187,N_2858,N_2573);
xor U3188 (N_3188,N_2064,N_2275);
nand U3189 (N_3189,N_2413,N_2514);
xor U3190 (N_3190,N_2419,N_2641);
xnor U3191 (N_3191,N_2357,N_2114);
nand U3192 (N_3192,N_2297,N_2107);
xnor U3193 (N_3193,N_2906,N_2438);
or U3194 (N_3194,N_2483,N_2903);
and U3195 (N_3195,N_2546,N_2998);
and U3196 (N_3196,N_2020,N_2346);
xnor U3197 (N_3197,N_2362,N_2363);
xor U3198 (N_3198,N_2791,N_2584);
xnor U3199 (N_3199,N_2412,N_2408);
or U3200 (N_3200,N_2782,N_2991);
xnor U3201 (N_3201,N_2818,N_2097);
nor U3202 (N_3202,N_2009,N_2677);
nor U3203 (N_3203,N_2809,N_2656);
nor U3204 (N_3204,N_2563,N_2108);
xor U3205 (N_3205,N_2006,N_2921);
or U3206 (N_3206,N_2916,N_2260);
and U3207 (N_3207,N_2211,N_2144);
nand U3208 (N_3208,N_2797,N_2036);
nand U3209 (N_3209,N_2772,N_2875);
and U3210 (N_3210,N_2802,N_2795);
and U3211 (N_3211,N_2651,N_2227);
or U3212 (N_3212,N_2843,N_2827);
nor U3213 (N_3213,N_2026,N_2970);
and U3214 (N_3214,N_2465,N_2058);
nand U3215 (N_3215,N_2033,N_2740);
xor U3216 (N_3216,N_2116,N_2318);
xor U3217 (N_3217,N_2411,N_2515);
nor U3218 (N_3218,N_2428,N_2197);
xor U3219 (N_3219,N_2360,N_2492);
and U3220 (N_3220,N_2920,N_2657);
xnor U3221 (N_3221,N_2048,N_2221);
and U3222 (N_3222,N_2662,N_2279);
and U3223 (N_3223,N_2457,N_2793);
nor U3224 (N_3224,N_2384,N_2704);
nor U3225 (N_3225,N_2706,N_2133);
or U3226 (N_3226,N_2359,N_2402);
nand U3227 (N_3227,N_2278,N_2041);
or U3228 (N_3228,N_2353,N_2096);
xnor U3229 (N_3229,N_2941,N_2172);
xor U3230 (N_3230,N_2194,N_2373);
xnor U3231 (N_3231,N_2436,N_2200);
or U3232 (N_3232,N_2321,N_2308);
and U3233 (N_3233,N_2490,N_2905);
or U3234 (N_3234,N_2974,N_2113);
or U3235 (N_3235,N_2248,N_2852);
and U3236 (N_3236,N_2622,N_2390);
nand U3237 (N_3237,N_2594,N_2671);
nor U3238 (N_3238,N_2554,N_2531);
or U3239 (N_3239,N_2826,N_2124);
nor U3240 (N_3240,N_2510,N_2709);
xnor U3241 (N_3241,N_2410,N_2085);
xnor U3242 (N_3242,N_2008,N_2882);
and U3243 (N_3243,N_2317,N_2979);
xnor U3244 (N_3244,N_2247,N_2231);
nor U3245 (N_3245,N_2687,N_2425);
nand U3246 (N_3246,N_2534,N_2517);
nand U3247 (N_3247,N_2824,N_2379);
and U3248 (N_3248,N_2292,N_2039);
nand U3249 (N_3249,N_2435,N_2558);
and U3250 (N_3250,N_2822,N_2711);
nand U3251 (N_3251,N_2062,N_2969);
and U3252 (N_3252,N_2647,N_2035);
xnor U3253 (N_3253,N_2836,N_2735);
or U3254 (N_3254,N_2276,N_2832);
nor U3255 (N_3255,N_2010,N_2023);
and U3256 (N_3256,N_2240,N_2908);
nand U3257 (N_3257,N_2475,N_2075);
and U3258 (N_3258,N_2566,N_2892);
and U3259 (N_3259,N_2996,N_2210);
and U3260 (N_3260,N_2029,N_2609);
nand U3261 (N_3261,N_2054,N_2066);
xor U3262 (N_3262,N_2174,N_2385);
or U3263 (N_3263,N_2263,N_2888);
nor U3264 (N_3264,N_2672,N_2592);
and U3265 (N_3265,N_2184,N_2714);
xnor U3266 (N_3266,N_2540,N_2375);
or U3267 (N_3267,N_2693,N_2294);
nand U3268 (N_3268,N_2866,N_2289);
or U3269 (N_3269,N_2658,N_2883);
and U3270 (N_3270,N_2620,N_2473);
or U3271 (N_3271,N_2471,N_2654);
nor U3272 (N_3272,N_2019,N_2751);
nor U3273 (N_3273,N_2806,N_2391);
or U3274 (N_3274,N_2611,N_2966);
xnor U3275 (N_3275,N_2865,N_2997);
nor U3276 (N_3276,N_2481,N_2060);
nor U3277 (N_3277,N_2917,N_2728);
nor U3278 (N_3278,N_2071,N_2214);
and U3279 (N_3279,N_2238,N_2732);
nand U3280 (N_3280,N_2474,N_2499);
nand U3281 (N_3281,N_2636,N_2674);
nor U3282 (N_3282,N_2277,N_2890);
and U3283 (N_3283,N_2142,N_2860);
and U3284 (N_3284,N_2004,N_2577);
nor U3285 (N_3285,N_2237,N_2511);
or U3286 (N_3286,N_2595,N_2545);
and U3287 (N_3287,N_2532,N_2032);
xnor U3288 (N_3288,N_2118,N_2233);
nor U3289 (N_3289,N_2053,N_2464);
nor U3290 (N_3290,N_2291,N_2642);
nand U3291 (N_3291,N_2244,N_2643);
nor U3292 (N_3292,N_2739,N_2090);
nor U3293 (N_3293,N_2675,N_2726);
or U3294 (N_3294,N_2288,N_2160);
xor U3295 (N_3295,N_2011,N_2507);
and U3296 (N_3296,N_2833,N_2980);
nor U3297 (N_3297,N_2472,N_2498);
nor U3298 (N_3298,N_2738,N_2506);
nand U3299 (N_3299,N_2853,N_2663);
nor U3300 (N_3300,N_2195,N_2153);
or U3301 (N_3301,N_2615,N_2597);
and U3302 (N_3302,N_2394,N_2823);
or U3303 (N_3303,N_2582,N_2171);
xnor U3304 (N_3304,N_2261,N_2426);
or U3305 (N_3305,N_2901,N_2623);
nand U3306 (N_3306,N_2867,N_2768);
and U3307 (N_3307,N_2325,N_2608);
nand U3308 (N_3308,N_2034,N_2667);
or U3309 (N_3309,N_2968,N_2117);
xor U3310 (N_3310,N_2350,N_2591);
nor U3311 (N_3311,N_2374,N_2388);
nand U3312 (N_3312,N_2168,N_2984);
or U3313 (N_3313,N_2722,N_2588);
nor U3314 (N_3314,N_2988,N_2841);
or U3315 (N_3315,N_2268,N_2670);
or U3316 (N_3316,N_2067,N_2708);
xnor U3317 (N_3317,N_2569,N_2769);
nor U3318 (N_3318,N_2756,N_2334);
nand U3319 (N_3319,N_2446,N_2796);
nand U3320 (N_3320,N_2570,N_2432);
nor U3321 (N_3321,N_2778,N_2629);
nor U3322 (N_3322,N_2236,N_2173);
xnor U3323 (N_3323,N_2170,N_2503);
and U3324 (N_3324,N_2521,N_2758);
and U3325 (N_3325,N_2530,N_2000);
xor U3326 (N_3326,N_2265,N_2127);
or U3327 (N_3327,N_2478,N_2931);
nand U3328 (N_3328,N_2690,N_2082);
nor U3329 (N_3329,N_2861,N_2817);
nor U3330 (N_3330,N_2911,N_2598);
or U3331 (N_3331,N_2111,N_2848);
nor U3332 (N_3332,N_2494,N_2417);
and U3333 (N_3333,N_2163,N_2396);
nor U3334 (N_3334,N_2717,N_2212);
nor U3335 (N_3335,N_2895,N_2789);
and U3336 (N_3336,N_2253,N_2269);
and U3337 (N_3337,N_2452,N_2954);
and U3338 (N_3338,N_2634,N_2030);
and U3339 (N_3339,N_2192,N_2673);
or U3340 (N_3340,N_2924,N_2816);
or U3341 (N_3341,N_2846,N_2305);
nand U3342 (N_3342,N_2347,N_2271);
xor U3343 (N_3343,N_2190,N_2933);
xor U3344 (N_3344,N_2188,N_2934);
xor U3345 (N_3345,N_2872,N_2103);
nor U3346 (N_3346,N_2044,N_2262);
nand U3347 (N_3347,N_2840,N_2856);
nand U3348 (N_3348,N_2710,N_2129);
xor U3349 (N_3349,N_2794,N_2196);
and U3350 (N_3350,N_2205,N_2730);
nand U3351 (N_3351,N_2459,N_2559);
nand U3352 (N_3352,N_2431,N_2328);
nor U3353 (N_3353,N_2106,N_2509);
nand U3354 (N_3354,N_2215,N_2736);
nand U3355 (N_3355,N_2283,N_2914);
nand U3356 (N_3356,N_2287,N_2792);
or U3357 (N_3357,N_2429,N_2330);
nand U3358 (N_3358,N_2230,N_2270);
nand U3359 (N_3359,N_2703,N_2028);
nand U3360 (N_3360,N_2799,N_2685);
nor U3361 (N_3361,N_2141,N_2254);
and U3362 (N_3362,N_2145,N_2580);
nand U3363 (N_3363,N_2805,N_2904);
and U3364 (N_3364,N_2343,N_2686);
nor U3365 (N_3365,N_2976,N_2387);
xnor U3366 (N_3366,N_2072,N_2392);
or U3367 (N_3367,N_2665,N_2716);
or U3368 (N_3368,N_2744,N_2909);
or U3369 (N_3369,N_2331,N_2080);
or U3370 (N_3370,N_2015,N_2522);
xnor U3371 (N_3371,N_2310,N_2299);
and U3372 (N_3372,N_2458,N_2076);
or U3373 (N_3373,N_2678,N_2637);
nand U3374 (N_3374,N_2406,N_2491);
nor U3375 (N_3375,N_2050,N_2043);
and U3376 (N_3376,N_2182,N_2495);
xor U3377 (N_3377,N_2899,N_2448);
and U3378 (N_3378,N_2978,N_2783);
and U3379 (N_3379,N_2272,N_2093);
and U3380 (N_3380,N_2045,N_2206);
nand U3381 (N_3381,N_2763,N_2919);
nor U3382 (N_3382,N_2679,N_2973);
nor U3383 (N_3383,N_2955,N_2528);
xor U3384 (N_3384,N_2844,N_2489);
nor U3385 (N_3385,N_2303,N_2523);
nand U3386 (N_3386,N_2947,N_2042);
xor U3387 (N_3387,N_2549,N_2886);
xnor U3388 (N_3388,N_2957,N_2928);
nor U3389 (N_3389,N_2542,N_2434);
or U3390 (N_3390,N_2741,N_2505);
nor U3391 (N_3391,N_2743,N_2239);
or U3392 (N_3392,N_2771,N_2327);
or U3393 (N_3393,N_2847,N_2203);
or U3394 (N_3394,N_2798,N_2536);
or U3395 (N_3395,N_2046,N_2579);
or U3396 (N_3396,N_2430,N_2223);
and U3397 (N_3397,N_2950,N_2165);
xor U3398 (N_3398,N_2158,N_2567);
nand U3399 (N_3399,N_2749,N_2228);
nand U3400 (N_3400,N_2296,N_2812);
nand U3401 (N_3401,N_2878,N_2378);
nand U3402 (N_3402,N_2433,N_2485);
nor U3403 (N_3403,N_2442,N_2516);
and U3404 (N_3404,N_2259,N_2087);
nor U3405 (N_3405,N_2737,N_2022);
or U3406 (N_3406,N_2601,N_2666);
nor U3407 (N_3407,N_2712,N_2208);
nand U3408 (N_3408,N_2956,N_2104);
or U3409 (N_3409,N_2607,N_2323);
nor U3410 (N_3410,N_2056,N_2100);
and U3411 (N_3411,N_2897,N_2314);
or U3412 (N_3412,N_2175,N_2870);
and U3413 (N_3413,N_2986,N_2676);
xor U3414 (N_3414,N_2780,N_2225);
nor U3415 (N_3415,N_2664,N_2242);
nand U3416 (N_3416,N_2351,N_2981);
or U3417 (N_3417,N_2880,N_2293);
nand U3418 (N_3418,N_2652,N_2187);
and U3419 (N_3419,N_2753,N_2893);
nor U3420 (N_3420,N_2149,N_2884);
nor U3421 (N_3421,N_2734,N_2927);
or U3422 (N_3422,N_2354,N_2808);
nor U3423 (N_3423,N_2444,N_2095);
nor U3424 (N_3424,N_2285,N_2788);
xor U3425 (N_3425,N_2079,N_2049);
and U3426 (N_3426,N_2251,N_2707);
and U3427 (N_3427,N_2777,N_2500);
nor U3428 (N_3428,N_2645,N_2501);
nand U3429 (N_3429,N_2773,N_2644);
or U3430 (N_3430,N_2776,N_2420);
nor U3431 (N_3431,N_2918,N_2746);
nor U3432 (N_3432,N_2094,N_2027);
or U3433 (N_3433,N_2972,N_2147);
nand U3434 (N_3434,N_2669,N_2868);
xor U3435 (N_3435,N_2377,N_2366);
and U3436 (N_3436,N_2774,N_2161);
and U3437 (N_3437,N_2120,N_2099);
nand U3438 (N_3438,N_2101,N_2073);
nand U3439 (N_3439,N_2619,N_2606);
xor U3440 (N_3440,N_2767,N_2179);
xnor U3441 (N_3441,N_2358,N_2721);
or U3442 (N_3442,N_2166,N_2138);
xor U3443 (N_3443,N_2092,N_2725);
and U3444 (N_3444,N_2855,N_2295);
xor U3445 (N_3445,N_2125,N_2863);
nor U3446 (N_3446,N_2477,N_2342);
and U3447 (N_3447,N_2839,N_2837);
nor U3448 (N_3448,N_2959,N_2167);
nor U3449 (N_3449,N_2222,N_2681);
xnor U3450 (N_3450,N_2733,N_2091);
nand U3451 (N_3451,N_2640,N_2476);
xnor U3452 (N_3452,N_2879,N_2626);
nand U3453 (N_3453,N_2538,N_2877);
nand U3454 (N_3454,N_2695,N_2112);
and U3455 (N_3455,N_2599,N_2720);
xnor U3456 (N_3456,N_2081,N_2849);
nand U3457 (N_3457,N_2126,N_2585);
xor U3458 (N_3458,N_2552,N_2368);
or U3459 (N_3459,N_2070,N_2975);
nand U3460 (N_3460,N_2544,N_2551);
and U3461 (N_3461,N_2264,N_2315);
nor U3462 (N_3462,N_2479,N_2587);
nand U3463 (N_3463,N_2132,N_2013);
and U3464 (N_3464,N_2176,N_2025);
or U3465 (N_3465,N_2320,N_2361);
and U3466 (N_3466,N_2232,N_2811);
nor U3467 (N_3467,N_2191,N_2801);
xnor U3468 (N_3468,N_2047,N_2115);
nor U3469 (N_3469,N_2593,N_2462);
nand U3470 (N_3470,N_2624,N_2156);
xor U3471 (N_3471,N_2508,N_2696);
xnor U3472 (N_3472,N_2146,N_2137);
nor U3473 (N_3473,N_2683,N_2828);
and U3474 (N_3474,N_2527,N_2418);
nor U3475 (N_3475,N_2162,N_2750);
or U3476 (N_3476,N_2987,N_2851);
nand U3477 (N_3477,N_2766,N_2065);
xnor U3478 (N_3478,N_2775,N_2140);
and U3479 (N_3479,N_2383,N_2659);
and U3480 (N_3480,N_2932,N_2134);
and U3481 (N_3481,N_2803,N_2699);
nor U3482 (N_3482,N_2831,N_2995);
nor U3483 (N_3483,N_2332,N_2164);
xor U3484 (N_3484,N_2369,N_2488);
and U3485 (N_3485,N_2694,N_2109);
and U3486 (N_3486,N_2701,N_2512);
xor U3487 (N_3487,N_2220,N_2193);
nor U3488 (N_3488,N_2639,N_2024);
nor U3489 (N_3489,N_2581,N_2063);
nand U3490 (N_3490,N_2083,N_2486);
or U3491 (N_3491,N_2437,N_2423);
and U3492 (N_3492,N_2915,N_2337);
or U3493 (N_3493,N_2648,N_2907);
and U3494 (N_3494,N_2017,N_2785);
xnor U3495 (N_3495,N_2800,N_2257);
nor U3496 (N_3496,N_2754,N_2568);
nand U3497 (N_3497,N_2589,N_2586);
nor U3498 (N_3498,N_2246,N_2110);
and U3499 (N_3499,N_2016,N_2649);
nand U3500 (N_3500,N_2272,N_2886);
or U3501 (N_3501,N_2843,N_2593);
nor U3502 (N_3502,N_2092,N_2121);
nor U3503 (N_3503,N_2363,N_2338);
xor U3504 (N_3504,N_2281,N_2635);
nand U3505 (N_3505,N_2736,N_2765);
nand U3506 (N_3506,N_2960,N_2915);
nand U3507 (N_3507,N_2494,N_2364);
and U3508 (N_3508,N_2037,N_2894);
xor U3509 (N_3509,N_2303,N_2878);
xor U3510 (N_3510,N_2440,N_2073);
nand U3511 (N_3511,N_2510,N_2879);
xor U3512 (N_3512,N_2049,N_2889);
xor U3513 (N_3513,N_2553,N_2391);
nand U3514 (N_3514,N_2655,N_2663);
xor U3515 (N_3515,N_2955,N_2584);
and U3516 (N_3516,N_2170,N_2340);
or U3517 (N_3517,N_2912,N_2821);
nand U3518 (N_3518,N_2075,N_2534);
or U3519 (N_3519,N_2213,N_2405);
and U3520 (N_3520,N_2507,N_2297);
xor U3521 (N_3521,N_2317,N_2415);
xnor U3522 (N_3522,N_2308,N_2804);
nand U3523 (N_3523,N_2051,N_2438);
and U3524 (N_3524,N_2870,N_2979);
and U3525 (N_3525,N_2800,N_2951);
or U3526 (N_3526,N_2077,N_2188);
xnor U3527 (N_3527,N_2713,N_2174);
nor U3528 (N_3528,N_2355,N_2906);
nor U3529 (N_3529,N_2287,N_2252);
nor U3530 (N_3530,N_2536,N_2467);
or U3531 (N_3531,N_2949,N_2506);
nor U3532 (N_3532,N_2507,N_2965);
and U3533 (N_3533,N_2083,N_2161);
nand U3534 (N_3534,N_2184,N_2838);
xor U3535 (N_3535,N_2576,N_2016);
nand U3536 (N_3536,N_2848,N_2824);
nand U3537 (N_3537,N_2082,N_2456);
xnor U3538 (N_3538,N_2636,N_2215);
and U3539 (N_3539,N_2977,N_2085);
or U3540 (N_3540,N_2677,N_2797);
xor U3541 (N_3541,N_2044,N_2679);
xor U3542 (N_3542,N_2359,N_2558);
or U3543 (N_3543,N_2596,N_2789);
and U3544 (N_3544,N_2423,N_2063);
xnor U3545 (N_3545,N_2937,N_2794);
nor U3546 (N_3546,N_2928,N_2203);
or U3547 (N_3547,N_2732,N_2818);
nand U3548 (N_3548,N_2008,N_2716);
and U3549 (N_3549,N_2566,N_2835);
and U3550 (N_3550,N_2109,N_2951);
or U3551 (N_3551,N_2945,N_2376);
xor U3552 (N_3552,N_2933,N_2979);
or U3553 (N_3553,N_2775,N_2856);
nand U3554 (N_3554,N_2235,N_2936);
xor U3555 (N_3555,N_2926,N_2994);
nor U3556 (N_3556,N_2585,N_2252);
and U3557 (N_3557,N_2906,N_2808);
xnor U3558 (N_3558,N_2348,N_2595);
or U3559 (N_3559,N_2862,N_2451);
xnor U3560 (N_3560,N_2740,N_2759);
nor U3561 (N_3561,N_2404,N_2811);
xnor U3562 (N_3562,N_2641,N_2566);
nor U3563 (N_3563,N_2643,N_2359);
nand U3564 (N_3564,N_2097,N_2389);
nand U3565 (N_3565,N_2604,N_2343);
nor U3566 (N_3566,N_2679,N_2582);
or U3567 (N_3567,N_2708,N_2008);
xor U3568 (N_3568,N_2344,N_2485);
and U3569 (N_3569,N_2547,N_2785);
nand U3570 (N_3570,N_2424,N_2522);
xor U3571 (N_3571,N_2020,N_2238);
or U3572 (N_3572,N_2176,N_2393);
and U3573 (N_3573,N_2324,N_2747);
xnor U3574 (N_3574,N_2511,N_2513);
nand U3575 (N_3575,N_2324,N_2111);
or U3576 (N_3576,N_2660,N_2052);
and U3577 (N_3577,N_2169,N_2529);
nand U3578 (N_3578,N_2949,N_2175);
xor U3579 (N_3579,N_2471,N_2736);
nor U3580 (N_3580,N_2124,N_2157);
xnor U3581 (N_3581,N_2154,N_2850);
nor U3582 (N_3582,N_2624,N_2412);
nand U3583 (N_3583,N_2044,N_2934);
or U3584 (N_3584,N_2055,N_2637);
nor U3585 (N_3585,N_2579,N_2599);
nor U3586 (N_3586,N_2626,N_2549);
nand U3587 (N_3587,N_2578,N_2574);
xnor U3588 (N_3588,N_2780,N_2499);
xor U3589 (N_3589,N_2351,N_2445);
and U3590 (N_3590,N_2406,N_2061);
nor U3591 (N_3591,N_2758,N_2455);
nor U3592 (N_3592,N_2971,N_2068);
nand U3593 (N_3593,N_2852,N_2471);
xor U3594 (N_3594,N_2467,N_2331);
nand U3595 (N_3595,N_2653,N_2997);
xnor U3596 (N_3596,N_2897,N_2648);
nor U3597 (N_3597,N_2238,N_2642);
or U3598 (N_3598,N_2573,N_2274);
nand U3599 (N_3599,N_2450,N_2542);
xnor U3600 (N_3600,N_2828,N_2285);
nand U3601 (N_3601,N_2377,N_2583);
xor U3602 (N_3602,N_2693,N_2944);
xor U3603 (N_3603,N_2153,N_2630);
and U3604 (N_3604,N_2981,N_2571);
nand U3605 (N_3605,N_2369,N_2408);
nor U3606 (N_3606,N_2102,N_2098);
nand U3607 (N_3607,N_2894,N_2011);
nor U3608 (N_3608,N_2589,N_2217);
xor U3609 (N_3609,N_2659,N_2281);
nand U3610 (N_3610,N_2331,N_2912);
or U3611 (N_3611,N_2228,N_2471);
nor U3612 (N_3612,N_2209,N_2297);
nand U3613 (N_3613,N_2846,N_2467);
and U3614 (N_3614,N_2314,N_2296);
nor U3615 (N_3615,N_2434,N_2088);
xor U3616 (N_3616,N_2264,N_2081);
nor U3617 (N_3617,N_2248,N_2302);
nor U3618 (N_3618,N_2250,N_2022);
and U3619 (N_3619,N_2354,N_2743);
xnor U3620 (N_3620,N_2569,N_2394);
and U3621 (N_3621,N_2534,N_2229);
nand U3622 (N_3622,N_2321,N_2814);
and U3623 (N_3623,N_2720,N_2637);
or U3624 (N_3624,N_2488,N_2572);
nor U3625 (N_3625,N_2865,N_2019);
nand U3626 (N_3626,N_2534,N_2174);
nor U3627 (N_3627,N_2426,N_2922);
or U3628 (N_3628,N_2826,N_2130);
xor U3629 (N_3629,N_2397,N_2902);
and U3630 (N_3630,N_2988,N_2295);
and U3631 (N_3631,N_2987,N_2058);
and U3632 (N_3632,N_2246,N_2951);
nand U3633 (N_3633,N_2550,N_2514);
xnor U3634 (N_3634,N_2521,N_2948);
and U3635 (N_3635,N_2249,N_2541);
and U3636 (N_3636,N_2720,N_2764);
and U3637 (N_3637,N_2264,N_2351);
and U3638 (N_3638,N_2512,N_2369);
xor U3639 (N_3639,N_2015,N_2592);
nand U3640 (N_3640,N_2301,N_2569);
xnor U3641 (N_3641,N_2769,N_2386);
or U3642 (N_3642,N_2056,N_2475);
xnor U3643 (N_3643,N_2634,N_2588);
nor U3644 (N_3644,N_2310,N_2642);
nand U3645 (N_3645,N_2841,N_2281);
and U3646 (N_3646,N_2225,N_2346);
nand U3647 (N_3647,N_2231,N_2712);
nand U3648 (N_3648,N_2494,N_2316);
nor U3649 (N_3649,N_2959,N_2667);
or U3650 (N_3650,N_2160,N_2715);
xor U3651 (N_3651,N_2111,N_2628);
nand U3652 (N_3652,N_2113,N_2991);
and U3653 (N_3653,N_2552,N_2687);
xnor U3654 (N_3654,N_2967,N_2636);
nor U3655 (N_3655,N_2417,N_2112);
or U3656 (N_3656,N_2747,N_2912);
nand U3657 (N_3657,N_2208,N_2211);
nor U3658 (N_3658,N_2804,N_2023);
xor U3659 (N_3659,N_2446,N_2851);
xor U3660 (N_3660,N_2807,N_2535);
and U3661 (N_3661,N_2872,N_2489);
nand U3662 (N_3662,N_2229,N_2398);
and U3663 (N_3663,N_2054,N_2185);
nand U3664 (N_3664,N_2980,N_2227);
and U3665 (N_3665,N_2054,N_2127);
nand U3666 (N_3666,N_2792,N_2510);
nand U3667 (N_3667,N_2164,N_2545);
or U3668 (N_3668,N_2861,N_2522);
nand U3669 (N_3669,N_2258,N_2240);
or U3670 (N_3670,N_2827,N_2929);
nor U3671 (N_3671,N_2708,N_2911);
and U3672 (N_3672,N_2835,N_2119);
and U3673 (N_3673,N_2835,N_2417);
or U3674 (N_3674,N_2557,N_2794);
nor U3675 (N_3675,N_2423,N_2226);
nand U3676 (N_3676,N_2578,N_2130);
nand U3677 (N_3677,N_2640,N_2772);
xor U3678 (N_3678,N_2350,N_2359);
nand U3679 (N_3679,N_2084,N_2183);
and U3680 (N_3680,N_2022,N_2618);
xnor U3681 (N_3681,N_2664,N_2508);
nor U3682 (N_3682,N_2199,N_2090);
or U3683 (N_3683,N_2539,N_2473);
and U3684 (N_3684,N_2885,N_2771);
or U3685 (N_3685,N_2579,N_2982);
xor U3686 (N_3686,N_2550,N_2558);
or U3687 (N_3687,N_2907,N_2276);
and U3688 (N_3688,N_2098,N_2308);
nor U3689 (N_3689,N_2142,N_2864);
and U3690 (N_3690,N_2657,N_2450);
or U3691 (N_3691,N_2162,N_2846);
nor U3692 (N_3692,N_2570,N_2917);
and U3693 (N_3693,N_2780,N_2286);
nor U3694 (N_3694,N_2545,N_2306);
xor U3695 (N_3695,N_2445,N_2111);
nor U3696 (N_3696,N_2662,N_2448);
nor U3697 (N_3697,N_2293,N_2906);
or U3698 (N_3698,N_2002,N_2548);
and U3699 (N_3699,N_2748,N_2243);
xnor U3700 (N_3700,N_2684,N_2824);
nand U3701 (N_3701,N_2437,N_2683);
xnor U3702 (N_3702,N_2006,N_2997);
xnor U3703 (N_3703,N_2711,N_2758);
or U3704 (N_3704,N_2761,N_2405);
and U3705 (N_3705,N_2569,N_2665);
and U3706 (N_3706,N_2900,N_2416);
nand U3707 (N_3707,N_2696,N_2021);
nand U3708 (N_3708,N_2041,N_2014);
and U3709 (N_3709,N_2407,N_2244);
or U3710 (N_3710,N_2152,N_2793);
or U3711 (N_3711,N_2300,N_2680);
nand U3712 (N_3712,N_2202,N_2080);
and U3713 (N_3713,N_2950,N_2922);
and U3714 (N_3714,N_2281,N_2760);
or U3715 (N_3715,N_2925,N_2541);
nor U3716 (N_3716,N_2395,N_2280);
nand U3717 (N_3717,N_2421,N_2618);
xor U3718 (N_3718,N_2870,N_2926);
xor U3719 (N_3719,N_2855,N_2448);
nand U3720 (N_3720,N_2885,N_2545);
and U3721 (N_3721,N_2477,N_2910);
nand U3722 (N_3722,N_2599,N_2435);
nor U3723 (N_3723,N_2338,N_2023);
or U3724 (N_3724,N_2483,N_2823);
nor U3725 (N_3725,N_2346,N_2948);
nor U3726 (N_3726,N_2488,N_2495);
nand U3727 (N_3727,N_2750,N_2010);
nand U3728 (N_3728,N_2867,N_2302);
or U3729 (N_3729,N_2945,N_2603);
nand U3730 (N_3730,N_2297,N_2711);
xnor U3731 (N_3731,N_2045,N_2394);
nand U3732 (N_3732,N_2096,N_2465);
or U3733 (N_3733,N_2153,N_2178);
nor U3734 (N_3734,N_2354,N_2735);
nand U3735 (N_3735,N_2031,N_2699);
nor U3736 (N_3736,N_2614,N_2290);
and U3737 (N_3737,N_2375,N_2959);
and U3738 (N_3738,N_2359,N_2395);
or U3739 (N_3739,N_2665,N_2007);
nor U3740 (N_3740,N_2804,N_2642);
and U3741 (N_3741,N_2614,N_2028);
xnor U3742 (N_3742,N_2281,N_2874);
nand U3743 (N_3743,N_2857,N_2087);
xnor U3744 (N_3744,N_2204,N_2901);
or U3745 (N_3745,N_2885,N_2433);
nand U3746 (N_3746,N_2460,N_2075);
xnor U3747 (N_3747,N_2197,N_2127);
xnor U3748 (N_3748,N_2747,N_2799);
nor U3749 (N_3749,N_2328,N_2581);
xnor U3750 (N_3750,N_2433,N_2828);
and U3751 (N_3751,N_2424,N_2951);
nor U3752 (N_3752,N_2494,N_2894);
nor U3753 (N_3753,N_2395,N_2781);
nand U3754 (N_3754,N_2869,N_2052);
xnor U3755 (N_3755,N_2544,N_2325);
nor U3756 (N_3756,N_2459,N_2472);
nand U3757 (N_3757,N_2715,N_2132);
nand U3758 (N_3758,N_2809,N_2101);
nor U3759 (N_3759,N_2201,N_2462);
and U3760 (N_3760,N_2481,N_2585);
nand U3761 (N_3761,N_2102,N_2166);
nand U3762 (N_3762,N_2709,N_2388);
nor U3763 (N_3763,N_2660,N_2965);
or U3764 (N_3764,N_2785,N_2370);
nand U3765 (N_3765,N_2728,N_2514);
xor U3766 (N_3766,N_2556,N_2474);
nand U3767 (N_3767,N_2723,N_2578);
and U3768 (N_3768,N_2312,N_2719);
or U3769 (N_3769,N_2153,N_2845);
nand U3770 (N_3770,N_2860,N_2103);
nor U3771 (N_3771,N_2485,N_2648);
or U3772 (N_3772,N_2742,N_2257);
nor U3773 (N_3773,N_2132,N_2050);
and U3774 (N_3774,N_2114,N_2638);
nor U3775 (N_3775,N_2253,N_2332);
and U3776 (N_3776,N_2997,N_2470);
nand U3777 (N_3777,N_2684,N_2268);
nand U3778 (N_3778,N_2661,N_2586);
or U3779 (N_3779,N_2868,N_2730);
nor U3780 (N_3780,N_2570,N_2367);
xor U3781 (N_3781,N_2696,N_2148);
nor U3782 (N_3782,N_2222,N_2818);
or U3783 (N_3783,N_2178,N_2742);
or U3784 (N_3784,N_2761,N_2290);
or U3785 (N_3785,N_2186,N_2388);
nand U3786 (N_3786,N_2303,N_2888);
xor U3787 (N_3787,N_2810,N_2247);
nand U3788 (N_3788,N_2590,N_2979);
nor U3789 (N_3789,N_2278,N_2540);
xnor U3790 (N_3790,N_2815,N_2739);
and U3791 (N_3791,N_2487,N_2147);
and U3792 (N_3792,N_2201,N_2748);
or U3793 (N_3793,N_2626,N_2412);
nand U3794 (N_3794,N_2812,N_2336);
nand U3795 (N_3795,N_2182,N_2191);
and U3796 (N_3796,N_2178,N_2935);
xor U3797 (N_3797,N_2274,N_2588);
nand U3798 (N_3798,N_2531,N_2788);
nor U3799 (N_3799,N_2405,N_2594);
and U3800 (N_3800,N_2407,N_2266);
or U3801 (N_3801,N_2242,N_2306);
xor U3802 (N_3802,N_2736,N_2744);
and U3803 (N_3803,N_2013,N_2986);
and U3804 (N_3804,N_2826,N_2345);
or U3805 (N_3805,N_2001,N_2592);
and U3806 (N_3806,N_2633,N_2901);
or U3807 (N_3807,N_2502,N_2542);
xor U3808 (N_3808,N_2498,N_2059);
or U3809 (N_3809,N_2055,N_2759);
nor U3810 (N_3810,N_2435,N_2965);
and U3811 (N_3811,N_2386,N_2105);
or U3812 (N_3812,N_2476,N_2250);
or U3813 (N_3813,N_2755,N_2942);
or U3814 (N_3814,N_2507,N_2839);
nand U3815 (N_3815,N_2181,N_2451);
nand U3816 (N_3816,N_2710,N_2759);
xnor U3817 (N_3817,N_2360,N_2560);
nand U3818 (N_3818,N_2352,N_2393);
nand U3819 (N_3819,N_2938,N_2776);
xor U3820 (N_3820,N_2933,N_2932);
xnor U3821 (N_3821,N_2979,N_2157);
nor U3822 (N_3822,N_2673,N_2903);
nor U3823 (N_3823,N_2881,N_2717);
and U3824 (N_3824,N_2943,N_2640);
and U3825 (N_3825,N_2242,N_2663);
nor U3826 (N_3826,N_2336,N_2801);
xor U3827 (N_3827,N_2409,N_2258);
and U3828 (N_3828,N_2641,N_2723);
and U3829 (N_3829,N_2700,N_2722);
nand U3830 (N_3830,N_2415,N_2840);
and U3831 (N_3831,N_2385,N_2532);
or U3832 (N_3832,N_2349,N_2679);
and U3833 (N_3833,N_2198,N_2560);
xor U3834 (N_3834,N_2804,N_2217);
or U3835 (N_3835,N_2108,N_2406);
xnor U3836 (N_3836,N_2802,N_2942);
and U3837 (N_3837,N_2134,N_2229);
and U3838 (N_3838,N_2941,N_2192);
nand U3839 (N_3839,N_2218,N_2887);
and U3840 (N_3840,N_2070,N_2405);
nor U3841 (N_3841,N_2810,N_2348);
nor U3842 (N_3842,N_2300,N_2917);
xor U3843 (N_3843,N_2296,N_2125);
or U3844 (N_3844,N_2253,N_2813);
nor U3845 (N_3845,N_2486,N_2432);
xor U3846 (N_3846,N_2625,N_2722);
nor U3847 (N_3847,N_2524,N_2351);
xnor U3848 (N_3848,N_2390,N_2091);
nand U3849 (N_3849,N_2630,N_2675);
nand U3850 (N_3850,N_2504,N_2130);
and U3851 (N_3851,N_2541,N_2013);
nor U3852 (N_3852,N_2798,N_2710);
and U3853 (N_3853,N_2833,N_2175);
nand U3854 (N_3854,N_2322,N_2286);
xnor U3855 (N_3855,N_2824,N_2694);
or U3856 (N_3856,N_2648,N_2300);
and U3857 (N_3857,N_2981,N_2947);
nor U3858 (N_3858,N_2112,N_2149);
xor U3859 (N_3859,N_2949,N_2870);
nor U3860 (N_3860,N_2931,N_2333);
nor U3861 (N_3861,N_2527,N_2289);
nor U3862 (N_3862,N_2285,N_2639);
xor U3863 (N_3863,N_2608,N_2349);
nand U3864 (N_3864,N_2546,N_2631);
nor U3865 (N_3865,N_2557,N_2579);
xor U3866 (N_3866,N_2611,N_2104);
and U3867 (N_3867,N_2816,N_2314);
xor U3868 (N_3868,N_2549,N_2830);
xor U3869 (N_3869,N_2407,N_2317);
and U3870 (N_3870,N_2876,N_2026);
xnor U3871 (N_3871,N_2873,N_2027);
or U3872 (N_3872,N_2916,N_2251);
and U3873 (N_3873,N_2810,N_2807);
nand U3874 (N_3874,N_2126,N_2520);
and U3875 (N_3875,N_2966,N_2279);
nor U3876 (N_3876,N_2696,N_2842);
or U3877 (N_3877,N_2313,N_2710);
or U3878 (N_3878,N_2044,N_2172);
xor U3879 (N_3879,N_2139,N_2545);
or U3880 (N_3880,N_2477,N_2888);
xor U3881 (N_3881,N_2933,N_2524);
or U3882 (N_3882,N_2220,N_2102);
and U3883 (N_3883,N_2945,N_2276);
nor U3884 (N_3884,N_2408,N_2315);
xor U3885 (N_3885,N_2885,N_2981);
or U3886 (N_3886,N_2187,N_2412);
nand U3887 (N_3887,N_2707,N_2340);
xnor U3888 (N_3888,N_2145,N_2656);
or U3889 (N_3889,N_2012,N_2064);
nor U3890 (N_3890,N_2295,N_2819);
xnor U3891 (N_3891,N_2033,N_2406);
nand U3892 (N_3892,N_2520,N_2778);
nor U3893 (N_3893,N_2399,N_2582);
nor U3894 (N_3894,N_2017,N_2574);
nand U3895 (N_3895,N_2931,N_2066);
or U3896 (N_3896,N_2449,N_2954);
nand U3897 (N_3897,N_2418,N_2563);
and U3898 (N_3898,N_2504,N_2693);
xnor U3899 (N_3899,N_2272,N_2234);
or U3900 (N_3900,N_2443,N_2080);
xnor U3901 (N_3901,N_2896,N_2359);
and U3902 (N_3902,N_2945,N_2764);
nand U3903 (N_3903,N_2085,N_2857);
and U3904 (N_3904,N_2191,N_2329);
nor U3905 (N_3905,N_2401,N_2126);
nor U3906 (N_3906,N_2208,N_2600);
xor U3907 (N_3907,N_2480,N_2943);
nand U3908 (N_3908,N_2881,N_2478);
and U3909 (N_3909,N_2136,N_2562);
nand U3910 (N_3910,N_2405,N_2734);
nand U3911 (N_3911,N_2117,N_2526);
nor U3912 (N_3912,N_2043,N_2059);
xor U3913 (N_3913,N_2001,N_2763);
or U3914 (N_3914,N_2686,N_2544);
xnor U3915 (N_3915,N_2830,N_2588);
xnor U3916 (N_3916,N_2671,N_2094);
xnor U3917 (N_3917,N_2315,N_2265);
or U3918 (N_3918,N_2877,N_2448);
xor U3919 (N_3919,N_2696,N_2840);
nor U3920 (N_3920,N_2285,N_2601);
nand U3921 (N_3921,N_2663,N_2067);
nand U3922 (N_3922,N_2714,N_2592);
nand U3923 (N_3923,N_2787,N_2829);
nor U3924 (N_3924,N_2364,N_2352);
nand U3925 (N_3925,N_2563,N_2207);
xnor U3926 (N_3926,N_2727,N_2488);
and U3927 (N_3927,N_2749,N_2778);
nand U3928 (N_3928,N_2952,N_2253);
and U3929 (N_3929,N_2800,N_2537);
xor U3930 (N_3930,N_2346,N_2191);
xnor U3931 (N_3931,N_2585,N_2427);
nor U3932 (N_3932,N_2320,N_2158);
nand U3933 (N_3933,N_2685,N_2188);
nor U3934 (N_3934,N_2038,N_2786);
nor U3935 (N_3935,N_2359,N_2053);
or U3936 (N_3936,N_2991,N_2686);
xnor U3937 (N_3937,N_2333,N_2977);
nand U3938 (N_3938,N_2286,N_2118);
or U3939 (N_3939,N_2092,N_2744);
xor U3940 (N_3940,N_2614,N_2475);
or U3941 (N_3941,N_2583,N_2745);
or U3942 (N_3942,N_2358,N_2226);
xnor U3943 (N_3943,N_2803,N_2732);
or U3944 (N_3944,N_2185,N_2998);
xnor U3945 (N_3945,N_2668,N_2459);
nand U3946 (N_3946,N_2587,N_2413);
nor U3947 (N_3947,N_2530,N_2930);
or U3948 (N_3948,N_2165,N_2318);
or U3949 (N_3949,N_2852,N_2643);
nand U3950 (N_3950,N_2208,N_2104);
or U3951 (N_3951,N_2837,N_2355);
and U3952 (N_3952,N_2466,N_2677);
nand U3953 (N_3953,N_2249,N_2068);
nor U3954 (N_3954,N_2474,N_2730);
or U3955 (N_3955,N_2737,N_2226);
or U3956 (N_3956,N_2943,N_2130);
or U3957 (N_3957,N_2782,N_2862);
xor U3958 (N_3958,N_2578,N_2647);
xor U3959 (N_3959,N_2694,N_2718);
nor U3960 (N_3960,N_2813,N_2295);
and U3961 (N_3961,N_2632,N_2436);
or U3962 (N_3962,N_2858,N_2813);
or U3963 (N_3963,N_2039,N_2366);
or U3964 (N_3964,N_2786,N_2084);
or U3965 (N_3965,N_2056,N_2907);
and U3966 (N_3966,N_2184,N_2124);
xor U3967 (N_3967,N_2836,N_2242);
xnor U3968 (N_3968,N_2540,N_2851);
and U3969 (N_3969,N_2443,N_2623);
xnor U3970 (N_3970,N_2978,N_2249);
nand U3971 (N_3971,N_2896,N_2046);
xnor U3972 (N_3972,N_2809,N_2750);
xnor U3973 (N_3973,N_2545,N_2526);
xor U3974 (N_3974,N_2065,N_2955);
nor U3975 (N_3975,N_2160,N_2520);
nand U3976 (N_3976,N_2039,N_2644);
nand U3977 (N_3977,N_2476,N_2502);
nand U3978 (N_3978,N_2055,N_2248);
xor U3979 (N_3979,N_2953,N_2291);
and U3980 (N_3980,N_2685,N_2371);
nand U3981 (N_3981,N_2862,N_2822);
xnor U3982 (N_3982,N_2835,N_2987);
and U3983 (N_3983,N_2538,N_2628);
nor U3984 (N_3984,N_2188,N_2702);
xor U3985 (N_3985,N_2216,N_2371);
or U3986 (N_3986,N_2355,N_2595);
or U3987 (N_3987,N_2406,N_2089);
and U3988 (N_3988,N_2062,N_2047);
xnor U3989 (N_3989,N_2783,N_2255);
or U3990 (N_3990,N_2866,N_2750);
nand U3991 (N_3991,N_2820,N_2721);
xnor U3992 (N_3992,N_2619,N_2699);
nand U3993 (N_3993,N_2745,N_2135);
xnor U3994 (N_3994,N_2460,N_2155);
xnor U3995 (N_3995,N_2722,N_2061);
nor U3996 (N_3996,N_2930,N_2146);
nor U3997 (N_3997,N_2922,N_2018);
nor U3998 (N_3998,N_2884,N_2293);
xor U3999 (N_3999,N_2518,N_2103);
xnor U4000 (N_4000,N_3188,N_3377);
nor U4001 (N_4001,N_3327,N_3579);
nor U4002 (N_4002,N_3111,N_3315);
nor U4003 (N_4003,N_3130,N_3737);
xor U4004 (N_4004,N_3128,N_3452);
or U4005 (N_4005,N_3797,N_3960);
or U4006 (N_4006,N_3904,N_3372);
or U4007 (N_4007,N_3056,N_3774);
nor U4008 (N_4008,N_3097,N_3385);
and U4009 (N_4009,N_3708,N_3662);
or U4010 (N_4010,N_3023,N_3608);
nand U4011 (N_4011,N_3302,N_3184);
or U4012 (N_4012,N_3927,N_3237);
and U4013 (N_4013,N_3576,N_3371);
nand U4014 (N_4014,N_3732,N_3709);
or U4015 (N_4015,N_3564,N_3101);
nor U4016 (N_4016,N_3654,N_3068);
nor U4017 (N_4017,N_3763,N_3031);
nor U4018 (N_4018,N_3383,N_3772);
nor U4019 (N_4019,N_3355,N_3767);
and U4020 (N_4020,N_3214,N_3690);
and U4021 (N_4021,N_3856,N_3438);
and U4022 (N_4022,N_3581,N_3081);
or U4023 (N_4023,N_3061,N_3476);
nand U4024 (N_4024,N_3403,N_3706);
and U4025 (N_4025,N_3109,N_3332);
nor U4026 (N_4026,N_3588,N_3011);
nand U4027 (N_4027,N_3387,N_3122);
xnor U4028 (N_4028,N_3168,N_3057);
and U4029 (N_4029,N_3202,N_3733);
nand U4030 (N_4030,N_3847,N_3508);
xnor U4031 (N_4031,N_3672,N_3204);
or U4032 (N_4032,N_3651,N_3653);
or U4033 (N_4033,N_3486,N_3255);
nor U4034 (N_4034,N_3765,N_3421);
nand U4035 (N_4035,N_3400,N_3726);
or U4036 (N_4036,N_3284,N_3343);
and U4037 (N_4037,N_3933,N_3474);
nand U4038 (N_4038,N_3936,N_3816);
and U4039 (N_4039,N_3905,N_3412);
nor U4040 (N_4040,N_3379,N_3034);
nand U4041 (N_4041,N_3606,N_3923);
nor U4042 (N_4042,N_3234,N_3192);
nor U4043 (N_4043,N_3578,N_3630);
or U4044 (N_4044,N_3511,N_3657);
and U4045 (N_4045,N_3752,N_3791);
nand U4046 (N_4046,N_3271,N_3328);
nand U4047 (N_4047,N_3118,N_3558);
nand U4048 (N_4048,N_3718,N_3829);
and U4049 (N_4049,N_3038,N_3303);
nand U4050 (N_4050,N_3992,N_3570);
xnor U4051 (N_4051,N_3205,N_3543);
and U4052 (N_4052,N_3523,N_3824);
or U4053 (N_4053,N_3888,N_3766);
xnor U4054 (N_4054,N_3203,N_3822);
and U4055 (N_4055,N_3114,N_3650);
nor U4056 (N_4056,N_3841,N_3739);
xnor U4057 (N_4057,N_3195,N_3404);
nand U4058 (N_4058,N_3585,N_3321);
xor U4059 (N_4059,N_3861,N_3643);
xnor U4060 (N_4060,N_3903,N_3539);
xor U4061 (N_4061,N_3574,N_3288);
or U4062 (N_4062,N_3730,N_3674);
and U4063 (N_4063,N_3591,N_3849);
or U4064 (N_4064,N_3838,N_3487);
nand U4065 (N_4065,N_3047,N_3125);
and U4066 (N_4066,N_3713,N_3595);
xor U4067 (N_4067,N_3473,N_3792);
nor U4068 (N_4068,N_3957,N_3796);
or U4069 (N_4069,N_3425,N_3871);
or U4070 (N_4070,N_3568,N_3013);
or U4071 (N_4071,N_3863,N_3663);
or U4072 (N_4072,N_3206,N_3330);
or U4073 (N_4073,N_3020,N_3700);
xnor U4074 (N_4074,N_3189,N_3333);
nand U4075 (N_4075,N_3426,N_3370);
xor U4076 (N_4076,N_3885,N_3670);
xnor U4077 (N_4077,N_3883,N_3074);
or U4078 (N_4078,N_3449,N_3457);
or U4079 (N_4079,N_3405,N_3665);
or U4080 (N_4080,N_3201,N_3605);
and U4081 (N_4081,N_3500,N_3235);
nand U4082 (N_4082,N_3433,N_3819);
nor U4083 (N_4083,N_3785,N_3636);
nor U4084 (N_4084,N_3602,N_3496);
or U4085 (N_4085,N_3021,N_3534);
xor U4086 (N_4086,N_3414,N_3399);
xor U4087 (N_4087,N_3624,N_3832);
or U4088 (N_4088,N_3760,N_3795);
xor U4089 (N_4089,N_3979,N_3880);
and U4090 (N_4090,N_3300,N_3734);
and U4091 (N_4091,N_3363,N_3727);
or U4092 (N_4092,N_3517,N_3912);
nand U4093 (N_4093,N_3768,N_3478);
nand U4094 (N_4094,N_3601,N_3095);
and U4095 (N_4095,N_3186,N_3617);
nand U4096 (N_4096,N_3563,N_3275);
xnor U4097 (N_4097,N_3108,N_3480);
nand U4098 (N_4098,N_3194,N_3110);
nor U4099 (N_4099,N_3398,N_3779);
nor U4100 (N_4100,N_3093,N_3169);
or U4101 (N_4101,N_3900,N_3054);
and U4102 (N_4102,N_3217,N_3806);
nand U4103 (N_4103,N_3682,N_3924);
nand U4104 (N_4104,N_3603,N_3975);
xor U4105 (N_4105,N_3022,N_3859);
xnor U4106 (N_4106,N_3540,N_3462);
nor U4107 (N_4107,N_3661,N_3287);
nor U4108 (N_4108,N_3466,N_3085);
and U4109 (N_4109,N_3613,N_3741);
xor U4110 (N_4110,N_3943,N_3036);
nor U4111 (N_4111,N_3515,N_3973);
and U4112 (N_4112,N_3178,N_3472);
nand U4113 (N_4113,N_3254,N_3917);
nand U4114 (N_4114,N_3974,N_3628);
and U4115 (N_4115,N_3793,N_3269);
and U4116 (N_4116,N_3535,N_3882);
nor U4117 (N_4117,N_3475,N_3876);
nand U4118 (N_4118,N_3483,N_3182);
nand U4119 (N_4119,N_3711,N_3986);
nor U4120 (N_4120,N_3375,N_3867);
and U4121 (N_4121,N_3348,N_3001);
and U4122 (N_4122,N_3507,N_3629);
xor U4123 (N_4123,N_3828,N_3865);
xor U4124 (N_4124,N_3135,N_3158);
nand U4125 (N_4125,N_3018,N_3336);
and U4126 (N_4126,N_3308,N_3143);
xor U4127 (N_4127,N_3609,N_3502);
and U4128 (N_4128,N_3889,N_3073);
and U4129 (N_4129,N_3304,N_3589);
and U4130 (N_4130,N_3921,N_3103);
or U4131 (N_4131,N_3864,N_3415);
xnor U4132 (N_4132,N_3391,N_3848);
xor U4133 (N_4133,N_3692,N_3242);
xnor U4134 (N_4134,N_3228,N_3075);
nor U4135 (N_4135,N_3631,N_3513);
and U4136 (N_4136,N_3544,N_3712);
or U4137 (N_4137,N_3744,N_3685);
nor U4138 (N_4138,N_3116,N_3091);
xnor U4139 (N_4139,N_3582,N_3612);
nor U4140 (N_4140,N_3440,N_3639);
or U4141 (N_4141,N_3532,N_3625);
nor U4142 (N_4142,N_3407,N_3925);
or U4143 (N_4143,N_3311,N_3614);
xor U4144 (N_4144,N_3196,N_3148);
or U4145 (N_4145,N_3331,N_3364);
and U4146 (N_4146,N_3185,N_3788);
xnor U4147 (N_4147,N_3469,N_3538);
or U4148 (N_4148,N_3843,N_3419);
xnor U4149 (N_4149,N_3362,N_3964);
xor U4150 (N_4150,N_3821,N_3569);
or U4151 (N_4151,N_3003,N_3839);
nor U4152 (N_4152,N_3669,N_3659);
xnor U4153 (N_4153,N_3257,N_3225);
or U4154 (N_4154,N_3504,N_3326);
xor U4155 (N_4155,N_3174,N_3844);
and U4156 (N_4156,N_3147,N_3969);
xnor U4157 (N_4157,N_3455,N_3928);
nand U4158 (N_4158,N_3716,N_3586);
and U4159 (N_4159,N_3966,N_3278);
nand U4160 (N_4160,N_3955,N_3159);
or U4161 (N_4161,N_3980,N_3037);
xor U4162 (N_4162,N_3113,N_3567);
and U4163 (N_4163,N_3120,N_3318);
xor U4164 (N_4164,N_3063,N_3825);
and U4165 (N_4165,N_3707,N_3655);
nand U4166 (N_4166,N_3067,N_3297);
and U4167 (N_4167,N_3157,N_3584);
xnor U4168 (N_4168,N_3347,N_3571);
and U4169 (N_4169,N_3922,N_3319);
xor U4170 (N_4170,N_3748,N_3627);
nor U4171 (N_4171,N_3557,N_3649);
and U4172 (N_4172,N_3820,N_3491);
xnor U4173 (N_4173,N_3423,N_3488);
and U4174 (N_4174,N_3547,N_3619);
nand U4175 (N_4175,N_3626,N_3256);
nand U4176 (N_4176,N_3652,N_3906);
nor U4177 (N_4177,N_3593,N_3698);
and U4178 (N_4178,N_3349,N_3756);
nand U4179 (N_4179,N_3002,N_3525);
xnor U4180 (N_4180,N_3673,N_3758);
or U4181 (N_4181,N_3528,N_3155);
nand U4182 (N_4182,N_3124,N_3675);
and U4183 (N_4183,N_3874,N_3990);
nor U4184 (N_4184,N_3080,N_3681);
nand U4185 (N_4185,N_3641,N_3505);
xnor U4186 (N_4186,N_3594,N_3704);
and U4187 (N_4187,N_3961,N_3325);
or U4188 (N_4188,N_3648,N_3434);
nor U4189 (N_4189,N_3810,N_3167);
or U4190 (N_4190,N_3890,N_3334);
nand U4191 (N_4191,N_3140,N_3222);
xor U4192 (N_4192,N_3241,N_3866);
nand U4193 (N_4193,N_3913,N_3039);
and U4194 (N_4194,N_3417,N_3647);
or U4195 (N_4195,N_3358,N_3497);
xor U4196 (N_4196,N_3944,N_3230);
nand U4197 (N_4197,N_3406,N_3644);
and U4198 (N_4198,N_3947,N_3549);
or U4199 (N_4199,N_3268,N_3247);
xor U4200 (N_4200,N_3703,N_3436);
xor U4201 (N_4201,N_3747,N_3294);
xor U4202 (N_4202,N_3658,N_3069);
nor U4203 (N_4203,N_3811,N_3954);
nand U4204 (N_4204,N_3762,N_3459);
nand U4205 (N_4205,N_3381,N_3561);
nand U4206 (N_4206,N_3442,N_3243);
or U4207 (N_4207,N_3410,N_3799);
or U4208 (N_4208,N_3723,N_3019);
nand U4209 (N_4209,N_3179,N_3078);
nor U4210 (N_4210,N_3123,N_3632);
and U4211 (N_4211,N_3076,N_3276);
nand U4212 (N_4212,N_3397,N_3615);
and U4213 (N_4213,N_3695,N_3638);
nor U4214 (N_4214,N_3531,N_3295);
and U4215 (N_4215,N_3025,N_3133);
nor U4216 (N_4216,N_3886,N_3060);
nand U4217 (N_4217,N_3721,N_3753);
nand U4218 (N_4218,N_3260,N_3320);
nor U4219 (N_4219,N_3006,N_3934);
nand U4220 (N_4220,N_3281,N_3450);
and U4221 (N_4221,N_3445,N_3142);
or U4222 (N_4222,N_3131,N_3552);
nor U4223 (N_4223,N_3117,N_3079);
and U4224 (N_4224,N_3596,N_3317);
nor U4225 (N_4225,N_3224,N_3240);
or U4226 (N_4226,N_3845,N_3495);
or U4227 (N_4227,N_3746,N_3789);
nor U4228 (N_4228,N_3471,N_3621);
xor U4229 (N_4229,N_3136,N_3312);
nand U4230 (N_4230,N_3678,N_3577);
nor U4231 (N_4231,N_3524,N_3066);
nor U4232 (N_4232,N_3164,N_3967);
nand U4233 (N_4233,N_3982,N_3181);
xnor U4234 (N_4234,N_3958,N_3464);
xnor U4235 (N_4235,N_3051,N_3467);
nand U4236 (N_4236,N_3378,N_3094);
nand U4237 (N_4237,N_3951,N_3351);
nor U4238 (N_4238,N_3842,N_3714);
nand U4239 (N_4239,N_3916,N_3808);
or U4240 (N_4240,N_3431,N_3520);
nand U4241 (N_4241,N_3139,N_3545);
or U4242 (N_4242,N_3536,N_3761);
nand U4243 (N_4243,N_3088,N_3899);
xor U4244 (N_4244,N_3699,N_3441);
or U4245 (N_4245,N_3776,N_3740);
xor U4246 (N_4246,N_3033,N_3770);
and U4247 (N_4247,N_3893,N_3942);
and U4248 (N_4248,N_3468,N_3562);
or U4249 (N_4249,N_3996,N_3245);
or U4250 (N_4250,N_3059,N_3213);
and U4251 (N_4251,N_3719,N_3233);
or U4252 (N_4252,N_3171,N_3454);
or U4253 (N_4253,N_3447,N_3800);
nor U4254 (N_4254,N_3679,N_3301);
xor U4255 (N_4255,N_3878,N_3208);
xnor U4256 (N_4256,N_3306,N_3231);
xor U4257 (N_4257,N_3892,N_3283);
xnor U4258 (N_4258,N_3046,N_3162);
nand U4259 (N_4259,N_3107,N_3742);
or U4260 (N_4260,N_3263,N_3451);
nand U4261 (N_4261,N_3322,N_3901);
xnor U4262 (N_4262,N_3052,N_3989);
xor U4263 (N_4263,N_3573,N_3814);
and U4264 (N_4264,N_3512,N_3553);
nor U4265 (N_4265,N_3161,N_3154);
or U4266 (N_4266,N_3953,N_3620);
xor U4267 (N_4267,N_3070,N_3548);
xor U4268 (N_4268,N_3494,N_3705);
or U4269 (N_4269,N_3015,N_3757);
or U4270 (N_4270,N_3367,N_3755);
or U4271 (N_4271,N_3272,N_3938);
nor U4272 (N_4272,N_3857,N_3823);
and U4273 (N_4273,N_3422,N_3945);
nand U4274 (N_4274,N_3198,N_3492);
xor U4275 (N_4275,N_3401,N_3265);
nand U4276 (N_4276,N_3702,N_3514);
nand U4277 (N_4277,N_3005,N_3259);
or U4278 (N_4278,N_3583,N_3873);
nor U4279 (N_4279,N_3600,N_3219);
or U4280 (N_4280,N_3394,N_3929);
nor U4281 (N_4281,N_3007,N_3868);
xor U4282 (N_4282,N_3270,N_3743);
nor U4283 (N_4283,N_3884,N_3910);
nand U4284 (N_4284,N_3780,N_3777);
and U4285 (N_4285,N_3072,N_3566);
or U4286 (N_4286,N_3926,N_3671);
xnor U4287 (N_4287,N_3855,N_3250);
xnor U4288 (N_4288,N_3369,N_3009);
or U4289 (N_4289,N_3754,N_3759);
and U4290 (N_4290,N_3533,N_3935);
nand U4291 (N_4291,N_3931,N_3813);
xnor U4292 (N_4292,N_3470,N_3830);
xor U4293 (N_4293,N_3251,N_3526);
or U4294 (N_4294,N_3994,N_3817);
or U4295 (N_4295,N_3798,N_3869);
nand U4296 (N_4296,N_3146,N_3309);
nand U4297 (N_4297,N_3127,N_3914);
nor U4298 (N_4298,N_3227,N_3911);
and U4299 (N_4299,N_3115,N_3106);
xor U4300 (N_4300,N_3393,N_3339);
and U4301 (N_4301,N_3390,N_3238);
and U4302 (N_4302,N_3887,N_3597);
xnor U4303 (N_4303,N_3190,N_3216);
nand U4304 (N_4304,N_3053,N_3236);
nand U4305 (N_4305,N_3771,N_3396);
nor U4306 (N_4306,N_3664,N_3968);
and U4307 (N_4307,N_3463,N_3645);
or U4308 (N_4308,N_3092,N_3411);
and U4309 (N_4309,N_3801,N_3089);
or U4310 (N_4310,N_3293,N_3720);
and U4311 (N_4311,N_3546,N_3805);
and U4312 (N_4312,N_3481,N_3909);
nor U4313 (N_4313,N_3689,N_3556);
or U4314 (N_4314,N_3999,N_3684);
nand U4315 (N_4315,N_3361,N_3342);
and U4316 (N_4316,N_3199,N_3879);
xor U4317 (N_4317,N_3853,N_3151);
nor U4318 (N_4318,N_3490,N_3289);
xor U4319 (N_4319,N_3919,N_3950);
nand U4320 (N_4320,N_3359,N_3509);
nor U4321 (N_4321,N_3728,N_3750);
and U4322 (N_4322,N_3144,N_3280);
nor U4323 (N_4323,N_3872,N_3338);
xnor U4324 (N_4324,N_3939,N_3498);
or U4325 (N_4325,N_3170,N_3392);
xor U4326 (N_4326,N_3261,N_3200);
nand U4327 (N_4327,N_3432,N_3232);
or U4328 (N_4328,N_3940,N_3668);
and U4329 (N_4329,N_3086,N_3132);
and U4330 (N_4330,N_3058,N_3465);
nor U4331 (N_4331,N_3489,N_3197);
xor U4332 (N_4332,N_3368,N_3995);
or U4333 (N_4333,N_3587,N_3292);
or U4334 (N_4334,N_3266,N_3264);
nand U4335 (N_4335,N_3177,N_3745);
or U4336 (N_4336,N_3042,N_3380);
nand U4337 (N_4337,N_3896,N_3781);
and U4338 (N_4338,N_3435,N_3282);
nor U4339 (N_4339,N_3693,N_3316);
or U4340 (N_4340,N_3104,N_3854);
or U4341 (N_4341,N_3642,N_3794);
nand U4342 (N_4342,N_3071,N_3701);
nor U4343 (N_4343,N_3386,N_3460);
or U4344 (N_4344,N_3376,N_3444);
xor U4345 (N_4345,N_3965,N_3035);
and U4346 (N_4346,N_3418,N_3804);
and U4347 (N_4347,N_3365,N_3751);
or U4348 (N_4348,N_3787,N_3784);
and U4349 (N_4349,N_3834,N_3313);
xnor U4350 (N_4350,N_3337,N_3898);
nand U4351 (N_4351,N_3191,N_3166);
or U4352 (N_4352,N_3895,N_3152);
or U4353 (N_4353,N_3027,N_3604);
nor U4354 (N_4354,N_3519,N_3985);
nand U4355 (N_4355,N_3978,N_3946);
or U4356 (N_4356,N_3004,N_3290);
or U4357 (N_4357,N_3000,N_3790);
and U4358 (N_4358,N_3215,N_3599);
nand U4359 (N_4359,N_3307,N_3738);
and U4360 (N_4360,N_3984,N_3150);
nand U4361 (N_4361,N_3437,N_3724);
nand U4362 (N_4362,N_3687,N_3062);
xor U4363 (N_4363,N_3439,N_3518);
and U4364 (N_4364,N_3948,N_3623);
nor U4365 (N_4365,N_3993,N_3285);
xnor U4366 (N_4366,N_3485,N_3356);
and U4367 (N_4367,N_3012,N_3210);
xnor U4368 (N_4368,N_3962,N_3350);
or U4369 (N_4369,N_3725,N_3346);
nand U4370 (N_4370,N_3640,N_3949);
nor U4371 (N_4371,N_3897,N_3807);
or U4372 (N_4372,N_3611,N_3050);
and U4373 (N_4373,N_3851,N_3860);
and U4374 (N_4374,N_3778,N_3024);
and U4375 (N_4375,N_3384,N_3501);
xor U4376 (N_4376,N_3055,N_3598);
nand U4377 (N_4377,N_3622,N_3881);
and U4378 (N_4378,N_3428,N_3134);
xor U4379 (N_4379,N_3683,N_3244);
nand U4380 (N_4380,N_3160,N_3279);
nand U4381 (N_4381,N_3017,N_3510);
and U4382 (N_4382,N_3920,N_3722);
nor U4383 (N_4383,N_3030,N_3220);
nor U4384 (N_4384,N_3360,N_3026);
and U4385 (N_4385,N_3082,N_3484);
or U4386 (N_4386,N_3499,N_3352);
nand U4387 (N_4387,N_3542,N_3559);
and U4388 (N_4388,N_3660,N_3065);
and U4389 (N_4389,N_3530,N_3666);
nor U4390 (N_4390,N_3987,N_3087);
nor U4391 (N_4391,N_3456,N_3835);
and U4392 (N_4392,N_3262,N_3218);
nand U4393 (N_4393,N_3555,N_3831);
or U4394 (N_4394,N_3253,N_3008);
nor U4395 (N_4395,N_3239,N_3341);
nand U4396 (N_4396,N_3374,N_3983);
xor U4397 (N_4397,N_3153,N_3044);
and U4398 (N_4398,N_3918,N_3782);
xnor U4399 (N_4399,N_3448,N_3775);
or U4400 (N_4400,N_3852,N_3691);
or U4401 (N_4401,N_3105,N_3715);
nand U4402 (N_4402,N_3634,N_3329);
nand U4403 (N_4403,N_3267,N_3305);
and U4404 (N_4404,N_3930,N_3633);
nand U4405 (N_4405,N_3064,N_3014);
xnor U4406 (N_4406,N_3656,N_3956);
nand U4407 (N_4407,N_3894,N_3100);
or U4408 (N_4408,N_3430,N_3786);
or U4409 (N_4409,N_3077,N_3667);
nor U4410 (N_4410,N_3453,N_3837);
xor U4411 (N_4411,N_3827,N_3090);
nor U4412 (N_4412,N_3163,N_3902);
or U4413 (N_4413,N_3972,N_3032);
xnor U4414 (N_4414,N_3096,N_3248);
nand U4415 (N_4415,N_3731,N_3610);
xnor U4416 (N_4416,N_3183,N_3043);
or U4417 (N_4417,N_3221,N_3840);
and U4418 (N_4418,N_3694,N_3395);
xnor U4419 (N_4419,N_3353,N_3141);
xnor U4420 (N_4420,N_3565,N_3335);
nand U4421 (N_4421,N_3382,N_3677);
nand U4422 (N_4422,N_3408,N_3029);
and U4423 (N_4423,N_3479,N_3314);
nor U4424 (N_4424,N_3907,N_3298);
or U4425 (N_4425,N_3915,N_3710);
and U4426 (N_4426,N_3818,N_3932);
nand U4427 (N_4427,N_3207,N_3554);
or U4428 (N_4428,N_3482,N_3252);
nor U4429 (N_4429,N_3580,N_3991);
nand U4430 (N_4430,N_3646,N_3413);
nor U4431 (N_4431,N_3815,N_3461);
and U4432 (N_4432,N_3175,N_3420);
and U4433 (N_4433,N_3875,N_3340);
nor U4434 (N_4434,N_3998,N_3607);
xnor U4435 (N_4435,N_3416,N_3697);
nor U4436 (N_4436,N_3084,N_3572);
or U4437 (N_4437,N_3590,N_3310);
xor U4438 (N_4438,N_3028,N_3041);
nor U4439 (N_4439,N_3212,N_3246);
or U4440 (N_4440,N_3971,N_3209);
and U4441 (N_4441,N_3959,N_3736);
nor U4442 (N_4442,N_3145,N_3891);
nand U4443 (N_4443,N_3126,N_3809);
xor U4444 (N_4444,N_3870,N_3592);
or U4445 (N_4445,N_3193,N_3286);
and U4446 (N_4446,N_3354,N_3223);
nand U4447 (N_4447,N_3119,N_3345);
xor U4448 (N_4448,N_3635,N_3970);
nand U4449 (N_4449,N_3291,N_3048);
nor U4450 (N_4450,N_3226,N_3783);
nand U4451 (N_4451,N_3997,N_3537);
and U4452 (N_4452,N_3560,N_3229);
xnor U4453 (N_4453,N_3862,N_3616);
xnor U4454 (N_4454,N_3098,N_3812);
or U4455 (N_4455,N_3274,N_3149);
and U4456 (N_4456,N_3258,N_3156);
or U4457 (N_4457,N_3366,N_3172);
xor U4458 (N_4458,N_3541,N_3388);
xor U4459 (N_4459,N_3802,N_3686);
nor U4460 (N_4460,N_3049,N_3173);
xor U4461 (N_4461,N_3273,N_3099);
nand U4462 (N_4462,N_3402,N_3277);
nor U4463 (N_4463,N_3764,N_3112);
and U4464 (N_4464,N_3696,N_3424);
nand U4465 (N_4465,N_3083,N_3010);
and U4466 (N_4466,N_3516,N_3323);
nand U4467 (N_4467,N_3981,N_3680);
and U4468 (N_4468,N_3550,N_3551);
nor U4469 (N_4469,N_3211,N_3102);
and U4470 (N_4470,N_3249,N_3522);
or U4471 (N_4471,N_3937,N_3129);
and U4472 (N_4472,N_3908,N_3803);
xor U4473 (N_4473,N_3846,N_3040);
or U4474 (N_4474,N_3688,N_3324);
or U4475 (N_4475,N_3717,N_3344);
or U4476 (N_4476,N_3296,N_3503);
or U4477 (N_4477,N_3575,N_3833);
xor U4478 (N_4478,N_3121,N_3187);
or U4479 (N_4479,N_3165,N_3976);
nand U4480 (N_4480,N_3138,N_3637);
nor U4481 (N_4481,N_3977,N_3521);
or U4482 (N_4482,N_3850,N_3527);
nor U4483 (N_4483,N_3443,N_3773);
nand U4484 (N_4484,N_3877,N_3180);
nand U4485 (N_4485,N_3373,N_3458);
nor U4486 (N_4486,N_3618,N_3858);
or U4487 (N_4487,N_3137,N_3735);
nand U4488 (N_4488,N_3529,N_3446);
or U4489 (N_4489,N_3836,N_3477);
nor U4490 (N_4490,N_3749,N_3409);
and U4491 (N_4491,N_3729,N_3299);
and U4492 (N_4492,N_3826,N_3357);
nand U4493 (N_4493,N_3769,N_3493);
nand U4494 (N_4494,N_3952,N_3988);
nor U4495 (N_4495,N_3506,N_3427);
nand U4496 (N_4496,N_3389,N_3941);
and U4497 (N_4497,N_3016,N_3429);
or U4498 (N_4498,N_3045,N_3676);
nor U4499 (N_4499,N_3176,N_3963);
nand U4500 (N_4500,N_3141,N_3079);
nor U4501 (N_4501,N_3256,N_3038);
xor U4502 (N_4502,N_3250,N_3835);
or U4503 (N_4503,N_3758,N_3843);
or U4504 (N_4504,N_3830,N_3215);
nor U4505 (N_4505,N_3035,N_3558);
nand U4506 (N_4506,N_3257,N_3747);
nand U4507 (N_4507,N_3134,N_3065);
or U4508 (N_4508,N_3685,N_3740);
xnor U4509 (N_4509,N_3990,N_3326);
nand U4510 (N_4510,N_3688,N_3468);
nand U4511 (N_4511,N_3283,N_3327);
and U4512 (N_4512,N_3701,N_3074);
xor U4513 (N_4513,N_3060,N_3992);
and U4514 (N_4514,N_3525,N_3265);
and U4515 (N_4515,N_3380,N_3861);
and U4516 (N_4516,N_3811,N_3894);
nand U4517 (N_4517,N_3828,N_3622);
and U4518 (N_4518,N_3546,N_3522);
or U4519 (N_4519,N_3081,N_3208);
or U4520 (N_4520,N_3315,N_3873);
nor U4521 (N_4521,N_3835,N_3514);
nand U4522 (N_4522,N_3520,N_3440);
and U4523 (N_4523,N_3756,N_3834);
or U4524 (N_4524,N_3571,N_3443);
xnor U4525 (N_4525,N_3190,N_3205);
xor U4526 (N_4526,N_3699,N_3976);
nor U4527 (N_4527,N_3794,N_3317);
nor U4528 (N_4528,N_3966,N_3472);
or U4529 (N_4529,N_3122,N_3252);
xnor U4530 (N_4530,N_3869,N_3679);
or U4531 (N_4531,N_3562,N_3407);
nand U4532 (N_4532,N_3439,N_3692);
xor U4533 (N_4533,N_3622,N_3533);
nand U4534 (N_4534,N_3470,N_3213);
nand U4535 (N_4535,N_3396,N_3114);
nand U4536 (N_4536,N_3864,N_3565);
xor U4537 (N_4537,N_3548,N_3735);
xor U4538 (N_4538,N_3443,N_3341);
nand U4539 (N_4539,N_3702,N_3637);
nand U4540 (N_4540,N_3872,N_3258);
xor U4541 (N_4541,N_3476,N_3121);
nor U4542 (N_4542,N_3565,N_3603);
xnor U4543 (N_4543,N_3754,N_3350);
nor U4544 (N_4544,N_3722,N_3746);
nand U4545 (N_4545,N_3781,N_3530);
nand U4546 (N_4546,N_3868,N_3134);
nand U4547 (N_4547,N_3231,N_3516);
nor U4548 (N_4548,N_3127,N_3347);
xor U4549 (N_4549,N_3425,N_3328);
and U4550 (N_4550,N_3135,N_3526);
xnor U4551 (N_4551,N_3341,N_3092);
xnor U4552 (N_4552,N_3797,N_3609);
nand U4553 (N_4553,N_3165,N_3496);
nor U4554 (N_4554,N_3928,N_3199);
or U4555 (N_4555,N_3982,N_3878);
xnor U4556 (N_4556,N_3720,N_3746);
or U4557 (N_4557,N_3502,N_3285);
nand U4558 (N_4558,N_3093,N_3392);
and U4559 (N_4559,N_3867,N_3663);
and U4560 (N_4560,N_3252,N_3085);
and U4561 (N_4561,N_3151,N_3251);
and U4562 (N_4562,N_3610,N_3443);
and U4563 (N_4563,N_3934,N_3064);
xor U4564 (N_4564,N_3950,N_3050);
nand U4565 (N_4565,N_3312,N_3414);
nand U4566 (N_4566,N_3636,N_3185);
or U4567 (N_4567,N_3855,N_3436);
and U4568 (N_4568,N_3795,N_3622);
xor U4569 (N_4569,N_3779,N_3129);
nor U4570 (N_4570,N_3192,N_3670);
nand U4571 (N_4571,N_3531,N_3046);
xnor U4572 (N_4572,N_3922,N_3978);
xnor U4573 (N_4573,N_3838,N_3868);
or U4574 (N_4574,N_3673,N_3802);
or U4575 (N_4575,N_3854,N_3663);
nand U4576 (N_4576,N_3599,N_3669);
or U4577 (N_4577,N_3861,N_3482);
or U4578 (N_4578,N_3947,N_3014);
nor U4579 (N_4579,N_3340,N_3822);
or U4580 (N_4580,N_3236,N_3010);
and U4581 (N_4581,N_3553,N_3256);
nor U4582 (N_4582,N_3553,N_3363);
xor U4583 (N_4583,N_3537,N_3293);
nor U4584 (N_4584,N_3923,N_3199);
and U4585 (N_4585,N_3451,N_3436);
nor U4586 (N_4586,N_3588,N_3585);
or U4587 (N_4587,N_3059,N_3561);
nor U4588 (N_4588,N_3125,N_3038);
nand U4589 (N_4589,N_3353,N_3473);
xor U4590 (N_4590,N_3516,N_3096);
xor U4591 (N_4591,N_3364,N_3010);
nor U4592 (N_4592,N_3845,N_3865);
and U4593 (N_4593,N_3839,N_3817);
nand U4594 (N_4594,N_3988,N_3989);
nand U4595 (N_4595,N_3151,N_3028);
nand U4596 (N_4596,N_3336,N_3406);
xor U4597 (N_4597,N_3139,N_3674);
and U4598 (N_4598,N_3520,N_3252);
nand U4599 (N_4599,N_3170,N_3029);
xor U4600 (N_4600,N_3574,N_3666);
and U4601 (N_4601,N_3349,N_3217);
xnor U4602 (N_4602,N_3920,N_3192);
xor U4603 (N_4603,N_3258,N_3765);
or U4604 (N_4604,N_3153,N_3282);
nand U4605 (N_4605,N_3325,N_3198);
or U4606 (N_4606,N_3650,N_3613);
xor U4607 (N_4607,N_3252,N_3917);
xnor U4608 (N_4608,N_3851,N_3733);
and U4609 (N_4609,N_3825,N_3680);
or U4610 (N_4610,N_3473,N_3999);
nand U4611 (N_4611,N_3791,N_3392);
or U4612 (N_4612,N_3218,N_3027);
nor U4613 (N_4613,N_3755,N_3270);
nor U4614 (N_4614,N_3906,N_3766);
and U4615 (N_4615,N_3253,N_3981);
nand U4616 (N_4616,N_3749,N_3765);
nand U4617 (N_4617,N_3990,N_3205);
and U4618 (N_4618,N_3381,N_3565);
or U4619 (N_4619,N_3629,N_3386);
or U4620 (N_4620,N_3858,N_3074);
nand U4621 (N_4621,N_3351,N_3833);
nor U4622 (N_4622,N_3763,N_3678);
xnor U4623 (N_4623,N_3071,N_3121);
or U4624 (N_4624,N_3035,N_3458);
and U4625 (N_4625,N_3851,N_3964);
nand U4626 (N_4626,N_3620,N_3569);
or U4627 (N_4627,N_3083,N_3411);
nor U4628 (N_4628,N_3840,N_3815);
nor U4629 (N_4629,N_3630,N_3444);
nand U4630 (N_4630,N_3779,N_3791);
and U4631 (N_4631,N_3600,N_3977);
and U4632 (N_4632,N_3990,N_3604);
nand U4633 (N_4633,N_3867,N_3021);
nand U4634 (N_4634,N_3531,N_3581);
and U4635 (N_4635,N_3943,N_3062);
nor U4636 (N_4636,N_3389,N_3163);
or U4637 (N_4637,N_3698,N_3127);
nand U4638 (N_4638,N_3014,N_3687);
xor U4639 (N_4639,N_3845,N_3012);
nor U4640 (N_4640,N_3722,N_3022);
nor U4641 (N_4641,N_3936,N_3931);
or U4642 (N_4642,N_3186,N_3005);
and U4643 (N_4643,N_3314,N_3339);
or U4644 (N_4644,N_3846,N_3253);
nand U4645 (N_4645,N_3644,N_3363);
or U4646 (N_4646,N_3254,N_3769);
or U4647 (N_4647,N_3369,N_3324);
or U4648 (N_4648,N_3431,N_3774);
nand U4649 (N_4649,N_3233,N_3514);
nand U4650 (N_4650,N_3807,N_3564);
nand U4651 (N_4651,N_3292,N_3637);
or U4652 (N_4652,N_3779,N_3783);
xnor U4653 (N_4653,N_3882,N_3689);
xor U4654 (N_4654,N_3926,N_3068);
xor U4655 (N_4655,N_3054,N_3379);
nor U4656 (N_4656,N_3331,N_3170);
nand U4657 (N_4657,N_3512,N_3562);
nor U4658 (N_4658,N_3032,N_3735);
nor U4659 (N_4659,N_3218,N_3064);
or U4660 (N_4660,N_3722,N_3366);
nor U4661 (N_4661,N_3908,N_3448);
or U4662 (N_4662,N_3123,N_3948);
nor U4663 (N_4663,N_3960,N_3907);
nand U4664 (N_4664,N_3895,N_3147);
xnor U4665 (N_4665,N_3286,N_3160);
and U4666 (N_4666,N_3577,N_3371);
or U4667 (N_4667,N_3503,N_3419);
xnor U4668 (N_4668,N_3600,N_3648);
or U4669 (N_4669,N_3802,N_3780);
nand U4670 (N_4670,N_3564,N_3941);
nor U4671 (N_4671,N_3205,N_3232);
xnor U4672 (N_4672,N_3750,N_3212);
or U4673 (N_4673,N_3522,N_3211);
nor U4674 (N_4674,N_3072,N_3724);
xor U4675 (N_4675,N_3648,N_3577);
nand U4676 (N_4676,N_3806,N_3718);
nor U4677 (N_4677,N_3123,N_3159);
or U4678 (N_4678,N_3657,N_3736);
nor U4679 (N_4679,N_3488,N_3174);
and U4680 (N_4680,N_3150,N_3252);
xor U4681 (N_4681,N_3441,N_3957);
nor U4682 (N_4682,N_3902,N_3127);
or U4683 (N_4683,N_3387,N_3251);
and U4684 (N_4684,N_3264,N_3023);
nand U4685 (N_4685,N_3515,N_3330);
nand U4686 (N_4686,N_3181,N_3509);
and U4687 (N_4687,N_3219,N_3016);
nand U4688 (N_4688,N_3285,N_3574);
xnor U4689 (N_4689,N_3266,N_3518);
xnor U4690 (N_4690,N_3004,N_3350);
nand U4691 (N_4691,N_3093,N_3341);
nor U4692 (N_4692,N_3774,N_3090);
or U4693 (N_4693,N_3518,N_3106);
xnor U4694 (N_4694,N_3582,N_3657);
nand U4695 (N_4695,N_3202,N_3977);
nor U4696 (N_4696,N_3816,N_3768);
nand U4697 (N_4697,N_3661,N_3285);
xnor U4698 (N_4698,N_3637,N_3878);
xor U4699 (N_4699,N_3156,N_3059);
xor U4700 (N_4700,N_3135,N_3977);
xnor U4701 (N_4701,N_3980,N_3458);
and U4702 (N_4702,N_3844,N_3595);
or U4703 (N_4703,N_3438,N_3942);
xor U4704 (N_4704,N_3991,N_3524);
and U4705 (N_4705,N_3031,N_3138);
nor U4706 (N_4706,N_3194,N_3166);
nand U4707 (N_4707,N_3658,N_3412);
nand U4708 (N_4708,N_3359,N_3389);
nand U4709 (N_4709,N_3506,N_3043);
or U4710 (N_4710,N_3856,N_3593);
or U4711 (N_4711,N_3366,N_3891);
and U4712 (N_4712,N_3552,N_3060);
nor U4713 (N_4713,N_3403,N_3615);
nor U4714 (N_4714,N_3545,N_3185);
xor U4715 (N_4715,N_3908,N_3058);
and U4716 (N_4716,N_3985,N_3616);
and U4717 (N_4717,N_3070,N_3687);
or U4718 (N_4718,N_3076,N_3348);
nand U4719 (N_4719,N_3361,N_3980);
and U4720 (N_4720,N_3095,N_3569);
or U4721 (N_4721,N_3275,N_3742);
and U4722 (N_4722,N_3052,N_3927);
or U4723 (N_4723,N_3999,N_3941);
xnor U4724 (N_4724,N_3852,N_3590);
xnor U4725 (N_4725,N_3309,N_3726);
nor U4726 (N_4726,N_3333,N_3734);
nand U4727 (N_4727,N_3412,N_3092);
and U4728 (N_4728,N_3942,N_3327);
or U4729 (N_4729,N_3627,N_3745);
nor U4730 (N_4730,N_3100,N_3711);
xor U4731 (N_4731,N_3368,N_3266);
and U4732 (N_4732,N_3432,N_3411);
nor U4733 (N_4733,N_3117,N_3196);
nor U4734 (N_4734,N_3557,N_3041);
and U4735 (N_4735,N_3229,N_3907);
and U4736 (N_4736,N_3130,N_3490);
nand U4737 (N_4737,N_3350,N_3940);
xor U4738 (N_4738,N_3386,N_3644);
nor U4739 (N_4739,N_3796,N_3038);
or U4740 (N_4740,N_3949,N_3214);
or U4741 (N_4741,N_3378,N_3499);
or U4742 (N_4742,N_3616,N_3458);
xor U4743 (N_4743,N_3588,N_3863);
and U4744 (N_4744,N_3405,N_3038);
xor U4745 (N_4745,N_3150,N_3158);
xor U4746 (N_4746,N_3053,N_3419);
or U4747 (N_4747,N_3074,N_3813);
nand U4748 (N_4748,N_3790,N_3711);
or U4749 (N_4749,N_3586,N_3900);
nand U4750 (N_4750,N_3250,N_3210);
nand U4751 (N_4751,N_3257,N_3506);
and U4752 (N_4752,N_3591,N_3995);
nor U4753 (N_4753,N_3999,N_3065);
xnor U4754 (N_4754,N_3529,N_3199);
nand U4755 (N_4755,N_3487,N_3304);
or U4756 (N_4756,N_3742,N_3622);
nand U4757 (N_4757,N_3954,N_3598);
or U4758 (N_4758,N_3876,N_3157);
nand U4759 (N_4759,N_3563,N_3579);
nand U4760 (N_4760,N_3235,N_3157);
nor U4761 (N_4761,N_3617,N_3029);
or U4762 (N_4762,N_3017,N_3774);
nor U4763 (N_4763,N_3409,N_3820);
nor U4764 (N_4764,N_3694,N_3098);
and U4765 (N_4765,N_3840,N_3317);
nor U4766 (N_4766,N_3369,N_3366);
nor U4767 (N_4767,N_3359,N_3156);
nand U4768 (N_4768,N_3522,N_3997);
xnor U4769 (N_4769,N_3058,N_3828);
or U4770 (N_4770,N_3519,N_3113);
nor U4771 (N_4771,N_3900,N_3951);
and U4772 (N_4772,N_3468,N_3728);
nor U4773 (N_4773,N_3737,N_3507);
nor U4774 (N_4774,N_3784,N_3502);
and U4775 (N_4775,N_3055,N_3106);
xor U4776 (N_4776,N_3216,N_3852);
nand U4777 (N_4777,N_3749,N_3891);
and U4778 (N_4778,N_3022,N_3032);
or U4779 (N_4779,N_3060,N_3245);
and U4780 (N_4780,N_3275,N_3900);
xor U4781 (N_4781,N_3814,N_3729);
and U4782 (N_4782,N_3190,N_3706);
and U4783 (N_4783,N_3933,N_3293);
xnor U4784 (N_4784,N_3492,N_3418);
nand U4785 (N_4785,N_3910,N_3443);
xnor U4786 (N_4786,N_3545,N_3926);
xnor U4787 (N_4787,N_3194,N_3590);
and U4788 (N_4788,N_3348,N_3257);
or U4789 (N_4789,N_3834,N_3726);
or U4790 (N_4790,N_3264,N_3443);
or U4791 (N_4791,N_3823,N_3895);
or U4792 (N_4792,N_3008,N_3639);
or U4793 (N_4793,N_3665,N_3674);
and U4794 (N_4794,N_3844,N_3292);
xnor U4795 (N_4795,N_3490,N_3717);
or U4796 (N_4796,N_3694,N_3542);
xor U4797 (N_4797,N_3034,N_3009);
or U4798 (N_4798,N_3948,N_3490);
and U4799 (N_4799,N_3179,N_3560);
nor U4800 (N_4800,N_3152,N_3938);
xor U4801 (N_4801,N_3182,N_3066);
xor U4802 (N_4802,N_3879,N_3440);
nand U4803 (N_4803,N_3108,N_3709);
or U4804 (N_4804,N_3854,N_3322);
xor U4805 (N_4805,N_3954,N_3848);
and U4806 (N_4806,N_3126,N_3122);
nor U4807 (N_4807,N_3791,N_3157);
nand U4808 (N_4808,N_3069,N_3854);
or U4809 (N_4809,N_3250,N_3704);
nor U4810 (N_4810,N_3321,N_3922);
nor U4811 (N_4811,N_3204,N_3093);
nand U4812 (N_4812,N_3657,N_3897);
nand U4813 (N_4813,N_3551,N_3375);
xnor U4814 (N_4814,N_3357,N_3949);
xor U4815 (N_4815,N_3898,N_3145);
or U4816 (N_4816,N_3245,N_3242);
or U4817 (N_4817,N_3470,N_3603);
or U4818 (N_4818,N_3453,N_3695);
nor U4819 (N_4819,N_3499,N_3528);
nor U4820 (N_4820,N_3681,N_3184);
or U4821 (N_4821,N_3180,N_3891);
nor U4822 (N_4822,N_3290,N_3434);
xor U4823 (N_4823,N_3243,N_3267);
and U4824 (N_4824,N_3318,N_3427);
or U4825 (N_4825,N_3263,N_3764);
nand U4826 (N_4826,N_3397,N_3542);
or U4827 (N_4827,N_3543,N_3780);
and U4828 (N_4828,N_3791,N_3655);
or U4829 (N_4829,N_3895,N_3607);
nand U4830 (N_4830,N_3919,N_3270);
and U4831 (N_4831,N_3847,N_3785);
nand U4832 (N_4832,N_3683,N_3952);
and U4833 (N_4833,N_3856,N_3038);
xnor U4834 (N_4834,N_3343,N_3415);
nor U4835 (N_4835,N_3578,N_3761);
nor U4836 (N_4836,N_3875,N_3154);
xor U4837 (N_4837,N_3443,N_3009);
xnor U4838 (N_4838,N_3870,N_3842);
or U4839 (N_4839,N_3249,N_3667);
or U4840 (N_4840,N_3160,N_3625);
and U4841 (N_4841,N_3878,N_3020);
xor U4842 (N_4842,N_3807,N_3870);
nor U4843 (N_4843,N_3934,N_3569);
and U4844 (N_4844,N_3919,N_3394);
nor U4845 (N_4845,N_3596,N_3468);
nor U4846 (N_4846,N_3312,N_3311);
or U4847 (N_4847,N_3913,N_3804);
and U4848 (N_4848,N_3984,N_3455);
and U4849 (N_4849,N_3905,N_3829);
nand U4850 (N_4850,N_3924,N_3465);
nand U4851 (N_4851,N_3734,N_3407);
nand U4852 (N_4852,N_3123,N_3307);
nand U4853 (N_4853,N_3636,N_3603);
or U4854 (N_4854,N_3265,N_3475);
and U4855 (N_4855,N_3141,N_3770);
or U4856 (N_4856,N_3223,N_3680);
xnor U4857 (N_4857,N_3368,N_3327);
nor U4858 (N_4858,N_3572,N_3964);
nand U4859 (N_4859,N_3204,N_3247);
and U4860 (N_4860,N_3575,N_3883);
nand U4861 (N_4861,N_3862,N_3773);
xnor U4862 (N_4862,N_3768,N_3094);
nand U4863 (N_4863,N_3404,N_3698);
nor U4864 (N_4864,N_3021,N_3990);
xnor U4865 (N_4865,N_3706,N_3160);
nand U4866 (N_4866,N_3054,N_3050);
nor U4867 (N_4867,N_3764,N_3434);
and U4868 (N_4868,N_3093,N_3785);
nand U4869 (N_4869,N_3599,N_3467);
or U4870 (N_4870,N_3449,N_3476);
and U4871 (N_4871,N_3105,N_3404);
nand U4872 (N_4872,N_3967,N_3795);
xor U4873 (N_4873,N_3088,N_3983);
and U4874 (N_4874,N_3744,N_3440);
xor U4875 (N_4875,N_3560,N_3235);
nor U4876 (N_4876,N_3566,N_3637);
or U4877 (N_4877,N_3581,N_3577);
or U4878 (N_4878,N_3459,N_3794);
nand U4879 (N_4879,N_3856,N_3686);
xnor U4880 (N_4880,N_3350,N_3904);
nor U4881 (N_4881,N_3006,N_3053);
and U4882 (N_4882,N_3619,N_3997);
and U4883 (N_4883,N_3798,N_3671);
nor U4884 (N_4884,N_3759,N_3592);
xor U4885 (N_4885,N_3689,N_3894);
or U4886 (N_4886,N_3158,N_3826);
nand U4887 (N_4887,N_3599,N_3406);
nor U4888 (N_4888,N_3520,N_3682);
and U4889 (N_4889,N_3467,N_3490);
nand U4890 (N_4890,N_3946,N_3465);
nand U4891 (N_4891,N_3042,N_3056);
nand U4892 (N_4892,N_3140,N_3711);
and U4893 (N_4893,N_3001,N_3241);
xor U4894 (N_4894,N_3391,N_3242);
and U4895 (N_4895,N_3223,N_3145);
and U4896 (N_4896,N_3324,N_3452);
xor U4897 (N_4897,N_3917,N_3800);
nand U4898 (N_4898,N_3098,N_3998);
nand U4899 (N_4899,N_3066,N_3478);
nor U4900 (N_4900,N_3441,N_3176);
xnor U4901 (N_4901,N_3300,N_3594);
nor U4902 (N_4902,N_3001,N_3445);
nor U4903 (N_4903,N_3039,N_3411);
nor U4904 (N_4904,N_3304,N_3307);
nor U4905 (N_4905,N_3769,N_3880);
xor U4906 (N_4906,N_3138,N_3928);
nor U4907 (N_4907,N_3905,N_3410);
or U4908 (N_4908,N_3454,N_3344);
and U4909 (N_4909,N_3261,N_3618);
or U4910 (N_4910,N_3676,N_3928);
xor U4911 (N_4911,N_3477,N_3633);
or U4912 (N_4912,N_3986,N_3829);
nand U4913 (N_4913,N_3472,N_3441);
and U4914 (N_4914,N_3439,N_3171);
xor U4915 (N_4915,N_3003,N_3957);
or U4916 (N_4916,N_3144,N_3956);
nand U4917 (N_4917,N_3603,N_3966);
or U4918 (N_4918,N_3193,N_3461);
and U4919 (N_4919,N_3644,N_3399);
nor U4920 (N_4920,N_3220,N_3884);
or U4921 (N_4921,N_3842,N_3974);
or U4922 (N_4922,N_3838,N_3018);
nand U4923 (N_4923,N_3431,N_3280);
and U4924 (N_4924,N_3519,N_3795);
nor U4925 (N_4925,N_3683,N_3559);
and U4926 (N_4926,N_3316,N_3295);
xor U4927 (N_4927,N_3585,N_3109);
nor U4928 (N_4928,N_3375,N_3452);
nand U4929 (N_4929,N_3369,N_3375);
xnor U4930 (N_4930,N_3964,N_3628);
xnor U4931 (N_4931,N_3454,N_3797);
nand U4932 (N_4932,N_3253,N_3167);
nor U4933 (N_4933,N_3236,N_3885);
nand U4934 (N_4934,N_3552,N_3010);
or U4935 (N_4935,N_3504,N_3332);
nand U4936 (N_4936,N_3702,N_3187);
xor U4937 (N_4937,N_3888,N_3188);
nor U4938 (N_4938,N_3730,N_3635);
and U4939 (N_4939,N_3405,N_3270);
or U4940 (N_4940,N_3475,N_3494);
or U4941 (N_4941,N_3692,N_3312);
or U4942 (N_4942,N_3730,N_3978);
xor U4943 (N_4943,N_3024,N_3399);
or U4944 (N_4944,N_3459,N_3413);
nand U4945 (N_4945,N_3214,N_3068);
nand U4946 (N_4946,N_3006,N_3285);
nor U4947 (N_4947,N_3458,N_3470);
nor U4948 (N_4948,N_3359,N_3797);
and U4949 (N_4949,N_3789,N_3435);
and U4950 (N_4950,N_3086,N_3850);
nand U4951 (N_4951,N_3136,N_3778);
and U4952 (N_4952,N_3437,N_3121);
nor U4953 (N_4953,N_3344,N_3288);
and U4954 (N_4954,N_3005,N_3623);
nor U4955 (N_4955,N_3112,N_3958);
nor U4956 (N_4956,N_3357,N_3730);
nor U4957 (N_4957,N_3914,N_3115);
xor U4958 (N_4958,N_3305,N_3127);
and U4959 (N_4959,N_3238,N_3131);
xor U4960 (N_4960,N_3076,N_3161);
xnor U4961 (N_4961,N_3329,N_3746);
or U4962 (N_4962,N_3396,N_3661);
nand U4963 (N_4963,N_3881,N_3828);
nand U4964 (N_4964,N_3678,N_3633);
xor U4965 (N_4965,N_3965,N_3765);
nor U4966 (N_4966,N_3872,N_3563);
xnor U4967 (N_4967,N_3610,N_3984);
nor U4968 (N_4968,N_3871,N_3006);
and U4969 (N_4969,N_3137,N_3869);
or U4970 (N_4970,N_3962,N_3597);
or U4971 (N_4971,N_3478,N_3322);
xnor U4972 (N_4972,N_3527,N_3798);
nand U4973 (N_4973,N_3715,N_3444);
xor U4974 (N_4974,N_3971,N_3728);
nor U4975 (N_4975,N_3870,N_3822);
nand U4976 (N_4976,N_3554,N_3132);
nand U4977 (N_4977,N_3112,N_3660);
nor U4978 (N_4978,N_3324,N_3849);
xnor U4979 (N_4979,N_3616,N_3380);
nor U4980 (N_4980,N_3726,N_3602);
and U4981 (N_4981,N_3667,N_3553);
nor U4982 (N_4982,N_3420,N_3280);
nor U4983 (N_4983,N_3626,N_3457);
xnor U4984 (N_4984,N_3983,N_3703);
or U4985 (N_4985,N_3019,N_3751);
nand U4986 (N_4986,N_3356,N_3166);
xnor U4987 (N_4987,N_3491,N_3796);
or U4988 (N_4988,N_3174,N_3112);
xor U4989 (N_4989,N_3372,N_3952);
or U4990 (N_4990,N_3728,N_3859);
or U4991 (N_4991,N_3759,N_3897);
nor U4992 (N_4992,N_3256,N_3600);
xnor U4993 (N_4993,N_3564,N_3593);
and U4994 (N_4994,N_3219,N_3618);
and U4995 (N_4995,N_3300,N_3185);
or U4996 (N_4996,N_3438,N_3206);
and U4997 (N_4997,N_3108,N_3946);
nand U4998 (N_4998,N_3934,N_3777);
nor U4999 (N_4999,N_3026,N_3474);
nand U5000 (N_5000,N_4582,N_4988);
nor U5001 (N_5001,N_4833,N_4766);
and U5002 (N_5002,N_4401,N_4596);
nand U5003 (N_5003,N_4884,N_4477);
nand U5004 (N_5004,N_4839,N_4705);
nor U5005 (N_5005,N_4269,N_4457);
nand U5006 (N_5006,N_4526,N_4784);
or U5007 (N_5007,N_4644,N_4449);
or U5008 (N_5008,N_4628,N_4516);
nand U5009 (N_5009,N_4267,N_4176);
or U5010 (N_5010,N_4216,N_4482);
nor U5011 (N_5011,N_4198,N_4320);
nor U5012 (N_5012,N_4575,N_4346);
or U5013 (N_5013,N_4723,N_4666);
and U5014 (N_5014,N_4037,N_4831);
and U5015 (N_5015,N_4060,N_4202);
and U5016 (N_5016,N_4057,N_4687);
xor U5017 (N_5017,N_4928,N_4150);
and U5018 (N_5018,N_4053,N_4740);
or U5019 (N_5019,N_4918,N_4563);
nand U5020 (N_5020,N_4820,N_4138);
nand U5021 (N_5021,N_4525,N_4901);
nand U5022 (N_5022,N_4545,N_4636);
nand U5023 (N_5023,N_4131,N_4388);
xor U5024 (N_5024,N_4682,N_4700);
xnor U5025 (N_5025,N_4667,N_4613);
or U5026 (N_5026,N_4837,N_4883);
and U5027 (N_5027,N_4913,N_4826);
nand U5028 (N_5028,N_4310,N_4830);
nor U5029 (N_5029,N_4409,N_4514);
nand U5030 (N_5030,N_4044,N_4009);
nor U5031 (N_5031,N_4195,N_4437);
nand U5032 (N_5032,N_4502,N_4219);
nand U5033 (N_5033,N_4121,N_4799);
nand U5034 (N_5034,N_4134,N_4810);
xnor U5035 (N_5035,N_4816,N_4846);
or U5036 (N_5036,N_4777,N_4112);
nand U5037 (N_5037,N_4709,N_4767);
nor U5038 (N_5038,N_4094,N_4424);
or U5039 (N_5039,N_4133,N_4298);
and U5040 (N_5040,N_4466,N_4370);
xor U5041 (N_5041,N_4908,N_4534);
nand U5042 (N_5042,N_4211,N_4435);
and U5043 (N_5043,N_4296,N_4841);
nand U5044 (N_5044,N_4220,N_4735);
or U5045 (N_5045,N_4379,N_4601);
and U5046 (N_5046,N_4077,N_4484);
and U5047 (N_5047,N_4556,N_4832);
or U5048 (N_5048,N_4641,N_4168);
nand U5049 (N_5049,N_4201,N_4270);
xor U5050 (N_5050,N_4209,N_4969);
nand U5051 (N_5051,N_4473,N_4172);
nand U5052 (N_5052,N_4366,N_4423);
nand U5053 (N_5053,N_4142,N_4371);
nand U5054 (N_5054,N_4452,N_4715);
and U5055 (N_5055,N_4807,N_4868);
nand U5056 (N_5056,N_4032,N_4660);
and U5057 (N_5057,N_4224,N_4471);
xor U5058 (N_5058,N_4994,N_4096);
nor U5059 (N_5059,N_4745,N_4809);
nand U5060 (N_5060,N_4936,N_4701);
nand U5061 (N_5061,N_4584,N_4113);
and U5062 (N_5062,N_4443,N_4998);
xnor U5063 (N_5063,N_4611,N_4204);
nand U5064 (N_5064,N_4271,N_4505);
or U5065 (N_5065,N_4690,N_4149);
xnor U5066 (N_5066,N_4532,N_4704);
nor U5067 (N_5067,N_4651,N_4865);
and U5068 (N_5068,N_4586,N_4965);
and U5069 (N_5069,N_4943,N_4670);
and U5070 (N_5070,N_4020,N_4529);
xnor U5071 (N_5071,N_4266,N_4001);
and U5072 (N_5072,N_4863,N_4402);
or U5073 (N_5073,N_4978,N_4173);
nor U5074 (N_5074,N_4265,N_4562);
or U5075 (N_5075,N_4671,N_4523);
and U5076 (N_5076,N_4903,N_4480);
nor U5077 (N_5077,N_4421,N_4025);
xnor U5078 (N_5078,N_4334,N_4742);
xnor U5079 (N_5079,N_4721,N_4243);
nand U5080 (N_5080,N_4987,N_4707);
nor U5081 (N_5081,N_4264,N_4823);
or U5082 (N_5082,N_4668,N_4245);
nand U5083 (N_5083,N_4227,N_4153);
xor U5084 (N_5084,N_4695,N_4445);
xnor U5085 (N_5085,N_4114,N_4862);
or U5086 (N_5086,N_4059,N_4256);
and U5087 (N_5087,N_4712,N_4045);
or U5088 (N_5088,N_4728,N_4738);
nand U5089 (N_5089,N_4536,N_4966);
xor U5090 (N_5090,N_4995,N_4842);
nand U5091 (N_5091,N_4981,N_4214);
and U5092 (N_5092,N_4018,N_4911);
nand U5093 (N_5093,N_4522,N_4447);
and U5094 (N_5094,N_4843,N_4039);
nand U5095 (N_5095,N_4249,N_4869);
and U5096 (N_5096,N_4308,N_4711);
or U5097 (N_5097,N_4576,N_4311);
or U5098 (N_5098,N_4864,N_4479);
and U5099 (N_5099,N_4905,N_4304);
and U5100 (N_5100,N_4193,N_4888);
and U5101 (N_5101,N_4789,N_4891);
nand U5102 (N_5102,N_4674,N_4254);
nand U5103 (N_5103,N_4467,N_4203);
xnor U5104 (N_5104,N_4947,N_4392);
nand U5105 (N_5105,N_4897,N_4182);
or U5106 (N_5106,N_4554,N_4827);
nand U5107 (N_5107,N_4364,N_4821);
or U5108 (N_5108,N_4898,N_4140);
xor U5109 (N_5109,N_4645,N_4907);
or U5110 (N_5110,N_4358,N_4323);
nand U5111 (N_5111,N_4836,N_4404);
and U5112 (N_5112,N_4231,N_4923);
or U5113 (N_5113,N_4188,N_4145);
nor U5114 (N_5114,N_4475,N_4159);
or U5115 (N_5115,N_4103,N_4946);
and U5116 (N_5116,N_4822,N_4210);
nor U5117 (N_5117,N_4335,N_4425);
and U5118 (N_5118,N_4034,N_4635);
or U5119 (N_5119,N_4253,N_4754);
xnor U5120 (N_5120,N_4881,N_4961);
or U5121 (N_5121,N_4250,N_4919);
and U5122 (N_5122,N_4438,N_4931);
nand U5123 (N_5123,N_4727,N_4314);
or U5124 (N_5124,N_4840,N_4079);
nor U5125 (N_5125,N_4024,N_4167);
nor U5126 (N_5126,N_4329,N_4436);
and U5127 (N_5127,N_4885,N_4819);
or U5128 (N_5128,N_4228,N_4110);
and U5129 (N_5129,N_4107,N_4893);
nor U5130 (N_5130,N_4647,N_4277);
or U5131 (N_5131,N_4458,N_4101);
nand U5132 (N_5132,N_4949,N_4190);
or U5133 (N_5133,N_4706,N_4515);
xnor U5134 (N_5134,N_4970,N_4147);
or U5135 (N_5135,N_4000,N_4128);
nand U5136 (N_5136,N_4415,N_4544);
or U5137 (N_5137,N_4504,N_4899);
and U5138 (N_5138,N_4261,N_4744);
nand U5139 (N_5139,N_4632,N_4280);
or U5140 (N_5140,N_4551,N_4708);
nor U5141 (N_5141,N_4681,N_4774);
or U5142 (N_5142,N_4200,N_4768);
xor U5143 (N_5143,N_4895,N_4360);
nand U5144 (N_5144,N_4629,N_4235);
nand U5145 (N_5145,N_4430,N_4794);
and U5146 (N_5146,N_4619,N_4866);
xor U5147 (N_5147,N_4796,N_4069);
nor U5148 (N_5148,N_4043,N_4495);
or U5149 (N_5149,N_4178,N_4410);
or U5150 (N_5150,N_4638,N_4130);
and U5151 (N_5151,N_4003,N_4603);
xnor U5152 (N_5152,N_4332,N_4143);
xor U5153 (N_5153,N_4456,N_4433);
and U5154 (N_5154,N_4263,N_4673);
nand U5155 (N_5155,N_4637,N_4412);
nand U5156 (N_5156,N_4073,N_4083);
or U5157 (N_5157,N_4325,N_4093);
and U5158 (N_5158,N_4353,N_4592);
and U5159 (N_5159,N_4717,N_4982);
nor U5160 (N_5160,N_4976,N_4012);
nor U5161 (N_5161,N_4450,N_4196);
and U5162 (N_5162,N_4086,N_4252);
and U5163 (N_5163,N_4500,N_4541);
and U5164 (N_5164,N_4815,N_4104);
or U5165 (N_5165,N_4860,N_4478);
nand U5166 (N_5166,N_4318,N_4848);
nand U5167 (N_5167,N_4382,N_4092);
or U5168 (N_5168,N_4071,N_4122);
and U5169 (N_5169,N_4274,N_4026);
nand U5170 (N_5170,N_4874,N_4236);
xor U5171 (N_5171,N_4278,N_4205);
nor U5172 (N_5172,N_4915,N_4411);
and U5173 (N_5173,N_4395,N_4446);
and U5174 (N_5174,N_4914,N_4572);
nand U5175 (N_5175,N_4646,N_4553);
xor U5176 (N_5176,N_4968,N_4782);
or U5177 (N_5177,N_4920,N_4950);
or U5178 (N_5178,N_4625,N_4959);
xnor U5179 (N_5179,N_4924,N_4187);
nand U5180 (N_5180,N_4129,N_4692);
nor U5181 (N_5181,N_4676,N_4569);
and U5182 (N_5182,N_4591,N_4088);
and U5183 (N_5183,N_4615,N_4791);
nor U5184 (N_5184,N_4369,N_4170);
xnor U5185 (N_5185,N_4238,N_4489);
and U5186 (N_5186,N_4564,N_4230);
xor U5187 (N_5187,N_4005,N_4896);
nand U5188 (N_5188,N_4599,N_4531);
nand U5189 (N_5189,N_4886,N_4416);
nor U5190 (N_5190,N_4349,N_4486);
xnor U5191 (N_5191,N_4028,N_4776);
nor U5192 (N_5192,N_4418,N_4558);
and U5193 (N_5193,N_4834,N_4922);
nand U5194 (N_5194,N_4702,N_4498);
and U5195 (N_5195,N_4180,N_4900);
nor U5196 (N_5196,N_4684,N_4055);
xnor U5197 (N_5197,N_4612,N_4503);
and U5198 (N_5198,N_4838,N_4882);
and U5199 (N_5199,N_4626,N_4019);
and U5200 (N_5200,N_4795,N_4460);
or U5201 (N_5201,N_4117,N_4521);
nand U5202 (N_5202,N_4483,N_4499);
xor U5203 (N_5203,N_4002,N_4533);
xor U5204 (N_5204,N_4488,N_4281);
nand U5205 (N_5205,N_4746,N_4474);
xor U5206 (N_5206,N_4260,N_4125);
nand U5207 (N_5207,N_4643,N_4123);
nand U5208 (N_5208,N_4307,N_4689);
and U5209 (N_5209,N_4105,N_4441);
xor U5210 (N_5210,N_4588,N_4455);
nor U5211 (N_5211,N_4621,N_4806);
nand U5212 (N_5212,N_4115,N_4313);
nor U5213 (N_5213,N_4889,N_4273);
xor U5214 (N_5214,N_4322,N_4930);
nor U5215 (N_5215,N_4546,N_4171);
and U5216 (N_5216,N_4878,N_4607);
or U5217 (N_5217,N_4381,N_4585);
and U5218 (N_5218,N_4539,N_4099);
nand U5219 (N_5219,N_4944,N_4528);
nand U5220 (N_5220,N_4547,N_4925);
nor U5221 (N_5221,N_4622,N_4972);
nand U5222 (N_5222,N_4511,N_4319);
xor U5223 (N_5223,N_4633,N_4952);
nand U5224 (N_5224,N_4679,N_4779);
nor U5225 (N_5225,N_4288,N_4075);
nor U5226 (N_5226,N_4858,N_4751);
nand U5227 (N_5227,N_4999,N_4461);
or U5228 (N_5228,N_4383,N_4800);
nor U5229 (N_5229,N_4036,N_4734);
and U5230 (N_5230,N_4783,N_4151);
xnor U5231 (N_5231,N_4760,N_4451);
nand U5232 (N_5232,N_4041,N_4747);
xor U5233 (N_5233,N_4297,N_4384);
nor U5234 (N_5234,N_4741,N_4778);
or U5235 (N_5235,N_4492,N_4470);
nor U5236 (N_5236,N_4165,N_4337);
xnor U5237 (N_5237,N_4251,N_4213);
xnor U5238 (N_5238,N_4589,N_4089);
and U5239 (N_5239,N_4653,N_4758);
or U5240 (N_5240,N_4669,N_4852);
or U5241 (N_5241,N_4377,N_4772);
and U5242 (N_5242,N_4971,N_4434);
nand U5243 (N_5243,N_4139,N_4752);
nand U5244 (N_5244,N_4067,N_4262);
nand U5245 (N_5245,N_4602,N_4697);
or U5246 (N_5246,N_4798,N_4387);
and U5247 (N_5247,N_4229,N_4835);
and U5248 (N_5248,N_4341,N_4517);
and U5249 (N_5249,N_4102,N_4127);
nand U5250 (N_5250,N_4007,N_4512);
xnor U5251 (N_5251,N_4773,N_4081);
nand U5252 (N_5252,N_4221,N_4465);
and U5253 (N_5253,N_4380,N_4469);
and U5254 (N_5254,N_4937,N_4743);
or U5255 (N_5255,N_4312,N_4141);
nand U5256 (N_5256,N_4340,N_4004);
or U5257 (N_5257,N_4080,N_4725);
nand U5258 (N_5258,N_4934,N_4351);
xnor U5259 (N_5259,N_4476,N_4485);
nor U5260 (N_5260,N_4400,N_4661);
and U5261 (N_5261,N_4552,N_4225);
and U5262 (N_5262,N_4775,N_4082);
and U5263 (N_5263,N_4010,N_4710);
or U5264 (N_5264,N_4166,N_4718);
xnor U5265 (N_5265,N_4194,N_4688);
nand U5266 (N_5266,N_4524,N_4716);
nor U5267 (N_5267,N_4570,N_4070);
or U5268 (N_5268,N_4406,N_4904);
and U5269 (N_5269,N_4493,N_4391);
and U5270 (N_5270,N_4283,N_4509);
or U5271 (N_5271,N_4954,N_4289);
and U5272 (N_5272,N_4605,N_4733);
and U5273 (N_5273,N_4973,N_4785);
xor U5274 (N_5274,N_4574,N_4355);
and U5275 (N_5275,N_4063,N_4303);
and U5276 (N_5276,N_4540,N_4111);
nand U5277 (N_5277,N_4126,N_4953);
or U5278 (N_5278,N_4136,N_4315);
and U5279 (N_5279,N_4013,N_4354);
and U5280 (N_5280,N_4109,N_4218);
nor U5281 (N_5281,N_4549,N_4805);
nand U5282 (N_5282,N_4336,N_4639);
or U5283 (N_5283,N_4964,N_4665);
nor U5284 (N_5284,N_4051,N_4124);
nor U5285 (N_5285,N_4282,N_4390);
nor U5286 (N_5286,N_4365,N_4958);
nand U5287 (N_5287,N_4581,N_4031);
nor U5288 (N_5288,N_4861,N_4120);
or U5289 (N_5289,N_4719,N_4156);
xnor U5290 (N_5290,N_4917,N_4787);
and U5291 (N_5291,N_4326,N_4975);
nor U5292 (N_5292,N_4508,N_4983);
or U5293 (N_5293,N_4825,N_4542);
nor U5294 (N_5294,N_4164,N_4650);
or U5295 (N_5295,N_4590,N_4640);
xnor U5296 (N_5296,N_4299,N_4372);
or U5297 (N_5297,N_4812,N_4426);
or U5298 (N_5298,N_4330,N_4792);
or U5299 (N_5299,N_4610,N_4560);
and U5300 (N_5300,N_4941,N_4763);
xnor U5301 (N_5301,N_4118,N_4685);
or U5302 (N_5302,N_4662,N_4146);
and U5303 (N_5303,N_4939,N_4916);
and U5304 (N_5304,N_4338,N_4955);
or U5305 (N_5305,N_4683,N_4921);
nor U5306 (N_5306,N_4356,N_4321);
and U5307 (N_5307,N_4873,N_4698);
nand U5308 (N_5308,N_4847,N_4246);
nand U5309 (N_5309,N_4659,N_4343);
and U5310 (N_5310,N_4068,N_4054);
nand U5311 (N_5311,N_4306,N_4248);
or U5312 (N_5312,N_4344,N_4163);
nor U5313 (N_5313,N_4023,N_4046);
xnor U5314 (N_5314,N_4394,N_4285);
nor U5315 (N_5315,N_4749,N_4030);
or U5316 (N_5316,N_4654,N_4872);
nand U5317 (N_5317,N_4573,N_4183);
xnor U5318 (N_5318,N_4957,N_4440);
and U5319 (N_5319,N_4510,N_4993);
nand U5320 (N_5320,N_4997,N_4902);
nand U5321 (N_5321,N_4407,N_4491);
or U5322 (N_5322,N_4977,N_4557);
nor U5323 (N_5323,N_4568,N_4604);
nor U5324 (N_5324,N_4960,N_4648);
nand U5325 (N_5325,N_4561,N_4595);
and U5326 (N_5326,N_4879,N_4880);
xor U5327 (N_5327,N_4513,N_4609);
and U5328 (N_5328,N_4212,N_4756);
or U5329 (N_5329,N_4011,N_4757);
nor U5330 (N_5330,N_4762,N_4696);
nand U5331 (N_5331,N_4148,N_4655);
nand U5332 (N_5332,N_4362,N_4694);
or U5333 (N_5333,N_4932,N_4630);
nor U5334 (N_5334,N_4929,N_4824);
or U5335 (N_5335,N_4061,N_4062);
xor U5336 (N_5336,N_4520,N_4597);
nor U5337 (N_5337,N_4287,N_4293);
nand U5338 (N_5338,N_4006,N_4593);
or U5339 (N_5339,N_4331,N_4518);
and U5340 (N_5340,N_4276,N_4234);
or U5341 (N_5341,N_4184,N_4255);
xnor U5342 (N_5342,N_4468,N_4890);
nor U5343 (N_5343,N_4571,N_4459);
and U5344 (N_5344,N_4771,N_4226);
nand U5345 (N_5345,N_4155,N_4162);
or U5346 (N_5346,N_4014,N_4040);
and U5347 (N_5347,N_4803,N_4286);
nor U5348 (N_5348,N_4686,N_4239);
xnor U5349 (N_5349,N_4186,N_4550);
nor U5350 (N_5350,N_4420,N_4714);
xnor U5351 (N_5351,N_4097,N_4295);
nor U5352 (N_5352,N_4979,N_4699);
nand U5353 (N_5353,N_4537,N_4462);
nand U5354 (N_5354,N_4577,N_4967);
or U5355 (N_5355,N_4066,N_4616);
nor U5356 (N_5356,N_4910,N_4802);
nand U5357 (N_5357,N_4813,N_4347);
nand U5358 (N_5358,N_4927,N_4814);
and U5359 (N_5359,N_4132,N_4948);
or U5360 (N_5360,N_4161,N_4399);
xnor U5361 (N_5361,N_4519,N_4207);
and U5362 (N_5362,N_4022,N_4828);
or U5363 (N_5363,N_4464,N_4021);
nor U5364 (N_5364,N_4317,N_4870);
nand U5365 (N_5365,N_4427,N_4962);
nand U5366 (N_5366,N_4567,N_4432);
xor U5367 (N_5367,N_4217,N_4631);
nand U5368 (N_5368,N_4854,N_4781);
nor U5369 (N_5369,N_4566,N_4678);
and U5370 (N_5370,N_4215,N_4652);
nor U5371 (N_5371,N_4853,N_4185);
nand U5372 (N_5372,N_4753,N_4675);
nor U5373 (N_5373,N_4750,N_4892);
and U5374 (N_5374,N_4877,N_4378);
and U5375 (N_5375,N_4078,N_4578);
xor U5376 (N_5376,N_4444,N_4691);
xor U5377 (N_5377,N_4851,N_4116);
and U5378 (N_5378,N_4240,N_4793);
and U5379 (N_5379,N_4199,N_4108);
or U5380 (N_5380,N_4015,N_4598);
nand U5381 (N_5381,N_4726,N_4414);
and U5382 (N_5382,N_4759,N_4780);
and U5383 (N_5383,N_4376,N_4845);
and U5384 (N_5384,N_4072,N_4087);
nor U5385 (N_5385,N_4487,N_4247);
xor U5386 (N_5386,N_4580,N_4618);
and U5387 (N_5387,N_4237,N_4453);
or U5388 (N_5388,N_4693,N_4986);
xor U5389 (N_5389,N_4100,N_4990);
nor U5390 (N_5390,N_4565,N_4137);
and U5391 (N_5391,N_4413,N_4876);
xor U5392 (N_5392,N_4175,N_4033);
nand U5393 (N_5393,N_4179,N_4048);
xnor U5394 (N_5394,N_4152,N_4984);
xor U5395 (N_5395,N_4909,N_4912);
nand U5396 (N_5396,N_4106,N_4906);
or U5397 (N_5397,N_4985,N_4206);
nand U5398 (N_5398,N_4333,N_4680);
or U5399 (N_5399,N_4940,N_4797);
or U5400 (N_5400,N_4594,N_4047);
or U5401 (N_5401,N_4790,N_4135);
nor U5402 (N_5402,N_4942,N_4084);
and U5403 (N_5403,N_4850,N_4016);
xor U5404 (N_5404,N_4027,N_4829);
or U5405 (N_5405,N_4405,N_4623);
xor U5406 (N_5406,N_4857,N_4098);
and U5407 (N_5407,N_4448,N_4309);
or U5408 (N_5408,N_4656,N_4494);
nor U5409 (N_5409,N_4535,N_4677);
or U5410 (N_5410,N_4974,N_4038);
nor U5411 (N_5411,N_4764,N_4454);
nand U5412 (N_5412,N_4339,N_4992);
and U5413 (N_5413,N_4703,N_4818);
xnor U5414 (N_5414,N_4042,N_4367);
xnor U5415 (N_5415,N_4350,N_4731);
nand U5416 (N_5416,N_4403,N_4272);
xnor U5417 (N_5417,N_4419,N_4801);
nor U5418 (N_5418,N_4357,N_4713);
nand U5419 (N_5419,N_4538,N_4770);
and U5420 (N_5420,N_4373,N_4617);
nand U5421 (N_5421,N_4634,N_4233);
and U5422 (N_5422,N_4472,N_4232);
nor U5423 (N_5423,N_4844,N_4490);
xnor U5424 (N_5424,N_4374,N_4649);
or U5425 (N_5425,N_4050,N_4730);
nand U5426 (N_5426,N_4608,N_4359);
and U5427 (N_5427,N_4189,N_4257);
and U5428 (N_5428,N_4951,N_4056);
or U5429 (N_5429,N_4739,N_4428);
nand U5430 (N_5430,N_4144,N_4658);
xor U5431 (N_5431,N_4157,N_4052);
nor U5432 (N_5432,N_4049,N_4393);
or U5433 (N_5433,N_4933,N_4191);
and U5434 (N_5434,N_4991,N_4761);
nor U5435 (N_5435,N_4368,N_4849);
xnor U5436 (N_5436,N_4158,N_4302);
nand U5437 (N_5437,N_4291,N_4284);
xnor U5438 (N_5438,N_4090,N_4555);
nand U5439 (N_5439,N_4624,N_4769);
or U5440 (N_5440,N_4095,N_4530);
nand U5441 (N_5441,N_4657,N_4808);
xnor U5442 (N_5442,N_4980,N_4279);
and U5443 (N_5443,N_4664,N_4497);
and U5444 (N_5444,N_4856,N_4804);
nor U5445 (N_5445,N_4956,N_4169);
nand U5446 (N_5446,N_4463,N_4290);
or U5447 (N_5447,N_4398,N_4672);
and U5448 (N_5448,N_4208,N_4259);
and U5449 (N_5449,N_4663,N_4543);
xor U5450 (N_5450,N_4065,N_4501);
and U5451 (N_5451,N_4408,N_4345);
nand U5452 (N_5452,N_4017,N_4222);
or U5453 (N_5453,N_4327,N_4305);
nor U5454 (N_5454,N_4342,N_4328);
nor U5455 (N_5455,N_4720,N_4064);
or U5456 (N_5456,N_4361,N_4788);
or U5457 (N_5457,N_4627,N_4765);
xnor U5458 (N_5458,N_4085,N_4348);
nor U5459 (N_5459,N_4363,N_4887);
and U5460 (N_5460,N_4008,N_4076);
or U5461 (N_5461,N_4268,N_4894);
nand U5462 (N_5462,N_4417,N_4507);
or U5463 (N_5463,N_4496,N_4755);
xnor U5464 (N_5464,N_4811,N_4935);
and U5465 (N_5465,N_4642,N_4963);
nand U5466 (N_5466,N_4292,N_4275);
nor U5467 (N_5467,N_4481,N_4736);
and U5468 (N_5468,N_4241,N_4729);
nand U5469 (N_5469,N_4871,N_4385);
or U5470 (N_5470,N_4091,N_4074);
xor U5471 (N_5471,N_4389,N_4396);
nand U5472 (N_5472,N_4375,N_4386);
nand U5473 (N_5473,N_4855,N_4748);
nor U5474 (N_5474,N_4301,N_4737);
and U5475 (N_5475,N_4119,N_4786);
nor U5476 (N_5476,N_4352,N_4732);
nand U5477 (N_5477,N_4527,N_4945);
xnor U5478 (N_5478,N_4316,N_4192);
or U5479 (N_5479,N_4579,N_4875);
nor U5480 (N_5480,N_4506,N_4559);
xnor U5481 (N_5481,N_4422,N_4867);
or U5482 (N_5482,N_4926,N_4242);
xnor U5483 (N_5483,N_4258,N_4724);
or U5484 (N_5484,N_4548,N_4300);
nand U5485 (N_5485,N_4197,N_4587);
nor U5486 (N_5486,N_4029,N_4429);
and U5487 (N_5487,N_4174,N_4431);
and U5488 (N_5488,N_4439,N_4244);
nand U5489 (N_5489,N_4294,N_4989);
nand U5490 (N_5490,N_4160,N_4442);
xnor U5491 (N_5491,N_4620,N_4996);
xnor U5492 (N_5492,N_4154,N_4324);
nor U5493 (N_5493,N_4583,N_4722);
nor U5494 (N_5494,N_4600,N_4397);
xor U5495 (N_5495,N_4817,N_4614);
or U5496 (N_5496,N_4181,N_4859);
nor U5497 (N_5497,N_4606,N_4938);
nand U5498 (N_5498,N_4058,N_4177);
nand U5499 (N_5499,N_4223,N_4035);
and U5500 (N_5500,N_4834,N_4545);
xor U5501 (N_5501,N_4034,N_4492);
xnor U5502 (N_5502,N_4003,N_4112);
or U5503 (N_5503,N_4199,N_4008);
nand U5504 (N_5504,N_4834,N_4717);
or U5505 (N_5505,N_4314,N_4762);
xnor U5506 (N_5506,N_4647,N_4893);
and U5507 (N_5507,N_4867,N_4895);
nand U5508 (N_5508,N_4419,N_4754);
xor U5509 (N_5509,N_4288,N_4533);
xnor U5510 (N_5510,N_4319,N_4728);
or U5511 (N_5511,N_4643,N_4445);
or U5512 (N_5512,N_4576,N_4450);
or U5513 (N_5513,N_4442,N_4346);
or U5514 (N_5514,N_4265,N_4836);
nand U5515 (N_5515,N_4140,N_4583);
xnor U5516 (N_5516,N_4317,N_4839);
nand U5517 (N_5517,N_4822,N_4778);
nor U5518 (N_5518,N_4749,N_4948);
and U5519 (N_5519,N_4554,N_4431);
and U5520 (N_5520,N_4421,N_4078);
nor U5521 (N_5521,N_4203,N_4631);
and U5522 (N_5522,N_4196,N_4604);
or U5523 (N_5523,N_4859,N_4646);
and U5524 (N_5524,N_4160,N_4735);
xor U5525 (N_5525,N_4715,N_4830);
nor U5526 (N_5526,N_4064,N_4270);
nand U5527 (N_5527,N_4998,N_4717);
nand U5528 (N_5528,N_4258,N_4480);
and U5529 (N_5529,N_4341,N_4067);
nor U5530 (N_5530,N_4628,N_4635);
xnor U5531 (N_5531,N_4294,N_4624);
and U5532 (N_5532,N_4527,N_4632);
nand U5533 (N_5533,N_4758,N_4629);
nand U5534 (N_5534,N_4233,N_4269);
nor U5535 (N_5535,N_4443,N_4484);
nand U5536 (N_5536,N_4970,N_4527);
nor U5537 (N_5537,N_4798,N_4669);
xor U5538 (N_5538,N_4596,N_4179);
nor U5539 (N_5539,N_4350,N_4856);
nor U5540 (N_5540,N_4966,N_4263);
nor U5541 (N_5541,N_4876,N_4830);
and U5542 (N_5542,N_4172,N_4318);
and U5543 (N_5543,N_4448,N_4557);
nor U5544 (N_5544,N_4566,N_4289);
and U5545 (N_5545,N_4310,N_4051);
and U5546 (N_5546,N_4058,N_4800);
nand U5547 (N_5547,N_4297,N_4193);
nor U5548 (N_5548,N_4651,N_4116);
nor U5549 (N_5549,N_4996,N_4345);
nand U5550 (N_5550,N_4322,N_4847);
or U5551 (N_5551,N_4449,N_4161);
nor U5552 (N_5552,N_4189,N_4450);
or U5553 (N_5553,N_4187,N_4489);
nor U5554 (N_5554,N_4803,N_4754);
and U5555 (N_5555,N_4095,N_4670);
xnor U5556 (N_5556,N_4771,N_4235);
nand U5557 (N_5557,N_4220,N_4502);
nor U5558 (N_5558,N_4059,N_4455);
nor U5559 (N_5559,N_4428,N_4770);
xnor U5560 (N_5560,N_4103,N_4549);
and U5561 (N_5561,N_4734,N_4625);
nor U5562 (N_5562,N_4543,N_4046);
and U5563 (N_5563,N_4440,N_4700);
nor U5564 (N_5564,N_4787,N_4869);
and U5565 (N_5565,N_4560,N_4137);
and U5566 (N_5566,N_4437,N_4767);
xor U5567 (N_5567,N_4497,N_4774);
nor U5568 (N_5568,N_4307,N_4946);
xor U5569 (N_5569,N_4777,N_4701);
nor U5570 (N_5570,N_4757,N_4933);
and U5571 (N_5571,N_4566,N_4089);
xor U5572 (N_5572,N_4491,N_4382);
xor U5573 (N_5573,N_4641,N_4831);
and U5574 (N_5574,N_4302,N_4872);
xor U5575 (N_5575,N_4572,N_4561);
and U5576 (N_5576,N_4184,N_4213);
and U5577 (N_5577,N_4044,N_4688);
xnor U5578 (N_5578,N_4556,N_4220);
or U5579 (N_5579,N_4738,N_4730);
xnor U5580 (N_5580,N_4785,N_4595);
and U5581 (N_5581,N_4834,N_4268);
xor U5582 (N_5582,N_4479,N_4788);
xnor U5583 (N_5583,N_4785,N_4626);
or U5584 (N_5584,N_4870,N_4635);
and U5585 (N_5585,N_4497,N_4854);
nor U5586 (N_5586,N_4445,N_4230);
nand U5587 (N_5587,N_4221,N_4267);
or U5588 (N_5588,N_4732,N_4170);
and U5589 (N_5589,N_4980,N_4331);
and U5590 (N_5590,N_4252,N_4176);
xnor U5591 (N_5591,N_4364,N_4657);
nor U5592 (N_5592,N_4395,N_4658);
or U5593 (N_5593,N_4835,N_4121);
nor U5594 (N_5594,N_4174,N_4557);
nor U5595 (N_5595,N_4809,N_4014);
nor U5596 (N_5596,N_4513,N_4634);
xor U5597 (N_5597,N_4007,N_4151);
and U5598 (N_5598,N_4909,N_4418);
nand U5599 (N_5599,N_4246,N_4736);
xnor U5600 (N_5600,N_4760,N_4974);
or U5601 (N_5601,N_4584,N_4019);
and U5602 (N_5602,N_4670,N_4902);
or U5603 (N_5603,N_4960,N_4755);
nor U5604 (N_5604,N_4380,N_4080);
and U5605 (N_5605,N_4202,N_4434);
xnor U5606 (N_5606,N_4141,N_4303);
xnor U5607 (N_5607,N_4773,N_4374);
xnor U5608 (N_5608,N_4513,N_4247);
nand U5609 (N_5609,N_4417,N_4027);
xnor U5610 (N_5610,N_4151,N_4723);
nor U5611 (N_5611,N_4061,N_4580);
nor U5612 (N_5612,N_4787,N_4543);
nor U5613 (N_5613,N_4922,N_4545);
nand U5614 (N_5614,N_4869,N_4178);
or U5615 (N_5615,N_4730,N_4614);
xor U5616 (N_5616,N_4434,N_4490);
or U5617 (N_5617,N_4972,N_4487);
and U5618 (N_5618,N_4583,N_4121);
or U5619 (N_5619,N_4781,N_4019);
xor U5620 (N_5620,N_4729,N_4296);
or U5621 (N_5621,N_4798,N_4386);
xor U5622 (N_5622,N_4704,N_4384);
nand U5623 (N_5623,N_4683,N_4767);
nand U5624 (N_5624,N_4416,N_4058);
xor U5625 (N_5625,N_4717,N_4009);
and U5626 (N_5626,N_4893,N_4727);
nor U5627 (N_5627,N_4766,N_4263);
and U5628 (N_5628,N_4597,N_4662);
and U5629 (N_5629,N_4400,N_4735);
or U5630 (N_5630,N_4024,N_4471);
xnor U5631 (N_5631,N_4011,N_4960);
nand U5632 (N_5632,N_4438,N_4916);
nand U5633 (N_5633,N_4985,N_4811);
and U5634 (N_5634,N_4177,N_4649);
and U5635 (N_5635,N_4174,N_4317);
nand U5636 (N_5636,N_4247,N_4052);
or U5637 (N_5637,N_4881,N_4893);
xor U5638 (N_5638,N_4748,N_4708);
nor U5639 (N_5639,N_4981,N_4578);
xor U5640 (N_5640,N_4900,N_4528);
or U5641 (N_5641,N_4333,N_4322);
and U5642 (N_5642,N_4682,N_4408);
nor U5643 (N_5643,N_4380,N_4906);
xnor U5644 (N_5644,N_4175,N_4454);
nor U5645 (N_5645,N_4339,N_4251);
or U5646 (N_5646,N_4834,N_4241);
and U5647 (N_5647,N_4900,N_4535);
and U5648 (N_5648,N_4691,N_4673);
and U5649 (N_5649,N_4718,N_4975);
nand U5650 (N_5650,N_4467,N_4284);
or U5651 (N_5651,N_4870,N_4984);
xor U5652 (N_5652,N_4583,N_4287);
nand U5653 (N_5653,N_4365,N_4831);
or U5654 (N_5654,N_4859,N_4416);
nand U5655 (N_5655,N_4734,N_4153);
or U5656 (N_5656,N_4542,N_4260);
xor U5657 (N_5657,N_4975,N_4521);
xnor U5658 (N_5658,N_4984,N_4571);
and U5659 (N_5659,N_4137,N_4341);
or U5660 (N_5660,N_4432,N_4912);
nand U5661 (N_5661,N_4779,N_4088);
and U5662 (N_5662,N_4731,N_4180);
nand U5663 (N_5663,N_4606,N_4590);
or U5664 (N_5664,N_4715,N_4338);
nand U5665 (N_5665,N_4974,N_4762);
nand U5666 (N_5666,N_4221,N_4810);
or U5667 (N_5667,N_4524,N_4603);
or U5668 (N_5668,N_4800,N_4019);
nand U5669 (N_5669,N_4937,N_4317);
xor U5670 (N_5670,N_4912,N_4194);
nand U5671 (N_5671,N_4994,N_4443);
nor U5672 (N_5672,N_4380,N_4173);
or U5673 (N_5673,N_4378,N_4172);
nand U5674 (N_5674,N_4300,N_4019);
and U5675 (N_5675,N_4102,N_4323);
xor U5676 (N_5676,N_4613,N_4649);
or U5677 (N_5677,N_4771,N_4730);
nor U5678 (N_5678,N_4286,N_4670);
nor U5679 (N_5679,N_4452,N_4042);
and U5680 (N_5680,N_4210,N_4633);
nand U5681 (N_5681,N_4863,N_4767);
or U5682 (N_5682,N_4765,N_4004);
nand U5683 (N_5683,N_4564,N_4859);
or U5684 (N_5684,N_4468,N_4505);
xor U5685 (N_5685,N_4323,N_4936);
or U5686 (N_5686,N_4203,N_4603);
nand U5687 (N_5687,N_4866,N_4800);
or U5688 (N_5688,N_4312,N_4609);
nor U5689 (N_5689,N_4830,N_4435);
and U5690 (N_5690,N_4494,N_4247);
and U5691 (N_5691,N_4762,N_4681);
and U5692 (N_5692,N_4491,N_4929);
nor U5693 (N_5693,N_4218,N_4058);
xor U5694 (N_5694,N_4323,N_4741);
and U5695 (N_5695,N_4998,N_4968);
and U5696 (N_5696,N_4118,N_4972);
nand U5697 (N_5697,N_4842,N_4591);
xnor U5698 (N_5698,N_4106,N_4721);
nand U5699 (N_5699,N_4707,N_4964);
and U5700 (N_5700,N_4147,N_4599);
or U5701 (N_5701,N_4238,N_4817);
nand U5702 (N_5702,N_4026,N_4145);
or U5703 (N_5703,N_4872,N_4246);
and U5704 (N_5704,N_4751,N_4140);
nor U5705 (N_5705,N_4405,N_4855);
nand U5706 (N_5706,N_4522,N_4103);
nor U5707 (N_5707,N_4951,N_4404);
and U5708 (N_5708,N_4939,N_4566);
nand U5709 (N_5709,N_4164,N_4614);
xnor U5710 (N_5710,N_4731,N_4624);
nand U5711 (N_5711,N_4446,N_4669);
and U5712 (N_5712,N_4568,N_4011);
xnor U5713 (N_5713,N_4736,N_4519);
xnor U5714 (N_5714,N_4364,N_4644);
or U5715 (N_5715,N_4481,N_4539);
xnor U5716 (N_5716,N_4853,N_4421);
or U5717 (N_5717,N_4707,N_4561);
nand U5718 (N_5718,N_4282,N_4620);
nor U5719 (N_5719,N_4308,N_4989);
nand U5720 (N_5720,N_4179,N_4940);
nor U5721 (N_5721,N_4187,N_4100);
or U5722 (N_5722,N_4462,N_4490);
xnor U5723 (N_5723,N_4213,N_4655);
xor U5724 (N_5724,N_4902,N_4080);
or U5725 (N_5725,N_4313,N_4158);
or U5726 (N_5726,N_4500,N_4912);
and U5727 (N_5727,N_4763,N_4354);
and U5728 (N_5728,N_4279,N_4937);
nor U5729 (N_5729,N_4613,N_4507);
and U5730 (N_5730,N_4350,N_4447);
nor U5731 (N_5731,N_4429,N_4219);
nor U5732 (N_5732,N_4853,N_4026);
nor U5733 (N_5733,N_4860,N_4888);
xor U5734 (N_5734,N_4996,N_4329);
xor U5735 (N_5735,N_4040,N_4491);
xor U5736 (N_5736,N_4839,N_4872);
or U5737 (N_5737,N_4314,N_4835);
xnor U5738 (N_5738,N_4298,N_4595);
and U5739 (N_5739,N_4706,N_4676);
or U5740 (N_5740,N_4802,N_4067);
and U5741 (N_5741,N_4187,N_4847);
and U5742 (N_5742,N_4167,N_4519);
and U5743 (N_5743,N_4417,N_4303);
nor U5744 (N_5744,N_4792,N_4129);
xnor U5745 (N_5745,N_4979,N_4758);
xnor U5746 (N_5746,N_4219,N_4419);
xor U5747 (N_5747,N_4406,N_4973);
or U5748 (N_5748,N_4625,N_4235);
or U5749 (N_5749,N_4262,N_4441);
and U5750 (N_5750,N_4184,N_4384);
or U5751 (N_5751,N_4372,N_4496);
nor U5752 (N_5752,N_4828,N_4431);
nor U5753 (N_5753,N_4854,N_4114);
or U5754 (N_5754,N_4894,N_4294);
nand U5755 (N_5755,N_4658,N_4252);
or U5756 (N_5756,N_4603,N_4954);
and U5757 (N_5757,N_4443,N_4749);
and U5758 (N_5758,N_4680,N_4637);
and U5759 (N_5759,N_4150,N_4163);
or U5760 (N_5760,N_4371,N_4424);
nor U5761 (N_5761,N_4839,N_4381);
nand U5762 (N_5762,N_4109,N_4532);
or U5763 (N_5763,N_4938,N_4740);
xor U5764 (N_5764,N_4877,N_4827);
or U5765 (N_5765,N_4416,N_4149);
and U5766 (N_5766,N_4395,N_4247);
and U5767 (N_5767,N_4671,N_4794);
nor U5768 (N_5768,N_4507,N_4702);
or U5769 (N_5769,N_4833,N_4620);
xor U5770 (N_5770,N_4659,N_4616);
or U5771 (N_5771,N_4393,N_4282);
or U5772 (N_5772,N_4881,N_4247);
and U5773 (N_5773,N_4143,N_4235);
xor U5774 (N_5774,N_4008,N_4083);
nor U5775 (N_5775,N_4051,N_4315);
nor U5776 (N_5776,N_4225,N_4537);
nor U5777 (N_5777,N_4218,N_4963);
xor U5778 (N_5778,N_4678,N_4348);
and U5779 (N_5779,N_4590,N_4004);
xnor U5780 (N_5780,N_4408,N_4555);
nand U5781 (N_5781,N_4920,N_4075);
nor U5782 (N_5782,N_4779,N_4790);
and U5783 (N_5783,N_4934,N_4867);
nand U5784 (N_5784,N_4210,N_4469);
nand U5785 (N_5785,N_4151,N_4434);
or U5786 (N_5786,N_4963,N_4104);
nor U5787 (N_5787,N_4316,N_4986);
nand U5788 (N_5788,N_4562,N_4750);
nand U5789 (N_5789,N_4865,N_4911);
and U5790 (N_5790,N_4766,N_4864);
nand U5791 (N_5791,N_4619,N_4540);
nand U5792 (N_5792,N_4635,N_4927);
nor U5793 (N_5793,N_4848,N_4567);
and U5794 (N_5794,N_4118,N_4259);
and U5795 (N_5795,N_4589,N_4240);
xor U5796 (N_5796,N_4328,N_4288);
and U5797 (N_5797,N_4786,N_4782);
xnor U5798 (N_5798,N_4993,N_4806);
xnor U5799 (N_5799,N_4140,N_4498);
or U5800 (N_5800,N_4513,N_4252);
or U5801 (N_5801,N_4456,N_4707);
and U5802 (N_5802,N_4281,N_4086);
nand U5803 (N_5803,N_4129,N_4706);
nand U5804 (N_5804,N_4078,N_4750);
nor U5805 (N_5805,N_4522,N_4111);
nand U5806 (N_5806,N_4613,N_4195);
nand U5807 (N_5807,N_4487,N_4401);
xor U5808 (N_5808,N_4033,N_4010);
nand U5809 (N_5809,N_4648,N_4624);
or U5810 (N_5810,N_4509,N_4359);
nand U5811 (N_5811,N_4631,N_4910);
and U5812 (N_5812,N_4704,N_4863);
or U5813 (N_5813,N_4440,N_4063);
xor U5814 (N_5814,N_4822,N_4879);
xnor U5815 (N_5815,N_4412,N_4623);
or U5816 (N_5816,N_4700,N_4034);
nor U5817 (N_5817,N_4978,N_4375);
nand U5818 (N_5818,N_4546,N_4319);
xor U5819 (N_5819,N_4529,N_4836);
xor U5820 (N_5820,N_4273,N_4838);
and U5821 (N_5821,N_4721,N_4278);
xnor U5822 (N_5822,N_4287,N_4619);
or U5823 (N_5823,N_4606,N_4868);
nand U5824 (N_5824,N_4946,N_4063);
nand U5825 (N_5825,N_4244,N_4130);
and U5826 (N_5826,N_4025,N_4932);
xnor U5827 (N_5827,N_4478,N_4187);
xor U5828 (N_5828,N_4572,N_4594);
or U5829 (N_5829,N_4622,N_4911);
or U5830 (N_5830,N_4531,N_4353);
nand U5831 (N_5831,N_4338,N_4701);
nand U5832 (N_5832,N_4178,N_4582);
or U5833 (N_5833,N_4713,N_4871);
nor U5834 (N_5834,N_4723,N_4695);
nor U5835 (N_5835,N_4406,N_4871);
or U5836 (N_5836,N_4081,N_4176);
or U5837 (N_5837,N_4537,N_4275);
or U5838 (N_5838,N_4660,N_4121);
nor U5839 (N_5839,N_4434,N_4765);
xor U5840 (N_5840,N_4597,N_4588);
xnor U5841 (N_5841,N_4450,N_4875);
nor U5842 (N_5842,N_4524,N_4329);
xor U5843 (N_5843,N_4492,N_4631);
and U5844 (N_5844,N_4553,N_4215);
nor U5845 (N_5845,N_4536,N_4336);
nor U5846 (N_5846,N_4981,N_4054);
or U5847 (N_5847,N_4538,N_4583);
xor U5848 (N_5848,N_4641,N_4871);
nand U5849 (N_5849,N_4129,N_4533);
or U5850 (N_5850,N_4648,N_4023);
or U5851 (N_5851,N_4242,N_4482);
xnor U5852 (N_5852,N_4936,N_4320);
or U5853 (N_5853,N_4321,N_4444);
nor U5854 (N_5854,N_4047,N_4131);
nor U5855 (N_5855,N_4007,N_4574);
or U5856 (N_5856,N_4823,N_4681);
nand U5857 (N_5857,N_4861,N_4963);
nand U5858 (N_5858,N_4778,N_4244);
xor U5859 (N_5859,N_4268,N_4166);
and U5860 (N_5860,N_4848,N_4418);
xor U5861 (N_5861,N_4055,N_4862);
or U5862 (N_5862,N_4240,N_4278);
or U5863 (N_5863,N_4886,N_4160);
or U5864 (N_5864,N_4808,N_4667);
nand U5865 (N_5865,N_4660,N_4313);
and U5866 (N_5866,N_4060,N_4125);
nor U5867 (N_5867,N_4083,N_4031);
xor U5868 (N_5868,N_4113,N_4632);
nand U5869 (N_5869,N_4467,N_4196);
nand U5870 (N_5870,N_4242,N_4622);
nor U5871 (N_5871,N_4290,N_4667);
or U5872 (N_5872,N_4854,N_4747);
or U5873 (N_5873,N_4109,N_4004);
or U5874 (N_5874,N_4298,N_4254);
nor U5875 (N_5875,N_4939,N_4789);
nor U5876 (N_5876,N_4254,N_4862);
nor U5877 (N_5877,N_4551,N_4568);
xnor U5878 (N_5878,N_4844,N_4733);
nand U5879 (N_5879,N_4745,N_4184);
and U5880 (N_5880,N_4199,N_4780);
or U5881 (N_5881,N_4546,N_4255);
nand U5882 (N_5882,N_4574,N_4328);
or U5883 (N_5883,N_4811,N_4980);
or U5884 (N_5884,N_4763,N_4696);
or U5885 (N_5885,N_4623,N_4977);
nand U5886 (N_5886,N_4750,N_4628);
xor U5887 (N_5887,N_4514,N_4202);
and U5888 (N_5888,N_4971,N_4972);
nor U5889 (N_5889,N_4070,N_4328);
or U5890 (N_5890,N_4072,N_4259);
nand U5891 (N_5891,N_4793,N_4453);
nor U5892 (N_5892,N_4846,N_4322);
nor U5893 (N_5893,N_4115,N_4783);
or U5894 (N_5894,N_4106,N_4130);
or U5895 (N_5895,N_4685,N_4221);
xor U5896 (N_5896,N_4824,N_4788);
nand U5897 (N_5897,N_4840,N_4241);
xor U5898 (N_5898,N_4741,N_4402);
xor U5899 (N_5899,N_4170,N_4638);
and U5900 (N_5900,N_4039,N_4925);
xor U5901 (N_5901,N_4300,N_4591);
and U5902 (N_5902,N_4783,N_4916);
and U5903 (N_5903,N_4445,N_4743);
nand U5904 (N_5904,N_4172,N_4603);
or U5905 (N_5905,N_4071,N_4521);
nand U5906 (N_5906,N_4206,N_4027);
nor U5907 (N_5907,N_4625,N_4523);
or U5908 (N_5908,N_4330,N_4850);
and U5909 (N_5909,N_4807,N_4598);
and U5910 (N_5910,N_4650,N_4072);
nor U5911 (N_5911,N_4213,N_4490);
or U5912 (N_5912,N_4336,N_4231);
xor U5913 (N_5913,N_4779,N_4848);
nor U5914 (N_5914,N_4416,N_4461);
and U5915 (N_5915,N_4856,N_4094);
or U5916 (N_5916,N_4348,N_4032);
xnor U5917 (N_5917,N_4908,N_4685);
nor U5918 (N_5918,N_4100,N_4093);
or U5919 (N_5919,N_4830,N_4285);
nor U5920 (N_5920,N_4406,N_4667);
xnor U5921 (N_5921,N_4069,N_4992);
or U5922 (N_5922,N_4590,N_4019);
nor U5923 (N_5923,N_4440,N_4401);
or U5924 (N_5924,N_4819,N_4763);
and U5925 (N_5925,N_4537,N_4603);
and U5926 (N_5926,N_4719,N_4307);
nor U5927 (N_5927,N_4757,N_4801);
xnor U5928 (N_5928,N_4849,N_4132);
or U5929 (N_5929,N_4744,N_4661);
xor U5930 (N_5930,N_4679,N_4379);
xnor U5931 (N_5931,N_4201,N_4680);
and U5932 (N_5932,N_4831,N_4361);
or U5933 (N_5933,N_4396,N_4781);
xor U5934 (N_5934,N_4572,N_4735);
nand U5935 (N_5935,N_4337,N_4627);
or U5936 (N_5936,N_4808,N_4020);
xor U5937 (N_5937,N_4818,N_4876);
and U5938 (N_5938,N_4306,N_4934);
and U5939 (N_5939,N_4779,N_4528);
nand U5940 (N_5940,N_4071,N_4959);
nor U5941 (N_5941,N_4281,N_4772);
nand U5942 (N_5942,N_4222,N_4433);
or U5943 (N_5943,N_4006,N_4322);
nor U5944 (N_5944,N_4776,N_4422);
or U5945 (N_5945,N_4411,N_4657);
and U5946 (N_5946,N_4508,N_4204);
nor U5947 (N_5947,N_4406,N_4082);
or U5948 (N_5948,N_4019,N_4972);
xor U5949 (N_5949,N_4741,N_4644);
and U5950 (N_5950,N_4013,N_4518);
xnor U5951 (N_5951,N_4683,N_4158);
nand U5952 (N_5952,N_4691,N_4921);
xor U5953 (N_5953,N_4001,N_4284);
xor U5954 (N_5954,N_4967,N_4206);
or U5955 (N_5955,N_4406,N_4476);
xnor U5956 (N_5956,N_4493,N_4909);
xor U5957 (N_5957,N_4127,N_4561);
xnor U5958 (N_5958,N_4023,N_4058);
or U5959 (N_5959,N_4091,N_4247);
xnor U5960 (N_5960,N_4819,N_4144);
or U5961 (N_5961,N_4001,N_4544);
xor U5962 (N_5962,N_4561,N_4642);
or U5963 (N_5963,N_4926,N_4985);
and U5964 (N_5964,N_4744,N_4758);
nand U5965 (N_5965,N_4059,N_4039);
or U5966 (N_5966,N_4622,N_4985);
nand U5967 (N_5967,N_4657,N_4980);
and U5968 (N_5968,N_4569,N_4727);
or U5969 (N_5969,N_4226,N_4393);
and U5970 (N_5970,N_4173,N_4218);
or U5971 (N_5971,N_4575,N_4801);
or U5972 (N_5972,N_4435,N_4725);
and U5973 (N_5973,N_4028,N_4467);
or U5974 (N_5974,N_4653,N_4808);
and U5975 (N_5975,N_4703,N_4505);
nor U5976 (N_5976,N_4035,N_4499);
and U5977 (N_5977,N_4178,N_4434);
xor U5978 (N_5978,N_4779,N_4627);
and U5979 (N_5979,N_4068,N_4763);
or U5980 (N_5980,N_4703,N_4211);
nand U5981 (N_5981,N_4511,N_4546);
nand U5982 (N_5982,N_4700,N_4797);
or U5983 (N_5983,N_4690,N_4960);
xnor U5984 (N_5984,N_4999,N_4297);
xnor U5985 (N_5985,N_4846,N_4715);
or U5986 (N_5986,N_4301,N_4615);
xnor U5987 (N_5987,N_4714,N_4991);
xnor U5988 (N_5988,N_4936,N_4371);
nand U5989 (N_5989,N_4976,N_4077);
and U5990 (N_5990,N_4060,N_4223);
xnor U5991 (N_5991,N_4092,N_4814);
and U5992 (N_5992,N_4546,N_4497);
xnor U5993 (N_5993,N_4821,N_4334);
nor U5994 (N_5994,N_4048,N_4010);
or U5995 (N_5995,N_4282,N_4800);
and U5996 (N_5996,N_4810,N_4674);
or U5997 (N_5997,N_4217,N_4718);
nand U5998 (N_5998,N_4565,N_4643);
nor U5999 (N_5999,N_4879,N_4618);
or U6000 (N_6000,N_5544,N_5181);
and U6001 (N_6001,N_5099,N_5106);
nor U6002 (N_6002,N_5180,N_5859);
or U6003 (N_6003,N_5906,N_5416);
xnor U6004 (N_6004,N_5741,N_5861);
nand U6005 (N_6005,N_5208,N_5693);
nor U6006 (N_6006,N_5471,N_5641);
and U6007 (N_6007,N_5549,N_5895);
or U6008 (N_6008,N_5989,N_5087);
xnor U6009 (N_6009,N_5766,N_5426);
nand U6010 (N_6010,N_5392,N_5232);
nor U6011 (N_6011,N_5311,N_5457);
and U6012 (N_6012,N_5004,N_5139);
and U6013 (N_6013,N_5753,N_5269);
xor U6014 (N_6014,N_5937,N_5639);
xor U6015 (N_6015,N_5170,N_5898);
xnor U6016 (N_6016,N_5039,N_5782);
xor U6017 (N_6017,N_5280,N_5955);
nor U6018 (N_6018,N_5108,N_5556);
and U6019 (N_6019,N_5899,N_5090);
nor U6020 (N_6020,N_5648,N_5680);
or U6021 (N_6021,N_5418,N_5671);
or U6022 (N_6022,N_5603,N_5963);
xor U6023 (N_6023,N_5456,N_5884);
or U6024 (N_6024,N_5797,N_5318);
and U6025 (N_6025,N_5515,N_5107);
nor U6026 (N_6026,N_5691,N_5427);
nand U6027 (N_6027,N_5351,N_5821);
xor U6028 (N_6028,N_5804,N_5966);
nand U6029 (N_6029,N_5529,N_5151);
and U6030 (N_6030,N_5740,N_5986);
and U6031 (N_6031,N_5612,N_5774);
and U6032 (N_6032,N_5074,N_5417);
and U6033 (N_6033,N_5422,N_5425);
nand U6034 (N_6034,N_5845,N_5564);
and U6035 (N_6035,N_5134,N_5551);
nor U6036 (N_6036,N_5993,N_5506);
xnor U6037 (N_6037,N_5485,N_5114);
or U6038 (N_6038,N_5300,N_5468);
nand U6039 (N_6039,N_5445,N_5027);
nand U6040 (N_6040,N_5721,N_5623);
nor U6041 (N_6041,N_5754,N_5032);
xor U6042 (N_6042,N_5540,N_5902);
xor U6043 (N_6043,N_5237,N_5781);
and U6044 (N_6044,N_5591,N_5281);
nand U6045 (N_6045,N_5524,N_5750);
or U6046 (N_6046,N_5562,N_5254);
nor U6047 (N_6047,N_5194,N_5361);
nor U6048 (N_6048,N_5917,N_5832);
xor U6049 (N_6049,N_5904,N_5408);
nor U6050 (N_6050,N_5923,N_5961);
or U6051 (N_6051,N_5119,N_5949);
and U6052 (N_6052,N_5589,N_5015);
and U6053 (N_6053,N_5203,N_5517);
or U6054 (N_6054,N_5795,N_5707);
or U6055 (N_6055,N_5331,N_5258);
nand U6056 (N_6056,N_5340,N_5465);
xor U6057 (N_6057,N_5089,N_5121);
and U6058 (N_6058,N_5251,N_5849);
xor U6059 (N_6059,N_5334,N_5950);
and U6060 (N_6060,N_5290,N_5244);
nor U6061 (N_6061,N_5373,N_5060);
or U6062 (N_6062,N_5262,N_5967);
nand U6063 (N_6063,N_5147,N_5588);
or U6064 (N_6064,N_5747,N_5609);
nand U6065 (N_6065,N_5135,N_5306);
or U6066 (N_6066,N_5379,N_5703);
xnor U6067 (N_6067,N_5935,N_5701);
or U6068 (N_6068,N_5994,N_5560);
xor U6069 (N_6069,N_5344,N_5620);
or U6070 (N_6070,N_5830,N_5856);
nand U6071 (N_6071,N_5828,N_5985);
xnor U6072 (N_6072,N_5679,N_5096);
and U6073 (N_6073,N_5948,N_5681);
nor U6074 (N_6074,N_5111,N_5778);
or U6075 (N_6075,N_5330,N_5532);
or U6076 (N_6076,N_5327,N_5137);
nor U6077 (N_6077,N_5548,N_5944);
nor U6078 (N_6078,N_5686,N_5077);
nor U6079 (N_6079,N_5525,N_5481);
nand U6080 (N_6080,N_5080,N_5836);
xor U6081 (N_6081,N_5055,N_5144);
and U6082 (N_6082,N_5382,N_5574);
xnor U6083 (N_6083,N_5822,N_5224);
or U6084 (N_6084,N_5505,N_5209);
nand U6085 (N_6085,N_5200,N_5761);
xor U6086 (N_6086,N_5067,N_5959);
or U6087 (N_6087,N_5850,N_5756);
and U6088 (N_6088,N_5875,N_5328);
nor U6089 (N_6089,N_5339,N_5837);
or U6090 (N_6090,N_5010,N_5195);
and U6091 (N_6091,N_5476,N_5855);
and U6092 (N_6092,N_5625,N_5267);
and U6093 (N_6093,N_5659,N_5829);
xnor U6094 (N_6094,N_5358,N_5307);
nor U6095 (N_6095,N_5854,N_5284);
nand U6096 (N_6096,N_5930,N_5050);
nor U6097 (N_6097,N_5889,N_5810);
xnor U6098 (N_6098,N_5784,N_5927);
xnor U6099 (N_6099,N_5263,N_5365);
nand U6100 (N_6100,N_5235,N_5653);
nand U6101 (N_6101,N_5593,N_5495);
or U6102 (N_6102,N_5780,N_5833);
xor U6103 (N_6103,N_5610,N_5891);
nand U6104 (N_6104,N_5720,N_5722);
xor U6105 (N_6105,N_5621,N_5957);
xor U6106 (N_6106,N_5903,N_5310);
and U6107 (N_6107,N_5744,N_5069);
and U6108 (N_6108,N_5678,N_5001);
xor U6109 (N_6109,N_5569,N_5186);
and U6110 (N_6110,N_5513,N_5697);
nand U6111 (N_6111,N_5853,N_5656);
and U6112 (N_6112,N_5557,N_5101);
or U6113 (N_6113,N_5072,N_5666);
xnor U6114 (N_6114,N_5030,N_5698);
xnor U6115 (N_6115,N_5768,N_5692);
and U6116 (N_6116,N_5599,N_5455);
and U6117 (N_6117,N_5897,N_5502);
and U6118 (N_6118,N_5940,N_5672);
nor U6119 (N_6119,N_5617,N_5199);
nor U6120 (N_6120,N_5584,N_5071);
and U6121 (N_6121,N_5304,N_5431);
xor U6122 (N_6122,N_5120,N_5522);
xor U6123 (N_6123,N_5185,N_5594);
nand U6124 (N_6124,N_5982,N_5025);
or U6125 (N_6125,N_5402,N_5226);
xor U6126 (N_6126,N_5138,N_5764);
and U6127 (N_6127,N_5397,N_5690);
xor U6128 (N_6128,N_5322,N_5894);
and U6129 (N_6129,N_5079,N_5969);
nand U6130 (N_6130,N_5393,N_5437);
nand U6131 (N_6131,N_5174,N_5458);
xnor U6132 (N_6132,N_5009,N_5265);
xor U6133 (N_6133,N_5978,N_5113);
xor U6134 (N_6134,N_5876,N_5215);
nand U6135 (N_6135,N_5865,N_5296);
nand U6136 (N_6136,N_5512,N_5813);
nand U6137 (N_6137,N_5511,N_5742);
xor U6138 (N_6138,N_5480,N_5825);
or U6139 (N_6139,N_5667,N_5913);
xor U6140 (N_6140,N_5916,N_5291);
and U6141 (N_6141,N_5933,N_5000);
or U6142 (N_6142,N_5858,N_5799);
xnor U6143 (N_6143,N_5790,N_5413);
xnor U6144 (N_6144,N_5595,N_5005);
nand U6145 (N_6145,N_5160,N_5758);
nand U6146 (N_6146,N_5530,N_5812);
nand U6147 (N_6147,N_5541,N_5173);
nand U6148 (N_6148,N_5081,N_5789);
nor U6149 (N_6149,N_5539,N_5708);
or U6150 (N_6150,N_5964,N_5839);
xnor U6151 (N_6151,N_5939,N_5775);
xnor U6152 (N_6152,N_5577,N_5806);
nand U6153 (N_6153,N_5951,N_5533);
nor U6154 (N_6154,N_5760,N_5862);
nand U6155 (N_6155,N_5439,N_5911);
or U6156 (N_6156,N_5559,N_5293);
xor U6157 (N_6157,N_5326,N_5622);
or U6158 (N_6158,N_5289,N_5410);
and U6159 (N_6159,N_5091,N_5364);
nand U6160 (N_6160,N_5662,N_5095);
xor U6161 (N_6161,N_5117,N_5676);
xor U6162 (N_6162,N_5857,N_5847);
nand U6163 (N_6163,N_5864,N_5872);
or U6164 (N_6164,N_5162,N_5110);
and U6165 (N_6165,N_5154,N_5367);
or U6166 (N_6166,N_5227,N_5257);
nor U6167 (N_6167,N_5273,N_5308);
nand U6168 (N_6168,N_5488,N_5268);
xor U6169 (N_6169,N_5632,N_5677);
or U6170 (N_6170,N_5924,N_5472);
or U6171 (N_6171,N_5256,N_5461);
or U6172 (N_6172,N_5424,N_5554);
nand U6173 (N_6173,N_5242,N_5236);
nand U6174 (N_6174,N_5757,N_5105);
and U6175 (N_6175,N_5246,N_5033);
or U6176 (N_6176,N_5570,N_5486);
nor U6177 (N_6177,N_5028,N_5870);
nor U6178 (N_6178,N_5454,N_5572);
and U6179 (N_6179,N_5316,N_5255);
nand U6180 (N_6180,N_5840,N_5996);
or U6181 (N_6181,N_5918,N_5348);
and U6182 (N_6182,N_5286,N_5968);
and U6183 (N_6183,N_5936,N_5156);
or U6184 (N_6184,N_5024,N_5088);
nand U6185 (N_6185,N_5163,N_5109);
and U6186 (N_6186,N_5211,N_5398);
xor U6187 (N_6187,N_5807,N_5718);
or U6188 (N_6188,N_5036,N_5355);
or U6189 (N_6189,N_5596,N_5018);
and U6190 (N_6190,N_5735,N_5746);
nand U6191 (N_6191,N_5563,N_5890);
or U6192 (N_6192,N_5919,N_5201);
xnor U6193 (N_6193,N_5523,N_5710);
nand U6194 (N_6194,N_5818,N_5491);
xnor U6195 (N_6195,N_5366,N_5886);
and U6196 (N_6196,N_5082,N_5571);
and U6197 (N_6197,N_5647,N_5448);
and U6198 (N_6198,N_5991,N_5315);
nand U6199 (N_6199,N_5483,N_5585);
xor U6200 (N_6200,N_5323,N_5630);
nor U6201 (N_6201,N_5216,N_5130);
nor U6202 (N_6202,N_5543,N_5479);
nor U6203 (N_6203,N_5401,N_5178);
or U6204 (N_6204,N_5992,N_5403);
nor U6205 (N_6205,N_5094,N_5078);
or U6206 (N_6206,N_5100,N_5451);
or U6207 (N_6207,N_5008,N_5576);
or U6208 (N_6208,N_5202,N_5343);
xnor U6209 (N_6209,N_5153,N_5534);
xor U6210 (N_6210,N_5006,N_5298);
nand U6211 (N_6211,N_5386,N_5664);
or U6212 (N_6212,N_5231,N_5925);
and U6213 (N_6213,N_5669,N_5827);
and U6214 (N_6214,N_5650,N_5792);
xor U6215 (N_6215,N_5976,N_5303);
nor U6216 (N_6216,N_5835,N_5145);
or U6217 (N_6217,N_5054,N_5282);
nand U6218 (N_6218,N_5363,N_5808);
or U6219 (N_6219,N_5467,N_5124);
nand U6220 (N_6220,N_5654,N_5507);
nor U6221 (N_6221,N_5558,N_5207);
and U6222 (N_6222,N_5044,N_5443);
nor U6223 (N_6223,N_5759,N_5352);
xnor U6224 (N_6224,N_5869,N_5083);
nor U6225 (N_6225,N_5466,N_5819);
xnor U6226 (N_6226,N_5706,N_5133);
nand U6227 (N_6227,N_5017,N_5682);
and U6228 (N_6228,N_5168,N_5779);
xnor U6229 (N_6229,N_5346,N_5934);
or U6230 (N_6230,N_5064,N_5843);
nor U6231 (N_6231,N_5673,N_5374);
nand U6232 (N_6232,N_5469,N_5212);
nor U6233 (N_6233,N_5527,N_5299);
and U6234 (N_6234,N_5482,N_5824);
or U6235 (N_6235,N_5245,N_5606);
or U6236 (N_6236,N_5449,N_5063);
nor U6237 (N_6237,N_5086,N_5520);
and U6238 (N_6238,N_5204,N_5118);
xnor U6239 (N_6239,N_5058,N_5724);
xnor U6240 (N_6240,N_5762,N_5056);
nor U6241 (N_6241,N_5689,N_5932);
nand U6242 (N_6242,N_5871,N_5016);
nor U6243 (N_6243,N_5128,N_5776);
or U6244 (N_6244,N_5148,N_5732);
xor U6245 (N_6245,N_5440,N_5247);
nand U6246 (N_6246,N_5019,N_5020);
xnor U6247 (N_6247,N_5419,N_5463);
nor U6248 (N_6248,N_5003,N_5140);
nor U6249 (N_6249,N_5749,N_5193);
xor U6250 (N_6250,N_5717,N_5504);
nor U6251 (N_6251,N_5941,N_5222);
nand U6252 (N_6252,N_5013,N_5979);
nand U6253 (N_6253,N_5002,N_5167);
nor U6254 (N_6254,N_5022,N_5369);
or U6255 (N_6255,N_5838,N_5047);
xnor U6256 (N_6256,N_5116,N_5550);
or U6257 (N_6257,N_5217,N_5730);
and U6258 (N_6258,N_5542,N_5997);
xor U6259 (N_6259,N_5040,N_5446);
xnor U6260 (N_6260,N_5498,N_5958);
or U6261 (N_6261,N_5954,N_5531);
nand U6262 (N_6262,N_5442,N_5947);
nand U6263 (N_6263,N_5319,N_5271);
xor U6264 (N_6264,N_5737,N_5910);
xnor U6265 (N_6265,N_5014,N_5191);
nand U6266 (N_6266,N_5125,N_5752);
xnor U6267 (N_6267,N_5070,N_5412);
and U6268 (N_6268,N_5687,N_5132);
xor U6269 (N_6269,N_5516,N_5977);
xor U6270 (N_6270,N_5399,N_5773);
and U6271 (N_6271,N_5210,N_5031);
nand U6272 (N_6272,N_5597,N_5566);
and U6273 (N_6273,N_5716,N_5474);
nand U6274 (N_6274,N_5608,N_5583);
nor U6275 (N_6275,N_5643,N_5092);
nand U6276 (N_6276,N_5763,N_5177);
or U6277 (N_6277,N_5183,N_5826);
and U6278 (N_6278,N_5868,N_5834);
and U6279 (N_6279,N_5360,N_5786);
nor U6280 (N_6280,N_5011,N_5149);
nor U6281 (N_6281,N_5592,N_5152);
or U6282 (N_6282,N_5394,N_5309);
nor U6283 (N_6283,N_5547,N_5179);
xnor U6284 (N_6284,N_5802,N_5526);
and U6285 (N_6285,N_5123,N_5473);
or U6286 (N_6286,N_5699,N_5433);
xor U6287 (N_6287,N_5823,N_5248);
nand U6288 (N_6288,N_5877,N_5312);
nor U6289 (N_6289,N_5026,N_5189);
xnor U6290 (N_6290,N_5801,N_5356);
nor U6291 (N_6291,N_5342,N_5912);
nor U6292 (N_6292,N_5127,N_5785);
nor U6293 (N_6293,N_5956,N_5450);
and U6294 (N_6294,N_5888,N_5990);
nand U6295 (N_6295,N_5863,N_5278);
nand U6296 (N_6296,N_5713,N_5415);
nand U6297 (N_6297,N_5892,N_5651);
or U6298 (N_6298,N_5743,N_5788);
nor U6299 (N_6299,N_5805,N_5464);
nor U6300 (N_6300,N_5143,N_5702);
xnor U6301 (N_6301,N_5261,N_5624);
and U6302 (N_6302,N_5860,N_5234);
and U6303 (N_6303,N_5605,N_5219);
or U6304 (N_6304,N_5301,N_5102);
and U6305 (N_6305,N_5377,N_5613);
xnor U6306 (N_6306,N_5841,N_5580);
xnor U6307 (N_6307,N_5921,N_5338);
and U6308 (N_6308,N_5809,N_5353);
and U6309 (N_6309,N_5965,N_5561);
xor U6310 (N_6310,N_5565,N_5171);
xor U6311 (N_6311,N_5674,N_5230);
nand U6312 (N_6312,N_5305,N_5484);
nand U6313 (N_6313,N_5783,N_5981);
nand U6314 (N_6314,N_5059,N_5734);
or U6315 (N_6315,N_5252,N_5980);
xor U6316 (N_6316,N_5052,N_5896);
and U6317 (N_6317,N_5586,N_5974);
xnor U6318 (N_6318,N_5973,N_5196);
or U6319 (N_6319,N_5368,N_5129);
nor U6320 (N_6320,N_5510,N_5395);
nor U6321 (N_6321,N_5453,N_5141);
and U6322 (N_6322,N_5545,N_5600);
nand U6323 (N_6323,N_5452,N_5514);
or U6324 (N_6324,N_5169,N_5611);
or U6325 (N_6325,N_5727,N_5260);
nand U6326 (N_6326,N_5731,N_5288);
nand U6327 (N_6327,N_5998,N_5384);
nor U6328 (N_6328,N_5279,N_5618);
nor U6329 (N_6329,N_5638,N_5695);
or U6330 (N_6330,N_5668,N_5509);
nor U6331 (N_6331,N_5385,N_5553);
or U6332 (N_6332,N_5378,N_5387);
xnor U6333 (N_6333,N_5112,N_5637);
or U6334 (N_6334,N_5842,N_5049);
nor U6335 (N_6335,N_5867,N_5400);
and U6336 (N_6336,N_5175,N_5815);
nor U6337 (N_6337,N_5700,N_5349);
or U6338 (N_6338,N_5844,N_5239);
xor U6339 (N_6339,N_5161,N_5444);
nor U6340 (N_6340,N_5811,N_5670);
xnor U6341 (N_6341,N_5928,N_5496);
xor U6342 (N_6342,N_5615,N_5259);
nor U6343 (N_6343,N_5568,N_5831);
or U6344 (N_6344,N_5614,N_5852);
xnor U6345 (N_6345,N_5640,N_5396);
nor U6346 (N_6346,N_5601,N_5885);
xnor U6347 (N_6347,N_5462,N_5057);
xor U6348 (N_6348,N_5053,N_5314);
or U6349 (N_6349,N_5158,N_5960);
nand U6350 (N_6350,N_5029,N_5430);
or U6351 (N_6351,N_5297,N_5249);
nand U6352 (N_6352,N_5694,N_5642);
nand U6353 (N_6353,N_5084,N_5240);
or U6354 (N_6354,N_5076,N_5223);
or U6355 (N_6355,N_5616,N_5893);
or U6356 (N_6356,N_5777,N_5205);
nand U6357 (N_6357,N_5946,N_5901);
nand U6358 (N_6358,N_5719,N_5987);
and U6359 (N_6359,N_5535,N_5920);
xnor U6360 (N_6360,N_5683,N_5213);
nor U6361 (N_6361,N_5705,N_5880);
xor U6362 (N_6362,N_5429,N_5733);
xor U6363 (N_6363,N_5283,N_5165);
and U6364 (N_6364,N_5492,N_5736);
and U6365 (N_6365,N_5848,N_5688);
xor U6366 (N_6366,N_5347,N_5073);
and U6367 (N_6367,N_5287,N_5851);
or U6368 (N_6368,N_5045,N_5441);
nand U6369 (N_6369,N_5391,N_5908);
nor U6370 (N_6370,N_5475,N_5122);
or U6371 (N_6371,N_5150,N_5942);
xor U6372 (N_6372,N_5329,N_5325);
nor U6373 (N_6373,N_5276,N_5602);
xor U6374 (N_6374,N_5729,N_5336);
nand U6375 (N_6375,N_5266,N_5626);
or U6376 (N_6376,N_5035,N_5627);
or U6377 (N_6377,N_5646,N_5988);
or U6378 (N_6378,N_5791,N_5975);
and U6379 (N_6379,N_5769,N_5350);
or U6380 (N_6380,N_5447,N_5164);
nand U6381 (N_6381,N_5995,N_5814);
nor U6382 (N_6382,N_5712,N_5907);
and U6383 (N_6383,N_5241,N_5587);
nor U6384 (N_6384,N_5633,N_5324);
nor U6385 (N_6385,N_5665,N_5389);
nand U6386 (N_6386,N_5414,N_5061);
xor U6387 (N_6387,N_5798,N_5537);
or U6388 (N_6388,N_5817,N_5816);
or U6389 (N_6389,N_5182,N_5800);
nand U6390 (N_6390,N_5218,N_5272);
or U6391 (N_6391,N_5136,N_5142);
xor U6392 (N_6392,N_5846,N_5984);
nor U6393 (N_6393,N_5909,N_5075);
nand U6394 (N_6394,N_5221,N_5172);
and U6395 (N_6395,N_5270,N_5065);
nor U6396 (N_6396,N_5380,N_5383);
nor U6397 (N_6397,N_5887,N_5404);
nand U6398 (N_6398,N_5157,N_5715);
or U6399 (N_6399,N_5709,N_5477);
nand U6400 (N_6400,N_5952,N_5772);
nor U6401 (N_6401,N_5264,N_5655);
nand U6402 (N_6402,N_5370,N_5335);
nor U6403 (N_6403,N_5787,N_5765);
xor U6404 (N_6404,N_5922,N_5362);
or U6405 (N_6405,N_5684,N_5629);
or U6406 (N_6406,N_5905,N_5376);
nor U6407 (N_6407,N_5657,N_5192);
or U6408 (N_6408,N_5423,N_5794);
nor U6409 (N_6409,N_5292,N_5745);
and U6410 (N_6410,N_5508,N_5098);
xor U6411 (N_6411,N_5972,N_5739);
xnor U6412 (N_6412,N_5598,N_5866);
or U6413 (N_6413,N_5728,N_5500);
nand U6414 (N_6414,N_5796,N_5337);
nor U6415 (N_6415,N_5714,N_5675);
xor U6416 (N_6416,N_5658,N_5214);
nand U6417 (N_6417,N_5007,N_5037);
or U6418 (N_6418,N_5652,N_5931);
and U6419 (N_6419,N_5190,N_5536);
nor U6420 (N_6420,N_5926,N_5711);
or U6421 (N_6421,N_5357,N_5751);
xnor U6422 (N_6422,N_5999,N_5704);
nor U6423 (N_6423,N_5436,N_5093);
nor U6424 (N_6424,N_5341,N_5197);
and U6425 (N_6425,N_5229,N_5793);
and U6426 (N_6426,N_5723,N_5405);
xnor U6427 (N_6427,N_5878,N_5159);
or U6428 (N_6428,N_5771,N_5220);
and U6429 (N_6429,N_5187,N_5051);
or U6430 (N_6430,N_5225,N_5938);
or U6431 (N_6431,N_5660,N_5490);
nor U6432 (N_6432,N_5277,N_5115);
nor U6433 (N_6433,N_5198,N_5929);
nand U6434 (N_6434,N_5478,N_5494);
nor U6435 (N_6435,N_5881,N_5188);
nand U6436 (N_6436,N_5636,N_5332);
xor U6437 (N_6437,N_5489,N_5883);
nor U6438 (N_6438,N_5275,N_5874);
xor U6439 (N_6439,N_5879,N_5645);
and U6440 (N_6440,N_5354,N_5253);
or U6441 (N_6441,N_5428,N_5206);
nor U6442 (N_6442,N_5943,N_5575);
xnor U6443 (N_6443,N_5233,N_5726);
nor U6444 (N_6444,N_5953,N_5493);
nand U6445 (N_6445,N_5914,N_5023);
or U6446 (N_6446,N_5435,N_5317);
nor U6447 (N_6447,N_5649,N_5238);
and U6448 (N_6448,N_5459,N_5770);
and U6449 (N_6449,N_5607,N_5528);
and U6450 (N_6450,N_5371,N_5915);
nor U6451 (N_6451,N_5390,N_5519);
or U6452 (N_6452,N_5166,N_5820);
xor U6453 (N_6453,N_5634,N_5685);
or U6454 (N_6454,N_5146,N_5126);
and U6455 (N_6455,N_5321,N_5501);
nand U6456 (N_6456,N_5274,N_5748);
xnor U6457 (N_6457,N_5411,N_5538);
nor U6458 (N_6458,N_5333,N_5041);
nand U6459 (N_6459,N_5628,N_5432);
or U6460 (N_6460,N_5803,N_5552);
and U6461 (N_6461,N_5250,N_5421);
nor U6462 (N_6462,N_5407,N_5313);
xor U6463 (N_6463,N_5503,N_5038);
nor U6464 (N_6464,N_5499,N_5176);
nand U6465 (N_6465,N_5155,N_5034);
nand U6466 (N_6466,N_5042,N_5104);
or U6467 (N_6467,N_5882,N_5381);
or U6468 (N_6468,N_5631,N_5578);
and U6469 (N_6469,N_5590,N_5945);
or U6470 (N_6470,N_5696,N_5012);
or U6471 (N_6471,N_5438,N_5184);
nor U6472 (N_6472,N_5573,N_5983);
nor U6473 (N_6473,N_5644,N_5767);
nor U6474 (N_6474,N_5295,N_5021);
and U6475 (N_6475,N_5873,N_5345);
xnor U6476 (N_6476,N_5097,N_5970);
nand U6477 (N_6477,N_5663,N_5555);
xnor U6478 (N_6478,N_5497,N_5320);
and U6479 (N_6479,N_5521,N_5579);
and U6480 (N_6480,N_5738,N_5487);
nor U6481 (N_6481,N_5066,N_5243);
or U6482 (N_6482,N_5062,N_5518);
xnor U6483 (N_6483,N_5302,N_5103);
or U6484 (N_6484,N_5619,N_5567);
nand U6485 (N_6485,N_5470,N_5582);
nor U6486 (N_6486,N_5604,N_5409);
or U6487 (N_6487,N_5085,N_5043);
nand U6488 (N_6488,N_5375,N_5372);
and U6489 (N_6489,N_5068,N_5755);
nor U6490 (N_6490,N_5046,N_5900);
nor U6491 (N_6491,N_5048,N_5962);
or U6492 (N_6492,N_5285,N_5725);
or U6493 (N_6493,N_5131,N_5460);
nand U6494 (N_6494,N_5546,N_5635);
and U6495 (N_6495,N_5228,N_5581);
or U6496 (N_6496,N_5434,N_5406);
xnor U6497 (N_6497,N_5359,N_5420);
nor U6498 (N_6498,N_5294,N_5388);
or U6499 (N_6499,N_5661,N_5971);
xor U6500 (N_6500,N_5936,N_5115);
or U6501 (N_6501,N_5143,N_5734);
and U6502 (N_6502,N_5949,N_5719);
nor U6503 (N_6503,N_5943,N_5664);
nor U6504 (N_6504,N_5861,N_5800);
and U6505 (N_6505,N_5238,N_5732);
xnor U6506 (N_6506,N_5350,N_5217);
nand U6507 (N_6507,N_5815,N_5287);
nand U6508 (N_6508,N_5192,N_5737);
or U6509 (N_6509,N_5344,N_5753);
nand U6510 (N_6510,N_5980,N_5236);
nand U6511 (N_6511,N_5066,N_5939);
or U6512 (N_6512,N_5936,N_5043);
xor U6513 (N_6513,N_5136,N_5645);
xor U6514 (N_6514,N_5292,N_5419);
nand U6515 (N_6515,N_5516,N_5183);
nor U6516 (N_6516,N_5791,N_5820);
xor U6517 (N_6517,N_5332,N_5415);
or U6518 (N_6518,N_5348,N_5526);
and U6519 (N_6519,N_5546,N_5619);
or U6520 (N_6520,N_5635,N_5041);
or U6521 (N_6521,N_5555,N_5928);
nand U6522 (N_6522,N_5898,N_5878);
or U6523 (N_6523,N_5804,N_5875);
nor U6524 (N_6524,N_5910,N_5719);
xor U6525 (N_6525,N_5605,N_5189);
xor U6526 (N_6526,N_5403,N_5305);
nor U6527 (N_6527,N_5337,N_5243);
xor U6528 (N_6528,N_5030,N_5421);
xor U6529 (N_6529,N_5360,N_5457);
nor U6530 (N_6530,N_5714,N_5629);
nor U6531 (N_6531,N_5579,N_5219);
nand U6532 (N_6532,N_5390,N_5541);
or U6533 (N_6533,N_5588,N_5553);
and U6534 (N_6534,N_5019,N_5201);
nand U6535 (N_6535,N_5396,N_5794);
and U6536 (N_6536,N_5031,N_5695);
nor U6537 (N_6537,N_5181,N_5724);
nand U6538 (N_6538,N_5093,N_5584);
nand U6539 (N_6539,N_5135,N_5339);
or U6540 (N_6540,N_5494,N_5134);
xnor U6541 (N_6541,N_5204,N_5751);
or U6542 (N_6542,N_5308,N_5612);
nor U6543 (N_6543,N_5695,N_5572);
xor U6544 (N_6544,N_5901,N_5922);
nand U6545 (N_6545,N_5132,N_5857);
xnor U6546 (N_6546,N_5620,N_5274);
and U6547 (N_6547,N_5005,N_5235);
nor U6548 (N_6548,N_5320,N_5890);
nor U6549 (N_6549,N_5959,N_5938);
nor U6550 (N_6550,N_5957,N_5099);
and U6551 (N_6551,N_5350,N_5279);
nor U6552 (N_6552,N_5445,N_5073);
nor U6553 (N_6553,N_5168,N_5225);
nand U6554 (N_6554,N_5067,N_5760);
nor U6555 (N_6555,N_5887,N_5085);
or U6556 (N_6556,N_5247,N_5621);
nand U6557 (N_6557,N_5967,N_5599);
and U6558 (N_6558,N_5270,N_5424);
nor U6559 (N_6559,N_5477,N_5943);
xor U6560 (N_6560,N_5477,N_5929);
nand U6561 (N_6561,N_5898,N_5104);
and U6562 (N_6562,N_5202,N_5264);
or U6563 (N_6563,N_5115,N_5673);
nand U6564 (N_6564,N_5514,N_5101);
xnor U6565 (N_6565,N_5527,N_5106);
and U6566 (N_6566,N_5197,N_5595);
nor U6567 (N_6567,N_5365,N_5646);
nand U6568 (N_6568,N_5570,N_5508);
xnor U6569 (N_6569,N_5089,N_5082);
or U6570 (N_6570,N_5617,N_5233);
xor U6571 (N_6571,N_5394,N_5729);
or U6572 (N_6572,N_5668,N_5174);
nor U6573 (N_6573,N_5436,N_5857);
nand U6574 (N_6574,N_5937,N_5566);
and U6575 (N_6575,N_5551,N_5165);
or U6576 (N_6576,N_5688,N_5871);
nor U6577 (N_6577,N_5178,N_5652);
xor U6578 (N_6578,N_5491,N_5829);
or U6579 (N_6579,N_5953,N_5480);
xnor U6580 (N_6580,N_5350,N_5851);
nand U6581 (N_6581,N_5292,N_5337);
xor U6582 (N_6582,N_5969,N_5315);
xnor U6583 (N_6583,N_5080,N_5592);
xnor U6584 (N_6584,N_5730,N_5095);
or U6585 (N_6585,N_5613,N_5669);
nor U6586 (N_6586,N_5064,N_5377);
or U6587 (N_6587,N_5855,N_5614);
xor U6588 (N_6588,N_5743,N_5953);
nand U6589 (N_6589,N_5235,N_5165);
nand U6590 (N_6590,N_5916,N_5617);
nand U6591 (N_6591,N_5699,N_5378);
xnor U6592 (N_6592,N_5549,N_5096);
nor U6593 (N_6593,N_5243,N_5463);
nand U6594 (N_6594,N_5716,N_5101);
nand U6595 (N_6595,N_5235,N_5617);
or U6596 (N_6596,N_5808,N_5312);
nand U6597 (N_6597,N_5533,N_5600);
nor U6598 (N_6598,N_5301,N_5863);
and U6599 (N_6599,N_5304,N_5986);
or U6600 (N_6600,N_5800,N_5863);
nor U6601 (N_6601,N_5328,N_5118);
or U6602 (N_6602,N_5831,N_5587);
xnor U6603 (N_6603,N_5541,N_5032);
nand U6604 (N_6604,N_5650,N_5253);
or U6605 (N_6605,N_5634,N_5049);
nand U6606 (N_6606,N_5766,N_5399);
and U6607 (N_6607,N_5720,N_5482);
xor U6608 (N_6608,N_5784,N_5306);
nand U6609 (N_6609,N_5148,N_5061);
and U6610 (N_6610,N_5861,N_5234);
nand U6611 (N_6611,N_5258,N_5958);
xor U6612 (N_6612,N_5796,N_5374);
and U6613 (N_6613,N_5946,N_5971);
nor U6614 (N_6614,N_5393,N_5481);
and U6615 (N_6615,N_5805,N_5976);
and U6616 (N_6616,N_5185,N_5169);
and U6617 (N_6617,N_5772,N_5620);
xor U6618 (N_6618,N_5162,N_5145);
nor U6619 (N_6619,N_5854,N_5061);
and U6620 (N_6620,N_5373,N_5179);
xor U6621 (N_6621,N_5927,N_5216);
xnor U6622 (N_6622,N_5633,N_5934);
xnor U6623 (N_6623,N_5168,N_5488);
or U6624 (N_6624,N_5103,N_5499);
or U6625 (N_6625,N_5554,N_5675);
nor U6626 (N_6626,N_5016,N_5711);
nand U6627 (N_6627,N_5032,N_5818);
nand U6628 (N_6628,N_5251,N_5263);
nor U6629 (N_6629,N_5914,N_5619);
nand U6630 (N_6630,N_5440,N_5707);
and U6631 (N_6631,N_5963,N_5018);
nor U6632 (N_6632,N_5419,N_5265);
xnor U6633 (N_6633,N_5653,N_5565);
xor U6634 (N_6634,N_5469,N_5109);
nand U6635 (N_6635,N_5094,N_5118);
and U6636 (N_6636,N_5481,N_5489);
nor U6637 (N_6637,N_5226,N_5670);
or U6638 (N_6638,N_5033,N_5512);
xor U6639 (N_6639,N_5120,N_5325);
nor U6640 (N_6640,N_5841,N_5072);
nand U6641 (N_6641,N_5929,N_5377);
xor U6642 (N_6642,N_5828,N_5546);
nand U6643 (N_6643,N_5047,N_5833);
nand U6644 (N_6644,N_5723,N_5910);
or U6645 (N_6645,N_5529,N_5688);
xnor U6646 (N_6646,N_5112,N_5852);
nand U6647 (N_6647,N_5670,N_5294);
or U6648 (N_6648,N_5617,N_5970);
nand U6649 (N_6649,N_5116,N_5344);
nor U6650 (N_6650,N_5781,N_5670);
xor U6651 (N_6651,N_5062,N_5816);
nand U6652 (N_6652,N_5582,N_5884);
or U6653 (N_6653,N_5326,N_5232);
and U6654 (N_6654,N_5580,N_5341);
nand U6655 (N_6655,N_5216,N_5967);
and U6656 (N_6656,N_5217,N_5222);
or U6657 (N_6657,N_5270,N_5585);
nand U6658 (N_6658,N_5461,N_5148);
or U6659 (N_6659,N_5546,N_5960);
or U6660 (N_6660,N_5633,N_5836);
and U6661 (N_6661,N_5250,N_5591);
or U6662 (N_6662,N_5886,N_5792);
nor U6663 (N_6663,N_5681,N_5796);
xnor U6664 (N_6664,N_5727,N_5776);
xor U6665 (N_6665,N_5634,N_5586);
nor U6666 (N_6666,N_5028,N_5720);
or U6667 (N_6667,N_5019,N_5128);
xnor U6668 (N_6668,N_5444,N_5976);
or U6669 (N_6669,N_5122,N_5730);
nand U6670 (N_6670,N_5249,N_5762);
and U6671 (N_6671,N_5271,N_5138);
or U6672 (N_6672,N_5713,N_5569);
or U6673 (N_6673,N_5237,N_5012);
nor U6674 (N_6674,N_5893,N_5921);
or U6675 (N_6675,N_5844,N_5678);
xor U6676 (N_6676,N_5260,N_5068);
or U6677 (N_6677,N_5190,N_5458);
and U6678 (N_6678,N_5581,N_5485);
xor U6679 (N_6679,N_5298,N_5093);
xor U6680 (N_6680,N_5279,N_5824);
nor U6681 (N_6681,N_5504,N_5468);
nor U6682 (N_6682,N_5983,N_5777);
xor U6683 (N_6683,N_5237,N_5535);
and U6684 (N_6684,N_5600,N_5133);
xnor U6685 (N_6685,N_5567,N_5736);
or U6686 (N_6686,N_5368,N_5916);
or U6687 (N_6687,N_5306,N_5436);
nor U6688 (N_6688,N_5639,N_5396);
nor U6689 (N_6689,N_5935,N_5722);
xnor U6690 (N_6690,N_5710,N_5992);
xnor U6691 (N_6691,N_5500,N_5413);
nand U6692 (N_6692,N_5729,N_5731);
and U6693 (N_6693,N_5418,N_5241);
xnor U6694 (N_6694,N_5440,N_5762);
or U6695 (N_6695,N_5967,N_5758);
xnor U6696 (N_6696,N_5653,N_5872);
or U6697 (N_6697,N_5951,N_5261);
nor U6698 (N_6698,N_5098,N_5555);
nand U6699 (N_6699,N_5537,N_5931);
nand U6700 (N_6700,N_5841,N_5009);
or U6701 (N_6701,N_5632,N_5404);
and U6702 (N_6702,N_5554,N_5261);
or U6703 (N_6703,N_5101,N_5728);
nand U6704 (N_6704,N_5716,N_5661);
xor U6705 (N_6705,N_5757,N_5661);
or U6706 (N_6706,N_5335,N_5617);
nand U6707 (N_6707,N_5631,N_5327);
or U6708 (N_6708,N_5823,N_5408);
nor U6709 (N_6709,N_5509,N_5539);
xor U6710 (N_6710,N_5588,N_5904);
nor U6711 (N_6711,N_5264,N_5642);
nor U6712 (N_6712,N_5106,N_5736);
and U6713 (N_6713,N_5087,N_5603);
xor U6714 (N_6714,N_5630,N_5230);
nor U6715 (N_6715,N_5895,N_5605);
nand U6716 (N_6716,N_5127,N_5310);
and U6717 (N_6717,N_5930,N_5615);
nand U6718 (N_6718,N_5554,N_5384);
nand U6719 (N_6719,N_5591,N_5103);
nand U6720 (N_6720,N_5591,N_5316);
nor U6721 (N_6721,N_5684,N_5033);
and U6722 (N_6722,N_5987,N_5606);
xor U6723 (N_6723,N_5592,N_5260);
or U6724 (N_6724,N_5427,N_5141);
nor U6725 (N_6725,N_5969,N_5722);
nand U6726 (N_6726,N_5113,N_5645);
or U6727 (N_6727,N_5388,N_5485);
and U6728 (N_6728,N_5110,N_5452);
nand U6729 (N_6729,N_5848,N_5678);
xnor U6730 (N_6730,N_5732,N_5301);
xnor U6731 (N_6731,N_5008,N_5598);
xor U6732 (N_6732,N_5589,N_5535);
xor U6733 (N_6733,N_5485,N_5817);
xor U6734 (N_6734,N_5270,N_5917);
nor U6735 (N_6735,N_5486,N_5383);
nor U6736 (N_6736,N_5152,N_5165);
and U6737 (N_6737,N_5093,N_5522);
or U6738 (N_6738,N_5380,N_5872);
xnor U6739 (N_6739,N_5416,N_5160);
or U6740 (N_6740,N_5696,N_5951);
nand U6741 (N_6741,N_5359,N_5457);
xor U6742 (N_6742,N_5336,N_5545);
and U6743 (N_6743,N_5488,N_5257);
xnor U6744 (N_6744,N_5794,N_5250);
or U6745 (N_6745,N_5645,N_5942);
or U6746 (N_6746,N_5752,N_5875);
or U6747 (N_6747,N_5186,N_5112);
or U6748 (N_6748,N_5250,N_5708);
nor U6749 (N_6749,N_5561,N_5667);
nor U6750 (N_6750,N_5182,N_5257);
or U6751 (N_6751,N_5706,N_5104);
xnor U6752 (N_6752,N_5953,N_5592);
nor U6753 (N_6753,N_5139,N_5640);
xnor U6754 (N_6754,N_5301,N_5896);
nand U6755 (N_6755,N_5545,N_5669);
nor U6756 (N_6756,N_5108,N_5763);
and U6757 (N_6757,N_5018,N_5586);
xnor U6758 (N_6758,N_5029,N_5823);
nor U6759 (N_6759,N_5798,N_5564);
and U6760 (N_6760,N_5002,N_5201);
nand U6761 (N_6761,N_5409,N_5690);
nor U6762 (N_6762,N_5442,N_5148);
nor U6763 (N_6763,N_5128,N_5147);
xor U6764 (N_6764,N_5026,N_5042);
xor U6765 (N_6765,N_5049,N_5880);
or U6766 (N_6766,N_5935,N_5801);
nor U6767 (N_6767,N_5997,N_5791);
nand U6768 (N_6768,N_5710,N_5365);
or U6769 (N_6769,N_5696,N_5425);
xnor U6770 (N_6770,N_5477,N_5765);
nand U6771 (N_6771,N_5053,N_5711);
nor U6772 (N_6772,N_5165,N_5968);
nand U6773 (N_6773,N_5092,N_5809);
nor U6774 (N_6774,N_5843,N_5308);
nand U6775 (N_6775,N_5942,N_5625);
and U6776 (N_6776,N_5917,N_5409);
and U6777 (N_6777,N_5031,N_5668);
or U6778 (N_6778,N_5224,N_5790);
or U6779 (N_6779,N_5411,N_5802);
xnor U6780 (N_6780,N_5654,N_5233);
nand U6781 (N_6781,N_5391,N_5060);
nor U6782 (N_6782,N_5989,N_5019);
nand U6783 (N_6783,N_5299,N_5147);
nand U6784 (N_6784,N_5254,N_5927);
nand U6785 (N_6785,N_5570,N_5242);
and U6786 (N_6786,N_5659,N_5054);
and U6787 (N_6787,N_5772,N_5118);
xnor U6788 (N_6788,N_5149,N_5489);
nand U6789 (N_6789,N_5419,N_5062);
or U6790 (N_6790,N_5447,N_5967);
nand U6791 (N_6791,N_5591,N_5453);
nor U6792 (N_6792,N_5317,N_5227);
or U6793 (N_6793,N_5608,N_5885);
nand U6794 (N_6794,N_5388,N_5646);
or U6795 (N_6795,N_5738,N_5423);
or U6796 (N_6796,N_5168,N_5938);
or U6797 (N_6797,N_5755,N_5326);
and U6798 (N_6798,N_5224,N_5593);
xnor U6799 (N_6799,N_5682,N_5492);
xnor U6800 (N_6800,N_5566,N_5343);
or U6801 (N_6801,N_5441,N_5024);
or U6802 (N_6802,N_5052,N_5950);
or U6803 (N_6803,N_5884,N_5033);
nor U6804 (N_6804,N_5318,N_5651);
xor U6805 (N_6805,N_5091,N_5990);
nand U6806 (N_6806,N_5230,N_5957);
xnor U6807 (N_6807,N_5454,N_5098);
xnor U6808 (N_6808,N_5755,N_5454);
or U6809 (N_6809,N_5163,N_5433);
nand U6810 (N_6810,N_5503,N_5762);
or U6811 (N_6811,N_5299,N_5737);
and U6812 (N_6812,N_5910,N_5888);
xnor U6813 (N_6813,N_5630,N_5189);
xor U6814 (N_6814,N_5511,N_5529);
nand U6815 (N_6815,N_5611,N_5052);
xnor U6816 (N_6816,N_5420,N_5791);
xnor U6817 (N_6817,N_5876,N_5816);
nor U6818 (N_6818,N_5462,N_5345);
nand U6819 (N_6819,N_5914,N_5044);
nor U6820 (N_6820,N_5705,N_5726);
or U6821 (N_6821,N_5500,N_5409);
nor U6822 (N_6822,N_5444,N_5574);
nand U6823 (N_6823,N_5522,N_5946);
and U6824 (N_6824,N_5351,N_5454);
and U6825 (N_6825,N_5969,N_5239);
and U6826 (N_6826,N_5900,N_5931);
xnor U6827 (N_6827,N_5101,N_5634);
nand U6828 (N_6828,N_5262,N_5308);
nor U6829 (N_6829,N_5010,N_5899);
and U6830 (N_6830,N_5653,N_5688);
and U6831 (N_6831,N_5287,N_5559);
xnor U6832 (N_6832,N_5322,N_5851);
xor U6833 (N_6833,N_5323,N_5539);
xnor U6834 (N_6834,N_5249,N_5059);
or U6835 (N_6835,N_5410,N_5653);
nor U6836 (N_6836,N_5366,N_5248);
nor U6837 (N_6837,N_5422,N_5640);
nand U6838 (N_6838,N_5811,N_5606);
and U6839 (N_6839,N_5908,N_5954);
or U6840 (N_6840,N_5569,N_5807);
and U6841 (N_6841,N_5870,N_5621);
nor U6842 (N_6842,N_5011,N_5929);
xnor U6843 (N_6843,N_5577,N_5674);
and U6844 (N_6844,N_5687,N_5967);
or U6845 (N_6845,N_5615,N_5699);
and U6846 (N_6846,N_5752,N_5282);
xnor U6847 (N_6847,N_5280,N_5651);
xnor U6848 (N_6848,N_5778,N_5352);
and U6849 (N_6849,N_5006,N_5026);
and U6850 (N_6850,N_5487,N_5632);
and U6851 (N_6851,N_5008,N_5092);
and U6852 (N_6852,N_5549,N_5985);
or U6853 (N_6853,N_5500,N_5862);
or U6854 (N_6854,N_5303,N_5491);
and U6855 (N_6855,N_5335,N_5754);
nor U6856 (N_6856,N_5470,N_5824);
xnor U6857 (N_6857,N_5066,N_5200);
or U6858 (N_6858,N_5732,N_5645);
nand U6859 (N_6859,N_5469,N_5987);
xnor U6860 (N_6860,N_5122,N_5703);
and U6861 (N_6861,N_5339,N_5280);
and U6862 (N_6862,N_5631,N_5535);
nand U6863 (N_6863,N_5690,N_5561);
nor U6864 (N_6864,N_5631,N_5719);
xor U6865 (N_6865,N_5882,N_5705);
or U6866 (N_6866,N_5384,N_5398);
and U6867 (N_6867,N_5724,N_5525);
nor U6868 (N_6868,N_5524,N_5362);
nor U6869 (N_6869,N_5145,N_5460);
or U6870 (N_6870,N_5406,N_5421);
or U6871 (N_6871,N_5943,N_5022);
nor U6872 (N_6872,N_5490,N_5925);
nor U6873 (N_6873,N_5278,N_5660);
or U6874 (N_6874,N_5674,N_5306);
and U6875 (N_6875,N_5606,N_5503);
nor U6876 (N_6876,N_5186,N_5901);
nand U6877 (N_6877,N_5614,N_5080);
and U6878 (N_6878,N_5279,N_5321);
nor U6879 (N_6879,N_5023,N_5261);
or U6880 (N_6880,N_5285,N_5568);
nand U6881 (N_6881,N_5153,N_5150);
and U6882 (N_6882,N_5163,N_5655);
nand U6883 (N_6883,N_5456,N_5334);
xnor U6884 (N_6884,N_5978,N_5642);
xnor U6885 (N_6885,N_5031,N_5864);
and U6886 (N_6886,N_5422,N_5141);
nand U6887 (N_6887,N_5502,N_5190);
nor U6888 (N_6888,N_5272,N_5327);
nand U6889 (N_6889,N_5712,N_5604);
xor U6890 (N_6890,N_5519,N_5281);
nor U6891 (N_6891,N_5922,N_5033);
xor U6892 (N_6892,N_5862,N_5884);
and U6893 (N_6893,N_5183,N_5836);
and U6894 (N_6894,N_5308,N_5647);
and U6895 (N_6895,N_5500,N_5819);
nand U6896 (N_6896,N_5608,N_5680);
nor U6897 (N_6897,N_5181,N_5029);
nor U6898 (N_6898,N_5482,N_5881);
nor U6899 (N_6899,N_5678,N_5100);
and U6900 (N_6900,N_5459,N_5581);
nand U6901 (N_6901,N_5868,N_5911);
and U6902 (N_6902,N_5483,N_5008);
nor U6903 (N_6903,N_5525,N_5318);
nand U6904 (N_6904,N_5852,N_5861);
or U6905 (N_6905,N_5251,N_5647);
xnor U6906 (N_6906,N_5387,N_5503);
xnor U6907 (N_6907,N_5514,N_5941);
nor U6908 (N_6908,N_5941,N_5424);
or U6909 (N_6909,N_5175,N_5499);
and U6910 (N_6910,N_5371,N_5443);
nor U6911 (N_6911,N_5193,N_5890);
and U6912 (N_6912,N_5834,N_5311);
xor U6913 (N_6913,N_5371,N_5409);
nor U6914 (N_6914,N_5976,N_5851);
or U6915 (N_6915,N_5199,N_5278);
xnor U6916 (N_6916,N_5612,N_5391);
nand U6917 (N_6917,N_5518,N_5138);
nand U6918 (N_6918,N_5589,N_5877);
or U6919 (N_6919,N_5053,N_5767);
xor U6920 (N_6920,N_5832,N_5796);
and U6921 (N_6921,N_5717,N_5175);
or U6922 (N_6922,N_5333,N_5967);
and U6923 (N_6923,N_5024,N_5822);
nor U6924 (N_6924,N_5334,N_5350);
and U6925 (N_6925,N_5175,N_5406);
and U6926 (N_6926,N_5313,N_5717);
nor U6927 (N_6927,N_5779,N_5726);
nand U6928 (N_6928,N_5556,N_5857);
nor U6929 (N_6929,N_5072,N_5078);
and U6930 (N_6930,N_5050,N_5343);
and U6931 (N_6931,N_5942,N_5749);
or U6932 (N_6932,N_5154,N_5388);
and U6933 (N_6933,N_5048,N_5357);
and U6934 (N_6934,N_5303,N_5857);
and U6935 (N_6935,N_5997,N_5490);
or U6936 (N_6936,N_5510,N_5268);
or U6937 (N_6937,N_5549,N_5810);
and U6938 (N_6938,N_5530,N_5782);
nand U6939 (N_6939,N_5387,N_5766);
or U6940 (N_6940,N_5628,N_5134);
nor U6941 (N_6941,N_5872,N_5771);
nor U6942 (N_6942,N_5405,N_5091);
xnor U6943 (N_6943,N_5502,N_5064);
or U6944 (N_6944,N_5857,N_5767);
and U6945 (N_6945,N_5175,N_5006);
or U6946 (N_6946,N_5508,N_5433);
xor U6947 (N_6947,N_5552,N_5061);
nand U6948 (N_6948,N_5687,N_5983);
and U6949 (N_6949,N_5129,N_5557);
nor U6950 (N_6950,N_5917,N_5783);
nor U6951 (N_6951,N_5264,N_5379);
nor U6952 (N_6952,N_5527,N_5176);
nor U6953 (N_6953,N_5870,N_5798);
nor U6954 (N_6954,N_5483,N_5454);
nand U6955 (N_6955,N_5606,N_5937);
nor U6956 (N_6956,N_5823,N_5152);
nor U6957 (N_6957,N_5737,N_5042);
nand U6958 (N_6958,N_5532,N_5998);
nand U6959 (N_6959,N_5975,N_5802);
nor U6960 (N_6960,N_5147,N_5627);
and U6961 (N_6961,N_5402,N_5244);
and U6962 (N_6962,N_5762,N_5775);
and U6963 (N_6963,N_5862,N_5299);
nand U6964 (N_6964,N_5116,N_5531);
or U6965 (N_6965,N_5478,N_5899);
nor U6966 (N_6966,N_5323,N_5641);
and U6967 (N_6967,N_5609,N_5752);
nand U6968 (N_6968,N_5145,N_5186);
xnor U6969 (N_6969,N_5333,N_5170);
and U6970 (N_6970,N_5056,N_5815);
nand U6971 (N_6971,N_5232,N_5441);
nor U6972 (N_6972,N_5257,N_5713);
and U6973 (N_6973,N_5063,N_5656);
and U6974 (N_6974,N_5337,N_5553);
and U6975 (N_6975,N_5621,N_5718);
nand U6976 (N_6976,N_5319,N_5010);
or U6977 (N_6977,N_5779,N_5197);
nand U6978 (N_6978,N_5595,N_5427);
xor U6979 (N_6979,N_5972,N_5647);
and U6980 (N_6980,N_5583,N_5814);
or U6981 (N_6981,N_5378,N_5800);
or U6982 (N_6982,N_5870,N_5861);
or U6983 (N_6983,N_5755,N_5318);
or U6984 (N_6984,N_5508,N_5763);
nand U6985 (N_6985,N_5872,N_5748);
nand U6986 (N_6986,N_5514,N_5047);
nand U6987 (N_6987,N_5320,N_5823);
nand U6988 (N_6988,N_5609,N_5870);
or U6989 (N_6989,N_5969,N_5283);
xor U6990 (N_6990,N_5930,N_5020);
nor U6991 (N_6991,N_5274,N_5405);
nor U6992 (N_6992,N_5388,N_5352);
nand U6993 (N_6993,N_5893,N_5872);
or U6994 (N_6994,N_5928,N_5825);
and U6995 (N_6995,N_5867,N_5013);
or U6996 (N_6996,N_5778,N_5073);
or U6997 (N_6997,N_5695,N_5759);
nand U6998 (N_6998,N_5082,N_5132);
nor U6999 (N_6999,N_5969,N_5349);
nor U7000 (N_7000,N_6793,N_6802);
xnor U7001 (N_7001,N_6570,N_6038);
xor U7002 (N_7002,N_6792,N_6691);
xnor U7003 (N_7003,N_6550,N_6747);
or U7004 (N_7004,N_6982,N_6578);
or U7005 (N_7005,N_6696,N_6619);
nor U7006 (N_7006,N_6751,N_6139);
and U7007 (N_7007,N_6147,N_6315);
nor U7008 (N_7008,N_6742,N_6372);
nand U7009 (N_7009,N_6137,N_6173);
xor U7010 (N_7010,N_6246,N_6429);
and U7011 (N_7011,N_6289,N_6073);
nand U7012 (N_7012,N_6718,N_6013);
and U7013 (N_7013,N_6974,N_6739);
and U7014 (N_7014,N_6381,N_6818);
xnor U7015 (N_7015,N_6897,N_6445);
xnor U7016 (N_7016,N_6942,N_6510);
and U7017 (N_7017,N_6489,N_6768);
or U7018 (N_7018,N_6437,N_6382);
or U7019 (N_7019,N_6957,N_6409);
or U7020 (N_7020,N_6842,N_6744);
nand U7021 (N_7021,N_6392,N_6106);
and U7022 (N_7022,N_6320,N_6646);
nor U7023 (N_7023,N_6324,N_6019);
xnor U7024 (N_7024,N_6254,N_6297);
and U7025 (N_7025,N_6209,N_6822);
xnor U7026 (N_7026,N_6090,N_6084);
xnor U7027 (N_7027,N_6155,N_6203);
xor U7028 (N_7028,N_6430,N_6117);
nand U7029 (N_7029,N_6538,N_6002);
and U7030 (N_7030,N_6357,N_6304);
xnor U7031 (N_7031,N_6714,N_6308);
nand U7032 (N_7032,N_6347,N_6699);
nor U7033 (N_7033,N_6984,N_6892);
or U7034 (N_7034,N_6956,N_6580);
nand U7035 (N_7035,N_6355,N_6815);
and U7036 (N_7036,N_6573,N_6423);
or U7037 (N_7037,N_6743,N_6218);
and U7038 (N_7038,N_6288,N_6303);
nand U7039 (N_7039,N_6681,N_6929);
nor U7040 (N_7040,N_6986,N_6804);
nor U7041 (N_7041,N_6583,N_6894);
or U7042 (N_7042,N_6260,N_6466);
and U7043 (N_7043,N_6647,N_6431);
nor U7044 (N_7044,N_6447,N_6458);
nor U7045 (N_7045,N_6734,N_6766);
or U7046 (N_7046,N_6459,N_6539);
and U7047 (N_7047,N_6018,N_6582);
or U7048 (N_7048,N_6505,N_6994);
or U7049 (N_7049,N_6448,N_6593);
nor U7050 (N_7050,N_6868,N_6726);
xnor U7051 (N_7051,N_6387,N_6206);
or U7052 (N_7052,N_6312,N_6270);
nand U7053 (N_7053,N_6835,N_6759);
xnor U7054 (N_7054,N_6735,N_6716);
nor U7055 (N_7055,N_6990,N_6074);
xor U7056 (N_7056,N_6152,N_6241);
and U7057 (N_7057,N_6700,N_6157);
and U7058 (N_7058,N_6677,N_6484);
xor U7059 (N_7059,N_6870,N_6008);
and U7060 (N_7060,N_6451,N_6778);
or U7061 (N_7061,N_6273,N_6220);
xnor U7062 (N_7062,N_6895,N_6888);
xor U7063 (N_7063,N_6454,N_6969);
or U7064 (N_7064,N_6980,N_6965);
nor U7065 (N_7065,N_6732,N_6258);
and U7066 (N_7066,N_6144,N_6380);
or U7067 (N_7067,N_6026,N_6032);
nor U7068 (N_7068,N_6029,N_6920);
and U7069 (N_7069,N_6690,N_6680);
nand U7070 (N_7070,N_6536,N_6577);
nand U7071 (N_7071,N_6648,N_6875);
and U7072 (N_7072,N_6444,N_6480);
nand U7073 (N_7073,N_6240,N_6396);
and U7074 (N_7074,N_6672,N_6323);
or U7075 (N_7075,N_6860,N_6419);
or U7076 (N_7076,N_6773,N_6050);
and U7077 (N_7077,N_6925,N_6350);
and U7078 (N_7078,N_6384,N_6615);
or U7079 (N_7079,N_6938,N_6821);
or U7080 (N_7080,N_6042,N_6841);
xnor U7081 (N_7081,N_6207,N_6356);
xor U7082 (N_7082,N_6330,N_6222);
nor U7083 (N_7083,N_6108,N_6611);
nand U7084 (N_7084,N_6671,N_6752);
xor U7085 (N_7085,N_6852,N_6488);
and U7086 (N_7086,N_6584,N_6004);
nand U7087 (N_7087,N_6941,N_6943);
nand U7088 (N_7088,N_6080,N_6478);
xnor U7089 (N_7089,N_6481,N_6632);
xor U7090 (N_7090,N_6238,N_6215);
nand U7091 (N_7091,N_6928,N_6418);
nand U7092 (N_7092,N_6039,N_6197);
nand U7093 (N_7093,N_6475,N_6493);
xor U7094 (N_7094,N_6406,N_6824);
and U7095 (N_7095,N_6118,N_6168);
nand U7096 (N_7096,N_6214,N_6398);
xnor U7097 (N_7097,N_6085,N_6282);
nor U7098 (N_7098,N_6736,N_6154);
nor U7099 (N_7099,N_6999,N_6464);
or U7100 (N_7100,N_6887,N_6721);
and U7101 (N_7101,N_6024,N_6201);
and U7102 (N_7102,N_6587,N_6031);
nor U7103 (N_7103,N_6693,N_6912);
nand U7104 (N_7104,N_6972,N_6257);
and U7105 (N_7105,N_6198,N_6194);
nor U7106 (N_7106,N_6377,N_6973);
or U7107 (N_7107,N_6015,N_6523);
xor U7108 (N_7108,N_6500,N_6914);
nand U7109 (N_7109,N_6666,N_6124);
nor U7110 (N_7110,N_6149,N_6182);
xnor U7111 (N_7111,N_6638,N_6623);
and U7112 (N_7112,N_6075,N_6760);
and U7113 (N_7113,N_6656,N_6286);
or U7114 (N_7114,N_6283,N_6809);
nor U7115 (N_7115,N_6176,N_6100);
nand U7116 (N_7116,N_6446,N_6335);
and U7117 (N_7117,N_6777,N_6053);
xor U7118 (N_7118,N_6056,N_6457);
and U7119 (N_7119,N_6810,N_6256);
and U7120 (N_7120,N_6813,N_6247);
nor U7121 (N_7121,N_6911,N_6263);
and U7122 (N_7122,N_6313,N_6307);
nor U7123 (N_7123,N_6939,N_6219);
xor U7124 (N_7124,N_6397,N_6132);
nor U7125 (N_7125,N_6959,N_6571);
xnor U7126 (N_7126,N_6055,N_6848);
nand U7127 (N_7127,N_6242,N_6131);
nand U7128 (N_7128,N_6153,N_6927);
nor U7129 (N_7129,N_6417,N_6688);
or U7130 (N_7130,N_6800,N_6715);
nor U7131 (N_7131,N_6618,N_6439);
and U7132 (N_7132,N_6295,N_6122);
and U7133 (N_7133,N_6245,N_6910);
or U7134 (N_7134,N_6280,N_6292);
nand U7135 (N_7135,N_6874,N_6299);
xor U7136 (N_7136,N_6436,N_6851);
or U7137 (N_7137,N_6798,N_6094);
nor U7138 (N_7138,N_6151,N_6613);
or U7139 (N_7139,N_6544,N_6180);
and U7140 (N_7140,N_6184,N_6087);
xor U7141 (N_7141,N_6937,N_6591);
xor U7142 (N_7142,N_6048,N_6903);
xnor U7143 (N_7143,N_6104,N_6059);
nor U7144 (N_7144,N_6170,N_6129);
or U7145 (N_7145,N_6685,N_6163);
and U7146 (N_7146,N_6027,N_6239);
or U7147 (N_7147,N_6373,N_6531);
and U7148 (N_7148,N_6595,N_6267);
and U7149 (N_7149,N_6713,N_6639);
nand U7150 (N_7150,N_6915,N_6044);
and U7151 (N_7151,N_6005,N_6158);
nand U7152 (N_7152,N_6322,N_6832);
or U7153 (N_7153,N_6694,N_6196);
and U7154 (N_7154,N_6820,N_6594);
xor U7155 (N_7155,N_6125,N_6511);
xnor U7156 (N_7156,N_6881,N_6088);
nand U7157 (N_7157,N_6856,N_6022);
xnor U7158 (N_7158,N_6390,N_6837);
and U7159 (N_7159,N_6195,N_6020);
xnor U7160 (N_7160,N_6248,N_6907);
or U7161 (N_7161,N_6827,N_6253);
or U7162 (N_7162,N_6609,N_6754);
xnor U7163 (N_7163,N_6068,N_6534);
and U7164 (N_7164,N_6425,N_6668);
and U7165 (N_7165,N_6797,N_6963);
nand U7166 (N_7166,N_6787,N_6831);
and U7167 (N_7167,N_6626,N_6641);
xnor U7168 (N_7168,N_6477,N_6733);
nand U7169 (N_7169,N_6816,N_6231);
xor U7170 (N_7170,N_6096,N_6495);
xnor U7171 (N_7171,N_6847,N_6169);
nand U7172 (N_7172,N_6949,N_6934);
nand U7173 (N_7173,N_6041,N_6670);
or U7174 (N_7174,N_6072,N_6551);
or U7175 (N_7175,N_6922,N_6443);
and U7176 (N_7176,N_6605,N_6424);
nand U7177 (N_7177,N_6530,N_6228);
and U7178 (N_7178,N_6097,N_6871);
nor U7179 (N_7179,N_6473,N_6730);
or U7180 (N_7180,N_6741,N_6617);
nand U7181 (N_7181,N_6187,N_6954);
and U7182 (N_7182,N_6364,N_6342);
nand U7183 (N_7183,N_6720,N_6634);
xnor U7184 (N_7184,N_6452,N_6692);
nor U7185 (N_7185,N_6208,N_6416);
or U7186 (N_7186,N_6405,N_6790);
nand U7187 (N_7187,N_6675,N_6853);
and U7188 (N_7188,N_6558,N_6255);
xor U7189 (N_7189,N_6555,N_6327);
or U7190 (N_7190,N_6134,N_6037);
xnor U7191 (N_7191,N_6082,N_6628);
nand U7192 (N_7192,N_6300,N_6596);
nand U7193 (N_7193,N_6866,N_6612);
xnor U7194 (N_7194,N_6470,N_6191);
and U7195 (N_7195,N_6917,N_6123);
and U7196 (N_7196,N_6794,N_6126);
and U7197 (N_7197,N_6805,N_6183);
or U7198 (N_7198,N_6045,N_6225);
nor U7199 (N_7199,N_6686,N_6078);
xor U7200 (N_7200,N_6230,N_6321);
and U7201 (N_7201,N_6047,N_6479);
nand U7202 (N_7202,N_6515,N_6368);
nand U7203 (N_7203,N_6723,N_6896);
nand U7204 (N_7204,N_6753,N_6375);
and U7205 (N_7205,N_6614,N_6119);
or U7206 (N_7206,N_6394,N_6636);
xnor U7207 (N_7207,N_6232,N_6876);
nand U7208 (N_7208,N_6621,N_6823);
nand U7209 (N_7209,N_6345,N_6360);
or U7210 (N_7210,N_6758,N_6052);
or U7211 (N_7211,N_6449,N_6236);
or U7212 (N_7212,N_6293,N_6003);
or U7213 (N_7213,N_6962,N_6838);
nor U7214 (N_7214,N_6947,N_6465);
nand U7215 (N_7215,N_6644,N_6058);
nand U7216 (N_7216,N_6784,N_6977);
and U7217 (N_7217,N_6834,N_6843);
or U7218 (N_7218,N_6991,N_6606);
nor U7219 (N_7219,N_6287,N_6918);
nand U7220 (N_7220,N_6262,N_6840);
and U7221 (N_7221,N_6395,N_6789);
xor U7222 (N_7222,N_6252,N_6844);
and U7223 (N_7223,N_6140,N_6537);
and U7224 (N_7224,N_6542,N_6676);
nor U7225 (N_7225,N_6998,N_6791);
or U7226 (N_7226,N_6305,N_6442);
xnor U7227 (N_7227,N_6358,N_6079);
xnor U7228 (N_7228,N_6565,N_6830);
nand U7229 (N_7229,N_6175,N_6376);
nand U7230 (N_7230,N_6642,N_6845);
xnor U7231 (N_7231,N_6143,N_6349);
and U7232 (N_7232,N_6036,N_6955);
nor U7233 (N_7233,N_6427,N_6795);
and U7234 (N_7234,N_6202,N_6547);
nand U7235 (N_7235,N_6878,N_6359);
and U7236 (N_7236,N_6598,N_6948);
xnor U7237 (N_7237,N_6265,N_6521);
nor U7238 (N_7238,N_6657,N_6487);
nor U7239 (N_7239,N_6924,N_6344);
nand U7240 (N_7240,N_6669,N_6340);
nor U7241 (N_7241,N_6828,N_6091);
nand U7242 (N_7242,N_6512,N_6251);
nand U7243 (N_7243,N_6640,N_6069);
nor U7244 (N_7244,N_6399,N_6826);
xnor U7245 (N_7245,N_6599,N_6568);
and U7246 (N_7246,N_6112,N_6127);
nand U7247 (N_7247,N_6908,N_6562);
nor U7248 (N_7248,N_6764,N_6334);
nor U7249 (N_7249,N_6105,N_6825);
and U7250 (N_7250,N_6362,N_6433);
and U7251 (N_7251,N_6520,N_6517);
nor U7252 (N_7252,N_6114,N_6796);
nor U7253 (N_7253,N_6077,N_6543);
or U7254 (N_7254,N_6979,N_6566);
nand U7255 (N_7255,N_6936,N_6412);
xor U7256 (N_7256,N_6585,N_6552);
and U7257 (N_7257,N_6627,N_6064);
nand U7258 (N_7258,N_6467,N_6331);
nor U7259 (N_7259,N_6574,N_6393);
xnor U7260 (N_7260,N_6710,N_6630);
and U7261 (N_7261,N_6223,N_6361);
nor U7262 (N_7262,N_6863,N_6066);
or U7263 (N_7263,N_6259,N_6785);
nand U7264 (N_7264,N_6498,N_6689);
nor U7265 (N_7265,N_6235,N_6607);
nor U7266 (N_7266,N_6659,N_6391);
nand U7267 (N_7267,N_6839,N_6325);
nor U7268 (N_7268,N_6033,N_6635);
and U7269 (N_7269,N_6142,N_6034);
nand U7270 (N_7270,N_6503,N_6775);
nor U7271 (N_7271,N_6643,N_6575);
nor U7272 (N_7272,N_6369,N_6040);
and U7273 (N_7273,N_6421,N_6237);
and U7274 (N_7274,N_6535,N_6211);
nand U7275 (N_7275,N_6490,N_6833);
nor U7276 (N_7276,N_6367,N_6148);
nand U7277 (N_7277,N_6755,N_6919);
or U7278 (N_7278,N_6001,N_6160);
or U7279 (N_7279,N_6712,N_6468);
or U7280 (N_7280,N_6946,N_6590);
nor U7281 (N_7281,N_6803,N_6179);
and U7282 (N_7282,N_6882,N_6704);
or U7283 (N_7283,N_6904,N_6886);
nor U7284 (N_7284,N_6185,N_6441);
nand U7285 (N_7285,N_6724,N_6210);
and U7286 (N_7286,N_6683,N_6109);
nor U7287 (N_7287,N_6276,N_6660);
and U7288 (N_7288,N_6654,N_6757);
nor U7289 (N_7289,N_6306,N_6243);
or U7290 (N_7290,N_6836,N_6093);
nand U7291 (N_7291,N_6099,N_6862);
and U7292 (N_7292,N_6563,N_6224);
and U7293 (N_7293,N_6859,N_6217);
or U7294 (N_7294,N_6318,N_6136);
or U7295 (N_7295,N_6885,N_6861);
nand U7296 (N_7296,N_6051,N_6291);
nand U7297 (N_7297,N_6389,N_6776);
and U7298 (N_7298,N_6961,N_6631);
or U7299 (N_7299,N_6597,N_6341);
nand U7300 (N_7300,N_6524,N_6738);
nor U7301 (N_7301,N_6450,N_6719);
nand U7302 (N_7302,N_6814,N_6199);
and U7303 (N_7303,N_6731,N_6701);
nor U7304 (N_7304,N_6592,N_6352);
xor U7305 (N_7305,N_6687,N_6801);
and U7306 (N_7306,N_6854,N_6649);
nor U7307 (N_7307,N_6435,N_6301);
nand U7308 (N_7308,N_6916,N_6604);
nor U7309 (N_7309,N_6684,N_6296);
and U7310 (N_7310,N_6411,N_6401);
xnor U7311 (N_7311,N_6788,N_6455);
and U7312 (N_7312,N_6576,N_6010);
and U7313 (N_7313,N_6983,N_6319);
and U7314 (N_7314,N_6966,N_6767);
xor U7315 (N_7315,N_6637,N_6165);
and U7316 (N_7316,N_6407,N_6346);
xor U7317 (N_7317,N_6930,N_6229);
nand U7318 (N_7318,N_6779,N_6111);
or U7319 (N_7319,N_6374,N_6332);
nor U7320 (N_7320,N_6200,N_6561);
and U7321 (N_7321,N_6933,N_6829);
nor U7322 (N_7322,N_6471,N_6279);
or U7323 (N_7323,N_6740,N_6522);
and U7324 (N_7324,N_6062,N_6549);
and U7325 (N_7325,N_6653,N_6438);
nand U7326 (N_7326,N_6532,N_6463);
and U7327 (N_7327,N_6817,N_6808);
or U7328 (N_7328,N_6309,N_6290);
and U7329 (N_7329,N_6261,N_6769);
and U7330 (N_7330,N_6770,N_6560);
nor U7331 (N_7331,N_6661,N_6378);
nand U7332 (N_7332,N_6996,N_6171);
or U7333 (N_7333,N_6932,N_6923);
and U7334 (N_7334,N_6899,N_6453);
nor U7335 (N_7335,N_6083,N_6501);
nand U7336 (N_7336,N_6216,N_6343);
or U7337 (N_7337,N_6130,N_6415);
and U7338 (N_7338,N_6940,N_6329);
and U7339 (N_7339,N_6095,N_6975);
and U7340 (N_7340,N_6909,N_6061);
or U7341 (N_7341,N_6128,N_6071);
xor U7342 (N_7342,N_6662,N_6205);
and U7343 (N_7343,N_6012,N_6545);
or U7344 (N_7344,N_6746,N_6750);
nor U7345 (N_7345,N_6705,N_6548);
or U7346 (N_7346,N_6120,N_6749);
nor U7347 (N_7347,N_6164,N_6278);
or U7348 (N_7348,N_6655,N_6610);
xnor U7349 (N_7349,N_6469,N_6586);
nand U7350 (N_7350,N_6772,N_6107);
nor U7351 (N_7351,N_6336,N_6021);
nor U7352 (N_7352,N_6101,N_6284);
nand U7353 (N_7353,N_6997,N_6978);
and U7354 (N_7354,N_6703,N_6460);
or U7355 (N_7355,N_6065,N_6951);
xor U7356 (N_7356,N_6000,N_6567);
nor U7357 (N_7357,N_6893,N_6366);
or U7358 (N_7358,N_6958,N_6529);
xnor U7359 (N_7359,N_6811,N_6492);
xnor U7360 (N_7360,N_6181,N_6633);
nor U7361 (N_7361,N_6275,N_6508);
or U7362 (N_7362,N_6855,N_6518);
or U7363 (N_7363,N_6900,N_6141);
nor U7364 (N_7364,N_6432,N_6076);
nand U7365 (N_7365,N_6509,N_6652);
nor U7366 (N_7366,N_6474,N_6428);
nor U7367 (N_7367,N_6608,N_6514);
xnor U7368 (N_7368,N_6926,N_6988);
and U7369 (N_7369,N_6227,N_6748);
and U7370 (N_7370,N_6858,N_6519);
xor U7371 (N_7371,N_6115,N_6277);
nor U7372 (N_7372,N_6968,N_6651);
or U7373 (N_7373,N_6023,N_6717);
xor U7374 (N_7374,N_6025,N_6440);
or U7375 (N_7375,N_6890,N_6186);
xor U7376 (N_7376,N_6167,N_6014);
and U7377 (N_7377,N_6673,N_6849);
and U7378 (N_7378,N_6883,N_6485);
xnor U7379 (N_7379,N_6906,N_6526);
or U7380 (N_7380,N_6317,N_6150);
and U7381 (N_7381,N_6133,N_6867);
and U7382 (N_7382,N_6159,N_6970);
nor U7383 (N_7383,N_6745,N_6365);
nand U7384 (N_7384,N_6113,N_6622);
and U7385 (N_7385,N_6650,N_6725);
or U7386 (N_7386,N_6880,N_6695);
and U7387 (N_7387,N_6889,N_6879);
nor U7388 (N_7388,N_6316,N_6891);
or U7389 (N_7389,N_6782,N_6281);
nor U7390 (N_7390,N_6935,N_6383);
and U7391 (N_7391,N_6172,N_6121);
nor U7392 (N_7392,N_6110,N_6326);
nand U7393 (N_7393,N_6188,N_6901);
nand U7394 (N_7394,N_6658,N_6645);
nor U7395 (N_7395,N_6337,N_6410);
or U7396 (N_7396,N_6995,N_6092);
nand U7397 (N_7397,N_6271,N_6952);
or U7398 (N_7398,N_6353,N_6884);
or U7399 (N_7399,N_6011,N_6385);
and U7400 (N_7400,N_6351,N_6212);
xnor U7401 (N_7401,N_6625,N_6553);
and U7402 (N_7402,N_6146,N_6402);
or U7403 (N_7403,N_6145,N_6070);
nor U7404 (N_7404,N_6913,N_6985);
xnor U7405 (N_7405,N_6310,N_6722);
nor U7406 (N_7406,N_6116,N_6992);
xor U7407 (N_7407,N_6006,N_6166);
nand U7408 (N_7408,N_6264,N_6572);
nor U7409 (N_7409,N_6422,N_6865);
nor U7410 (N_7410,N_6976,N_6945);
or U7411 (N_7411,N_6494,N_6426);
xor U7412 (N_7412,N_6872,N_6348);
or U7413 (N_7413,N_6063,N_6799);
nor U7414 (N_7414,N_6667,N_6981);
xnor U7415 (N_7415,N_6679,N_6763);
xor U7416 (N_7416,N_6098,N_6192);
nor U7417 (N_7417,N_6204,N_6496);
and U7418 (N_7418,N_6971,N_6602);
or U7419 (N_7419,N_6781,N_6476);
xor U7420 (N_7420,N_6363,N_6371);
and U7421 (N_7421,N_6483,N_6864);
or U7422 (N_7422,N_6629,N_6302);
nand U7423 (N_7423,N_6274,N_6761);
nand U7424 (N_7424,N_6328,N_6806);
nand U7425 (N_7425,N_6786,N_6589);
and U7426 (N_7426,N_6054,N_6103);
nand U7427 (N_7427,N_6780,N_6221);
nor U7428 (N_7428,N_6162,N_6850);
nand U7429 (N_7429,N_6456,N_6921);
nand U7430 (N_7430,N_6771,N_6017);
or U7431 (N_7431,N_6482,N_6727);
nand U7432 (N_7432,N_6190,N_6783);
or U7433 (N_7433,N_6461,N_6525);
nand U7434 (N_7434,N_6472,N_6386);
nor U7435 (N_7435,N_6035,N_6857);
nand U7436 (N_7436,N_6601,N_6314);
xor U7437 (N_7437,N_6707,N_6507);
nor U7438 (N_7438,N_6665,N_6413);
or U7439 (N_7439,N_6603,N_6388);
and U7440 (N_7440,N_6819,N_6138);
nand U7441 (N_7441,N_6737,N_6765);
and U7442 (N_7442,N_6953,N_6135);
nor U7443 (N_7443,N_6504,N_6339);
nor U7444 (N_7444,N_6311,N_6564);
nand U7445 (N_7445,N_6728,N_6193);
and U7446 (N_7446,N_6931,N_6226);
and U7447 (N_7447,N_6902,N_6379);
nor U7448 (N_7448,N_6729,N_6964);
xor U7449 (N_7449,N_6081,N_6400);
nand U7450 (N_7450,N_6016,N_6403);
nor U7451 (N_7451,N_6569,N_6007);
nand U7452 (N_7452,N_6462,N_6967);
xor U7453 (N_7453,N_6499,N_6028);
xnor U7454 (N_7454,N_6404,N_6497);
nand U7455 (N_7455,N_6950,N_6960);
or U7456 (N_7456,N_6709,N_6579);
nor U7457 (N_7457,N_6556,N_6756);
xor U7458 (N_7458,N_6294,N_6674);
nand U7459 (N_7459,N_6269,N_6702);
xnor U7460 (N_7460,N_6414,N_6102);
nor U7461 (N_7461,N_6774,N_6812);
and U7462 (N_7462,N_6009,N_6533);
xnor U7463 (N_7463,N_6711,N_6559);
or U7464 (N_7464,N_6898,N_6057);
nor U7465 (N_7465,N_6354,N_6541);
nand U7466 (N_7466,N_6491,N_6333);
xor U7467 (N_7467,N_6156,N_6616);
nor U7468 (N_7468,N_6664,N_6060);
nor U7469 (N_7469,N_6506,N_6298);
nand U7470 (N_7470,N_6043,N_6502);
nor U7471 (N_7471,N_6408,N_6989);
or U7472 (N_7472,N_6869,N_6486);
xor U7473 (N_7473,N_6516,N_6268);
xnor U7474 (N_7474,N_6234,N_6513);
or U7475 (N_7475,N_6581,N_6067);
or U7476 (N_7476,N_6046,N_6189);
xor U7477 (N_7477,N_6233,N_6554);
nor U7478 (N_7478,N_6338,N_6161);
xor U7479 (N_7479,N_6249,N_6086);
xnor U7480 (N_7480,N_6272,N_6807);
and U7481 (N_7481,N_6624,N_6682);
nand U7482 (N_7482,N_6546,N_6178);
and U7483 (N_7483,N_6540,N_6846);
or U7484 (N_7484,N_6213,N_6588);
nand U7485 (N_7485,N_6993,N_6944);
xnor U7486 (N_7486,N_6177,N_6420);
nor U7487 (N_7487,N_6678,N_6285);
xnor U7488 (N_7488,N_6600,N_6697);
xor U7489 (N_7489,N_6663,N_6434);
nand U7490 (N_7490,N_6873,N_6528);
and U7491 (N_7491,N_6905,N_6527);
nand U7492 (N_7492,N_6877,N_6706);
and U7493 (N_7493,N_6049,N_6708);
or U7494 (N_7494,N_6174,N_6244);
or U7495 (N_7495,N_6266,N_6987);
nor U7496 (N_7496,N_6620,N_6370);
nand U7497 (N_7497,N_6030,N_6250);
nand U7498 (N_7498,N_6557,N_6762);
or U7499 (N_7499,N_6698,N_6089);
nand U7500 (N_7500,N_6470,N_6118);
and U7501 (N_7501,N_6025,N_6680);
or U7502 (N_7502,N_6430,N_6001);
nand U7503 (N_7503,N_6058,N_6116);
and U7504 (N_7504,N_6460,N_6640);
and U7505 (N_7505,N_6406,N_6970);
or U7506 (N_7506,N_6321,N_6902);
nor U7507 (N_7507,N_6643,N_6274);
xnor U7508 (N_7508,N_6397,N_6043);
and U7509 (N_7509,N_6179,N_6205);
nand U7510 (N_7510,N_6878,N_6118);
or U7511 (N_7511,N_6427,N_6028);
and U7512 (N_7512,N_6414,N_6479);
nand U7513 (N_7513,N_6817,N_6356);
nand U7514 (N_7514,N_6715,N_6416);
xnor U7515 (N_7515,N_6273,N_6430);
and U7516 (N_7516,N_6037,N_6570);
nand U7517 (N_7517,N_6956,N_6842);
xor U7518 (N_7518,N_6421,N_6051);
nand U7519 (N_7519,N_6332,N_6413);
or U7520 (N_7520,N_6307,N_6795);
and U7521 (N_7521,N_6561,N_6986);
nand U7522 (N_7522,N_6653,N_6446);
or U7523 (N_7523,N_6877,N_6350);
or U7524 (N_7524,N_6549,N_6179);
xor U7525 (N_7525,N_6303,N_6089);
nor U7526 (N_7526,N_6641,N_6274);
nand U7527 (N_7527,N_6206,N_6094);
and U7528 (N_7528,N_6127,N_6011);
or U7529 (N_7529,N_6485,N_6038);
or U7530 (N_7530,N_6574,N_6694);
xnor U7531 (N_7531,N_6507,N_6120);
and U7532 (N_7532,N_6014,N_6940);
xor U7533 (N_7533,N_6666,N_6956);
xnor U7534 (N_7534,N_6586,N_6991);
nand U7535 (N_7535,N_6764,N_6217);
and U7536 (N_7536,N_6716,N_6857);
and U7537 (N_7537,N_6466,N_6634);
nor U7538 (N_7538,N_6066,N_6810);
nor U7539 (N_7539,N_6595,N_6970);
xor U7540 (N_7540,N_6721,N_6762);
xnor U7541 (N_7541,N_6453,N_6457);
or U7542 (N_7542,N_6575,N_6196);
xnor U7543 (N_7543,N_6275,N_6873);
nor U7544 (N_7544,N_6041,N_6089);
xor U7545 (N_7545,N_6346,N_6223);
and U7546 (N_7546,N_6479,N_6031);
nand U7547 (N_7547,N_6161,N_6125);
nor U7548 (N_7548,N_6027,N_6580);
nand U7549 (N_7549,N_6045,N_6250);
nor U7550 (N_7550,N_6769,N_6428);
and U7551 (N_7551,N_6899,N_6637);
and U7552 (N_7552,N_6529,N_6880);
and U7553 (N_7553,N_6959,N_6910);
or U7554 (N_7554,N_6746,N_6801);
and U7555 (N_7555,N_6961,N_6534);
or U7556 (N_7556,N_6620,N_6802);
xor U7557 (N_7557,N_6766,N_6454);
nand U7558 (N_7558,N_6194,N_6195);
nand U7559 (N_7559,N_6267,N_6789);
xnor U7560 (N_7560,N_6954,N_6487);
nand U7561 (N_7561,N_6323,N_6304);
nor U7562 (N_7562,N_6144,N_6137);
nand U7563 (N_7563,N_6130,N_6153);
nor U7564 (N_7564,N_6053,N_6292);
nand U7565 (N_7565,N_6295,N_6010);
nand U7566 (N_7566,N_6289,N_6175);
nand U7567 (N_7567,N_6850,N_6403);
and U7568 (N_7568,N_6734,N_6786);
nand U7569 (N_7569,N_6823,N_6714);
nor U7570 (N_7570,N_6712,N_6412);
nor U7571 (N_7571,N_6848,N_6904);
xnor U7572 (N_7572,N_6826,N_6243);
xor U7573 (N_7573,N_6034,N_6160);
and U7574 (N_7574,N_6165,N_6285);
and U7575 (N_7575,N_6333,N_6279);
and U7576 (N_7576,N_6288,N_6172);
and U7577 (N_7577,N_6824,N_6982);
xor U7578 (N_7578,N_6045,N_6147);
and U7579 (N_7579,N_6366,N_6155);
nor U7580 (N_7580,N_6258,N_6612);
or U7581 (N_7581,N_6348,N_6336);
or U7582 (N_7582,N_6548,N_6896);
and U7583 (N_7583,N_6690,N_6169);
nor U7584 (N_7584,N_6116,N_6100);
and U7585 (N_7585,N_6514,N_6628);
or U7586 (N_7586,N_6168,N_6236);
nand U7587 (N_7587,N_6394,N_6497);
nand U7588 (N_7588,N_6782,N_6764);
or U7589 (N_7589,N_6788,N_6745);
nand U7590 (N_7590,N_6588,N_6492);
xor U7591 (N_7591,N_6534,N_6959);
xnor U7592 (N_7592,N_6919,N_6553);
or U7593 (N_7593,N_6673,N_6639);
or U7594 (N_7594,N_6048,N_6972);
nand U7595 (N_7595,N_6679,N_6376);
nand U7596 (N_7596,N_6027,N_6500);
or U7597 (N_7597,N_6543,N_6190);
xor U7598 (N_7598,N_6463,N_6152);
and U7599 (N_7599,N_6956,N_6374);
nor U7600 (N_7600,N_6306,N_6485);
nor U7601 (N_7601,N_6853,N_6417);
and U7602 (N_7602,N_6939,N_6299);
and U7603 (N_7603,N_6323,N_6174);
and U7604 (N_7604,N_6623,N_6495);
or U7605 (N_7605,N_6286,N_6327);
nor U7606 (N_7606,N_6600,N_6582);
or U7607 (N_7607,N_6033,N_6428);
or U7608 (N_7608,N_6878,N_6413);
and U7609 (N_7609,N_6921,N_6522);
xor U7610 (N_7610,N_6206,N_6534);
and U7611 (N_7611,N_6689,N_6758);
nor U7612 (N_7612,N_6359,N_6855);
nor U7613 (N_7613,N_6993,N_6560);
and U7614 (N_7614,N_6401,N_6757);
xnor U7615 (N_7615,N_6882,N_6981);
or U7616 (N_7616,N_6186,N_6893);
nor U7617 (N_7617,N_6326,N_6217);
or U7618 (N_7618,N_6933,N_6232);
nand U7619 (N_7619,N_6748,N_6172);
and U7620 (N_7620,N_6619,N_6484);
xor U7621 (N_7621,N_6310,N_6645);
or U7622 (N_7622,N_6820,N_6337);
or U7623 (N_7623,N_6180,N_6824);
nand U7624 (N_7624,N_6991,N_6651);
or U7625 (N_7625,N_6410,N_6027);
nand U7626 (N_7626,N_6302,N_6512);
xor U7627 (N_7627,N_6542,N_6104);
nand U7628 (N_7628,N_6453,N_6018);
xnor U7629 (N_7629,N_6319,N_6976);
xor U7630 (N_7630,N_6574,N_6276);
nand U7631 (N_7631,N_6204,N_6577);
nor U7632 (N_7632,N_6813,N_6135);
nor U7633 (N_7633,N_6656,N_6840);
or U7634 (N_7634,N_6972,N_6170);
and U7635 (N_7635,N_6996,N_6178);
xor U7636 (N_7636,N_6216,N_6147);
nor U7637 (N_7637,N_6424,N_6650);
xor U7638 (N_7638,N_6029,N_6527);
nand U7639 (N_7639,N_6015,N_6747);
nand U7640 (N_7640,N_6667,N_6640);
or U7641 (N_7641,N_6113,N_6851);
and U7642 (N_7642,N_6714,N_6734);
and U7643 (N_7643,N_6442,N_6883);
xor U7644 (N_7644,N_6699,N_6547);
xnor U7645 (N_7645,N_6635,N_6868);
nor U7646 (N_7646,N_6914,N_6343);
xnor U7647 (N_7647,N_6234,N_6236);
and U7648 (N_7648,N_6636,N_6488);
nor U7649 (N_7649,N_6203,N_6017);
or U7650 (N_7650,N_6418,N_6073);
nand U7651 (N_7651,N_6695,N_6408);
or U7652 (N_7652,N_6959,N_6965);
xor U7653 (N_7653,N_6015,N_6605);
nand U7654 (N_7654,N_6777,N_6837);
or U7655 (N_7655,N_6667,N_6704);
and U7656 (N_7656,N_6406,N_6275);
nor U7657 (N_7657,N_6622,N_6746);
nand U7658 (N_7658,N_6904,N_6983);
nand U7659 (N_7659,N_6299,N_6018);
nand U7660 (N_7660,N_6140,N_6653);
xor U7661 (N_7661,N_6620,N_6055);
nor U7662 (N_7662,N_6587,N_6033);
and U7663 (N_7663,N_6832,N_6790);
nor U7664 (N_7664,N_6009,N_6719);
xor U7665 (N_7665,N_6834,N_6112);
nor U7666 (N_7666,N_6808,N_6887);
and U7667 (N_7667,N_6398,N_6944);
nor U7668 (N_7668,N_6406,N_6522);
nor U7669 (N_7669,N_6593,N_6874);
or U7670 (N_7670,N_6263,N_6921);
or U7671 (N_7671,N_6661,N_6275);
or U7672 (N_7672,N_6336,N_6450);
nor U7673 (N_7673,N_6677,N_6435);
nand U7674 (N_7674,N_6094,N_6149);
nor U7675 (N_7675,N_6844,N_6042);
and U7676 (N_7676,N_6869,N_6907);
nand U7677 (N_7677,N_6706,N_6800);
nor U7678 (N_7678,N_6721,N_6980);
nor U7679 (N_7679,N_6341,N_6668);
nor U7680 (N_7680,N_6642,N_6432);
nor U7681 (N_7681,N_6405,N_6566);
nand U7682 (N_7682,N_6719,N_6299);
nand U7683 (N_7683,N_6315,N_6782);
nand U7684 (N_7684,N_6748,N_6173);
or U7685 (N_7685,N_6167,N_6246);
nand U7686 (N_7686,N_6798,N_6613);
nor U7687 (N_7687,N_6016,N_6578);
or U7688 (N_7688,N_6446,N_6398);
and U7689 (N_7689,N_6970,N_6507);
xnor U7690 (N_7690,N_6099,N_6298);
nand U7691 (N_7691,N_6831,N_6911);
and U7692 (N_7692,N_6240,N_6715);
nand U7693 (N_7693,N_6992,N_6137);
xor U7694 (N_7694,N_6839,N_6866);
and U7695 (N_7695,N_6220,N_6861);
nor U7696 (N_7696,N_6630,N_6928);
or U7697 (N_7697,N_6010,N_6899);
and U7698 (N_7698,N_6978,N_6811);
nand U7699 (N_7699,N_6613,N_6394);
nor U7700 (N_7700,N_6768,N_6219);
nor U7701 (N_7701,N_6737,N_6194);
nand U7702 (N_7702,N_6777,N_6407);
nor U7703 (N_7703,N_6373,N_6505);
xor U7704 (N_7704,N_6887,N_6323);
nand U7705 (N_7705,N_6934,N_6289);
and U7706 (N_7706,N_6289,N_6112);
nor U7707 (N_7707,N_6842,N_6301);
xnor U7708 (N_7708,N_6009,N_6649);
nor U7709 (N_7709,N_6740,N_6084);
xor U7710 (N_7710,N_6486,N_6176);
nor U7711 (N_7711,N_6264,N_6196);
and U7712 (N_7712,N_6937,N_6941);
nand U7713 (N_7713,N_6161,N_6413);
nand U7714 (N_7714,N_6352,N_6781);
nand U7715 (N_7715,N_6875,N_6389);
xor U7716 (N_7716,N_6383,N_6393);
nor U7717 (N_7717,N_6319,N_6459);
xor U7718 (N_7718,N_6391,N_6322);
nand U7719 (N_7719,N_6903,N_6137);
xor U7720 (N_7720,N_6912,N_6169);
nor U7721 (N_7721,N_6132,N_6970);
nor U7722 (N_7722,N_6155,N_6458);
or U7723 (N_7723,N_6645,N_6339);
and U7724 (N_7724,N_6445,N_6418);
or U7725 (N_7725,N_6763,N_6169);
nor U7726 (N_7726,N_6103,N_6882);
or U7727 (N_7727,N_6340,N_6759);
nor U7728 (N_7728,N_6002,N_6371);
xor U7729 (N_7729,N_6111,N_6303);
nor U7730 (N_7730,N_6686,N_6185);
and U7731 (N_7731,N_6709,N_6535);
or U7732 (N_7732,N_6282,N_6588);
nor U7733 (N_7733,N_6224,N_6050);
or U7734 (N_7734,N_6106,N_6926);
nor U7735 (N_7735,N_6420,N_6402);
or U7736 (N_7736,N_6132,N_6497);
or U7737 (N_7737,N_6200,N_6204);
or U7738 (N_7738,N_6392,N_6821);
or U7739 (N_7739,N_6769,N_6078);
and U7740 (N_7740,N_6999,N_6578);
nor U7741 (N_7741,N_6456,N_6557);
xor U7742 (N_7742,N_6722,N_6148);
or U7743 (N_7743,N_6132,N_6511);
xnor U7744 (N_7744,N_6266,N_6946);
or U7745 (N_7745,N_6617,N_6315);
nor U7746 (N_7746,N_6376,N_6362);
nor U7747 (N_7747,N_6302,N_6266);
and U7748 (N_7748,N_6163,N_6482);
xnor U7749 (N_7749,N_6873,N_6430);
nand U7750 (N_7750,N_6236,N_6056);
xor U7751 (N_7751,N_6171,N_6795);
nand U7752 (N_7752,N_6998,N_6990);
nand U7753 (N_7753,N_6420,N_6026);
nor U7754 (N_7754,N_6120,N_6034);
xor U7755 (N_7755,N_6557,N_6693);
or U7756 (N_7756,N_6985,N_6271);
nand U7757 (N_7757,N_6506,N_6131);
nor U7758 (N_7758,N_6128,N_6539);
nor U7759 (N_7759,N_6521,N_6671);
xnor U7760 (N_7760,N_6719,N_6287);
and U7761 (N_7761,N_6042,N_6767);
or U7762 (N_7762,N_6473,N_6882);
xor U7763 (N_7763,N_6089,N_6485);
and U7764 (N_7764,N_6338,N_6631);
nor U7765 (N_7765,N_6414,N_6715);
nor U7766 (N_7766,N_6462,N_6234);
xor U7767 (N_7767,N_6891,N_6837);
nor U7768 (N_7768,N_6755,N_6278);
xnor U7769 (N_7769,N_6421,N_6533);
and U7770 (N_7770,N_6457,N_6798);
nand U7771 (N_7771,N_6034,N_6266);
xor U7772 (N_7772,N_6771,N_6055);
xnor U7773 (N_7773,N_6120,N_6083);
nand U7774 (N_7774,N_6195,N_6508);
nor U7775 (N_7775,N_6466,N_6067);
xor U7776 (N_7776,N_6174,N_6170);
nand U7777 (N_7777,N_6140,N_6528);
nor U7778 (N_7778,N_6969,N_6028);
nand U7779 (N_7779,N_6896,N_6373);
nand U7780 (N_7780,N_6436,N_6218);
and U7781 (N_7781,N_6811,N_6729);
xor U7782 (N_7782,N_6693,N_6983);
and U7783 (N_7783,N_6842,N_6577);
and U7784 (N_7784,N_6718,N_6003);
xor U7785 (N_7785,N_6430,N_6002);
xnor U7786 (N_7786,N_6641,N_6414);
xor U7787 (N_7787,N_6021,N_6359);
xor U7788 (N_7788,N_6726,N_6373);
and U7789 (N_7789,N_6235,N_6028);
or U7790 (N_7790,N_6915,N_6971);
or U7791 (N_7791,N_6125,N_6638);
and U7792 (N_7792,N_6383,N_6514);
nor U7793 (N_7793,N_6531,N_6259);
or U7794 (N_7794,N_6654,N_6388);
nor U7795 (N_7795,N_6557,N_6628);
and U7796 (N_7796,N_6761,N_6276);
and U7797 (N_7797,N_6310,N_6026);
nand U7798 (N_7798,N_6170,N_6330);
nor U7799 (N_7799,N_6152,N_6600);
and U7800 (N_7800,N_6294,N_6090);
nand U7801 (N_7801,N_6381,N_6284);
or U7802 (N_7802,N_6469,N_6014);
nor U7803 (N_7803,N_6995,N_6583);
and U7804 (N_7804,N_6016,N_6502);
xor U7805 (N_7805,N_6075,N_6429);
or U7806 (N_7806,N_6012,N_6285);
and U7807 (N_7807,N_6942,N_6700);
xnor U7808 (N_7808,N_6978,N_6841);
and U7809 (N_7809,N_6809,N_6980);
nand U7810 (N_7810,N_6929,N_6696);
and U7811 (N_7811,N_6422,N_6594);
and U7812 (N_7812,N_6727,N_6535);
or U7813 (N_7813,N_6196,N_6240);
or U7814 (N_7814,N_6113,N_6085);
and U7815 (N_7815,N_6327,N_6613);
nor U7816 (N_7816,N_6383,N_6119);
and U7817 (N_7817,N_6609,N_6481);
xor U7818 (N_7818,N_6316,N_6253);
and U7819 (N_7819,N_6332,N_6158);
xor U7820 (N_7820,N_6915,N_6547);
nand U7821 (N_7821,N_6862,N_6646);
nor U7822 (N_7822,N_6900,N_6111);
and U7823 (N_7823,N_6168,N_6101);
nand U7824 (N_7824,N_6788,N_6466);
and U7825 (N_7825,N_6989,N_6873);
nand U7826 (N_7826,N_6880,N_6957);
or U7827 (N_7827,N_6058,N_6369);
and U7828 (N_7828,N_6706,N_6995);
or U7829 (N_7829,N_6104,N_6338);
xor U7830 (N_7830,N_6750,N_6086);
xor U7831 (N_7831,N_6282,N_6520);
or U7832 (N_7832,N_6858,N_6686);
or U7833 (N_7833,N_6995,N_6961);
nand U7834 (N_7834,N_6197,N_6334);
nand U7835 (N_7835,N_6871,N_6855);
nor U7836 (N_7836,N_6446,N_6342);
and U7837 (N_7837,N_6904,N_6175);
nor U7838 (N_7838,N_6132,N_6163);
xnor U7839 (N_7839,N_6446,N_6020);
nor U7840 (N_7840,N_6666,N_6078);
and U7841 (N_7841,N_6126,N_6637);
nor U7842 (N_7842,N_6775,N_6334);
xor U7843 (N_7843,N_6119,N_6041);
xor U7844 (N_7844,N_6530,N_6952);
and U7845 (N_7845,N_6223,N_6208);
or U7846 (N_7846,N_6824,N_6130);
xnor U7847 (N_7847,N_6524,N_6822);
nor U7848 (N_7848,N_6453,N_6382);
or U7849 (N_7849,N_6364,N_6489);
and U7850 (N_7850,N_6397,N_6219);
nor U7851 (N_7851,N_6817,N_6218);
and U7852 (N_7852,N_6977,N_6688);
or U7853 (N_7853,N_6024,N_6439);
nand U7854 (N_7854,N_6590,N_6535);
or U7855 (N_7855,N_6239,N_6381);
and U7856 (N_7856,N_6875,N_6169);
nand U7857 (N_7857,N_6414,N_6522);
or U7858 (N_7858,N_6813,N_6236);
and U7859 (N_7859,N_6430,N_6221);
or U7860 (N_7860,N_6901,N_6916);
and U7861 (N_7861,N_6703,N_6923);
nor U7862 (N_7862,N_6008,N_6342);
nor U7863 (N_7863,N_6840,N_6129);
nor U7864 (N_7864,N_6326,N_6983);
nor U7865 (N_7865,N_6981,N_6621);
nor U7866 (N_7866,N_6373,N_6751);
nor U7867 (N_7867,N_6624,N_6984);
or U7868 (N_7868,N_6339,N_6651);
or U7869 (N_7869,N_6331,N_6776);
nor U7870 (N_7870,N_6774,N_6230);
and U7871 (N_7871,N_6273,N_6246);
or U7872 (N_7872,N_6886,N_6462);
xnor U7873 (N_7873,N_6339,N_6890);
or U7874 (N_7874,N_6852,N_6228);
or U7875 (N_7875,N_6476,N_6761);
nor U7876 (N_7876,N_6578,N_6658);
and U7877 (N_7877,N_6349,N_6478);
and U7878 (N_7878,N_6730,N_6369);
nor U7879 (N_7879,N_6605,N_6197);
or U7880 (N_7880,N_6212,N_6489);
or U7881 (N_7881,N_6579,N_6855);
or U7882 (N_7882,N_6664,N_6993);
xor U7883 (N_7883,N_6398,N_6572);
and U7884 (N_7884,N_6032,N_6945);
xor U7885 (N_7885,N_6831,N_6929);
nand U7886 (N_7886,N_6265,N_6308);
nor U7887 (N_7887,N_6388,N_6464);
xor U7888 (N_7888,N_6391,N_6613);
and U7889 (N_7889,N_6290,N_6635);
nand U7890 (N_7890,N_6940,N_6969);
or U7891 (N_7891,N_6385,N_6616);
or U7892 (N_7892,N_6486,N_6078);
xnor U7893 (N_7893,N_6615,N_6113);
nand U7894 (N_7894,N_6391,N_6557);
nor U7895 (N_7895,N_6556,N_6212);
xor U7896 (N_7896,N_6987,N_6470);
nand U7897 (N_7897,N_6167,N_6033);
nor U7898 (N_7898,N_6250,N_6918);
nor U7899 (N_7899,N_6096,N_6415);
or U7900 (N_7900,N_6487,N_6998);
nand U7901 (N_7901,N_6487,N_6975);
or U7902 (N_7902,N_6088,N_6160);
nand U7903 (N_7903,N_6912,N_6332);
xnor U7904 (N_7904,N_6345,N_6525);
xor U7905 (N_7905,N_6939,N_6449);
xnor U7906 (N_7906,N_6527,N_6244);
and U7907 (N_7907,N_6346,N_6564);
nand U7908 (N_7908,N_6945,N_6841);
nand U7909 (N_7909,N_6310,N_6554);
or U7910 (N_7910,N_6643,N_6671);
xnor U7911 (N_7911,N_6148,N_6528);
nand U7912 (N_7912,N_6868,N_6454);
xnor U7913 (N_7913,N_6533,N_6300);
nor U7914 (N_7914,N_6931,N_6545);
xnor U7915 (N_7915,N_6053,N_6665);
nor U7916 (N_7916,N_6121,N_6222);
nor U7917 (N_7917,N_6105,N_6502);
xor U7918 (N_7918,N_6105,N_6328);
nand U7919 (N_7919,N_6945,N_6538);
nor U7920 (N_7920,N_6345,N_6542);
nor U7921 (N_7921,N_6469,N_6536);
or U7922 (N_7922,N_6205,N_6233);
and U7923 (N_7923,N_6773,N_6556);
and U7924 (N_7924,N_6677,N_6308);
nor U7925 (N_7925,N_6327,N_6855);
xor U7926 (N_7926,N_6662,N_6309);
and U7927 (N_7927,N_6287,N_6271);
and U7928 (N_7928,N_6895,N_6371);
and U7929 (N_7929,N_6003,N_6693);
xnor U7930 (N_7930,N_6641,N_6003);
or U7931 (N_7931,N_6006,N_6806);
xnor U7932 (N_7932,N_6258,N_6940);
or U7933 (N_7933,N_6711,N_6694);
nor U7934 (N_7934,N_6602,N_6734);
and U7935 (N_7935,N_6656,N_6452);
or U7936 (N_7936,N_6450,N_6435);
xor U7937 (N_7937,N_6591,N_6432);
and U7938 (N_7938,N_6010,N_6484);
xor U7939 (N_7939,N_6785,N_6408);
or U7940 (N_7940,N_6817,N_6664);
or U7941 (N_7941,N_6048,N_6700);
or U7942 (N_7942,N_6359,N_6890);
nor U7943 (N_7943,N_6995,N_6271);
nand U7944 (N_7944,N_6287,N_6470);
nand U7945 (N_7945,N_6856,N_6796);
and U7946 (N_7946,N_6214,N_6651);
or U7947 (N_7947,N_6879,N_6060);
nand U7948 (N_7948,N_6173,N_6309);
nor U7949 (N_7949,N_6790,N_6821);
and U7950 (N_7950,N_6141,N_6879);
xnor U7951 (N_7951,N_6625,N_6883);
or U7952 (N_7952,N_6220,N_6176);
and U7953 (N_7953,N_6715,N_6665);
nor U7954 (N_7954,N_6591,N_6255);
or U7955 (N_7955,N_6060,N_6745);
or U7956 (N_7956,N_6884,N_6253);
nand U7957 (N_7957,N_6943,N_6511);
and U7958 (N_7958,N_6195,N_6676);
xnor U7959 (N_7959,N_6550,N_6027);
nor U7960 (N_7960,N_6318,N_6694);
and U7961 (N_7961,N_6034,N_6576);
xnor U7962 (N_7962,N_6345,N_6903);
or U7963 (N_7963,N_6944,N_6629);
nor U7964 (N_7964,N_6775,N_6201);
xnor U7965 (N_7965,N_6306,N_6837);
and U7966 (N_7966,N_6438,N_6451);
nor U7967 (N_7967,N_6260,N_6892);
and U7968 (N_7968,N_6073,N_6541);
and U7969 (N_7969,N_6597,N_6025);
xor U7970 (N_7970,N_6370,N_6477);
or U7971 (N_7971,N_6517,N_6943);
and U7972 (N_7972,N_6883,N_6036);
nand U7973 (N_7973,N_6932,N_6987);
xnor U7974 (N_7974,N_6407,N_6434);
and U7975 (N_7975,N_6051,N_6122);
nand U7976 (N_7976,N_6606,N_6643);
or U7977 (N_7977,N_6871,N_6749);
nand U7978 (N_7978,N_6551,N_6348);
xnor U7979 (N_7979,N_6793,N_6073);
or U7980 (N_7980,N_6043,N_6532);
or U7981 (N_7981,N_6398,N_6598);
and U7982 (N_7982,N_6932,N_6913);
nor U7983 (N_7983,N_6947,N_6341);
xnor U7984 (N_7984,N_6673,N_6846);
nand U7985 (N_7985,N_6285,N_6284);
or U7986 (N_7986,N_6612,N_6213);
nand U7987 (N_7987,N_6176,N_6151);
nand U7988 (N_7988,N_6130,N_6639);
nand U7989 (N_7989,N_6342,N_6586);
nor U7990 (N_7990,N_6461,N_6650);
and U7991 (N_7991,N_6179,N_6605);
or U7992 (N_7992,N_6894,N_6747);
nor U7993 (N_7993,N_6911,N_6107);
nand U7994 (N_7994,N_6425,N_6151);
or U7995 (N_7995,N_6023,N_6437);
nor U7996 (N_7996,N_6467,N_6066);
xor U7997 (N_7997,N_6078,N_6286);
and U7998 (N_7998,N_6878,N_6781);
nor U7999 (N_7999,N_6606,N_6956);
nor U8000 (N_8000,N_7719,N_7335);
or U8001 (N_8001,N_7988,N_7153);
or U8002 (N_8002,N_7194,N_7385);
or U8003 (N_8003,N_7122,N_7108);
xor U8004 (N_8004,N_7818,N_7678);
nand U8005 (N_8005,N_7279,N_7535);
or U8006 (N_8006,N_7317,N_7869);
and U8007 (N_8007,N_7872,N_7050);
nand U8008 (N_8008,N_7713,N_7854);
xor U8009 (N_8009,N_7570,N_7145);
nand U8010 (N_8010,N_7039,N_7073);
nor U8011 (N_8011,N_7697,N_7051);
and U8012 (N_8012,N_7498,N_7646);
nand U8013 (N_8013,N_7307,N_7421);
xnor U8014 (N_8014,N_7972,N_7846);
nand U8015 (N_8015,N_7209,N_7827);
nor U8016 (N_8016,N_7769,N_7847);
xor U8017 (N_8017,N_7837,N_7605);
nand U8018 (N_8018,N_7264,N_7033);
xnor U8019 (N_8019,N_7926,N_7034);
nand U8020 (N_8020,N_7090,N_7329);
and U8021 (N_8021,N_7565,N_7306);
xnor U8022 (N_8022,N_7688,N_7579);
and U8023 (N_8023,N_7990,N_7223);
xnor U8024 (N_8024,N_7799,N_7763);
nand U8025 (N_8025,N_7971,N_7836);
nor U8026 (N_8026,N_7301,N_7013);
and U8027 (N_8027,N_7916,N_7734);
nor U8028 (N_8028,N_7158,N_7685);
xor U8029 (N_8029,N_7442,N_7466);
or U8030 (N_8030,N_7114,N_7155);
and U8031 (N_8031,N_7654,N_7290);
nand U8032 (N_8032,N_7035,N_7345);
xnor U8033 (N_8033,N_7377,N_7183);
xor U8034 (N_8034,N_7124,N_7800);
nor U8035 (N_8035,N_7206,N_7299);
xnor U8036 (N_8036,N_7427,N_7705);
and U8037 (N_8037,N_7957,N_7341);
xor U8038 (N_8038,N_7499,N_7454);
and U8039 (N_8039,N_7361,N_7426);
and U8040 (N_8040,N_7067,N_7208);
nor U8041 (N_8041,N_7105,N_7464);
nor U8042 (N_8042,N_7875,N_7046);
xor U8043 (N_8043,N_7251,N_7865);
or U8044 (N_8044,N_7729,N_7011);
nor U8045 (N_8045,N_7627,N_7227);
nor U8046 (N_8046,N_7031,N_7230);
nor U8047 (N_8047,N_7075,N_7337);
nand U8048 (N_8048,N_7170,N_7536);
or U8049 (N_8049,N_7977,N_7541);
or U8050 (N_8050,N_7524,N_7282);
or U8051 (N_8051,N_7140,N_7446);
or U8052 (N_8052,N_7045,N_7178);
and U8053 (N_8053,N_7042,N_7802);
xnor U8054 (N_8054,N_7908,N_7984);
or U8055 (N_8055,N_7581,N_7101);
nand U8056 (N_8056,N_7473,N_7297);
and U8057 (N_8057,N_7505,N_7249);
nand U8058 (N_8058,N_7512,N_7631);
and U8059 (N_8059,N_7597,N_7455);
xor U8060 (N_8060,N_7168,N_7439);
and U8061 (N_8061,N_7816,N_7423);
or U8062 (N_8062,N_7861,N_7344);
xor U8063 (N_8063,N_7923,N_7870);
or U8064 (N_8064,N_7970,N_7723);
or U8065 (N_8065,N_7893,N_7028);
and U8066 (N_8066,N_7214,N_7741);
nor U8067 (N_8067,N_7475,N_7416);
or U8068 (N_8068,N_7761,N_7089);
nor U8069 (N_8069,N_7559,N_7259);
and U8070 (N_8070,N_7691,N_7386);
nand U8071 (N_8071,N_7112,N_7213);
and U8072 (N_8072,N_7720,N_7815);
and U8073 (N_8073,N_7997,N_7954);
and U8074 (N_8074,N_7702,N_7975);
xnor U8075 (N_8075,N_7138,N_7623);
or U8076 (N_8076,N_7400,N_7233);
and U8077 (N_8077,N_7195,N_7468);
and U8078 (N_8078,N_7628,N_7561);
or U8079 (N_8079,N_7822,N_7521);
nor U8080 (N_8080,N_7405,N_7185);
xor U8081 (N_8081,N_7117,N_7128);
nand U8082 (N_8082,N_7991,N_7576);
or U8083 (N_8083,N_7292,N_7929);
or U8084 (N_8084,N_7146,N_7538);
nand U8085 (N_8085,N_7774,N_7196);
or U8086 (N_8086,N_7120,N_7712);
nand U8087 (N_8087,N_7103,N_7891);
and U8088 (N_8088,N_7071,N_7392);
and U8089 (N_8089,N_7900,N_7030);
xor U8090 (N_8090,N_7969,N_7298);
or U8091 (N_8091,N_7668,N_7266);
nor U8092 (N_8092,N_7490,N_7435);
and U8093 (N_8093,N_7281,N_7346);
and U8094 (N_8094,N_7932,N_7116);
nand U8095 (N_8095,N_7488,N_7353);
nor U8096 (N_8096,N_7171,N_7229);
xnor U8097 (N_8097,N_7210,N_7789);
and U8098 (N_8098,N_7440,N_7722);
nand U8099 (N_8099,N_7135,N_7636);
xnor U8100 (N_8100,N_7692,N_7895);
or U8101 (N_8101,N_7874,N_7262);
nor U8102 (N_8102,N_7326,N_7772);
nand U8103 (N_8103,N_7767,N_7620);
xor U8104 (N_8104,N_7617,N_7857);
or U8105 (N_8105,N_7265,N_7660);
nor U8106 (N_8106,N_7912,N_7083);
nor U8107 (N_8107,N_7193,N_7612);
and U8108 (N_8108,N_7023,N_7513);
and U8109 (N_8109,N_7411,N_7658);
or U8110 (N_8110,N_7580,N_7432);
nor U8111 (N_8111,N_7642,N_7111);
nor U8112 (N_8112,N_7684,N_7533);
and U8113 (N_8113,N_7902,N_7037);
or U8114 (N_8114,N_7302,N_7630);
or U8115 (N_8115,N_7064,N_7609);
or U8116 (N_8116,N_7093,N_7425);
and U8117 (N_8117,N_7755,N_7843);
and U8118 (N_8118,N_7157,N_7129);
and U8119 (N_8119,N_7441,N_7629);
and U8120 (N_8120,N_7644,N_7821);
or U8121 (N_8121,N_7563,N_7086);
nand U8122 (N_8122,N_7958,N_7504);
nor U8123 (N_8123,N_7389,N_7598);
or U8124 (N_8124,N_7635,N_7322);
nor U8125 (N_8125,N_7167,N_7974);
or U8126 (N_8126,N_7608,N_7358);
and U8127 (N_8127,N_7234,N_7641);
nand U8128 (N_8128,N_7921,N_7502);
or U8129 (N_8129,N_7099,N_7291);
and U8130 (N_8130,N_7825,N_7364);
and U8131 (N_8131,N_7731,N_7191);
and U8132 (N_8132,N_7324,N_7829);
and U8133 (N_8133,N_7169,N_7881);
xor U8134 (N_8134,N_7492,N_7496);
nand U8135 (N_8135,N_7607,N_7283);
xnor U8136 (N_8136,N_7651,N_7764);
nor U8137 (N_8137,N_7689,N_7486);
nor U8138 (N_8138,N_7239,N_7321);
xnor U8139 (N_8139,N_7733,N_7342);
xnor U8140 (N_8140,N_7257,N_7380);
nand U8141 (N_8141,N_7500,N_7632);
nand U8142 (N_8142,N_7901,N_7029);
nor U8143 (N_8143,N_7469,N_7069);
or U8144 (N_8144,N_7832,N_7671);
and U8145 (N_8145,N_7225,N_7550);
or U8146 (N_8146,N_7773,N_7918);
and U8147 (N_8147,N_7357,N_7296);
nor U8148 (N_8148,N_7395,N_7606);
and U8149 (N_8149,N_7087,N_7255);
or U8150 (N_8150,N_7394,N_7396);
nor U8151 (N_8151,N_7333,N_7066);
xor U8152 (N_8152,N_7373,N_7241);
and U8153 (N_8153,N_7273,N_7638);
xor U8154 (N_8154,N_7156,N_7352);
nand U8155 (N_8155,N_7928,N_7624);
nor U8156 (N_8156,N_7819,N_7205);
or U8157 (N_8157,N_7005,N_7882);
or U8158 (N_8158,N_7663,N_7586);
xnor U8159 (N_8159,N_7445,N_7978);
nor U8160 (N_8160,N_7422,N_7770);
xor U8161 (N_8161,N_7163,N_7634);
nand U8162 (N_8162,N_7061,N_7211);
and U8163 (N_8163,N_7759,N_7188);
and U8164 (N_8164,N_7845,N_7009);
nand U8165 (N_8165,N_7784,N_7104);
or U8166 (N_8166,N_7058,N_7224);
nand U8167 (N_8167,N_7313,N_7278);
or U8168 (N_8168,N_7704,N_7740);
nand U8169 (N_8169,N_7993,N_7760);
xor U8170 (N_8170,N_7899,N_7068);
or U8171 (N_8171,N_7700,N_7022);
nor U8172 (N_8172,N_7976,N_7369);
nand U8173 (N_8173,N_7952,N_7359);
xor U8174 (N_8174,N_7650,N_7356);
or U8175 (N_8175,N_7786,N_7657);
and U8176 (N_8176,N_7231,N_7556);
nor U8177 (N_8177,N_7433,N_7388);
xnor U8178 (N_8178,N_7826,N_7983);
xnor U8179 (N_8179,N_7938,N_7840);
nand U8180 (N_8180,N_7849,N_7949);
and U8181 (N_8181,N_7244,N_7094);
and U8182 (N_8182,N_7735,N_7300);
xnor U8183 (N_8183,N_7714,N_7944);
or U8184 (N_8184,N_7177,N_7510);
or U8185 (N_8185,N_7746,N_7235);
nor U8186 (N_8186,N_7184,N_7247);
xor U8187 (N_8187,N_7621,N_7343);
nor U8188 (N_8188,N_7830,N_7232);
or U8189 (N_8189,N_7002,N_7522);
nor U8190 (N_8190,N_7525,N_7543);
and U8191 (N_8191,N_7820,N_7771);
and U8192 (N_8192,N_7176,N_7238);
or U8193 (N_8193,N_7478,N_7204);
or U8194 (N_8194,N_7675,N_7626);
nand U8195 (N_8195,N_7043,N_7665);
and U8196 (N_8196,N_7413,N_7943);
nor U8197 (N_8197,N_7085,N_7012);
nor U8198 (N_8198,N_7980,N_7165);
nor U8199 (N_8199,N_7384,N_7387);
or U8200 (N_8200,N_7507,N_7765);
or U8201 (N_8201,N_7240,N_7611);
xor U8202 (N_8202,N_7141,N_7057);
xor U8203 (N_8203,N_7744,N_7585);
xor U8204 (N_8204,N_7986,N_7964);
and U8205 (N_8205,N_7564,N_7319);
nor U8206 (N_8206,N_7633,N_7372);
and U8207 (N_8207,N_7109,N_7877);
nor U8208 (N_8208,N_7001,N_7062);
nand U8209 (N_8209,N_7798,N_7474);
nand U8210 (N_8210,N_7973,N_7271);
nor U8211 (N_8211,N_7708,N_7399);
xnor U8212 (N_8212,N_7180,N_7070);
nand U8213 (N_8213,N_7796,N_7715);
and U8214 (N_8214,N_7376,N_7202);
xnor U8215 (N_8215,N_7219,N_7886);
nor U8216 (N_8216,N_7850,N_7197);
or U8217 (N_8217,N_7339,N_7573);
and U8218 (N_8218,N_7593,N_7560);
nor U8219 (N_8219,N_7936,N_7887);
or U8220 (N_8220,N_7098,N_7925);
xnor U8221 (N_8221,N_7753,N_7501);
nor U8222 (N_8222,N_7587,N_7792);
or U8223 (N_8223,N_7458,N_7709);
or U8224 (N_8224,N_7019,N_7443);
and U8225 (N_8225,N_7000,N_7123);
nand U8226 (N_8226,N_7788,N_7477);
and U8227 (N_8227,N_7495,N_7088);
nor U8228 (N_8228,N_7817,N_7481);
nor U8229 (N_8229,N_7595,N_7010);
and U8230 (N_8230,N_7780,N_7467);
nor U8231 (N_8231,N_7452,N_7397);
xnor U8232 (N_8232,N_7876,N_7200);
nand U8233 (N_8233,N_7718,N_7737);
nor U8234 (N_8234,N_7429,N_7250);
nand U8235 (N_8235,N_7998,N_7097);
and U8236 (N_8236,N_7574,N_7212);
xnor U8237 (N_8237,N_7749,N_7055);
nor U8238 (N_8238,N_7553,N_7252);
or U8239 (N_8239,N_7618,N_7268);
nand U8240 (N_8240,N_7331,N_7428);
nor U8241 (N_8241,N_7577,N_7834);
nor U8242 (N_8242,N_7965,N_7742);
nand U8243 (N_8243,N_7898,N_7732);
nor U8244 (N_8244,N_7750,N_7937);
xor U8245 (N_8245,N_7431,N_7340);
or U8246 (N_8246,N_7007,N_7215);
and U8247 (N_8247,N_7332,N_7132);
nand U8248 (N_8248,N_7126,N_7717);
xnor U8249 (N_8249,N_7785,N_7690);
and U8250 (N_8250,N_7025,N_7226);
nor U8251 (N_8251,N_7520,N_7878);
xnor U8252 (N_8252,N_7189,N_7160);
nand U8253 (N_8253,N_7269,N_7640);
and U8254 (N_8254,N_7182,N_7602);
nand U8255 (N_8255,N_7444,N_7059);
xor U8256 (N_8256,N_7221,N_7531);
and U8257 (N_8257,N_7866,N_7894);
nand U8258 (N_8258,N_7381,N_7924);
xnor U8259 (N_8259,N_7693,N_7933);
xnor U8260 (N_8260,N_7653,N_7448);
xnor U8261 (N_8261,N_7649,N_7511);
and U8262 (N_8262,N_7904,N_7806);
nor U8263 (N_8263,N_7575,N_7953);
xor U8264 (N_8264,N_7776,N_7032);
nand U8265 (N_8265,N_7303,N_7884);
or U8266 (N_8266,N_7979,N_7917);
or U8267 (N_8267,N_7562,N_7048);
and U8268 (N_8268,N_7447,N_7681);
or U8269 (N_8269,N_7325,N_7179);
nor U8270 (N_8270,N_7453,N_7318);
nor U8271 (N_8271,N_7615,N_7551);
nor U8272 (N_8272,N_7151,N_7508);
nor U8273 (N_8273,N_7961,N_7838);
nand U8274 (N_8274,N_7076,N_7679);
xnor U8275 (N_8275,N_7885,N_7787);
nand U8276 (N_8276,N_7643,N_7027);
and U8277 (N_8277,N_7537,N_7142);
and U8278 (N_8278,N_7102,N_7438);
xnor U8279 (N_8279,N_7664,N_7054);
xor U8280 (N_8280,N_7809,N_7354);
or U8281 (N_8281,N_7567,N_7794);
or U8282 (N_8282,N_7106,N_7078);
xnor U8283 (N_8283,N_7981,N_7020);
nor U8284 (N_8284,N_7107,N_7967);
xor U8285 (N_8285,N_7462,N_7880);
xnor U8286 (N_8286,N_7552,N_7727);
nand U8287 (N_8287,N_7777,N_7828);
nor U8288 (N_8288,N_7187,N_7320);
nand U8289 (N_8289,N_7152,N_7349);
nand U8290 (N_8290,N_7616,N_7436);
nor U8291 (N_8291,N_7758,N_7338);
xor U8292 (N_8292,N_7148,N_7379);
nor U8293 (N_8293,N_7154,N_7201);
or U8294 (N_8294,N_7940,N_7793);
nand U8295 (N_8295,N_7748,N_7256);
xnor U8296 (N_8296,N_7418,N_7941);
nand U8297 (N_8297,N_7582,N_7639);
xor U8298 (N_8298,N_7049,N_7987);
xnor U8299 (N_8299,N_7267,N_7736);
nor U8300 (N_8300,N_7619,N_7962);
and U8301 (N_8301,N_7931,N_7844);
nand U8302 (N_8302,N_7589,N_7738);
nand U8303 (N_8303,N_7757,N_7645);
nand U8304 (N_8304,N_7222,N_7412);
nor U8305 (N_8305,N_7368,N_7018);
nand U8306 (N_8306,N_7280,N_7724);
nand U8307 (N_8307,N_7417,N_7515);
nand U8308 (N_8308,N_7779,N_7790);
nand U8309 (N_8309,N_7960,N_7610);
and U8310 (N_8310,N_7014,N_7754);
xnor U8311 (N_8311,N_7237,N_7483);
and U8312 (N_8312,N_7420,N_7082);
nand U8313 (N_8313,N_7601,N_7519);
and U8314 (N_8314,N_7192,N_7778);
nor U8315 (N_8315,N_7622,N_7041);
nor U8316 (N_8316,N_7166,N_7127);
nor U8317 (N_8317,N_7532,N_7311);
or U8318 (N_8318,N_7270,N_7137);
xor U8319 (N_8319,N_7698,N_7853);
nor U8320 (N_8320,N_7021,N_7999);
and U8321 (N_8321,N_7457,N_7930);
xnor U8322 (N_8322,N_7801,N_7347);
and U8323 (N_8323,N_7131,N_7591);
nor U8324 (N_8324,N_7285,N_7695);
and U8325 (N_8325,N_7922,N_7781);
nor U8326 (N_8326,N_7371,N_7476);
xnor U8327 (N_8327,N_7424,N_7355);
nor U8328 (N_8328,N_7246,N_7903);
and U8329 (N_8329,N_7831,N_7963);
or U8330 (N_8330,N_7751,N_7888);
nand U8331 (N_8331,N_7275,N_7430);
and U8332 (N_8332,N_7451,N_7277);
nor U8333 (N_8333,N_7701,N_7756);
or U8334 (N_8334,N_7889,N_7336);
nor U8335 (N_8335,N_7951,N_7295);
nor U8336 (N_8336,N_7008,N_7110);
xor U8337 (N_8337,N_7803,N_7766);
or U8338 (N_8338,N_7548,N_7004);
nor U8339 (N_8339,N_7811,N_7047);
xor U8340 (N_8340,N_7666,N_7599);
and U8341 (N_8341,N_7568,N_7398);
nand U8342 (N_8342,N_7220,N_7557);
xnor U8343 (N_8343,N_7228,N_7015);
xnor U8344 (N_8344,N_7017,N_7175);
and U8345 (N_8345,N_7402,N_7841);
xor U8346 (N_8346,N_7968,N_7199);
and U8347 (N_8347,N_7079,N_7945);
xor U8348 (N_8348,N_7040,N_7648);
xor U8349 (N_8349,N_7286,N_7527);
or U8350 (N_8350,N_7897,N_7118);
or U8351 (N_8351,N_7711,N_7330);
or U8352 (N_8352,N_7456,N_7024);
nand U8353 (N_8353,N_7600,N_7378);
nor U8354 (N_8354,N_7948,N_7092);
or U8355 (N_8355,N_7044,N_7450);
nand U8356 (N_8356,N_7253,N_7946);
xor U8357 (N_8357,N_7860,N_7683);
and U8358 (N_8358,N_7652,N_7489);
and U8359 (N_8359,N_7125,N_7762);
nor U8360 (N_8360,N_7487,N_7804);
nor U8361 (N_8361,N_7216,N_7494);
or U8362 (N_8362,N_7374,N_7686);
or U8363 (N_8363,N_7725,N_7540);
xnor U8364 (N_8364,N_7879,N_7314);
and U8365 (N_8365,N_7484,N_7470);
xnor U8366 (N_8366,N_7419,N_7710);
nand U8367 (N_8367,N_7065,N_7544);
nor U8368 (N_8368,N_7393,N_7437);
and U8369 (N_8369,N_7207,N_7592);
nand U8370 (N_8370,N_7864,N_7588);
and U8371 (N_8371,N_7217,N_7161);
and U8372 (N_8372,N_7913,N_7939);
and U8373 (N_8373,N_7479,N_7056);
nand U8374 (N_8374,N_7036,N_7471);
xor U8375 (N_8375,N_7835,N_7375);
and U8376 (N_8376,N_7382,N_7687);
xor U8377 (N_8377,N_7254,N_7308);
or U8378 (N_8378,N_7294,N_7143);
and U8379 (N_8379,N_7003,N_7366);
nand U8380 (N_8380,N_7465,N_7289);
xnor U8381 (N_8381,N_7542,N_7909);
or U8382 (N_8382,N_7842,N_7350);
or U8383 (N_8383,N_7309,N_7706);
or U8384 (N_8384,N_7613,N_7081);
and U8385 (N_8385,N_7914,N_7316);
and U8386 (N_8386,N_7288,N_7530);
nor U8387 (N_8387,N_7873,N_7583);
nand U8388 (N_8388,N_7172,N_7721);
nand U8389 (N_8389,N_7074,N_7674);
and U8390 (N_8390,N_7121,N_7328);
or U8391 (N_8391,N_7404,N_7461);
nor U8392 (N_8392,N_7323,N_7673);
and U8393 (N_8393,N_7995,N_7287);
or U8394 (N_8394,N_7572,N_7449);
nor U8395 (N_8395,N_7672,N_7401);
nor U8396 (N_8396,N_7365,N_7383);
and U8397 (N_8397,N_7994,N_7839);
or U8398 (N_8398,N_7186,N_7578);
xor U8399 (N_8399,N_7824,N_7862);
or U8400 (N_8400,N_7584,N_7805);
xor U8401 (N_8401,N_7258,N_7463);
nand U8402 (N_8402,N_7680,N_7647);
nand U8403 (N_8403,N_7966,N_7096);
xor U8404 (N_8404,N_7833,N_7915);
and U8405 (N_8405,N_7119,N_7659);
nand U8406 (N_8406,N_7077,N_7173);
and U8407 (N_8407,N_7752,N_7662);
and U8408 (N_8408,N_7934,N_7813);
nand U8409 (N_8409,N_7670,N_7667);
and U8410 (N_8410,N_7315,N_7115);
and U8411 (N_8411,N_7539,N_7408);
nand U8412 (N_8412,N_7590,N_7919);
nor U8413 (N_8413,N_7414,N_7669);
or U8414 (N_8414,N_7677,N_7276);
nand U8415 (N_8415,N_7390,N_7569);
nor U8416 (N_8416,N_7703,N_7528);
xnor U8417 (N_8417,N_7006,N_7768);
or U8418 (N_8418,N_7482,N_7149);
xnor U8419 (N_8419,N_7682,N_7996);
xnor U8420 (N_8420,N_7808,N_7848);
nor U8421 (N_8421,N_7775,N_7852);
nor U8422 (N_8422,N_7676,N_7038);
or U8423 (N_8423,N_7855,N_7514);
xnor U8424 (N_8424,N_7053,N_7360);
and U8425 (N_8425,N_7989,N_7858);
nand U8426 (N_8426,N_7284,N_7518);
xor U8427 (N_8427,N_7871,N_7243);
nand U8428 (N_8428,N_7026,N_7956);
and U8429 (N_8429,N_7526,N_7459);
xnor U8430 (N_8430,N_7992,N_7245);
or U8431 (N_8431,N_7745,N_7959);
nand U8432 (N_8432,N_7707,N_7910);
and U8433 (N_8433,N_7982,N_7955);
nand U8434 (N_8434,N_7950,N_7555);
nand U8435 (N_8435,N_7134,N_7743);
nand U8436 (N_8436,N_7716,N_7625);
xnor U8437 (N_8437,N_7367,N_7812);
and U8438 (N_8438,N_7485,N_7304);
nor U8439 (N_8439,N_7868,N_7236);
or U8440 (N_8440,N_7503,N_7272);
nand U8441 (N_8441,N_7164,N_7596);
xnor U8442 (N_8442,N_7133,N_7144);
nand U8443 (N_8443,N_7517,N_7203);
or U8444 (N_8444,N_7472,N_7883);
xor U8445 (N_8445,N_7529,N_7095);
nor U8446 (N_8446,N_7571,N_7546);
nor U8447 (N_8447,N_7370,N_7867);
xnor U8448 (N_8448,N_7136,N_7016);
and U8449 (N_8449,N_7174,N_7791);
xnor U8450 (N_8450,N_7558,N_7797);
and U8451 (N_8451,N_7890,N_7351);
or U8452 (N_8452,N_7656,N_7905);
xnor U8453 (N_8453,N_7523,N_7150);
or U8454 (N_8454,N_7147,N_7493);
xnor U8455 (N_8455,N_7554,N_7814);
nor U8456 (N_8456,N_7604,N_7549);
or U8457 (N_8457,N_7863,N_7927);
nand U8458 (N_8458,N_7728,N_7263);
xnor U8459 (N_8459,N_7407,N_7130);
and U8460 (N_8460,N_7661,N_7614);
nand U8461 (N_8461,N_7509,N_7739);
nor U8462 (N_8462,N_7409,N_7060);
nand U8463 (N_8463,N_7547,N_7699);
or U8464 (N_8464,N_7594,N_7274);
nand U8465 (N_8465,N_7261,N_7334);
or U8466 (N_8466,N_7892,N_7545);
xor U8467 (N_8467,N_7906,N_7730);
xnor U8468 (N_8468,N_7603,N_7497);
or U8469 (N_8469,N_7312,N_7516);
nor U8470 (N_8470,N_7305,N_7139);
nor U8471 (N_8471,N_7480,N_7851);
and U8472 (N_8472,N_7696,N_7491);
and U8473 (N_8473,N_7985,N_7460);
or U8474 (N_8474,N_7362,N_7859);
and U8475 (N_8475,N_7566,N_7807);
nor U8476 (N_8476,N_7942,N_7260);
or U8477 (N_8477,N_7434,N_7795);
xnor U8478 (N_8478,N_7242,N_7823);
and U8479 (N_8479,N_7218,N_7159);
nand U8480 (N_8480,N_7084,N_7637);
and U8481 (N_8481,N_7248,N_7162);
nand U8482 (N_8482,N_7091,N_7935);
nor U8483 (N_8483,N_7190,N_7410);
nor U8484 (N_8484,N_7415,N_7391);
xnor U8485 (N_8485,N_7403,N_7896);
and U8486 (N_8486,N_7072,N_7327);
or U8487 (N_8487,N_7363,N_7747);
nand U8488 (N_8488,N_7080,N_7534);
nor U8489 (N_8489,N_7198,N_7947);
and U8490 (N_8490,N_7506,N_7694);
and U8491 (N_8491,N_7113,N_7911);
or U8492 (N_8492,N_7052,N_7856);
nor U8493 (N_8493,N_7406,N_7810);
and U8494 (N_8494,N_7907,N_7310);
nand U8495 (N_8495,N_7782,N_7920);
or U8496 (N_8496,N_7293,N_7783);
nand U8497 (N_8497,N_7655,N_7100);
nand U8498 (N_8498,N_7063,N_7348);
nor U8499 (N_8499,N_7726,N_7181);
xnor U8500 (N_8500,N_7942,N_7209);
nor U8501 (N_8501,N_7568,N_7887);
and U8502 (N_8502,N_7919,N_7034);
nand U8503 (N_8503,N_7805,N_7743);
nand U8504 (N_8504,N_7474,N_7913);
nor U8505 (N_8505,N_7796,N_7855);
nor U8506 (N_8506,N_7350,N_7675);
nand U8507 (N_8507,N_7122,N_7439);
nor U8508 (N_8508,N_7490,N_7649);
nand U8509 (N_8509,N_7801,N_7414);
nor U8510 (N_8510,N_7403,N_7261);
xnor U8511 (N_8511,N_7470,N_7902);
or U8512 (N_8512,N_7080,N_7170);
nor U8513 (N_8513,N_7915,N_7111);
or U8514 (N_8514,N_7813,N_7392);
xor U8515 (N_8515,N_7311,N_7679);
or U8516 (N_8516,N_7858,N_7299);
xor U8517 (N_8517,N_7496,N_7429);
and U8518 (N_8518,N_7867,N_7458);
and U8519 (N_8519,N_7851,N_7367);
xor U8520 (N_8520,N_7688,N_7293);
xor U8521 (N_8521,N_7493,N_7133);
xor U8522 (N_8522,N_7199,N_7830);
nor U8523 (N_8523,N_7749,N_7000);
xor U8524 (N_8524,N_7268,N_7643);
nand U8525 (N_8525,N_7224,N_7504);
and U8526 (N_8526,N_7903,N_7906);
nand U8527 (N_8527,N_7784,N_7679);
nand U8528 (N_8528,N_7268,N_7654);
or U8529 (N_8529,N_7431,N_7595);
or U8530 (N_8530,N_7953,N_7156);
xor U8531 (N_8531,N_7121,N_7379);
and U8532 (N_8532,N_7432,N_7839);
nand U8533 (N_8533,N_7010,N_7520);
nor U8534 (N_8534,N_7556,N_7230);
nor U8535 (N_8535,N_7208,N_7825);
and U8536 (N_8536,N_7514,N_7143);
nor U8537 (N_8537,N_7871,N_7792);
xnor U8538 (N_8538,N_7802,N_7283);
nand U8539 (N_8539,N_7363,N_7569);
or U8540 (N_8540,N_7383,N_7212);
or U8541 (N_8541,N_7730,N_7740);
nand U8542 (N_8542,N_7248,N_7750);
or U8543 (N_8543,N_7992,N_7526);
nand U8544 (N_8544,N_7000,N_7317);
nor U8545 (N_8545,N_7837,N_7247);
nand U8546 (N_8546,N_7124,N_7102);
nand U8547 (N_8547,N_7548,N_7527);
nand U8548 (N_8548,N_7407,N_7205);
nor U8549 (N_8549,N_7542,N_7491);
xnor U8550 (N_8550,N_7284,N_7645);
or U8551 (N_8551,N_7688,N_7444);
nand U8552 (N_8552,N_7527,N_7589);
or U8553 (N_8553,N_7025,N_7848);
or U8554 (N_8554,N_7775,N_7771);
and U8555 (N_8555,N_7059,N_7463);
nor U8556 (N_8556,N_7954,N_7188);
and U8557 (N_8557,N_7768,N_7631);
and U8558 (N_8558,N_7624,N_7206);
nor U8559 (N_8559,N_7566,N_7436);
or U8560 (N_8560,N_7726,N_7951);
and U8561 (N_8561,N_7303,N_7741);
nor U8562 (N_8562,N_7044,N_7679);
nor U8563 (N_8563,N_7874,N_7733);
or U8564 (N_8564,N_7536,N_7090);
xor U8565 (N_8565,N_7322,N_7758);
nor U8566 (N_8566,N_7739,N_7158);
nand U8567 (N_8567,N_7419,N_7260);
and U8568 (N_8568,N_7425,N_7360);
nor U8569 (N_8569,N_7824,N_7302);
or U8570 (N_8570,N_7939,N_7269);
nor U8571 (N_8571,N_7656,N_7663);
nand U8572 (N_8572,N_7113,N_7063);
and U8573 (N_8573,N_7247,N_7149);
and U8574 (N_8574,N_7410,N_7267);
and U8575 (N_8575,N_7863,N_7125);
or U8576 (N_8576,N_7478,N_7743);
or U8577 (N_8577,N_7645,N_7312);
and U8578 (N_8578,N_7731,N_7593);
xnor U8579 (N_8579,N_7156,N_7929);
nor U8580 (N_8580,N_7350,N_7949);
nor U8581 (N_8581,N_7844,N_7606);
nand U8582 (N_8582,N_7999,N_7935);
or U8583 (N_8583,N_7547,N_7386);
nand U8584 (N_8584,N_7354,N_7797);
nor U8585 (N_8585,N_7146,N_7846);
nand U8586 (N_8586,N_7976,N_7320);
xnor U8587 (N_8587,N_7405,N_7712);
nor U8588 (N_8588,N_7992,N_7081);
or U8589 (N_8589,N_7597,N_7341);
or U8590 (N_8590,N_7164,N_7173);
xor U8591 (N_8591,N_7171,N_7452);
nor U8592 (N_8592,N_7005,N_7344);
and U8593 (N_8593,N_7543,N_7739);
or U8594 (N_8594,N_7298,N_7402);
nand U8595 (N_8595,N_7432,N_7395);
nand U8596 (N_8596,N_7765,N_7371);
nand U8597 (N_8597,N_7329,N_7696);
and U8598 (N_8598,N_7714,N_7364);
and U8599 (N_8599,N_7740,N_7257);
or U8600 (N_8600,N_7421,N_7985);
nor U8601 (N_8601,N_7699,N_7422);
xnor U8602 (N_8602,N_7025,N_7752);
and U8603 (N_8603,N_7149,N_7726);
or U8604 (N_8604,N_7273,N_7285);
nand U8605 (N_8605,N_7163,N_7417);
xor U8606 (N_8606,N_7784,N_7374);
nand U8607 (N_8607,N_7741,N_7103);
nand U8608 (N_8608,N_7680,N_7201);
nor U8609 (N_8609,N_7080,N_7307);
or U8610 (N_8610,N_7847,N_7387);
or U8611 (N_8611,N_7761,N_7987);
xnor U8612 (N_8612,N_7043,N_7018);
nor U8613 (N_8613,N_7171,N_7258);
or U8614 (N_8614,N_7931,N_7705);
and U8615 (N_8615,N_7426,N_7859);
nand U8616 (N_8616,N_7328,N_7239);
nand U8617 (N_8617,N_7992,N_7881);
xnor U8618 (N_8618,N_7053,N_7139);
xor U8619 (N_8619,N_7529,N_7350);
nor U8620 (N_8620,N_7358,N_7469);
nor U8621 (N_8621,N_7794,N_7181);
xnor U8622 (N_8622,N_7810,N_7846);
or U8623 (N_8623,N_7788,N_7327);
or U8624 (N_8624,N_7267,N_7051);
nor U8625 (N_8625,N_7424,N_7480);
xnor U8626 (N_8626,N_7335,N_7559);
or U8627 (N_8627,N_7340,N_7324);
nand U8628 (N_8628,N_7737,N_7556);
and U8629 (N_8629,N_7501,N_7158);
nand U8630 (N_8630,N_7346,N_7750);
nand U8631 (N_8631,N_7195,N_7044);
or U8632 (N_8632,N_7027,N_7204);
or U8633 (N_8633,N_7902,N_7418);
xnor U8634 (N_8634,N_7771,N_7165);
or U8635 (N_8635,N_7662,N_7650);
nand U8636 (N_8636,N_7718,N_7138);
nand U8637 (N_8637,N_7901,N_7171);
xor U8638 (N_8638,N_7189,N_7724);
or U8639 (N_8639,N_7975,N_7588);
nand U8640 (N_8640,N_7199,N_7624);
xnor U8641 (N_8641,N_7962,N_7404);
and U8642 (N_8642,N_7230,N_7403);
nor U8643 (N_8643,N_7640,N_7965);
nor U8644 (N_8644,N_7517,N_7467);
and U8645 (N_8645,N_7911,N_7382);
xnor U8646 (N_8646,N_7820,N_7562);
nor U8647 (N_8647,N_7271,N_7656);
nor U8648 (N_8648,N_7820,N_7920);
nand U8649 (N_8649,N_7717,N_7932);
nor U8650 (N_8650,N_7536,N_7368);
xnor U8651 (N_8651,N_7231,N_7272);
nand U8652 (N_8652,N_7663,N_7154);
or U8653 (N_8653,N_7312,N_7484);
and U8654 (N_8654,N_7512,N_7537);
and U8655 (N_8655,N_7604,N_7459);
xnor U8656 (N_8656,N_7985,N_7447);
and U8657 (N_8657,N_7335,N_7761);
xor U8658 (N_8658,N_7878,N_7085);
or U8659 (N_8659,N_7927,N_7740);
nand U8660 (N_8660,N_7348,N_7622);
nand U8661 (N_8661,N_7848,N_7885);
and U8662 (N_8662,N_7613,N_7723);
or U8663 (N_8663,N_7981,N_7887);
nand U8664 (N_8664,N_7732,N_7617);
xor U8665 (N_8665,N_7859,N_7476);
and U8666 (N_8666,N_7903,N_7701);
or U8667 (N_8667,N_7992,N_7671);
nor U8668 (N_8668,N_7335,N_7286);
or U8669 (N_8669,N_7817,N_7698);
nor U8670 (N_8670,N_7005,N_7220);
xor U8671 (N_8671,N_7265,N_7020);
or U8672 (N_8672,N_7341,N_7196);
nand U8673 (N_8673,N_7530,N_7693);
and U8674 (N_8674,N_7850,N_7133);
and U8675 (N_8675,N_7212,N_7061);
nand U8676 (N_8676,N_7728,N_7848);
nor U8677 (N_8677,N_7065,N_7390);
and U8678 (N_8678,N_7533,N_7672);
xnor U8679 (N_8679,N_7212,N_7887);
or U8680 (N_8680,N_7866,N_7870);
or U8681 (N_8681,N_7382,N_7702);
or U8682 (N_8682,N_7399,N_7180);
nand U8683 (N_8683,N_7383,N_7523);
xnor U8684 (N_8684,N_7089,N_7485);
xor U8685 (N_8685,N_7443,N_7838);
and U8686 (N_8686,N_7779,N_7201);
or U8687 (N_8687,N_7723,N_7700);
or U8688 (N_8688,N_7509,N_7222);
nand U8689 (N_8689,N_7205,N_7014);
or U8690 (N_8690,N_7677,N_7911);
or U8691 (N_8691,N_7296,N_7374);
or U8692 (N_8692,N_7208,N_7439);
and U8693 (N_8693,N_7203,N_7743);
nand U8694 (N_8694,N_7187,N_7958);
nand U8695 (N_8695,N_7853,N_7764);
or U8696 (N_8696,N_7067,N_7821);
and U8697 (N_8697,N_7507,N_7619);
xor U8698 (N_8698,N_7485,N_7537);
nand U8699 (N_8699,N_7118,N_7299);
xnor U8700 (N_8700,N_7755,N_7587);
and U8701 (N_8701,N_7886,N_7113);
and U8702 (N_8702,N_7767,N_7585);
or U8703 (N_8703,N_7667,N_7436);
and U8704 (N_8704,N_7203,N_7840);
xor U8705 (N_8705,N_7020,N_7629);
nor U8706 (N_8706,N_7993,N_7077);
nand U8707 (N_8707,N_7668,N_7736);
nand U8708 (N_8708,N_7119,N_7082);
nor U8709 (N_8709,N_7006,N_7949);
nor U8710 (N_8710,N_7404,N_7062);
and U8711 (N_8711,N_7930,N_7052);
nand U8712 (N_8712,N_7302,N_7174);
or U8713 (N_8713,N_7616,N_7530);
xor U8714 (N_8714,N_7676,N_7967);
and U8715 (N_8715,N_7686,N_7491);
and U8716 (N_8716,N_7037,N_7522);
xor U8717 (N_8717,N_7161,N_7350);
nor U8718 (N_8718,N_7225,N_7056);
xnor U8719 (N_8719,N_7301,N_7164);
or U8720 (N_8720,N_7706,N_7374);
xor U8721 (N_8721,N_7623,N_7867);
and U8722 (N_8722,N_7884,N_7262);
and U8723 (N_8723,N_7455,N_7185);
nor U8724 (N_8724,N_7632,N_7358);
nor U8725 (N_8725,N_7984,N_7976);
or U8726 (N_8726,N_7355,N_7760);
and U8727 (N_8727,N_7835,N_7582);
or U8728 (N_8728,N_7178,N_7674);
nor U8729 (N_8729,N_7393,N_7050);
or U8730 (N_8730,N_7260,N_7723);
xor U8731 (N_8731,N_7273,N_7445);
nor U8732 (N_8732,N_7966,N_7789);
xor U8733 (N_8733,N_7769,N_7592);
xnor U8734 (N_8734,N_7763,N_7579);
nor U8735 (N_8735,N_7179,N_7191);
and U8736 (N_8736,N_7193,N_7076);
or U8737 (N_8737,N_7929,N_7796);
or U8738 (N_8738,N_7294,N_7091);
xnor U8739 (N_8739,N_7147,N_7175);
or U8740 (N_8740,N_7276,N_7233);
and U8741 (N_8741,N_7837,N_7827);
xor U8742 (N_8742,N_7075,N_7207);
xor U8743 (N_8743,N_7711,N_7561);
nor U8744 (N_8744,N_7207,N_7541);
nor U8745 (N_8745,N_7391,N_7041);
nand U8746 (N_8746,N_7729,N_7547);
xor U8747 (N_8747,N_7174,N_7756);
xor U8748 (N_8748,N_7964,N_7320);
nand U8749 (N_8749,N_7414,N_7290);
or U8750 (N_8750,N_7240,N_7273);
xnor U8751 (N_8751,N_7733,N_7181);
nand U8752 (N_8752,N_7409,N_7734);
nand U8753 (N_8753,N_7631,N_7051);
nor U8754 (N_8754,N_7489,N_7852);
nand U8755 (N_8755,N_7358,N_7113);
nor U8756 (N_8756,N_7003,N_7626);
or U8757 (N_8757,N_7124,N_7243);
nand U8758 (N_8758,N_7389,N_7247);
xor U8759 (N_8759,N_7666,N_7699);
nand U8760 (N_8760,N_7833,N_7539);
nor U8761 (N_8761,N_7375,N_7908);
and U8762 (N_8762,N_7068,N_7460);
and U8763 (N_8763,N_7584,N_7532);
nor U8764 (N_8764,N_7400,N_7314);
nor U8765 (N_8765,N_7653,N_7982);
and U8766 (N_8766,N_7002,N_7986);
or U8767 (N_8767,N_7594,N_7130);
nand U8768 (N_8768,N_7658,N_7887);
xnor U8769 (N_8769,N_7147,N_7291);
and U8770 (N_8770,N_7726,N_7967);
nand U8771 (N_8771,N_7613,N_7376);
and U8772 (N_8772,N_7771,N_7794);
nand U8773 (N_8773,N_7965,N_7867);
xnor U8774 (N_8774,N_7380,N_7493);
nand U8775 (N_8775,N_7448,N_7462);
or U8776 (N_8776,N_7057,N_7528);
or U8777 (N_8777,N_7024,N_7317);
and U8778 (N_8778,N_7207,N_7390);
and U8779 (N_8779,N_7635,N_7068);
nand U8780 (N_8780,N_7209,N_7768);
nand U8781 (N_8781,N_7116,N_7905);
nand U8782 (N_8782,N_7117,N_7470);
and U8783 (N_8783,N_7901,N_7291);
and U8784 (N_8784,N_7691,N_7770);
and U8785 (N_8785,N_7648,N_7109);
nand U8786 (N_8786,N_7093,N_7765);
and U8787 (N_8787,N_7709,N_7289);
nand U8788 (N_8788,N_7976,N_7971);
xnor U8789 (N_8789,N_7916,N_7892);
nor U8790 (N_8790,N_7158,N_7249);
xnor U8791 (N_8791,N_7985,N_7362);
or U8792 (N_8792,N_7357,N_7358);
nand U8793 (N_8793,N_7840,N_7174);
or U8794 (N_8794,N_7355,N_7133);
and U8795 (N_8795,N_7261,N_7581);
nand U8796 (N_8796,N_7454,N_7648);
xnor U8797 (N_8797,N_7922,N_7713);
nand U8798 (N_8798,N_7881,N_7618);
nor U8799 (N_8799,N_7103,N_7752);
nor U8800 (N_8800,N_7505,N_7295);
or U8801 (N_8801,N_7516,N_7131);
nand U8802 (N_8802,N_7712,N_7858);
xor U8803 (N_8803,N_7648,N_7092);
nor U8804 (N_8804,N_7412,N_7634);
nor U8805 (N_8805,N_7132,N_7154);
or U8806 (N_8806,N_7216,N_7992);
xor U8807 (N_8807,N_7336,N_7800);
or U8808 (N_8808,N_7023,N_7049);
xnor U8809 (N_8809,N_7545,N_7122);
or U8810 (N_8810,N_7916,N_7014);
nor U8811 (N_8811,N_7255,N_7279);
nor U8812 (N_8812,N_7914,N_7958);
or U8813 (N_8813,N_7758,N_7992);
xnor U8814 (N_8814,N_7189,N_7478);
or U8815 (N_8815,N_7961,N_7013);
and U8816 (N_8816,N_7189,N_7555);
nor U8817 (N_8817,N_7386,N_7182);
and U8818 (N_8818,N_7847,N_7985);
or U8819 (N_8819,N_7325,N_7301);
nand U8820 (N_8820,N_7344,N_7742);
nand U8821 (N_8821,N_7613,N_7060);
or U8822 (N_8822,N_7246,N_7664);
nand U8823 (N_8823,N_7581,N_7608);
and U8824 (N_8824,N_7411,N_7732);
and U8825 (N_8825,N_7658,N_7725);
or U8826 (N_8826,N_7328,N_7452);
and U8827 (N_8827,N_7383,N_7038);
nor U8828 (N_8828,N_7943,N_7341);
or U8829 (N_8829,N_7921,N_7419);
or U8830 (N_8830,N_7498,N_7336);
nor U8831 (N_8831,N_7751,N_7315);
or U8832 (N_8832,N_7043,N_7762);
xnor U8833 (N_8833,N_7581,N_7661);
or U8834 (N_8834,N_7598,N_7778);
nor U8835 (N_8835,N_7476,N_7005);
and U8836 (N_8836,N_7304,N_7966);
xnor U8837 (N_8837,N_7919,N_7319);
nand U8838 (N_8838,N_7517,N_7682);
and U8839 (N_8839,N_7188,N_7323);
or U8840 (N_8840,N_7848,N_7426);
nand U8841 (N_8841,N_7997,N_7517);
nor U8842 (N_8842,N_7004,N_7528);
nor U8843 (N_8843,N_7805,N_7950);
and U8844 (N_8844,N_7813,N_7946);
or U8845 (N_8845,N_7509,N_7041);
nand U8846 (N_8846,N_7335,N_7627);
or U8847 (N_8847,N_7687,N_7783);
xnor U8848 (N_8848,N_7692,N_7260);
nor U8849 (N_8849,N_7221,N_7043);
or U8850 (N_8850,N_7366,N_7207);
nand U8851 (N_8851,N_7541,N_7382);
nand U8852 (N_8852,N_7633,N_7461);
nor U8853 (N_8853,N_7134,N_7195);
and U8854 (N_8854,N_7894,N_7570);
nand U8855 (N_8855,N_7118,N_7333);
xnor U8856 (N_8856,N_7950,N_7316);
nor U8857 (N_8857,N_7148,N_7192);
xnor U8858 (N_8858,N_7635,N_7820);
nor U8859 (N_8859,N_7412,N_7843);
nor U8860 (N_8860,N_7935,N_7901);
and U8861 (N_8861,N_7467,N_7705);
and U8862 (N_8862,N_7842,N_7677);
xnor U8863 (N_8863,N_7311,N_7151);
nand U8864 (N_8864,N_7356,N_7798);
nand U8865 (N_8865,N_7231,N_7781);
and U8866 (N_8866,N_7441,N_7555);
or U8867 (N_8867,N_7920,N_7348);
nand U8868 (N_8868,N_7430,N_7952);
and U8869 (N_8869,N_7553,N_7643);
nor U8870 (N_8870,N_7082,N_7046);
and U8871 (N_8871,N_7335,N_7326);
or U8872 (N_8872,N_7870,N_7331);
and U8873 (N_8873,N_7878,N_7661);
or U8874 (N_8874,N_7922,N_7170);
and U8875 (N_8875,N_7583,N_7671);
nand U8876 (N_8876,N_7846,N_7766);
nor U8877 (N_8877,N_7161,N_7682);
xor U8878 (N_8878,N_7781,N_7001);
nand U8879 (N_8879,N_7744,N_7521);
and U8880 (N_8880,N_7685,N_7045);
and U8881 (N_8881,N_7442,N_7629);
or U8882 (N_8882,N_7299,N_7291);
nor U8883 (N_8883,N_7638,N_7709);
xor U8884 (N_8884,N_7811,N_7822);
and U8885 (N_8885,N_7697,N_7030);
nand U8886 (N_8886,N_7013,N_7318);
and U8887 (N_8887,N_7641,N_7688);
xor U8888 (N_8888,N_7817,N_7912);
or U8889 (N_8889,N_7335,N_7989);
and U8890 (N_8890,N_7587,N_7889);
nand U8891 (N_8891,N_7262,N_7740);
nor U8892 (N_8892,N_7114,N_7408);
nor U8893 (N_8893,N_7032,N_7676);
nand U8894 (N_8894,N_7010,N_7961);
or U8895 (N_8895,N_7252,N_7842);
or U8896 (N_8896,N_7621,N_7278);
nand U8897 (N_8897,N_7075,N_7810);
nand U8898 (N_8898,N_7598,N_7283);
nor U8899 (N_8899,N_7109,N_7341);
and U8900 (N_8900,N_7458,N_7456);
xor U8901 (N_8901,N_7244,N_7223);
nand U8902 (N_8902,N_7531,N_7944);
nand U8903 (N_8903,N_7374,N_7453);
or U8904 (N_8904,N_7157,N_7770);
or U8905 (N_8905,N_7850,N_7697);
and U8906 (N_8906,N_7191,N_7431);
or U8907 (N_8907,N_7287,N_7065);
nand U8908 (N_8908,N_7170,N_7660);
and U8909 (N_8909,N_7802,N_7476);
nor U8910 (N_8910,N_7636,N_7614);
nand U8911 (N_8911,N_7455,N_7408);
nor U8912 (N_8912,N_7178,N_7115);
xnor U8913 (N_8913,N_7724,N_7092);
nand U8914 (N_8914,N_7546,N_7442);
nand U8915 (N_8915,N_7441,N_7072);
and U8916 (N_8916,N_7291,N_7188);
and U8917 (N_8917,N_7766,N_7547);
or U8918 (N_8918,N_7218,N_7557);
and U8919 (N_8919,N_7450,N_7956);
and U8920 (N_8920,N_7688,N_7668);
xor U8921 (N_8921,N_7352,N_7667);
and U8922 (N_8922,N_7717,N_7203);
or U8923 (N_8923,N_7327,N_7346);
nor U8924 (N_8924,N_7579,N_7278);
nor U8925 (N_8925,N_7215,N_7706);
nand U8926 (N_8926,N_7561,N_7807);
or U8927 (N_8927,N_7413,N_7258);
nor U8928 (N_8928,N_7066,N_7202);
nor U8929 (N_8929,N_7815,N_7150);
or U8930 (N_8930,N_7512,N_7613);
or U8931 (N_8931,N_7865,N_7171);
xnor U8932 (N_8932,N_7196,N_7809);
and U8933 (N_8933,N_7033,N_7481);
or U8934 (N_8934,N_7895,N_7140);
nand U8935 (N_8935,N_7472,N_7688);
xnor U8936 (N_8936,N_7858,N_7053);
nand U8937 (N_8937,N_7757,N_7344);
or U8938 (N_8938,N_7973,N_7692);
xnor U8939 (N_8939,N_7182,N_7450);
nand U8940 (N_8940,N_7294,N_7227);
and U8941 (N_8941,N_7548,N_7043);
xor U8942 (N_8942,N_7346,N_7330);
nand U8943 (N_8943,N_7702,N_7007);
xor U8944 (N_8944,N_7463,N_7646);
nand U8945 (N_8945,N_7677,N_7979);
xnor U8946 (N_8946,N_7402,N_7513);
nor U8947 (N_8947,N_7468,N_7667);
nand U8948 (N_8948,N_7528,N_7973);
or U8949 (N_8949,N_7342,N_7332);
nand U8950 (N_8950,N_7798,N_7720);
and U8951 (N_8951,N_7832,N_7176);
and U8952 (N_8952,N_7369,N_7233);
nor U8953 (N_8953,N_7225,N_7523);
nand U8954 (N_8954,N_7564,N_7552);
or U8955 (N_8955,N_7421,N_7350);
xor U8956 (N_8956,N_7160,N_7861);
nand U8957 (N_8957,N_7400,N_7971);
or U8958 (N_8958,N_7727,N_7977);
nor U8959 (N_8959,N_7402,N_7196);
and U8960 (N_8960,N_7070,N_7122);
and U8961 (N_8961,N_7859,N_7890);
xor U8962 (N_8962,N_7256,N_7764);
and U8963 (N_8963,N_7700,N_7102);
nor U8964 (N_8964,N_7155,N_7635);
nor U8965 (N_8965,N_7321,N_7688);
and U8966 (N_8966,N_7693,N_7841);
xor U8967 (N_8967,N_7226,N_7911);
and U8968 (N_8968,N_7316,N_7041);
nand U8969 (N_8969,N_7154,N_7577);
xor U8970 (N_8970,N_7108,N_7402);
nand U8971 (N_8971,N_7495,N_7081);
xor U8972 (N_8972,N_7562,N_7852);
and U8973 (N_8973,N_7794,N_7992);
or U8974 (N_8974,N_7036,N_7878);
nor U8975 (N_8975,N_7619,N_7601);
or U8976 (N_8976,N_7839,N_7325);
nand U8977 (N_8977,N_7351,N_7766);
xnor U8978 (N_8978,N_7821,N_7812);
and U8979 (N_8979,N_7017,N_7995);
or U8980 (N_8980,N_7502,N_7764);
or U8981 (N_8981,N_7622,N_7691);
nor U8982 (N_8982,N_7602,N_7286);
nor U8983 (N_8983,N_7802,N_7796);
nor U8984 (N_8984,N_7768,N_7889);
nand U8985 (N_8985,N_7279,N_7696);
nor U8986 (N_8986,N_7828,N_7832);
nor U8987 (N_8987,N_7154,N_7887);
xor U8988 (N_8988,N_7516,N_7667);
and U8989 (N_8989,N_7021,N_7587);
xnor U8990 (N_8990,N_7652,N_7997);
nand U8991 (N_8991,N_7118,N_7759);
and U8992 (N_8992,N_7585,N_7248);
nand U8993 (N_8993,N_7842,N_7508);
or U8994 (N_8994,N_7182,N_7941);
or U8995 (N_8995,N_7037,N_7078);
nor U8996 (N_8996,N_7994,N_7348);
nor U8997 (N_8997,N_7322,N_7324);
xor U8998 (N_8998,N_7342,N_7464);
nand U8999 (N_8999,N_7451,N_7504);
nor U9000 (N_9000,N_8458,N_8208);
or U9001 (N_9001,N_8845,N_8413);
nand U9002 (N_9002,N_8793,N_8888);
xor U9003 (N_9003,N_8966,N_8117);
nand U9004 (N_9004,N_8906,N_8228);
and U9005 (N_9005,N_8852,N_8249);
nor U9006 (N_9006,N_8119,N_8680);
nor U9007 (N_9007,N_8003,N_8835);
nor U9008 (N_9008,N_8843,N_8272);
xnor U9009 (N_9009,N_8085,N_8187);
and U9010 (N_9010,N_8065,N_8275);
nor U9011 (N_9011,N_8593,N_8647);
nand U9012 (N_9012,N_8252,N_8039);
or U9013 (N_9013,N_8436,N_8859);
nor U9014 (N_9014,N_8253,N_8712);
and U9015 (N_9015,N_8974,N_8659);
or U9016 (N_9016,N_8081,N_8388);
and U9017 (N_9017,N_8056,N_8274);
or U9018 (N_9018,N_8491,N_8842);
xor U9019 (N_9019,N_8507,N_8692);
or U9020 (N_9020,N_8131,N_8070);
or U9021 (N_9021,N_8244,N_8331);
or U9022 (N_9022,N_8213,N_8876);
or U9023 (N_9023,N_8444,N_8041);
and U9024 (N_9024,N_8433,N_8267);
or U9025 (N_9025,N_8754,N_8541);
xor U9026 (N_9026,N_8828,N_8989);
or U9027 (N_9027,N_8199,N_8320);
and U9028 (N_9028,N_8701,N_8600);
xnor U9029 (N_9029,N_8172,N_8094);
nor U9030 (N_9030,N_8024,N_8072);
and U9031 (N_9031,N_8825,N_8457);
nand U9032 (N_9032,N_8245,N_8711);
nand U9033 (N_9033,N_8751,N_8703);
nor U9034 (N_9034,N_8202,N_8145);
xor U9035 (N_9035,N_8561,N_8690);
or U9036 (N_9036,N_8826,N_8585);
or U9037 (N_9037,N_8391,N_8919);
or U9038 (N_9038,N_8717,N_8519);
xnor U9039 (N_9039,N_8494,N_8053);
nor U9040 (N_9040,N_8424,N_8903);
nand U9041 (N_9041,N_8667,N_8300);
nand U9042 (N_9042,N_8222,N_8995);
nand U9043 (N_9043,N_8753,N_8658);
xor U9044 (N_9044,N_8184,N_8892);
nand U9045 (N_9045,N_8881,N_8676);
xnor U9046 (N_9046,N_8018,N_8908);
and U9047 (N_9047,N_8454,N_8231);
nor U9048 (N_9048,N_8428,N_8955);
xnor U9049 (N_9049,N_8582,N_8517);
nor U9050 (N_9050,N_8084,N_8833);
nand U9051 (N_9051,N_8653,N_8118);
nand U9052 (N_9052,N_8087,N_8720);
xnor U9053 (N_9053,N_8130,N_8101);
nand U9054 (N_9054,N_8339,N_8716);
or U9055 (N_9055,N_8107,N_8029);
nand U9056 (N_9056,N_8788,N_8277);
xor U9057 (N_9057,N_8031,N_8856);
xnor U9058 (N_9058,N_8235,N_8013);
or U9059 (N_9059,N_8884,N_8104);
or U9060 (N_9060,N_8142,N_8971);
or U9061 (N_9061,N_8322,N_8488);
or U9062 (N_9062,N_8838,N_8465);
and U9063 (N_9063,N_8344,N_8779);
or U9064 (N_9064,N_8907,N_8451);
xnor U9065 (N_9065,N_8103,N_8991);
nand U9066 (N_9066,N_8347,N_8550);
nand U9067 (N_9067,N_8940,N_8067);
nor U9068 (N_9068,N_8238,N_8006);
or U9069 (N_9069,N_8257,N_8318);
and U9070 (N_9070,N_8951,N_8448);
nor U9071 (N_9071,N_8446,N_8193);
nand U9072 (N_9072,N_8891,N_8401);
xnor U9073 (N_9073,N_8564,N_8254);
nand U9074 (N_9074,N_8863,N_8175);
or U9075 (N_9075,N_8399,N_8250);
xnor U9076 (N_9076,N_8742,N_8513);
xnor U9077 (N_9077,N_8981,N_8821);
and U9078 (N_9078,N_8261,N_8894);
or U9079 (N_9079,N_8189,N_8468);
nand U9080 (N_9080,N_8554,N_8850);
or U9081 (N_9081,N_8303,N_8707);
xnor U9082 (N_9082,N_8555,N_8675);
xnor U9083 (N_9083,N_8030,N_8663);
xnor U9084 (N_9084,N_8594,N_8325);
or U9085 (N_9085,N_8738,N_8535);
nand U9086 (N_9086,N_8719,N_8950);
xor U9087 (N_9087,N_8048,N_8122);
nor U9088 (N_9088,N_8196,N_8452);
or U9089 (N_9089,N_8141,N_8326);
and U9090 (N_9090,N_8685,N_8670);
and U9091 (N_9091,N_8755,N_8483);
nand U9092 (N_9092,N_8882,N_8607);
nand U9093 (N_9093,N_8480,N_8918);
nor U9094 (N_9094,N_8686,N_8233);
xnor U9095 (N_9095,N_8410,N_8724);
nand U9096 (N_9096,N_8419,N_8800);
nor U9097 (N_9097,N_8167,N_8210);
nand U9098 (N_9098,N_8999,N_8774);
xnor U9099 (N_9099,N_8256,N_8740);
nand U9100 (N_9100,N_8731,N_8666);
nor U9101 (N_9101,N_8571,N_8434);
nor U9102 (N_9102,N_8460,N_8808);
xor U9103 (N_9103,N_8425,N_8371);
nor U9104 (N_9104,N_8350,N_8080);
nand U9105 (N_9105,N_8781,N_8660);
nor U9106 (N_9106,N_8022,N_8572);
nand U9107 (N_9107,N_8563,N_8962);
nor U9108 (N_9108,N_8931,N_8602);
xnor U9109 (N_9109,N_8886,N_8185);
and U9110 (N_9110,N_8694,N_8083);
or U9111 (N_9111,N_8289,N_8035);
or U9112 (N_9112,N_8920,N_8477);
nand U9113 (N_9113,N_8033,N_8832);
or U9114 (N_9114,N_8916,N_8868);
and U9115 (N_9115,N_8327,N_8551);
and U9116 (N_9116,N_8552,N_8363);
or U9117 (N_9117,N_8534,N_8416);
and U9118 (N_9118,N_8569,N_8043);
or U9119 (N_9119,N_8268,N_8725);
xnor U9120 (N_9120,N_8062,N_8171);
nand U9121 (N_9121,N_8100,N_8328);
nand U9122 (N_9122,N_8759,N_8890);
or U9123 (N_9123,N_8664,N_8049);
nand U9124 (N_9124,N_8467,N_8713);
or U9125 (N_9125,N_8179,N_8540);
xor U9126 (N_9126,N_8040,N_8099);
and U9127 (N_9127,N_8234,N_8158);
xor U9128 (N_9128,N_8830,N_8478);
or U9129 (N_9129,N_8678,N_8873);
nand U9130 (N_9130,N_8217,N_8190);
and U9131 (N_9131,N_8246,N_8127);
or U9132 (N_9132,N_8381,N_8736);
and U9133 (N_9133,N_8046,N_8878);
or U9134 (N_9134,N_8064,N_8626);
xor U9135 (N_9135,N_8329,N_8744);
and U9136 (N_9136,N_8956,N_8204);
nand U9137 (N_9137,N_8604,N_8829);
or U9138 (N_9138,N_8503,N_8005);
xor U9139 (N_9139,N_8216,N_8532);
nand U9140 (N_9140,N_8575,N_8773);
or U9141 (N_9141,N_8687,N_8591);
nor U9142 (N_9142,N_8605,N_8314);
nor U9143 (N_9143,N_8449,N_8285);
nor U9144 (N_9144,N_8586,N_8954);
nor U9145 (N_9145,N_8553,N_8105);
or U9146 (N_9146,N_8521,N_8426);
nor U9147 (N_9147,N_8522,N_8967);
xor U9148 (N_9148,N_8927,N_8596);
or U9149 (N_9149,N_8860,N_8455);
xnor U9150 (N_9150,N_8932,N_8290);
nand U9151 (N_9151,N_8936,N_8674);
xnor U9152 (N_9152,N_8164,N_8182);
nand U9153 (N_9153,N_8269,N_8128);
nand U9154 (N_9154,N_8902,N_8473);
nand U9155 (N_9155,N_8078,N_8750);
nand U9156 (N_9156,N_8840,N_8224);
nor U9157 (N_9157,N_8370,N_8054);
nor U9158 (N_9158,N_8476,N_8437);
xor U9159 (N_9159,N_8923,N_8728);
or U9160 (N_9160,N_8806,N_8620);
nand U9161 (N_9161,N_8296,N_8549);
xnor U9162 (N_9162,N_8114,N_8280);
and U9163 (N_9163,N_8851,N_8215);
and U9164 (N_9164,N_8823,N_8362);
and U9165 (N_9165,N_8527,N_8125);
xnor U9166 (N_9166,N_8622,N_8461);
and U9167 (N_9167,N_8095,N_8952);
xnor U9168 (N_9168,N_8870,N_8520);
xnor U9169 (N_9169,N_8153,N_8565);
and U9170 (N_9170,N_8258,N_8163);
or U9171 (N_9171,N_8349,N_8079);
nor U9172 (N_9172,N_8273,N_8559);
xor U9173 (N_9173,N_8038,N_8696);
or U9174 (N_9174,N_8021,N_8880);
xor U9175 (N_9175,N_8305,N_8389);
xor U9176 (N_9176,N_8542,N_8827);
or U9177 (N_9177,N_8479,N_8803);
or U9178 (N_9178,N_8661,N_8722);
xor U9179 (N_9179,N_8695,N_8775);
nand U9180 (N_9180,N_8963,N_8338);
nor U9181 (N_9181,N_8140,N_8609);
nor U9182 (N_9182,N_8778,N_8760);
nand U9183 (N_9183,N_8718,N_8342);
nand U9184 (N_9184,N_8901,N_8904);
or U9185 (N_9185,N_8421,N_8510);
nor U9186 (N_9186,N_8621,N_8001);
and U9187 (N_9187,N_8983,N_8980);
and U9188 (N_9188,N_8058,N_8688);
nand U9189 (N_9189,N_8822,N_8945);
and U9190 (N_9190,N_8443,N_8914);
nand U9191 (N_9191,N_8958,N_8787);
xor U9192 (N_9192,N_8734,N_8283);
nand U9193 (N_9193,N_8281,N_8921);
xnor U9194 (N_9194,N_8929,N_8197);
and U9195 (N_9195,N_8745,N_8402);
xnor U9196 (N_9196,N_8807,N_8323);
nand U9197 (N_9197,N_8608,N_8797);
xor U9198 (N_9198,N_8059,N_8198);
or U9199 (N_9199,N_8612,N_8986);
nor U9200 (N_9200,N_8867,N_8544);
nor U9201 (N_9201,N_8294,N_8450);
nor U9202 (N_9202,N_8743,N_8340);
or U9203 (N_9203,N_8993,N_8547);
and U9204 (N_9204,N_8293,N_8581);
nand U9205 (N_9205,N_8149,N_8351);
or U9206 (N_9206,N_8475,N_8073);
nand U9207 (N_9207,N_8935,N_8108);
nor U9208 (N_9208,N_8166,N_8236);
nand U9209 (N_9209,N_8221,N_8247);
nand U9210 (N_9210,N_8648,N_8885);
and U9211 (N_9211,N_8764,N_8982);
or U9212 (N_9212,N_8007,N_8530);
and U9213 (N_9213,N_8627,N_8960);
and U9214 (N_9214,N_8637,N_8543);
nor U9215 (N_9215,N_8313,N_8700);
nor U9216 (N_9216,N_8137,N_8050);
and U9217 (N_9217,N_8404,N_8353);
and U9218 (N_9218,N_8495,N_8590);
nand U9219 (N_9219,N_8211,N_8506);
nor U9220 (N_9220,N_8136,N_8174);
and U9221 (N_9221,N_8384,N_8849);
and U9222 (N_9222,N_8802,N_8577);
and U9223 (N_9223,N_8156,N_8133);
xor U9224 (N_9224,N_8749,N_8203);
or U9225 (N_9225,N_8368,N_8372);
and U9226 (N_9226,N_8490,N_8933);
or U9227 (N_9227,N_8223,N_8299);
nor U9228 (N_9228,N_8529,N_8899);
nor U9229 (N_9229,N_8086,N_8624);
nand U9230 (N_9230,N_8943,N_8629);
nor U9231 (N_9231,N_8889,N_8191);
or U9232 (N_9232,N_8330,N_8747);
or U9233 (N_9233,N_8964,N_8599);
xnor U9234 (N_9234,N_8486,N_8017);
nand U9235 (N_9235,N_8106,N_8387);
and U9236 (N_9236,N_8896,N_8205);
and U9237 (N_9237,N_8589,N_8409);
or U9238 (N_9238,N_8335,N_8898);
nor U9239 (N_9239,N_8580,N_8874);
xor U9240 (N_9240,N_8592,N_8343);
nor U9241 (N_9241,N_8111,N_8855);
nand U9242 (N_9242,N_8310,N_8028);
nand U9243 (N_9243,N_8456,N_8518);
xnor U9244 (N_9244,N_8741,N_8121);
nor U9245 (N_9245,N_8809,N_8699);
xor U9246 (N_9246,N_8287,N_8373);
nor U9247 (N_9247,N_8110,N_8804);
xnor U9248 (N_9248,N_8308,N_8459);
or U9249 (N_9249,N_8525,N_8218);
nor U9250 (N_9250,N_8509,N_8173);
or U9251 (N_9251,N_8445,N_8500);
xnor U9252 (N_9252,N_8422,N_8392);
and U9253 (N_9253,N_8727,N_8374);
nor U9254 (N_9254,N_8973,N_8297);
and U9255 (N_9255,N_8656,N_8789);
nand U9256 (N_9256,N_8498,N_8526);
xnor U9257 (N_9257,N_8536,N_8192);
or U9258 (N_9258,N_8706,N_8390);
and U9259 (N_9259,N_8771,N_8533);
nand U9260 (N_9260,N_8034,N_8008);
or U9261 (N_9261,N_8630,N_8897);
nand U9262 (N_9262,N_8587,N_8693);
nand U9263 (N_9263,N_8412,N_8237);
and U9264 (N_9264,N_8776,N_8143);
xnor U9265 (N_9265,N_8523,N_8306);
nor U9266 (N_9266,N_8777,N_8669);
nand U9267 (N_9267,N_8464,N_8207);
or U9268 (N_9268,N_8922,N_8463);
xnor U9269 (N_9269,N_8866,N_8044);
and U9270 (N_9270,N_8912,N_8655);
nor U9271 (N_9271,N_8097,N_8438);
xnor U9272 (N_9272,N_8440,N_8453);
or U9273 (N_9273,N_8435,N_8834);
nand U9274 (N_9274,N_8934,N_8492);
nor U9275 (N_9275,N_8093,N_8474);
nand U9276 (N_9276,N_8255,N_8579);
and U9277 (N_9277,N_8841,N_8977);
xor U9278 (N_9278,N_8528,N_8248);
nor U9279 (N_9279,N_8472,N_8423);
xnor U9280 (N_9280,N_8970,N_8721);
xor U9281 (N_9281,N_8767,N_8004);
nor U9282 (N_9282,N_8795,N_8790);
and U9283 (N_9283,N_8176,N_8641);
and U9284 (N_9284,N_8139,N_8023);
nand U9285 (N_9285,N_8194,N_8941);
nor U9286 (N_9286,N_8937,N_8628);
xnor U9287 (N_9287,N_8784,N_8801);
nand U9288 (N_9288,N_8066,N_8877);
or U9289 (N_9289,N_8766,N_8161);
or U9290 (N_9290,N_8691,N_8109);
nor U9291 (N_9291,N_8848,N_8756);
nand U9292 (N_9292,N_8987,N_8539);
or U9293 (N_9293,N_8279,N_8853);
xor U9294 (N_9294,N_8124,N_8762);
or U9295 (N_9295,N_8112,N_8872);
and U9296 (N_9296,N_8824,N_8232);
and U9297 (N_9297,N_8225,N_8051);
or U9298 (N_9298,N_8869,N_8505);
or U9299 (N_9299,N_8016,N_8015);
nand U9300 (N_9300,N_8415,N_8556);
or U9301 (N_9301,N_8811,N_8441);
and U9302 (N_9302,N_8733,N_8512);
nor U9303 (N_9303,N_8566,N_8961);
and U9304 (N_9304,N_8689,N_8606);
nand U9305 (N_9305,N_8625,N_8430);
and U9306 (N_9306,N_8671,N_8113);
nor U9307 (N_9307,N_8180,N_8150);
nor U9308 (N_9308,N_8188,N_8568);
nor U9309 (N_9309,N_8643,N_8546);
xnor U9310 (N_9310,N_8905,N_8386);
xnor U9311 (N_9311,N_8729,N_8770);
or U9312 (N_9312,N_8270,N_8155);
xor U9313 (N_9313,N_8610,N_8146);
or U9314 (N_9314,N_8662,N_8939);
and U9315 (N_9315,N_8574,N_8515);
nand U9316 (N_9316,N_8096,N_8411);
and U9317 (N_9317,N_8723,N_8276);
or U9318 (N_9318,N_8996,N_8361);
nor U9319 (N_9319,N_8011,N_8915);
nand U9320 (N_9320,N_8603,N_8262);
or U9321 (N_9321,N_8944,N_8241);
xor U9322 (N_9322,N_8684,N_8705);
and U9323 (N_9323,N_8836,N_8168);
nor U9324 (N_9324,N_8780,N_8497);
xor U9325 (N_9325,N_8427,N_8036);
xnor U9326 (N_9326,N_8469,N_8082);
nand U9327 (N_9327,N_8938,N_8408);
nor U9328 (N_9328,N_8375,N_8129);
nand U9329 (N_9329,N_8239,N_8861);
nor U9330 (N_9330,N_8466,N_8900);
or U9331 (N_9331,N_8814,N_8893);
xnor U9332 (N_9332,N_8407,N_8895);
nand U9333 (N_9333,N_8414,N_8649);
or U9334 (N_9334,N_8639,N_8615);
and U9335 (N_9335,N_8794,N_8047);
or U9336 (N_9336,N_8052,N_8924);
or U9337 (N_9337,N_8442,N_8668);
nand U9338 (N_9338,N_8364,N_8819);
nor U9339 (N_9339,N_8489,N_8926);
and U9340 (N_9340,N_8682,N_8484);
or U9341 (N_9341,N_8617,N_8346);
nand U9342 (N_9342,N_8352,N_8854);
and U9343 (N_9343,N_8910,N_8169);
nor U9344 (N_9344,N_8965,N_8969);
or U9345 (N_9345,N_8948,N_8366);
or U9346 (N_9346,N_8000,N_8014);
nand U9347 (N_9347,N_8292,N_8462);
nand U9348 (N_9348,N_8644,N_8200);
nor U9349 (N_9349,N_8160,N_8786);
or U9350 (N_9350,N_8672,N_8116);
xnor U9351 (N_9351,N_8432,N_8398);
nor U9352 (N_9352,N_8077,N_8730);
or U9353 (N_9353,N_8165,N_8799);
or U9354 (N_9354,N_8831,N_8162);
or U9355 (N_9355,N_8531,N_8930);
nor U9356 (N_9356,N_8487,N_8642);
xor U9357 (N_9357,N_8504,N_8883);
nand U9358 (N_9358,N_8925,N_8220);
or U9359 (N_9359,N_8076,N_8037);
xnor U9360 (N_9360,N_8514,N_8345);
nand U9361 (N_9361,N_8714,N_8061);
and U9362 (N_9362,N_8471,N_8988);
nor U9363 (N_9363,N_8282,N_8357);
nor U9364 (N_9364,N_8012,N_8301);
and U9365 (N_9365,N_8942,N_8508);
xor U9366 (N_9366,N_8002,N_8321);
and U9367 (N_9367,N_8702,N_8619);
and U9368 (N_9368,N_8382,N_8286);
nor U9369 (N_9369,N_8025,N_8482);
or U9370 (N_9370,N_8772,N_8406);
nand U9371 (N_9371,N_8214,N_8148);
and U9372 (N_9372,N_8154,N_8356);
nand U9373 (N_9373,N_8126,N_8377);
nor U9374 (N_9374,N_8511,N_8151);
and U9375 (N_9375,N_8735,N_8481);
nor U9376 (N_9376,N_8710,N_8708);
and U9377 (N_9377,N_8545,N_8646);
and U9378 (N_9378,N_8578,N_8618);
and U9379 (N_9379,N_8645,N_8858);
and U9380 (N_9380,N_8369,N_8847);
nand U9381 (N_9381,N_8757,N_8560);
and U9382 (N_9382,N_8673,N_8635);
nor U9383 (N_9383,N_8782,N_8844);
and U9384 (N_9384,N_8752,N_8206);
nand U9385 (N_9385,N_8812,N_8769);
nor U9386 (N_9386,N_8573,N_8379);
nand U9387 (N_9387,N_8132,N_8557);
or U9388 (N_9388,N_8677,N_8558);
nand U9389 (N_9389,N_8229,N_8324);
nor U9390 (N_9390,N_8020,N_8470);
xnor U9391 (N_9391,N_8857,N_8651);
and U9392 (N_9392,N_8336,N_8997);
nand U9393 (N_9393,N_8820,N_8360);
nor U9394 (N_9394,N_8309,N_8726);
or U9395 (N_9395,N_8312,N_8201);
and U9396 (N_9396,N_8665,N_8538);
nor U9397 (N_9397,N_8611,N_8638);
xnor U9398 (N_9398,N_8177,N_8144);
nor U9399 (N_9399,N_8697,N_8068);
and U9400 (N_9400,N_8953,N_8123);
xor U9401 (N_9401,N_8209,N_8266);
xor U9402 (N_9402,N_8698,N_8818);
nor U9403 (N_9403,N_8798,N_8737);
and U9404 (N_9404,N_8791,N_8613);
or U9405 (N_9405,N_8887,N_8588);
and U9406 (N_9406,N_8746,N_8975);
nor U9407 (N_9407,N_8763,N_8075);
and U9408 (N_9408,N_8102,N_8385);
nand U9409 (N_9409,N_8055,N_8992);
xor U9410 (N_9410,N_8298,N_8976);
nor U9411 (N_9411,N_8524,N_8758);
and U9412 (N_9412,N_8378,N_8597);
and U9413 (N_9413,N_8367,N_8354);
nand U9414 (N_9414,N_8748,N_8315);
and U9415 (N_9415,N_8317,N_8288);
xnor U9416 (N_9416,N_8178,N_8816);
or U9417 (N_9417,N_8420,N_8623);
or U9418 (N_9418,N_8501,N_8089);
xnor U9419 (N_9419,N_8380,N_8447);
and U9420 (N_9420,N_8650,N_8226);
nor U9421 (N_9421,N_8365,N_8091);
nand U9422 (N_9422,N_8271,N_8957);
xnor U9423 (N_9423,N_8978,N_8092);
nand U9424 (N_9424,N_8251,N_8355);
xnor U9425 (N_9425,N_8376,N_8537);
nand U9426 (N_9426,N_8994,N_8567);
xor U9427 (N_9427,N_8010,N_8260);
nand U9428 (N_9428,N_8761,N_8098);
xnor U9429 (N_9429,N_8640,N_8295);
nand U9430 (N_9430,N_8071,N_8946);
and U9431 (N_9431,N_8418,N_8088);
or U9432 (N_9432,N_8074,N_8732);
and U9433 (N_9433,N_8243,N_8636);
xnor U9434 (N_9434,N_8333,N_8595);
and U9435 (N_9435,N_8120,N_8431);
or U9436 (N_9436,N_8348,N_8429);
nand U9437 (N_9437,N_8026,N_8278);
or U9438 (N_9438,N_8739,N_8291);
or U9439 (N_9439,N_8968,N_8496);
xor U9440 (N_9440,N_8947,N_8583);
and U9441 (N_9441,N_8069,N_8709);
nor U9442 (N_9442,N_8042,N_8383);
or U9443 (N_9443,N_8334,N_8186);
or U9444 (N_9444,N_8715,N_8159);
xor U9445 (N_9445,N_8959,N_8359);
xor U9446 (N_9446,N_8631,N_8400);
nor U9447 (N_9447,N_8240,N_8304);
xnor U9448 (N_9448,N_8439,N_8397);
nand U9449 (N_9449,N_8704,N_8307);
and U9450 (N_9450,N_8990,N_8570);
or U9451 (N_9451,N_8019,N_8837);
nand U9452 (N_9452,N_8810,N_8485);
nand U9453 (N_9453,N_8316,N_8032);
and U9454 (N_9454,N_8393,N_8768);
or U9455 (N_9455,N_8060,N_8057);
nand U9456 (N_9456,N_8633,N_8634);
xor U9457 (N_9457,N_8516,N_8548);
nor U9458 (N_9458,N_8792,N_8063);
nand U9459 (N_9459,N_8783,N_8871);
and U9460 (N_9460,N_8183,N_8115);
xor U9461 (N_9461,N_8212,N_8598);
nor U9462 (N_9462,N_8949,N_8817);
or U9463 (N_9463,N_8417,N_8027);
xor U9464 (N_9464,N_8805,N_8864);
xnor U9465 (N_9465,N_8311,N_8395);
nand U9466 (N_9466,N_8928,N_8138);
xnor U9467 (N_9467,N_8584,N_8135);
xnor U9468 (N_9468,N_8576,N_8601);
nor U9469 (N_9469,N_8265,N_8865);
or U9470 (N_9470,N_8839,N_8396);
nand U9471 (N_9471,N_8170,N_8230);
and U9472 (N_9472,N_8862,N_8332);
xnor U9473 (N_9473,N_8813,N_8219);
nand U9474 (N_9474,N_8909,N_8654);
or U9475 (N_9475,N_8998,N_8616);
nor U9476 (N_9476,N_8875,N_8652);
and U9477 (N_9477,N_8815,N_8341);
nor U9478 (N_9478,N_8614,N_8911);
and U9479 (N_9479,N_8493,N_8259);
nor U9480 (N_9480,N_8284,N_8134);
xnor U9481 (N_9481,N_8242,N_8683);
nand U9482 (N_9482,N_8337,N_8319);
nand U9483 (N_9483,N_8227,N_8681);
xnor U9484 (N_9484,N_8657,N_8263);
and U9485 (N_9485,N_8045,N_8403);
or U9486 (N_9486,N_8846,N_8765);
xor U9487 (N_9487,N_8152,N_8499);
xor U9488 (N_9488,N_8562,N_8502);
or U9489 (N_9489,N_8181,N_8632);
nor U9490 (N_9490,N_8157,N_8879);
nand U9491 (N_9491,N_8264,N_8984);
xor U9492 (N_9492,N_8796,N_8679);
xor U9493 (N_9493,N_8394,N_8302);
xnor U9494 (N_9494,N_8358,N_8972);
nor U9495 (N_9495,N_8917,N_8405);
nand U9496 (N_9496,N_8979,N_8090);
and U9497 (N_9497,N_8985,N_8913);
nand U9498 (N_9498,N_8147,N_8785);
and U9499 (N_9499,N_8195,N_8009);
nand U9500 (N_9500,N_8629,N_8980);
xnor U9501 (N_9501,N_8654,N_8787);
xnor U9502 (N_9502,N_8244,N_8673);
and U9503 (N_9503,N_8638,N_8930);
or U9504 (N_9504,N_8562,N_8929);
nor U9505 (N_9505,N_8851,N_8806);
nand U9506 (N_9506,N_8070,N_8455);
xor U9507 (N_9507,N_8438,N_8612);
and U9508 (N_9508,N_8940,N_8583);
or U9509 (N_9509,N_8418,N_8996);
nand U9510 (N_9510,N_8158,N_8903);
nand U9511 (N_9511,N_8565,N_8639);
and U9512 (N_9512,N_8831,N_8401);
nor U9513 (N_9513,N_8505,N_8720);
or U9514 (N_9514,N_8765,N_8236);
xor U9515 (N_9515,N_8037,N_8681);
and U9516 (N_9516,N_8019,N_8048);
and U9517 (N_9517,N_8610,N_8289);
and U9518 (N_9518,N_8815,N_8032);
or U9519 (N_9519,N_8194,N_8043);
nand U9520 (N_9520,N_8819,N_8800);
nand U9521 (N_9521,N_8110,N_8024);
xor U9522 (N_9522,N_8075,N_8620);
nand U9523 (N_9523,N_8431,N_8046);
xor U9524 (N_9524,N_8877,N_8377);
or U9525 (N_9525,N_8360,N_8393);
or U9526 (N_9526,N_8873,N_8074);
nand U9527 (N_9527,N_8454,N_8751);
or U9528 (N_9528,N_8736,N_8756);
or U9529 (N_9529,N_8568,N_8450);
xnor U9530 (N_9530,N_8232,N_8961);
and U9531 (N_9531,N_8011,N_8672);
nand U9532 (N_9532,N_8152,N_8935);
or U9533 (N_9533,N_8386,N_8942);
xor U9534 (N_9534,N_8331,N_8708);
nor U9535 (N_9535,N_8032,N_8840);
xnor U9536 (N_9536,N_8488,N_8460);
or U9537 (N_9537,N_8193,N_8136);
nand U9538 (N_9538,N_8855,N_8538);
nor U9539 (N_9539,N_8346,N_8818);
and U9540 (N_9540,N_8296,N_8976);
xor U9541 (N_9541,N_8068,N_8651);
nand U9542 (N_9542,N_8649,N_8420);
or U9543 (N_9543,N_8156,N_8754);
and U9544 (N_9544,N_8735,N_8247);
xor U9545 (N_9545,N_8779,N_8584);
nor U9546 (N_9546,N_8539,N_8054);
and U9547 (N_9547,N_8159,N_8112);
nand U9548 (N_9548,N_8546,N_8297);
nand U9549 (N_9549,N_8777,N_8013);
and U9550 (N_9550,N_8921,N_8719);
nand U9551 (N_9551,N_8558,N_8907);
or U9552 (N_9552,N_8381,N_8164);
xnor U9553 (N_9553,N_8891,N_8193);
xnor U9554 (N_9554,N_8449,N_8461);
and U9555 (N_9555,N_8170,N_8082);
or U9556 (N_9556,N_8033,N_8318);
and U9557 (N_9557,N_8667,N_8549);
nand U9558 (N_9558,N_8433,N_8071);
nand U9559 (N_9559,N_8687,N_8630);
nand U9560 (N_9560,N_8154,N_8646);
and U9561 (N_9561,N_8652,N_8614);
and U9562 (N_9562,N_8597,N_8573);
and U9563 (N_9563,N_8374,N_8316);
nand U9564 (N_9564,N_8827,N_8284);
or U9565 (N_9565,N_8165,N_8201);
nor U9566 (N_9566,N_8976,N_8339);
xnor U9567 (N_9567,N_8088,N_8487);
and U9568 (N_9568,N_8270,N_8400);
nand U9569 (N_9569,N_8287,N_8031);
nor U9570 (N_9570,N_8201,N_8023);
xor U9571 (N_9571,N_8078,N_8058);
nand U9572 (N_9572,N_8055,N_8592);
nand U9573 (N_9573,N_8069,N_8099);
nor U9574 (N_9574,N_8124,N_8099);
nor U9575 (N_9575,N_8945,N_8236);
nand U9576 (N_9576,N_8130,N_8928);
and U9577 (N_9577,N_8294,N_8253);
xnor U9578 (N_9578,N_8792,N_8352);
xnor U9579 (N_9579,N_8039,N_8168);
or U9580 (N_9580,N_8788,N_8559);
nand U9581 (N_9581,N_8638,N_8818);
or U9582 (N_9582,N_8117,N_8668);
or U9583 (N_9583,N_8358,N_8494);
xnor U9584 (N_9584,N_8063,N_8163);
nand U9585 (N_9585,N_8006,N_8637);
or U9586 (N_9586,N_8264,N_8808);
xnor U9587 (N_9587,N_8583,N_8730);
or U9588 (N_9588,N_8802,N_8764);
and U9589 (N_9589,N_8694,N_8158);
or U9590 (N_9590,N_8950,N_8653);
nand U9591 (N_9591,N_8896,N_8583);
nor U9592 (N_9592,N_8436,N_8535);
nor U9593 (N_9593,N_8881,N_8072);
nand U9594 (N_9594,N_8724,N_8752);
and U9595 (N_9595,N_8741,N_8006);
and U9596 (N_9596,N_8747,N_8951);
nand U9597 (N_9597,N_8382,N_8025);
nand U9598 (N_9598,N_8740,N_8105);
nor U9599 (N_9599,N_8633,N_8184);
nor U9600 (N_9600,N_8216,N_8421);
and U9601 (N_9601,N_8969,N_8218);
or U9602 (N_9602,N_8834,N_8940);
nand U9603 (N_9603,N_8749,N_8685);
and U9604 (N_9604,N_8620,N_8993);
nor U9605 (N_9605,N_8722,N_8145);
xor U9606 (N_9606,N_8486,N_8494);
nand U9607 (N_9607,N_8321,N_8703);
or U9608 (N_9608,N_8346,N_8507);
xor U9609 (N_9609,N_8013,N_8270);
nand U9610 (N_9610,N_8472,N_8345);
nor U9611 (N_9611,N_8313,N_8865);
xnor U9612 (N_9612,N_8516,N_8318);
and U9613 (N_9613,N_8732,N_8239);
and U9614 (N_9614,N_8040,N_8031);
xor U9615 (N_9615,N_8825,N_8515);
and U9616 (N_9616,N_8370,N_8621);
xor U9617 (N_9617,N_8151,N_8759);
nand U9618 (N_9618,N_8064,N_8811);
or U9619 (N_9619,N_8943,N_8400);
nand U9620 (N_9620,N_8899,N_8108);
nand U9621 (N_9621,N_8023,N_8278);
xnor U9622 (N_9622,N_8911,N_8141);
nor U9623 (N_9623,N_8507,N_8451);
xor U9624 (N_9624,N_8915,N_8288);
or U9625 (N_9625,N_8157,N_8079);
and U9626 (N_9626,N_8775,N_8983);
nand U9627 (N_9627,N_8648,N_8495);
nand U9628 (N_9628,N_8306,N_8679);
nand U9629 (N_9629,N_8095,N_8732);
xor U9630 (N_9630,N_8014,N_8933);
or U9631 (N_9631,N_8662,N_8647);
and U9632 (N_9632,N_8264,N_8605);
and U9633 (N_9633,N_8120,N_8114);
xor U9634 (N_9634,N_8541,N_8035);
nand U9635 (N_9635,N_8775,N_8350);
or U9636 (N_9636,N_8856,N_8448);
or U9637 (N_9637,N_8624,N_8310);
nor U9638 (N_9638,N_8421,N_8017);
xor U9639 (N_9639,N_8440,N_8025);
nand U9640 (N_9640,N_8434,N_8413);
xor U9641 (N_9641,N_8670,N_8147);
nand U9642 (N_9642,N_8599,N_8186);
or U9643 (N_9643,N_8889,N_8729);
and U9644 (N_9644,N_8619,N_8986);
and U9645 (N_9645,N_8547,N_8802);
or U9646 (N_9646,N_8400,N_8424);
and U9647 (N_9647,N_8988,N_8500);
and U9648 (N_9648,N_8402,N_8998);
nor U9649 (N_9649,N_8630,N_8525);
nand U9650 (N_9650,N_8664,N_8972);
and U9651 (N_9651,N_8227,N_8656);
nand U9652 (N_9652,N_8375,N_8037);
xnor U9653 (N_9653,N_8830,N_8937);
nor U9654 (N_9654,N_8652,N_8679);
and U9655 (N_9655,N_8594,N_8520);
or U9656 (N_9656,N_8573,N_8691);
nor U9657 (N_9657,N_8395,N_8813);
xnor U9658 (N_9658,N_8912,N_8558);
nand U9659 (N_9659,N_8429,N_8400);
xnor U9660 (N_9660,N_8238,N_8656);
nand U9661 (N_9661,N_8438,N_8833);
and U9662 (N_9662,N_8592,N_8487);
or U9663 (N_9663,N_8545,N_8206);
and U9664 (N_9664,N_8874,N_8325);
nand U9665 (N_9665,N_8232,N_8034);
xor U9666 (N_9666,N_8127,N_8041);
and U9667 (N_9667,N_8548,N_8691);
or U9668 (N_9668,N_8853,N_8851);
xnor U9669 (N_9669,N_8458,N_8189);
or U9670 (N_9670,N_8788,N_8104);
xnor U9671 (N_9671,N_8812,N_8823);
nor U9672 (N_9672,N_8154,N_8112);
and U9673 (N_9673,N_8989,N_8899);
nor U9674 (N_9674,N_8984,N_8288);
xor U9675 (N_9675,N_8950,N_8911);
and U9676 (N_9676,N_8845,N_8772);
nor U9677 (N_9677,N_8052,N_8674);
and U9678 (N_9678,N_8660,N_8361);
and U9679 (N_9679,N_8184,N_8216);
nand U9680 (N_9680,N_8471,N_8164);
nand U9681 (N_9681,N_8116,N_8572);
nor U9682 (N_9682,N_8080,N_8204);
nand U9683 (N_9683,N_8322,N_8259);
nand U9684 (N_9684,N_8457,N_8520);
xor U9685 (N_9685,N_8582,N_8912);
and U9686 (N_9686,N_8941,N_8220);
nand U9687 (N_9687,N_8673,N_8834);
or U9688 (N_9688,N_8658,N_8721);
nor U9689 (N_9689,N_8402,N_8583);
xor U9690 (N_9690,N_8156,N_8015);
xor U9691 (N_9691,N_8456,N_8273);
or U9692 (N_9692,N_8567,N_8004);
nor U9693 (N_9693,N_8702,N_8023);
and U9694 (N_9694,N_8546,N_8772);
xor U9695 (N_9695,N_8882,N_8786);
nor U9696 (N_9696,N_8646,N_8263);
xnor U9697 (N_9697,N_8257,N_8042);
or U9698 (N_9698,N_8780,N_8251);
xnor U9699 (N_9699,N_8194,N_8781);
xnor U9700 (N_9700,N_8196,N_8985);
and U9701 (N_9701,N_8691,N_8503);
xnor U9702 (N_9702,N_8308,N_8974);
and U9703 (N_9703,N_8359,N_8566);
nand U9704 (N_9704,N_8904,N_8761);
xnor U9705 (N_9705,N_8589,N_8897);
and U9706 (N_9706,N_8213,N_8979);
nand U9707 (N_9707,N_8743,N_8387);
xor U9708 (N_9708,N_8417,N_8960);
or U9709 (N_9709,N_8524,N_8202);
or U9710 (N_9710,N_8411,N_8622);
xor U9711 (N_9711,N_8075,N_8706);
or U9712 (N_9712,N_8158,N_8548);
nor U9713 (N_9713,N_8199,N_8368);
and U9714 (N_9714,N_8594,N_8530);
nand U9715 (N_9715,N_8268,N_8256);
nand U9716 (N_9716,N_8338,N_8528);
nand U9717 (N_9717,N_8148,N_8864);
or U9718 (N_9718,N_8655,N_8689);
and U9719 (N_9719,N_8330,N_8432);
xor U9720 (N_9720,N_8278,N_8413);
and U9721 (N_9721,N_8945,N_8264);
nand U9722 (N_9722,N_8589,N_8670);
xor U9723 (N_9723,N_8663,N_8348);
xor U9724 (N_9724,N_8061,N_8827);
or U9725 (N_9725,N_8694,N_8117);
and U9726 (N_9726,N_8215,N_8281);
or U9727 (N_9727,N_8307,N_8154);
xnor U9728 (N_9728,N_8244,N_8556);
nand U9729 (N_9729,N_8005,N_8497);
nand U9730 (N_9730,N_8809,N_8563);
and U9731 (N_9731,N_8323,N_8914);
and U9732 (N_9732,N_8699,N_8760);
nand U9733 (N_9733,N_8832,N_8517);
nand U9734 (N_9734,N_8730,N_8151);
xnor U9735 (N_9735,N_8153,N_8198);
nand U9736 (N_9736,N_8743,N_8859);
nor U9737 (N_9737,N_8528,N_8548);
xnor U9738 (N_9738,N_8068,N_8083);
nor U9739 (N_9739,N_8465,N_8870);
xor U9740 (N_9740,N_8815,N_8720);
nor U9741 (N_9741,N_8018,N_8655);
or U9742 (N_9742,N_8201,N_8740);
nor U9743 (N_9743,N_8329,N_8968);
and U9744 (N_9744,N_8049,N_8942);
and U9745 (N_9745,N_8690,N_8704);
nand U9746 (N_9746,N_8560,N_8095);
nor U9747 (N_9747,N_8348,N_8810);
and U9748 (N_9748,N_8414,N_8634);
xnor U9749 (N_9749,N_8365,N_8025);
xnor U9750 (N_9750,N_8954,N_8618);
and U9751 (N_9751,N_8627,N_8208);
xor U9752 (N_9752,N_8921,N_8372);
nor U9753 (N_9753,N_8243,N_8532);
and U9754 (N_9754,N_8480,N_8166);
nor U9755 (N_9755,N_8620,N_8531);
and U9756 (N_9756,N_8388,N_8849);
xnor U9757 (N_9757,N_8751,N_8130);
nand U9758 (N_9758,N_8634,N_8850);
nand U9759 (N_9759,N_8169,N_8020);
nand U9760 (N_9760,N_8359,N_8739);
nand U9761 (N_9761,N_8812,N_8920);
nand U9762 (N_9762,N_8387,N_8084);
or U9763 (N_9763,N_8104,N_8990);
or U9764 (N_9764,N_8070,N_8169);
nor U9765 (N_9765,N_8253,N_8711);
nand U9766 (N_9766,N_8897,N_8825);
nor U9767 (N_9767,N_8600,N_8522);
nor U9768 (N_9768,N_8401,N_8337);
xnor U9769 (N_9769,N_8503,N_8434);
or U9770 (N_9770,N_8752,N_8897);
or U9771 (N_9771,N_8277,N_8310);
xnor U9772 (N_9772,N_8707,N_8692);
or U9773 (N_9773,N_8748,N_8420);
xor U9774 (N_9774,N_8016,N_8949);
and U9775 (N_9775,N_8346,N_8915);
xnor U9776 (N_9776,N_8177,N_8621);
and U9777 (N_9777,N_8439,N_8402);
nand U9778 (N_9778,N_8460,N_8526);
nand U9779 (N_9779,N_8940,N_8240);
or U9780 (N_9780,N_8601,N_8889);
nand U9781 (N_9781,N_8623,N_8746);
nand U9782 (N_9782,N_8224,N_8704);
nand U9783 (N_9783,N_8178,N_8371);
or U9784 (N_9784,N_8608,N_8335);
nand U9785 (N_9785,N_8297,N_8458);
xor U9786 (N_9786,N_8377,N_8589);
or U9787 (N_9787,N_8313,N_8895);
nor U9788 (N_9788,N_8972,N_8668);
nand U9789 (N_9789,N_8775,N_8582);
xnor U9790 (N_9790,N_8539,N_8044);
nor U9791 (N_9791,N_8984,N_8747);
or U9792 (N_9792,N_8835,N_8647);
nand U9793 (N_9793,N_8244,N_8268);
nand U9794 (N_9794,N_8383,N_8565);
xor U9795 (N_9795,N_8958,N_8658);
nor U9796 (N_9796,N_8757,N_8931);
nor U9797 (N_9797,N_8715,N_8601);
nand U9798 (N_9798,N_8935,N_8790);
nor U9799 (N_9799,N_8419,N_8521);
and U9800 (N_9800,N_8735,N_8514);
and U9801 (N_9801,N_8111,N_8225);
or U9802 (N_9802,N_8210,N_8425);
xor U9803 (N_9803,N_8012,N_8415);
and U9804 (N_9804,N_8112,N_8360);
xor U9805 (N_9805,N_8351,N_8100);
nand U9806 (N_9806,N_8768,N_8439);
or U9807 (N_9807,N_8019,N_8641);
nand U9808 (N_9808,N_8142,N_8067);
or U9809 (N_9809,N_8105,N_8096);
nand U9810 (N_9810,N_8463,N_8849);
nand U9811 (N_9811,N_8638,N_8712);
or U9812 (N_9812,N_8889,N_8433);
or U9813 (N_9813,N_8453,N_8377);
nand U9814 (N_9814,N_8953,N_8835);
nor U9815 (N_9815,N_8848,N_8740);
or U9816 (N_9816,N_8667,N_8045);
nor U9817 (N_9817,N_8405,N_8747);
nor U9818 (N_9818,N_8701,N_8402);
or U9819 (N_9819,N_8748,N_8261);
and U9820 (N_9820,N_8692,N_8866);
nand U9821 (N_9821,N_8936,N_8201);
nor U9822 (N_9822,N_8595,N_8343);
or U9823 (N_9823,N_8238,N_8277);
nand U9824 (N_9824,N_8507,N_8526);
nor U9825 (N_9825,N_8886,N_8250);
xnor U9826 (N_9826,N_8441,N_8753);
and U9827 (N_9827,N_8467,N_8692);
xnor U9828 (N_9828,N_8586,N_8074);
nor U9829 (N_9829,N_8890,N_8343);
xnor U9830 (N_9830,N_8722,N_8175);
xnor U9831 (N_9831,N_8175,N_8349);
nor U9832 (N_9832,N_8665,N_8825);
and U9833 (N_9833,N_8237,N_8764);
or U9834 (N_9834,N_8530,N_8040);
nor U9835 (N_9835,N_8220,N_8210);
nor U9836 (N_9836,N_8096,N_8006);
nand U9837 (N_9837,N_8044,N_8465);
xnor U9838 (N_9838,N_8850,N_8264);
nand U9839 (N_9839,N_8653,N_8422);
or U9840 (N_9840,N_8738,N_8744);
nand U9841 (N_9841,N_8225,N_8186);
xnor U9842 (N_9842,N_8943,N_8470);
nor U9843 (N_9843,N_8614,N_8499);
xor U9844 (N_9844,N_8371,N_8206);
and U9845 (N_9845,N_8230,N_8277);
and U9846 (N_9846,N_8918,N_8424);
nor U9847 (N_9847,N_8221,N_8915);
xnor U9848 (N_9848,N_8738,N_8616);
nor U9849 (N_9849,N_8383,N_8367);
xnor U9850 (N_9850,N_8685,N_8986);
nor U9851 (N_9851,N_8584,N_8033);
nor U9852 (N_9852,N_8992,N_8940);
xnor U9853 (N_9853,N_8255,N_8439);
xnor U9854 (N_9854,N_8962,N_8953);
and U9855 (N_9855,N_8577,N_8406);
and U9856 (N_9856,N_8858,N_8788);
or U9857 (N_9857,N_8529,N_8671);
xnor U9858 (N_9858,N_8963,N_8446);
or U9859 (N_9859,N_8814,N_8178);
nand U9860 (N_9860,N_8300,N_8466);
nor U9861 (N_9861,N_8286,N_8198);
and U9862 (N_9862,N_8092,N_8378);
or U9863 (N_9863,N_8982,N_8836);
nor U9864 (N_9864,N_8312,N_8785);
and U9865 (N_9865,N_8056,N_8069);
nor U9866 (N_9866,N_8806,N_8594);
xor U9867 (N_9867,N_8562,N_8196);
nor U9868 (N_9868,N_8418,N_8843);
nand U9869 (N_9869,N_8695,N_8968);
nand U9870 (N_9870,N_8344,N_8456);
nand U9871 (N_9871,N_8395,N_8111);
nand U9872 (N_9872,N_8801,N_8836);
xnor U9873 (N_9873,N_8577,N_8427);
xor U9874 (N_9874,N_8713,N_8404);
nand U9875 (N_9875,N_8272,N_8763);
or U9876 (N_9876,N_8970,N_8224);
and U9877 (N_9877,N_8448,N_8323);
or U9878 (N_9878,N_8233,N_8890);
xnor U9879 (N_9879,N_8513,N_8854);
and U9880 (N_9880,N_8825,N_8470);
nor U9881 (N_9881,N_8073,N_8174);
xor U9882 (N_9882,N_8854,N_8160);
or U9883 (N_9883,N_8429,N_8697);
or U9884 (N_9884,N_8898,N_8084);
and U9885 (N_9885,N_8620,N_8909);
and U9886 (N_9886,N_8379,N_8776);
nand U9887 (N_9887,N_8297,N_8690);
nor U9888 (N_9888,N_8143,N_8595);
nand U9889 (N_9889,N_8719,N_8824);
nand U9890 (N_9890,N_8393,N_8002);
nand U9891 (N_9891,N_8432,N_8395);
and U9892 (N_9892,N_8985,N_8244);
nor U9893 (N_9893,N_8692,N_8185);
nor U9894 (N_9894,N_8679,N_8138);
nand U9895 (N_9895,N_8503,N_8402);
xor U9896 (N_9896,N_8757,N_8285);
nand U9897 (N_9897,N_8022,N_8441);
nand U9898 (N_9898,N_8063,N_8284);
nor U9899 (N_9899,N_8585,N_8293);
and U9900 (N_9900,N_8195,N_8856);
or U9901 (N_9901,N_8513,N_8350);
nand U9902 (N_9902,N_8358,N_8253);
nand U9903 (N_9903,N_8069,N_8184);
or U9904 (N_9904,N_8955,N_8905);
nand U9905 (N_9905,N_8464,N_8753);
xor U9906 (N_9906,N_8134,N_8834);
nor U9907 (N_9907,N_8224,N_8275);
nand U9908 (N_9908,N_8465,N_8457);
or U9909 (N_9909,N_8436,N_8904);
nand U9910 (N_9910,N_8779,N_8523);
or U9911 (N_9911,N_8267,N_8412);
nor U9912 (N_9912,N_8648,N_8372);
xnor U9913 (N_9913,N_8378,N_8030);
xnor U9914 (N_9914,N_8620,N_8106);
xnor U9915 (N_9915,N_8610,N_8194);
and U9916 (N_9916,N_8400,N_8865);
xor U9917 (N_9917,N_8877,N_8499);
xnor U9918 (N_9918,N_8778,N_8627);
nand U9919 (N_9919,N_8833,N_8132);
or U9920 (N_9920,N_8805,N_8082);
nor U9921 (N_9921,N_8227,N_8152);
and U9922 (N_9922,N_8966,N_8309);
nor U9923 (N_9923,N_8160,N_8191);
or U9924 (N_9924,N_8069,N_8140);
nand U9925 (N_9925,N_8560,N_8690);
nand U9926 (N_9926,N_8770,N_8824);
nand U9927 (N_9927,N_8834,N_8197);
or U9928 (N_9928,N_8082,N_8366);
or U9929 (N_9929,N_8903,N_8238);
nand U9930 (N_9930,N_8197,N_8645);
or U9931 (N_9931,N_8049,N_8539);
or U9932 (N_9932,N_8136,N_8763);
or U9933 (N_9933,N_8497,N_8467);
and U9934 (N_9934,N_8731,N_8018);
nor U9935 (N_9935,N_8987,N_8012);
nor U9936 (N_9936,N_8578,N_8072);
nor U9937 (N_9937,N_8330,N_8181);
and U9938 (N_9938,N_8315,N_8318);
nor U9939 (N_9939,N_8851,N_8816);
xnor U9940 (N_9940,N_8248,N_8435);
nor U9941 (N_9941,N_8415,N_8798);
xnor U9942 (N_9942,N_8414,N_8778);
or U9943 (N_9943,N_8037,N_8052);
nand U9944 (N_9944,N_8798,N_8331);
and U9945 (N_9945,N_8289,N_8385);
and U9946 (N_9946,N_8285,N_8876);
nand U9947 (N_9947,N_8458,N_8649);
xor U9948 (N_9948,N_8782,N_8402);
nand U9949 (N_9949,N_8809,N_8774);
xnor U9950 (N_9950,N_8668,N_8680);
nor U9951 (N_9951,N_8467,N_8075);
nand U9952 (N_9952,N_8788,N_8218);
nand U9953 (N_9953,N_8593,N_8592);
xnor U9954 (N_9954,N_8087,N_8352);
or U9955 (N_9955,N_8280,N_8619);
nand U9956 (N_9956,N_8176,N_8126);
nor U9957 (N_9957,N_8061,N_8629);
or U9958 (N_9958,N_8898,N_8255);
nand U9959 (N_9959,N_8930,N_8182);
xor U9960 (N_9960,N_8134,N_8568);
xor U9961 (N_9961,N_8241,N_8699);
xor U9962 (N_9962,N_8649,N_8622);
or U9963 (N_9963,N_8173,N_8327);
xnor U9964 (N_9964,N_8472,N_8962);
nand U9965 (N_9965,N_8015,N_8458);
and U9966 (N_9966,N_8271,N_8889);
nand U9967 (N_9967,N_8361,N_8978);
nand U9968 (N_9968,N_8711,N_8328);
and U9969 (N_9969,N_8448,N_8544);
or U9970 (N_9970,N_8746,N_8665);
nor U9971 (N_9971,N_8895,N_8120);
nor U9972 (N_9972,N_8787,N_8080);
and U9973 (N_9973,N_8011,N_8675);
nor U9974 (N_9974,N_8162,N_8782);
and U9975 (N_9975,N_8603,N_8713);
and U9976 (N_9976,N_8209,N_8761);
and U9977 (N_9977,N_8603,N_8222);
xor U9978 (N_9978,N_8741,N_8656);
nand U9979 (N_9979,N_8461,N_8333);
xnor U9980 (N_9980,N_8849,N_8049);
and U9981 (N_9981,N_8328,N_8257);
nand U9982 (N_9982,N_8508,N_8610);
xnor U9983 (N_9983,N_8282,N_8435);
nand U9984 (N_9984,N_8735,N_8475);
or U9985 (N_9985,N_8037,N_8796);
and U9986 (N_9986,N_8192,N_8277);
xnor U9987 (N_9987,N_8488,N_8348);
xor U9988 (N_9988,N_8076,N_8276);
xnor U9989 (N_9989,N_8430,N_8330);
nor U9990 (N_9990,N_8977,N_8890);
nor U9991 (N_9991,N_8711,N_8620);
nand U9992 (N_9992,N_8268,N_8299);
and U9993 (N_9993,N_8005,N_8858);
and U9994 (N_9994,N_8106,N_8867);
nor U9995 (N_9995,N_8626,N_8150);
nor U9996 (N_9996,N_8402,N_8106);
nand U9997 (N_9997,N_8310,N_8223);
or U9998 (N_9998,N_8486,N_8615);
and U9999 (N_9999,N_8662,N_8351);
xor U10000 (N_10000,N_9793,N_9927);
xnor U10001 (N_10001,N_9578,N_9689);
or U10002 (N_10002,N_9328,N_9008);
nor U10003 (N_10003,N_9105,N_9033);
nor U10004 (N_10004,N_9762,N_9907);
or U10005 (N_10005,N_9076,N_9056);
nand U10006 (N_10006,N_9016,N_9479);
and U10007 (N_10007,N_9298,N_9232);
or U10008 (N_10008,N_9525,N_9398);
or U10009 (N_10009,N_9204,N_9724);
xnor U10010 (N_10010,N_9528,N_9219);
nand U10011 (N_10011,N_9338,N_9668);
xnor U10012 (N_10012,N_9455,N_9249);
and U10013 (N_10013,N_9471,N_9753);
nor U10014 (N_10014,N_9655,N_9878);
xnor U10015 (N_10015,N_9199,N_9406);
xor U10016 (N_10016,N_9480,N_9586);
nand U10017 (N_10017,N_9997,N_9703);
nand U10018 (N_10018,N_9962,N_9353);
xor U10019 (N_10019,N_9392,N_9553);
xor U10020 (N_10020,N_9032,N_9855);
nand U10021 (N_10021,N_9048,N_9501);
or U10022 (N_10022,N_9014,N_9215);
nand U10023 (N_10023,N_9568,N_9978);
xnor U10024 (N_10024,N_9991,N_9229);
nand U10025 (N_10025,N_9102,N_9601);
xnor U10026 (N_10026,N_9859,N_9325);
nor U10027 (N_10027,N_9567,N_9630);
and U10028 (N_10028,N_9660,N_9323);
nor U10029 (N_10029,N_9582,N_9696);
and U10030 (N_10030,N_9576,N_9504);
or U10031 (N_10031,N_9900,N_9626);
nand U10032 (N_10032,N_9852,N_9468);
nand U10033 (N_10033,N_9449,N_9632);
xnor U10034 (N_10034,N_9972,N_9517);
xnor U10035 (N_10035,N_9333,N_9983);
nand U10036 (N_10036,N_9691,N_9025);
xor U10037 (N_10037,N_9915,N_9269);
nor U10038 (N_10038,N_9585,N_9144);
xor U10039 (N_10039,N_9417,N_9286);
or U10040 (N_10040,N_9295,N_9395);
and U10041 (N_10041,N_9268,N_9506);
nand U10042 (N_10042,N_9542,N_9709);
or U10043 (N_10043,N_9075,N_9986);
and U10044 (N_10044,N_9861,N_9796);
nand U10045 (N_10045,N_9231,N_9133);
xor U10046 (N_10046,N_9721,N_9513);
nor U10047 (N_10047,N_9264,N_9957);
or U10048 (N_10048,N_9875,N_9397);
nand U10049 (N_10049,N_9018,N_9457);
xnor U10050 (N_10050,N_9136,N_9499);
nand U10051 (N_10051,N_9013,N_9639);
nand U10052 (N_10052,N_9519,N_9967);
xor U10053 (N_10053,N_9924,N_9839);
nand U10054 (N_10054,N_9718,N_9532);
and U10055 (N_10055,N_9277,N_9055);
nor U10056 (N_10056,N_9556,N_9867);
or U10057 (N_10057,N_9917,N_9384);
and U10058 (N_10058,N_9717,N_9943);
and U10059 (N_10059,N_9066,N_9091);
nor U10060 (N_10060,N_9431,N_9699);
or U10061 (N_10061,N_9386,N_9176);
or U10062 (N_10062,N_9217,N_9625);
xor U10063 (N_10063,N_9308,N_9040);
and U10064 (N_10064,N_9090,N_9147);
and U10065 (N_10065,N_9970,N_9421);
xor U10066 (N_10066,N_9562,N_9493);
and U10067 (N_10067,N_9291,N_9099);
or U10068 (N_10068,N_9732,N_9862);
nor U10069 (N_10069,N_9330,N_9830);
and U10070 (N_10070,N_9694,N_9111);
nor U10071 (N_10071,N_9110,N_9530);
and U10072 (N_10072,N_9445,N_9824);
nor U10073 (N_10073,N_9038,N_9987);
nor U10074 (N_10074,N_9448,N_9754);
or U10075 (N_10075,N_9423,N_9591);
and U10076 (N_10076,N_9171,N_9916);
and U10077 (N_10077,N_9010,N_9363);
and U10078 (N_10078,N_9408,N_9122);
or U10079 (N_10079,N_9460,N_9758);
and U10080 (N_10080,N_9311,N_9736);
nand U10081 (N_10081,N_9258,N_9175);
nand U10082 (N_10082,N_9009,N_9463);
nor U10083 (N_10083,N_9939,N_9496);
xor U10084 (N_10084,N_9690,N_9677);
nor U10085 (N_10085,N_9918,N_9054);
nand U10086 (N_10086,N_9058,N_9404);
and U10087 (N_10087,N_9287,N_9557);
nor U10088 (N_10088,N_9139,N_9913);
and U10089 (N_10089,N_9934,N_9383);
or U10090 (N_10090,N_9096,N_9597);
and U10091 (N_10091,N_9821,N_9263);
nand U10092 (N_10092,N_9604,N_9451);
nor U10093 (N_10093,N_9687,N_9920);
nor U10094 (N_10094,N_9117,N_9946);
or U10095 (N_10095,N_9738,N_9419);
nor U10096 (N_10096,N_9940,N_9174);
or U10097 (N_10097,N_9304,N_9609);
and U10098 (N_10098,N_9168,N_9202);
or U10099 (N_10099,N_9926,N_9870);
xnor U10100 (N_10100,N_9743,N_9605);
nand U10101 (N_10101,N_9886,N_9871);
xor U10102 (N_10102,N_9512,N_9848);
xor U10103 (N_10103,N_9728,N_9294);
or U10104 (N_10104,N_9279,N_9800);
xor U10105 (N_10105,N_9617,N_9619);
xor U10106 (N_10106,N_9465,N_9869);
nor U10107 (N_10107,N_9389,N_9780);
nor U10108 (N_10108,N_9108,N_9831);
or U10109 (N_10109,N_9890,N_9078);
or U10110 (N_10110,N_9046,N_9931);
nor U10111 (N_10111,N_9554,N_9845);
and U10112 (N_10112,N_9674,N_9317);
nor U10113 (N_10113,N_9146,N_9923);
nor U10114 (N_10114,N_9012,N_9563);
and U10115 (N_10115,N_9245,N_9148);
nand U10116 (N_10116,N_9782,N_9836);
nor U10117 (N_10117,N_9274,N_9372);
nand U10118 (N_10118,N_9807,N_9067);
xnor U10119 (N_10119,N_9297,N_9739);
xor U10120 (N_10120,N_9726,N_9080);
nor U10121 (N_10121,N_9187,N_9273);
and U10122 (N_10122,N_9705,N_9347);
nor U10123 (N_10123,N_9158,N_9949);
or U10124 (N_10124,N_9220,N_9252);
or U10125 (N_10125,N_9050,N_9153);
nor U10126 (N_10126,N_9536,N_9675);
xor U10127 (N_10127,N_9921,N_9053);
and U10128 (N_10128,N_9321,N_9894);
nand U10129 (N_10129,N_9095,N_9785);
or U10130 (N_10130,N_9896,N_9107);
and U10131 (N_10131,N_9768,N_9786);
nor U10132 (N_10132,N_9827,N_9082);
xnor U10133 (N_10133,N_9874,N_9779);
nor U10134 (N_10134,N_9706,N_9692);
xnor U10135 (N_10135,N_9285,N_9879);
nand U10136 (N_10136,N_9611,N_9093);
xor U10137 (N_10137,N_9310,N_9633);
nor U10138 (N_10138,N_9209,N_9276);
xor U10139 (N_10139,N_9747,N_9369);
and U10140 (N_10140,N_9128,N_9381);
nor U10141 (N_10141,N_9531,N_9529);
nor U10142 (N_10142,N_9198,N_9239);
or U10143 (N_10143,N_9378,N_9461);
and U10144 (N_10144,N_9180,N_9631);
nor U10145 (N_10145,N_9284,N_9283);
nor U10146 (N_10146,N_9343,N_9505);
nor U10147 (N_10147,N_9545,N_9261);
or U10148 (N_10148,N_9935,N_9334);
or U10149 (N_10149,N_9620,N_9841);
nand U10150 (N_10150,N_9169,N_9248);
xor U10151 (N_10151,N_9805,N_9769);
or U10152 (N_10152,N_9079,N_9322);
and U10153 (N_10153,N_9956,N_9643);
nor U10154 (N_10154,N_9897,N_9524);
nor U10155 (N_10155,N_9974,N_9751);
xnor U10156 (N_10156,N_9316,N_9233);
xor U10157 (N_10157,N_9351,N_9784);
xor U10158 (N_10158,N_9045,N_9968);
nor U10159 (N_10159,N_9925,N_9003);
and U10160 (N_10160,N_9037,N_9083);
nand U10161 (N_10161,N_9550,N_9394);
and U10162 (N_10162,N_9436,N_9179);
xnor U10163 (N_10163,N_9906,N_9314);
and U10164 (N_10164,N_9100,N_9701);
or U10165 (N_10165,N_9636,N_9755);
nor U10166 (N_10166,N_9382,N_9627);
xnor U10167 (N_10167,N_9339,N_9256);
or U10168 (N_10168,N_9422,N_9434);
nand U10169 (N_10169,N_9326,N_9470);
nand U10170 (N_10170,N_9977,N_9905);
or U10171 (N_10171,N_9558,N_9760);
xnor U10172 (N_10172,N_9663,N_9300);
and U10173 (N_10173,N_9534,N_9729);
and U10174 (N_10174,N_9646,N_9988);
nor U10175 (N_10175,N_9002,N_9484);
or U10176 (N_10176,N_9137,N_9188);
nor U10177 (N_10177,N_9789,N_9998);
nor U10178 (N_10178,N_9361,N_9764);
nand U10179 (N_10179,N_9464,N_9355);
nor U10180 (N_10180,N_9425,N_9380);
nor U10181 (N_10181,N_9892,N_9370);
and U10182 (N_10182,N_9610,N_9603);
or U10183 (N_10183,N_9613,N_9833);
nor U10184 (N_10184,N_9126,N_9723);
xnor U10185 (N_10185,N_9811,N_9642);
xor U10186 (N_10186,N_9345,N_9645);
nand U10187 (N_10187,N_9662,N_9376);
xnor U10188 (N_10188,N_9930,N_9600);
nor U10189 (N_10189,N_9490,N_9569);
or U10190 (N_10190,N_9227,N_9544);
xor U10191 (N_10191,N_9428,N_9893);
or U10192 (N_10192,N_9961,N_9882);
xnor U10193 (N_10193,N_9963,N_9608);
nor U10194 (N_10194,N_9362,N_9001);
nand U10195 (N_10195,N_9292,N_9246);
or U10196 (N_10196,N_9981,N_9863);
nor U10197 (N_10197,N_9192,N_9942);
and U10198 (N_10198,N_9062,N_9026);
and U10199 (N_10199,N_9856,N_9659);
and U10200 (N_10200,N_9522,N_9710);
and U10201 (N_10201,N_9735,N_9685);
nand U10202 (N_10202,N_9938,N_9145);
nand U10203 (N_10203,N_9748,N_9681);
or U10204 (N_10204,N_9481,N_9621);
and U10205 (N_10205,N_9123,N_9388);
or U10206 (N_10206,N_9570,N_9864);
nand U10207 (N_10207,N_9750,N_9731);
or U10208 (N_10208,N_9899,N_9801);
and U10209 (N_10209,N_9377,N_9432);
xnor U10210 (N_10210,N_9167,N_9443);
xnor U10211 (N_10211,N_9761,N_9098);
and U10212 (N_10212,N_9344,N_9656);
and U10213 (N_10213,N_9476,N_9876);
or U10214 (N_10214,N_9358,N_9103);
nor U10215 (N_10215,N_9527,N_9958);
or U10216 (N_10216,N_9004,N_9795);
and U10217 (N_10217,N_9329,N_9759);
xnor U10218 (N_10218,N_9073,N_9520);
nor U10219 (N_10219,N_9085,N_9120);
nand U10220 (N_10220,N_9475,N_9510);
nand U10221 (N_10221,N_9777,N_9737);
xnor U10222 (N_10222,N_9488,N_9820);
xnor U10223 (N_10223,N_9757,N_9944);
xnor U10224 (N_10224,N_9223,N_9666);
or U10225 (N_10225,N_9473,N_9135);
and U10226 (N_10226,N_9230,N_9022);
or U10227 (N_10227,N_9390,N_9965);
nor U10228 (N_10228,N_9088,N_9995);
nor U10229 (N_10229,N_9034,N_9684);
and U10230 (N_10230,N_9799,N_9400);
nand U10231 (N_10231,N_9023,N_9672);
and U10232 (N_10232,N_9057,N_9819);
nor U10233 (N_10233,N_9368,N_9036);
xnor U10234 (N_10234,N_9812,N_9669);
nor U10235 (N_10235,N_9776,N_9772);
xor U10236 (N_10236,N_9224,N_9584);
nor U10237 (N_10237,N_9638,N_9301);
nor U10238 (N_10238,N_9156,N_9828);
xnor U10239 (N_10239,N_9028,N_9679);
xnor U10240 (N_10240,N_9980,N_9733);
and U10241 (N_10241,N_9700,N_9265);
nor U10242 (N_10242,N_9106,N_9447);
or U10243 (N_10243,N_9590,N_9410);
nand U10244 (N_10244,N_9719,N_9551);
nand U10245 (N_10245,N_9722,N_9213);
and U10246 (N_10246,N_9832,N_9409);
and U10247 (N_10247,N_9971,N_9740);
or U10248 (N_10248,N_9933,N_9132);
or U10249 (N_10249,N_9212,N_9420);
xor U10250 (N_10250,N_9500,N_9730);
or U10251 (N_10251,N_9727,N_9515);
or U10252 (N_10252,N_9251,N_9216);
and U10253 (N_10253,N_9911,N_9664);
nor U10254 (N_10254,N_9714,N_9068);
nand U10255 (N_10255,N_9708,N_9296);
nand U10256 (N_10256,N_9453,N_9454);
and U10257 (N_10257,N_9596,N_9086);
and U10258 (N_10258,N_9975,N_9313);
nor U10259 (N_10259,N_9868,N_9161);
nor U10260 (N_10260,N_9673,N_9838);
or U10261 (N_10261,N_9650,N_9887);
and U10262 (N_10262,N_9952,N_9507);
and U10263 (N_10263,N_9902,N_9257);
nor U10264 (N_10264,N_9290,N_9131);
and U10265 (N_10265,N_9797,N_9541);
nor U10266 (N_10266,N_9798,N_9170);
nor U10267 (N_10267,N_9307,N_9725);
xor U10268 (N_10268,N_9910,N_9825);
nor U10269 (N_10269,N_9020,N_9680);
and U10270 (N_10270,N_9477,N_9280);
xnor U10271 (N_10271,N_9883,N_9052);
xor U10272 (N_10272,N_9282,N_9514);
nor U10273 (N_10273,N_9474,N_9024);
and U10274 (N_10274,N_9686,N_9482);
nor U10275 (N_10275,N_9393,N_9564);
xor U10276 (N_10276,N_9077,N_9275);
or U10277 (N_10277,N_9342,N_9140);
and U10278 (N_10278,N_9462,N_9486);
nor U10279 (N_10279,N_9458,N_9561);
nand U10280 (N_10280,N_9787,N_9337);
and U10281 (N_10281,N_9155,N_9509);
xor U10282 (N_10282,N_9379,N_9624);
nand U10283 (N_10283,N_9396,N_9191);
xnor U10284 (N_10284,N_9456,N_9485);
and U10285 (N_10285,N_9640,N_9190);
or U10286 (N_10286,N_9982,N_9305);
and U10287 (N_10287,N_9773,N_9616);
and U10288 (N_10288,N_9403,N_9109);
xor U10289 (N_10289,N_9994,N_9047);
nor U10290 (N_10290,N_9592,N_9255);
nor U10291 (N_10291,N_9788,N_9872);
or U10292 (N_10292,N_9629,N_9823);
and U10293 (N_10293,N_9165,N_9654);
or U10294 (N_10294,N_9895,N_9637);
nand U10295 (N_10295,N_9041,N_9649);
nand U10296 (N_10296,N_9498,N_9884);
and U10297 (N_10297,N_9070,N_9152);
xor U10298 (N_10298,N_9060,N_9164);
and U10299 (N_10299,N_9712,N_9985);
and U10300 (N_10300,N_9332,N_9612);
nand U10301 (N_10301,N_9092,N_9118);
xnor U10302 (N_10302,N_9319,N_9818);
or U10303 (N_10303,N_9698,N_9635);
nor U10304 (N_10304,N_9955,N_9702);
or U10305 (N_10305,N_9221,N_9929);
nand U10306 (N_10306,N_9440,N_9424);
nand U10307 (N_10307,N_9163,N_9356);
xnor U10308 (N_10308,N_9559,N_9149);
xnor U10309 (N_10309,N_9017,N_9483);
nor U10310 (N_10310,N_9201,N_9948);
nand U10311 (N_10311,N_9150,N_9006);
nand U10312 (N_10312,N_9452,N_9250);
or U10313 (N_10313,N_9492,N_9115);
and U10314 (N_10314,N_9973,N_9318);
or U10315 (N_10315,N_9157,N_9734);
xor U10316 (N_10316,N_9803,N_9683);
nand U10317 (N_10317,N_9976,N_9826);
or U10318 (N_10318,N_9951,N_9954);
nor U10319 (N_10319,N_9543,N_9303);
xnor U10320 (N_10320,N_9502,N_9267);
or U10321 (N_10321,N_9346,N_9244);
nor U10322 (N_10322,N_9427,N_9181);
and U10323 (N_10323,N_9763,N_9840);
xnor U10324 (N_10324,N_9535,N_9270);
or U10325 (N_10325,N_9540,N_9450);
nand U10326 (N_10326,N_9143,N_9309);
or U10327 (N_10327,N_9352,N_9713);
and U10328 (N_10328,N_9580,N_9237);
and U10329 (N_10329,N_9950,N_9278);
nor U10330 (N_10330,N_9589,N_9439);
xor U10331 (N_10331,N_9588,N_9587);
nand U10332 (N_10332,N_9097,N_9446);
nor U10333 (N_10333,N_9555,N_9411);
xor U10334 (N_10334,N_9072,N_9908);
and U10335 (N_10335,N_9089,N_9953);
nor U10336 (N_10336,N_9288,N_9430);
and U10337 (N_10337,N_9682,N_9720);
nor U10338 (N_10338,N_9716,N_9129);
xnor U10339 (N_10339,N_9348,N_9546);
and U10340 (N_10340,N_9043,N_9770);
nor U10341 (N_10341,N_9593,N_9922);
nor U10342 (N_10342,N_9829,N_9566);
and U10343 (N_10343,N_9774,N_9375);
nand U10344 (N_10344,N_9491,N_9005);
xor U10345 (N_10345,N_9966,N_9945);
nand U10346 (N_10346,N_9560,N_9628);
nand U10347 (N_10347,N_9266,N_9183);
nor U10348 (N_10348,N_9865,N_9087);
nor U10349 (N_10349,N_9113,N_9808);
or U10350 (N_10350,N_9813,N_9315);
nor U10351 (N_10351,N_9299,N_9121);
nor U10352 (N_10352,N_9162,N_9860);
and U10353 (N_10353,N_9151,N_9741);
and U10354 (N_10354,N_9011,N_9577);
nor U10355 (N_10355,N_9416,N_9615);
or U10356 (N_10356,N_9472,N_9039);
xnor U10357 (N_10357,N_9693,N_9327);
and U10358 (N_10358,N_9990,N_9240);
and U10359 (N_10359,N_9027,N_9651);
xor U10360 (N_10360,N_9196,N_9324);
and U10361 (N_10361,N_9206,N_9804);
xor U10362 (N_10362,N_9790,N_9467);
and U10363 (N_10363,N_9766,N_9853);
xnor U10364 (N_10364,N_9749,N_9644);
nor U10365 (N_10365,N_9418,N_9007);
and U10366 (N_10366,N_9594,N_9602);
or U10367 (N_10367,N_9842,N_9194);
or U10368 (N_10368,N_9360,N_9247);
and U10369 (N_10369,N_9433,N_9814);
or U10370 (N_10370,N_9238,N_9579);
or U10371 (N_10371,N_9573,N_9441);
nor U10372 (N_10372,N_9197,N_9996);
nand U10373 (N_10373,N_9866,N_9401);
xnor U10374 (N_10374,N_9837,N_9225);
nand U10375 (N_10375,N_9847,N_9494);
xor U10376 (N_10376,N_9021,N_9834);
and U10377 (N_10377,N_9349,N_9665);
nor U10378 (N_10378,N_9200,N_9172);
nand U10379 (N_10379,N_9426,N_9262);
and U10380 (N_10380,N_9516,N_9399);
xnor U10381 (N_10381,N_9160,N_9341);
and U10382 (N_10382,N_9336,N_9335);
nor U10383 (N_10383,N_9574,N_9858);
nor U10384 (N_10384,N_9112,N_9081);
nand U10385 (N_10385,N_9539,N_9189);
nor U10386 (N_10386,N_9909,N_9815);
and U10387 (N_10387,N_9667,N_9029);
xor U10388 (N_10388,N_9989,N_9312);
nor U10389 (N_10389,N_9391,N_9993);
nor U10390 (N_10390,N_9688,N_9402);
nand U10391 (N_10391,N_9159,N_9648);
or U10392 (N_10392,N_9794,N_9742);
nand U10393 (N_10393,N_9241,N_9849);
or U10394 (N_10394,N_9671,N_9177);
nand U10395 (N_10395,N_9901,N_9444);
nor U10396 (N_10396,N_9538,N_9243);
nand U10397 (N_10397,N_9548,N_9289);
and U10398 (N_10398,N_9822,N_9138);
or U10399 (N_10399,N_9094,N_9063);
or U10400 (N_10400,N_9130,N_9571);
nand U10401 (N_10401,N_9850,N_9186);
xor U10402 (N_10402,N_9806,N_9653);
nor U10403 (N_10403,N_9623,N_9331);
nor U10404 (N_10404,N_9969,N_9914);
and U10405 (N_10405,N_9413,N_9599);
nand U10406 (N_10406,N_9715,N_9792);
nand U10407 (N_10407,N_9781,N_9125);
or U10408 (N_10408,N_9373,N_9676);
nand U10409 (N_10409,N_9697,N_9959);
xnor U10410 (N_10410,N_9178,N_9412);
or U10411 (N_10411,N_9365,N_9134);
or U10412 (N_10412,N_9984,N_9208);
and U10413 (N_10413,N_9835,N_9964);
nor U10414 (N_10414,N_9891,N_9218);
nand U10415 (N_10415,N_9614,N_9104);
xor U10416 (N_10416,N_9260,N_9817);
or U10417 (N_10417,N_9873,N_9521);
xnor U10418 (N_10418,N_9254,N_9116);
xnor U10419 (N_10419,N_9783,N_9704);
and U10420 (N_10420,N_9359,N_9438);
and U10421 (N_10421,N_9802,N_9881);
xor U10422 (N_10422,N_9071,N_9992);
and U10423 (N_10423,N_9366,N_9302);
nand U10424 (N_10424,N_9607,N_9320);
and U10425 (N_10425,N_9854,N_9889);
nand U10426 (N_10426,N_9166,N_9809);
and U10427 (N_10427,N_9019,N_9407);
nor U10428 (N_10428,N_9572,N_9101);
and U10429 (N_10429,N_9124,N_9778);
xnor U10430 (N_10430,N_9466,N_9707);
xor U10431 (N_10431,N_9414,N_9919);
xor U10432 (N_10432,N_9767,N_9000);
xor U10433 (N_10433,N_9618,N_9652);
or U10434 (N_10434,N_9880,N_9661);
xnor U10435 (N_10435,N_9552,N_9435);
and U10436 (N_10436,N_9888,N_9184);
nand U10437 (N_10437,N_9069,N_9015);
nor U10438 (N_10438,N_9928,N_9084);
nand U10439 (N_10439,N_9647,N_9581);
nor U10440 (N_10440,N_9222,N_9903);
xnor U10441 (N_10441,N_9234,N_9657);
and U10442 (N_10442,N_9658,N_9371);
xnor U10443 (N_10443,N_9415,N_9745);
and U10444 (N_10444,N_9207,N_9670);
or U10445 (N_10445,N_9752,N_9364);
nor U10446 (N_10446,N_9547,N_9306);
or U10447 (N_10447,N_9526,N_9442);
and U10448 (N_10448,N_9044,N_9523);
nand U10449 (N_10449,N_9960,N_9979);
nor U10450 (N_10450,N_9203,N_9583);
and U10451 (N_10451,N_9746,N_9059);
or U10452 (N_10452,N_9695,N_9641);
nand U10453 (N_10453,N_9374,N_9182);
nand U10454 (N_10454,N_9511,N_9429);
xor U10455 (N_10455,N_9357,N_9478);
nand U10456 (N_10456,N_9904,N_9193);
and U10457 (N_10457,N_9503,N_9127);
xor U10458 (N_10458,N_9771,N_9898);
or U10459 (N_10459,N_9253,N_9765);
nor U10460 (N_10460,N_9775,N_9912);
nor U10461 (N_10461,N_9756,N_9851);
and U10462 (N_10462,N_9235,N_9051);
nor U10463 (N_10463,N_9214,N_9367);
nor U10464 (N_10464,N_9487,N_9350);
and U10465 (N_10465,N_9210,N_9340);
nand U10466 (N_10466,N_9226,N_9937);
xnor U10467 (N_10467,N_9064,N_9537);
or U10468 (N_10468,N_9272,N_9065);
nand U10469 (N_10469,N_9387,N_9049);
xnor U10470 (N_10470,N_9857,N_9242);
nand U10471 (N_10471,N_9114,N_9154);
nor U10472 (N_10472,N_9495,N_9293);
nand U10473 (N_10473,N_9622,N_9606);
or U10474 (N_10474,N_9549,N_9843);
or U10475 (N_10475,N_9459,N_9354);
or U10476 (N_10476,N_9405,N_9119);
nand U10477 (N_10477,N_9195,N_9565);
nor U10478 (N_10478,N_9598,N_9385);
xnor U10479 (N_10479,N_9185,N_9061);
nor U10480 (N_10480,N_9595,N_9281);
nand U10481 (N_10481,N_9844,N_9205);
and U10482 (N_10482,N_9885,N_9437);
nand U10483 (N_10483,N_9035,N_9259);
nor U10484 (N_10484,N_9031,N_9877);
and U10485 (N_10485,N_9271,N_9678);
nor U10486 (N_10486,N_9489,N_9947);
nor U10487 (N_10487,N_9936,N_9236);
and U10488 (N_10488,N_9634,N_9142);
or U10489 (N_10489,N_9932,N_9211);
xnor U10490 (N_10490,N_9469,N_9711);
nand U10491 (N_10491,N_9518,N_9173);
or U10492 (N_10492,N_9074,N_9497);
nand U10493 (N_10493,N_9575,N_9030);
xor U10494 (N_10494,N_9999,N_9810);
xnor U10495 (N_10495,N_9941,N_9816);
nand U10496 (N_10496,N_9744,N_9228);
xnor U10497 (N_10497,N_9141,N_9846);
nand U10498 (N_10498,N_9533,N_9042);
nor U10499 (N_10499,N_9508,N_9791);
nor U10500 (N_10500,N_9261,N_9942);
nand U10501 (N_10501,N_9387,N_9345);
nor U10502 (N_10502,N_9580,N_9412);
and U10503 (N_10503,N_9430,N_9462);
nand U10504 (N_10504,N_9389,N_9820);
xor U10505 (N_10505,N_9011,N_9926);
or U10506 (N_10506,N_9777,N_9906);
nand U10507 (N_10507,N_9175,N_9620);
nor U10508 (N_10508,N_9942,N_9960);
and U10509 (N_10509,N_9834,N_9669);
xor U10510 (N_10510,N_9962,N_9186);
nand U10511 (N_10511,N_9774,N_9541);
or U10512 (N_10512,N_9170,N_9456);
and U10513 (N_10513,N_9605,N_9575);
nand U10514 (N_10514,N_9416,N_9934);
and U10515 (N_10515,N_9179,N_9312);
or U10516 (N_10516,N_9581,N_9339);
nand U10517 (N_10517,N_9633,N_9420);
or U10518 (N_10518,N_9834,N_9775);
xnor U10519 (N_10519,N_9700,N_9711);
nand U10520 (N_10520,N_9057,N_9444);
nor U10521 (N_10521,N_9065,N_9823);
nand U10522 (N_10522,N_9361,N_9834);
or U10523 (N_10523,N_9092,N_9212);
or U10524 (N_10524,N_9672,N_9254);
xnor U10525 (N_10525,N_9238,N_9267);
or U10526 (N_10526,N_9663,N_9029);
nand U10527 (N_10527,N_9808,N_9948);
xnor U10528 (N_10528,N_9761,N_9039);
or U10529 (N_10529,N_9838,N_9338);
and U10530 (N_10530,N_9529,N_9179);
or U10531 (N_10531,N_9250,N_9341);
xor U10532 (N_10532,N_9871,N_9219);
nand U10533 (N_10533,N_9585,N_9171);
nor U10534 (N_10534,N_9438,N_9988);
nand U10535 (N_10535,N_9720,N_9358);
nor U10536 (N_10536,N_9576,N_9819);
or U10537 (N_10537,N_9423,N_9334);
nand U10538 (N_10538,N_9708,N_9170);
nor U10539 (N_10539,N_9593,N_9413);
nand U10540 (N_10540,N_9751,N_9455);
or U10541 (N_10541,N_9857,N_9047);
nor U10542 (N_10542,N_9089,N_9164);
and U10543 (N_10543,N_9898,N_9511);
xnor U10544 (N_10544,N_9434,N_9303);
nand U10545 (N_10545,N_9833,N_9238);
and U10546 (N_10546,N_9195,N_9529);
and U10547 (N_10547,N_9289,N_9903);
or U10548 (N_10548,N_9427,N_9378);
or U10549 (N_10549,N_9224,N_9371);
and U10550 (N_10550,N_9560,N_9040);
or U10551 (N_10551,N_9309,N_9639);
and U10552 (N_10552,N_9744,N_9599);
xor U10553 (N_10553,N_9876,N_9953);
nor U10554 (N_10554,N_9985,N_9987);
xnor U10555 (N_10555,N_9601,N_9717);
nor U10556 (N_10556,N_9983,N_9610);
and U10557 (N_10557,N_9341,N_9604);
xor U10558 (N_10558,N_9219,N_9238);
xnor U10559 (N_10559,N_9628,N_9873);
nor U10560 (N_10560,N_9163,N_9812);
or U10561 (N_10561,N_9870,N_9174);
nand U10562 (N_10562,N_9693,N_9656);
xnor U10563 (N_10563,N_9567,N_9942);
xor U10564 (N_10564,N_9620,N_9110);
nor U10565 (N_10565,N_9676,N_9021);
or U10566 (N_10566,N_9964,N_9022);
nor U10567 (N_10567,N_9619,N_9310);
nand U10568 (N_10568,N_9180,N_9426);
or U10569 (N_10569,N_9592,N_9266);
and U10570 (N_10570,N_9694,N_9411);
nor U10571 (N_10571,N_9792,N_9837);
or U10572 (N_10572,N_9037,N_9145);
nor U10573 (N_10573,N_9566,N_9626);
nand U10574 (N_10574,N_9309,N_9977);
and U10575 (N_10575,N_9793,N_9998);
and U10576 (N_10576,N_9772,N_9794);
nand U10577 (N_10577,N_9072,N_9502);
and U10578 (N_10578,N_9348,N_9228);
xnor U10579 (N_10579,N_9206,N_9189);
and U10580 (N_10580,N_9852,N_9314);
nand U10581 (N_10581,N_9934,N_9345);
nor U10582 (N_10582,N_9079,N_9952);
and U10583 (N_10583,N_9165,N_9225);
nor U10584 (N_10584,N_9672,N_9835);
or U10585 (N_10585,N_9470,N_9823);
nand U10586 (N_10586,N_9131,N_9514);
nor U10587 (N_10587,N_9646,N_9401);
and U10588 (N_10588,N_9663,N_9500);
or U10589 (N_10589,N_9363,N_9551);
nand U10590 (N_10590,N_9983,N_9806);
and U10591 (N_10591,N_9241,N_9124);
xnor U10592 (N_10592,N_9854,N_9456);
and U10593 (N_10593,N_9002,N_9383);
nor U10594 (N_10594,N_9719,N_9485);
nand U10595 (N_10595,N_9125,N_9970);
nor U10596 (N_10596,N_9260,N_9008);
xor U10597 (N_10597,N_9998,N_9887);
nor U10598 (N_10598,N_9253,N_9109);
xor U10599 (N_10599,N_9030,N_9477);
or U10600 (N_10600,N_9045,N_9746);
and U10601 (N_10601,N_9823,N_9897);
nand U10602 (N_10602,N_9756,N_9426);
or U10603 (N_10603,N_9920,N_9908);
nor U10604 (N_10604,N_9718,N_9751);
or U10605 (N_10605,N_9811,N_9420);
or U10606 (N_10606,N_9614,N_9955);
nand U10607 (N_10607,N_9933,N_9905);
xnor U10608 (N_10608,N_9977,N_9575);
xor U10609 (N_10609,N_9644,N_9630);
and U10610 (N_10610,N_9306,N_9971);
xnor U10611 (N_10611,N_9457,N_9733);
or U10612 (N_10612,N_9668,N_9073);
nand U10613 (N_10613,N_9279,N_9958);
xnor U10614 (N_10614,N_9711,N_9298);
or U10615 (N_10615,N_9154,N_9778);
nand U10616 (N_10616,N_9956,N_9063);
nor U10617 (N_10617,N_9371,N_9815);
nor U10618 (N_10618,N_9238,N_9186);
nand U10619 (N_10619,N_9992,N_9023);
or U10620 (N_10620,N_9054,N_9683);
xor U10621 (N_10621,N_9001,N_9408);
nand U10622 (N_10622,N_9509,N_9419);
or U10623 (N_10623,N_9819,N_9171);
and U10624 (N_10624,N_9856,N_9741);
and U10625 (N_10625,N_9930,N_9818);
or U10626 (N_10626,N_9324,N_9304);
or U10627 (N_10627,N_9155,N_9953);
nor U10628 (N_10628,N_9926,N_9146);
and U10629 (N_10629,N_9899,N_9963);
nor U10630 (N_10630,N_9025,N_9150);
nor U10631 (N_10631,N_9333,N_9443);
nor U10632 (N_10632,N_9984,N_9313);
or U10633 (N_10633,N_9741,N_9658);
or U10634 (N_10634,N_9206,N_9508);
xor U10635 (N_10635,N_9214,N_9928);
nor U10636 (N_10636,N_9259,N_9059);
nor U10637 (N_10637,N_9283,N_9020);
or U10638 (N_10638,N_9721,N_9713);
xor U10639 (N_10639,N_9265,N_9985);
nand U10640 (N_10640,N_9398,N_9533);
nor U10641 (N_10641,N_9906,N_9401);
nand U10642 (N_10642,N_9260,N_9053);
and U10643 (N_10643,N_9457,N_9344);
and U10644 (N_10644,N_9941,N_9957);
or U10645 (N_10645,N_9098,N_9467);
nand U10646 (N_10646,N_9097,N_9451);
or U10647 (N_10647,N_9638,N_9019);
nand U10648 (N_10648,N_9858,N_9041);
nor U10649 (N_10649,N_9494,N_9477);
nor U10650 (N_10650,N_9745,N_9724);
xnor U10651 (N_10651,N_9013,N_9544);
nor U10652 (N_10652,N_9017,N_9466);
xor U10653 (N_10653,N_9438,N_9168);
nor U10654 (N_10654,N_9322,N_9651);
nor U10655 (N_10655,N_9327,N_9830);
and U10656 (N_10656,N_9192,N_9605);
nand U10657 (N_10657,N_9009,N_9613);
and U10658 (N_10658,N_9744,N_9469);
nor U10659 (N_10659,N_9842,N_9642);
xor U10660 (N_10660,N_9658,N_9282);
xor U10661 (N_10661,N_9110,N_9955);
and U10662 (N_10662,N_9040,N_9419);
and U10663 (N_10663,N_9560,N_9441);
xor U10664 (N_10664,N_9697,N_9760);
and U10665 (N_10665,N_9257,N_9432);
nor U10666 (N_10666,N_9605,N_9878);
nand U10667 (N_10667,N_9843,N_9672);
xnor U10668 (N_10668,N_9513,N_9967);
and U10669 (N_10669,N_9262,N_9965);
nand U10670 (N_10670,N_9710,N_9244);
nor U10671 (N_10671,N_9970,N_9607);
and U10672 (N_10672,N_9041,N_9833);
nand U10673 (N_10673,N_9085,N_9226);
nor U10674 (N_10674,N_9326,N_9780);
or U10675 (N_10675,N_9312,N_9204);
or U10676 (N_10676,N_9037,N_9990);
nand U10677 (N_10677,N_9023,N_9830);
or U10678 (N_10678,N_9450,N_9494);
nand U10679 (N_10679,N_9425,N_9156);
or U10680 (N_10680,N_9785,N_9175);
or U10681 (N_10681,N_9358,N_9223);
xnor U10682 (N_10682,N_9403,N_9793);
or U10683 (N_10683,N_9890,N_9023);
or U10684 (N_10684,N_9277,N_9282);
xor U10685 (N_10685,N_9673,N_9979);
nand U10686 (N_10686,N_9951,N_9244);
or U10687 (N_10687,N_9678,N_9673);
or U10688 (N_10688,N_9966,N_9289);
nand U10689 (N_10689,N_9955,N_9667);
or U10690 (N_10690,N_9378,N_9544);
nand U10691 (N_10691,N_9802,N_9297);
nor U10692 (N_10692,N_9873,N_9362);
and U10693 (N_10693,N_9746,N_9969);
nand U10694 (N_10694,N_9795,N_9367);
nand U10695 (N_10695,N_9191,N_9717);
and U10696 (N_10696,N_9329,N_9130);
and U10697 (N_10697,N_9983,N_9868);
nor U10698 (N_10698,N_9378,N_9901);
nand U10699 (N_10699,N_9610,N_9427);
nor U10700 (N_10700,N_9230,N_9597);
nand U10701 (N_10701,N_9925,N_9063);
xnor U10702 (N_10702,N_9864,N_9248);
and U10703 (N_10703,N_9077,N_9543);
nand U10704 (N_10704,N_9215,N_9054);
or U10705 (N_10705,N_9135,N_9083);
or U10706 (N_10706,N_9929,N_9030);
or U10707 (N_10707,N_9361,N_9418);
xor U10708 (N_10708,N_9455,N_9610);
nor U10709 (N_10709,N_9097,N_9370);
xor U10710 (N_10710,N_9747,N_9235);
or U10711 (N_10711,N_9854,N_9133);
xor U10712 (N_10712,N_9504,N_9554);
and U10713 (N_10713,N_9961,N_9060);
nand U10714 (N_10714,N_9825,N_9727);
xnor U10715 (N_10715,N_9594,N_9651);
nand U10716 (N_10716,N_9596,N_9008);
xnor U10717 (N_10717,N_9314,N_9294);
nand U10718 (N_10718,N_9910,N_9618);
or U10719 (N_10719,N_9764,N_9067);
or U10720 (N_10720,N_9427,N_9426);
or U10721 (N_10721,N_9715,N_9620);
nor U10722 (N_10722,N_9470,N_9459);
nand U10723 (N_10723,N_9772,N_9488);
or U10724 (N_10724,N_9335,N_9346);
and U10725 (N_10725,N_9731,N_9789);
nand U10726 (N_10726,N_9178,N_9535);
nand U10727 (N_10727,N_9728,N_9808);
and U10728 (N_10728,N_9581,N_9386);
nor U10729 (N_10729,N_9340,N_9680);
nor U10730 (N_10730,N_9441,N_9094);
and U10731 (N_10731,N_9530,N_9327);
or U10732 (N_10732,N_9260,N_9386);
nor U10733 (N_10733,N_9244,N_9814);
and U10734 (N_10734,N_9226,N_9815);
nand U10735 (N_10735,N_9561,N_9638);
nand U10736 (N_10736,N_9047,N_9525);
nand U10737 (N_10737,N_9977,N_9877);
nand U10738 (N_10738,N_9261,N_9178);
nand U10739 (N_10739,N_9256,N_9006);
xor U10740 (N_10740,N_9196,N_9205);
nor U10741 (N_10741,N_9598,N_9965);
and U10742 (N_10742,N_9510,N_9343);
nor U10743 (N_10743,N_9376,N_9734);
and U10744 (N_10744,N_9334,N_9061);
nand U10745 (N_10745,N_9385,N_9805);
xnor U10746 (N_10746,N_9915,N_9767);
nor U10747 (N_10747,N_9908,N_9783);
nor U10748 (N_10748,N_9199,N_9570);
nand U10749 (N_10749,N_9784,N_9758);
and U10750 (N_10750,N_9302,N_9427);
nand U10751 (N_10751,N_9445,N_9941);
or U10752 (N_10752,N_9071,N_9725);
and U10753 (N_10753,N_9604,N_9222);
nand U10754 (N_10754,N_9993,N_9769);
or U10755 (N_10755,N_9501,N_9287);
nand U10756 (N_10756,N_9620,N_9650);
nand U10757 (N_10757,N_9327,N_9117);
or U10758 (N_10758,N_9681,N_9315);
nor U10759 (N_10759,N_9264,N_9215);
or U10760 (N_10760,N_9543,N_9523);
or U10761 (N_10761,N_9089,N_9079);
xnor U10762 (N_10762,N_9222,N_9602);
and U10763 (N_10763,N_9193,N_9770);
and U10764 (N_10764,N_9682,N_9046);
nor U10765 (N_10765,N_9422,N_9229);
nor U10766 (N_10766,N_9199,N_9072);
nor U10767 (N_10767,N_9046,N_9844);
nand U10768 (N_10768,N_9553,N_9738);
nor U10769 (N_10769,N_9663,N_9562);
nor U10770 (N_10770,N_9940,N_9012);
nor U10771 (N_10771,N_9530,N_9053);
or U10772 (N_10772,N_9858,N_9697);
xor U10773 (N_10773,N_9125,N_9788);
nand U10774 (N_10774,N_9305,N_9948);
nor U10775 (N_10775,N_9407,N_9409);
and U10776 (N_10776,N_9172,N_9194);
or U10777 (N_10777,N_9879,N_9818);
and U10778 (N_10778,N_9003,N_9246);
nand U10779 (N_10779,N_9764,N_9732);
nand U10780 (N_10780,N_9196,N_9928);
nand U10781 (N_10781,N_9484,N_9448);
nand U10782 (N_10782,N_9211,N_9612);
or U10783 (N_10783,N_9341,N_9708);
xor U10784 (N_10784,N_9767,N_9320);
xor U10785 (N_10785,N_9399,N_9296);
nand U10786 (N_10786,N_9309,N_9510);
and U10787 (N_10787,N_9909,N_9715);
and U10788 (N_10788,N_9139,N_9198);
and U10789 (N_10789,N_9806,N_9493);
nor U10790 (N_10790,N_9415,N_9993);
nand U10791 (N_10791,N_9933,N_9594);
nand U10792 (N_10792,N_9641,N_9476);
and U10793 (N_10793,N_9365,N_9588);
nor U10794 (N_10794,N_9541,N_9421);
or U10795 (N_10795,N_9153,N_9708);
xnor U10796 (N_10796,N_9141,N_9095);
and U10797 (N_10797,N_9927,N_9357);
and U10798 (N_10798,N_9044,N_9243);
and U10799 (N_10799,N_9920,N_9738);
nand U10800 (N_10800,N_9991,N_9504);
nor U10801 (N_10801,N_9833,N_9636);
or U10802 (N_10802,N_9387,N_9579);
and U10803 (N_10803,N_9983,N_9033);
nor U10804 (N_10804,N_9456,N_9123);
xnor U10805 (N_10805,N_9372,N_9541);
or U10806 (N_10806,N_9421,N_9370);
or U10807 (N_10807,N_9913,N_9914);
and U10808 (N_10808,N_9176,N_9537);
or U10809 (N_10809,N_9455,N_9314);
xnor U10810 (N_10810,N_9569,N_9939);
and U10811 (N_10811,N_9906,N_9542);
xor U10812 (N_10812,N_9889,N_9708);
or U10813 (N_10813,N_9092,N_9073);
nand U10814 (N_10814,N_9751,N_9825);
xor U10815 (N_10815,N_9023,N_9419);
or U10816 (N_10816,N_9977,N_9614);
xor U10817 (N_10817,N_9831,N_9946);
and U10818 (N_10818,N_9376,N_9208);
nand U10819 (N_10819,N_9155,N_9732);
nor U10820 (N_10820,N_9340,N_9274);
or U10821 (N_10821,N_9970,N_9426);
or U10822 (N_10822,N_9805,N_9378);
xnor U10823 (N_10823,N_9313,N_9454);
nand U10824 (N_10824,N_9644,N_9379);
or U10825 (N_10825,N_9954,N_9069);
nand U10826 (N_10826,N_9044,N_9248);
or U10827 (N_10827,N_9757,N_9922);
and U10828 (N_10828,N_9087,N_9031);
xor U10829 (N_10829,N_9355,N_9806);
nand U10830 (N_10830,N_9013,N_9888);
nor U10831 (N_10831,N_9373,N_9989);
or U10832 (N_10832,N_9171,N_9542);
nor U10833 (N_10833,N_9606,N_9428);
and U10834 (N_10834,N_9071,N_9239);
nand U10835 (N_10835,N_9283,N_9709);
nor U10836 (N_10836,N_9600,N_9980);
and U10837 (N_10837,N_9578,N_9564);
xor U10838 (N_10838,N_9336,N_9593);
or U10839 (N_10839,N_9263,N_9164);
or U10840 (N_10840,N_9874,N_9879);
and U10841 (N_10841,N_9315,N_9639);
nand U10842 (N_10842,N_9216,N_9851);
or U10843 (N_10843,N_9036,N_9422);
and U10844 (N_10844,N_9314,N_9304);
or U10845 (N_10845,N_9364,N_9648);
nor U10846 (N_10846,N_9877,N_9758);
xnor U10847 (N_10847,N_9398,N_9164);
nand U10848 (N_10848,N_9300,N_9468);
nand U10849 (N_10849,N_9171,N_9591);
nor U10850 (N_10850,N_9094,N_9323);
xnor U10851 (N_10851,N_9365,N_9904);
nor U10852 (N_10852,N_9035,N_9932);
or U10853 (N_10853,N_9371,N_9761);
or U10854 (N_10854,N_9293,N_9893);
nand U10855 (N_10855,N_9503,N_9029);
or U10856 (N_10856,N_9380,N_9773);
nor U10857 (N_10857,N_9645,N_9431);
nand U10858 (N_10858,N_9477,N_9379);
xnor U10859 (N_10859,N_9641,N_9346);
nor U10860 (N_10860,N_9042,N_9299);
nor U10861 (N_10861,N_9014,N_9230);
and U10862 (N_10862,N_9998,N_9362);
nand U10863 (N_10863,N_9409,N_9675);
or U10864 (N_10864,N_9077,N_9645);
or U10865 (N_10865,N_9893,N_9964);
or U10866 (N_10866,N_9083,N_9741);
nand U10867 (N_10867,N_9318,N_9684);
nor U10868 (N_10868,N_9179,N_9651);
or U10869 (N_10869,N_9401,N_9605);
or U10870 (N_10870,N_9482,N_9225);
and U10871 (N_10871,N_9607,N_9183);
or U10872 (N_10872,N_9124,N_9921);
and U10873 (N_10873,N_9725,N_9646);
nor U10874 (N_10874,N_9478,N_9418);
or U10875 (N_10875,N_9405,N_9130);
or U10876 (N_10876,N_9371,N_9812);
nand U10877 (N_10877,N_9762,N_9711);
xnor U10878 (N_10878,N_9324,N_9101);
nor U10879 (N_10879,N_9144,N_9902);
nor U10880 (N_10880,N_9400,N_9147);
nor U10881 (N_10881,N_9135,N_9154);
or U10882 (N_10882,N_9082,N_9375);
or U10883 (N_10883,N_9296,N_9840);
nand U10884 (N_10884,N_9444,N_9120);
or U10885 (N_10885,N_9787,N_9416);
or U10886 (N_10886,N_9098,N_9496);
and U10887 (N_10887,N_9168,N_9327);
or U10888 (N_10888,N_9619,N_9990);
nand U10889 (N_10889,N_9698,N_9706);
nor U10890 (N_10890,N_9345,N_9216);
nor U10891 (N_10891,N_9155,N_9607);
nand U10892 (N_10892,N_9335,N_9647);
nor U10893 (N_10893,N_9460,N_9815);
or U10894 (N_10894,N_9413,N_9092);
or U10895 (N_10895,N_9082,N_9941);
xor U10896 (N_10896,N_9196,N_9654);
xor U10897 (N_10897,N_9228,N_9351);
nor U10898 (N_10898,N_9791,N_9115);
or U10899 (N_10899,N_9817,N_9238);
and U10900 (N_10900,N_9885,N_9684);
nand U10901 (N_10901,N_9204,N_9922);
and U10902 (N_10902,N_9272,N_9915);
nand U10903 (N_10903,N_9771,N_9278);
nand U10904 (N_10904,N_9605,N_9651);
nor U10905 (N_10905,N_9553,N_9420);
or U10906 (N_10906,N_9687,N_9430);
nor U10907 (N_10907,N_9523,N_9408);
and U10908 (N_10908,N_9924,N_9141);
nor U10909 (N_10909,N_9547,N_9456);
and U10910 (N_10910,N_9019,N_9402);
and U10911 (N_10911,N_9433,N_9985);
nor U10912 (N_10912,N_9114,N_9223);
xor U10913 (N_10913,N_9341,N_9824);
nor U10914 (N_10914,N_9971,N_9541);
nor U10915 (N_10915,N_9732,N_9018);
xnor U10916 (N_10916,N_9238,N_9945);
nand U10917 (N_10917,N_9770,N_9744);
nor U10918 (N_10918,N_9369,N_9468);
or U10919 (N_10919,N_9877,N_9175);
nor U10920 (N_10920,N_9225,N_9286);
and U10921 (N_10921,N_9937,N_9155);
or U10922 (N_10922,N_9842,N_9500);
xor U10923 (N_10923,N_9189,N_9420);
or U10924 (N_10924,N_9755,N_9969);
or U10925 (N_10925,N_9317,N_9692);
or U10926 (N_10926,N_9312,N_9890);
xor U10927 (N_10927,N_9902,N_9638);
xor U10928 (N_10928,N_9877,N_9033);
nand U10929 (N_10929,N_9529,N_9434);
nand U10930 (N_10930,N_9530,N_9583);
or U10931 (N_10931,N_9455,N_9839);
or U10932 (N_10932,N_9205,N_9955);
xnor U10933 (N_10933,N_9099,N_9101);
nor U10934 (N_10934,N_9445,N_9516);
and U10935 (N_10935,N_9144,N_9361);
and U10936 (N_10936,N_9912,N_9891);
nand U10937 (N_10937,N_9296,N_9368);
nand U10938 (N_10938,N_9122,N_9343);
and U10939 (N_10939,N_9549,N_9056);
or U10940 (N_10940,N_9861,N_9270);
nor U10941 (N_10941,N_9506,N_9641);
nor U10942 (N_10942,N_9637,N_9420);
nand U10943 (N_10943,N_9374,N_9040);
xor U10944 (N_10944,N_9260,N_9093);
nor U10945 (N_10945,N_9163,N_9626);
nor U10946 (N_10946,N_9576,N_9898);
nor U10947 (N_10947,N_9239,N_9492);
or U10948 (N_10948,N_9798,N_9888);
and U10949 (N_10949,N_9507,N_9926);
xor U10950 (N_10950,N_9350,N_9438);
nand U10951 (N_10951,N_9143,N_9985);
nand U10952 (N_10952,N_9236,N_9304);
nand U10953 (N_10953,N_9767,N_9475);
nor U10954 (N_10954,N_9711,N_9992);
nand U10955 (N_10955,N_9138,N_9594);
nor U10956 (N_10956,N_9795,N_9383);
xnor U10957 (N_10957,N_9853,N_9814);
or U10958 (N_10958,N_9922,N_9814);
xnor U10959 (N_10959,N_9262,N_9717);
nor U10960 (N_10960,N_9921,N_9575);
xnor U10961 (N_10961,N_9867,N_9326);
nor U10962 (N_10962,N_9993,N_9941);
xnor U10963 (N_10963,N_9679,N_9863);
nor U10964 (N_10964,N_9224,N_9019);
xnor U10965 (N_10965,N_9635,N_9874);
and U10966 (N_10966,N_9012,N_9503);
xnor U10967 (N_10967,N_9776,N_9360);
xor U10968 (N_10968,N_9584,N_9140);
nand U10969 (N_10969,N_9900,N_9839);
xor U10970 (N_10970,N_9084,N_9903);
and U10971 (N_10971,N_9902,N_9593);
nand U10972 (N_10972,N_9919,N_9260);
xor U10973 (N_10973,N_9740,N_9196);
nor U10974 (N_10974,N_9848,N_9539);
nand U10975 (N_10975,N_9731,N_9921);
and U10976 (N_10976,N_9092,N_9932);
or U10977 (N_10977,N_9061,N_9455);
nand U10978 (N_10978,N_9822,N_9430);
xor U10979 (N_10979,N_9359,N_9949);
xor U10980 (N_10980,N_9423,N_9141);
xor U10981 (N_10981,N_9646,N_9641);
or U10982 (N_10982,N_9521,N_9463);
and U10983 (N_10983,N_9708,N_9558);
nor U10984 (N_10984,N_9127,N_9553);
nor U10985 (N_10985,N_9712,N_9745);
nor U10986 (N_10986,N_9843,N_9440);
nor U10987 (N_10987,N_9682,N_9963);
and U10988 (N_10988,N_9791,N_9973);
nand U10989 (N_10989,N_9415,N_9198);
nor U10990 (N_10990,N_9688,N_9161);
or U10991 (N_10991,N_9858,N_9644);
or U10992 (N_10992,N_9285,N_9633);
nor U10993 (N_10993,N_9274,N_9859);
xnor U10994 (N_10994,N_9278,N_9782);
nand U10995 (N_10995,N_9699,N_9020);
nor U10996 (N_10996,N_9132,N_9370);
nor U10997 (N_10997,N_9772,N_9630);
nand U10998 (N_10998,N_9827,N_9001);
or U10999 (N_10999,N_9491,N_9702);
nor U11000 (N_11000,N_10042,N_10315);
and U11001 (N_11001,N_10988,N_10407);
or U11002 (N_11002,N_10531,N_10076);
nor U11003 (N_11003,N_10183,N_10369);
nor U11004 (N_11004,N_10336,N_10921);
and U11005 (N_11005,N_10473,N_10895);
nor U11006 (N_11006,N_10200,N_10532);
and U11007 (N_11007,N_10801,N_10897);
nand U11008 (N_11008,N_10789,N_10162);
or U11009 (N_11009,N_10491,N_10421);
xnor U11010 (N_11010,N_10535,N_10630);
nand U11011 (N_11011,N_10140,N_10341);
nor U11012 (N_11012,N_10793,N_10425);
nand U11013 (N_11013,N_10869,N_10609);
xnor U11014 (N_11014,N_10119,N_10301);
nand U11015 (N_11015,N_10134,N_10956);
xor U11016 (N_11016,N_10181,N_10114);
xor U11017 (N_11017,N_10035,N_10733);
nand U11018 (N_11018,N_10252,N_10154);
nor U11019 (N_11019,N_10802,N_10120);
nand U11020 (N_11020,N_10461,N_10937);
nand U11021 (N_11021,N_10322,N_10554);
nor U11022 (N_11022,N_10659,N_10146);
nand U11023 (N_11023,N_10914,N_10069);
or U11024 (N_11024,N_10562,N_10040);
or U11025 (N_11025,N_10863,N_10185);
nand U11026 (N_11026,N_10498,N_10163);
xnor U11027 (N_11027,N_10688,N_10691);
nor U11028 (N_11028,N_10221,N_10822);
and U11029 (N_11029,N_10884,N_10788);
xnor U11030 (N_11030,N_10215,N_10497);
and U11031 (N_11031,N_10063,N_10036);
nand U11032 (N_11032,N_10482,N_10084);
or U11033 (N_11033,N_10826,N_10928);
nor U11034 (N_11034,N_10334,N_10957);
xnor U11035 (N_11035,N_10792,N_10285);
or U11036 (N_11036,N_10397,N_10318);
nand U11037 (N_11037,N_10774,N_10777);
xor U11038 (N_11038,N_10664,N_10748);
xnor U11039 (N_11039,N_10817,N_10098);
nand U11040 (N_11040,N_10027,N_10573);
nor U11041 (N_11041,N_10402,N_10850);
xor U11042 (N_11042,N_10606,N_10833);
nand U11043 (N_11043,N_10392,N_10130);
or U11044 (N_11044,N_10949,N_10809);
or U11045 (N_11045,N_10700,N_10601);
and U11046 (N_11046,N_10842,N_10616);
nor U11047 (N_11047,N_10489,N_10441);
or U11048 (N_11048,N_10864,N_10852);
nand U11049 (N_11049,N_10682,N_10198);
and U11050 (N_11050,N_10583,N_10180);
nand U11051 (N_11051,N_10654,N_10759);
or U11052 (N_11052,N_10045,N_10079);
or U11053 (N_11053,N_10212,N_10074);
xor U11054 (N_11054,N_10634,N_10553);
and U11055 (N_11055,N_10712,N_10480);
xor U11056 (N_11056,N_10560,N_10250);
xor U11057 (N_11057,N_10060,N_10575);
xnor U11058 (N_11058,N_10718,N_10039);
xor U11059 (N_11059,N_10605,N_10373);
xor U11060 (N_11060,N_10874,N_10371);
nor U11061 (N_11061,N_10326,N_10339);
and U11062 (N_11062,N_10711,N_10579);
or U11063 (N_11063,N_10628,N_10739);
xor U11064 (N_11064,N_10086,N_10526);
nand U11065 (N_11065,N_10727,N_10751);
and U11066 (N_11066,N_10451,N_10219);
nand U11067 (N_11067,N_10176,N_10106);
and U11068 (N_11068,N_10910,N_10135);
nor U11069 (N_11069,N_10061,N_10885);
nor U11070 (N_11070,N_10071,N_10843);
nand U11071 (N_11071,N_10714,N_10851);
or U11072 (N_11072,N_10433,N_10624);
and U11073 (N_11073,N_10314,N_10249);
and U11074 (N_11074,N_10379,N_10115);
nand U11075 (N_11075,N_10358,N_10158);
nor U11076 (N_11076,N_10048,N_10354);
nor U11077 (N_11077,N_10993,N_10858);
and U11078 (N_11078,N_10552,N_10933);
and U11079 (N_11079,N_10348,N_10335);
or U11080 (N_11080,N_10983,N_10656);
and U11081 (N_11081,N_10429,N_10089);
nand U11082 (N_11082,N_10149,N_10930);
or U11083 (N_11083,N_10571,N_10267);
nor U11084 (N_11084,N_10830,N_10588);
nor U11085 (N_11085,N_10184,N_10383);
xor U11086 (N_11086,N_10104,N_10686);
nand U11087 (N_11087,N_10598,N_10331);
nor U11088 (N_11088,N_10617,N_10368);
nor U11089 (N_11089,N_10168,N_10906);
nor U11090 (N_11090,N_10772,N_10935);
and U11091 (N_11091,N_10641,N_10110);
nor U11092 (N_11092,N_10235,N_10567);
nand U11093 (N_11093,N_10475,N_10723);
and U11094 (N_11094,N_10139,N_10595);
or U11095 (N_11095,N_10078,N_10261);
nor U11096 (N_11096,N_10838,N_10478);
nor U11097 (N_11097,N_10345,N_10224);
and U11098 (N_11098,N_10907,N_10969);
xor U11099 (N_11099,N_10298,N_10380);
xor U11100 (N_11100,N_10931,N_10097);
or U11101 (N_11101,N_10195,N_10898);
xnor U11102 (N_11102,N_10259,N_10513);
nand U11103 (N_11103,N_10753,N_10619);
or U11104 (N_11104,N_10414,N_10205);
or U11105 (N_11105,N_10924,N_10702);
or U11106 (N_11106,N_10133,N_10343);
and U11107 (N_11107,N_10613,N_10502);
xnor U11108 (N_11108,N_10389,N_10964);
xor U11109 (N_11109,N_10961,N_10465);
nor U11110 (N_11110,N_10207,N_10716);
nand U11111 (N_11111,N_10776,N_10311);
nand U11112 (N_11112,N_10481,N_10799);
nand U11113 (N_11113,N_10600,N_10735);
nor U11114 (N_11114,N_10410,N_10829);
or U11115 (N_11115,N_10728,N_10364);
nor U11116 (N_11116,N_10750,N_10277);
xor U11117 (N_11117,N_10965,N_10627);
and U11118 (N_11118,N_10746,N_10291);
nand U11119 (N_11119,N_10680,N_10679);
nor U11120 (N_11120,N_10674,N_10888);
nor U11121 (N_11121,N_10398,N_10941);
nand U11122 (N_11122,N_10860,N_10378);
xor U11123 (N_11123,N_10237,N_10846);
nor U11124 (N_11124,N_10572,N_10155);
nand U11125 (N_11125,N_10811,N_10596);
nand U11126 (N_11126,N_10515,N_10443);
and U11127 (N_11127,N_10954,N_10059);
xnor U11128 (N_11128,N_10943,N_10761);
or U11129 (N_11129,N_10555,N_10032);
nand U11130 (N_11130,N_10859,N_10376);
nor U11131 (N_11131,N_10775,N_10282);
xnor U11132 (N_11132,N_10058,N_10156);
nand U11133 (N_11133,N_10747,N_10835);
or U11134 (N_11134,N_10033,N_10883);
nand U11135 (N_11135,N_10960,N_10516);
or U11136 (N_11136,N_10824,N_10740);
or U11137 (N_11137,N_10743,N_10289);
nand U11138 (N_11138,N_10026,N_10268);
xor U11139 (N_11139,N_10657,N_10137);
and U11140 (N_11140,N_10002,N_10503);
nand U11141 (N_11141,N_10096,N_10161);
and U11142 (N_11142,N_10985,N_10464);
and U11143 (N_11143,N_10297,N_10790);
and U11144 (N_11144,N_10019,N_10785);
or U11145 (N_11145,N_10646,N_10794);
nand U11146 (N_11146,N_10390,N_10153);
nor U11147 (N_11147,N_10132,N_10187);
nor U11148 (N_11148,N_10210,N_10952);
or U11149 (N_11149,N_10206,N_10584);
and U11150 (N_11150,N_10013,N_10675);
nor U11151 (N_11151,N_10881,N_10493);
nor U11152 (N_11152,N_10085,N_10043);
xnor U11153 (N_11153,N_10338,N_10666);
xnor U11154 (N_11154,N_10321,N_10868);
nand U11155 (N_11155,N_10903,N_10696);
xor U11156 (N_11156,N_10866,N_10342);
nand U11157 (N_11157,N_10847,N_10430);
xnor U11158 (N_11158,N_10182,N_10405);
and U11159 (N_11159,N_10091,N_10370);
or U11160 (N_11160,N_10795,N_10099);
and U11161 (N_11161,N_10468,N_10107);
and U11162 (N_11162,N_10064,N_10934);
and U11163 (N_11163,N_10521,N_10056);
and U11164 (N_11164,N_10328,N_10360);
xor U11165 (N_11165,N_10418,N_10442);
and U11166 (N_11166,N_10999,N_10530);
nor U11167 (N_11167,N_10170,N_10455);
xor U11168 (N_11168,N_10239,N_10891);
nor U11169 (N_11169,N_10900,N_10982);
nand U11170 (N_11170,N_10118,N_10971);
xnor U11171 (N_11171,N_10361,N_10963);
and U11172 (N_11172,N_10485,N_10953);
nand U11173 (N_11173,N_10703,N_10265);
or U11174 (N_11174,N_10916,N_10009);
and U11175 (N_11175,N_10672,N_10220);
xor U11176 (N_11176,N_10626,N_10568);
nand U11177 (N_11177,N_10787,N_10917);
nand U11178 (N_11178,N_10055,N_10668);
nor U11179 (N_11179,N_10142,N_10100);
nand U11180 (N_11180,N_10374,N_10412);
nand U11181 (N_11181,N_10255,N_10940);
and U11182 (N_11182,N_10003,N_10523);
nand U11183 (N_11183,N_10528,N_10642);
nand U11184 (N_11184,N_10209,N_10236);
and U11185 (N_11185,N_10208,N_10806);
nor U11186 (N_11186,N_10367,N_10266);
nand U11187 (N_11187,N_10340,N_10403);
and U11188 (N_11188,N_10658,N_10426);
or U11189 (N_11189,N_10808,N_10016);
or U11190 (N_11190,N_10710,N_10014);
nor U11191 (N_11191,N_10660,N_10165);
or U11192 (N_11192,N_10292,N_10362);
xnor U11193 (N_11193,N_10452,N_10427);
nand U11194 (N_11194,N_10175,N_10823);
or U11195 (N_11195,N_10186,N_10512);
or U11196 (N_11196,N_10223,N_10986);
nand U11197 (N_11197,N_10325,N_10505);
xnor U11198 (N_11198,N_10857,N_10484);
or U11199 (N_11199,N_10307,N_10196);
nor U11200 (N_11200,N_10088,N_10745);
and U11201 (N_11201,N_10251,N_10438);
or U11202 (N_11202,N_10446,N_10872);
and U11203 (N_11203,N_10507,N_10669);
xnor U11204 (N_11204,N_10677,N_10462);
and U11205 (N_11205,N_10545,N_10603);
nor U11206 (N_11206,N_10765,N_10254);
nand U11207 (N_11207,N_10225,N_10877);
and U11208 (N_11208,N_10839,N_10030);
and U11209 (N_11209,N_10768,N_10477);
nand U11210 (N_11210,N_10457,N_10730);
xnor U11211 (N_11211,N_10721,N_10000);
or U11212 (N_11212,N_10913,N_10984);
and U11213 (N_11213,N_10814,N_10537);
or U11214 (N_11214,N_10923,N_10695);
nand U11215 (N_11215,N_10798,N_10976);
or U11216 (N_11216,N_10066,N_10729);
nand U11217 (N_11217,N_10580,N_10705);
or U11218 (N_11218,N_10350,N_10226);
or U11219 (N_11219,N_10440,N_10428);
nor U11220 (N_11220,N_10582,N_10749);
and U11221 (N_11221,N_10529,N_10391);
nand U11222 (N_11222,N_10919,N_10577);
and U11223 (N_11223,N_10661,N_10889);
and U11224 (N_11224,N_10001,N_10275);
xnor U11225 (N_11225,N_10278,N_10692);
nand U11226 (N_11226,N_10308,N_10676);
xnor U11227 (N_11227,N_10458,N_10681);
nor U11228 (N_11228,N_10166,N_10122);
nand U11229 (N_11229,N_10887,N_10262);
nor U11230 (N_11230,N_10217,N_10356);
or U11231 (N_11231,N_10805,N_10241);
nor U11232 (N_11232,N_10294,N_10720);
and U11233 (N_11233,N_10296,N_10796);
or U11234 (N_11234,N_10509,N_10243);
and U11235 (N_11235,N_10434,N_10770);
nand U11236 (N_11236,N_10570,N_10757);
nand U11237 (N_11237,N_10202,N_10604);
nand U11238 (N_11238,N_10621,N_10966);
or U11239 (N_11239,N_10432,N_10150);
and U11240 (N_11240,N_10848,N_10693);
xnor U11241 (N_11241,N_10422,N_10612);
nand U11242 (N_11242,N_10652,N_10488);
or U11243 (N_11243,N_10145,N_10673);
and U11244 (N_11244,N_10786,N_10593);
xor U11245 (N_11245,N_10062,N_10707);
nor U11246 (N_11246,N_10445,N_10270);
or U11247 (N_11247,N_10147,N_10853);
or U11248 (N_11248,N_10229,N_10346);
and U11249 (N_11249,N_10645,N_10920);
or U11250 (N_11250,N_10093,N_10247);
nand U11251 (N_11251,N_10722,N_10831);
xor U11252 (N_11252,N_10047,N_10663);
and U11253 (N_11253,N_10527,N_10385);
and U11254 (N_11254,N_10274,N_10494);
or U11255 (N_11255,N_10944,N_10670);
nand U11256 (N_11256,N_10594,N_10581);
or U11257 (N_11257,N_10375,N_10886);
xor U11258 (N_11258,N_10908,N_10077);
nor U11259 (N_11259,N_10685,N_10447);
xnor U11260 (N_11260,N_10306,N_10544);
xnor U11261 (N_11261,N_10193,N_10233);
or U11262 (N_11262,N_10312,N_10766);
or U11263 (N_11263,N_10736,N_10500);
nor U11264 (N_11264,N_10317,N_10929);
xor U11265 (N_11265,N_10649,N_10726);
nand U11266 (N_11266,N_10420,N_10615);
or U11267 (N_11267,N_10762,N_10015);
and U11268 (N_11268,N_10448,N_10994);
and U11269 (N_11269,N_10901,N_10576);
and U11270 (N_11270,N_10067,N_10836);
xnor U11271 (N_11271,N_10978,N_10618);
xnor U11272 (N_11272,N_10893,N_10820);
and U11273 (N_11273,N_10607,N_10813);
or U11274 (N_11274,N_10347,N_10591);
nor U11275 (N_11275,N_10939,N_10017);
nor U11276 (N_11276,N_10539,N_10495);
xnor U11277 (N_11277,N_10393,N_10540);
xnor U11278 (N_11278,N_10499,N_10810);
nand U11279 (N_11279,N_10138,N_10684);
or U11280 (N_11280,N_10011,N_10911);
and U11281 (N_11281,N_10525,N_10875);
nor U11282 (N_11282,N_10754,N_10372);
and U11283 (N_11283,N_10199,N_10556);
nand U11284 (N_11284,N_10201,N_10053);
or U11285 (N_11285,N_10087,N_10651);
or U11286 (N_11286,N_10821,N_10123);
or U11287 (N_11287,N_10942,N_10037);
or U11288 (N_11288,N_10044,N_10510);
nand U11289 (N_11289,N_10778,N_10483);
nand U11290 (N_11290,N_10102,N_10173);
nor U11291 (N_11291,N_10396,N_10041);
and U11292 (N_11292,N_10989,N_10366);
nand U11293 (N_11293,N_10968,N_10126);
or U11294 (N_11294,N_10713,N_10611);
nand U11295 (N_11295,N_10293,N_10807);
and U11296 (N_11296,N_10424,N_10644);
nor U11297 (N_11297,N_10861,N_10948);
and U11298 (N_11298,N_10980,N_10678);
nor U11299 (N_11299,N_10330,N_10648);
nand U11300 (N_11300,N_10622,N_10918);
nand U11301 (N_11301,N_10052,N_10637);
nand U11302 (N_11302,N_10784,N_10511);
or U11303 (N_11303,N_10951,N_10141);
or U11304 (N_11304,N_10541,N_10479);
xor U11305 (N_11305,N_10408,N_10234);
and U11306 (N_11306,N_10862,N_10231);
or U11307 (N_11307,N_10319,N_10734);
xor U11308 (N_11308,N_10534,N_10671);
nor U11309 (N_11309,N_10188,N_10463);
and U11310 (N_11310,N_10629,N_10871);
and U11311 (N_11311,N_10082,N_10365);
xor U11312 (N_11312,N_10073,N_10812);
nor U11313 (N_11313,N_10998,N_10417);
nor U11314 (N_11314,N_10894,N_10882);
nand U11315 (N_11315,N_10228,N_10771);
or U11316 (N_11316,N_10909,N_10625);
nor U11317 (N_11317,N_10218,N_10697);
or U11318 (N_11318,N_10466,N_10880);
xnor U11319 (N_11319,N_10992,N_10873);
nand U11320 (N_11320,N_10599,N_10551);
xnor U11321 (N_11321,N_10631,N_10117);
or U11322 (N_11322,N_10431,N_10548);
nand U11323 (N_11323,N_10271,N_10470);
and U11324 (N_11324,N_10148,N_10837);
xnor U11325 (N_11325,N_10590,N_10204);
nor U11326 (N_11326,N_10962,N_10709);
and U11327 (N_11327,N_10159,N_10213);
and U11328 (N_11328,N_10349,N_10151);
and U11329 (N_11329,N_10113,N_10890);
xor U11330 (N_11330,N_10737,N_10804);
and U11331 (N_11331,N_10870,N_10245);
nand U11332 (N_11332,N_10967,N_10828);
or U11333 (N_11333,N_10021,N_10051);
and U11334 (N_11334,N_10756,N_10487);
nor U11335 (N_11335,N_10004,N_10701);
and U11336 (N_11336,N_10057,N_10844);
nor U11337 (N_11337,N_10549,N_10996);
and U11338 (N_11338,N_10423,N_10955);
and U11339 (N_11339,N_10501,N_10409);
or U11340 (N_11340,N_10496,N_10781);
nand U11341 (N_11341,N_10018,N_10263);
nor U11342 (N_11342,N_10344,N_10623);
xor U11343 (N_11343,N_10127,N_10633);
nor U11344 (N_11344,N_10782,N_10995);
nand U11345 (N_11345,N_10300,N_10116);
nor U11346 (N_11346,N_10103,N_10359);
or U11347 (N_11347,N_10460,N_10650);
nor U11348 (N_11348,N_10172,N_10327);
xor U11349 (N_11349,N_10602,N_10449);
nand U11350 (N_11350,N_10932,N_10111);
nand U11351 (N_11351,N_10827,N_10387);
xnor U11352 (N_11352,N_10474,N_10230);
nand U11353 (N_11353,N_10081,N_10284);
xnor U11354 (N_11354,N_10302,N_10744);
nor U11355 (N_11355,N_10467,N_10101);
xor U11356 (N_11356,N_10610,N_10550);
nor U11357 (N_11357,N_10717,N_10471);
and U11358 (N_11358,N_10905,N_10492);
xnor U11359 (N_11359,N_10958,N_10049);
and U11360 (N_11360,N_10783,N_10286);
or U11361 (N_11361,N_10006,N_10879);
or U11362 (N_11362,N_10401,N_10972);
nand U11363 (N_11363,N_10171,N_10276);
and U11364 (N_11364,N_10586,N_10760);
or U11365 (N_11365,N_10272,N_10620);
xnor U11366 (N_11366,N_10752,N_10856);
xor U11367 (N_11367,N_10108,N_10504);
xnor U11368 (N_11368,N_10197,N_10936);
or U11369 (N_11369,N_10324,N_10357);
and U11370 (N_11370,N_10981,N_10453);
or U11371 (N_11371,N_10258,N_10520);
or U11372 (N_11372,N_10769,N_10090);
and U11373 (N_11373,N_10436,N_10022);
nand U11374 (N_11374,N_10143,N_10028);
and U11375 (N_11375,N_10416,N_10855);
xnor U11376 (N_11376,N_10012,N_10095);
or U11377 (N_11377,N_10557,N_10411);
or U11378 (N_11378,N_10518,N_10456);
nand U11379 (N_11379,N_10922,N_10506);
and U11380 (N_11380,N_10585,N_10260);
or U11381 (N_11381,N_10708,N_10072);
nand U11382 (N_11382,N_10136,N_10508);
or U11383 (N_11383,N_10394,N_10899);
or U11384 (N_11384,N_10203,N_10083);
and U11385 (N_11385,N_10818,N_10945);
and U11386 (N_11386,N_10815,N_10105);
and U11387 (N_11387,N_10987,N_10587);
or U11388 (N_11388,N_10240,N_10608);
and U11389 (N_11389,N_10636,N_10164);
and U11390 (N_11390,N_10316,N_10382);
and U11391 (N_11391,N_10192,N_10667);
and U11392 (N_11392,N_10538,N_10564);
and U11393 (N_11393,N_10732,N_10386);
nor U11394 (N_11394,N_10803,N_10635);
nor U11395 (N_11395,N_10329,N_10283);
and U11396 (N_11396,N_10699,N_10706);
xnor U11397 (N_11397,N_10938,N_10832);
and U11398 (N_11398,N_10337,N_10303);
and U11399 (N_11399,N_10310,N_10991);
nand U11400 (N_11400,N_10112,N_10758);
and U11401 (N_11401,N_10773,N_10522);
or U11402 (N_11402,N_10476,N_10640);
xor U11403 (N_11403,N_10947,N_10253);
nor U11404 (N_11404,N_10242,N_10194);
or U11405 (N_11405,N_10280,N_10975);
nand U11406 (N_11406,N_10400,N_10065);
nand U11407 (N_11407,N_10574,N_10323);
and U11408 (N_11408,N_10121,N_10742);
nor U11409 (N_11409,N_10977,N_10320);
nor U11410 (N_11410,N_10313,N_10524);
or U11411 (N_11411,N_10912,N_10309);
nand U11412 (N_11412,N_10388,N_10264);
nand U11413 (N_11413,N_10517,N_10160);
and U11414 (N_11414,N_10287,N_10174);
and U11415 (N_11415,N_10486,N_10381);
nor U11416 (N_11416,N_10655,N_10780);
xnor U11417 (N_11417,N_10566,N_10269);
and U11418 (N_11418,N_10689,N_10819);
nand U11419 (N_11419,N_10273,N_10189);
nor U11420 (N_11420,N_10915,N_10169);
or U11421 (N_11421,N_10377,N_10005);
nand U11422 (N_11422,N_10597,N_10878);
nor U11423 (N_11423,N_10970,N_10514);
nand U11424 (N_11424,N_10020,N_10959);
and U11425 (N_11425,N_10238,N_10070);
or U11426 (N_11426,N_10638,N_10926);
and U11427 (N_11427,N_10248,N_10413);
or U11428 (N_11428,N_10854,N_10643);
or U11429 (N_11429,N_10279,N_10865);
xor U11430 (N_11430,N_10904,N_10450);
and U11431 (N_11431,N_10214,N_10244);
and U11432 (N_11432,N_10876,N_10216);
nand U11433 (N_11433,N_10469,N_10825);
or U11434 (N_11434,N_10351,N_10288);
xor U11435 (N_11435,N_10800,N_10867);
or U11436 (N_11436,N_10724,N_10179);
and U11437 (N_11437,N_10536,N_10764);
and U11438 (N_11438,N_10419,N_10395);
xor U11439 (N_11439,N_10925,N_10589);
or U11440 (N_11440,N_10472,N_10025);
or U11441 (N_11441,N_10054,N_10738);
nor U11442 (N_11442,N_10845,N_10257);
nand U11443 (N_11443,N_10979,N_10834);
xnor U11444 (N_11444,N_10731,N_10694);
nor U11445 (N_11445,N_10896,N_10653);
nand U11446 (N_11446,N_10816,N_10592);
nand U11447 (N_11447,N_10211,N_10719);
nand U11448 (N_11448,N_10565,N_10755);
nand U11449 (N_11449,N_10352,N_10129);
nand U11450 (N_11450,N_10125,N_10007);
nor U11451 (N_11451,N_10791,N_10715);
and U11452 (N_11452,N_10167,N_10191);
or U11453 (N_11453,N_10152,N_10665);
and U11454 (N_11454,N_10190,N_10632);
and U11455 (N_11455,N_10068,N_10290);
xor U11456 (N_11456,N_10333,N_10038);
and U11457 (N_11457,N_10973,N_10704);
or U11458 (N_11458,N_10406,N_10841);
nand U11459 (N_11459,N_10010,N_10384);
or U11460 (N_11460,N_10454,N_10144);
xor U11461 (N_11461,N_10698,N_10974);
or U11462 (N_11462,N_10797,N_10543);
and U11463 (N_11463,N_10767,N_10533);
nand U11464 (N_11464,N_10990,N_10256);
nor U11465 (N_11465,N_10563,N_10415);
or U11466 (N_11466,N_10950,N_10295);
or U11467 (N_11467,N_10178,N_10542);
nor U11468 (N_11468,N_10779,N_10569);
and U11469 (N_11469,N_10662,N_10490);
or U11470 (N_11470,N_10687,N_10614);
or U11471 (N_11471,N_10094,N_10222);
nor U11472 (N_11472,N_10034,N_10092);
nand U11473 (N_11473,N_10299,N_10639);
and U11474 (N_11474,N_10399,N_10741);
nor U11475 (N_11475,N_10459,N_10075);
xor U11476 (N_11476,N_10023,N_10177);
and U11477 (N_11477,N_10031,N_10332);
nor U11478 (N_11478,N_10547,N_10437);
and U11479 (N_11479,N_10559,N_10849);
xnor U11480 (N_11480,N_10683,N_10128);
and U11481 (N_11481,N_10546,N_10444);
or U11482 (N_11482,N_10578,N_10404);
nand U11483 (N_11483,N_10046,N_10725);
or U11484 (N_11484,N_10435,N_10281);
and U11485 (N_11485,N_10008,N_10157);
nand U11486 (N_11486,N_10080,N_10927);
xor U11487 (N_11487,N_10561,N_10519);
nand U11488 (N_11488,N_10353,N_10232);
and U11489 (N_11489,N_10946,N_10227);
or U11490 (N_11490,N_10131,N_10109);
nor U11491 (N_11491,N_10246,N_10355);
and U11492 (N_11492,N_10558,N_10304);
nor U11493 (N_11493,N_10029,N_10892);
and U11494 (N_11494,N_10050,N_10305);
xnor U11495 (N_11495,N_10363,N_10439);
nor U11496 (N_11496,N_10763,N_10997);
nand U11497 (N_11497,N_10690,N_10124);
nor U11498 (N_11498,N_10902,N_10024);
and U11499 (N_11499,N_10840,N_10647);
and U11500 (N_11500,N_10483,N_10454);
or U11501 (N_11501,N_10373,N_10832);
nand U11502 (N_11502,N_10410,N_10755);
nor U11503 (N_11503,N_10808,N_10674);
nor U11504 (N_11504,N_10841,N_10394);
or U11505 (N_11505,N_10829,N_10926);
and U11506 (N_11506,N_10034,N_10273);
and U11507 (N_11507,N_10087,N_10287);
nor U11508 (N_11508,N_10283,N_10644);
or U11509 (N_11509,N_10919,N_10708);
nand U11510 (N_11510,N_10087,N_10604);
and U11511 (N_11511,N_10425,N_10787);
nand U11512 (N_11512,N_10383,N_10349);
or U11513 (N_11513,N_10378,N_10256);
nand U11514 (N_11514,N_10267,N_10570);
nor U11515 (N_11515,N_10502,N_10456);
or U11516 (N_11516,N_10671,N_10581);
or U11517 (N_11517,N_10454,N_10894);
and U11518 (N_11518,N_10354,N_10946);
nand U11519 (N_11519,N_10907,N_10569);
nand U11520 (N_11520,N_10048,N_10193);
nand U11521 (N_11521,N_10920,N_10766);
xnor U11522 (N_11522,N_10945,N_10990);
and U11523 (N_11523,N_10418,N_10030);
nand U11524 (N_11524,N_10005,N_10542);
nand U11525 (N_11525,N_10899,N_10166);
xor U11526 (N_11526,N_10225,N_10960);
xnor U11527 (N_11527,N_10448,N_10031);
nand U11528 (N_11528,N_10945,N_10778);
xor U11529 (N_11529,N_10773,N_10422);
and U11530 (N_11530,N_10162,N_10819);
nand U11531 (N_11531,N_10378,N_10191);
xnor U11532 (N_11532,N_10681,N_10839);
nand U11533 (N_11533,N_10841,N_10490);
xor U11534 (N_11534,N_10008,N_10666);
nor U11535 (N_11535,N_10753,N_10435);
nor U11536 (N_11536,N_10918,N_10470);
nand U11537 (N_11537,N_10944,N_10608);
or U11538 (N_11538,N_10432,N_10668);
xor U11539 (N_11539,N_10356,N_10760);
nand U11540 (N_11540,N_10965,N_10859);
and U11541 (N_11541,N_10557,N_10575);
nand U11542 (N_11542,N_10818,N_10957);
or U11543 (N_11543,N_10071,N_10915);
or U11544 (N_11544,N_10564,N_10994);
nor U11545 (N_11545,N_10342,N_10466);
and U11546 (N_11546,N_10294,N_10189);
xor U11547 (N_11547,N_10860,N_10402);
nand U11548 (N_11548,N_10177,N_10182);
or U11549 (N_11549,N_10057,N_10881);
xor U11550 (N_11550,N_10071,N_10880);
xor U11551 (N_11551,N_10091,N_10016);
and U11552 (N_11552,N_10147,N_10652);
xor U11553 (N_11553,N_10967,N_10991);
xnor U11554 (N_11554,N_10136,N_10026);
nor U11555 (N_11555,N_10696,N_10129);
nor U11556 (N_11556,N_10134,N_10860);
and U11557 (N_11557,N_10588,N_10214);
nor U11558 (N_11558,N_10633,N_10774);
xnor U11559 (N_11559,N_10716,N_10746);
and U11560 (N_11560,N_10350,N_10070);
or U11561 (N_11561,N_10402,N_10016);
nand U11562 (N_11562,N_10820,N_10947);
nor U11563 (N_11563,N_10435,N_10716);
nand U11564 (N_11564,N_10407,N_10119);
and U11565 (N_11565,N_10300,N_10176);
nand U11566 (N_11566,N_10539,N_10756);
xor U11567 (N_11567,N_10445,N_10033);
and U11568 (N_11568,N_10963,N_10035);
nand U11569 (N_11569,N_10378,N_10795);
nand U11570 (N_11570,N_10345,N_10557);
nor U11571 (N_11571,N_10303,N_10619);
or U11572 (N_11572,N_10688,N_10295);
xor U11573 (N_11573,N_10094,N_10249);
xor U11574 (N_11574,N_10729,N_10949);
nor U11575 (N_11575,N_10564,N_10112);
nand U11576 (N_11576,N_10809,N_10158);
nor U11577 (N_11577,N_10888,N_10162);
and U11578 (N_11578,N_10073,N_10402);
xnor U11579 (N_11579,N_10609,N_10839);
or U11580 (N_11580,N_10932,N_10495);
nor U11581 (N_11581,N_10385,N_10516);
and U11582 (N_11582,N_10753,N_10185);
and U11583 (N_11583,N_10202,N_10167);
or U11584 (N_11584,N_10968,N_10727);
nand U11585 (N_11585,N_10307,N_10368);
and U11586 (N_11586,N_10322,N_10231);
xor U11587 (N_11587,N_10430,N_10054);
and U11588 (N_11588,N_10768,N_10849);
nor U11589 (N_11589,N_10799,N_10644);
nor U11590 (N_11590,N_10670,N_10123);
and U11591 (N_11591,N_10745,N_10216);
or U11592 (N_11592,N_10796,N_10048);
nand U11593 (N_11593,N_10050,N_10332);
or U11594 (N_11594,N_10808,N_10620);
xor U11595 (N_11595,N_10234,N_10268);
or U11596 (N_11596,N_10702,N_10162);
xnor U11597 (N_11597,N_10107,N_10436);
and U11598 (N_11598,N_10130,N_10285);
or U11599 (N_11599,N_10041,N_10077);
nor U11600 (N_11600,N_10231,N_10295);
nand U11601 (N_11601,N_10637,N_10064);
nand U11602 (N_11602,N_10407,N_10360);
nand U11603 (N_11603,N_10400,N_10464);
nor U11604 (N_11604,N_10618,N_10191);
or U11605 (N_11605,N_10236,N_10918);
or U11606 (N_11606,N_10188,N_10985);
xnor U11607 (N_11607,N_10336,N_10281);
or U11608 (N_11608,N_10822,N_10149);
nor U11609 (N_11609,N_10988,N_10870);
xnor U11610 (N_11610,N_10453,N_10546);
xor U11611 (N_11611,N_10562,N_10758);
and U11612 (N_11612,N_10393,N_10898);
and U11613 (N_11613,N_10242,N_10424);
or U11614 (N_11614,N_10877,N_10794);
xor U11615 (N_11615,N_10859,N_10611);
or U11616 (N_11616,N_10122,N_10957);
and U11617 (N_11617,N_10770,N_10975);
nand U11618 (N_11618,N_10913,N_10832);
xnor U11619 (N_11619,N_10490,N_10221);
or U11620 (N_11620,N_10966,N_10193);
xnor U11621 (N_11621,N_10294,N_10871);
nand U11622 (N_11622,N_10285,N_10051);
or U11623 (N_11623,N_10763,N_10064);
or U11624 (N_11624,N_10632,N_10400);
or U11625 (N_11625,N_10708,N_10355);
nand U11626 (N_11626,N_10391,N_10375);
or U11627 (N_11627,N_10607,N_10787);
nor U11628 (N_11628,N_10683,N_10597);
nor U11629 (N_11629,N_10530,N_10292);
xor U11630 (N_11630,N_10385,N_10758);
xor U11631 (N_11631,N_10037,N_10908);
and U11632 (N_11632,N_10257,N_10181);
nand U11633 (N_11633,N_10105,N_10678);
and U11634 (N_11634,N_10133,N_10336);
nor U11635 (N_11635,N_10194,N_10687);
nor U11636 (N_11636,N_10452,N_10540);
xor U11637 (N_11637,N_10291,N_10180);
nor U11638 (N_11638,N_10900,N_10049);
nand U11639 (N_11639,N_10950,N_10523);
nor U11640 (N_11640,N_10258,N_10945);
xor U11641 (N_11641,N_10449,N_10173);
xnor U11642 (N_11642,N_10343,N_10748);
or U11643 (N_11643,N_10195,N_10668);
or U11644 (N_11644,N_10421,N_10378);
and U11645 (N_11645,N_10963,N_10951);
nor U11646 (N_11646,N_10215,N_10878);
xor U11647 (N_11647,N_10357,N_10369);
nand U11648 (N_11648,N_10097,N_10552);
or U11649 (N_11649,N_10216,N_10041);
and U11650 (N_11650,N_10245,N_10551);
xor U11651 (N_11651,N_10891,N_10263);
xor U11652 (N_11652,N_10073,N_10827);
nor U11653 (N_11653,N_10816,N_10713);
nand U11654 (N_11654,N_10635,N_10381);
xor U11655 (N_11655,N_10251,N_10612);
and U11656 (N_11656,N_10713,N_10164);
and U11657 (N_11657,N_10650,N_10673);
nand U11658 (N_11658,N_10053,N_10247);
nor U11659 (N_11659,N_10938,N_10395);
nand U11660 (N_11660,N_10166,N_10681);
and U11661 (N_11661,N_10583,N_10382);
and U11662 (N_11662,N_10176,N_10098);
nand U11663 (N_11663,N_10010,N_10742);
xnor U11664 (N_11664,N_10463,N_10097);
and U11665 (N_11665,N_10385,N_10761);
xor U11666 (N_11666,N_10628,N_10173);
nor U11667 (N_11667,N_10830,N_10061);
nor U11668 (N_11668,N_10246,N_10133);
xor U11669 (N_11669,N_10202,N_10966);
and U11670 (N_11670,N_10524,N_10038);
xnor U11671 (N_11671,N_10326,N_10201);
xor U11672 (N_11672,N_10400,N_10688);
or U11673 (N_11673,N_10704,N_10887);
nor U11674 (N_11674,N_10125,N_10934);
nand U11675 (N_11675,N_10874,N_10824);
or U11676 (N_11676,N_10381,N_10827);
nor U11677 (N_11677,N_10119,N_10773);
or U11678 (N_11678,N_10789,N_10870);
or U11679 (N_11679,N_10567,N_10723);
nor U11680 (N_11680,N_10329,N_10946);
xor U11681 (N_11681,N_10537,N_10154);
or U11682 (N_11682,N_10109,N_10084);
nor U11683 (N_11683,N_10338,N_10633);
nor U11684 (N_11684,N_10215,N_10563);
and U11685 (N_11685,N_10094,N_10599);
nand U11686 (N_11686,N_10864,N_10506);
nor U11687 (N_11687,N_10690,N_10270);
and U11688 (N_11688,N_10974,N_10023);
xor U11689 (N_11689,N_10479,N_10910);
nand U11690 (N_11690,N_10562,N_10992);
nand U11691 (N_11691,N_10883,N_10453);
or U11692 (N_11692,N_10564,N_10135);
nand U11693 (N_11693,N_10123,N_10792);
and U11694 (N_11694,N_10965,N_10021);
xor U11695 (N_11695,N_10963,N_10229);
xnor U11696 (N_11696,N_10633,N_10118);
or U11697 (N_11697,N_10974,N_10424);
nor U11698 (N_11698,N_10772,N_10894);
xnor U11699 (N_11699,N_10150,N_10902);
or U11700 (N_11700,N_10339,N_10596);
nor U11701 (N_11701,N_10473,N_10220);
nor U11702 (N_11702,N_10121,N_10636);
and U11703 (N_11703,N_10818,N_10492);
nand U11704 (N_11704,N_10294,N_10644);
nor U11705 (N_11705,N_10747,N_10783);
xor U11706 (N_11706,N_10767,N_10212);
and U11707 (N_11707,N_10706,N_10906);
and U11708 (N_11708,N_10259,N_10005);
nor U11709 (N_11709,N_10054,N_10259);
or U11710 (N_11710,N_10686,N_10756);
xnor U11711 (N_11711,N_10153,N_10671);
nand U11712 (N_11712,N_10189,N_10337);
or U11713 (N_11713,N_10460,N_10482);
and U11714 (N_11714,N_10592,N_10571);
xnor U11715 (N_11715,N_10682,N_10375);
or U11716 (N_11716,N_10390,N_10590);
and U11717 (N_11717,N_10839,N_10981);
or U11718 (N_11718,N_10580,N_10121);
and U11719 (N_11719,N_10918,N_10471);
nand U11720 (N_11720,N_10639,N_10204);
and U11721 (N_11721,N_10020,N_10916);
nor U11722 (N_11722,N_10532,N_10012);
and U11723 (N_11723,N_10335,N_10712);
nor U11724 (N_11724,N_10096,N_10234);
or U11725 (N_11725,N_10687,N_10591);
nor U11726 (N_11726,N_10053,N_10143);
or U11727 (N_11727,N_10538,N_10513);
xor U11728 (N_11728,N_10319,N_10134);
or U11729 (N_11729,N_10904,N_10782);
xor U11730 (N_11730,N_10302,N_10603);
and U11731 (N_11731,N_10649,N_10305);
and U11732 (N_11732,N_10548,N_10493);
or U11733 (N_11733,N_10911,N_10906);
nand U11734 (N_11734,N_10940,N_10589);
or U11735 (N_11735,N_10655,N_10991);
or U11736 (N_11736,N_10539,N_10318);
and U11737 (N_11737,N_10156,N_10407);
and U11738 (N_11738,N_10914,N_10010);
nand U11739 (N_11739,N_10331,N_10232);
nor U11740 (N_11740,N_10846,N_10169);
xnor U11741 (N_11741,N_10603,N_10178);
or U11742 (N_11742,N_10523,N_10228);
nand U11743 (N_11743,N_10119,N_10389);
and U11744 (N_11744,N_10181,N_10686);
nand U11745 (N_11745,N_10014,N_10251);
nor U11746 (N_11746,N_10299,N_10823);
nor U11747 (N_11747,N_10198,N_10441);
or U11748 (N_11748,N_10368,N_10635);
nand U11749 (N_11749,N_10155,N_10083);
xnor U11750 (N_11750,N_10831,N_10545);
or U11751 (N_11751,N_10779,N_10573);
nand U11752 (N_11752,N_10475,N_10173);
nor U11753 (N_11753,N_10005,N_10264);
xnor U11754 (N_11754,N_10824,N_10732);
xor U11755 (N_11755,N_10765,N_10444);
nand U11756 (N_11756,N_10762,N_10955);
and U11757 (N_11757,N_10211,N_10934);
xor U11758 (N_11758,N_10240,N_10171);
and U11759 (N_11759,N_10509,N_10810);
or U11760 (N_11760,N_10422,N_10672);
nor U11761 (N_11761,N_10051,N_10546);
nand U11762 (N_11762,N_10008,N_10952);
and U11763 (N_11763,N_10668,N_10001);
xnor U11764 (N_11764,N_10820,N_10840);
or U11765 (N_11765,N_10935,N_10717);
nor U11766 (N_11766,N_10431,N_10116);
and U11767 (N_11767,N_10339,N_10609);
and U11768 (N_11768,N_10445,N_10208);
and U11769 (N_11769,N_10712,N_10860);
and U11770 (N_11770,N_10907,N_10548);
or U11771 (N_11771,N_10534,N_10861);
and U11772 (N_11772,N_10220,N_10934);
nand U11773 (N_11773,N_10535,N_10992);
and U11774 (N_11774,N_10087,N_10534);
nand U11775 (N_11775,N_10281,N_10473);
nor U11776 (N_11776,N_10086,N_10570);
xnor U11777 (N_11777,N_10758,N_10955);
nand U11778 (N_11778,N_10640,N_10343);
or U11779 (N_11779,N_10322,N_10240);
nor U11780 (N_11780,N_10245,N_10655);
nor U11781 (N_11781,N_10123,N_10650);
or U11782 (N_11782,N_10543,N_10390);
nand U11783 (N_11783,N_10568,N_10861);
nor U11784 (N_11784,N_10166,N_10948);
xnor U11785 (N_11785,N_10725,N_10773);
nor U11786 (N_11786,N_10919,N_10762);
nand U11787 (N_11787,N_10088,N_10099);
and U11788 (N_11788,N_10882,N_10926);
and U11789 (N_11789,N_10795,N_10931);
nor U11790 (N_11790,N_10725,N_10292);
and U11791 (N_11791,N_10101,N_10243);
nand U11792 (N_11792,N_10890,N_10287);
nand U11793 (N_11793,N_10040,N_10928);
xnor U11794 (N_11794,N_10265,N_10841);
xor U11795 (N_11795,N_10783,N_10594);
or U11796 (N_11796,N_10366,N_10361);
and U11797 (N_11797,N_10621,N_10857);
nand U11798 (N_11798,N_10662,N_10364);
and U11799 (N_11799,N_10271,N_10767);
nor U11800 (N_11800,N_10502,N_10328);
and U11801 (N_11801,N_10726,N_10214);
and U11802 (N_11802,N_10757,N_10744);
or U11803 (N_11803,N_10059,N_10304);
and U11804 (N_11804,N_10302,N_10690);
and U11805 (N_11805,N_10876,N_10326);
or U11806 (N_11806,N_10889,N_10110);
or U11807 (N_11807,N_10546,N_10735);
nand U11808 (N_11808,N_10953,N_10158);
xnor U11809 (N_11809,N_10742,N_10360);
or U11810 (N_11810,N_10626,N_10822);
or U11811 (N_11811,N_10691,N_10586);
nand U11812 (N_11812,N_10437,N_10385);
nor U11813 (N_11813,N_10211,N_10803);
or U11814 (N_11814,N_10308,N_10601);
xnor U11815 (N_11815,N_10629,N_10301);
and U11816 (N_11816,N_10856,N_10983);
and U11817 (N_11817,N_10156,N_10369);
xor U11818 (N_11818,N_10931,N_10588);
or U11819 (N_11819,N_10503,N_10550);
or U11820 (N_11820,N_10247,N_10436);
or U11821 (N_11821,N_10856,N_10775);
nand U11822 (N_11822,N_10296,N_10788);
xor U11823 (N_11823,N_10486,N_10404);
or U11824 (N_11824,N_10749,N_10554);
and U11825 (N_11825,N_10085,N_10440);
xor U11826 (N_11826,N_10370,N_10447);
nor U11827 (N_11827,N_10463,N_10493);
and U11828 (N_11828,N_10934,N_10377);
and U11829 (N_11829,N_10901,N_10732);
xnor U11830 (N_11830,N_10674,N_10689);
xnor U11831 (N_11831,N_10745,N_10606);
nand U11832 (N_11832,N_10748,N_10396);
nor U11833 (N_11833,N_10956,N_10994);
xor U11834 (N_11834,N_10320,N_10454);
nor U11835 (N_11835,N_10224,N_10601);
nor U11836 (N_11836,N_10556,N_10376);
or U11837 (N_11837,N_10093,N_10070);
nand U11838 (N_11838,N_10940,N_10485);
or U11839 (N_11839,N_10680,N_10209);
xor U11840 (N_11840,N_10274,N_10414);
and U11841 (N_11841,N_10258,N_10552);
and U11842 (N_11842,N_10432,N_10396);
nor U11843 (N_11843,N_10888,N_10310);
and U11844 (N_11844,N_10705,N_10677);
nand U11845 (N_11845,N_10911,N_10085);
and U11846 (N_11846,N_10442,N_10370);
xnor U11847 (N_11847,N_10524,N_10613);
or U11848 (N_11848,N_10553,N_10766);
or U11849 (N_11849,N_10199,N_10899);
or U11850 (N_11850,N_10850,N_10878);
nand U11851 (N_11851,N_10633,N_10618);
nor U11852 (N_11852,N_10952,N_10970);
or U11853 (N_11853,N_10491,N_10602);
nor U11854 (N_11854,N_10530,N_10546);
xor U11855 (N_11855,N_10753,N_10624);
and U11856 (N_11856,N_10676,N_10934);
or U11857 (N_11857,N_10338,N_10815);
xor U11858 (N_11858,N_10337,N_10370);
nand U11859 (N_11859,N_10133,N_10694);
nor U11860 (N_11860,N_10069,N_10469);
or U11861 (N_11861,N_10535,N_10113);
xor U11862 (N_11862,N_10152,N_10196);
or U11863 (N_11863,N_10507,N_10326);
xor U11864 (N_11864,N_10001,N_10784);
and U11865 (N_11865,N_10788,N_10786);
and U11866 (N_11866,N_10886,N_10153);
and U11867 (N_11867,N_10641,N_10049);
nor U11868 (N_11868,N_10877,N_10718);
or U11869 (N_11869,N_10268,N_10677);
nor U11870 (N_11870,N_10431,N_10412);
or U11871 (N_11871,N_10756,N_10903);
xnor U11872 (N_11872,N_10138,N_10194);
nor U11873 (N_11873,N_10673,N_10806);
nand U11874 (N_11874,N_10286,N_10423);
or U11875 (N_11875,N_10125,N_10332);
or U11876 (N_11876,N_10670,N_10538);
or U11877 (N_11877,N_10029,N_10900);
or U11878 (N_11878,N_10930,N_10722);
xor U11879 (N_11879,N_10827,N_10633);
or U11880 (N_11880,N_10391,N_10245);
nand U11881 (N_11881,N_10358,N_10641);
nand U11882 (N_11882,N_10154,N_10838);
and U11883 (N_11883,N_10196,N_10051);
or U11884 (N_11884,N_10154,N_10935);
and U11885 (N_11885,N_10933,N_10311);
xnor U11886 (N_11886,N_10897,N_10878);
xnor U11887 (N_11887,N_10332,N_10758);
nand U11888 (N_11888,N_10135,N_10429);
or U11889 (N_11889,N_10796,N_10944);
nor U11890 (N_11890,N_10936,N_10858);
or U11891 (N_11891,N_10280,N_10882);
xor U11892 (N_11892,N_10933,N_10273);
nor U11893 (N_11893,N_10851,N_10786);
and U11894 (N_11894,N_10238,N_10428);
nand U11895 (N_11895,N_10326,N_10770);
and U11896 (N_11896,N_10713,N_10854);
or U11897 (N_11897,N_10997,N_10480);
xor U11898 (N_11898,N_10777,N_10129);
xnor U11899 (N_11899,N_10142,N_10728);
and U11900 (N_11900,N_10153,N_10712);
nor U11901 (N_11901,N_10929,N_10575);
nand U11902 (N_11902,N_10196,N_10649);
xnor U11903 (N_11903,N_10178,N_10593);
xnor U11904 (N_11904,N_10450,N_10313);
nand U11905 (N_11905,N_10386,N_10859);
and U11906 (N_11906,N_10288,N_10437);
and U11907 (N_11907,N_10522,N_10568);
or U11908 (N_11908,N_10841,N_10762);
nor U11909 (N_11909,N_10359,N_10880);
nand U11910 (N_11910,N_10459,N_10486);
xor U11911 (N_11911,N_10106,N_10599);
or U11912 (N_11912,N_10240,N_10095);
or U11913 (N_11913,N_10256,N_10971);
xnor U11914 (N_11914,N_10051,N_10984);
xor U11915 (N_11915,N_10601,N_10321);
xor U11916 (N_11916,N_10511,N_10421);
nor U11917 (N_11917,N_10798,N_10244);
xnor U11918 (N_11918,N_10914,N_10933);
nor U11919 (N_11919,N_10058,N_10491);
or U11920 (N_11920,N_10458,N_10753);
and U11921 (N_11921,N_10561,N_10886);
nand U11922 (N_11922,N_10310,N_10788);
nor U11923 (N_11923,N_10237,N_10860);
or U11924 (N_11924,N_10081,N_10212);
and U11925 (N_11925,N_10230,N_10298);
nor U11926 (N_11926,N_10852,N_10242);
and U11927 (N_11927,N_10703,N_10465);
nand U11928 (N_11928,N_10753,N_10674);
or U11929 (N_11929,N_10940,N_10043);
nand U11930 (N_11930,N_10209,N_10451);
and U11931 (N_11931,N_10978,N_10357);
nor U11932 (N_11932,N_10533,N_10272);
xor U11933 (N_11933,N_10476,N_10375);
or U11934 (N_11934,N_10238,N_10487);
and U11935 (N_11935,N_10803,N_10579);
nand U11936 (N_11936,N_10905,N_10765);
or U11937 (N_11937,N_10960,N_10810);
and U11938 (N_11938,N_10418,N_10231);
nand U11939 (N_11939,N_10443,N_10460);
nor U11940 (N_11940,N_10769,N_10949);
xor U11941 (N_11941,N_10632,N_10331);
xor U11942 (N_11942,N_10369,N_10611);
or U11943 (N_11943,N_10358,N_10860);
nand U11944 (N_11944,N_10417,N_10196);
or U11945 (N_11945,N_10479,N_10838);
and U11946 (N_11946,N_10751,N_10614);
nor U11947 (N_11947,N_10118,N_10968);
and U11948 (N_11948,N_10285,N_10007);
and U11949 (N_11949,N_10333,N_10928);
and U11950 (N_11950,N_10398,N_10536);
xnor U11951 (N_11951,N_10194,N_10009);
and U11952 (N_11952,N_10793,N_10696);
and U11953 (N_11953,N_10455,N_10656);
or U11954 (N_11954,N_10569,N_10325);
or U11955 (N_11955,N_10372,N_10115);
and U11956 (N_11956,N_10511,N_10215);
and U11957 (N_11957,N_10694,N_10122);
nand U11958 (N_11958,N_10429,N_10783);
and U11959 (N_11959,N_10737,N_10134);
or U11960 (N_11960,N_10849,N_10285);
and U11961 (N_11961,N_10084,N_10091);
nand U11962 (N_11962,N_10390,N_10421);
and U11963 (N_11963,N_10923,N_10069);
xor U11964 (N_11964,N_10074,N_10038);
nor U11965 (N_11965,N_10213,N_10247);
xnor U11966 (N_11966,N_10649,N_10572);
and U11967 (N_11967,N_10244,N_10591);
xor U11968 (N_11968,N_10952,N_10178);
nor U11969 (N_11969,N_10090,N_10791);
or U11970 (N_11970,N_10776,N_10903);
and U11971 (N_11971,N_10209,N_10149);
nor U11972 (N_11972,N_10174,N_10409);
and U11973 (N_11973,N_10526,N_10782);
nor U11974 (N_11974,N_10186,N_10394);
or U11975 (N_11975,N_10832,N_10996);
nor U11976 (N_11976,N_10121,N_10557);
and U11977 (N_11977,N_10441,N_10588);
or U11978 (N_11978,N_10873,N_10920);
nand U11979 (N_11979,N_10073,N_10768);
nor U11980 (N_11980,N_10869,N_10821);
nand U11981 (N_11981,N_10200,N_10042);
or U11982 (N_11982,N_10178,N_10514);
nand U11983 (N_11983,N_10522,N_10099);
nor U11984 (N_11984,N_10153,N_10782);
nor U11985 (N_11985,N_10744,N_10644);
nand U11986 (N_11986,N_10037,N_10953);
nor U11987 (N_11987,N_10801,N_10668);
xnor U11988 (N_11988,N_10257,N_10037);
or U11989 (N_11989,N_10467,N_10426);
nor U11990 (N_11990,N_10166,N_10171);
and U11991 (N_11991,N_10084,N_10727);
nor U11992 (N_11992,N_10409,N_10446);
nor U11993 (N_11993,N_10119,N_10191);
and U11994 (N_11994,N_10843,N_10671);
or U11995 (N_11995,N_10740,N_10101);
nor U11996 (N_11996,N_10014,N_10831);
or U11997 (N_11997,N_10345,N_10409);
nor U11998 (N_11998,N_10684,N_10373);
and U11999 (N_11999,N_10404,N_10901);
and U12000 (N_12000,N_11071,N_11441);
xor U12001 (N_12001,N_11721,N_11252);
nor U12002 (N_12002,N_11643,N_11970);
or U12003 (N_12003,N_11817,N_11410);
or U12004 (N_12004,N_11029,N_11450);
xnor U12005 (N_12005,N_11737,N_11820);
nand U12006 (N_12006,N_11086,N_11860);
nand U12007 (N_12007,N_11492,N_11982);
nand U12008 (N_12008,N_11113,N_11420);
or U12009 (N_12009,N_11364,N_11907);
xor U12010 (N_12010,N_11800,N_11581);
nor U12011 (N_12011,N_11514,N_11310);
nand U12012 (N_12012,N_11210,N_11749);
xnor U12013 (N_12013,N_11444,N_11783);
nor U12014 (N_12014,N_11690,N_11255);
nand U12015 (N_12015,N_11742,N_11774);
or U12016 (N_12016,N_11223,N_11657);
or U12017 (N_12017,N_11107,N_11259);
nor U12018 (N_12018,N_11767,N_11801);
or U12019 (N_12019,N_11173,N_11438);
and U12020 (N_12020,N_11597,N_11156);
nand U12021 (N_12021,N_11862,N_11031);
nand U12022 (N_12022,N_11475,N_11595);
nand U12023 (N_12023,N_11773,N_11389);
nand U12024 (N_12024,N_11286,N_11279);
nor U12025 (N_12025,N_11529,N_11530);
and U12026 (N_12026,N_11566,N_11160);
nand U12027 (N_12027,N_11798,N_11846);
nor U12028 (N_12028,N_11495,N_11466);
nor U12029 (N_12029,N_11004,N_11046);
nor U12030 (N_12030,N_11946,N_11732);
xnor U12031 (N_12031,N_11938,N_11047);
and U12032 (N_12032,N_11165,N_11283);
xor U12033 (N_12033,N_11250,N_11082);
nand U12034 (N_12034,N_11640,N_11261);
nor U12035 (N_12035,N_11207,N_11292);
xor U12036 (N_12036,N_11991,N_11873);
nor U12037 (N_12037,N_11952,N_11013);
xnor U12038 (N_12038,N_11079,N_11404);
nor U12039 (N_12039,N_11992,N_11848);
or U12040 (N_12040,N_11921,N_11758);
nor U12041 (N_12041,N_11795,N_11022);
nand U12042 (N_12042,N_11069,N_11367);
or U12043 (N_12043,N_11141,N_11018);
xnor U12044 (N_12044,N_11356,N_11414);
xor U12045 (N_12045,N_11028,N_11456);
xnor U12046 (N_12046,N_11186,N_11646);
and U12047 (N_12047,N_11620,N_11203);
nand U12048 (N_12048,N_11779,N_11053);
xor U12049 (N_12049,N_11890,N_11642);
nor U12050 (N_12050,N_11672,N_11975);
nor U12051 (N_12051,N_11519,N_11592);
nor U12052 (N_12052,N_11469,N_11666);
or U12053 (N_12053,N_11096,N_11854);
nand U12054 (N_12054,N_11139,N_11825);
xor U12055 (N_12055,N_11934,N_11927);
or U12056 (N_12056,N_11987,N_11818);
nand U12057 (N_12057,N_11338,N_11589);
and U12058 (N_12058,N_11370,N_11949);
nand U12059 (N_12059,N_11502,N_11813);
nand U12060 (N_12060,N_11211,N_11533);
nand U12061 (N_12061,N_11020,N_11346);
or U12062 (N_12062,N_11014,N_11659);
xor U12063 (N_12063,N_11948,N_11608);
xor U12064 (N_12064,N_11451,N_11521);
or U12065 (N_12065,N_11467,N_11781);
or U12066 (N_12066,N_11075,N_11163);
xnor U12067 (N_12067,N_11078,N_11696);
nor U12068 (N_12068,N_11751,N_11000);
nand U12069 (N_12069,N_11663,N_11169);
or U12070 (N_12070,N_11710,N_11049);
xor U12071 (N_12071,N_11081,N_11726);
and U12072 (N_12072,N_11723,N_11147);
and U12073 (N_12073,N_11912,N_11677);
xnor U12074 (N_12074,N_11043,N_11319);
xor U12075 (N_12075,N_11480,N_11145);
nand U12076 (N_12076,N_11740,N_11650);
or U12077 (N_12077,N_11164,N_11309);
nand U12078 (N_12078,N_11233,N_11808);
xnor U12079 (N_12079,N_11812,N_11264);
nor U12080 (N_12080,N_11586,N_11605);
or U12081 (N_12081,N_11419,N_11428);
or U12082 (N_12082,N_11962,N_11501);
xor U12083 (N_12083,N_11457,N_11702);
nor U12084 (N_12084,N_11357,N_11598);
and U12085 (N_12085,N_11509,N_11058);
nor U12086 (N_12086,N_11285,N_11562);
and U12087 (N_12087,N_11613,N_11228);
and U12088 (N_12088,N_11778,N_11603);
nor U12089 (N_12089,N_11709,N_11688);
or U12090 (N_12090,N_11877,N_11072);
nand U12091 (N_12091,N_11220,N_11988);
nand U12092 (N_12092,N_11615,N_11093);
and U12093 (N_12093,N_11254,N_11488);
or U12094 (N_12094,N_11601,N_11131);
or U12095 (N_12095,N_11746,N_11926);
nand U12096 (N_12096,N_11477,N_11833);
xor U12097 (N_12097,N_11504,N_11590);
or U12098 (N_12098,N_11656,N_11627);
nor U12099 (N_12099,N_11424,N_11231);
and U12100 (N_12100,N_11409,N_11771);
xnor U12101 (N_12101,N_11426,N_11112);
nor U12102 (N_12102,N_11070,N_11685);
and U12103 (N_12103,N_11077,N_11832);
and U12104 (N_12104,N_11528,N_11225);
and U12105 (N_12105,N_11911,N_11277);
or U12106 (N_12106,N_11236,N_11744);
and U12107 (N_12107,N_11258,N_11671);
and U12108 (N_12108,N_11960,N_11755);
or U12109 (N_12109,N_11101,N_11303);
or U12110 (N_12110,N_11632,N_11388);
nand U12111 (N_12111,N_11221,N_11700);
or U12112 (N_12112,N_11995,N_11161);
xnor U12113 (N_12113,N_11707,N_11397);
xor U12114 (N_12114,N_11675,N_11644);
xnor U12115 (N_12115,N_11994,N_11224);
nand U12116 (N_12116,N_11734,N_11212);
or U12117 (N_12117,N_11869,N_11799);
nand U12118 (N_12118,N_11035,N_11246);
nor U12119 (N_12119,N_11287,N_11323);
and U12120 (N_12120,N_11859,N_11454);
and U12121 (N_12121,N_11826,N_11447);
and U12122 (N_12122,N_11315,N_11340);
or U12123 (N_12123,N_11136,N_11146);
nor U12124 (N_12124,N_11684,N_11980);
and U12125 (N_12125,N_11312,N_11114);
nor U12126 (N_12126,N_11507,N_11193);
xnor U12127 (N_12127,N_11459,N_11120);
nor U12128 (N_12128,N_11554,N_11371);
xor U12129 (N_12129,N_11443,N_11032);
and U12130 (N_12130,N_11009,N_11302);
nand U12131 (N_12131,N_11669,N_11683);
and U12132 (N_12132,N_11856,N_11768);
and U12133 (N_12133,N_11490,N_11953);
xor U12134 (N_12134,N_11660,N_11494);
nor U12135 (N_12135,N_11919,N_11025);
and U12136 (N_12136,N_11850,N_11213);
and U12137 (N_12137,N_11940,N_11793);
nor U12138 (N_12138,N_11840,N_11133);
xor U12139 (N_12139,N_11652,N_11244);
or U12140 (N_12140,N_11928,N_11943);
nor U12141 (N_12141,N_11234,N_11347);
or U12142 (N_12142,N_11325,N_11378);
or U12143 (N_12143,N_11532,N_11068);
nor U12144 (N_12144,N_11753,N_11423);
nand U12145 (N_12145,N_11824,N_11416);
or U12146 (N_12146,N_11485,N_11355);
or U12147 (N_12147,N_11366,N_11117);
nand U12148 (N_12148,N_11422,N_11819);
nand U12149 (N_12149,N_11052,N_11587);
or U12150 (N_12150,N_11574,N_11321);
xor U12151 (N_12151,N_11008,N_11674);
and U12152 (N_12152,N_11573,N_11855);
nand U12153 (N_12153,N_11730,N_11332);
and U12154 (N_12154,N_11769,N_11089);
nand U12155 (N_12155,N_11406,N_11476);
and U12156 (N_12156,N_11522,N_11472);
nor U12157 (N_12157,N_11142,N_11654);
and U12158 (N_12158,N_11174,N_11331);
nand U12159 (N_12159,N_11864,N_11048);
and U12160 (N_12160,N_11026,N_11358);
xnor U12161 (N_12161,N_11513,N_11549);
nor U12162 (N_12162,N_11750,N_11842);
nor U12163 (N_12163,N_11963,N_11119);
or U12164 (N_12164,N_11874,N_11491);
or U12165 (N_12165,N_11373,N_11993);
nor U12166 (N_12166,N_11903,N_11922);
or U12167 (N_12167,N_11439,N_11568);
nor U12168 (N_12168,N_11508,N_11293);
nor U12169 (N_12169,N_11788,N_11350);
xor U12170 (N_12170,N_11839,N_11716);
and U12171 (N_12171,N_11636,N_11741);
nor U12172 (N_12172,N_11056,N_11074);
and U12173 (N_12173,N_11875,N_11230);
xor U12174 (N_12174,N_11455,N_11421);
and U12175 (N_12175,N_11628,N_11695);
xnor U12176 (N_12176,N_11841,N_11253);
nand U12177 (N_12177,N_11924,N_11239);
nor U12178 (N_12178,N_11761,N_11896);
or U12179 (N_12179,N_11094,N_11735);
nand U12180 (N_12180,N_11296,N_11999);
and U12181 (N_12181,N_11055,N_11904);
nor U12182 (N_12182,N_11204,N_11381);
nand U12183 (N_12183,N_11898,N_11481);
xor U12184 (N_12184,N_11852,N_11065);
and U12185 (N_12185,N_11238,N_11602);
or U12186 (N_12186,N_11973,N_11604);
nand U12187 (N_12187,N_11007,N_11941);
or U12188 (N_12188,N_11555,N_11205);
or U12189 (N_12189,N_11158,N_11470);
and U12190 (N_12190,N_11412,N_11775);
nor U12191 (N_12191,N_11437,N_11564);
or U12192 (N_12192,N_11442,N_11834);
nand U12193 (N_12193,N_11499,N_11436);
nand U12194 (N_12194,N_11757,N_11405);
and U12195 (N_12195,N_11823,N_11708);
or U12196 (N_12196,N_11351,N_11944);
nand U12197 (N_12197,N_11937,N_11914);
and U12198 (N_12198,N_11376,N_11967);
xnor U12199 (N_12199,N_11493,N_11929);
nor U12200 (N_12200,N_11128,N_11731);
xor U12201 (N_12201,N_11593,N_11104);
and U12202 (N_12202,N_11698,N_11301);
or U12203 (N_12203,N_11140,N_11092);
xor U12204 (N_12204,N_11809,N_11111);
and U12205 (N_12205,N_11900,N_11617);
and U12206 (N_12206,N_11237,N_11348);
and U12207 (N_12207,N_11282,N_11427);
xor U12208 (N_12208,N_11512,N_11118);
and U12209 (N_12209,N_11676,N_11951);
xnor U12210 (N_12210,N_11251,N_11167);
nor U12211 (N_12211,N_11541,N_11782);
or U12212 (N_12212,N_11382,N_11594);
xor U12213 (N_12213,N_11393,N_11317);
nor U12214 (N_12214,N_11059,N_11042);
xor U12215 (N_12215,N_11762,N_11106);
xor U12216 (N_12216,N_11016,N_11314);
xor U12217 (N_12217,N_11473,N_11027);
nand U12218 (N_12218,N_11387,N_11369);
xnor U12219 (N_12219,N_11484,N_11263);
nand U12220 (N_12220,N_11998,N_11330);
nand U12221 (N_12221,N_11242,N_11956);
nor U12222 (N_12222,N_11284,N_11905);
nand U12223 (N_12223,N_11226,N_11538);
or U12224 (N_12224,N_11379,N_11343);
nor U12225 (N_12225,N_11844,N_11085);
nand U12226 (N_12226,N_11445,N_11648);
xor U12227 (N_12227,N_11959,N_11634);
and U12228 (N_12228,N_11882,N_11308);
nand U12229 (N_12229,N_11712,N_11316);
or U12230 (N_12230,N_11720,N_11395);
and U12231 (N_12231,N_11784,N_11171);
xor U12232 (N_12232,N_11961,N_11958);
and U12233 (N_12233,N_11763,N_11127);
nor U12234 (N_12234,N_11184,N_11017);
nor U12235 (N_12235,N_11232,N_11516);
nand U12236 (N_12236,N_11638,N_11610);
nand U12237 (N_12237,N_11247,N_11327);
nor U12238 (N_12238,N_11827,N_11517);
xor U12239 (N_12239,N_11972,N_11468);
xnor U12240 (N_12240,N_11614,N_11265);
xor U12241 (N_12241,N_11354,N_11401);
or U12242 (N_12242,N_11828,N_11816);
nand U12243 (N_12243,N_11403,N_11334);
and U12244 (N_12244,N_11155,N_11913);
xor U12245 (N_12245,N_11197,N_11449);
and U12246 (N_12246,N_11429,N_11015);
nand U12247 (N_12247,N_11578,N_11333);
nor U12248 (N_12248,N_11130,N_11985);
or U12249 (N_12249,N_11374,N_11122);
nor U12250 (N_12250,N_11915,N_11010);
and U12251 (N_12251,N_11489,N_11372);
nand U12252 (N_12252,N_11157,N_11526);
and U12253 (N_12253,N_11872,N_11979);
nand U12254 (N_12254,N_11137,N_11545);
nand U12255 (N_12255,N_11288,N_11125);
and U12256 (N_12256,N_11881,N_11002);
xor U12257 (N_12257,N_11148,N_11706);
or U12258 (N_12258,N_11460,N_11486);
nand U12259 (N_12259,N_11363,N_11005);
nand U12260 (N_12260,N_11571,N_11425);
and U12261 (N_12261,N_11407,N_11630);
nor U12262 (N_12262,N_11728,N_11968);
and U12263 (N_12263,N_11889,N_11599);
and U12264 (N_12264,N_11715,N_11876);
xor U12265 (N_12265,N_11318,N_11668);
and U12266 (N_12266,N_11135,N_11273);
and U12267 (N_12267,N_11097,N_11479);
nand U12268 (N_12268,N_11083,N_11011);
and U12269 (N_12269,N_11849,N_11543);
nor U12270 (N_12270,N_11670,N_11150);
xnor U12271 (N_12271,N_11266,N_11458);
or U12272 (N_12272,N_11714,N_11006);
and U12273 (N_12273,N_11152,N_11548);
xor U12274 (N_12274,N_11129,N_11352);
xor U12275 (N_12275,N_11787,N_11531);
and U12276 (N_12276,N_11368,N_11899);
xor U12277 (N_12277,N_11192,N_11342);
xor U12278 (N_12278,N_11115,N_11766);
and U12279 (N_12279,N_11756,N_11618);
xor U12280 (N_12280,N_11123,N_11153);
nand U12281 (N_12281,N_11099,N_11391);
and U12282 (N_12282,N_11496,N_11645);
nand U12283 (N_12283,N_11084,N_11339);
nor U12284 (N_12284,N_11430,N_11159);
nor U12285 (N_12285,N_11177,N_11718);
or U12286 (N_12286,N_11815,N_11932);
xor U12287 (N_12287,N_11694,N_11465);
and U12288 (N_12288,N_11544,N_11188);
or U12289 (N_12289,N_11910,N_11474);
nand U12290 (N_12290,N_11754,N_11478);
or U12291 (N_12291,N_11229,N_11134);
nand U12292 (N_12292,N_11144,N_11747);
nand U12293 (N_12293,N_11736,N_11858);
or U12294 (N_12294,N_11066,N_11176);
or U12295 (N_12295,N_11448,N_11704);
nand U12296 (N_12296,N_11377,N_11933);
or U12297 (N_12297,N_11745,N_11743);
nand U12298 (N_12298,N_11966,N_11196);
xnor U12299 (N_12299,N_11579,N_11341);
xnor U12300 (N_12300,N_11390,N_11701);
xor U12301 (N_12301,N_11727,N_11981);
and U12302 (N_12302,N_11996,N_11440);
and U12303 (N_12303,N_11765,N_11322);
and U12304 (N_12304,N_11520,N_11691);
or U12305 (N_12305,N_11182,N_11785);
nand U12306 (N_12306,N_11661,N_11299);
or U12307 (N_12307,N_11971,N_11984);
or U12308 (N_12308,N_11076,N_11681);
nand U12309 (N_12309,N_11621,N_11845);
xor U12310 (N_12310,N_11415,N_11609);
and U12311 (N_12311,N_11777,N_11311);
or U12312 (N_12312,N_11344,N_11064);
xnor U12313 (N_12313,N_11651,N_11965);
nor U12314 (N_12314,N_11585,N_11090);
xnor U12315 (N_12315,N_11619,N_11281);
xor U12316 (N_12316,N_11471,N_11655);
nor U12317 (N_12317,N_11616,N_11664);
xnor U12318 (N_12318,N_11738,N_11417);
or U12319 (N_12319,N_11591,N_11584);
or U12320 (N_12320,N_11446,N_11611);
nand U12321 (N_12321,N_11256,N_11917);
nand U12322 (N_12322,N_11073,N_11957);
nor U12323 (N_12323,N_11091,N_11306);
nand U12324 (N_12324,N_11304,N_11558);
or U12325 (N_12325,N_11974,N_11892);
and U12326 (N_12326,N_11143,N_11262);
or U12327 (N_12327,N_11983,N_11300);
nor U12328 (N_12328,N_11969,N_11868);
or U12329 (N_12329,N_11780,N_11891);
nand U12330 (N_12330,N_11623,N_11853);
or U12331 (N_12331,N_11452,N_11271);
or U12332 (N_12332,N_11183,N_11977);
xor U12333 (N_12333,N_11362,N_11518);
or U12334 (N_12334,N_11087,N_11879);
xor U12335 (N_12335,N_11794,N_11198);
xnor U12336 (N_12336,N_11556,N_11003);
and U12337 (N_12337,N_11189,N_11375);
or U12338 (N_12338,N_11897,N_11653);
nor U12339 (N_12339,N_11673,N_11039);
or U12340 (N_12340,N_11553,N_11240);
nor U12341 (N_12341,N_11567,N_11641);
or U12342 (N_12342,N_11583,N_11515);
or U12343 (N_12343,N_11705,N_11209);
nand U12344 (N_12344,N_11699,N_11936);
and U12345 (N_12345,N_11098,N_11386);
nor U12346 (N_12346,N_11569,N_11510);
xnor U12347 (N_12347,N_11103,N_11108);
xnor U12348 (N_12348,N_11215,N_11976);
nor U12349 (N_12349,N_11267,N_11217);
nor U12350 (N_12350,N_11887,N_11249);
or U12351 (N_12351,N_11418,N_11525);
xor U12352 (N_12352,N_11733,N_11384);
nand U12353 (N_12353,N_11760,N_11649);
nor U12354 (N_12354,N_11622,N_11606);
and U12355 (N_12355,N_11878,N_11829);
and U12356 (N_12356,N_11194,N_11639);
and U12357 (N_12357,N_11222,N_11863);
and U12358 (N_12358,N_11739,N_11637);
nor U12359 (N_12359,N_11682,N_11550);
xor U12360 (N_12360,N_11866,N_11524);
nand U12361 (N_12361,N_11180,N_11885);
and U12362 (N_12362,N_11539,N_11294);
and U12363 (N_12363,N_11206,N_11320);
and U12364 (N_12364,N_11770,N_11433);
nand U12365 (N_12365,N_11811,N_11792);
nand U12366 (N_12366,N_11498,N_11202);
nor U12367 (N_12367,N_11274,N_11551);
or U12368 (N_12368,N_11324,N_11270);
xor U12369 (N_12369,N_11132,N_11200);
or U12370 (N_12370,N_11124,N_11764);
xnor U12371 (N_12371,N_11797,N_11349);
xor U12372 (N_12372,N_11001,N_11038);
nand U12373 (N_12373,N_11665,N_11464);
nor U12374 (N_12374,N_11463,N_11930);
or U12375 (N_12375,N_11431,N_11275);
nand U12376 (N_12376,N_11462,N_11523);
and U12377 (N_12377,N_11034,N_11298);
xnor U12378 (N_12378,N_11552,N_11278);
or U12379 (N_12379,N_11235,N_11686);
and U12380 (N_12380,N_11810,N_11804);
nor U12381 (N_12381,N_11759,N_11580);
nor U12382 (N_12382,N_11453,N_11088);
nor U12383 (N_12383,N_11483,N_11057);
or U12384 (N_12384,N_11260,N_11893);
xnor U12385 (N_12385,N_11612,N_11729);
nor U12386 (N_12386,N_11280,N_11191);
and U12387 (N_12387,N_11776,N_11434);
nand U12388 (N_12388,N_11990,N_11162);
xnor U12389 (N_12389,N_11679,N_11385);
nor U12390 (N_12390,N_11095,N_11843);
and U12391 (N_12391,N_11717,N_11693);
or U12392 (N_12392,N_11527,N_11045);
nor U12393 (N_12393,N_11432,N_11631);
or U12394 (N_12394,N_11772,N_11208);
or U12395 (N_12395,N_11337,N_11536);
nand U12396 (N_12396,N_11506,N_11557);
nand U12397 (N_12397,N_11154,N_11080);
nand U12398 (N_12398,N_11019,N_11178);
and U12399 (N_12399,N_11870,N_11044);
nand U12400 (N_12400,N_11786,N_11021);
nor U12401 (N_12401,N_11942,N_11577);
nand U12402 (N_12402,N_11814,N_11269);
or U12403 (N_12403,N_11884,N_11396);
nor U12404 (N_12404,N_11713,N_11647);
or U12405 (N_12405,N_11487,N_11678);
nor U12406 (N_12406,N_11600,N_11964);
xnor U12407 (N_12407,N_11170,N_11201);
xor U12408 (N_12408,N_11790,N_11109);
xor U12409 (N_12409,N_11116,N_11181);
or U12410 (N_12410,N_11482,N_11245);
and U12411 (N_12411,N_11110,N_11172);
nor U12412 (N_12412,N_11326,N_11138);
and U12413 (N_12413,N_11955,N_11289);
nor U12414 (N_12414,N_11680,N_11305);
and U12415 (N_12415,N_11805,N_11168);
nand U12416 (N_12416,N_11361,N_11945);
nand U12417 (N_12417,N_11796,N_11625);
or U12418 (N_12418,N_11947,N_11692);
nand U12419 (N_12419,N_11313,N_11497);
xor U12420 (N_12420,N_11883,N_11121);
and U12421 (N_12421,N_11307,N_11923);
or U12422 (N_12422,N_11540,N_11175);
nor U12423 (N_12423,N_11040,N_11821);
or U12424 (N_12424,N_11335,N_11689);
or U12425 (N_12425,N_11561,N_11570);
nand U12426 (N_12426,N_11791,N_11576);
xor U12427 (N_12427,N_11328,N_11582);
nand U12428 (N_12428,N_11803,N_11986);
and U12429 (N_12429,N_11394,N_11997);
xor U12430 (N_12430,N_11888,N_11916);
nor U12431 (N_12431,N_11752,N_11719);
nand U12432 (N_12432,N_11037,N_11257);
and U12433 (N_12433,N_11703,N_11906);
and U12434 (N_12434,N_11575,N_11500);
nand U12435 (N_12435,N_11607,N_11711);
xor U12436 (N_12436,N_11051,N_11241);
or U12437 (N_12437,N_11216,N_11272);
and U12438 (N_12438,N_11836,N_11297);
nand U12439 (N_12439,N_11830,N_11725);
nand U12440 (N_12440,N_11151,N_11100);
xnor U12441 (N_12441,N_11291,N_11511);
nor U12442 (N_12442,N_11435,N_11925);
xor U12443 (N_12443,N_11054,N_11149);
xnor U12444 (N_12444,N_11629,N_11935);
nor U12445 (N_12445,N_11722,N_11248);
and U12446 (N_12446,N_11534,N_11023);
xnor U12447 (N_12447,N_11662,N_11067);
xor U12448 (N_12448,N_11360,N_11806);
nand U12449 (N_12449,N_11954,N_11380);
nand U12450 (N_12450,N_11041,N_11989);
xnor U12451 (N_12451,N_11918,N_11886);
xor U12452 (N_12452,N_11748,N_11847);
nand U12453 (N_12453,N_11398,N_11353);
or U12454 (N_12454,N_11822,N_11894);
and U12455 (N_12455,N_11542,N_11588);
or U12456 (N_12456,N_11030,N_11295);
or U12457 (N_12457,N_11195,N_11939);
nor U12458 (N_12458,N_11802,N_11199);
or U12459 (N_12459,N_11413,N_11461);
and U12460 (N_12460,N_11724,N_11851);
or U12461 (N_12461,N_11909,N_11187);
xnor U12462 (N_12462,N_11880,N_11871);
nand U12463 (N_12463,N_11102,N_11667);
xnor U12464 (N_12464,N_11895,N_11179);
and U12465 (N_12465,N_11902,N_11276);
and U12466 (N_12466,N_11063,N_11061);
xor U12467 (N_12467,N_11624,N_11978);
and U12468 (N_12468,N_11565,N_11336);
and U12469 (N_12469,N_11359,N_11901);
nand U12470 (N_12470,N_11857,N_11033);
and U12471 (N_12471,N_11062,N_11329);
or U12472 (N_12472,N_11290,N_11867);
nand U12473 (N_12473,N_11626,N_11503);
or U12474 (N_12474,N_11920,N_11547);
nand U12475 (N_12475,N_11535,N_11635);
and U12476 (N_12476,N_11012,N_11227);
xor U12477 (N_12477,N_11658,N_11835);
and U12478 (N_12478,N_11190,N_11908);
xor U12479 (N_12479,N_11861,N_11505);
nand U12480 (N_12480,N_11036,N_11837);
and U12481 (N_12481,N_11383,N_11365);
xnor U12482 (N_12482,N_11789,N_11399);
xnor U12483 (N_12483,N_11392,N_11563);
xor U12484 (N_12484,N_11214,N_11697);
nand U12485 (N_12485,N_11105,N_11402);
nor U12486 (N_12486,N_11950,N_11838);
nand U12487 (N_12487,N_11596,N_11345);
nand U12488 (N_12488,N_11060,N_11218);
nand U12489 (N_12489,N_11408,N_11865);
nand U12490 (N_12490,N_11546,N_11024);
or U12491 (N_12491,N_11126,N_11807);
xor U12492 (N_12492,N_11166,N_11687);
nor U12493 (N_12493,N_11400,N_11560);
nand U12494 (N_12494,N_11572,N_11243);
xnor U12495 (N_12495,N_11559,N_11185);
or U12496 (N_12496,N_11411,N_11268);
nand U12497 (N_12497,N_11219,N_11633);
nor U12498 (N_12498,N_11931,N_11537);
and U12499 (N_12499,N_11831,N_11050);
nor U12500 (N_12500,N_11164,N_11910);
nor U12501 (N_12501,N_11036,N_11712);
and U12502 (N_12502,N_11007,N_11719);
nand U12503 (N_12503,N_11778,N_11654);
or U12504 (N_12504,N_11026,N_11495);
xor U12505 (N_12505,N_11053,N_11197);
xnor U12506 (N_12506,N_11405,N_11340);
and U12507 (N_12507,N_11367,N_11997);
and U12508 (N_12508,N_11740,N_11561);
nand U12509 (N_12509,N_11468,N_11949);
nand U12510 (N_12510,N_11396,N_11373);
nand U12511 (N_12511,N_11949,N_11323);
nor U12512 (N_12512,N_11522,N_11984);
xor U12513 (N_12513,N_11822,N_11221);
nand U12514 (N_12514,N_11066,N_11776);
and U12515 (N_12515,N_11691,N_11185);
nand U12516 (N_12516,N_11210,N_11242);
xnor U12517 (N_12517,N_11936,N_11735);
xnor U12518 (N_12518,N_11394,N_11732);
nor U12519 (N_12519,N_11272,N_11798);
nor U12520 (N_12520,N_11750,N_11101);
nand U12521 (N_12521,N_11510,N_11088);
and U12522 (N_12522,N_11665,N_11273);
nor U12523 (N_12523,N_11922,N_11445);
nand U12524 (N_12524,N_11709,N_11369);
xnor U12525 (N_12525,N_11684,N_11473);
nor U12526 (N_12526,N_11660,N_11613);
or U12527 (N_12527,N_11364,N_11416);
nand U12528 (N_12528,N_11285,N_11517);
and U12529 (N_12529,N_11578,N_11817);
nand U12530 (N_12530,N_11415,N_11632);
and U12531 (N_12531,N_11871,N_11238);
nor U12532 (N_12532,N_11054,N_11423);
or U12533 (N_12533,N_11490,N_11907);
and U12534 (N_12534,N_11174,N_11253);
nand U12535 (N_12535,N_11868,N_11741);
xor U12536 (N_12536,N_11351,N_11430);
xnor U12537 (N_12537,N_11060,N_11628);
xor U12538 (N_12538,N_11433,N_11118);
xor U12539 (N_12539,N_11032,N_11688);
nand U12540 (N_12540,N_11903,N_11192);
or U12541 (N_12541,N_11145,N_11140);
or U12542 (N_12542,N_11621,N_11462);
and U12543 (N_12543,N_11719,N_11296);
nand U12544 (N_12544,N_11868,N_11624);
xor U12545 (N_12545,N_11374,N_11824);
nand U12546 (N_12546,N_11215,N_11327);
nand U12547 (N_12547,N_11948,N_11883);
or U12548 (N_12548,N_11364,N_11818);
xor U12549 (N_12549,N_11011,N_11731);
xor U12550 (N_12550,N_11604,N_11030);
nand U12551 (N_12551,N_11154,N_11111);
or U12552 (N_12552,N_11946,N_11344);
nor U12553 (N_12553,N_11566,N_11129);
or U12554 (N_12554,N_11812,N_11876);
and U12555 (N_12555,N_11016,N_11511);
nor U12556 (N_12556,N_11304,N_11862);
and U12557 (N_12557,N_11598,N_11789);
or U12558 (N_12558,N_11670,N_11172);
nand U12559 (N_12559,N_11147,N_11515);
or U12560 (N_12560,N_11214,N_11499);
nand U12561 (N_12561,N_11877,N_11922);
xnor U12562 (N_12562,N_11765,N_11030);
nand U12563 (N_12563,N_11053,N_11495);
nor U12564 (N_12564,N_11645,N_11700);
xor U12565 (N_12565,N_11516,N_11536);
xnor U12566 (N_12566,N_11413,N_11379);
and U12567 (N_12567,N_11067,N_11408);
and U12568 (N_12568,N_11460,N_11069);
or U12569 (N_12569,N_11949,N_11372);
nand U12570 (N_12570,N_11530,N_11331);
xnor U12571 (N_12571,N_11872,N_11571);
or U12572 (N_12572,N_11764,N_11013);
nor U12573 (N_12573,N_11836,N_11197);
nor U12574 (N_12574,N_11212,N_11808);
or U12575 (N_12575,N_11088,N_11701);
or U12576 (N_12576,N_11566,N_11903);
nand U12577 (N_12577,N_11020,N_11878);
or U12578 (N_12578,N_11972,N_11030);
xnor U12579 (N_12579,N_11664,N_11148);
nor U12580 (N_12580,N_11329,N_11310);
or U12581 (N_12581,N_11518,N_11655);
xor U12582 (N_12582,N_11253,N_11099);
or U12583 (N_12583,N_11796,N_11507);
xnor U12584 (N_12584,N_11477,N_11575);
nand U12585 (N_12585,N_11703,N_11942);
nand U12586 (N_12586,N_11731,N_11013);
and U12587 (N_12587,N_11653,N_11661);
nor U12588 (N_12588,N_11710,N_11006);
or U12589 (N_12589,N_11877,N_11096);
and U12590 (N_12590,N_11926,N_11032);
nand U12591 (N_12591,N_11251,N_11159);
xnor U12592 (N_12592,N_11548,N_11185);
nand U12593 (N_12593,N_11354,N_11006);
nor U12594 (N_12594,N_11757,N_11577);
nand U12595 (N_12595,N_11632,N_11826);
xor U12596 (N_12596,N_11225,N_11675);
and U12597 (N_12597,N_11632,N_11304);
or U12598 (N_12598,N_11791,N_11059);
nand U12599 (N_12599,N_11595,N_11757);
or U12600 (N_12600,N_11096,N_11112);
nand U12601 (N_12601,N_11381,N_11348);
xnor U12602 (N_12602,N_11026,N_11157);
or U12603 (N_12603,N_11438,N_11287);
or U12604 (N_12604,N_11705,N_11528);
nor U12605 (N_12605,N_11706,N_11640);
nand U12606 (N_12606,N_11179,N_11566);
and U12607 (N_12607,N_11180,N_11473);
xnor U12608 (N_12608,N_11512,N_11580);
xor U12609 (N_12609,N_11795,N_11945);
nor U12610 (N_12610,N_11075,N_11788);
xnor U12611 (N_12611,N_11142,N_11148);
and U12612 (N_12612,N_11816,N_11615);
nor U12613 (N_12613,N_11259,N_11757);
and U12614 (N_12614,N_11169,N_11494);
or U12615 (N_12615,N_11337,N_11837);
or U12616 (N_12616,N_11300,N_11302);
xnor U12617 (N_12617,N_11194,N_11551);
nor U12618 (N_12618,N_11428,N_11534);
xor U12619 (N_12619,N_11138,N_11523);
and U12620 (N_12620,N_11539,N_11130);
and U12621 (N_12621,N_11604,N_11850);
xor U12622 (N_12622,N_11364,N_11606);
or U12623 (N_12623,N_11811,N_11374);
nand U12624 (N_12624,N_11607,N_11493);
or U12625 (N_12625,N_11013,N_11060);
or U12626 (N_12626,N_11319,N_11706);
or U12627 (N_12627,N_11374,N_11737);
or U12628 (N_12628,N_11787,N_11902);
nor U12629 (N_12629,N_11745,N_11139);
and U12630 (N_12630,N_11806,N_11540);
xnor U12631 (N_12631,N_11067,N_11816);
nor U12632 (N_12632,N_11129,N_11107);
and U12633 (N_12633,N_11676,N_11973);
and U12634 (N_12634,N_11662,N_11240);
and U12635 (N_12635,N_11053,N_11383);
xor U12636 (N_12636,N_11030,N_11609);
xor U12637 (N_12637,N_11211,N_11382);
nand U12638 (N_12638,N_11010,N_11956);
xor U12639 (N_12639,N_11854,N_11878);
nand U12640 (N_12640,N_11620,N_11438);
or U12641 (N_12641,N_11373,N_11268);
or U12642 (N_12642,N_11795,N_11875);
or U12643 (N_12643,N_11889,N_11977);
xor U12644 (N_12644,N_11329,N_11671);
nor U12645 (N_12645,N_11428,N_11696);
nand U12646 (N_12646,N_11957,N_11600);
nor U12647 (N_12647,N_11435,N_11454);
xnor U12648 (N_12648,N_11363,N_11287);
nor U12649 (N_12649,N_11387,N_11249);
and U12650 (N_12650,N_11221,N_11782);
or U12651 (N_12651,N_11836,N_11360);
and U12652 (N_12652,N_11256,N_11403);
nand U12653 (N_12653,N_11431,N_11727);
or U12654 (N_12654,N_11132,N_11103);
or U12655 (N_12655,N_11716,N_11325);
nand U12656 (N_12656,N_11310,N_11581);
and U12657 (N_12657,N_11576,N_11008);
nor U12658 (N_12658,N_11010,N_11382);
xnor U12659 (N_12659,N_11592,N_11103);
nand U12660 (N_12660,N_11179,N_11579);
and U12661 (N_12661,N_11479,N_11633);
or U12662 (N_12662,N_11915,N_11357);
nand U12663 (N_12663,N_11965,N_11810);
or U12664 (N_12664,N_11824,N_11550);
nor U12665 (N_12665,N_11714,N_11032);
nor U12666 (N_12666,N_11572,N_11173);
xnor U12667 (N_12667,N_11804,N_11140);
nand U12668 (N_12668,N_11766,N_11397);
nand U12669 (N_12669,N_11774,N_11655);
nand U12670 (N_12670,N_11731,N_11421);
or U12671 (N_12671,N_11808,N_11881);
or U12672 (N_12672,N_11921,N_11945);
or U12673 (N_12673,N_11997,N_11007);
nand U12674 (N_12674,N_11602,N_11295);
xor U12675 (N_12675,N_11503,N_11825);
and U12676 (N_12676,N_11008,N_11301);
nor U12677 (N_12677,N_11515,N_11135);
nor U12678 (N_12678,N_11241,N_11313);
and U12679 (N_12679,N_11308,N_11584);
nand U12680 (N_12680,N_11230,N_11423);
and U12681 (N_12681,N_11310,N_11742);
and U12682 (N_12682,N_11017,N_11113);
and U12683 (N_12683,N_11150,N_11216);
or U12684 (N_12684,N_11835,N_11384);
and U12685 (N_12685,N_11993,N_11871);
or U12686 (N_12686,N_11753,N_11576);
xor U12687 (N_12687,N_11276,N_11454);
nand U12688 (N_12688,N_11743,N_11963);
nor U12689 (N_12689,N_11573,N_11323);
and U12690 (N_12690,N_11563,N_11633);
xnor U12691 (N_12691,N_11322,N_11313);
or U12692 (N_12692,N_11329,N_11642);
nand U12693 (N_12693,N_11256,N_11916);
xnor U12694 (N_12694,N_11191,N_11062);
xor U12695 (N_12695,N_11551,N_11076);
nand U12696 (N_12696,N_11694,N_11741);
or U12697 (N_12697,N_11402,N_11320);
or U12698 (N_12698,N_11749,N_11332);
xor U12699 (N_12699,N_11853,N_11450);
nor U12700 (N_12700,N_11442,N_11357);
nor U12701 (N_12701,N_11059,N_11803);
nor U12702 (N_12702,N_11424,N_11726);
and U12703 (N_12703,N_11842,N_11758);
nand U12704 (N_12704,N_11417,N_11419);
nor U12705 (N_12705,N_11267,N_11786);
and U12706 (N_12706,N_11523,N_11693);
or U12707 (N_12707,N_11513,N_11027);
and U12708 (N_12708,N_11174,N_11970);
xor U12709 (N_12709,N_11686,N_11975);
xor U12710 (N_12710,N_11421,N_11309);
xor U12711 (N_12711,N_11363,N_11060);
nor U12712 (N_12712,N_11628,N_11098);
xnor U12713 (N_12713,N_11554,N_11961);
xnor U12714 (N_12714,N_11860,N_11250);
or U12715 (N_12715,N_11770,N_11398);
nor U12716 (N_12716,N_11856,N_11211);
xnor U12717 (N_12717,N_11864,N_11428);
and U12718 (N_12718,N_11777,N_11438);
and U12719 (N_12719,N_11216,N_11960);
nor U12720 (N_12720,N_11484,N_11258);
nor U12721 (N_12721,N_11695,N_11594);
nor U12722 (N_12722,N_11958,N_11145);
or U12723 (N_12723,N_11699,N_11325);
xor U12724 (N_12724,N_11678,N_11453);
xnor U12725 (N_12725,N_11869,N_11240);
xor U12726 (N_12726,N_11834,N_11994);
or U12727 (N_12727,N_11520,N_11029);
or U12728 (N_12728,N_11591,N_11653);
or U12729 (N_12729,N_11631,N_11238);
nand U12730 (N_12730,N_11480,N_11194);
or U12731 (N_12731,N_11827,N_11730);
xor U12732 (N_12732,N_11594,N_11189);
or U12733 (N_12733,N_11870,N_11111);
nor U12734 (N_12734,N_11285,N_11811);
nand U12735 (N_12735,N_11345,N_11492);
or U12736 (N_12736,N_11633,N_11138);
or U12737 (N_12737,N_11324,N_11026);
nand U12738 (N_12738,N_11299,N_11219);
nand U12739 (N_12739,N_11324,N_11284);
nand U12740 (N_12740,N_11529,N_11458);
xor U12741 (N_12741,N_11725,N_11804);
nor U12742 (N_12742,N_11916,N_11220);
or U12743 (N_12743,N_11655,N_11202);
or U12744 (N_12744,N_11444,N_11240);
or U12745 (N_12745,N_11676,N_11330);
xnor U12746 (N_12746,N_11416,N_11660);
and U12747 (N_12747,N_11941,N_11279);
xnor U12748 (N_12748,N_11783,N_11959);
and U12749 (N_12749,N_11417,N_11518);
xor U12750 (N_12750,N_11395,N_11003);
xor U12751 (N_12751,N_11750,N_11922);
nor U12752 (N_12752,N_11057,N_11313);
or U12753 (N_12753,N_11097,N_11462);
or U12754 (N_12754,N_11330,N_11264);
nand U12755 (N_12755,N_11582,N_11300);
xor U12756 (N_12756,N_11624,N_11269);
nand U12757 (N_12757,N_11401,N_11266);
xor U12758 (N_12758,N_11975,N_11903);
xor U12759 (N_12759,N_11920,N_11691);
nor U12760 (N_12760,N_11848,N_11220);
xor U12761 (N_12761,N_11428,N_11307);
and U12762 (N_12762,N_11801,N_11089);
or U12763 (N_12763,N_11030,N_11587);
or U12764 (N_12764,N_11714,N_11058);
xor U12765 (N_12765,N_11318,N_11615);
or U12766 (N_12766,N_11058,N_11410);
nor U12767 (N_12767,N_11354,N_11229);
nor U12768 (N_12768,N_11552,N_11762);
nand U12769 (N_12769,N_11450,N_11286);
nand U12770 (N_12770,N_11393,N_11770);
or U12771 (N_12771,N_11199,N_11777);
nor U12772 (N_12772,N_11372,N_11685);
or U12773 (N_12773,N_11073,N_11022);
nor U12774 (N_12774,N_11097,N_11093);
nand U12775 (N_12775,N_11882,N_11416);
and U12776 (N_12776,N_11128,N_11038);
nand U12777 (N_12777,N_11586,N_11809);
and U12778 (N_12778,N_11402,N_11596);
xor U12779 (N_12779,N_11260,N_11594);
or U12780 (N_12780,N_11190,N_11563);
xor U12781 (N_12781,N_11821,N_11335);
nand U12782 (N_12782,N_11990,N_11404);
nand U12783 (N_12783,N_11263,N_11121);
and U12784 (N_12784,N_11722,N_11280);
xor U12785 (N_12785,N_11365,N_11764);
nand U12786 (N_12786,N_11624,N_11503);
and U12787 (N_12787,N_11177,N_11581);
nand U12788 (N_12788,N_11307,N_11715);
xnor U12789 (N_12789,N_11371,N_11070);
nand U12790 (N_12790,N_11447,N_11098);
or U12791 (N_12791,N_11455,N_11616);
xnor U12792 (N_12792,N_11834,N_11246);
or U12793 (N_12793,N_11498,N_11780);
and U12794 (N_12794,N_11152,N_11552);
or U12795 (N_12795,N_11272,N_11689);
nor U12796 (N_12796,N_11194,N_11635);
and U12797 (N_12797,N_11055,N_11724);
xor U12798 (N_12798,N_11341,N_11756);
xor U12799 (N_12799,N_11002,N_11047);
xnor U12800 (N_12800,N_11388,N_11541);
and U12801 (N_12801,N_11624,N_11165);
and U12802 (N_12802,N_11165,N_11356);
xnor U12803 (N_12803,N_11498,N_11723);
or U12804 (N_12804,N_11599,N_11746);
nand U12805 (N_12805,N_11491,N_11887);
xnor U12806 (N_12806,N_11945,N_11053);
nor U12807 (N_12807,N_11150,N_11699);
and U12808 (N_12808,N_11260,N_11067);
nor U12809 (N_12809,N_11230,N_11705);
or U12810 (N_12810,N_11539,N_11837);
nand U12811 (N_12811,N_11535,N_11966);
nand U12812 (N_12812,N_11660,N_11814);
or U12813 (N_12813,N_11138,N_11752);
and U12814 (N_12814,N_11399,N_11424);
nor U12815 (N_12815,N_11831,N_11357);
nor U12816 (N_12816,N_11164,N_11951);
nand U12817 (N_12817,N_11466,N_11479);
or U12818 (N_12818,N_11419,N_11677);
nand U12819 (N_12819,N_11536,N_11844);
nor U12820 (N_12820,N_11950,N_11002);
or U12821 (N_12821,N_11510,N_11634);
nand U12822 (N_12822,N_11714,N_11077);
xor U12823 (N_12823,N_11171,N_11403);
and U12824 (N_12824,N_11845,N_11810);
nor U12825 (N_12825,N_11568,N_11863);
xor U12826 (N_12826,N_11832,N_11023);
nand U12827 (N_12827,N_11004,N_11190);
or U12828 (N_12828,N_11084,N_11344);
nor U12829 (N_12829,N_11430,N_11929);
and U12830 (N_12830,N_11646,N_11060);
xnor U12831 (N_12831,N_11818,N_11113);
or U12832 (N_12832,N_11961,N_11046);
nand U12833 (N_12833,N_11914,N_11338);
or U12834 (N_12834,N_11925,N_11554);
or U12835 (N_12835,N_11425,N_11560);
nor U12836 (N_12836,N_11306,N_11622);
xnor U12837 (N_12837,N_11670,N_11626);
and U12838 (N_12838,N_11521,N_11582);
or U12839 (N_12839,N_11331,N_11649);
and U12840 (N_12840,N_11775,N_11639);
or U12841 (N_12841,N_11471,N_11934);
or U12842 (N_12842,N_11088,N_11753);
and U12843 (N_12843,N_11179,N_11147);
nor U12844 (N_12844,N_11348,N_11719);
nor U12845 (N_12845,N_11198,N_11664);
nand U12846 (N_12846,N_11160,N_11979);
xor U12847 (N_12847,N_11867,N_11546);
xor U12848 (N_12848,N_11766,N_11373);
xor U12849 (N_12849,N_11784,N_11760);
or U12850 (N_12850,N_11978,N_11540);
nand U12851 (N_12851,N_11210,N_11557);
or U12852 (N_12852,N_11676,N_11887);
and U12853 (N_12853,N_11596,N_11394);
nand U12854 (N_12854,N_11740,N_11194);
nor U12855 (N_12855,N_11389,N_11783);
and U12856 (N_12856,N_11172,N_11566);
nand U12857 (N_12857,N_11811,N_11307);
or U12858 (N_12858,N_11966,N_11754);
or U12859 (N_12859,N_11776,N_11656);
or U12860 (N_12860,N_11950,N_11598);
or U12861 (N_12861,N_11917,N_11984);
xnor U12862 (N_12862,N_11564,N_11307);
nor U12863 (N_12863,N_11842,N_11314);
xor U12864 (N_12864,N_11826,N_11932);
xor U12865 (N_12865,N_11134,N_11009);
nand U12866 (N_12866,N_11617,N_11677);
or U12867 (N_12867,N_11326,N_11406);
or U12868 (N_12868,N_11328,N_11823);
nand U12869 (N_12869,N_11652,N_11788);
xnor U12870 (N_12870,N_11761,N_11533);
and U12871 (N_12871,N_11954,N_11699);
nor U12872 (N_12872,N_11462,N_11456);
nand U12873 (N_12873,N_11874,N_11324);
nor U12874 (N_12874,N_11181,N_11236);
xnor U12875 (N_12875,N_11912,N_11361);
or U12876 (N_12876,N_11899,N_11621);
or U12877 (N_12877,N_11120,N_11863);
and U12878 (N_12878,N_11288,N_11413);
nand U12879 (N_12879,N_11176,N_11061);
or U12880 (N_12880,N_11954,N_11011);
or U12881 (N_12881,N_11133,N_11124);
and U12882 (N_12882,N_11417,N_11190);
xnor U12883 (N_12883,N_11367,N_11204);
nand U12884 (N_12884,N_11243,N_11613);
or U12885 (N_12885,N_11856,N_11958);
or U12886 (N_12886,N_11776,N_11144);
nor U12887 (N_12887,N_11993,N_11628);
xnor U12888 (N_12888,N_11754,N_11544);
nor U12889 (N_12889,N_11510,N_11788);
and U12890 (N_12890,N_11341,N_11167);
nand U12891 (N_12891,N_11831,N_11306);
and U12892 (N_12892,N_11851,N_11385);
and U12893 (N_12893,N_11263,N_11156);
and U12894 (N_12894,N_11536,N_11576);
or U12895 (N_12895,N_11450,N_11225);
nor U12896 (N_12896,N_11564,N_11462);
nand U12897 (N_12897,N_11298,N_11257);
and U12898 (N_12898,N_11958,N_11848);
nor U12899 (N_12899,N_11197,N_11725);
nor U12900 (N_12900,N_11183,N_11454);
or U12901 (N_12901,N_11754,N_11811);
and U12902 (N_12902,N_11161,N_11141);
or U12903 (N_12903,N_11865,N_11129);
or U12904 (N_12904,N_11677,N_11073);
and U12905 (N_12905,N_11125,N_11117);
xnor U12906 (N_12906,N_11316,N_11941);
nor U12907 (N_12907,N_11618,N_11641);
or U12908 (N_12908,N_11337,N_11556);
xor U12909 (N_12909,N_11708,N_11990);
nor U12910 (N_12910,N_11825,N_11851);
nand U12911 (N_12911,N_11972,N_11714);
nand U12912 (N_12912,N_11320,N_11689);
xnor U12913 (N_12913,N_11772,N_11757);
and U12914 (N_12914,N_11046,N_11363);
xor U12915 (N_12915,N_11995,N_11654);
nor U12916 (N_12916,N_11400,N_11350);
and U12917 (N_12917,N_11560,N_11655);
nand U12918 (N_12918,N_11266,N_11172);
xnor U12919 (N_12919,N_11220,N_11120);
nor U12920 (N_12920,N_11821,N_11855);
xnor U12921 (N_12921,N_11904,N_11723);
xor U12922 (N_12922,N_11280,N_11847);
xor U12923 (N_12923,N_11553,N_11290);
or U12924 (N_12924,N_11161,N_11803);
xor U12925 (N_12925,N_11329,N_11087);
nor U12926 (N_12926,N_11550,N_11500);
xnor U12927 (N_12927,N_11516,N_11412);
xnor U12928 (N_12928,N_11459,N_11753);
nand U12929 (N_12929,N_11896,N_11174);
or U12930 (N_12930,N_11503,N_11995);
xnor U12931 (N_12931,N_11110,N_11835);
and U12932 (N_12932,N_11219,N_11112);
and U12933 (N_12933,N_11327,N_11554);
and U12934 (N_12934,N_11658,N_11426);
and U12935 (N_12935,N_11480,N_11783);
and U12936 (N_12936,N_11849,N_11301);
nor U12937 (N_12937,N_11147,N_11657);
and U12938 (N_12938,N_11069,N_11143);
and U12939 (N_12939,N_11547,N_11141);
nand U12940 (N_12940,N_11275,N_11069);
xnor U12941 (N_12941,N_11889,N_11750);
xnor U12942 (N_12942,N_11235,N_11672);
nand U12943 (N_12943,N_11445,N_11601);
and U12944 (N_12944,N_11270,N_11282);
or U12945 (N_12945,N_11574,N_11994);
nand U12946 (N_12946,N_11821,N_11826);
nand U12947 (N_12947,N_11247,N_11718);
xor U12948 (N_12948,N_11546,N_11726);
or U12949 (N_12949,N_11231,N_11281);
or U12950 (N_12950,N_11288,N_11066);
nand U12951 (N_12951,N_11537,N_11814);
xor U12952 (N_12952,N_11524,N_11713);
xor U12953 (N_12953,N_11671,N_11630);
nand U12954 (N_12954,N_11700,N_11183);
nand U12955 (N_12955,N_11928,N_11079);
xnor U12956 (N_12956,N_11845,N_11613);
or U12957 (N_12957,N_11003,N_11995);
and U12958 (N_12958,N_11319,N_11501);
nand U12959 (N_12959,N_11468,N_11521);
or U12960 (N_12960,N_11724,N_11185);
and U12961 (N_12961,N_11186,N_11279);
xor U12962 (N_12962,N_11071,N_11105);
or U12963 (N_12963,N_11875,N_11118);
nor U12964 (N_12964,N_11758,N_11283);
nand U12965 (N_12965,N_11698,N_11088);
or U12966 (N_12966,N_11554,N_11277);
xnor U12967 (N_12967,N_11562,N_11741);
xor U12968 (N_12968,N_11166,N_11418);
or U12969 (N_12969,N_11253,N_11083);
xnor U12970 (N_12970,N_11252,N_11785);
or U12971 (N_12971,N_11051,N_11073);
nor U12972 (N_12972,N_11176,N_11312);
nand U12973 (N_12973,N_11241,N_11424);
nor U12974 (N_12974,N_11518,N_11018);
nor U12975 (N_12975,N_11012,N_11737);
and U12976 (N_12976,N_11694,N_11609);
nand U12977 (N_12977,N_11930,N_11059);
nor U12978 (N_12978,N_11828,N_11378);
or U12979 (N_12979,N_11212,N_11341);
and U12980 (N_12980,N_11321,N_11299);
nand U12981 (N_12981,N_11570,N_11075);
xor U12982 (N_12982,N_11511,N_11490);
nor U12983 (N_12983,N_11126,N_11938);
nor U12984 (N_12984,N_11741,N_11014);
and U12985 (N_12985,N_11998,N_11262);
xnor U12986 (N_12986,N_11197,N_11163);
xor U12987 (N_12987,N_11493,N_11420);
and U12988 (N_12988,N_11896,N_11650);
or U12989 (N_12989,N_11590,N_11215);
xnor U12990 (N_12990,N_11767,N_11034);
or U12991 (N_12991,N_11600,N_11852);
and U12992 (N_12992,N_11316,N_11300);
nand U12993 (N_12993,N_11107,N_11532);
xnor U12994 (N_12994,N_11922,N_11690);
nand U12995 (N_12995,N_11646,N_11774);
nand U12996 (N_12996,N_11041,N_11452);
nor U12997 (N_12997,N_11139,N_11797);
xnor U12998 (N_12998,N_11674,N_11931);
and U12999 (N_12999,N_11156,N_11185);
xor U13000 (N_13000,N_12390,N_12608);
xor U13001 (N_13001,N_12598,N_12404);
xnor U13002 (N_13002,N_12457,N_12983);
nor U13003 (N_13003,N_12539,N_12820);
xnor U13004 (N_13004,N_12321,N_12059);
nand U13005 (N_13005,N_12900,N_12196);
xor U13006 (N_13006,N_12437,N_12065);
or U13007 (N_13007,N_12728,N_12462);
and U13008 (N_13008,N_12541,N_12170);
and U13009 (N_13009,N_12612,N_12101);
and U13010 (N_13010,N_12543,N_12007);
nor U13011 (N_13011,N_12154,N_12791);
nor U13012 (N_13012,N_12155,N_12459);
nand U13013 (N_13013,N_12160,N_12409);
nor U13014 (N_13014,N_12184,N_12267);
nand U13015 (N_13015,N_12412,N_12518);
nor U13016 (N_13016,N_12291,N_12873);
xnor U13017 (N_13017,N_12723,N_12715);
nand U13018 (N_13018,N_12069,N_12511);
xnor U13019 (N_13019,N_12684,N_12617);
nor U13020 (N_13020,N_12984,N_12794);
xor U13021 (N_13021,N_12052,N_12844);
nand U13022 (N_13022,N_12968,N_12148);
or U13023 (N_13023,N_12955,N_12597);
and U13024 (N_13024,N_12137,N_12956);
nand U13025 (N_13025,N_12254,N_12329);
or U13026 (N_13026,N_12717,N_12009);
and U13027 (N_13027,N_12907,N_12330);
and U13028 (N_13028,N_12100,N_12662);
xor U13029 (N_13029,N_12484,N_12058);
nand U13030 (N_13030,N_12492,N_12536);
nand U13031 (N_13031,N_12111,N_12013);
nand U13032 (N_13032,N_12062,N_12260);
xor U13033 (N_13033,N_12736,N_12950);
nand U13034 (N_13034,N_12520,N_12737);
nor U13035 (N_13035,N_12243,N_12802);
xnor U13036 (N_13036,N_12314,N_12633);
nor U13037 (N_13037,N_12132,N_12050);
xor U13038 (N_13038,N_12772,N_12837);
and U13039 (N_13039,N_12973,N_12708);
and U13040 (N_13040,N_12877,N_12215);
nand U13041 (N_13041,N_12825,N_12578);
or U13042 (N_13042,N_12366,N_12290);
nor U13043 (N_13043,N_12925,N_12121);
nand U13044 (N_13044,N_12713,N_12171);
xnor U13045 (N_13045,N_12566,N_12257);
xor U13046 (N_13046,N_12821,N_12088);
and U13047 (N_13047,N_12851,N_12710);
and U13048 (N_13048,N_12365,N_12867);
nor U13049 (N_13049,N_12336,N_12174);
and U13050 (N_13050,N_12053,N_12250);
nor U13051 (N_13051,N_12477,N_12860);
xor U13052 (N_13052,N_12951,N_12341);
nand U13053 (N_13053,N_12831,N_12881);
nand U13054 (N_13054,N_12226,N_12252);
nor U13055 (N_13055,N_12754,N_12005);
nand U13056 (N_13056,N_12351,N_12985);
and U13057 (N_13057,N_12553,N_12836);
nand U13058 (N_13058,N_12499,N_12392);
or U13059 (N_13059,N_12919,N_12472);
xnor U13060 (N_13060,N_12027,N_12730);
or U13061 (N_13061,N_12380,N_12691);
and U13062 (N_13062,N_12859,N_12335);
nor U13063 (N_13063,N_12300,N_12440);
xnor U13064 (N_13064,N_12194,N_12638);
nand U13065 (N_13065,N_12699,N_12533);
and U13066 (N_13066,N_12507,N_12204);
xor U13067 (N_13067,N_12209,N_12508);
xor U13068 (N_13068,N_12588,N_12210);
or U13069 (N_13069,N_12281,N_12022);
xor U13070 (N_13070,N_12373,N_12678);
or U13071 (N_13071,N_12915,N_12801);
nand U13072 (N_13072,N_12021,N_12839);
nand U13073 (N_13073,N_12482,N_12724);
or U13074 (N_13074,N_12145,N_12406);
and U13075 (N_13075,N_12077,N_12671);
and U13076 (N_13076,N_12669,N_12551);
nand U13077 (N_13077,N_12786,N_12695);
xor U13078 (N_13078,N_12244,N_12400);
xnor U13079 (N_13079,N_12475,N_12656);
or U13080 (N_13080,N_12063,N_12562);
xnor U13081 (N_13081,N_12080,N_12711);
xor U13082 (N_13082,N_12041,N_12767);
nor U13083 (N_13083,N_12014,N_12239);
nand U13084 (N_13084,N_12283,N_12810);
and U13085 (N_13085,N_12670,N_12777);
xor U13086 (N_13086,N_12486,N_12299);
nor U13087 (N_13087,N_12798,N_12719);
nand U13088 (N_13088,N_12413,N_12641);
nor U13089 (N_13089,N_12033,N_12208);
xor U13090 (N_13090,N_12428,N_12378);
xor U13091 (N_13091,N_12280,N_12074);
nand U13092 (N_13092,N_12618,N_12948);
and U13093 (N_13093,N_12850,N_12161);
nand U13094 (N_13094,N_12784,N_12932);
nor U13095 (N_13095,N_12743,N_12371);
nor U13096 (N_13096,N_12085,N_12538);
or U13097 (N_13097,N_12768,N_12975);
or U13098 (N_13098,N_12510,N_12572);
xor U13099 (N_13099,N_12939,N_12377);
and U13100 (N_13100,N_12098,N_12011);
nand U13101 (N_13101,N_12523,N_12957);
xnor U13102 (N_13102,N_12549,N_12481);
and U13103 (N_13103,N_12463,N_12112);
nor U13104 (N_13104,N_12981,N_12182);
nor U13105 (N_13105,N_12411,N_12124);
xnor U13106 (N_13106,N_12513,N_12941);
nand U13107 (N_13107,N_12202,N_12187);
nand U13108 (N_13108,N_12331,N_12151);
and U13109 (N_13109,N_12782,N_12376);
xnor U13110 (N_13110,N_12363,N_12527);
xor U13111 (N_13111,N_12658,N_12185);
or U13112 (N_13112,N_12740,N_12640);
nand U13113 (N_13113,N_12158,N_12342);
or U13114 (N_13114,N_12051,N_12231);
nand U13115 (N_13115,N_12067,N_12890);
or U13116 (N_13116,N_12195,N_12055);
xnor U13117 (N_13117,N_12675,N_12201);
and U13118 (N_13118,N_12189,N_12455);
xor U13119 (N_13119,N_12333,N_12593);
nand U13120 (N_13120,N_12259,N_12808);
nor U13121 (N_13121,N_12910,N_12928);
nor U13122 (N_13122,N_12417,N_12146);
and U13123 (N_13123,N_12624,N_12266);
and U13124 (N_13124,N_12426,N_12150);
or U13125 (N_13125,N_12255,N_12230);
xnor U13126 (N_13126,N_12694,N_12275);
xnor U13127 (N_13127,N_12103,N_12176);
or U13128 (N_13128,N_12285,N_12357);
nor U13129 (N_13129,N_12131,N_12781);
nand U13130 (N_13130,N_12680,N_12653);
nand U13131 (N_13131,N_12010,N_12651);
nand U13132 (N_13132,N_12173,N_12727);
xnor U13133 (N_13133,N_12245,N_12818);
nand U13134 (N_13134,N_12256,N_12563);
xor U13135 (N_13135,N_12094,N_12198);
xnor U13136 (N_13136,N_12749,N_12017);
or U13137 (N_13137,N_12625,N_12620);
nor U13138 (N_13138,N_12097,N_12963);
nand U13139 (N_13139,N_12739,N_12912);
nor U13140 (N_13140,N_12982,N_12388);
nor U13141 (N_13141,N_12944,N_12138);
and U13142 (N_13142,N_12278,N_12323);
or U13143 (N_13143,N_12630,N_12833);
nor U13144 (N_13144,N_12594,N_12164);
nand U13145 (N_13145,N_12092,N_12470);
or U13146 (N_13146,N_12940,N_12992);
or U13147 (N_13147,N_12435,N_12468);
nor U13148 (N_13148,N_12502,N_12519);
or U13149 (N_13149,N_12505,N_12346);
xnor U13150 (N_13150,N_12863,N_12812);
and U13151 (N_13151,N_12783,N_12886);
xor U13152 (N_13152,N_12689,N_12071);
or U13153 (N_13153,N_12571,N_12676);
or U13154 (N_13154,N_12576,N_12908);
and U13155 (N_13155,N_12815,N_12762);
nand U13156 (N_13156,N_12157,N_12679);
and U13157 (N_13157,N_12993,N_12605);
or U13158 (N_13158,N_12177,N_12497);
xnor U13159 (N_13159,N_12879,N_12354);
or U13160 (N_13160,N_12466,N_12780);
and U13161 (N_13161,N_12116,N_12707);
and U13162 (N_13162,N_12193,N_12590);
nand U13163 (N_13163,N_12089,N_12035);
nor U13164 (N_13164,N_12232,N_12644);
xnor U13165 (N_13165,N_12720,N_12800);
xor U13166 (N_13166,N_12596,N_12504);
and U13167 (N_13167,N_12733,N_12672);
xor U13168 (N_13168,N_12805,N_12073);
and U13169 (N_13169,N_12872,N_12978);
nor U13170 (N_13170,N_12967,N_12826);
xnor U13171 (N_13171,N_12445,N_12178);
or U13172 (N_13172,N_12129,N_12359);
nor U13173 (N_13173,N_12034,N_12559);
nor U13174 (N_13174,N_12828,N_12474);
nand U13175 (N_13175,N_12407,N_12238);
nand U13176 (N_13176,N_12084,N_12582);
and U13177 (N_13177,N_12082,N_12652);
xnor U13178 (N_13178,N_12251,N_12569);
nor U13179 (N_13179,N_12667,N_12473);
nor U13180 (N_13180,N_12169,N_12337);
nor U13181 (N_13181,N_12483,N_12424);
or U13182 (N_13182,N_12528,N_12319);
or U13183 (N_13183,N_12580,N_12235);
nand U13184 (N_13184,N_12199,N_12374);
xor U13185 (N_13185,N_12382,N_12313);
or U13186 (N_13186,N_12494,N_12954);
nor U13187 (N_13187,N_12722,N_12835);
nand U13188 (N_13188,N_12126,N_12862);
and U13189 (N_13189,N_12990,N_12353);
nor U13190 (N_13190,N_12396,N_12343);
or U13191 (N_13191,N_12522,N_12107);
nor U13192 (N_13192,N_12642,N_12159);
xnor U13193 (N_13193,N_12287,N_12217);
or U13194 (N_13194,N_12056,N_12712);
nor U13195 (N_13195,N_12690,N_12247);
and U13196 (N_13196,N_12852,N_12697);
xor U13197 (N_13197,N_12842,N_12935);
and U13198 (N_13198,N_12262,N_12276);
or U13199 (N_13199,N_12156,N_12619);
and U13200 (N_13200,N_12449,N_12813);
and U13201 (N_13201,N_12627,N_12289);
nor U13202 (N_13202,N_12431,N_12391);
and U13203 (N_13203,N_12930,N_12047);
nor U13204 (N_13204,N_12205,N_12264);
nand U13205 (N_13205,N_12261,N_12586);
or U13206 (N_13206,N_12921,N_12222);
nor U13207 (N_13207,N_12296,N_12996);
or U13208 (N_13208,N_12302,N_12856);
nor U13209 (N_13209,N_12503,N_12478);
nor U13210 (N_13210,N_12600,N_12583);
or U13211 (N_13211,N_12393,N_12905);
xnor U13212 (N_13212,N_12420,N_12358);
nor U13213 (N_13213,N_12240,N_12488);
or U13214 (N_13214,N_12143,N_12175);
xnor U13215 (N_13215,N_12534,N_12911);
or U13216 (N_13216,N_12628,N_12493);
nand U13217 (N_13217,N_12414,N_12514);
and U13218 (N_13218,N_12117,N_12105);
nand U13219 (N_13219,N_12004,N_12415);
xnor U13220 (N_13220,N_12725,N_12423);
xnor U13221 (N_13221,N_12030,N_12855);
xor U13222 (N_13222,N_12344,N_12854);
nor U13223 (N_13223,N_12368,N_12292);
or U13224 (N_13224,N_12109,N_12375);
nand U13225 (N_13225,N_12726,N_12946);
or U13226 (N_13226,N_12634,N_12848);
nor U13227 (N_13227,N_12830,N_12183);
or U13228 (N_13228,N_12495,N_12626);
or U13229 (N_13229,N_12748,N_12362);
nor U13230 (N_13230,N_12448,N_12003);
or U13231 (N_13231,N_12389,N_12229);
and U13232 (N_13232,N_12308,N_12914);
or U13233 (N_13233,N_12703,N_12552);
and U13234 (N_13234,N_12309,N_12585);
or U13235 (N_13235,N_12076,N_12949);
nand U13236 (N_13236,N_12405,N_12714);
and U13237 (N_13237,N_12961,N_12153);
or U13238 (N_13238,N_12326,N_12370);
nor U13239 (N_13239,N_12937,N_12874);
and U13240 (N_13240,N_12698,N_12091);
and U13241 (N_13241,N_12168,N_12896);
or U13242 (N_13242,N_12347,N_12603);
xor U13243 (N_13243,N_12803,N_12995);
nand U13244 (N_13244,N_12310,N_12303);
nand U13245 (N_13245,N_12904,N_12249);
or U13246 (N_13246,N_12115,N_12757);
and U13247 (N_13247,N_12688,N_12832);
and U13248 (N_13248,N_12870,N_12847);
nand U13249 (N_13249,N_12660,N_12338);
or U13250 (N_13250,N_12899,N_12755);
and U13251 (N_13251,N_12573,N_12408);
or U13252 (N_13252,N_12364,N_12685);
nor U13253 (N_13253,N_12491,N_12057);
nand U13254 (N_13254,N_12643,N_12425);
and U13255 (N_13255,N_12064,N_12386);
xor U13256 (N_13256,N_12316,N_12324);
xnor U13257 (N_13257,N_12632,N_12958);
nand U13258 (N_13258,N_12927,N_12970);
or U13259 (N_13259,N_12043,N_12273);
nor U13260 (N_13260,N_12317,N_12123);
and U13261 (N_13261,N_12891,N_12804);
or U13262 (N_13262,N_12467,N_12019);
or U13263 (N_13263,N_12133,N_12384);
xnor U13264 (N_13264,N_12277,N_12433);
nor U13265 (N_13265,N_12190,N_12540);
and U13266 (N_13266,N_12040,N_12785);
nand U13267 (N_13267,N_12796,N_12997);
nand U13268 (N_13268,N_12942,N_12165);
and U13269 (N_13269,N_12284,N_12769);
nor U13270 (N_13270,N_12451,N_12339);
xnor U13271 (N_13271,N_12480,N_12136);
xnor U13272 (N_13272,N_12090,N_12795);
nand U13273 (N_13273,N_12306,N_12295);
xnor U13274 (N_13274,N_12489,N_12361);
or U13275 (N_13275,N_12427,N_12648);
xor U13276 (N_13276,N_12381,N_12422);
xnor U13277 (N_13277,N_12456,N_12673);
nand U13278 (N_13278,N_12227,N_12207);
nand U13279 (N_13279,N_12591,N_12840);
or U13280 (N_13280,N_12248,N_12841);
and U13281 (N_13281,N_12152,N_12923);
and U13282 (N_13282,N_12735,N_12977);
or U13283 (N_13283,N_12438,N_12677);
nand U13284 (N_13284,N_12631,N_12587);
nand U13285 (N_13285,N_12635,N_12203);
and U13286 (N_13286,N_12696,N_12385);
and U13287 (N_13287,N_12530,N_12895);
or U13288 (N_13288,N_12766,N_12060);
xor U13289 (N_13289,N_12788,N_12403);
or U13290 (N_13290,N_12853,N_12501);
xnor U13291 (N_13291,N_12212,N_12687);
nor U13292 (N_13292,N_12721,N_12953);
xnor U13293 (N_13293,N_12750,N_12646);
nand U13294 (N_13294,N_12924,N_12966);
or U13295 (N_13295,N_12599,N_12139);
nor U13296 (N_13296,N_12716,N_12779);
nor U13297 (N_13297,N_12824,N_12607);
nor U13298 (N_13298,N_12500,N_12888);
and U13299 (N_13299,N_12998,N_12016);
xor U13300 (N_13300,N_12629,N_12379);
nor U13301 (N_13301,N_12332,N_12130);
nor U13302 (N_13302,N_12621,N_12054);
nor U13303 (N_13303,N_12294,N_12147);
or U13304 (N_13304,N_12356,N_12926);
and U13305 (N_13305,N_12845,N_12272);
and U13306 (N_13306,N_12241,N_12706);
and U13307 (N_13307,N_12452,N_12464);
and U13308 (N_13308,N_12893,N_12061);
nor U13309 (N_13309,N_12086,N_12246);
or U13310 (N_13310,N_12668,N_12418);
xor U13311 (N_13311,N_12218,N_12439);
or U13312 (N_13312,N_12929,N_12799);
xnor U13313 (N_13313,N_12221,N_12809);
nor U13314 (N_13314,N_12894,N_12979);
and U13315 (N_13315,N_12823,N_12297);
xor U13316 (N_13316,N_12142,N_12609);
or U13317 (N_13317,N_12592,N_12616);
and U13318 (N_13318,N_12535,N_12988);
or U13319 (N_13319,N_12118,N_12878);
or U13320 (N_13320,N_12038,N_12729);
xor U13321 (N_13321,N_12991,N_12807);
nand U13322 (N_13322,N_12869,N_12490);
xor U13323 (N_13323,N_12328,N_12102);
and U13324 (N_13324,N_12686,N_12570);
nor U13325 (N_13325,N_12134,N_12738);
nor U13326 (N_13326,N_12223,N_12663);
xnor U13327 (N_13327,N_12399,N_12846);
xor U13328 (N_13328,N_12402,N_12545);
xor U13329 (N_13329,N_12301,N_12253);
and U13330 (N_13330,N_12775,N_12270);
nand U13331 (N_13331,N_12647,N_12623);
nor U13332 (N_13332,N_12681,N_12822);
nand U13333 (N_13333,N_12446,N_12037);
nand U13334 (N_13334,N_12293,N_12564);
nor U13335 (N_13335,N_12104,N_12471);
or U13336 (N_13336,N_12318,N_12601);
and U13337 (N_13337,N_12884,N_12320);
nor U13338 (N_13338,N_12745,N_12880);
or U13339 (N_13339,N_12485,N_12465);
nor U13340 (N_13340,N_12233,N_12920);
and U13341 (N_13341,N_12188,N_12352);
or U13342 (N_13342,N_12135,N_12649);
and U13343 (N_13343,N_12072,N_12565);
and U13344 (N_13344,N_12447,N_12639);
xor U13345 (N_13345,N_12849,N_12305);
nor U13346 (N_13346,N_12348,N_12093);
xnor U13347 (N_13347,N_12700,N_12555);
and U13348 (N_13348,N_12959,N_12122);
xor U13349 (N_13349,N_12015,N_12312);
and U13350 (N_13350,N_12219,N_12611);
nand U13351 (N_13351,N_12546,N_12531);
or U13352 (N_13352,N_12816,N_12980);
nor U13353 (N_13353,N_12454,N_12692);
nor U13354 (N_13354,N_12225,N_12263);
nand U13355 (N_13355,N_12683,N_12443);
or U13356 (N_13356,N_12661,N_12524);
xnor U13357 (N_13357,N_12216,N_12797);
or U13358 (N_13358,N_12001,N_12568);
nor U13359 (N_13359,N_12211,N_12416);
or U13360 (N_13360,N_12179,N_12974);
nor U13361 (N_13361,N_12916,N_12584);
or U13362 (N_13362,N_12498,N_12934);
xor U13363 (N_13363,N_12141,N_12909);
xnor U13364 (N_13364,N_12577,N_12023);
nand U13365 (N_13365,N_12410,N_12018);
nor U13366 (N_13366,N_12875,N_12645);
and U13367 (N_13367,N_12114,N_12561);
nor U13368 (N_13368,N_12224,N_12106);
and U13369 (N_13369,N_12560,N_12327);
nor U13370 (N_13370,N_12311,N_12945);
xnor U13371 (N_13371,N_12008,N_12206);
nor U13372 (N_13372,N_12602,N_12614);
and U13373 (N_13373,N_12265,N_12012);
and U13374 (N_13374,N_12039,N_12044);
xor U13375 (N_13375,N_12322,N_12127);
or U13376 (N_13376,N_12771,N_12657);
nor U13377 (N_13377,N_12989,N_12355);
nand U13378 (N_13378,N_12972,N_12579);
and U13379 (N_13379,N_12119,N_12025);
xnor U13380 (N_13380,N_12237,N_12838);
nor U13381 (N_13381,N_12819,N_12049);
and U13382 (N_13382,N_12655,N_12479);
or U13383 (N_13383,N_12702,N_12476);
and U13384 (N_13384,N_12436,N_12761);
and U13385 (N_13385,N_12718,N_12242);
xnor U13386 (N_13386,N_12458,N_12163);
nand U13387 (N_13387,N_12971,N_12931);
xnor U13388 (N_13388,N_12774,N_12020);
or U13389 (N_13389,N_12704,N_12705);
nand U13390 (N_13390,N_12637,N_12120);
and U13391 (N_13391,N_12140,N_12360);
nor U13392 (N_13392,N_12394,N_12747);
nand U13393 (N_13393,N_12889,N_12834);
and U13394 (N_13394,N_12734,N_12192);
nor U13395 (N_13395,N_12763,N_12885);
nor U13396 (N_13396,N_12567,N_12434);
and U13397 (N_13397,N_12024,N_12753);
nand U13398 (N_13398,N_12334,N_12764);
nand U13399 (N_13399,N_12172,N_12913);
or U13400 (N_13400,N_12419,N_12048);
or U13401 (N_13401,N_12550,N_12081);
nand U13402 (N_13402,N_12078,N_12397);
and U13403 (N_13403,N_12487,N_12516);
and U13404 (N_13404,N_12922,N_12269);
xnor U13405 (N_13405,N_12751,N_12087);
xor U13406 (N_13406,N_12066,N_12271);
or U13407 (N_13407,N_12228,N_12960);
and U13408 (N_13408,N_12773,N_12843);
nand U13409 (N_13409,N_12031,N_12028);
and U13410 (N_13410,N_12181,N_12682);
nor U13411 (N_13411,N_12383,N_12595);
xnor U13412 (N_13412,N_12110,N_12936);
or U13413 (N_13413,N_12636,N_12046);
nor U13414 (N_13414,N_12986,N_12918);
and U13415 (N_13415,N_12898,N_12315);
or U13416 (N_13416,N_12864,N_12026);
xor U13417 (N_13417,N_12108,N_12298);
nor U13418 (N_13418,N_12674,N_12079);
and U13419 (N_13419,N_12547,N_12000);
and U13420 (N_13420,N_12180,N_12191);
nand U13421 (N_13421,N_12964,N_12792);
or U13422 (N_13422,N_12162,N_12529);
and U13423 (N_13423,N_12515,N_12128);
xor U13424 (N_13424,N_12654,N_12613);
and U13425 (N_13425,N_12200,N_12892);
or U13426 (N_13426,N_12962,N_12906);
and U13427 (N_13427,N_12075,N_12744);
xnor U13428 (N_13428,N_12943,N_12917);
or U13429 (N_13429,N_12307,N_12701);
nand U13430 (N_13430,N_12268,N_12902);
or U13431 (N_13431,N_12282,N_12901);
or U13432 (N_13432,N_12537,N_12793);
xor U13433 (N_13433,N_12526,N_12589);
or U13434 (N_13434,N_12665,N_12525);
nor U13435 (N_13435,N_12969,N_12756);
or U13436 (N_13436,N_12758,N_12166);
or U13437 (N_13437,N_12113,N_12532);
nor U13438 (N_13438,N_12350,N_12125);
xnor U13439 (N_13439,N_12096,N_12778);
nor U13440 (N_13440,N_12395,N_12857);
or U13441 (N_13441,N_12461,N_12994);
or U13442 (N_13442,N_12236,N_12469);
or U13443 (N_13443,N_12544,N_12167);
nor U13444 (N_13444,N_12036,N_12548);
and U13445 (N_13445,N_12770,N_12759);
nand U13446 (N_13446,N_12421,N_12650);
or U13447 (N_13447,N_12610,N_12325);
and U13448 (N_13448,N_12517,N_12938);
or U13449 (N_13449,N_12509,N_12542);
and U13450 (N_13450,N_12398,N_12790);
xnor U13451 (N_13451,N_12866,N_12622);
xor U13452 (N_13452,N_12045,N_12387);
or U13453 (N_13453,N_12876,N_12868);
or U13454 (N_13454,N_12042,N_12442);
and U13455 (N_13455,N_12430,N_12947);
xnor U13456 (N_13456,N_12987,N_12760);
nor U13457 (N_13457,N_12976,N_12095);
nand U13458 (N_13458,N_12732,N_12731);
nand U13459 (N_13459,N_12444,N_12817);
and U13460 (N_13460,N_12234,N_12693);
nand U13461 (N_13461,N_12861,N_12002);
xor U13462 (N_13462,N_12742,N_12554);
nand U13463 (N_13463,N_12070,N_12068);
and U13464 (N_13464,N_12664,N_12933);
and U13465 (N_13465,N_12372,N_12741);
xor U13466 (N_13466,N_12214,N_12186);
and U13467 (N_13467,N_12882,N_12197);
nand U13468 (N_13468,N_12441,N_12709);
and U13469 (N_13469,N_12099,N_12258);
nand U13470 (N_13470,N_12220,N_12558);
nand U13471 (N_13471,N_12369,N_12032);
xor U13472 (N_13472,N_12345,N_12083);
xor U13473 (N_13473,N_12811,N_12897);
xor U13474 (N_13474,N_12829,N_12659);
nand U13475 (N_13475,N_12776,N_12367);
and U13476 (N_13476,N_12460,N_12858);
or U13477 (N_13477,N_12887,N_12765);
nand U13478 (N_13478,N_12752,N_12666);
or U13479 (N_13479,N_12274,N_12006);
nor U13480 (N_13480,N_12574,N_12581);
nor U13481 (N_13481,N_12279,N_12787);
nor U13482 (N_13482,N_12149,N_12304);
nor U13483 (N_13483,N_12286,N_12506);
nand U13484 (N_13484,N_12557,N_12556);
xor U13485 (N_13485,N_12450,N_12512);
and U13486 (N_13486,N_12453,N_12903);
xnor U13487 (N_13487,N_12521,N_12806);
nor U13488 (N_13488,N_12746,N_12288);
and U13489 (N_13489,N_12865,N_12349);
or U13490 (N_13490,N_12606,N_12789);
nor U13491 (N_13491,N_12604,N_12999);
and U13492 (N_13492,N_12814,N_12496);
or U13493 (N_13493,N_12965,N_12429);
xor U13494 (N_13494,N_12144,N_12401);
and U13495 (N_13495,N_12952,N_12213);
xor U13496 (N_13496,N_12575,N_12340);
and U13497 (N_13497,N_12827,N_12432);
nand U13498 (N_13498,N_12871,N_12883);
nor U13499 (N_13499,N_12029,N_12615);
nand U13500 (N_13500,N_12466,N_12079);
and U13501 (N_13501,N_12209,N_12886);
xor U13502 (N_13502,N_12771,N_12173);
nor U13503 (N_13503,N_12263,N_12213);
or U13504 (N_13504,N_12100,N_12526);
xor U13505 (N_13505,N_12955,N_12917);
nor U13506 (N_13506,N_12619,N_12979);
or U13507 (N_13507,N_12282,N_12096);
xnor U13508 (N_13508,N_12031,N_12507);
and U13509 (N_13509,N_12345,N_12358);
nand U13510 (N_13510,N_12388,N_12899);
and U13511 (N_13511,N_12526,N_12887);
and U13512 (N_13512,N_12593,N_12580);
xnor U13513 (N_13513,N_12660,N_12468);
xor U13514 (N_13514,N_12410,N_12534);
nand U13515 (N_13515,N_12889,N_12590);
and U13516 (N_13516,N_12398,N_12558);
nor U13517 (N_13517,N_12038,N_12060);
nand U13518 (N_13518,N_12016,N_12404);
and U13519 (N_13519,N_12507,N_12623);
nand U13520 (N_13520,N_12834,N_12075);
nand U13521 (N_13521,N_12620,N_12450);
or U13522 (N_13522,N_12093,N_12392);
or U13523 (N_13523,N_12756,N_12629);
and U13524 (N_13524,N_12983,N_12253);
and U13525 (N_13525,N_12000,N_12030);
nor U13526 (N_13526,N_12834,N_12763);
nor U13527 (N_13527,N_12884,N_12999);
nor U13528 (N_13528,N_12639,N_12308);
nand U13529 (N_13529,N_12176,N_12969);
or U13530 (N_13530,N_12524,N_12149);
nor U13531 (N_13531,N_12359,N_12695);
and U13532 (N_13532,N_12149,N_12162);
xor U13533 (N_13533,N_12434,N_12854);
or U13534 (N_13534,N_12098,N_12552);
nor U13535 (N_13535,N_12853,N_12468);
and U13536 (N_13536,N_12766,N_12642);
and U13537 (N_13537,N_12315,N_12263);
nor U13538 (N_13538,N_12070,N_12262);
nand U13539 (N_13539,N_12643,N_12406);
or U13540 (N_13540,N_12001,N_12803);
nand U13541 (N_13541,N_12989,N_12001);
nand U13542 (N_13542,N_12275,N_12971);
and U13543 (N_13543,N_12325,N_12422);
nand U13544 (N_13544,N_12136,N_12466);
or U13545 (N_13545,N_12259,N_12189);
or U13546 (N_13546,N_12144,N_12240);
nor U13547 (N_13547,N_12692,N_12782);
nand U13548 (N_13548,N_12182,N_12116);
and U13549 (N_13549,N_12660,N_12454);
and U13550 (N_13550,N_12778,N_12984);
nand U13551 (N_13551,N_12163,N_12354);
or U13552 (N_13552,N_12021,N_12593);
nor U13553 (N_13553,N_12128,N_12568);
nand U13554 (N_13554,N_12977,N_12207);
nor U13555 (N_13555,N_12666,N_12565);
xnor U13556 (N_13556,N_12874,N_12154);
nor U13557 (N_13557,N_12504,N_12678);
and U13558 (N_13558,N_12170,N_12841);
and U13559 (N_13559,N_12683,N_12141);
and U13560 (N_13560,N_12471,N_12349);
and U13561 (N_13561,N_12013,N_12449);
or U13562 (N_13562,N_12947,N_12219);
and U13563 (N_13563,N_12692,N_12142);
nor U13564 (N_13564,N_12563,N_12622);
and U13565 (N_13565,N_12207,N_12455);
xor U13566 (N_13566,N_12941,N_12592);
nor U13567 (N_13567,N_12884,N_12428);
and U13568 (N_13568,N_12812,N_12190);
or U13569 (N_13569,N_12133,N_12879);
nand U13570 (N_13570,N_12213,N_12442);
or U13571 (N_13571,N_12391,N_12264);
nor U13572 (N_13572,N_12162,N_12013);
nor U13573 (N_13573,N_12737,N_12257);
xnor U13574 (N_13574,N_12607,N_12881);
or U13575 (N_13575,N_12181,N_12759);
nand U13576 (N_13576,N_12400,N_12705);
xor U13577 (N_13577,N_12767,N_12692);
or U13578 (N_13578,N_12238,N_12572);
and U13579 (N_13579,N_12471,N_12765);
or U13580 (N_13580,N_12297,N_12279);
nor U13581 (N_13581,N_12393,N_12128);
or U13582 (N_13582,N_12706,N_12609);
nor U13583 (N_13583,N_12536,N_12441);
and U13584 (N_13584,N_12505,N_12971);
xor U13585 (N_13585,N_12243,N_12879);
and U13586 (N_13586,N_12734,N_12603);
and U13587 (N_13587,N_12738,N_12032);
nand U13588 (N_13588,N_12397,N_12721);
nand U13589 (N_13589,N_12688,N_12510);
and U13590 (N_13590,N_12089,N_12157);
nor U13591 (N_13591,N_12507,N_12461);
and U13592 (N_13592,N_12193,N_12136);
or U13593 (N_13593,N_12821,N_12033);
xnor U13594 (N_13594,N_12760,N_12705);
nor U13595 (N_13595,N_12034,N_12623);
xnor U13596 (N_13596,N_12079,N_12594);
or U13597 (N_13597,N_12310,N_12872);
and U13598 (N_13598,N_12802,N_12238);
and U13599 (N_13599,N_12411,N_12628);
xnor U13600 (N_13600,N_12042,N_12585);
and U13601 (N_13601,N_12285,N_12091);
nor U13602 (N_13602,N_12967,N_12787);
nand U13603 (N_13603,N_12034,N_12715);
nor U13604 (N_13604,N_12083,N_12035);
nand U13605 (N_13605,N_12322,N_12804);
or U13606 (N_13606,N_12085,N_12554);
nand U13607 (N_13607,N_12989,N_12432);
nand U13608 (N_13608,N_12180,N_12864);
nand U13609 (N_13609,N_12315,N_12948);
nor U13610 (N_13610,N_12269,N_12500);
nand U13611 (N_13611,N_12576,N_12756);
and U13612 (N_13612,N_12485,N_12505);
and U13613 (N_13613,N_12817,N_12504);
and U13614 (N_13614,N_12632,N_12363);
or U13615 (N_13615,N_12020,N_12127);
or U13616 (N_13616,N_12346,N_12741);
or U13617 (N_13617,N_12298,N_12480);
nor U13618 (N_13618,N_12752,N_12761);
or U13619 (N_13619,N_12943,N_12298);
xor U13620 (N_13620,N_12192,N_12895);
nor U13621 (N_13621,N_12654,N_12335);
xor U13622 (N_13622,N_12843,N_12034);
nand U13623 (N_13623,N_12041,N_12919);
nor U13624 (N_13624,N_12892,N_12433);
and U13625 (N_13625,N_12982,N_12282);
and U13626 (N_13626,N_12645,N_12001);
and U13627 (N_13627,N_12380,N_12954);
and U13628 (N_13628,N_12285,N_12027);
nand U13629 (N_13629,N_12653,N_12764);
nor U13630 (N_13630,N_12395,N_12031);
xnor U13631 (N_13631,N_12257,N_12210);
xnor U13632 (N_13632,N_12954,N_12220);
and U13633 (N_13633,N_12506,N_12741);
or U13634 (N_13634,N_12799,N_12861);
nand U13635 (N_13635,N_12462,N_12123);
nor U13636 (N_13636,N_12276,N_12136);
nand U13637 (N_13637,N_12471,N_12115);
or U13638 (N_13638,N_12790,N_12517);
nand U13639 (N_13639,N_12958,N_12565);
or U13640 (N_13640,N_12783,N_12671);
nor U13641 (N_13641,N_12997,N_12041);
nand U13642 (N_13642,N_12051,N_12778);
and U13643 (N_13643,N_12583,N_12227);
xor U13644 (N_13644,N_12181,N_12510);
and U13645 (N_13645,N_12196,N_12449);
xnor U13646 (N_13646,N_12962,N_12747);
and U13647 (N_13647,N_12395,N_12605);
or U13648 (N_13648,N_12494,N_12847);
xnor U13649 (N_13649,N_12844,N_12782);
or U13650 (N_13650,N_12142,N_12405);
and U13651 (N_13651,N_12088,N_12528);
or U13652 (N_13652,N_12146,N_12144);
or U13653 (N_13653,N_12315,N_12729);
or U13654 (N_13654,N_12724,N_12152);
nand U13655 (N_13655,N_12165,N_12228);
xor U13656 (N_13656,N_12346,N_12121);
nand U13657 (N_13657,N_12793,N_12728);
xnor U13658 (N_13658,N_12796,N_12896);
nor U13659 (N_13659,N_12467,N_12457);
xor U13660 (N_13660,N_12711,N_12844);
or U13661 (N_13661,N_12481,N_12218);
xnor U13662 (N_13662,N_12667,N_12394);
nand U13663 (N_13663,N_12283,N_12873);
and U13664 (N_13664,N_12328,N_12662);
nor U13665 (N_13665,N_12753,N_12401);
or U13666 (N_13666,N_12801,N_12972);
xor U13667 (N_13667,N_12442,N_12460);
and U13668 (N_13668,N_12438,N_12569);
and U13669 (N_13669,N_12363,N_12868);
nand U13670 (N_13670,N_12366,N_12126);
and U13671 (N_13671,N_12086,N_12647);
nor U13672 (N_13672,N_12950,N_12362);
and U13673 (N_13673,N_12596,N_12279);
nor U13674 (N_13674,N_12577,N_12228);
and U13675 (N_13675,N_12184,N_12060);
nand U13676 (N_13676,N_12963,N_12547);
nor U13677 (N_13677,N_12509,N_12321);
nand U13678 (N_13678,N_12829,N_12081);
nand U13679 (N_13679,N_12168,N_12351);
xor U13680 (N_13680,N_12216,N_12511);
nand U13681 (N_13681,N_12318,N_12091);
and U13682 (N_13682,N_12500,N_12842);
xnor U13683 (N_13683,N_12681,N_12152);
nor U13684 (N_13684,N_12467,N_12826);
xnor U13685 (N_13685,N_12700,N_12158);
xor U13686 (N_13686,N_12698,N_12656);
and U13687 (N_13687,N_12377,N_12299);
or U13688 (N_13688,N_12005,N_12472);
and U13689 (N_13689,N_12475,N_12644);
xor U13690 (N_13690,N_12183,N_12540);
xor U13691 (N_13691,N_12161,N_12990);
or U13692 (N_13692,N_12072,N_12327);
and U13693 (N_13693,N_12522,N_12019);
xnor U13694 (N_13694,N_12937,N_12913);
or U13695 (N_13695,N_12438,N_12425);
and U13696 (N_13696,N_12373,N_12913);
nor U13697 (N_13697,N_12741,N_12338);
xnor U13698 (N_13698,N_12998,N_12178);
nand U13699 (N_13699,N_12328,N_12534);
nand U13700 (N_13700,N_12740,N_12755);
or U13701 (N_13701,N_12871,N_12668);
and U13702 (N_13702,N_12064,N_12125);
xnor U13703 (N_13703,N_12393,N_12114);
and U13704 (N_13704,N_12193,N_12522);
and U13705 (N_13705,N_12942,N_12591);
nor U13706 (N_13706,N_12610,N_12078);
xor U13707 (N_13707,N_12594,N_12745);
xor U13708 (N_13708,N_12237,N_12737);
or U13709 (N_13709,N_12223,N_12062);
or U13710 (N_13710,N_12245,N_12183);
or U13711 (N_13711,N_12627,N_12797);
and U13712 (N_13712,N_12869,N_12948);
nor U13713 (N_13713,N_12079,N_12309);
xnor U13714 (N_13714,N_12303,N_12998);
nor U13715 (N_13715,N_12860,N_12432);
xor U13716 (N_13716,N_12933,N_12634);
nand U13717 (N_13717,N_12242,N_12304);
nand U13718 (N_13718,N_12526,N_12319);
xnor U13719 (N_13719,N_12341,N_12660);
nor U13720 (N_13720,N_12105,N_12821);
xnor U13721 (N_13721,N_12483,N_12701);
xnor U13722 (N_13722,N_12874,N_12943);
nor U13723 (N_13723,N_12171,N_12625);
nand U13724 (N_13724,N_12028,N_12354);
nor U13725 (N_13725,N_12364,N_12921);
nand U13726 (N_13726,N_12551,N_12426);
or U13727 (N_13727,N_12871,N_12546);
nand U13728 (N_13728,N_12044,N_12483);
nor U13729 (N_13729,N_12295,N_12077);
nand U13730 (N_13730,N_12585,N_12449);
nand U13731 (N_13731,N_12993,N_12488);
nor U13732 (N_13732,N_12075,N_12334);
nand U13733 (N_13733,N_12219,N_12852);
nand U13734 (N_13734,N_12319,N_12765);
nand U13735 (N_13735,N_12659,N_12388);
nor U13736 (N_13736,N_12523,N_12603);
xnor U13737 (N_13737,N_12352,N_12379);
nor U13738 (N_13738,N_12573,N_12679);
nand U13739 (N_13739,N_12085,N_12237);
nor U13740 (N_13740,N_12433,N_12829);
and U13741 (N_13741,N_12702,N_12837);
nor U13742 (N_13742,N_12107,N_12132);
nor U13743 (N_13743,N_12274,N_12950);
nor U13744 (N_13744,N_12857,N_12664);
nor U13745 (N_13745,N_12104,N_12983);
xor U13746 (N_13746,N_12704,N_12975);
nand U13747 (N_13747,N_12199,N_12418);
nand U13748 (N_13748,N_12655,N_12212);
and U13749 (N_13749,N_12936,N_12120);
and U13750 (N_13750,N_12606,N_12346);
nor U13751 (N_13751,N_12859,N_12464);
nand U13752 (N_13752,N_12489,N_12384);
nor U13753 (N_13753,N_12827,N_12510);
xnor U13754 (N_13754,N_12484,N_12551);
nand U13755 (N_13755,N_12364,N_12032);
nand U13756 (N_13756,N_12814,N_12606);
nor U13757 (N_13757,N_12869,N_12923);
nand U13758 (N_13758,N_12957,N_12395);
nor U13759 (N_13759,N_12508,N_12918);
or U13760 (N_13760,N_12258,N_12628);
nand U13761 (N_13761,N_12482,N_12337);
nor U13762 (N_13762,N_12478,N_12024);
nor U13763 (N_13763,N_12382,N_12663);
and U13764 (N_13764,N_12051,N_12947);
and U13765 (N_13765,N_12077,N_12100);
or U13766 (N_13766,N_12995,N_12548);
and U13767 (N_13767,N_12163,N_12809);
and U13768 (N_13768,N_12341,N_12616);
or U13769 (N_13769,N_12937,N_12825);
nand U13770 (N_13770,N_12326,N_12319);
nand U13771 (N_13771,N_12054,N_12928);
nand U13772 (N_13772,N_12878,N_12634);
xor U13773 (N_13773,N_12144,N_12311);
nand U13774 (N_13774,N_12806,N_12366);
nor U13775 (N_13775,N_12652,N_12396);
and U13776 (N_13776,N_12941,N_12828);
and U13777 (N_13777,N_12242,N_12040);
nor U13778 (N_13778,N_12262,N_12856);
xnor U13779 (N_13779,N_12112,N_12817);
nor U13780 (N_13780,N_12645,N_12856);
nor U13781 (N_13781,N_12930,N_12524);
nor U13782 (N_13782,N_12077,N_12587);
xor U13783 (N_13783,N_12733,N_12416);
and U13784 (N_13784,N_12338,N_12159);
or U13785 (N_13785,N_12016,N_12030);
nor U13786 (N_13786,N_12484,N_12140);
nor U13787 (N_13787,N_12346,N_12403);
and U13788 (N_13788,N_12026,N_12187);
and U13789 (N_13789,N_12727,N_12219);
xnor U13790 (N_13790,N_12978,N_12141);
nand U13791 (N_13791,N_12449,N_12333);
and U13792 (N_13792,N_12042,N_12095);
or U13793 (N_13793,N_12984,N_12251);
xnor U13794 (N_13794,N_12345,N_12837);
xnor U13795 (N_13795,N_12228,N_12152);
nand U13796 (N_13796,N_12721,N_12997);
nor U13797 (N_13797,N_12736,N_12039);
xnor U13798 (N_13798,N_12080,N_12273);
and U13799 (N_13799,N_12194,N_12326);
xnor U13800 (N_13800,N_12504,N_12975);
xnor U13801 (N_13801,N_12557,N_12756);
nor U13802 (N_13802,N_12084,N_12344);
nor U13803 (N_13803,N_12887,N_12787);
nor U13804 (N_13804,N_12284,N_12854);
xnor U13805 (N_13805,N_12154,N_12266);
xor U13806 (N_13806,N_12617,N_12922);
xnor U13807 (N_13807,N_12172,N_12383);
and U13808 (N_13808,N_12623,N_12791);
xor U13809 (N_13809,N_12209,N_12699);
or U13810 (N_13810,N_12860,N_12963);
and U13811 (N_13811,N_12602,N_12586);
nor U13812 (N_13812,N_12322,N_12077);
xnor U13813 (N_13813,N_12459,N_12228);
and U13814 (N_13814,N_12401,N_12463);
nand U13815 (N_13815,N_12818,N_12806);
nor U13816 (N_13816,N_12184,N_12523);
xnor U13817 (N_13817,N_12505,N_12288);
and U13818 (N_13818,N_12507,N_12938);
or U13819 (N_13819,N_12122,N_12932);
nand U13820 (N_13820,N_12336,N_12467);
and U13821 (N_13821,N_12348,N_12978);
xnor U13822 (N_13822,N_12568,N_12434);
xnor U13823 (N_13823,N_12855,N_12035);
nand U13824 (N_13824,N_12196,N_12625);
or U13825 (N_13825,N_12278,N_12108);
or U13826 (N_13826,N_12242,N_12565);
nor U13827 (N_13827,N_12804,N_12398);
or U13828 (N_13828,N_12580,N_12883);
and U13829 (N_13829,N_12048,N_12112);
nand U13830 (N_13830,N_12685,N_12457);
or U13831 (N_13831,N_12205,N_12638);
and U13832 (N_13832,N_12298,N_12915);
or U13833 (N_13833,N_12491,N_12915);
xor U13834 (N_13834,N_12350,N_12778);
nand U13835 (N_13835,N_12664,N_12887);
xor U13836 (N_13836,N_12628,N_12390);
xor U13837 (N_13837,N_12570,N_12028);
nor U13838 (N_13838,N_12829,N_12477);
and U13839 (N_13839,N_12984,N_12805);
and U13840 (N_13840,N_12940,N_12990);
xor U13841 (N_13841,N_12161,N_12181);
and U13842 (N_13842,N_12218,N_12848);
or U13843 (N_13843,N_12329,N_12169);
or U13844 (N_13844,N_12725,N_12102);
or U13845 (N_13845,N_12254,N_12375);
nor U13846 (N_13846,N_12259,N_12057);
nand U13847 (N_13847,N_12723,N_12147);
and U13848 (N_13848,N_12420,N_12034);
xnor U13849 (N_13849,N_12005,N_12792);
and U13850 (N_13850,N_12986,N_12216);
and U13851 (N_13851,N_12974,N_12222);
and U13852 (N_13852,N_12258,N_12749);
nand U13853 (N_13853,N_12745,N_12900);
xnor U13854 (N_13854,N_12942,N_12903);
or U13855 (N_13855,N_12408,N_12710);
or U13856 (N_13856,N_12104,N_12715);
or U13857 (N_13857,N_12959,N_12807);
or U13858 (N_13858,N_12995,N_12261);
and U13859 (N_13859,N_12221,N_12857);
and U13860 (N_13860,N_12521,N_12920);
or U13861 (N_13861,N_12632,N_12038);
or U13862 (N_13862,N_12440,N_12031);
and U13863 (N_13863,N_12593,N_12450);
nand U13864 (N_13864,N_12276,N_12779);
or U13865 (N_13865,N_12808,N_12880);
nand U13866 (N_13866,N_12168,N_12918);
xor U13867 (N_13867,N_12974,N_12340);
or U13868 (N_13868,N_12828,N_12014);
or U13869 (N_13869,N_12120,N_12214);
nor U13870 (N_13870,N_12090,N_12309);
nand U13871 (N_13871,N_12141,N_12455);
or U13872 (N_13872,N_12390,N_12615);
nand U13873 (N_13873,N_12078,N_12789);
nand U13874 (N_13874,N_12404,N_12209);
and U13875 (N_13875,N_12551,N_12893);
and U13876 (N_13876,N_12838,N_12046);
and U13877 (N_13877,N_12193,N_12000);
nand U13878 (N_13878,N_12955,N_12713);
nand U13879 (N_13879,N_12596,N_12063);
or U13880 (N_13880,N_12513,N_12381);
xor U13881 (N_13881,N_12416,N_12032);
nand U13882 (N_13882,N_12480,N_12858);
and U13883 (N_13883,N_12271,N_12891);
xnor U13884 (N_13884,N_12076,N_12490);
nor U13885 (N_13885,N_12575,N_12546);
nand U13886 (N_13886,N_12878,N_12361);
nand U13887 (N_13887,N_12567,N_12628);
or U13888 (N_13888,N_12556,N_12824);
nor U13889 (N_13889,N_12087,N_12687);
xor U13890 (N_13890,N_12864,N_12341);
and U13891 (N_13891,N_12933,N_12564);
or U13892 (N_13892,N_12230,N_12947);
and U13893 (N_13893,N_12853,N_12340);
nor U13894 (N_13894,N_12043,N_12775);
nor U13895 (N_13895,N_12920,N_12612);
xor U13896 (N_13896,N_12957,N_12923);
or U13897 (N_13897,N_12464,N_12760);
and U13898 (N_13898,N_12127,N_12433);
or U13899 (N_13899,N_12229,N_12070);
or U13900 (N_13900,N_12800,N_12124);
nand U13901 (N_13901,N_12456,N_12617);
nand U13902 (N_13902,N_12724,N_12552);
nand U13903 (N_13903,N_12613,N_12808);
nor U13904 (N_13904,N_12890,N_12173);
and U13905 (N_13905,N_12089,N_12301);
and U13906 (N_13906,N_12683,N_12526);
nand U13907 (N_13907,N_12504,N_12483);
or U13908 (N_13908,N_12572,N_12621);
nand U13909 (N_13909,N_12909,N_12155);
nand U13910 (N_13910,N_12260,N_12472);
and U13911 (N_13911,N_12786,N_12623);
nand U13912 (N_13912,N_12559,N_12697);
or U13913 (N_13913,N_12029,N_12854);
xor U13914 (N_13914,N_12763,N_12439);
nand U13915 (N_13915,N_12478,N_12763);
nor U13916 (N_13916,N_12150,N_12177);
nand U13917 (N_13917,N_12305,N_12541);
and U13918 (N_13918,N_12105,N_12518);
and U13919 (N_13919,N_12799,N_12580);
nor U13920 (N_13920,N_12143,N_12353);
xor U13921 (N_13921,N_12574,N_12214);
or U13922 (N_13922,N_12823,N_12285);
or U13923 (N_13923,N_12226,N_12791);
nand U13924 (N_13924,N_12731,N_12322);
or U13925 (N_13925,N_12714,N_12225);
xnor U13926 (N_13926,N_12193,N_12190);
nand U13927 (N_13927,N_12736,N_12668);
or U13928 (N_13928,N_12056,N_12285);
nand U13929 (N_13929,N_12493,N_12564);
nand U13930 (N_13930,N_12661,N_12038);
nand U13931 (N_13931,N_12897,N_12586);
nand U13932 (N_13932,N_12111,N_12137);
xor U13933 (N_13933,N_12334,N_12716);
nor U13934 (N_13934,N_12265,N_12086);
or U13935 (N_13935,N_12287,N_12117);
or U13936 (N_13936,N_12547,N_12935);
nor U13937 (N_13937,N_12415,N_12400);
and U13938 (N_13938,N_12808,N_12587);
or U13939 (N_13939,N_12403,N_12903);
nand U13940 (N_13940,N_12426,N_12690);
nor U13941 (N_13941,N_12755,N_12162);
or U13942 (N_13942,N_12552,N_12536);
nand U13943 (N_13943,N_12980,N_12939);
and U13944 (N_13944,N_12018,N_12300);
nand U13945 (N_13945,N_12816,N_12146);
and U13946 (N_13946,N_12558,N_12944);
and U13947 (N_13947,N_12536,N_12438);
nand U13948 (N_13948,N_12740,N_12357);
and U13949 (N_13949,N_12130,N_12610);
and U13950 (N_13950,N_12715,N_12579);
and U13951 (N_13951,N_12313,N_12531);
nor U13952 (N_13952,N_12474,N_12132);
nor U13953 (N_13953,N_12274,N_12668);
or U13954 (N_13954,N_12708,N_12238);
xor U13955 (N_13955,N_12403,N_12163);
or U13956 (N_13956,N_12171,N_12627);
and U13957 (N_13957,N_12323,N_12400);
or U13958 (N_13958,N_12467,N_12369);
or U13959 (N_13959,N_12304,N_12760);
xnor U13960 (N_13960,N_12924,N_12066);
nand U13961 (N_13961,N_12685,N_12370);
and U13962 (N_13962,N_12039,N_12398);
nor U13963 (N_13963,N_12009,N_12758);
and U13964 (N_13964,N_12706,N_12541);
or U13965 (N_13965,N_12193,N_12267);
or U13966 (N_13966,N_12574,N_12955);
nand U13967 (N_13967,N_12562,N_12091);
and U13968 (N_13968,N_12099,N_12530);
xnor U13969 (N_13969,N_12368,N_12726);
and U13970 (N_13970,N_12563,N_12375);
xnor U13971 (N_13971,N_12539,N_12769);
xnor U13972 (N_13972,N_12385,N_12712);
xor U13973 (N_13973,N_12858,N_12657);
and U13974 (N_13974,N_12783,N_12263);
xor U13975 (N_13975,N_12059,N_12908);
or U13976 (N_13976,N_12973,N_12787);
or U13977 (N_13977,N_12329,N_12722);
nor U13978 (N_13978,N_12312,N_12436);
nand U13979 (N_13979,N_12508,N_12889);
nor U13980 (N_13980,N_12691,N_12665);
or U13981 (N_13981,N_12267,N_12741);
or U13982 (N_13982,N_12790,N_12576);
nor U13983 (N_13983,N_12429,N_12476);
xor U13984 (N_13984,N_12288,N_12743);
nand U13985 (N_13985,N_12272,N_12929);
or U13986 (N_13986,N_12163,N_12708);
nand U13987 (N_13987,N_12060,N_12457);
nor U13988 (N_13988,N_12308,N_12580);
nand U13989 (N_13989,N_12130,N_12465);
nand U13990 (N_13990,N_12165,N_12502);
xnor U13991 (N_13991,N_12045,N_12912);
or U13992 (N_13992,N_12694,N_12373);
or U13993 (N_13993,N_12301,N_12727);
nand U13994 (N_13994,N_12414,N_12133);
xnor U13995 (N_13995,N_12834,N_12385);
xor U13996 (N_13996,N_12738,N_12652);
nor U13997 (N_13997,N_12408,N_12252);
and U13998 (N_13998,N_12910,N_12448);
nor U13999 (N_13999,N_12635,N_12202);
and U14000 (N_14000,N_13529,N_13986);
nand U14001 (N_14001,N_13457,N_13209);
nand U14002 (N_14002,N_13689,N_13709);
or U14003 (N_14003,N_13364,N_13941);
or U14004 (N_14004,N_13748,N_13952);
nand U14005 (N_14005,N_13257,N_13517);
and U14006 (N_14006,N_13006,N_13357);
or U14007 (N_14007,N_13383,N_13452);
nand U14008 (N_14008,N_13755,N_13855);
nand U14009 (N_14009,N_13439,N_13682);
xor U14010 (N_14010,N_13353,N_13697);
nand U14011 (N_14011,N_13750,N_13976);
xnor U14012 (N_14012,N_13679,N_13226);
and U14013 (N_14013,N_13417,N_13983);
and U14014 (N_14014,N_13822,N_13639);
xor U14015 (N_14015,N_13892,N_13898);
nand U14016 (N_14016,N_13631,N_13603);
nand U14017 (N_14017,N_13445,N_13670);
xor U14018 (N_14018,N_13746,N_13740);
nand U14019 (N_14019,N_13914,N_13859);
nand U14020 (N_14020,N_13723,N_13481);
and U14021 (N_14021,N_13791,N_13165);
nand U14022 (N_14022,N_13195,N_13024);
and U14023 (N_14023,N_13212,N_13292);
nand U14024 (N_14024,N_13395,N_13358);
nor U14025 (N_14025,N_13695,N_13271);
or U14026 (N_14026,N_13554,N_13479);
nand U14027 (N_14027,N_13985,N_13034);
nand U14028 (N_14028,N_13122,N_13926);
or U14029 (N_14029,N_13132,N_13575);
nor U14030 (N_14030,N_13542,N_13798);
or U14031 (N_14031,N_13522,N_13373);
xor U14032 (N_14032,N_13907,N_13050);
xnor U14033 (N_14033,N_13728,N_13393);
nand U14034 (N_14034,N_13090,N_13704);
or U14035 (N_14035,N_13662,N_13778);
or U14036 (N_14036,N_13903,N_13675);
nor U14037 (N_14037,N_13298,N_13724);
and U14038 (N_14038,N_13375,N_13780);
nor U14039 (N_14039,N_13538,N_13945);
and U14040 (N_14040,N_13366,N_13158);
nand U14041 (N_14041,N_13912,N_13726);
or U14042 (N_14042,N_13478,N_13772);
and U14043 (N_14043,N_13063,N_13411);
or U14044 (N_14044,N_13000,N_13003);
or U14045 (N_14045,N_13541,N_13011);
nand U14046 (N_14046,N_13716,N_13207);
and U14047 (N_14047,N_13362,N_13115);
nand U14048 (N_14048,N_13534,N_13141);
or U14049 (N_14049,N_13921,N_13066);
xnor U14050 (N_14050,N_13964,N_13918);
xnor U14051 (N_14051,N_13137,N_13973);
xor U14052 (N_14052,N_13064,N_13618);
or U14053 (N_14053,N_13763,N_13727);
and U14054 (N_14054,N_13301,N_13101);
nor U14055 (N_14055,N_13518,N_13140);
nand U14056 (N_14056,N_13502,N_13228);
or U14057 (N_14057,N_13218,N_13312);
or U14058 (N_14058,N_13845,N_13749);
or U14059 (N_14059,N_13107,N_13640);
or U14060 (N_14060,N_13835,N_13203);
and U14061 (N_14061,N_13299,N_13084);
and U14062 (N_14062,N_13744,N_13787);
or U14063 (N_14063,N_13131,N_13192);
nor U14064 (N_14064,N_13832,N_13237);
or U14065 (N_14065,N_13863,N_13570);
nand U14066 (N_14066,N_13551,N_13036);
xor U14067 (N_14067,N_13110,N_13546);
nor U14068 (N_14068,N_13747,N_13255);
or U14069 (N_14069,N_13556,N_13118);
or U14070 (N_14070,N_13136,N_13611);
xor U14071 (N_14071,N_13595,N_13437);
or U14072 (N_14072,N_13114,N_13410);
xor U14073 (N_14073,N_13079,N_13632);
and U14074 (N_14074,N_13854,N_13719);
or U14075 (N_14075,N_13865,N_13974);
nand U14076 (N_14076,N_13615,N_13537);
nand U14077 (N_14077,N_13174,N_13217);
and U14078 (N_14078,N_13351,N_13069);
nand U14079 (N_14079,N_13324,N_13241);
nor U14080 (N_14080,N_13329,N_13039);
xnor U14081 (N_14081,N_13198,N_13026);
nor U14082 (N_14082,N_13499,N_13577);
xor U14083 (N_14083,N_13206,N_13049);
xnor U14084 (N_14084,N_13042,N_13380);
nor U14085 (N_14085,N_13369,N_13968);
nand U14086 (N_14086,N_13394,N_13608);
nand U14087 (N_14087,N_13055,N_13743);
xnor U14088 (N_14088,N_13497,N_13071);
xor U14089 (N_14089,N_13216,N_13360);
xnor U14090 (N_14090,N_13852,N_13438);
nor U14091 (N_14091,N_13381,N_13046);
nor U14092 (N_14092,N_13932,N_13571);
xnor U14093 (N_14093,N_13599,N_13967);
and U14094 (N_14094,N_13509,N_13978);
and U14095 (N_14095,N_13630,N_13665);
and U14096 (N_14096,N_13619,N_13593);
nor U14097 (N_14097,N_13045,N_13899);
or U14098 (N_14098,N_13935,N_13103);
nor U14099 (N_14099,N_13532,N_13947);
xnor U14100 (N_14100,N_13188,N_13955);
or U14101 (N_14101,N_13235,N_13458);
nand U14102 (N_14102,N_13247,N_13792);
or U14103 (N_14103,N_13104,N_13939);
and U14104 (N_14104,N_13475,N_13781);
or U14105 (N_14105,N_13076,N_13105);
xnor U14106 (N_14106,N_13738,N_13576);
nand U14107 (N_14107,N_13594,N_13685);
and U14108 (N_14108,N_13664,N_13225);
nor U14109 (N_14109,N_13702,N_13688);
nand U14110 (N_14110,N_13193,N_13521);
nand U14111 (N_14111,N_13233,N_13182);
xnor U14112 (N_14112,N_13923,N_13568);
xor U14113 (N_14113,N_13591,N_13988);
nand U14114 (N_14114,N_13982,N_13490);
and U14115 (N_14115,N_13672,N_13960);
and U14116 (N_14116,N_13334,N_13092);
nor U14117 (N_14117,N_13906,N_13585);
nor U14118 (N_14118,N_13184,N_13120);
nor U14119 (N_14119,N_13460,N_13562);
nor U14120 (N_14120,N_13784,N_13501);
nand U14121 (N_14121,N_13590,N_13732);
and U14122 (N_14122,N_13266,N_13229);
xor U14123 (N_14123,N_13548,N_13651);
nor U14124 (N_14124,N_13442,N_13572);
xnor U14125 (N_14125,N_13646,N_13493);
nand U14126 (N_14126,N_13937,N_13513);
nor U14127 (N_14127,N_13256,N_13302);
nor U14128 (N_14128,N_13370,N_13459);
or U14129 (N_14129,N_13290,N_13403);
nor U14130 (N_14130,N_13773,N_13809);
xnor U14131 (N_14131,N_13344,N_13837);
nand U14132 (N_14132,N_13032,N_13396);
or U14133 (N_14133,N_13453,N_13155);
or U14134 (N_14134,N_13663,N_13645);
and U14135 (N_14135,N_13963,N_13149);
or U14136 (N_14136,N_13520,N_13994);
and U14137 (N_14137,N_13346,N_13068);
nand U14138 (N_14138,N_13189,N_13965);
and U14139 (N_14139,N_13349,N_13187);
nand U14140 (N_14140,N_13087,N_13525);
nand U14141 (N_14141,N_13762,N_13082);
or U14142 (N_14142,N_13156,N_13638);
nand U14143 (N_14143,N_13721,N_13860);
xnor U14144 (N_14144,N_13836,N_13566);
and U14145 (N_14145,N_13875,N_13339);
or U14146 (N_14146,N_13074,N_13151);
nor U14147 (N_14147,N_13236,N_13494);
xor U14148 (N_14148,N_13816,N_13486);
nand U14149 (N_14149,N_13191,N_13023);
and U14150 (N_14150,N_13928,N_13461);
nor U14151 (N_14151,N_13119,N_13751);
nor U14152 (N_14152,N_13504,N_13143);
and U14153 (N_14153,N_13249,N_13589);
nand U14154 (N_14154,N_13943,N_13760);
and U14155 (N_14155,N_13356,N_13839);
nand U14156 (N_14156,N_13936,N_13678);
xor U14157 (N_14157,N_13588,N_13673);
nor U14158 (N_14158,N_13083,N_13392);
nand U14159 (N_14159,N_13909,N_13065);
and U14160 (N_14160,N_13560,N_13433);
nand U14161 (N_14161,N_13029,N_13372);
xnor U14162 (N_14162,N_13880,N_13549);
and U14163 (N_14163,N_13774,N_13205);
nor U14164 (N_14164,N_13345,N_13680);
and U14165 (N_14165,N_13861,N_13086);
or U14166 (N_14166,N_13020,N_13598);
and U14167 (N_14167,N_13954,N_13862);
nand U14168 (N_14168,N_13498,N_13031);
and U14169 (N_14169,N_13070,N_13626);
nand U14170 (N_14170,N_13950,N_13674);
nor U14171 (N_14171,N_13367,N_13268);
xor U14172 (N_14172,N_13060,N_13322);
nand U14173 (N_14173,N_13145,N_13113);
or U14174 (N_14174,N_13328,N_13843);
nor U14175 (N_14175,N_13240,N_13866);
nor U14176 (N_14176,N_13088,N_13850);
nand U14177 (N_14177,N_13765,N_13647);
nor U14178 (N_14178,N_13876,N_13758);
nand U14179 (N_14179,N_13484,N_13172);
xnor U14180 (N_14180,N_13467,N_13788);
or U14181 (N_14181,N_13223,N_13482);
nand U14182 (N_14182,N_13783,N_13095);
xnor U14183 (N_14183,N_13425,N_13842);
xor U14184 (N_14184,N_13007,N_13642);
xnor U14185 (N_14185,N_13872,N_13833);
nor U14186 (N_14186,N_13824,N_13102);
and U14187 (N_14187,N_13446,N_13934);
nor U14188 (N_14188,N_13582,N_13186);
or U14189 (N_14189,N_13014,N_13953);
nor U14190 (N_14190,N_13736,N_13530);
xor U14191 (N_14191,N_13756,N_13430);
and U14192 (N_14192,N_13879,N_13354);
nor U14193 (N_14193,N_13305,N_13896);
xor U14194 (N_14194,N_13600,N_13777);
or U14195 (N_14195,N_13869,N_13797);
nand U14196 (N_14196,N_13179,N_13279);
and U14197 (N_14197,N_13735,N_13098);
xnor U14198 (N_14198,N_13733,N_13013);
nand U14199 (N_14199,N_13807,N_13818);
nor U14200 (N_14200,N_13359,N_13831);
nand U14201 (N_14201,N_13810,N_13146);
nand U14202 (N_14202,N_13966,N_13867);
and U14203 (N_14203,N_13224,N_13757);
or U14204 (N_14204,N_13480,N_13227);
and U14205 (N_14205,N_13821,N_13707);
or U14206 (N_14206,N_13243,N_13905);
or U14207 (N_14207,N_13160,N_13303);
nand U14208 (N_14208,N_13270,N_13093);
xor U14209 (N_14209,N_13667,N_13213);
xor U14210 (N_14210,N_13164,N_13462);
or U14211 (N_14211,N_13483,N_13385);
nand U14212 (N_14212,N_13715,N_13340);
nand U14213 (N_14213,N_13668,N_13379);
nor U14214 (N_14214,N_13676,N_13081);
nand U14215 (N_14215,N_13288,N_13691);
and U14216 (N_14216,N_13811,N_13776);
and U14217 (N_14217,N_13620,N_13979);
nand U14218 (N_14218,N_13157,N_13434);
and U14219 (N_14219,N_13489,N_13264);
nand U14220 (N_14220,N_13913,N_13658);
and U14221 (N_14221,N_13782,N_13725);
nor U14222 (N_14222,N_13469,N_13201);
nor U14223 (N_14223,N_13769,N_13210);
nand U14224 (N_14224,N_13406,N_13565);
nand U14225 (N_14225,N_13655,N_13150);
nand U14226 (N_14226,N_13830,N_13038);
nand U14227 (N_14227,N_13730,N_13002);
nor U14228 (N_14228,N_13258,N_13786);
or U14229 (N_14229,N_13190,N_13316);
and U14230 (N_14230,N_13096,N_13687);
xnor U14231 (N_14231,N_13610,N_13993);
and U14232 (N_14232,N_13827,N_13882);
or U14233 (N_14233,N_13717,N_13705);
and U14234 (N_14234,N_13503,N_13550);
and U14235 (N_14235,N_13848,N_13838);
nand U14236 (N_14236,N_13222,N_13106);
and U14237 (N_14237,N_13531,N_13286);
xnor U14238 (N_14238,N_13016,N_13643);
nor U14239 (N_14239,N_13699,N_13168);
or U14240 (N_14240,N_13564,N_13901);
or U14241 (N_14241,N_13825,N_13614);
xor U14242 (N_14242,N_13309,N_13408);
or U14243 (N_14243,N_13500,N_13443);
or U14244 (N_14244,N_13278,N_13251);
or U14245 (N_14245,N_13547,N_13390);
nor U14246 (N_14246,N_13857,N_13789);
nand U14247 (N_14247,N_13890,N_13111);
and U14248 (N_14248,N_13826,N_13265);
and U14249 (N_14249,N_13720,N_13922);
nor U14250 (N_14250,N_13802,N_13931);
xor U14251 (N_14251,N_13180,N_13904);
nand U14252 (N_14252,N_13327,N_13183);
or U14253 (N_14253,N_13874,N_13269);
and U14254 (N_14254,N_13634,N_13061);
or U14255 (N_14255,N_13121,N_13887);
xnor U14256 (N_14256,N_13378,N_13561);
xor U14257 (N_14257,N_13819,N_13753);
nor U14258 (N_14258,N_13167,N_13741);
nand U14259 (N_14259,N_13371,N_13488);
nand U14260 (N_14260,N_13677,N_13796);
nand U14261 (N_14261,N_13515,N_13424);
nor U14262 (N_14262,N_13889,N_13075);
nor U14263 (N_14263,N_13109,N_13181);
and U14264 (N_14264,N_13427,N_13628);
xnor U14265 (N_14265,N_13051,N_13545);
and U14266 (N_14266,N_13621,N_13972);
or U14267 (N_14267,N_13771,N_13812);
nand U14268 (N_14268,N_13464,N_13980);
xnor U14269 (N_14269,N_13117,N_13868);
and U14270 (N_14270,N_13078,N_13250);
xnor U14271 (N_14271,N_13731,N_13397);
and U14272 (N_14272,N_13536,N_13466);
nor U14273 (N_14273,N_13770,N_13262);
nand U14274 (N_14274,N_13514,N_13019);
nand U14275 (N_14275,N_13130,N_13178);
nand U14276 (N_14276,N_13559,N_13535);
nand U14277 (N_14277,N_13660,N_13737);
or U14278 (N_14278,N_13281,N_13888);
nor U14279 (N_14279,N_13388,N_13350);
nand U14280 (N_14280,N_13477,N_13295);
nor U14281 (N_14281,N_13124,N_13175);
nand U14282 (N_14282,N_13592,N_13745);
or U14283 (N_14283,N_13790,N_13176);
nand U14284 (N_14284,N_13659,N_13202);
and U14285 (N_14285,N_13315,N_13277);
nor U14286 (N_14286,N_13808,N_13300);
nor U14287 (N_14287,N_13170,N_13123);
xnor U14288 (N_14288,N_13806,N_13920);
and U14289 (N_14289,N_13873,N_13558);
and U14290 (N_14290,N_13929,N_13048);
nand U14291 (N_14291,N_13420,N_13942);
xor U14292 (N_14292,N_13915,N_13847);
xor U14293 (N_14293,N_13169,N_13470);
nor U14294 (N_14294,N_13455,N_13764);
nand U14295 (N_14295,N_13597,N_13519);
nand U14296 (N_14296,N_13259,N_13239);
xor U14297 (N_14297,N_13230,N_13030);
nor U14298 (N_14298,N_13428,N_13254);
xor U14299 (N_14299,N_13204,N_13989);
xnor U14300 (N_14300,N_13047,N_13219);
nand U14301 (N_14301,N_13584,N_13895);
and U14302 (N_14302,N_13948,N_13636);
nand U14303 (N_14303,N_13871,N_13563);
and U14304 (N_14304,N_13252,N_13690);
xor U14305 (N_14305,N_13449,N_13194);
nand U14306 (N_14306,N_13799,N_13841);
xnor U14307 (N_14307,N_13512,N_13581);
nor U14308 (N_14308,N_13524,N_13919);
and U14309 (N_14309,N_13996,N_13402);
or U14310 (N_14310,N_13569,N_13669);
nand U14311 (N_14311,N_13692,N_13984);
and U14312 (N_14312,N_13331,N_13293);
nor U14313 (N_14313,N_13804,N_13275);
xnor U14314 (N_14314,N_13714,N_13413);
or U14315 (N_14315,N_13991,N_13527);
nor U14316 (N_14316,N_13294,N_13418);
nand U14317 (N_14317,N_13800,N_13080);
nand U14318 (N_14318,N_13035,N_13507);
or U14319 (N_14319,N_13633,N_13429);
xnor U14320 (N_14320,N_13846,N_13607);
or U14321 (N_14321,N_13085,N_13089);
xnor U14322 (N_14322,N_13539,N_13291);
or U14323 (N_14323,N_13508,N_13694);
nand U14324 (N_14324,N_13422,N_13077);
or U14325 (N_14325,N_13058,N_13033);
and U14326 (N_14326,N_13606,N_13648);
and U14327 (N_14327,N_13491,N_13352);
and U14328 (N_14328,N_13917,N_13883);
nand U14329 (N_14329,N_13511,N_13273);
xnor U14330 (N_14330,N_13612,N_13742);
nor U14331 (N_14331,N_13289,N_13635);
or U14332 (N_14332,N_13557,N_13405);
nand U14333 (N_14333,N_13056,N_13552);
nor U14334 (N_14334,N_13336,N_13766);
nand U14335 (N_14335,N_13423,N_13386);
nor U14336 (N_14336,N_13173,N_13400);
and U14337 (N_14337,N_13116,N_13355);
nor U14338 (N_14338,N_13649,N_13220);
or U14339 (N_14339,N_13037,N_13998);
nor U14340 (N_14340,N_13997,N_13686);
or U14341 (N_14341,N_13543,N_13981);
xnor U14342 (N_14342,N_13125,N_13759);
and U14343 (N_14343,N_13496,N_13043);
xor U14344 (N_14344,N_13573,N_13706);
and U14345 (N_14345,N_13959,N_13404);
nor U14346 (N_14346,N_13415,N_13886);
xnor U14347 (N_14347,N_13465,N_13091);
xor U14348 (N_14348,N_13933,N_13267);
and U14349 (N_14349,N_13199,N_13384);
nand U14350 (N_14350,N_13703,N_13701);
nand U14351 (N_14351,N_13399,N_13849);
nor U14352 (N_14352,N_13793,N_13656);
xnor U14353 (N_14353,N_13574,N_13062);
and U14354 (N_14354,N_13473,N_13661);
nand U14355 (N_14355,N_13368,N_13779);
or U14356 (N_14356,N_13700,N_13244);
or U14357 (N_14357,N_13280,N_13326);
nand U14358 (N_14358,N_13341,N_13492);
or U14359 (N_14359,N_13127,N_13314);
nor U14360 (N_14360,N_13285,N_13197);
nand U14361 (N_14361,N_13944,N_13583);
xor U14362 (N_14362,N_13987,N_13159);
or U14363 (N_14363,N_13977,N_13834);
nor U14364 (N_14364,N_13739,N_13946);
nor U14365 (N_14365,N_13586,N_13625);
nor U14366 (N_14366,N_13153,N_13208);
and U14367 (N_14367,N_13363,N_13310);
xor U14368 (N_14368,N_13343,N_13185);
nor U14369 (N_14369,N_13495,N_13803);
or U14370 (N_14370,N_13067,N_13696);
and U14371 (N_14371,N_13940,N_13617);
xnor U14372 (N_14372,N_13870,N_13698);
xor U14373 (N_14373,N_13108,N_13468);
and U14374 (N_14374,N_13627,N_13580);
xor U14375 (N_14375,N_13094,N_13387);
nand U14376 (N_14376,N_13604,N_13112);
nand U14377 (N_14377,N_13684,N_13021);
nand U14378 (N_14378,N_13284,N_13053);
or U14379 (N_14379,N_13601,N_13485);
xor U14380 (N_14380,N_13908,N_13801);
or U14381 (N_14381,N_13949,N_13001);
nor U14382 (N_14382,N_13487,N_13794);
and U14383 (N_14383,N_13938,N_13337);
or U14384 (N_14384,N_13320,N_13957);
xnor U14385 (N_14385,N_13318,N_13272);
or U14386 (N_14386,N_13924,N_13693);
and U14387 (N_14387,N_13805,N_13450);
or U14388 (N_14388,N_13711,N_13958);
and U14389 (N_14389,N_13099,N_13474);
or U14390 (N_14390,N_13260,N_13377);
and U14391 (N_14391,N_13856,N_13283);
nand U14392 (N_14392,N_13444,N_13040);
nand U14393 (N_14393,N_13729,N_13814);
or U14394 (N_14394,N_13313,N_13374);
nor U14395 (N_14395,N_13894,N_13027);
or U14396 (N_14396,N_13100,N_13995);
nor U14397 (N_14397,N_13022,N_13059);
or U14398 (N_14398,N_13657,N_13897);
nor U14399 (N_14399,N_13927,N_13376);
xor U14400 (N_14400,N_13414,N_13829);
nand U14401 (N_14401,N_13505,N_13962);
nor U14402 (N_14402,N_13523,N_13813);
nor U14403 (N_14403,N_13454,N_13555);
and U14404 (N_14404,N_13348,N_13718);
nor U14405 (N_14405,N_13416,N_13389);
or U14406 (N_14406,N_13162,N_13884);
and U14407 (N_14407,N_13891,N_13602);
and U14408 (N_14408,N_13332,N_13544);
nand U14409 (N_14409,N_13881,N_13163);
or U14410 (N_14410,N_13054,N_13274);
nand U14411 (N_14411,N_13005,N_13910);
or U14412 (N_14412,N_13767,N_13330);
xor U14413 (N_14413,N_13307,N_13177);
or U14414 (N_14414,N_13166,N_13238);
nand U14415 (N_14415,N_13161,N_13623);
or U14416 (N_14416,N_13347,N_13009);
or U14417 (N_14417,N_13154,N_13893);
nand U14418 (N_14418,N_13231,N_13421);
and U14419 (N_14419,N_13456,N_13282);
xnor U14420 (N_14420,N_13133,N_13605);
and U14421 (N_14421,N_13025,N_13900);
nand U14422 (N_14422,N_13671,N_13681);
xnor U14423 (N_14423,N_13015,N_13097);
and U14424 (N_14424,N_13877,N_13072);
xor U14425 (N_14425,N_13992,N_13409);
xnor U14426 (N_14426,N_13010,N_13510);
and U14427 (N_14427,N_13925,N_13472);
and U14428 (N_14428,N_13683,N_13956);
xor U14429 (N_14429,N_13419,N_13596);
nand U14430 (N_14430,N_13142,N_13578);
xor U14431 (N_14431,N_13028,N_13232);
or U14432 (N_14432,N_13815,N_13234);
xnor U14433 (N_14433,N_13644,N_13253);
xor U14434 (N_14434,N_13245,N_13448);
or U14435 (N_14435,N_13930,N_13044);
nand U14436 (N_14436,N_13436,N_13817);
nor U14437 (N_14437,N_13975,N_13840);
and U14438 (N_14438,N_13752,N_13629);
nand U14439 (N_14439,N_13382,N_13306);
or U14440 (N_14440,N_13311,N_13785);
or U14441 (N_14441,N_13248,N_13654);
and U14442 (N_14442,N_13325,N_13135);
xor U14443 (N_14443,N_13317,N_13533);
nand U14444 (N_14444,N_13319,N_13221);
and U14445 (N_14445,N_13795,N_13057);
or U14446 (N_14446,N_13553,N_13171);
and U14447 (N_14447,N_13018,N_13214);
and U14448 (N_14448,N_13435,N_13653);
or U14449 (N_14449,N_13622,N_13471);
and U14450 (N_14450,N_13969,N_13878);
and U14451 (N_14451,N_13246,N_13323);
and U14452 (N_14452,N_13853,N_13754);
nand U14453 (N_14453,N_13858,N_13333);
xnor U14454 (N_14454,N_13616,N_13579);
nor U14455 (N_14455,N_13722,N_13708);
or U14456 (N_14456,N_13641,N_13276);
nand U14457 (N_14457,N_13526,N_13304);
and U14458 (N_14458,N_13263,N_13666);
nand U14459 (N_14459,N_13823,N_13287);
and U14460 (N_14460,N_13447,N_13012);
or U14461 (N_14461,N_13775,N_13540);
nor U14462 (N_14462,N_13261,N_13851);
nor U14463 (N_14463,N_13321,N_13008);
and U14464 (N_14464,N_13999,N_13147);
nor U14465 (N_14465,N_13139,N_13391);
or U14466 (N_14466,N_13308,N_13609);
nor U14467 (N_14467,N_13134,N_13426);
or U14468 (N_14468,N_13637,N_13242);
or U14469 (N_14469,N_13463,N_13587);
nand U14470 (N_14470,N_13431,N_13970);
and U14471 (N_14471,N_13361,N_13129);
and U14472 (N_14472,N_13624,N_13451);
or U14473 (N_14473,N_13844,N_13916);
nand U14474 (N_14474,N_13200,N_13017);
xor U14475 (N_14475,N_13296,N_13407);
nor U14476 (N_14476,N_13073,N_13398);
and U14477 (N_14477,N_13516,N_13148);
and U14478 (N_14478,N_13211,N_13528);
or U14479 (N_14479,N_13885,N_13004);
nand U14480 (N_14480,N_13820,N_13432);
or U14481 (N_14481,N_13650,N_13567);
xnor U14482 (N_14482,N_13713,N_13412);
xor U14483 (N_14483,N_13128,N_13126);
nor U14484 (N_14484,N_13951,N_13710);
xor U14485 (N_14485,N_13144,N_13041);
or U14486 (N_14486,N_13768,N_13138);
and U14487 (N_14487,N_13971,N_13297);
nor U14488 (N_14488,N_13152,N_13215);
xor U14489 (N_14489,N_13342,N_13734);
or U14490 (N_14490,N_13712,N_13990);
and U14491 (N_14491,N_13902,N_13401);
nand U14492 (N_14492,N_13911,N_13961);
or U14493 (N_14493,N_13335,N_13052);
and U14494 (N_14494,N_13476,N_13613);
or U14495 (N_14495,N_13864,N_13338);
and U14496 (N_14496,N_13828,N_13365);
nand U14497 (N_14497,N_13440,N_13761);
or U14498 (N_14498,N_13506,N_13196);
xor U14499 (N_14499,N_13652,N_13441);
xnor U14500 (N_14500,N_13324,N_13149);
or U14501 (N_14501,N_13084,N_13991);
xnor U14502 (N_14502,N_13643,N_13164);
xnor U14503 (N_14503,N_13225,N_13703);
and U14504 (N_14504,N_13947,N_13691);
nand U14505 (N_14505,N_13353,N_13035);
or U14506 (N_14506,N_13635,N_13403);
and U14507 (N_14507,N_13732,N_13525);
nand U14508 (N_14508,N_13493,N_13283);
or U14509 (N_14509,N_13378,N_13878);
nand U14510 (N_14510,N_13046,N_13123);
or U14511 (N_14511,N_13037,N_13720);
xnor U14512 (N_14512,N_13685,N_13052);
or U14513 (N_14513,N_13557,N_13654);
xor U14514 (N_14514,N_13099,N_13612);
or U14515 (N_14515,N_13043,N_13189);
xor U14516 (N_14516,N_13722,N_13948);
and U14517 (N_14517,N_13507,N_13858);
xor U14518 (N_14518,N_13385,N_13650);
nor U14519 (N_14519,N_13696,N_13035);
nand U14520 (N_14520,N_13727,N_13181);
nand U14521 (N_14521,N_13969,N_13599);
and U14522 (N_14522,N_13028,N_13557);
and U14523 (N_14523,N_13495,N_13150);
xor U14524 (N_14524,N_13068,N_13156);
nand U14525 (N_14525,N_13907,N_13332);
nor U14526 (N_14526,N_13599,N_13901);
or U14527 (N_14527,N_13415,N_13345);
nand U14528 (N_14528,N_13687,N_13244);
nand U14529 (N_14529,N_13131,N_13263);
nor U14530 (N_14530,N_13509,N_13497);
nor U14531 (N_14531,N_13130,N_13585);
nand U14532 (N_14532,N_13046,N_13947);
and U14533 (N_14533,N_13853,N_13997);
nand U14534 (N_14534,N_13689,N_13732);
or U14535 (N_14535,N_13392,N_13061);
nor U14536 (N_14536,N_13711,N_13370);
or U14537 (N_14537,N_13476,N_13423);
xor U14538 (N_14538,N_13327,N_13779);
and U14539 (N_14539,N_13077,N_13963);
xor U14540 (N_14540,N_13530,N_13977);
and U14541 (N_14541,N_13362,N_13490);
nand U14542 (N_14542,N_13123,N_13059);
nor U14543 (N_14543,N_13139,N_13378);
or U14544 (N_14544,N_13442,N_13186);
xnor U14545 (N_14545,N_13900,N_13185);
nand U14546 (N_14546,N_13558,N_13709);
and U14547 (N_14547,N_13917,N_13445);
and U14548 (N_14548,N_13628,N_13282);
or U14549 (N_14549,N_13053,N_13610);
nand U14550 (N_14550,N_13924,N_13083);
nor U14551 (N_14551,N_13167,N_13102);
and U14552 (N_14552,N_13232,N_13472);
or U14553 (N_14553,N_13631,N_13814);
nor U14554 (N_14554,N_13876,N_13862);
or U14555 (N_14555,N_13252,N_13827);
nand U14556 (N_14556,N_13938,N_13126);
nor U14557 (N_14557,N_13657,N_13462);
and U14558 (N_14558,N_13494,N_13654);
and U14559 (N_14559,N_13855,N_13524);
nor U14560 (N_14560,N_13801,N_13790);
xnor U14561 (N_14561,N_13396,N_13566);
and U14562 (N_14562,N_13564,N_13328);
xnor U14563 (N_14563,N_13601,N_13591);
nor U14564 (N_14564,N_13435,N_13219);
and U14565 (N_14565,N_13457,N_13847);
and U14566 (N_14566,N_13368,N_13160);
xor U14567 (N_14567,N_13962,N_13006);
or U14568 (N_14568,N_13544,N_13092);
or U14569 (N_14569,N_13627,N_13317);
nand U14570 (N_14570,N_13466,N_13152);
nand U14571 (N_14571,N_13776,N_13269);
nor U14572 (N_14572,N_13824,N_13621);
nor U14573 (N_14573,N_13538,N_13588);
or U14574 (N_14574,N_13671,N_13289);
or U14575 (N_14575,N_13928,N_13129);
and U14576 (N_14576,N_13922,N_13635);
or U14577 (N_14577,N_13834,N_13798);
nand U14578 (N_14578,N_13514,N_13008);
nand U14579 (N_14579,N_13999,N_13706);
and U14580 (N_14580,N_13100,N_13894);
xnor U14581 (N_14581,N_13682,N_13258);
and U14582 (N_14582,N_13791,N_13067);
nor U14583 (N_14583,N_13250,N_13926);
nand U14584 (N_14584,N_13587,N_13404);
nand U14585 (N_14585,N_13651,N_13501);
xnor U14586 (N_14586,N_13953,N_13580);
and U14587 (N_14587,N_13210,N_13858);
nand U14588 (N_14588,N_13881,N_13204);
nor U14589 (N_14589,N_13311,N_13096);
nor U14590 (N_14590,N_13492,N_13343);
xnor U14591 (N_14591,N_13316,N_13135);
nand U14592 (N_14592,N_13883,N_13562);
and U14593 (N_14593,N_13639,N_13934);
or U14594 (N_14594,N_13363,N_13081);
nand U14595 (N_14595,N_13447,N_13836);
nor U14596 (N_14596,N_13370,N_13588);
and U14597 (N_14597,N_13214,N_13550);
and U14598 (N_14598,N_13146,N_13463);
and U14599 (N_14599,N_13286,N_13516);
nor U14600 (N_14600,N_13651,N_13191);
nor U14601 (N_14601,N_13135,N_13582);
or U14602 (N_14602,N_13439,N_13797);
nor U14603 (N_14603,N_13102,N_13547);
nand U14604 (N_14604,N_13420,N_13241);
or U14605 (N_14605,N_13821,N_13266);
or U14606 (N_14606,N_13764,N_13403);
nand U14607 (N_14607,N_13134,N_13558);
nand U14608 (N_14608,N_13565,N_13672);
nand U14609 (N_14609,N_13731,N_13049);
and U14610 (N_14610,N_13091,N_13836);
or U14611 (N_14611,N_13494,N_13851);
xnor U14612 (N_14612,N_13070,N_13190);
xor U14613 (N_14613,N_13457,N_13758);
nand U14614 (N_14614,N_13249,N_13659);
nor U14615 (N_14615,N_13174,N_13442);
nand U14616 (N_14616,N_13649,N_13943);
or U14617 (N_14617,N_13856,N_13157);
nand U14618 (N_14618,N_13022,N_13844);
nand U14619 (N_14619,N_13487,N_13983);
xor U14620 (N_14620,N_13777,N_13703);
xor U14621 (N_14621,N_13002,N_13868);
nand U14622 (N_14622,N_13804,N_13237);
nor U14623 (N_14623,N_13182,N_13655);
and U14624 (N_14624,N_13283,N_13550);
and U14625 (N_14625,N_13825,N_13443);
nor U14626 (N_14626,N_13049,N_13808);
or U14627 (N_14627,N_13614,N_13312);
xor U14628 (N_14628,N_13860,N_13097);
nand U14629 (N_14629,N_13524,N_13842);
xor U14630 (N_14630,N_13782,N_13249);
and U14631 (N_14631,N_13201,N_13164);
and U14632 (N_14632,N_13046,N_13979);
or U14633 (N_14633,N_13131,N_13295);
nor U14634 (N_14634,N_13067,N_13061);
or U14635 (N_14635,N_13371,N_13184);
or U14636 (N_14636,N_13396,N_13027);
nand U14637 (N_14637,N_13284,N_13119);
xnor U14638 (N_14638,N_13064,N_13436);
or U14639 (N_14639,N_13483,N_13861);
nor U14640 (N_14640,N_13089,N_13585);
or U14641 (N_14641,N_13166,N_13788);
nor U14642 (N_14642,N_13039,N_13046);
or U14643 (N_14643,N_13543,N_13808);
or U14644 (N_14644,N_13964,N_13808);
nand U14645 (N_14645,N_13496,N_13598);
or U14646 (N_14646,N_13298,N_13431);
nand U14647 (N_14647,N_13697,N_13646);
xnor U14648 (N_14648,N_13870,N_13967);
nand U14649 (N_14649,N_13150,N_13615);
nor U14650 (N_14650,N_13321,N_13715);
nor U14651 (N_14651,N_13943,N_13624);
nand U14652 (N_14652,N_13993,N_13869);
and U14653 (N_14653,N_13957,N_13216);
or U14654 (N_14654,N_13563,N_13695);
and U14655 (N_14655,N_13900,N_13883);
or U14656 (N_14656,N_13331,N_13861);
nand U14657 (N_14657,N_13527,N_13721);
xnor U14658 (N_14658,N_13694,N_13855);
or U14659 (N_14659,N_13645,N_13736);
or U14660 (N_14660,N_13815,N_13210);
nor U14661 (N_14661,N_13495,N_13366);
nand U14662 (N_14662,N_13513,N_13922);
xor U14663 (N_14663,N_13700,N_13239);
or U14664 (N_14664,N_13115,N_13147);
nand U14665 (N_14665,N_13525,N_13043);
nand U14666 (N_14666,N_13769,N_13692);
nand U14667 (N_14667,N_13779,N_13004);
nor U14668 (N_14668,N_13473,N_13045);
xor U14669 (N_14669,N_13092,N_13529);
xor U14670 (N_14670,N_13605,N_13625);
xor U14671 (N_14671,N_13841,N_13742);
xor U14672 (N_14672,N_13120,N_13589);
nor U14673 (N_14673,N_13770,N_13106);
and U14674 (N_14674,N_13156,N_13126);
nor U14675 (N_14675,N_13350,N_13051);
and U14676 (N_14676,N_13776,N_13649);
or U14677 (N_14677,N_13399,N_13453);
or U14678 (N_14678,N_13149,N_13457);
nor U14679 (N_14679,N_13102,N_13335);
nand U14680 (N_14680,N_13004,N_13536);
or U14681 (N_14681,N_13848,N_13258);
or U14682 (N_14682,N_13437,N_13506);
xnor U14683 (N_14683,N_13462,N_13357);
nor U14684 (N_14684,N_13150,N_13018);
nand U14685 (N_14685,N_13988,N_13487);
nand U14686 (N_14686,N_13844,N_13459);
nor U14687 (N_14687,N_13239,N_13121);
nor U14688 (N_14688,N_13430,N_13814);
nand U14689 (N_14689,N_13688,N_13400);
nand U14690 (N_14690,N_13594,N_13821);
nor U14691 (N_14691,N_13638,N_13228);
and U14692 (N_14692,N_13796,N_13843);
nand U14693 (N_14693,N_13043,N_13317);
and U14694 (N_14694,N_13275,N_13835);
nor U14695 (N_14695,N_13298,N_13964);
nor U14696 (N_14696,N_13557,N_13691);
and U14697 (N_14697,N_13616,N_13840);
xor U14698 (N_14698,N_13607,N_13035);
and U14699 (N_14699,N_13586,N_13990);
nor U14700 (N_14700,N_13428,N_13207);
and U14701 (N_14701,N_13064,N_13341);
and U14702 (N_14702,N_13513,N_13184);
and U14703 (N_14703,N_13740,N_13593);
nand U14704 (N_14704,N_13647,N_13613);
nand U14705 (N_14705,N_13206,N_13379);
nor U14706 (N_14706,N_13846,N_13256);
and U14707 (N_14707,N_13961,N_13665);
or U14708 (N_14708,N_13551,N_13179);
nor U14709 (N_14709,N_13630,N_13994);
nand U14710 (N_14710,N_13805,N_13698);
or U14711 (N_14711,N_13997,N_13359);
and U14712 (N_14712,N_13156,N_13528);
nand U14713 (N_14713,N_13013,N_13936);
nand U14714 (N_14714,N_13135,N_13214);
nand U14715 (N_14715,N_13864,N_13363);
xnor U14716 (N_14716,N_13736,N_13808);
or U14717 (N_14717,N_13588,N_13237);
and U14718 (N_14718,N_13980,N_13078);
and U14719 (N_14719,N_13954,N_13680);
nor U14720 (N_14720,N_13635,N_13282);
nand U14721 (N_14721,N_13352,N_13490);
xnor U14722 (N_14722,N_13098,N_13836);
nand U14723 (N_14723,N_13211,N_13566);
and U14724 (N_14724,N_13318,N_13922);
nand U14725 (N_14725,N_13405,N_13162);
or U14726 (N_14726,N_13127,N_13571);
nor U14727 (N_14727,N_13972,N_13292);
nor U14728 (N_14728,N_13438,N_13305);
and U14729 (N_14729,N_13699,N_13777);
nor U14730 (N_14730,N_13356,N_13949);
or U14731 (N_14731,N_13104,N_13247);
nand U14732 (N_14732,N_13970,N_13756);
xnor U14733 (N_14733,N_13738,N_13438);
xnor U14734 (N_14734,N_13760,N_13438);
nor U14735 (N_14735,N_13003,N_13767);
nor U14736 (N_14736,N_13103,N_13958);
xor U14737 (N_14737,N_13661,N_13937);
or U14738 (N_14738,N_13193,N_13060);
nand U14739 (N_14739,N_13694,N_13437);
nor U14740 (N_14740,N_13080,N_13790);
nor U14741 (N_14741,N_13043,N_13307);
nor U14742 (N_14742,N_13476,N_13207);
and U14743 (N_14743,N_13518,N_13331);
nor U14744 (N_14744,N_13300,N_13772);
nor U14745 (N_14745,N_13818,N_13257);
nand U14746 (N_14746,N_13915,N_13793);
or U14747 (N_14747,N_13791,N_13377);
nand U14748 (N_14748,N_13367,N_13808);
nor U14749 (N_14749,N_13530,N_13555);
xor U14750 (N_14750,N_13818,N_13451);
and U14751 (N_14751,N_13425,N_13642);
nor U14752 (N_14752,N_13642,N_13271);
and U14753 (N_14753,N_13606,N_13617);
and U14754 (N_14754,N_13339,N_13678);
and U14755 (N_14755,N_13843,N_13043);
xnor U14756 (N_14756,N_13917,N_13533);
nor U14757 (N_14757,N_13091,N_13853);
or U14758 (N_14758,N_13402,N_13425);
or U14759 (N_14759,N_13484,N_13933);
nor U14760 (N_14760,N_13418,N_13257);
and U14761 (N_14761,N_13771,N_13669);
nor U14762 (N_14762,N_13944,N_13614);
and U14763 (N_14763,N_13056,N_13081);
or U14764 (N_14764,N_13984,N_13373);
nand U14765 (N_14765,N_13357,N_13113);
nand U14766 (N_14766,N_13798,N_13073);
or U14767 (N_14767,N_13495,N_13572);
and U14768 (N_14768,N_13091,N_13064);
nor U14769 (N_14769,N_13502,N_13827);
or U14770 (N_14770,N_13072,N_13903);
nor U14771 (N_14771,N_13802,N_13423);
nor U14772 (N_14772,N_13938,N_13919);
nor U14773 (N_14773,N_13458,N_13493);
nand U14774 (N_14774,N_13923,N_13861);
xor U14775 (N_14775,N_13340,N_13316);
nand U14776 (N_14776,N_13656,N_13197);
nor U14777 (N_14777,N_13036,N_13344);
and U14778 (N_14778,N_13193,N_13817);
and U14779 (N_14779,N_13167,N_13190);
or U14780 (N_14780,N_13829,N_13167);
or U14781 (N_14781,N_13615,N_13840);
or U14782 (N_14782,N_13212,N_13180);
and U14783 (N_14783,N_13569,N_13740);
and U14784 (N_14784,N_13634,N_13138);
or U14785 (N_14785,N_13245,N_13492);
nand U14786 (N_14786,N_13311,N_13753);
or U14787 (N_14787,N_13662,N_13710);
nand U14788 (N_14788,N_13156,N_13339);
nand U14789 (N_14789,N_13580,N_13592);
or U14790 (N_14790,N_13613,N_13299);
and U14791 (N_14791,N_13074,N_13623);
or U14792 (N_14792,N_13495,N_13590);
and U14793 (N_14793,N_13472,N_13150);
or U14794 (N_14794,N_13759,N_13672);
nor U14795 (N_14795,N_13165,N_13486);
or U14796 (N_14796,N_13027,N_13251);
and U14797 (N_14797,N_13637,N_13669);
and U14798 (N_14798,N_13057,N_13740);
xor U14799 (N_14799,N_13572,N_13240);
or U14800 (N_14800,N_13298,N_13797);
xor U14801 (N_14801,N_13734,N_13996);
or U14802 (N_14802,N_13397,N_13816);
nand U14803 (N_14803,N_13093,N_13148);
nand U14804 (N_14804,N_13141,N_13175);
or U14805 (N_14805,N_13559,N_13002);
nor U14806 (N_14806,N_13192,N_13744);
or U14807 (N_14807,N_13190,N_13047);
xnor U14808 (N_14808,N_13054,N_13065);
nor U14809 (N_14809,N_13269,N_13369);
and U14810 (N_14810,N_13724,N_13951);
and U14811 (N_14811,N_13837,N_13438);
xnor U14812 (N_14812,N_13635,N_13534);
and U14813 (N_14813,N_13532,N_13829);
or U14814 (N_14814,N_13046,N_13205);
or U14815 (N_14815,N_13946,N_13306);
and U14816 (N_14816,N_13796,N_13685);
or U14817 (N_14817,N_13652,N_13290);
or U14818 (N_14818,N_13603,N_13103);
nor U14819 (N_14819,N_13844,N_13177);
nor U14820 (N_14820,N_13343,N_13348);
and U14821 (N_14821,N_13266,N_13877);
xnor U14822 (N_14822,N_13408,N_13834);
and U14823 (N_14823,N_13785,N_13880);
nand U14824 (N_14824,N_13558,N_13150);
nand U14825 (N_14825,N_13560,N_13283);
and U14826 (N_14826,N_13450,N_13208);
or U14827 (N_14827,N_13260,N_13877);
xnor U14828 (N_14828,N_13253,N_13040);
or U14829 (N_14829,N_13982,N_13977);
nor U14830 (N_14830,N_13218,N_13493);
xnor U14831 (N_14831,N_13131,N_13576);
nor U14832 (N_14832,N_13295,N_13014);
nor U14833 (N_14833,N_13322,N_13833);
nand U14834 (N_14834,N_13299,N_13573);
and U14835 (N_14835,N_13720,N_13497);
nand U14836 (N_14836,N_13707,N_13567);
nor U14837 (N_14837,N_13945,N_13061);
xor U14838 (N_14838,N_13750,N_13930);
xnor U14839 (N_14839,N_13765,N_13412);
or U14840 (N_14840,N_13617,N_13189);
and U14841 (N_14841,N_13212,N_13107);
xor U14842 (N_14842,N_13850,N_13992);
nor U14843 (N_14843,N_13233,N_13121);
nor U14844 (N_14844,N_13393,N_13773);
and U14845 (N_14845,N_13442,N_13947);
and U14846 (N_14846,N_13006,N_13735);
and U14847 (N_14847,N_13492,N_13148);
xnor U14848 (N_14848,N_13846,N_13115);
xor U14849 (N_14849,N_13321,N_13878);
xor U14850 (N_14850,N_13849,N_13129);
xor U14851 (N_14851,N_13637,N_13941);
nor U14852 (N_14852,N_13027,N_13243);
xor U14853 (N_14853,N_13094,N_13345);
nor U14854 (N_14854,N_13112,N_13735);
xor U14855 (N_14855,N_13667,N_13233);
nor U14856 (N_14856,N_13109,N_13558);
xor U14857 (N_14857,N_13048,N_13889);
and U14858 (N_14858,N_13679,N_13479);
and U14859 (N_14859,N_13459,N_13245);
or U14860 (N_14860,N_13154,N_13678);
nand U14861 (N_14861,N_13389,N_13320);
and U14862 (N_14862,N_13851,N_13366);
xor U14863 (N_14863,N_13054,N_13594);
xnor U14864 (N_14864,N_13021,N_13843);
or U14865 (N_14865,N_13994,N_13366);
nor U14866 (N_14866,N_13255,N_13751);
or U14867 (N_14867,N_13099,N_13273);
nand U14868 (N_14868,N_13365,N_13525);
and U14869 (N_14869,N_13931,N_13978);
xnor U14870 (N_14870,N_13533,N_13508);
nand U14871 (N_14871,N_13256,N_13391);
xnor U14872 (N_14872,N_13981,N_13090);
xor U14873 (N_14873,N_13530,N_13178);
or U14874 (N_14874,N_13616,N_13224);
nor U14875 (N_14875,N_13106,N_13801);
nor U14876 (N_14876,N_13972,N_13315);
xnor U14877 (N_14877,N_13347,N_13355);
nand U14878 (N_14878,N_13554,N_13198);
nand U14879 (N_14879,N_13387,N_13291);
and U14880 (N_14880,N_13187,N_13403);
nand U14881 (N_14881,N_13572,N_13812);
and U14882 (N_14882,N_13034,N_13801);
nand U14883 (N_14883,N_13660,N_13516);
xnor U14884 (N_14884,N_13106,N_13602);
xnor U14885 (N_14885,N_13346,N_13764);
xnor U14886 (N_14886,N_13159,N_13047);
or U14887 (N_14887,N_13425,N_13116);
or U14888 (N_14888,N_13078,N_13971);
nand U14889 (N_14889,N_13965,N_13646);
or U14890 (N_14890,N_13446,N_13601);
and U14891 (N_14891,N_13385,N_13899);
nor U14892 (N_14892,N_13218,N_13222);
nor U14893 (N_14893,N_13794,N_13415);
or U14894 (N_14894,N_13762,N_13289);
xnor U14895 (N_14895,N_13839,N_13610);
xnor U14896 (N_14896,N_13376,N_13574);
and U14897 (N_14897,N_13020,N_13448);
nand U14898 (N_14898,N_13645,N_13529);
nor U14899 (N_14899,N_13888,N_13072);
or U14900 (N_14900,N_13742,N_13752);
or U14901 (N_14901,N_13111,N_13573);
and U14902 (N_14902,N_13496,N_13035);
nand U14903 (N_14903,N_13855,N_13973);
and U14904 (N_14904,N_13201,N_13182);
nand U14905 (N_14905,N_13974,N_13094);
nor U14906 (N_14906,N_13028,N_13220);
and U14907 (N_14907,N_13032,N_13375);
and U14908 (N_14908,N_13920,N_13360);
and U14909 (N_14909,N_13405,N_13241);
nand U14910 (N_14910,N_13437,N_13504);
xor U14911 (N_14911,N_13562,N_13984);
xnor U14912 (N_14912,N_13052,N_13602);
and U14913 (N_14913,N_13906,N_13542);
nor U14914 (N_14914,N_13830,N_13993);
and U14915 (N_14915,N_13040,N_13307);
nand U14916 (N_14916,N_13707,N_13374);
nor U14917 (N_14917,N_13888,N_13736);
nand U14918 (N_14918,N_13920,N_13343);
and U14919 (N_14919,N_13851,N_13773);
xnor U14920 (N_14920,N_13122,N_13951);
nand U14921 (N_14921,N_13211,N_13270);
or U14922 (N_14922,N_13742,N_13043);
nand U14923 (N_14923,N_13529,N_13483);
and U14924 (N_14924,N_13144,N_13092);
and U14925 (N_14925,N_13294,N_13076);
nand U14926 (N_14926,N_13695,N_13632);
nor U14927 (N_14927,N_13558,N_13166);
nand U14928 (N_14928,N_13840,N_13665);
nor U14929 (N_14929,N_13029,N_13401);
or U14930 (N_14930,N_13077,N_13294);
xor U14931 (N_14931,N_13695,N_13077);
xnor U14932 (N_14932,N_13284,N_13457);
and U14933 (N_14933,N_13039,N_13097);
nand U14934 (N_14934,N_13464,N_13535);
xnor U14935 (N_14935,N_13124,N_13290);
or U14936 (N_14936,N_13479,N_13867);
or U14937 (N_14937,N_13943,N_13701);
xor U14938 (N_14938,N_13193,N_13870);
nand U14939 (N_14939,N_13759,N_13816);
and U14940 (N_14940,N_13579,N_13368);
and U14941 (N_14941,N_13364,N_13778);
xor U14942 (N_14942,N_13368,N_13540);
nand U14943 (N_14943,N_13365,N_13756);
xor U14944 (N_14944,N_13645,N_13078);
or U14945 (N_14945,N_13805,N_13328);
nand U14946 (N_14946,N_13722,N_13880);
or U14947 (N_14947,N_13129,N_13844);
and U14948 (N_14948,N_13965,N_13738);
or U14949 (N_14949,N_13813,N_13632);
or U14950 (N_14950,N_13724,N_13416);
nor U14951 (N_14951,N_13647,N_13066);
xnor U14952 (N_14952,N_13461,N_13831);
xnor U14953 (N_14953,N_13497,N_13020);
or U14954 (N_14954,N_13353,N_13995);
and U14955 (N_14955,N_13342,N_13951);
nand U14956 (N_14956,N_13072,N_13193);
or U14957 (N_14957,N_13308,N_13904);
or U14958 (N_14958,N_13643,N_13637);
or U14959 (N_14959,N_13114,N_13610);
xnor U14960 (N_14960,N_13804,N_13726);
nor U14961 (N_14961,N_13661,N_13242);
and U14962 (N_14962,N_13728,N_13563);
nand U14963 (N_14963,N_13865,N_13357);
and U14964 (N_14964,N_13022,N_13471);
nor U14965 (N_14965,N_13211,N_13851);
and U14966 (N_14966,N_13722,N_13763);
xor U14967 (N_14967,N_13484,N_13743);
xnor U14968 (N_14968,N_13398,N_13504);
nor U14969 (N_14969,N_13579,N_13102);
xor U14970 (N_14970,N_13008,N_13277);
or U14971 (N_14971,N_13719,N_13743);
nor U14972 (N_14972,N_13344,N_13172);
or U14973 (N_14973,N_13476,N_13166);
nor U14974 (N_14974,N_13999,N_13968);
nor U14975 (N_14975,N_13138,N_13058);
or U14976 (N_14976,N_13170,N_13248);
or U14977 (N_14977,N_13425,N_13185);
and U14978 (N_14978,N_13046,N_13461);
and U14979 (N_14979,N_13618,N_13278);
nand U14980 (N_14980,N_13140,N_13639);
nand U14981 (N_14981,N_13195,N_13194);
nand U14982 (N_14982,N_13930,N_13936);
xor U14983 (N_14983,N_13550,N_13351);
xnor U14984 (N_14984,N_13183,N_13149);
nand U14985 (N_14985,N_13820,N_13528);
and U14986 (N_14986,N_13829,N_13579);
or U14987 (N_14987,N_13056,N_13085);
nor U14988 (N_14988,N_13410,N_13301);
or U14989 (N_14989,N_13392,N_13553);
nor U14990 (N_14990,N_13007,N_13459);
and U14991 (N_14991,N_13877,N_13792);
or U14992 (N_14992,N_13322,N_13935);
xnor U14993 (N_14993,N_13449,N_13427);
and U14994 (N_14994,N_13915,N_13834);
xor U14995 (N_14995,N_13425,N_13929);
and U14996 (N_14996,N_13842,N_13435);
or U14997 (N_14997,N_13359,N_13447);
nand U14998 (N_14998,N_13808,N_13496);
nor U14999 (N_14999,N_13177,N_13472);
or U15000 (N_15000,N_14461,N_14323);
and U15001 (N_15001,N_14072,N_14659);
nand U15002 (N_15002,N_14830,N_14357);
xor U15003 (N_15003,N_14044,N_14681);
or U15004 (N_15004,N_14180,N_14256);
nor U15005 (N_15005,N_14413,N_14941);
nand U15006 (N_15006,N_14593,N_14492);
nand U15007 (N_15007,N_14149,N_14460);
xor U15008 (N_15008,N_14902,N_14817);
nand U15009 (N_15009,N_14863,N_14721);
nand U15010 (N_15010,N_14932,N_14799);
or U15011 (N_15011,N_14995,N_14914);
or U15012 (N_15012,N_14478,N_14561);
nor U15013 (N_15013,N_14582,N_14675);
and U15014 (N_15014,N_14191,N_14209);
xnor U15015 (N_15015,N_14848,N_14885);
and U15016 (N_15016,N_14345,N_14882);
and U15017 (N_15017,N_14510,N_14815);
nor U15018 (N_15018,N_14971,N_14860);
nor U15019 (N_15019,N_14155,N_14532);
and U15020 (N_15020,N_14019,N_14497);
or U15021 (N_15021,N_14583,N_14741);
nand U15022 (N_15022,N_14810,N_14168);
nor U15023 (N_15023,N_14321,N_14097);
and U15024 (N_15024,N_14515,N_14785);
or U15025 (N_15025,N_14813,N_14892);
xor U15026 (N_15026,N_14259,N_14333);
xor U15027 (N_15027,N_14748,N_14753);
or U15028 (N_15028,N_14327,N_14551);
or U15029 (N_15029,N_14276,N_14852);
and U15030 (N_15030,N_14416,N_14189);
nor U15031 (N_15031,N_14513,N_14747);
or U15032 (N_15032,N_14875,N_14338);
xnor U15033 (N_15033,N_14722,N_14030);
or U15034 (N_15034,N_14847,N_14490);
nand U15035 (N_15035,N_14027,N_14322);
nor U15036 (N_15036,N_14074,N_14867);
or U15037 (N_15037,N_14636,N_14969);
nand U15038 (N_15038,N_14405,N_14639);
nor U15039 (N_15039,N_14621,N_14265);
xor U15040 (N_15040,N_14238,N_14226);
or U15041 (N_15041,N_14433,N_14602);
nor U15042 (N_15042,N_14887,N_14175);
xor U15043 (N_15043,N_14518,N_14505);
nand U15044 (N_15044,N_14397,N_14279);
or U15045 (N_15045,N_14751,N_14884);
nand U15046 (N_15046,N_14542,N_14300);
and U15047 (N_15047,N_14701,N_14579);
nor U15048 (N_15048,N_14800,N_14543);
and U15049 (N_15049,N_14126,N_14438);
xnor U15050 (N_15050,N_14428,N_14060);
or U15051 (N_15051,N_14704,N_14371);
and U15052 (N_15052,N_14408,N_14444);
nor U15053 (N_15053,N_14893,N_14352);
nand U15054 (N_15054,N_14267,N_14114);
and U15055 (N_15055,N_14698,N_14919);
xor U15056 (N_15056,N_14319,N_14609);
nand U15057 (N_15057,N_14504,N_14784);
and U15058 (N_15058,N_14950,N_14295);
nor U15059 (N_15059,N_14101,N_14253);
nor U15060 (N_15060,N_14682,N_14442);
nand U15061 (N_15061,N_14630,N_14156);
nor U15062 (N_15062,N_14744,N_14911);
nor U15063 (N_15063,N_14084,N_14772);
and U15064 (N_15064,N_14576,N_14217);
nand U15065 (N_15065,N_14767,N_14344);
xnor U15066 (N_15066,N_14528,N_14177);
and U15067 (N_15067,N_14961,N_14261);
or U15068 (N_15068,N_14945,N_14263);
nand U15069 (N_15069,N_14029,N_14110);
xor U15070 (N_15070,N_14764,N_14953);
nand U15071 (N_15071,N_14720,N_14173);
nor U15072 (N_15072,N_14890,N_14834);
xor U15073 (N_15073,N_14994,N_14182);
or U15074 (N_15074,N_14017,N_14003);
xnor U15075 (N_15075,N_14805,N_14018);
or U15076 (N_15076,N_14394,N_14700);
xnor U15077 (N_15077,N_14844,N_14568);
and U15078 (N_15078,N_14475,N_14250);
nand U15079 (N_15079,N_14788,N_14752);
or U15080 (N_15080,N_14880,N_14098);
xor U15081 (N_15081,N_14087,N_14973);
xnor U15082 (N_15082,N_14610,N_14100);
nor U15083 (N_15083,N_14757,N_14904);
xor U15084 (N_15084,N_14021,N_14996);
or U15085 (N_15085,N_14917,N_14999);
nor U15086 (N_15086,N_14674,N_14496);
nor U15087 (N_15087,N_14640,N_14251);
and U15088 (N_15088,N_14872,N_14968);
or U15089 (N_15089,N_14960,N_14529);
or U15090 (N_15090,N_14467,N_14943);
nor U15091 (N_15091,N_14270,N_14680);
xnor U15092 (N_15092,N_14679,N_14913);
nor U15093 (N_15093,N_14071,N_14476);
nor U15094 (N_15094,N_14427,N_14735);
nor U15095 (N_15095,N_14443,N_14678);
and U15096 (N_15096,N_14170,N_14174);
nand U15097 (N_15097,N_14311,N_14406);
nor U15098 (N_15098,N_14131,N_14690);
and U15099 (N_15099,N_14749,N_14124);
xor U15100 (N_15100,N_14506,N_14448);
and U15101 (N_15101,N_14082,N_14203);
or U15102 (N_15102,N_14703,N_14570);
nand U15103 (N_15103,N_14934,N_14358);
or U15104 (N_15104,N_14755,N_14694);
xnor U15105 (N_15105,N_14670,N_14618);
nand U15106 (N_15106,N_14667,N_14555);
or U15107 (N_15107,N_14992,N_14857);
nor U15108 (N_15108,N_14676,N_14435);
xor U15109 (N_15109,N_14851,N_14056);
nand U15110 (N_15110,N_14033,N_14920);
or U15111 (N_15111,N_14395,N_14828);
xor U15112 (N_15112,N_14137,N_14318);
and U15113 (N_15113,N_14502,N_14252);
nand U15114 (N_15114,N_14717,N_14424);
xnor U15115 (N_15115,N_14669,N_14736);
or U15116 (N_15116,N_14468,N_14310);
nand U15117 (N_15117,N_14449,N_14092);
nand U15118 (N_15118,N_14835,N_14485);
nand U15119 (N_15119,N_14465,N_14944);
and U15120 (N_15120,N_14500,N_14373);
or U15121 (N_15121,N_14967,N_14545);
or U15122 (N_15122,N_14858,N_14556);
and U15123 (N_15123,N_14931,N_14199);
and U15124 (N_15124,N_14819,N_14483);
and U15125 (N_15125,N_14574,N_14301);
nand U15126 (N_15126,N_14009,N_14959);
nand U15127 (N_15127,N_14070,N_14275);
xor U15128 (N_15128,N_14763,N_14878);
xor U15129 (N_15129,N_14981,N_14566);
nand U15130 (N_15130,N_14894,N_14011);
or U15131 (N_15131,N_14268,N_14601);
or U15132 (N_15132,N_14974,N_14787);
nor U15133 (N_15133,N_14487,N_14160);
nor U15134 (N_15134,N_14620,N_14419);
xor U15135 (N_15135,N_14525,N_14530);
xor U15136 (N_15136,N_14000,N_14255);
nand U15137 (N_15137,N_14043,N_14673);
nor U15138 (N_15138,N_14606,N_14329);
and U15139 (N_15139,N_14888,N_14103);
or U15140 (N_15140,N_14269,N_14775);
xor U15141 (N_15141,N_14184,N_14808);
nand U15142 (N_15142,N_14796,N_14198);
nand U15143 (N_15143,N_14112,N_14164);
xor U15144 (N_15144,N_14061,N_14527);
nand U15145 (N_15145,N_14861,N_14624);
or U15146 (N_15146,N_14647,N_14572);
xor U15147 (N_15147,N_14598,N_14133);
xor U15148 (N_15148,N_14942,N_14113);
nand U15149 (N_15149,N_14993,N_14140);
and U15150 (N_15150,N_14446,N_14066);
nand U15151 (N_15151,N_14782,N_14454);
or U15152 (N_15152,N_14531,N_14372);
and U15153 (N_15153,N_14053,N_14615);
nor U15154 (N_15154,N_14010,N_14425);
and U15155 (N_15155,N_14686,N_14392);
xnor U15156 (N_15156,N_14672,N_14874);
xor U15157 (N_15157,N_14708,N_14190);
nand U15158 (N_15158,N_14022,N_14738);
nand U15159 (N_15159,N_14626,N_14991);
xnor U15160 (N_15160,N_14035,N_14305);
xnor U15161 (N_15161,N_14325,N_14462);
nand U15162 (N_15162,N_14638,N_14871);
nor U15163 (N_15163,N_14432,N_14348);
and U15164 (N_15164,N_14907,N_14554);
nor U15165 (N_15165,N_14864,N_14109);
nor U15166 (N_15166,N_14731,N_14258);
xnor U15167 (N_15167,N_14289,N_14334);
nor U15168 (N_15168,N_14613,N_14507);
nor U15169 (N_15169,N_14115,N_14916);
or U15170 (N_15170,N_14662,N_14347);
or U15171 (N_15171,N_14565,N_14577);
or U15172 (N_15172,N_14227,N_14692);
xnor U15173 (N_15173,N_14280,N_14687);
or U15174 (N_15174,N_14353,N_14644);
nor U15175 (N_15175,N_14288,N_14363);
and U15176 (N_15176,N_14415,N_14926);
nand U15177 (N_15177,N_14240,N_14211);
nand U15178 (N_15178,N_14656,N_14377);
nor U15179 (N_15179,N_14266,N_14158);
or U15180 (N_15180,N_14599,N_14223);
nor U15181 (N_15181,N_14277,N_14336);
nand U15182 (N_15182,N_14645,N_14842);
nand U15183 (N_15183,N_14723,N_14459);
xnor U15184 (N_15184,N_14151,N_14648);
and U15185 (N_15185,N_14273,N_14023);
nand U15186 (N_15186,N_14936,N_14845);
xor U15187 (N_15187,N_14059,N_14829);
xor U15188 (N_15188,N_14564,N_14470);
xor U15189 (N_15189,N_14396,N_14099);
nor U15190 (N_15190,N_14612,N_14575);
nand U15191 (N_15191,N_14776,N_14388);
nor U15192 (N_15192,N_14581,N_14411);
and U15193 (N_15193,N_14924,N_14458);
and U15194 (N_15194,N_14024,N_14308);
or U15195 (N_15195,N_14984,N_14883);
and U15196 (N_15196,N_14290,N_14052);
xnor U15197 (N_15197,N_14452,N_14351);
and U15198 (N_15198,N_14997,N_14355);
nand U15199 (N_15199,N_14798,N_14412);
xnor U15200 (N_15200,N_14380,N_14517);
xor U15201 (N_15201,N_14341,N_14797);
or U15202 (N_15202,N_14282,N_14856);
nand U15203 (N_15203,N_14865,N_14144);
nor U15204 (N_15204,N_14237,N_14039);
nor U15205 (N_15205,N_14886,N_14132);
and U15206 (N_15206,N_14376,N_14816);
nand U15207 (N_15207,N_14578,N_14786);
xor U15208 (N_15208,N_14324,N_14939);
and U15209 (N_15209,N_14370,N_14331);
nand U15210 (N_15210,N_14135,N_14759);
or U15211 (N_15211,N_14417,N_14434);
xnor U15212 (N_15212,N_14185,N_14756);
and U15213 (N_15213,N_14095,N_14604);
or U15214 (N_15214,N_14063,N_14096);
and U15215 (N_15215,N_14595,N_14054);
nand U15216 (N_15216,N_14702,N_14105);
and U15217 (N_15217,N_14779,N_14143);
and U15218 (N_15218,N_14548,N_14938);
or U15219 (N_15219,N_14794,N_14627);
or U15220 (N_15220,N_14724,N_14387);
xor U15221 (N_15221,N_14389,N_14557);
and U15222 (N_15222,N_14827,N_14479);
xnor U15223 (N_15223,N_14439,N_14012);
or U15224 (N_15224,N_14119,N_14509);
and U15225 (N_15225,N_14422,N_14008);
nand U15226 (N_15226,N_14982,N_14730);
and U15227 (N_15227,N_14512,N_14309);
nand U15228 (N_15228,N_14495,N_14711);
nand U15229 (N_15229,N_14150,N_14803);
nand U15230 (N_15230,N_14716,N_14014);
or U15231 (N_15231,N_14026,N_14078);
nor U15232 (N_15232,N_14418,N_14846);
nand U15233 (N_15233,N_14218,N_14117);
or U15234 (N_15234,N_14623,N_14503);
or U15235 (N_15235,N_14818,N_14278);
xor U15236 (N_15236,N_14773,N_14243);
and U15237 (N_15237,N_14127,N_14873);
nand U15238 (N_15238,N_14954,N_14034);
or U15239 (N_15239,N_14677,N_14225);
nand U15240 (N_15240,N_14360,N_14048);
nor U15241 (N_15241,N_14544,N_14130);
xor U15242 (N_15242,N_14178,N_14589);
xor U15243 (N_15243,N_14165,N_14332);
or U15244 (N_15244,N_14866,N_14657);
nand U15245 (N_15245,N_14665,N_14603);
or U15246 (N_15246,N_14129,N_14346);
xor U15247 (N_15247,N_14952,N_14949);
or U15248 (N_15248,N_14963,N_14364);
nand U15249 (N_15249,N_14366,N_14743);
xor U15250 (N_15250,N_14036,N_14391);
nor U15251 (N_15251,N_14712,N_14868);
nand U15252 (N_15252,N_14286,N_14608);
nor U15253 (N_15253,N_14652,N_14409);
nor U15254 (N_15254,N_14660,N_14854);
xor U15255 (N_15255,N_14760,N_14732);
nor U15256 (N_15256,N_14002,N_14075);
nor U15257 (N_15257,N_14713,N_14783);
xor U15258 (N_15258,N_14629,N_14220);
and U15259 (N_15259,N_14634,N_14134);
or U15260 (N_15260,N_14838,N_14795);
or U15261 (N_15261,N_14474,N_14482);
and U15262 (N_15262,N_14912,N_14016);
nand U15263 (N_15263,N_14342,N_14314);
or U15264 (N_15264,N_14725,N_14306);
nand U15265 (N_15265,N_14718,N_14069);
and U15266 (N_15266,N_14777,N_14445);
xor U15267 (N_15267,N_14966,N_14451);
and U15268 (N_15268,N_14186,N_14354);
xor U15269 (N_15269,N_14141,N_14293);
nand U15270 (N_15270,N_14316,N_14244);
nor U15271 (N_15271,N_14402,N_14368);
and U15272 (N_15272,N_14403,N_14539);
nand U15273 (N_15273,N_14849,N_14549);
and U15274 (N_15274,N_14421,N_14179);
xnor U15275 (N_15275,N_14343,N_14375);
xor U15276 (N_15276,N_14921,N_14274);
xor U15277 (N_15277,N_14121,N_14242);
or U15278 (N_15278,N_14356,N_14754);
nand U15279 (N_15279,N_14330,N_14699);
nor U15280 (N_15280,N_14869,N_14384);
nor U15281 (N_15281,N_14664,N_14614);
and U15282 (N_15282,N_14107,N_14567);
or U15283 (N_15283,N_14840,N_14005);
nor U15284 (N_15284,N_14862,N_14637);
xor U15285 (N_15285,N_14560,N_14654);
xnor U15286 (N_15286,N_14216,N_14559);
or U15287 (N_15287,N_14970,N_14200);
xor U15288 (N_15288,N_14622,N_14688);
nor U15289 (N_15289,N_14284,N_14207);
nor U15290 (N_15290,N_14933,N_14666);
and U15291 (N_15291,N_14315,N_14522);
nor U15292 (N_15292,N_14705,N_14239);
nor U15293 (N_15293,N_14457,N_14587);
xor U15294 (N_15294,N_14958,N_14778);
xnor U15295 (N_15295,N_14247,N_14312);
xor U15296 (N_15296,N_14616,N_14015);
nand U15297 (N_15297,N_14617,N_14025);
or U15298 (N_15298,N_14249,N_14596);
or U15299 (N_15299,N_14167,N_14983);
and U15300 (N_15300,N_14832,N_14208);
nor U15301 (N_15301,N_14927,N_14379);
and U15302 (N_15302,N_14440,N_14147);
nand U15303 (N_15303,N_14770,N_14139);
and U15304 (N_15304,N_14154,N_14349);
nor U15305 (N_15305,N_14369,N_14739);
xnor U15306 (N_15306,N_14740,N_14714);
nand U15307 (N_15307,N_14374,N_14766);
and U15308 (N_15308,N_14812,N_14298);
and U15309 (N_15309,N_14940,N_14441);
xor U15310 (N_15310,N_14195,N_14987);
and U15311 (N_15311,N_14192,N_14196);
xor U15312 (N_15312,N_14317,N_14965);
nand U15313 (N_15313,N_14588,N_14520);
xnor U15314 (N_15314,N_14853,N_14597);
xnor U15315 (N_15315,N_14401,N_14859);
xnor U15316 (N_15316,N_14047,N_14076);
xnor U15317 (N_15317,N_14163,N_14161);
xor U15318 (N_15318,N_14068,N_14801);
or U15319 (N_15319,N_14594,N_14042);
xor U15320 (N_15320,N_14745,N_14715);
and U15321 (N_15321,N_14536,N_14480);
nor U15322 (N_15322,N_14643,N_14836);
xnor U15323 (N_15323,N_14929,N_14706);
nor U15324 (N_15324,N_14655,N_14550);
xnor U15325 (N_15325,N_14447,N_14264);
nand U15326 (N_15326,N_14563,N_14436);
nand U15327 (N_15327,N_14635,N_14399);
and U15328 (N_15328,N_14359,N_14260);
or U15329 (N_15329,N_14906,N_14386);
xor U15330 (N_15330,N_14526,N_14918);
or U15331 (N_15331,N_14962,N_14214);
nand U15332 (N_15332,N_14651,N_14108);
or U15333 (N_15333,N_14839,N_14946);
and U15334 (N_15334,N_14841,N_14407);
nand U15335 (N_15335,N_14224,N_14058);
nand U15336 (N_15336,N_14650,N_14899);
or U15337 (N_15337,N_14085,N_14233);
and U15338 (N_15338,N_14511,N_14262);
nand U15339 (N_15339,N_14197,N_14206);
xor U15340 (N_15340,N_14737,N_14695);
and U15341 (N_15341,N_14925,N_14619);
and U15342 (N_15342,N_14294,N_14326);
nand U15343 (N_15343,N_14245,N_14055);
nor U15344 (N_15344,N_14296,N_14398);
nor U15345 (N_15345,N_14145,N_14361);
nor U15346 (N_15346,N_14928,N_14083);
or U15347 (N_15347,N_14814,N_14683);
nand U15348 (N_15348,N_14820,N_14453);
xnor U15349 (N_15349,N_14727,N_14248);
nor U15350 (N_15350,N_14535,N_14001);
and U15351 (N_15351,N_14937,N_14758);
xor U15352 (N_15352,N_14205,N_14877);
xnor U15353 (N_15353,N_14091,N_14481);
and U15354 (N_15354,N_14930,N_14335);
xnor U15355 (N_15355,N_14106,N_14313);
xor U15356 (N_15356,N_14663,N_14172);
or U15357 (N_15357,N_14896,N_14230);
xor U15358 (N_15358,N_14519,N_14881);
and U15359 (N_15359,N_14146,N_14585);
xor U15360 (N_15360,N_14494,N_14302);
or U15361 (N_15361,N_14508,N_14607);
nor U15362 (N_15362,N_14235,N_14553);
or U15363 (N_15363,N_14383,N_14685);
and U15364 (N_15364,N_14390,N_14210);
xor U15365 (N_15365,N_14304,N_14988);
and U15366 (N_15366,N_14989,N_14824);
nand U15367 (N_15367,N_14032,N_14537);
nand U15368 (N_15368,N_14790,N_14693);
xor U15369 (N_15369,N_14891,N_14328);
and U15370 (N_15370,N_14089,N_14957);
or U15371 (N_15371,N_14037,N_14123);
nor U15372 (N_15372,N_14120,N_14649);
and U15373 (N_15373,N_14285,N_14013);
nor U15374 (N_15374,N_14420,N_14792);
nand U15375 (N_15375,N_14562,N_14696);
nand U15376 (N_15376,N_14291,N_14094);
xnor U15377 (N_15377,N_14362,N_14488);
xor U15378 (N_15378,N_14236,N_14762);
and U15379 (N_15379,N_14153,N_14534);
and U15380 (N_15380,N_14771,N_14558);
or U15381 (N_15381,N_14498,N_14365);
xor U15382 (N_15382,N_14437,N_14837);
or U15383 (N_15383,N_14985,N_14283);
nand U15384 (N_15384,N_14631,N_14978);
xnor U15385 (N_15385,N_14793,N_14804);
nand U15386 (N_15386,N_14051,N_14118);
and U15387 (N_15387,N_14975,N_14908);
nand U15388 (N_15388,N_14472,N_14590);
xnor U15389 (N_15389,N_14499,N_14229);
or U15390 (N_15390,N_14125,N_14935);
nor U15391 (N_15391,N_14547,N_14004);
nor U15392 (N_15392,N_14947,N_14876);
and U15393 (N_15393,N_14761,N_14430);
and U15394 (N_15394,N_14031,N_14050);
xor U15395 (N_15395,N_14948,N_14768);
or U15396 (N_15396,N_14922,N_14122);
nand U15397 (N_15397,N_14990,N_14455);
nand U15398 (N_15398,N_14769,N_14552);
nand U15399 (N_15399,N_14489,N_14806);
or U15400 (N_15400,N_14972,N_14956);
xor U15401 (N_15401,N_14750,N_14188);
xnor U15402 (N_15402,N_14429,N_14102);
xor U15403 (N_15403,N_14471,N_14213);
nand U15404 (N_15404,N_14831,N_14524);
and U15405 (N_15405,N_14215,N_14337);
and U15406 (N_15406,N_14514,N_14710);
and U15407 (N_15407,N_14774,N_14791);
or U15408 (N_15408,N_14400,N_14909);
xnor U15409 (N_15409,N_14231,N_14040);
nor U15410 (N_15410,N_14584,N_14658);
and U15411 (N_15411,N_14905,N_14986);
nand U15412 (N_15412,N_14642,N_14697);
or U15413 (N_15413,N_14915,N_14038);
xor U15414 (N_15414,N_14426,N_14671);
and U15415 (N_15415,N_14668,N_14569);
or U15416 (N_15416,N_14684,N_14028);
and U15417 (N_15417,N_14297,N_14951);
and U15418 (N_15418,N_14628,N_14726);
xnor U15419 (N_15419,N_14212,N_14350);
nand U15420 (N_15420,N_14491,N_14385);
nor U15421 (N_15421,N_14709,N_14065);
or U15422 (N_15422,N_14661,N_14166);
nor U15423 (N_15423,N_14340,N_14728);
and U15424 (N_15424,N_14171,N_14073);
nor U15425 (N_15425,N_14592,N_14580);
and U15426 (N_15426,N_14707,N_14691);
nor U15427 (N_15427,N_14181,N_14006);
xor U15428 (N_15428,N_14469,N_14466);
nor U15429 (N_15429,N_14546,N_14641);
nand U15430 (N_15430,N_14605,N_14201);
or U15431 (N_15431,N_14104,N_14923);
xor U15432 (N_15432,N_14802,N_14222);
and U15433 (N_15433,N_14281,N_14646);
or U15434 (N_15434,N_14378,N_14228);
or U15435 (N_15435,N_14964,N_14538);
xor U15436 (N_15436,N_14271,N_14142);
nor U15437 (N_15437,N_14367,N_14746);
nand U15438 (N_15438,N_14600,N_14254);
nor U15439 (N_15439,N_14116,N_14232);
and U15440 (N_15440,N_14910,N_14781);
or U15441 (N_15441,N_14955,N_14573);
xor U15442 (N_15442,N_14414,N_14879);
and U15443 (N_15443,N_14523,N_14611);
xnor U15444 (N_15444,N_14850,N_14111);
nand U15445 (N_15445,N_14020,N_14041);
and U15446 (N_15446,N_14571,N_14895);
and U15447 (N_15447,N_14077,N_14625);
xnor U15448 (N_15448,N_14093,N_14272);
and U15449 (N_15449,N_14241,N_14176);
nand U15450 (N_15450,N_14183,N_14067);
nand U15451 (N_15451,N_14079,N_14257);
and U15452 (N_15452,N_14410,N_14979);
or U15453 (N_15453,N_14521,N_14632);
nor U15454 (N_15454,N_14136,N_14221);
xnor U15455 (N_15455,N_14734,N_14540);
xnor U15456 (N_15456,N_14823,N_14733);
nand U15457 (N_15457,N_14825,N_14187);
or U15458 (N_15458,N_14809,N_14138);
or U15459 (N_15459,N_14423,N_14090);
nand U15460 (N_15460,N_14516,N_14486);
nor U15461 (N_15461,N_14477,N_14404);
nand U15462 (N_15462,N_14080,N_14431);
xnor U15463 (N_15463,N_14339,N_14689);
nand U15464 (N_15464,N_14780,N_14193);
or U15465 (N_15465,N_14586,N_14897);
and U15466 (N_15466,N_14541,N_14900);
and U15467 (N_15467,N_14046,N_14889);
and U15468 (N_15468,N_14307,N_14765);
nor U15469 (N_15469,N_14493,N_14219);
nand U15470 (N_15470,N_14484,N_14501);
nand U15471 (N_15471,N_14870,N_14903);
or U15472 (N_15472,N_14807,N_14162);
xnor U15473 (N_15473,N_14148,N_14287);
nor U15474 (N_15474,N_14826,N_14152);
nor U15475 (N_15475,N_14976,N_14202);
xor U15476 (N_15476,N_14789,N_14450);
xnor U15477 (N_15477,N_14064,N_14591);
xor U15478 (N_15478,N_14292,N_14719);
nor U15479 (N_15479,N_14007,N_14898);
nor U15480 (N_15480,N_14320,N_14246);
nor U15481 (N_15481,N_14980,N_14088);
nor U15482 (N_15482,N_14128,N_14533);
nand U15483 (N_15483,N_14049,N_14057);
or U15484 (N_15484,N_14381,N_14463);
or U15485 (N_15485,N_14633,N_14081);
nor U15486 (N_15486,N_14303,N_14843);
nor U15487 (N_15487,N_14234,N_14821);
xor U15488 (N_15488,N_14729,N_14855);
nor U15489 (N_15489,N_14382,N_14045);
nor U15490 (N_15490,N_14833,N_14086);
nand U15491 (N_15491,N_14977,N_14998);
nand U15492 (N_15492,N_14204,N_14194);
and U15493 (N_15493,N_14473,N_14456);
nor U15494 (N_15494,N_14811,N_14742);
xor U15495 (N_15495,N_14822,N_14393);
and U15496 (N_15496,N_14169,N_14901);
and U15497 (N_15497,N_14062,N_14653);
or U15498 (N_15498,N_14159,N_14464);
xnor U15499 (N_15499,N_14157,N_14299);
nand U15500 (N_15500,N_14490,N_14577);
and U15501 (N_15501,N_14052,N_14001);
nand U15502 (N_15502,N_14804,N_14478);
xor U15503 (N_15503,N_14318,N_14954);
or U15504 (N_15504,N_14354,N_14794);
or U15505 (N_15505,N_14968,N_14442);
xnor U15506 (N_15506,N_14071,N_14703);
nor U15507 (N_15507,N_14584,N_14947);
nand U15508 (N_15508,N_14631,N_14042);
and U15509 (N_15509,N_14763,N_14384);
nand U15510 (N_15510,N_14111,N_14935);
nand U15511 (N_15511,N_14823,N_14427);
or U15512 (N_15512,N_14217,N_14692);
and U15513 (N_15513,N_14843,N_14126);
xor U15514 (N_15514,N_14077,N_14017);
nor U15515 (N_15515,N_14208,N_14412);
and U15516 (N_15516,N_14370,N_14477);
and U15517 (N_15517,N_14974,N_14039);
or U15518 (N_15518,N_14416,N_14330);
or U15519 (N_15519,N_14326,N_14027);
or U15520 (N_15520,N_14722,N_14513);
nor U15521 (N_15521,N_14559,N_14697);
nand U15522 (N_15522,N_14786,N_14926);
or U15523 (N_15523,N_14178,N_14767);
nor U15524 (N_15524,N_14387,N_14149);
and U15525 (N_15525,N_14106,N_14545);
and U15526 (N_15526,N_14980,N_14580);
nor U15527 (N_15527,N_14089,N_14023);
nor U15528 (N_15528,N_14027,N_14437);
nor U15529 (N_15529,N_14616,N_14032);
xor U15530 (N_15530,N_14339,N_14290);
and U15531 (N_15531,N_14431,N_14141);
and U15532 (N_15532,N_14076,N_14036);
nand U15533 (N_15533,N_14319,N_14619);
xor U15534 (N_15534,N_14676,N_14247);
xnor U15535 (N_15535,N_14405,N_14592);
nand U15536 (N_15536,N_14799,N_14212);
nand U15537 (N_15537,N_14465,N_14136);
and U15538 (N_15538,N_14887,N_14233);
or U15539 (N_15539,N_14030,N_14755);
or U15540 (N_15540,N_14804,N_14055);
or U15541 (N_15541,N_14060,N_14306);
or U15542 (N_15542,N_14726,N_14346);
xor U15543 (N_15543,N_14126,N_14925);
or U15544 (N_15544,N_14206,N_14334);
and U15545 (N_15545,N_14062,N_14076);
or U15546 (N_15546,N_14083,N_14336);
xor U15547 (N_15547,N_14204,N_14629);
nand U15548 (N_15548,N_14003,N_14556);
nand U15549 (N_15549,N_14423,N_14771);
and U15550 (N_15550,N_14741,N_14641);
xor U15551 (N_15551,N_14162,N_14524);
nor U15552 (N_15552,N_14087,N_14083);
and U15553 (N_15553,N_14593,N_14080);
or U15554 (N_15554,N_14258,N_14282);
nor U15555 (N_15555,N_14571,N_14465);
nand U15556 (N_15556,N_14004,N_14419);
nand U15557 (N_15557,N_14434,N_14164);
nor U15558 (N_15558,N_14145,N_14881);
nand U15559 (N_15559,N_14682,N_14515);
xnor U15560 (N_15560,N_14669,N_14441);
and U15561 (N_15561,N_14898,N_14753);
nor U15562 (N_15562,N_14009,N_14544);
and U15563 (N_15563,N_14764,N_14105);
and U15564 (N_15564,N_14444,N_14748);
or U15565 (N_15565,N_14124,N_14527);
nand U15566 (N_15566,N_14006,N_14489);
nor U15567 (N_15567,N_14117,N_14957);
or U15568 (N_15568,N_14175,N_14897);
xnor U15569 (N_15569,N_14638,N_14841);
nor U15570 (N_15570,N_14798,N_14004);
xnor U15571 (N_15571,N_14646,N_14288);
nand U15572 (N_15572,N_14521,N_14779);
xor U15573 (N_15573,N_14904,N_14515);
and U15574 (N_15574,N_14475,N_14783);
nor U15575 (N_15575,N_14911,N_14758);
and U15576 (N_15576,N_14996,N_14976);
xnor U15577 (N_15577,N_14712,N_14391);
or U15578 (N_15578,N_14948,N_14211);
or U15579 (N_15579,N_14325,N_14297);
or U15580 (N_15580,N_14340,N_14739);
nor U15581 (N_15581,N_14040,N_14671);
nor U15582 (N_15582,N_14607,N_14891);
xor U15583 (N_15583,N_14338,N_14442);
xnor U15584 (N_15584,N_14539,N_14680);
nand U15585 (N_15585,N_14803,N_14585);
xnor U15586 (N_15586,N_14918,N_14625);
nand U15587 (N_15587,N_14512,N_14823);
nor U15588 (N_15588,N_14695,N_14175);
and U15589 (N_15589,N_14509,N_14750);
nor U15590 (N_15590,N_14625,N_14062);
and U15591 (N_15591,N_14877,N_14298);
or U15592 (N_15592,N_14383,N_14359);
xor U15593 (N_15593,N_14473,N_14248);
and U15594 (N_15594,N_14511,N_14773);
nor U15595 (N_15595,N_14447,N_14486);
xor U15596 (N_15596,N_14186,N_14365);
and U15597 (N_15597,N_14057,N_14829);
xor U15598 (N_15598,N_14047,N_14797);
nor U15599 (N_15599,N_14973,N_14729);
nand U15600 (N_15600,N_14188,N_14812);
xnor U15601 (N_15601,N_14167,N_14889);
xnor U15602 (N_15602,N_14083,N_14330);
xor U15603 (N_15603,N_14162,N_14113);
nand U15604 (N_15604,N_14603,N_14474);
and U15605 (N_15605,N_14776,N_14046);
nand U15606 (N_15606,N_14042,N_14218);
nor U15607 (N_15607,N_14854,N_14116);
nand U15608 (N_15608,N_14311,N_14863);
nand U15609 (N_15609,N_14615,N_14542);
nor U15610 (N_15610,N_14464,N_14822);
xnor U15611 (N_15611,N_14605,N_14047);
and U15612 (N_15612,N_14528,N_14737);
and U15613 (N_15613,N_14169,N_14919);
nand U15614 (N_15614,N_14342,N_14794);
nor U15615 (N_15615,N_14415,N_14255);
and U15616 (N_15616,N_14843,N_14362);
nor U15617 (N_15617,N_14340,N_14135);
or U15618 (N_15618,N_14755,N_14645);
nor U15619 (N_15619,N_14741,N_14508);
xnor U15620 (N_15620,N_14885,N_14632);
nand U15621 (N_15621,N_14952,N_14006);
nor U15622 (N_15622,N_14718,N_14526);
or U15623 (N_15623,N_14727,N_14368);
or U15624 (N_15624,N_14211,N_14994);
nand U15625 (N_15625,N_14814,N_14628);
or U15626 (N_15626,N_14444,N_14485);
or U15627 (N_15627,N_14340,N_14247);
and U15628 (N_15628,N_14458,N_14813);
or U15629 (N_15629,N_14037,N_14418);
nand U15630 (N_15630,N_14207,N_14480);
nor U15631 (N_15631,N_14795,N_14875);
nor U15632 (N_15632,N_14652,N_14266);
or U15633 (N_15633,N_14178,N_14350);
xor U15634 (N_15634,N_14253,N_14817);
nand U15635 (N_15635,N_14882,N_14425);
and U15636 (N_15636,N_14572,N_14226);
nand U15637 (N_15637,N_14938,N_14667);
nor U15638 (N_15638,N_14946,N_14628);
or U15639 (N_15639,N_14528,N_14458);
nand U15640 (N_15640,N_14045,N_14104);
nand U15641 (N_15641,N_14773,N_14590);
or U15642 (N_15642,N_14473,N_14756);
and U15643 (N_15643,N_14647,N_14478);
or U15644 (N_15644,N_14087,N_14044);
nor U15645 (N_15645,N_14795,N_14798);
nand U15646 (N_15646,N_14655,N_14561);
nor U15647 (N_15647,N_14164,N_14481);
nand U15648 (N_15648,N_14764,N_14867);
nor U15649 (N_15649,N_14029,N_14825);
or U15650 (N_15650,N_14371,N_14364);
or U15651 (N_15651,N_14645,N_14202);
or U15652 (N_15652,N_14336,N_14945);
and U15653 (N_15653,N_14251,N_14233);
or U15654 (N_15654,N_14253,N_14968);
and U15655 (N_15655,N_14527,N_14962);
and U15656 (N_15656,N_14527,N_14111);
xor U15657 (N_15657,N_14431,N_14531);
or U15658 (N_15658,N_14225,N_14632);
nor U15659 (N_15659,N_14173,N_14605);
or U15660 (N_15660,N_14388,N_14818);
xor U15661 (N_15661,N_14300,N_14025);
or U15662 (N_15662,N_14943,N_14988);
nand U15663 (N_15663,N_14132,N_14205);
or U15664 (N_15664,N_14226,N_14587);
and U15665 (N_15665,N_14774,N_14590);
and U15666 (N_15666,N_14674,N_14910);
xnor U15667 (N_15667,N_14157,N_14339);
and U15668 (N_15668,N_14039,N_14597);
nor U15669 (N_15669,N_14448,N_14791);
nand U15670 (N_15670,N_14980,N_14474);
nor U15671 (N_15671,N_14992,N_14149);
and U15672 (N_15672,N_14431,N_14982);
nor U15673 (N_15673,N_14714,N_14907);
nor U15674 (N_15674,N_14896,N_14647);
nor U15675 (N_15675,N_14546,N_14589);
nor U15676 (N_15676,N_14170,N_14658);
or U15677 (N_15677,N_14148,N_14847);
and U15678 (N_15678,N_14359,N_14882);
or U15679 (N_15679,N_14454,N_14425);
xor U15680 (N_15680,N_14989,N_14356);
xnor U15681 (N_15681,N_14182,N_14329);
nor U15682 (N_15682,N_14537,N_14217);
or U15683 (N_15683,N_14077,N_14307);
nand U15684 (N_15684,N_14973,N_14892);
xnor U15685 (N_15685,N_14173,N_14488);
and U15686 (N_15686,N_14287,N_14501);
or U15687 (N_15687,N_14784,N_14738);
or U15688 (N_15688,N_14222,N_14454);
and U15689 (N_15689,N_14875,N_14446);
nand U15690 (N_15690,N_14129,N_14035);
or U15691 (N_15691,N_14755,N_14154);
xor U15692 (N_15692,N_14973,N_14787);
nand U15693 (N_15693,N_14047,N_14832);
nand U15694 (N_15694,N_14176,N_14953);
nor U15695 (N_15695,N_14844,N_14201);
nand U15696 (N_15696,N_14591,N_14044);
nand U15697 (N_15697,N_14576,N_14278);
and U15698 (N_15698,N_14294,N_14638);
xnor U15699 (N_15699,N_14058,N_14977);
xor U15700 (N_15700,N_14893,N_14758);
xor U15701 (N_15701,N_14494,N_14942);
nor U15702 (N_15702,N_14471,N_14377);
nand U15703 (N_15703,N_14985,N_14702);
or U15704 (N_15704,N_14884,N_14661);
or U15705 (N_15705,N_14357,N_14403);
nor U15706 (N_15706,N_14321,N_14815);
and U15707 (N_15707,N_14952,N_14819);
and U15708 (N_15708,N_14999,N_14785);
and U15709 (N_15709,N_14266,N_14648);
nor U15710 (N_15710,N_14464,N_14999);
nor U15711 (N_15711,N_14325,N_14111);
nand U15712 (N_15712,N_14246,N_14881);
xnor U15713 (N_15713,N_14777,N_14062);
or U15714 (N_15714,N_14715,N_14361);
and U15715 (N_15715,N_14545,N_14779);
and U15716 (N_15716,N_14590,N_14199);
nand U15717 (N_15717,N_14208,N_14925);
or U15718 (N_15718,N_14059,N_14135);
and U15719 (N_15719,N_14151,N_14712);
xor U15720 (N_15720,N_14116,N_14405);
and U15721 (N_15721,N_14055,N_14510);
and U15722 (N_15722,N_14642,N_14734);
and U15723 (N_15723,N_14974,N_14713);
xnor U15724 (N_15724,N_14153,N_14868);
xor U15725 (N_15725,N_14490,N_14397);
nor U15726 (N_15726,N_14824,N_14947);
nor U15727 (N_15727,N_14975,N_14069);
and U15728 (N_15728,N_14656,N_14849);
and U15729 (N_15729,N_14764,N_14532);
and U15730 (N_15730,N_14003,N_14283);
nand U15731 (N_15731,N_14517,N_14444);
or U15732 (N_15732,N_14296,N_14373);
xor U15733 (N_15733,N_14185,N_14617);
xnor U15734 (N_15734,N_14901,N_14290);
nand U15735 (N_15735,N_14939,N_14800);
or U15736 (N_15736,N_14177,N_14455);
and U15737 (N_15737,N_14488,N_14796);
or U15738 (N_15738,N_14175,N_14298);
nand U15739 (N_15739,N_14503,N_14511);
or U15740 (N_15740,N_14593,N_14112);
nand U15741 (N_15741,N_14203,N_14880);
nor U15742 (N_15742,N_14167,N_14043);
and U15743 (N_15743,N_14500,N_14793);
or U15744 (N_15744,N_14272,N_14686);
xnor U15745 (N_15745,N_14960,N_14056);
or U15746 (N_15746,N_14903,N_14958);
nor U15747 (N_15747,N_14067,N_14380);
nand U15748 (N_15748,N_14414,N_14359);
and U15749 (N_15749,N_14454,N_14359);
and U15750 (N_15750,N_14955,N_14329);
xor U15751 (N_15751,N_14965,N_14535);
xnor U15752 (N_15752,N_14934,N_14250);
nor U15753 (N_15753,N_14667,N_14048);
nor U15754 (N_15754,N_14884,N_14637);
or U15755 (N_15755,N_14335,N_14524);
nor U15756 (N_15756,N_14963,N_14598);
nor U15757 (N_15757,N_14686,N_14343);
or U15758 (N_15758,N_14167,N_14463);
xnor U15759 (N_15759,N_14011,N_14216);
xor U15760 (N_15760,N_14030,N_14714);
nand U15761 (N_15761,N_14415,N_14121);
or U15762 (N_15762,N_14773,N_14484);
and U15763 (N_15763,N_14055,N_14777);
and U15764 (N_15764,N_14207,N_14693);
nor U15765 (N_15765,N_14461,N_14566);
xor U15766 (N_15766,N_14133,N_14596);
nor U15767 (N_15767,N_14941,N_14243);
xor U15768 (N_15768,N_14272,N_14580);
or U15769 (N_15769,N_14543,N_14053);
xnor U15770 (N_15770,N_14330,N_14417);
or U15771 (N_15771,N_14811,N_14151);
and U15772 (N_15772,N_14147,N_14394);
nand U15773 (N_15773,N_14055,N_14680);
nor U15774 (N_15774,N_14418,N_14632);
nand U15775 (N_15775,N_14740,N_14310);
and U15776 (N_15776,N_14983,N_14229);
and U15777 (N_15777,N_14005,N_14919);
nor U15778 (N_15778,N_14089,N_14250);
nor U15779 (N_15779,N_14364,N_14681);
or U15780 (N_15780,N_14036,N_14678);
xor U15781 (N_15781,N_14105,N_14693);
nand U15782 (N_15782,N_14013,N_14437);
and U15783 (N_15783,N_14662,N_14579);
nand U15784 (N_15784,N_14061,N_14988);
and U15785 (N_15785,N_14084,N_14913);
or U15786 (N_15786,N_14439,N_14339);
xnor U15787 (N_15787,N_14934,N_14909);
and U15788 (N_15788,N_14897,N_14356);
xnor U15789 (N_15789,N_14996,N_14787);
nor U15790 (N_15790,N_14490,N_14464);
or U15791 (N_15791,N_14294,N_14221);
and U15792 (N_15792,N_14838,N_14864);
nor U15793 (N_15793,N_14532,N_14379);
xnor U15794 (N_15794,N_14547,N_14167);
nand U15795 (N_15795,N_14901,N_14371);
nand U15796 (N_15796,N_14248,N_14793);
nor U15797 (N_15797,N_14594,N_14429);
xnor U15798 (N_15798,N_14973,N_14038);
xnor U15799 (N_15799,N_14098,N_14632);
or U15800 (N_15800,N_14302,N_14896);
nor U15801 (N_15801,N_14495,N_14712);
and U15802 (N_15802,N_14287,N_14606);
nor U15803 (N_15803,N_14352,N_14192);
or U15804 (N_15804,N_14770,N_14091);
or U15805 (N_15805,N_14561,N_14973);
and U15806 (N_15806,N_14940,N_14880);
xnor U15807 (N_15807,N_14105,N_14814);
or U15808 (N_15808,N_14724,N_14854);
nor U15809 (N_15809,N_14981,N_14366);
or U15810 (N_15810,N_14983,N_14981);
nand U15811 (N_15811,N_14156,N_14559);
nor U15812 (N_15812,N_14315,N_14276);
nand U15813 (N_15813,N_14730,N_14036);
nor U15814 (N_15814,N_14453,N_14708);
nor U15815 (N_15815,N_14448,N_14351);
nor U15816 (N_15816,N_14334,N_14347);
nor U15817 (N_15817,N_14096,N_14094);
or U15818 (N_15818,N_14559,N_14303);
or U15819 (N_15819,N_14714,N_14598);
xor U15820 (N_15820,N_14197,N_14292);
or U15821 (N_15821,N_14130,N_14321);
or U15822 (N_15822,N_14292,N_14337);
or U15823 (N_15823,N_14911,N_14057);
nand U15824 (N_15824,N_14490,N_14652);
xnor U15825 (N_15825,N_14806,N_14594);
xnor U15826 (N_15826,N_14517,N_14676);
nor U15827 (N_15827,N_14722,N_14680);
and U15828 (N_15828,N_14111,N_14516);
or U15829 (N_15829,N_14401,N_14927);
nand U15830 (N_15830,N_14387,N_14876);
nor U15831 (N_15831,N_14293,N_14351);
nand U15832 (N_15832,N_14638,N_14225);
xor U15833 (N_15833,N_14077,N_14676);
nor U15834 (N_15834,N_14322,N_14727);
nand U15835 (N_15835,N_14038,N_14102);
or U15836 (N_15836,N_14735,N_14675);
nand U15837 (N_15837,N_14421,N_14343);
nand U15838 (N_15838,N_14131,N_14134);
xnor U15839 (N_15839,N_14142,N_14321);
and U15840 (N_15840,N_14086,N_14900);
xor U15841 (N_15841,N_14716,N_14084);
or U15842 (N_15842,N_14427,N_14739);
or U15843 (N_15843,N_14536,N_14084);
xor U15844 (N_15844,N_14661,N_14920);
or U15845 (N_15845,N_14397,N_14657);
xor U15846 (N_15846,N_14603,N_14925);
nor U15847 (N_15847,N_14770,N_14621);
nand U15848 (N_15848,N_14525,N_14709);
nand U15849 (N_15849,N_14629,N_14518);
or U15850 (N_15850,N_14639,N_14726);
and U15851 (N_15851,N_14843,N_14616);
and U15852 (N_15852,N_14940,N_14496);
nand U15853 (N_15853,N_14351,N_14682);
xor U15854 (N_15854,N_14141,N_14702);
and U15855 (N_15855,N_14670,N_14011);
or U15856 (N_15856,N_14502,N_14603);
or U15857 (N_15857,N_14188,N_14235);
or U15858 (N_15858,N_14415,N_14573);
xor U15859 (N_15859,N_14924,N_14752);
xor U15860 (N_15860,N_14030,N_14992);
or U15861 (N_15861,N_14506,N_14538);
and U15862 (N_15862,N_14678,N_14848);
nor U15863 (N_15863,N_14399,N_14155);
and U15864 (N_15864,N_14967,N_14660);
nand U15865 (N_15865,N_14748,N_14459);
and U15866 (N_15866,N_14868,N_14876);
and U15867 (N_15867,N_14107,N_14027);
or U15868 (N_15868,N_14179,N_14430);
nor U15869 (N_15869,N_14192,N_14441);
nand U15870 (N_15870,N_14988,N_14278);
nand U15871 (N_15871,N_14700,N_14706);
or U15872 (N_15872,N_14885,N_14024);
xor U15873 (N_15873,N_14620,N_14006);
nor U15874 (N_15874,N_14635,N_14043);
nand U15875 (N_15875,N_14970,N_14797);
nand U15876 (N_15876,N_14595,N_14050);
xor U15877 (N_15877,N_14978,N_14637);
and U15878 (N_15878,N_14286,N_14052);
and U15879 (N_15879,N_14672,N_14653);
or U15880 (N_15880,N_14511,N_14751);
nor U15881 (N_15881,N_14442,N_14589);
or U15882 (N_15882,N_14927,N_14836);
or U15883 (N_15883,N_14706,N_14820);
xor U15884 (N_15884,N_14681,N_14624);
nand U15885 (N_15885,N_14042,N_14548);
xnor U15886 (N_15886,N_14323,N_14463);
nand U15887 (N_15887,N_14042,N_14525);
and U15888 (N_15888,N_14899,N_14428);
nand U15889 (N_15889,N_14513,N_14164);
nor U15890 (N_15890,N_14273,N_14703);
and U15891 (N_15891,N_14597,N_14046);
xor U15892 (N_15892,N_14195,N_14991);
or U15893 (N_15893,N_14908,N_14486);
or U15894 (N_15894,N_14247,N_14171);
and U15895 (N_15895,N_14510,N_14171);
xor U15896 (N_15896,N_14746,N_14596);
or U15897 (N_15897,N_14700,N_14306);
nand U15898 (N_15898,N_14940,N_14244);
and U15899 (N_15899,N_14229,N_14381);
xor U15900 (N_15900,N_14002,N_14557);
xnor U15901 (N_15901,N_14695,N_14479);
and U15902 (N_15902,N_14448,N_14312);
nand U15903 (N_15903,N_14537,N_14136);
nand U15904 (N_15904,N_14053,N_14712);
and U15905 (N_15905,N_14384,N_14235);
nor U15906 (N_15906,N_14950,N_14594);
and U15907 (N_15907,N_14404,N_14303);
or U15908 (N_15908,N_14973,N_14746);
nor U15909 (N_15909,N_14500,N_14453);
nand U15910 (N_15910,N_14014,N_14266);
nor U15911 (N_15911,N_14175,N_14656);
nor U15912 (N_15912,N_14633,N_14274);
nand U15913 (N_15913,N_14267,N_14018);
nor U15914 (N_15914,N_14466,N_14677);
or U15915 (N_15915,N_14311,N_14894);
nor U15916 (N_15916,N_14628,N_14596);
nand U15917 (N_15917,N_14872,N_14749);
and U15918 (N_15918,N_14028,N_14516);
nand U15919 (N_15919,N_14376,N_14132);
xor U15920 (N_15920,N_14949,N_14436);
nand U15921 (N_15921,N_14040,N_14392);
nor U15922 (N_15922,N_14802,N_14429);
or U15923 (N_15923,N_14301,N_14763);
or U15924 (N_15924,N_14345,N_14605);
or U15925 (N_15925,N_14053,N_14290);
and U15926 (N_15926,N_14718,N_14926);
and U15927 (N_15927,N_14022,N_14497);
xnor U15928 (N_15928,N_14907,N_14429);
nand U15929 (N_15929,N_14448,N_14853);
or U15930 (N_15930,N_14133,N_14048);
nand U15931 (N_15931,N_14419,N_14166);
nand U15932 (N_15932,N_14655,N_14040);
or U15933 (N_15933,N_14182,N_14217);
nor U15934 (N_15934,N_14520,N_14954);
xor U15935 (N_15935,N_14850,N_14986);
and U15936 (N_15936,N_14436,N_14278);
nand U15937 (N_15937,N_14567,N_14422);
xnor U15938 (N_15938,N_14107,N_14317);
and U15939 (N_15939,N_14838,N_14575);
nor U15940 (N_15940,N_14962,N_14947);
or U15941 (N_15941,N_14794,N_14240);
xnor U15942 (N_15942,N_14600,N_14549);
nand U15943 (N_15943,N_14873,N_14158);
xor U15944 (N_15944,N_14590,N_14881);
and U15945 (N_15945,N_14709,N_14105);
and U15946 (N_15946,N_14928,N_14709);
or U15947 (N_15947,N_14723,N_14745);
or U15948 (N_15948,N_14477,N_14272);
and U15949 (N_15949,N_14004,N_14074);
or U15950 (N_15950,N_14546,N_14192);
xnor U15951 (N_15951,N_14163,N_14680);
xnor U15952 (N_15952,N_14613,N_14897);
nor U15953 (N_15953,N_14891,N_14276);
xor U15954 (N_15954,N_14717,N_14715);
xor U15955 (N_15955,N_14490,N_14835);
nor U15956 (N_15956,N_14225,N_14496);
and U15957 (N_15957,N_14119,N_14477);
xnor U15958 (N_15958,N_14423,N_14736);
or U15959 (N_15959,N_14962,N_14046);
nand U15960 (N_15960,N_14076,N_14931);
or U15961 (N_15961,N_14010,N_14693);
or U15962 (N_15962,N_14848,N_14760);
and U15963 (N_15963,N_14778,N_14878);
and U15964 (N_15964,N_14022,N_14052);
xor U15965 (N_15965,N_14079,N_14471);
nor U15966 (N_15966,N_14495,N_14927);
and U15967 (N_15967,N_14944,N_14119);
nand U15968 (N_15968,N_14284,N_14609);
xnor U15969 (N_15969,N_14199,N_14749);
or U15970 (N_15970,N_14538,N_14114);
xor U15971 (N_15971,N_14242,N_14178);
or U15972 (N_15972,N_14510,N_14101);
xnor U15973 (N_15973,N_14493,N_14797);
or U15974 (N_15974,N_14938,N_14460);
or U15975 (N_15975,N_14043,N_14630);
or U15976 (N_15976,N_14775,N_14386);
and U15977 (N_15977,N_14561,N_14720);
xnor U15978 (N_15978,N_14841,N_14477);
or U15979 (N_15979,N_14548,N_14032);
nand U15980 (N_15980,N_14624,N_14925);
or U15981 (N_15981,N_14292,N_14059);
nor U15982 (N_15982,N_14357,N_14131);
nor U15983 (N_15983,N_14071,N_14576);
and U15984 (N_15984,N_14088,N_14204);
xnor U15985 (N_15985,N_14803,N_14818);
and U15986 (N_15986,N_14294,N_14478);
nand U15987 (N_15987,N_14918,N_14493);
xnor U15988 (N_15988,N_14604,N_14829);
and U15989 (N_15989,N_14998,N_14560);
and U15990 (N_15990,N_14369,N_14149);
nor U15991 (N_15991,N_14779,N_14187);
or U15992 (N_15992,N_14254,N_14696);
nand U15993 (N_15993,N_14452,N_14033);
and U15994 (N_15994,N_14216,N_14789);
xor U15995 (N_15995,N_14846,N_14803);
xor U15996 (N_15996,N_14105,N_14498);
xor U15997 (N_15997,N_14657,N_14586);
nor U15998 (N_15998,N_14832,N_14577);
nor U15999 (N_15999,N_14701,N_14900);
xnor U16000 (N_16000,N_15973,N_15750);
nand U16001 (N_16001,N_15134,N_15563);
nand U16002 (N_16002,N_15039,N_15330);
xor U16003 (N_16003,N_15608,N_15775);
nand U16004 (N_16004,N_15206,N_15865);
xnor U16005 (N_16005,N_15731,N_15263);
and U16006 (N_16006,N_15370,N_15672);
nor U16007 (N_16007,N_15689,N_15985);
nor U16008 (N_16008,N_15296,N_15033);
xnor U16009 (N_16009,N_15368,N_15711);
nor U16010 (N_16010,N_15778,N_15416);
and U16011 (N_16011,N_15746,N_15025);
nor U16012 (N_16012,N_15958,N_15496);
and U16013 (N_16013,N_15392,N_15990);
and U16014 (N_16014,N_15571,N_15361);
nand U16015 (N_16015,N_15446,N_15929);
nor U16016 (N_16016,N_15120,N_15481);
and U16017 (N_16017,N_15139,N_15908);
nor U16018 (N_16018,N_15310,N_15472);
nand U16019 (N_16019,N_15390,N_15708);
and U16020 (N_16020,N_15900,N_15680);
nand U16021 (N_16021,N_15088,N_15534);
xnor U16022 (N_16022,N_15270,N_15986);
xor U16023 (N_16023,N_15308,N_15739);
nor U16024 (N_16024,N_15628,N_15381);
and U16025 (N_16025,N_15597,N_15029);
xor U16026 (N_16026,N_15523,N_15978);
nand U16027 (N_16027,N_15452,N_15465);
and U16028 (N_16028,N_15313,N_15433);
xor U16029 (N_16029,N_15283,N_15478);
nor U16030 (N_16030,N_15982,N_15076);
or U16031 (N_16031,N_15826,N_15605);
or U16032 (N_16032,N_15410,N_15871);
or U16033 (N_16033,N_15664,N_15437);
or U16034 (N_16034,N_15801,N_15273);
xnor U16035 (N_16035,N_15227,N_15872);
xnor U16036 (N_16036,N_15339,N_15143);
xor U16037 (N_16037,N_15742,N_15524);
or U16038 (N_16038,N_15972,N_15948);
and U16039 (N_16039,N_15526,N_15618);
and U16040 (N_16040,N_15650,N_15773);
or U16041 (N_16041,N_15189,N_15841);
xor U16042 (N_16042,N_15312,N_15417);
and U16043 (N_16043,N_15629,N_15464);
xor U16044 (N_16044,N_15490,N_15087);
and U16045 (N_16045,N_15549,N_15516);
nor U16046 (N_16046,N_15503,N_15401);
nor U16047 (N_16047,N_15395,N_15558);
or U16048 (N_16048,N_15870,N_15694);
nor U16049 (N_16049,N_15202,N_15645);
xor U16050 (N_16050,N_15073,N_15554);
xor U16051 (N_16051,N_15585,N_15696);
or U16052 (N_16052,N_15583,N_15819);
nor U16053 (N_16053,N_15932,N_15808);
nand U16054 (N_16054,N_15574,N_15068);
or U16055 (N_16055,N_15935,N_15785);
nor U16056 (N_16056,N_15107,N_15041);
nand U16057 (N_16057,N_15665,N_15001);
nor U16058 (N_16058,N_15745,N_15250);
nand U16059 (N_16059,N_15406,N_15910);
nand U16060 (N_16060,N_15722,N_15561);
or U16061 (N_16061,N_15705,N_15700);
and U16062 (N_16062,N_15324,N_15649);
xor U16063 (N_16063,N_15881,N_15164);
nor U16064 (N_16064,N_15850,N_15196);
nor U16065 (N_16065,N_15514,N_15853);
xnor U16066 (N_16066,N_15166,N_15398);
nand U16067 (N_16067,N_15342,N_15971);
or U16068 (N_16068,N_15764,N_15765);
nor U16069 (N_16069,N_15170,N_15737);
or U16070 (N_16070,N_15440,N_15993);
xnor U16071 (N_16071,N_15385,N_15444);
or U16072 (N_16072,N_15805,N_15060);
nand U16073 (N_16073,N_15278,N_15412);
nor U16074 (N_16074,N_15218,N_15100);
nor U16075 (N_16075,N_15491,N_15732);
or U16076 (N_16076,N_15506,N_15083);
nand U16077 (N_16077,N_15615,N_15197);
xor U16078 (N_16078,N_15579,N_15424);
nor U16079 (N_16079,N_15316,N_15955);
nor U16080 (N_16080,N_15432,N_15251);
nand U16081 (N_16081,N_15034,N_15695);
xnor U16082 (N_16082,N_15415,N_15710);
nand U16083 (N_16083,N_15353,N_15787);
nor U16084 (N_16084,N_15008,N_15822);
nor U16085 (N_16085,N_15866,N_15730);
or U16086 (N_16086,N_15341,N_15484);
nor U16087 (N_16087,N_15788,N_15726);
xor U16088 (N_16088,N_15428,N_15755);
nor U16089 (N_16089,N_15640,N_15691);
nor U16090 (N_16090,N_15631,N_15169);
or U16091 (N_16091,N_15586,N_15109);
and U16092 (N_16092,N_15847,N_15079);
nor U16093 (N_16093,N_15272,N_15002);
xnor U16094 (N_16094,N_15494,N_15223);
or U16095 (N_16095,N_15630,N_15091);
xor U16096 (N_16096,N_15821,N_15714);
xor U16097 (N_16097,N_15147,N_15204);
nand U16098 (N_16098,N_15936,N_15727);
xnor U16099 (N_16099,N_15889,N_15358);
xnor U16100 (N_16100,N_15386,N_15243);
or U16101 (N_16101,N_15562,N_15280);
xor U16102 (N_16102,N_15566,N_15954);
xor U16103 (N_16103,N_15071,N_15208);
or U16104 (N_16104,N_15102,N_15125);
xor U16105 (N_16105,N_15212,N_15620);
xnor U16106 (N_16106,N_15048,N_15167);
xnor U16107 (N_16107,N_15413,N_15439);
and U16108 (N_16108,N_15776,N_15944);
xor U16109 (N_16109,N_15816,N_15837);
nand U16110 (N_16110,N_15876,N_15698);
nor U16111 (N_16111,N_15019,N_15303);
or U16112 (N_16112,N_15565,N_15262);
xor U16113 (N_16113,N_15495,N_15610);
nor U16114 (N_16114,N_15824,N_15422);
nor U16115 (N_16115,N_15090,N_15271);
and U16116 (N_16116,N_15797,N_15789);
xor U16117 (N_16117,N_15364,N_15895);
or U16118 (N_16118,N_15111,N_15298);
and U16119 (N_16119,N_15892,N_15857);
or U16120 (N_16120,N_15219,N_15854);
and U16121 (N_16121,N_15477,N_15532);
nand U16122 (N_16122,N_15687,N_15080);
nand U16123 (N_16123,N_15456,N_15753);
nand U16124 (N_16124,N_15930,N_15793);
nand U16125 (N_16125,N_15810,N_15114);
and U16126 (N_16126,N_15966,N_15836);
and U16127 (N_16127,N_15814,N_15177);
nand U16128 (N_16128,N_15355,N_15551);
nor U16129 (N_16129,N_15180,N_15724);
nand U16130 (N_16130,N_15407,N_15042);
or U16131 (N_16131,N_15337,N_15688);
or U16132 (N_16132,N_15072,N_15252);
xor U16133 (N_16133,N_15749,N_15338);
or U16134 (N_16134,N_15307,N_15423);
nand U16135 (N_16135,N_15183,N_15927);
or U16136 (N_16136,N_15205,N_15969);
or U16137 (N_16137,N_15149,N_15301);
and U16138 (N_16138,N_15030,N_15634);
or U16139 (N_16139,N_15659,N_15064);
or U16140 (N_16140,N_15038,N_15633);
xnor U16141 (N_16141,N_15233,N_15885);
or U16142 (N_16142,N_15720,N_15425);
or U16143 (N_16143,N_15480,N_15070);
or U16144 (N_16144,N_15614,N_15903);
or U16145 (N_16145,N_15146,N_15589);
and U16146 (N_16146,N_15774,N_15455);
and U16147 (N_16147,N_15352,N_15616);
nand U16148 (N_16148,N_15598,N_15128);
nand U16149 (N_16149,N_15811,N_15334);
or U16150 (N_16150,N_15241,N_15917);
nor U16151 (N_16151,N_15040,N_15284);
nand U16152 (N_16152,N_15124,N_15254);
and U16153 (N_16153,N_15117,N_15305);
and U16154 (N_16154,N_15436,N_15158);
nor U16155 (N_16155,N_15926,N_15832);
nand U16156 (N_16156,N_15264,N_15825);
nand U16157 (N_16157,N_15427,N_15581);
or U16158 (N_16158,N_15995,N_15479);
nor U16159 (N_16159,N_15093,N_15609);
nand U16160 (N_16160,N_15289,N_15131);
nor U16161 (N_16161,N_15913,N_15260);
nor U16162 (N_16162,N_15539,N_15976);
xor U16163 (N_16163,N_15956,N_15999);
nor U16164 (N_16164,N_15621,N_15611);
xor U16165 (N_16165,N_15098,N_15568);
and U16166 (N_16166,N_15396,N_15624);
nand U16167 (N_16167,N_15367,N_15761);
nand U16168 (N_16168,N_15584,N_15096);
nor U16169 (N_16169,N_15962,N_15528);
nand U16170 (N_16170,N_15894,N_15261);
nand U16171 (N_16171,N_15815,N_15031);
and U16172 (N_16172,N_15855,N_15522);
xor U16173 (N_16173,N_15319,N_15820);
nand U16174 (N_16174,N_15372,N_15757);
xor U16175 (N_16175,N_15809,N_15612);
nand U16176 (N_16176,N_15763,N_15045);
nor U16177 (N_16177,N_15201,N_15709);
or U16178 (N_16178,N_15601,N_15545);
xor U16179 (N_16179,N_15914,N_15943);
nor U16180 (N_16180,N_15759,N_15781);
or U16181 (N_16181,N_15046,N_15302);
nand U16182 (N_16182,N_15660,N_15622);
nand U16183 (N_16183,N_15741,N_15678);
nor U16184 (N_16184,N_15987,N_15642);
nor U16185 (N_16185,N_15207,N_15572);
xnor U16186 (N_16186,N_15027,N_15178);
or U16187 (N_16187,N_15964,N_15460);
and U16188 (N_16188,N_15663,N_15834);
and U16189 (N_16189,N_15105,N_15486);
nand U16190 (N_16190,N_15487,N_15285);
or U16191 (N_16191,N_15101,N_15179);
or U16192 (N_16192,N_15356,N_15662);
nor U16193 (N_16193,N_15823,N_15217);
xnor U16194 (N_16194,N_15081,N_15553);
or U16195 (N_16195,N_15383,N_15783);
nor U16196 (N_16196,N_15991,N_15963);
or U16197 (N_16197,N_15023,N_15018);
or U16198 (N_16198,N_15276,N_15915);
or U16199 (N_16199,N_15151,N_15475);
nor U16200 (N_16200,N_15216,N_15320);
nor U16201 (N_16201,N_15132,N_15258);
and U16202 (N_16202,N_15391,N_15028);
nor U16203 (N_16203,N_15235,N_15074);
and U16204 (N_16204,N_15454,N_15968);
or U16205 (N_16205,N_15559,N_15552);
nand U16206 (N_16206,N_15239,N_15032);
nand U16207 (N_16207,N_15082,N_15403);
nand U16208 (N_16208,N_15902,N_15118);
and U16209 (N_16209,N_15817,N_15807);
nand U16210 (N_16210,N_15156,N_15378);
or U16211 (N_16211,N_15875,N_15803);
or U16212 (N_16212,N_15482,N_15666);
and U16213 (N_16213,N_15225,N_15136);
nor U16214 (N_16214,N_15248,N_15861);
nand U16215 (N_16215,N_15668,N_15014);
xor U16216 (N_16216,N_15468,N_15186);
xor U16217 (N_16217,N_15744,N_15097);
or U16218 (N_16218,N_15939,N_15512);
or U16219 (N_16219,N_15162,N_15141);
nand U16220 (N_16220,N_15343,N_15671);
and U16221 (N_16221,N_15362,N_15473);
nor U16222 (N_16222,N_15144,N_15347);
and U16223 (N_16223,N_15443,N_15508);
and U16224 (N_16224,N_15379,N_15573);
nand U16225 (N_16225,N_15268,N_15654);
or U16226 (N_16226,N_15013,N_15901);
and U16227 (N_16227,N_15684,N_15004);
nand U16228 (N_16228,N_15527,N_15920);
nand U16229 (N_16229,N_15828,N_15474);
nor U16230 (N_16230,N_15288,N_15960);
xor U16231 (N_16231,N_15274,N_15569);
and U16232 (N_16232,N_15537,N_15835);
xor U16233 (N_16233,N_15287,N_15992);
nand U16234 (N_16234,N_15214,N_15838);
and U16235 (N_16235,N_15582,N_15595);
and U16236 (N_16236,N_15829,N_15981);
or U16237 (N_16237,N_15122,N_15716);
or U16238 (N_16238,N_15844,N_15348);
and U16239 (N_16239,N_15578,N_15193);
and U16240 (N_16240,N_15500,N_15567);
xor U16241 (N_16241,N_15632,N_15556);
and U16242 (N_16242,N_15904,N_15215);
nor U16243 (N_16243,N_15542,N_15931);
and U16244 (N_16244,N_15536,N_15269);
and U16245 (N_16245,N_15898,N_15845);
or U16246 (N_16246,N_15617,N_15951);
nor U16247 (N_16247,N_15770,N_15492);
nor U16248 (N_16248,N_15376,N_15674);
or U16249 (N_16249,N_15326,N_15232);
xnor U16250 (N_16250,N_15110,N_15648);
nand U16251 (N_16251,N_15445,N_15513);
nor U16252 (N_16252,N_15575,N_15676);
or U16253 (N_16253,N_15728,N_15505);
nor U16254 (N_16254,N_15723,N_15967);
or U16255 (N_16255,N_15106,N_15497);
or U16256 (N_16256,N_15719,N_15300);
and U16257 (N_16257,N_15449,N_15812);
or U16258 (N_16258,N_15952,N_15880);
xor U16259 (N_16259,N_15600,N_15485);
nand U16260 (N_16260,N_15588,N_15418);
nor U16261 (N_16261,N_15488,N_15521);
or U16262 (N_16262,N_15246,N_15957);
xnor U16263 (N_16263,N_15380,N_15762);
nand U16264 (N_16264,N_15056,N_15044);
or U16265 (N_16265,N_15063,N_15461);
or U16266 (N_16266,N_15290,N_15813);
nand U16267 (N_16267,N_15603,N_15275);
and U16268 (N_16268,N_15796,N_15831);
nand U16269 (N_16269,N_15113,N_15509);
nand U16270 (N_16270,N_15743,N_15493);
xnor U16271 (N_16271,N_15161,N_15667);
xnor U16272 (N_16272,N_15007,N_15069);
nor U16273 (N_16273,N_15476,N_15721);
and U16274 (N_16274,N_15245,N_15409);
or U16275 (N_16275,N_15546,N_15682);
nand U16276 (N_16276,N_15679,N_15635);
and U16277 (N_16277,N_15345,N_15644);
nand U16278 (N_16278,N_15129,N_15555);
and U16279 (N_16279,N_15525,N_15365);
nor U16280 (N_16280,N_15863,N_15818);
nand U16281 (N_16281,N_15230,N_15085);
xor U16282 (N_16282,N_15874,N_15879);
nor U16283 (N_16283,N_15692,N_15108);
nor U16284 (N_16284,N_15827,N_15655);
and U16285 (N_16285,N_15411,N_15923);
and U16286 (N_16286,N_15893,N_15800);
nor U16287 (N_16287,N_15171,N_15974);
and U16288 (N_16288,N_15909,N_15947);
or U16289 (N_16289,N_15231,N_15518);
or U16290 (N_16290,N_15035,N_15849);
and U16291 (N_16291,N_15145,N_15697);
xor U16292 (N_16292,N_15184,N_15317);
nand U16293 (N_16293,N_15733,N_15606);
xnor U16294 (N_16294,N_15115,N_15602);
nor U16295 (N_16295,N_15388,N_15699);
nand U16296 (N_16296,N_15771,N_15344);
nand U16297 (N_16297,N_15751,N_15089);
xnor U16298 (N_16298,N_15587,N_15195);
xor U16299 (N_16299,N_15123,N_15061);
and U16300 (N_16300,N_15942,N_15349);
nor U16301 (N_16301,N_15483,N_15519);
and U16302 (N_16302,N_15191,N_15596);
and U16303 (N_16303,N_15883,N_15306);
and U16304 (N_16304,N_15627,N_15099);
nand U16305 (N_16305,N_15237,N_15703);
or U16306 (N_16306,N_15229,N_15658);
nor U16307 (N_16307,N_15053,N_15541);
xnor U16308 (N_16308,N_15511,N_15389);
nand U16309 (N_16309,N_15983,N_15938);
and U16310 (N_16310,N_15921,N_15086);
or U16311 (N_16311,N_15159,N_15127);
or U16312 (N_16312,N_15176,N_15661);
xnor U16313 (N_16313,N_15138,N_15980);
and U16314 (N_16314,N_15848,N_15150);
xnor U16315 (N_16315,N_15154,N_15092);
xnor U16316 (N_16316,N_15458,N_15222);
nand U16317 (N_16317,N_15238,N_15887);
nand U16318 (N_16318,N_15095,N_15256);
nand U16319 (N_16319,N_15209,N_15314);
nand U16320 (N_16320,N_15540,N_15673);
xnor U16321 (N_16321,N_15970,N_15447);
nand U16322 (N_16322,N_15408,N_15340);
or U16323 (N_16323,N_15188,N_15160);
xor U16324 (N_16324,N_15802,N_15538);
nor U16325 (N_16325,N_15979,N_15897);
nor U16326 (N_16326,N_15414,N_15748);
xnor U16327 (N_16327,N_15840,N_15756);
nand U16328 (N_16328,N_15804,N_15471);
nand U16329 (N_16329,N_15639,N_15321);
nand U16330 (N_16330,N_15000,N_15005);
nor U16331 (N_16331,N_15112,N_15148);
and U16332 (N_16332,N_15707,N_15557);
xnor U16333 (N_16333,N_15940,N_15405);
or U16334 (N_16334,N_15911,N_15760);
and U16335 (N_16335,N_15058,N_15706);
nand U16336 (N_16336,N_15309,N_15282);
or U16337 (N_16337,N_15846,N_15182);
nor U16338 (N_16338,N_15419,N_15140);
and U16339 (N_16339,N_15036,N_15366);
xnor U16340 (N_16340,N_15591,N_15011);
nor U16341 (N_16341,N_15996,N_15426);
xnor U16342 (N_16342,N_15043,N_15255);
nand U16343 (N_16343,N_15357,N_15886);
or U16344 (N_16344,N_15890,N_15501);
and U16345 (N_16345,N_15856,N_15022);
xnor U16346 (N_16346,N_15564,N_15758);
nor U16347 (N_16347,N_15172,N_15020);
nor U16348 (N_16348,N_15470,N_15448);
or U16349 (N_16349,N_15950,N_15713);
nand U16350 (N_16350,N_15806,N_15953);
nor U16351 (N_16351,N_15067,N_15830);
nand U16352 (N_16352,N_15626,N_15946);
nand U16353 (N_16353,N_15941,N_15402);
nand U16354 (N_16354,N_15693,N_15531);
and U16355 (N_16355,N_15729,N_15015);
or U16356 (N_16356,N_15675,N_15651);
nand U16357 (N_16357,N_15860,N_15520);
nand U16358 (N_16358,N_15299,N_15570);
xor U16359 (N_16359,N_15924,N_15747);
or U16360 (N_16360,N_15194,N_15322);
nand U16361 (N_16361,N_15670,N_15442);
nor U16362 (N_16362,N_15234,N_15594);
nor U16363 (N_16363,N_15734,N_15690);
nor U16364 (N_16364,N_15152,N_15717);
xnor U16365 (N_16365,N_15315,N_15281);
nand U16366 (N_16366,N_15641,N_15686);
nand U16367 (N_16367,N_15346,N_15049);
xnor U16368 (N_16368,N_15653,N_15293);
xor U16369 (N_16369,N_15989,N_15790);
xnor U16370 (N_16370,N_15604,N_15244);
or U16371 (N_16371,N_15163,N_15652);
nand U16372 (N_16372,N_15017,N_15153);
nor U16373 (N_16373,N_15135,N_15257);
xnor U16374 (N_16374,N_15752,N_15062);
and U16375 (N_16375,N_15187,N_15899);
nor U16376 (N_16376,N_15200,N_15577);
and U16377 (N_16377,N_15791,N_15965);
nor U16378 (N_16378,N_15259,N_15155);
nor U16379 (N_16379,N_15777,N_15253);
nor U16380 (N_16380,N_15051,N_15685);
xor U16381 (N_16381,N_15772,N_15451);
and U16382 (N_16382,N_15780,N_15798);
or U16383 (N_16383,N_15643,N_15740);
nand U16384 (N_16384,N_15453,N_15121);
or U16385 (N_16385,N_15906,N_15912);
nor U16386 (N_16386,N_15323,N_15363);
and U16387 (N_16387,N_15590,N_15236);
xor U16388 (N_16388,N_15794,N_15350);
or U16389 (N_16389,N_15210,N_15116);
xnor U16390 (N_16390,N_15226,N_15701);
nor U16391 (N_16391,N_15718,N_15467);
nand U16392 (N_16392,N_15174,N_15997);
xnor U16393 (N_16393,N_15533,N_15012);
nand U16394 (N_16394,N_15869,N_15977);
xnor U16395 (N_16395,N_15351,N_15499);
nand U16396 (N_16396,N_15400,N_15548);
nor U16397 (N_16397,N_15291,N_15429);
nor U16398 (N_16398,N_15374,N_15868);
xnor U16399 (N_16399,N_15387,N_15457);
and U16400 (N_16400,N_15373,N_15371);
or U16401 (N_16401,N_15438,N_15421);
xnor U16402 (N_16402,N_15420,N_15199);
and U16403 (N_16403,N_15434,N_15656);
xnor U16404 (N_16404,N_15333,N_15304);
nand U16405 (N_16405,N_15896,N_15286);
xor U16406 (N_16406,N_15712,N_15404);
nor U16407 (N_16407,N_15833,N_15297);
nor U16408 (N_16408,N_15021,N_15327);
nor U16409 (N_16409,N_15599,N_15852);
xnor U16410 (N_16410,N_15959,N_15735);
nor U16411 (N_16411,N_15318,N_15619);
or U16412 (N_16412,N_15295,N_15576);
or U16413 (N_16413,N_15916,N_15329);
xor U16414 (N_16414,N_15625,N_15715);
nand U16415 (N_16415,N_15441,N_15075);
and U16416 (N_16416,N_15066,N_15779);
nor U16417 (N_16417,N_15873,N_15907);
nand U16418 (N_16418,N_15328,N_15228);
and U16419 (N_16419,N_15242,N_15360);
and U16420 (N_16420,N_15173,N_15240);
xnor U16421 (N_16421,N_15047,N_15862);
xor U16422 (N_16422,N_15016,N_15037);
and U16423 (N_16423,N_15126,N_15623);
xnor U16424 (N_16424,N_15504,N_15384);
xnor U16425 (N_16425,N_15009,N_15613);
and U16426 (N_16426,N_15767,N_15078);
or U16427 (N_16427,N_15736,N_15399);
and U16428 (N_16428,N_15462,N_15725);
nor U16429 (N_16429,N_15266,N_15331);
and U16430 (N_16430,N_15325,N_15249);
xnor U16431 (N_16431,N_15369,N_15463);
xnor U16432 (N_16432,N_15975,N_15130);
or U16433 (N_16433,N_15919,N_15891);
nor U16434 (N_16434,N_15277,N_15637);
nor U16435 (N_16435,N_15882,N_15190);
nor U16436 (N_16436,N_15181,N_15933);
xor U16437 (N_16437,N_15247,N_15221);
and U16438 (N_16438,N_15292,N_15133);
and U16439 (N_16439,N_15198,N_15510);
nand U16440 (N_16440,N_15646,N_15677);
nand U16441 (N_16441,N_15766,N_15311);
and U16442 (N_16442,N_15168,N_15768);
nor U16443 (N_16443,N_15961,N_15795);
xnor U16444 (N_16444,N_15435,N_15683);
or U16445 (N_16445,N_15430,N_15165);
or U16446 (N_16446,N_15104,N_15592);
xor U16447 (N_16447,N_15265,N_15945);
or U16448 (N_16448,N_15024,N_15026);
and U16449 (N_16449,N_15203,N_15431);
xnor U16450 (N_16450,N_15084,N_15784);
nor U16451 (N_16451,N_15050,N_15636);
nor U16452 (N_16452,N_15354,N_15657);
nand U16453 (N_16453,N_15843,N_15375);
and U16454 (N_16454,N_15517,N_15335);
or U16455 (N_16455,N_15185,N_15103);
nor U16456 (N_16456,N_15055,N_15382);
nand U16457 (N_16457,N_15858,N_15878);
xor U16458 (N_16458,N_15175,N_15934);
and U16459 (N_16459,N_15593,N_15786);
nor U16460 (N_16460,N_15459,N_15754);
xnor U16461 (N_16461,N_15535,N_15998);
nor U16462 (N_16462,N_15450,N_15397);
nand U16463 (N_16463,N_15884,N_15332);
or U16464 (N_16464,N_15769,N_15213);
or U16465 (N_16465,N_15864,N_15647);
and U16466 (N_16466,N_15119,N_15529);
nand U16467 (N_16467,N_15003,N_15065);
nand U16468 (N_16468,N_15543,N_15782);
nand U16469 (N_16469,N_15192,N_15502);
nand U16470 (N_16470,N_15137,N_15547);
nor U16471 (N_16471,N_15792,N_15851);
or U16472 (N_16472,N_15054,N_15738);
nor U16473 (N_16473,N_15550,N_15842);
nand U16474 (N_16474,N_15839,N_15638);
or U16475 (N_16475,N_15607,N_15220);
xor U16476 (N_16476,N_15157,N_15515);
nor U16477 (N_16477,N_15336,N_15294);
nand U16478 (N_16478,N_15211,N_15669);
or U16479 (N_16479,N_15544,N_15918);
nand U16480 (N_16480,N_15704,N_15949);
or U16481 (N_16481,N_15530,N_15988);
or U16482 (N_16482,N_15507,N_15888);
nand U16483 (N_16483,N_15393,N_15867);
xor U16484 (N_16484,N_15359,N_15469);
or U16485 (N_16485,N_15925,N_15994);
and U16486 (N_16486,N_15142,N_15466);
nor U16487 (N_16487,N_15052,N_15928);
nand U16488 (N_16488,N_15006,N_15681);
or U16489 (N_16489,N_15394,N_15279);
and U16490 (N_16490,N_15377,N_15489);
or U16491 (N_16491,N_15922,N_15877);
nor U16492 (N_16492,N_15859,N_15224);
xnor U16493 (N_16493,N_15057,N_15498);
xor U16494 (N_16494,N_15094,N_15560);
xnor U16495 (N_16495,N_15937,N_15905);
nand U16496 (N_16496,N_15984,N_15077);
or U16497 (N_16497,N_15267,N_15799);
nor U16498 (N_16498,N_15010,N_15702);
nor U16499 (N_16499,N_15580,N_15059);
nand U16500 (N_16500,N_15838,N_15802);
and U16501 (N_16501,N_15932,N_15259);
nand U16502 (N_16502,N_15018,N_15204);
xor U16503 (N_16503,N_15509,N_15088);
or U16504 (N_16504,N_15541,N_15006);
nand U16505 (N_16505,N_15237,N_15584);
or U16506 (N_16506,N_15837,N_15365);
or U16507 (N_16507,N_15531,N_15483);
xnor U16508 (N_16508,N_15377,N_15526);
or U16509 (N_16509,N_15589,N_15055);
nand U16510 (N_16510,N_15509,N_15574);
nand U16511 (N_16511,N_15172,N_15957);
and U16512 (N_16512,N_15672,N_15769);
and U16513 (N_16513,N_15189,N_15888);
or U16514 (N_16514,N_15794,N_15765);
xor U16515 (N_16515,N_15234,N_15498);
xnor U16516 (N_16516,N_15356,N_15166);
xnor U16517 (N_16517,N_15807,N_15402);
and U16518 (N_16518,N_15191,N_15823);
nand U16519 (N_16519,N_15688,N_15360);
nor U16520 (N_16520,N_15902,N_15991);
nand U16521 (N_16521,N_15128,N_15800);
and U16522 (N_16522,N_15542,N_15879);
nor U16523 (N_16523,N_15161,N_15651);
and U16524 (N_16524,N_15952,N_15368);
nor U16525 (N_16525,N_15968,N_15310);
or U16526 (N_16526,N_15876,N_15099);
or U16527 (N_16527,N_15930,N_15858);
and U16528 (N_16528,N_15383,N_15453);
xnor U16529 (N_16529,N_15439,N_15485);
nor U16530 (N_16530,N_15616,N_15541);
and U16531 (N_16531,N_15717,N_15081);
xor U16532 (N_16532,N_15020,N_15398);
xnor U16533 (N_16533,N_15273,N_15987);
nand U16534 (N_16534,N_15968,N_15551);
or U16535 (N_16535,N_15927,N_15428);
and U16536 (N_16536,N_15522,N_15736);
xnor U16537 (N_16537,N_15230,N_15358);
xor U16538 (N_16538,N_15491,N_15712);
nor U16539 (N_16539,N_15674,N_15941);
nor U16540 (N_16540,N_15599,N_15413);
and U16541 (N_16541,N_15667,N_15023);
nor U16542 (N_16542,N_15235,N_15897);
or U16543 (N_16543,N_15222,N_15673);
and U16544 (N_16544,N_15647,N_15441);
nor U16545 (N_16545,N_15856,N_15014);
or U16546 (N_16546,N_15553,N_15215);
or U16547 (N_16547,N_15152,N_15470);
or U16548 (N_16548,N_15439,N_15262);
xnor U16549 (N_16549,N_15065,N_15396);
nor U16550 (N_16550,N_15909,N_15179);
and U16551 (N_16551,N_15560,N_15301);
and U16552 (N_16552,N_15419,N_15252);
xnor U16553 (N_16553,N_15400,N_15212);
nand U16554 (N_16554,N_15078,N_15942);
and U16555 (N_16555,N_15698,N_15799);
xnor U16556 (N_16556,N_15624,N_15289);
or U16557 (N_16557,N_15728,N_15036);
nor U16558 (N_16558,N_15286,N_15074);
or U16559 (N_16559,N_15627,N_15947);
nor U16560 (N_16560,N_15403,N_15123);
and U16561 (N_16561,N_15314,N_15120);
xor U16562 (N_16562,N_15996,N_15112);
and U16563 (N_16563,N_15486,N_15991);
or U16564 (N_16564,N_15008,N_15833);
xnor U16565 (N_16565,N_15840,N_15438);
nand U16566 (N_16566,N_15506,N_15913);
nor U16567 (N_16567,N_15768,N_15625);
xnor U16568 (N_16568,N_15382,N_15957);
xnor U16569 (N_16569,N_15471,N_15839);
or U16570 (N_16570,N_15987,N_15654);
nor U16571 (N_16571,N_15057,N_15625);
nand U16572 (N_16572,N_15622,N_15906);
nand U16573 (N_16573,N_15733,N_15624);
nor U16574 (N_16574,N_15526,N_15813);
or U16575 (N_16575,N_15421,N_15413);
and U16576 (N_16576,N_15623,N_15711);
xor U16577 (N_16577,N_15029,N_15355);
and U16578 (N_16578,N_15177,N_15480);
xor U16579 (N_16579,N_15948,N_15191);
xnor U16580 (N_16580,N_15987,N_15942);
nor U16581 (N_16581,N_15200,N_15516);
xnor U16582 (N_16582,N_15171,N_15831);
nor U16583 (N_16583,N_15247,N_15451);
or U16584 (N_16584,N_15431,N_15029);
xnor U16585 (N_16585,N_15511,N_15561);
or U16586 (N_16586,N_15944,N_15716);
and U16587 (N_16587,N_15077,N_15808);
nand U16588 (N_16588,N_15063,N_15232);
or U16589 (N_16589,N_15891,N_15815);
or U16590 (N_16590,N_15288,N_15369);
xor U16591 (N_16591,N_15621,N_15315);
or U16592 (N_16592,N_15139,N_15842);
nor U16593 (N_16593,N_15805,N_15019);
nand U16594 (N_16594,N_15142,N_15273);
and U16595 (N_16595,N_15847,N_15941);
nand U16596 (N_16596,N_15432,N_15285);
xnor U16597 (N_16597,N_15490,N_15581);
and U16598 (N_16598,N_15738,N_15178);
and U16599 (N_16599,N_15610,N_15400);
nor U16600 (N_16600,N_15497,N_15102);
nand U16601 (N_16601,N_15567,N_15004);
nor U16602 (N_16602,N_15374,N_15234);
or U16603 (N_16603,N_15291,N_15184);
and U16604 (N_16604,N_15283,N_15221);
xor U16605 (N_16605,N_15928,N_15413);
xnor U16606 (N_16606,N_15040,N_15236);
or U16607 (N_16607,N_15583,N_15346);
nand U16608 (N_16608,N_15300,N_15747);
and U16609 (N_16609,N_15433,N_15992);
and U16610 (N_16610,N_15482,N_15946);
nand U16611 (N_16611,N_15602,N_15802);
nand U16612 (N_16612,N_15317,N_15629);
nor U16613 (N_16613,N_15731,N_15819);
nand U16614 (N_16614,N_15665,N_15305);
nand U16615 (N_16615,N_15225,N_15185);
nand U16616 (N_16616,N_15153,N_15601);
nand U16617 (N_16617,N_15463,N_15212);
nand U16618 (N_16618,N_15548,N_15016);
and U16619 (N_16619,N_15805,N_15650);
nand U16620 (N_16620,N_15951,N_15453);
and U16621 (N_16621,N_15525,N_15428);
xor U16622 (N_16622,N_15352,N_15433);
nand U16623 (N_16623,N_15964,N_15272);
nor U16624 (N_16624,N_15870,N_15799);
nor U16625 (N_16625,N_15670,N_15245);
and U16626 (N_16626,N_15620,N_15165);
nor U16627 (N_16627,N_15792,N_15881);
nor U16628 (N_16628,N_15913,N_15119);
nand U16629 (N_16629,N_15309,N_15005);
xnor U16630 (N_16630,N_15194,N_15466);
xor U16631 (N_16631,N_15286,N_15292);
xor U16632 (N_16632,N_15663,N_15425);
nand U16633 (N_16633,N_15690,N_15695);
xor U16634 (N_16634,N_15971,N_15403);
nor U16635 (N_16635,N_15177,N_15048);
nor U16636 (N_16636,N_15480,N_15806);
and U16637 (N_16637,N_15526,N_15933);
or U16638 (N_16638,N_15175,N_15774);
and U16639 (N_16639,N_15286,N_15252);
or U16640 (N_16640,N_15874,N_15345);
xnor U16641 (N_16641,N_15834,N_15130);
and U16642 (N_16642,N_15603,N_15339);
xnor U16643 (N_16643,N_15204,N_15200);
and U16644 (N_16644,N_15431,N_15223);
and U16645 (N_16645,N_15627,N_15605);
and U16646 (N_16646,N_15991,N_15840);
nor U16647 (N_16647,N_15323,N_15980);
xor U16648 (N_16648,N_15645,N_15919);
nor U16649 (N_16649,N_15920,N_15662);
or U16650 (N_16650,N_15969,N_15347);
or U16651 (N_16651,N_15294,N_15717);
xnor U16652 (N_16652,N_15512,N_15097);
xor U16653 (N_16653,N_15877,N_15826);
nor U16654 (N_16654,N_15042,N_15275);
and U16655 (N_16655,N_15416,N_15127);
nor U16656 (N_16656,N_15335,N_15313);
xnor U16657 (N_16657,N_15290,N_15804);
xnor U16658 (N_16658,N_15664,N_15484);
xnor U16659 (N_16659,N_15436,N_15985);
nand U16660 (N_16660,N_15979,N_15700);
nor U16661 (N_16661,N_15495,N_15134);
or U16662 (N_16662,N_15092,N_15743);
nor U16663 (N_16663,N_15293,N_15329);
nor U16664 (N_16664,N_15587,N_15156);
nor U16665 (N_16665,N_15234,N_15217);
and U16666 (N_16666,N_15136,N_15162);
xnor U16667 (N_16667,N_15898,N_15307);
nor U16668 (N_16668,N_15085,N_15772);
and U16669 (N_16669,N_15313,N_15463);
nor U16670 (N_16670,N_15458,N_15647);
nor U16671 (N_16671,N_15576,N_15586);
xor U16672 (N_16672,N_15950,N_15936);
nand U16673 (N_16673,N_15107,N_15314);
or U16674 (N_16674,N_15556,N_15744);
xnor U16675 (N_16675,N_15043,N_15491);
xnor U16676 (N_16676,N_15482,N_15133);
or U16677 (N_16677,N_15530,N_15604);
xor U16678 (N_16678,N_15826,N_15264);
xnor U16679 (N_16679,N_15017,N_15708);
or U16680 (N_16680,N_15098,N_15078);
nor U16681 (N_16681,N_15810,N_15423);
xnor U16682 (N_16682,N_15401,N_15086);
and U16683 (N_16683,N_15697,N_15626);
or U16684 (N_16684,N_15434,N_15271);
nand U16685 (N_16685,N_15683,N_15801);
xor U16686 (N_16686,N_15978,N_15892);
nor U16687 (N_16687,N_15962,N_15510);
nor U16688 (N_16688,N_15160,N_15493);
and U16689 (N_16689,N_15838,N_15472);
nor U16690 (N_16690,N_15250,N_15340);
nand U16691 (N_16691,N_15200,N_15664);
nand U16692 (N_16692,N_15908,N_15117);
xnor U16693 (N_16693,N_15347,N_15249);
nor U16694 (N_16694,N_15049,N_15071);
nor U16695 (N_16695,N_15986,N_15006);
nand U16696 (N_16696,N_15629,N_15573);
and U16697 (N_16697,N_15568,N_15813);
and U16698 (N_16698,N_15576,N_15519);
and U16699 (N_16699,N_15323,N_15235);
and U16700 (N_16700,N_15470,N_15729);
nor U16701 (N_16701,N_15955,N_15180);
xnor U16702 (N_16702,N_15550,N_15407);
xnor U16703 (N_16703,N_15759,N_15475);
nor U16704 (N_16704,N_15278,N_15726);
xnor U16705 (N_16705,N_15469,N_15712);
xor U16706 (N_16706,N_15322,N_15815);
and U16707 (N_16707,N_15210,N_15176);
and U16708 (N_16708,N_15455,N_15134);
xor U16709 (N_16709,N_15817,N_15341);
nand U16710 (N_16710,N_15442,N_15576);
nand U16711 (N_16711,N_15150,N_15294);
xnor U16712 (N_16712,N_15534,N_15265);
nand U16713 (N_16713,N_15564,N_15632);
nand U16714 (N_16714,N_15144,N_15329);
xor U16715 (N_16715,N_15175,N_15213);
or U16716 (N_16716,N_15055,N_15351);
or U16717 (N_16717,N_15226,N_15887);
nor U16718 (N_16718,N_15883,N_15108);
nand U16719 (N_16719,N_15310,N_15269);
and U16720 (N_16720,N_15164,N_15105);
xnor U16721 (N_16721,N_15733,N_15684);
and U16722 (N_16722,N_15067,N_15436);
xor U16723 (N_16723,N_15003,N_15626);
or U16724 (N_16724,N_15193,N_15836);
or U16725 (N_16725,N_15454,N_15631);
or U16726 (N_16726,N_15359,N_15367);
xnor U16727 (N_16727,N_15784,N_15467);
or U16728 (N_16728,N_15235,N_15890);
nand U16729 (N_16729,N_15689,N_15015);
nand U16730 (N_16730,N_15858,N_15540);
and U16731 (N_16731,N_15623,N_15650);
nor U16732 (N_16732,N_15412,N_15997);
xor U16733 (N_16733,N_15394,N_15862);
xnor U16734 (N_16734,N_15139,N_15800);
and U16735 (N_16735,N_15615,N_15135);
or U16736 (N_16736,N_15473,N_15498);
xor U16737 (N_16737,N_15271,N_15104);
or U16738 (N_16738,N_15636,N_15195);
nor U16739 (N_16739,N_15876,N_15085);
or U16740 (N_16740,N_15919,N_15844);
xor U16741 (N_16741,N_15407,N_15118);
nand U16742 (N_16742,N_15901,N_15357);
nand U16743 (N_16743,N_15579,N_15119);
nand U16744 (N_16744,N_15088,N_15724);
xnor U16745 (N_16745,N_15746,N_15722);
nand U16746 (N_16746,N_15555,N_15361);
xor U16747 (N_16747,N_15471,N_15273);
xor U16748 (N_16748,N_15883,N_15580);
xor U16749 (N_16749,N_15399,N_15675);
nor U16750 (N_16750,N_15543,N_15370);
or U16751 (N_16751,N_15609,N_15479);
or U16752 (N_16752,N_15591,N_15610);
nor U16753 (N_16753,N_15420,N_15820);
nor U16754 (N_16754,N_15031,N_15287);
and U16755 (N_16755,N_15564,N_15760);
or U16756 (N_16756,N_15953,N_15751);
or U16757 (N_16757,N_15017,N_15298);
and U16758 (N_16758,N_15214,N_15718);
and U16759 (N_16759,N_15123,N_15989);
and U16760 (N_16760,N_15971,N_15178);
nand U16761 (N_16761,N_15401,N_15904);
nor U16762 (N_16762,N_15078,N_15388);
xnor U16763 (N_16763,N_15570,N_15215);
and U16764 (N_16764,N_15454,N_15844);
nor U16765 (N_16765,N_15020,N_15655);
or U16766 (N_16766,N_15712,N_15693);
nor U16767 (N_16767,N_15369,N_15217);
nor U16768 (N_16768,N_15104,N_15423);
and U16769 (N_16769,N_15058,N_15059);
nor U16770 (N_16770,N_15023,N_15828);
nand U16771 (N_16771,N_15036,N_15292);
and U16772 (N_16772,N_15658,N_15789);
nor U16773 (N_16773,N_15229,N_15937);
nand U16774 (N_16774,N_15160,N_15231);
nor U16775 (N_16775,N_15773,N_15869);
nand U16776 (N_16776,N_15799,N_15578);
nand U16777 (N_16777,N_15372,N_15014);
nand U16778 (N_16778,N_15610,N_15987);
nor U16779 (N_16779,N_15412,N_15718);
nand U16780 (N_16780,N_15836,N_15977);
or U16781 (N_16781,N_15757,N_15118);
or U16782 (N_16782,N_15480,N_15066);
nand U16783 (N_16783,N_15093,N_15135);
nor U16784 (N_16784,N_15712,N_15061);
nor U16785 (N_16785,N_15501,N_15744);
or U16786 (N_16786,N_15645,N_15948);
and U16787 (N_16787,N_15484,N_15168);
or U16788 (N_16788,N_15849,N_15013);
nor U16789 (N_16789,N_15015,N_15473);
nand U16790 (N_16790,N_15443,N_15726);
and U16791 (N_16791,N_15349,N_15899);
or U16792 (N_16792,N_15797,N_15292);
xor U16793 (N_16793,N_15544,N_15482);
or U16794 (N_16794,N_15596,N_15866);
and U16795 (N_16795,N_15100,N_15136);
or U16796 (N_16796,N_15364,N_15838);
and U16797 (N_16797,N_15751,N_15163);
or U16798 (N_16798,N_15674,N_15514);
nor U16799 (N_16799,N_15341,N_15803);
xnor U16800 (N_16800,N_15515,N_15013);
or U16801 (N_16801,N_15191,N_15379);
nand U16802 (N_16802,N_15149,N_15677);
xnor U16803 (N_16803,N_15578,N_15446);
nand U16804 (N_16804,N_15496,N_15151);
xor U16805 (N_16805,N_15693,N_15467);
or U16806 (N_16806,N_15429,N_15670);
and U16807 (N_16807,N_15489,N_15469);
or U16808 (N_16808,N_15018,N_15167);
nor U16809 (N_16809,N_15145,N_15511);
nor U16810 (N_16810,N_15628,N_15182);
xnor U16811 (N_16811,N_15052,N_15572);
and U16812 (N_16812,N_15129,N_15882);
xnor U16813 (N_16813,N_15219,N_15798);
or U16814 (N_16814,N_15365,N_15340);
or U16815 (N_16815,N_15671,N_15467);
xor U16816 (N_16816,N_15780,N_15746);
and U16817 (N_16817,N_15850,N_15956);
or U16818 (N_16818,N_15615,N_15544);
or U16819 (N_16819,N_15090,N_15349);
and U16820 (N_16820,N_15950,N_15603);
nor U16821 (N_16821,N_15867,N_15669);
nor U16822 (N_16822,N_15586,N_15141);
xnor U16823 (N_16823,N_15242,N_15307);
and U16824 (N_16824,N_15838,N_15038);
and U16825 (N_16825,N_15829,N_15888);
nor U16826 (N_16826,N_15867,N_15923);
nand U16827 (N_16827,N_15872,N_15584);
and U16828 (N_16828,N_15108,N_15296);
or U16829 (N_16829,N_15495,N_15072);
xnor U16830 (N_16830,N_15552,N_15410);
xor U16831 (N_16831,N_15124,N_15292);
nor U16832 (N_16832,N_15050,N_15499);
nand U16833 (N_16833,N_15868,N_15418);
or U16834 (N_16834,N_15261,N_15981);
and U16835 (N_16835,N_15422,N_15118);
nor U16836 (N_16836,N_15112,N_15563);
and U16837 (N_16837,N_15701,N_15000);
or U16838 (N_16838,N_15766,N_15058);
nand U16839 (N_16839,N_15956,N_15792);
nor U16840 (N_16840,N_15753,N_15171);
xor U16841 (N_16841,N_15643,N_15793);
nand U16842 (N_16842,N_15735,N_15464);
nand U16843 (N_16843,N_15009,N_15218);
xnor U16844 (N_16844,N_15199,N_15149);
and U16845 (N_16845,N_15674,N_15633);
or U16846 (N_16846,N_15111,N_15408);
and U16847 (N_16847,N_15635,N_15349);
nor U16848 (N_16848,N_15313,N_15621);
xor U16849 (N_16849,N_15420,N_15919);
nand U16850 (N_16850,N_15149,N_15179);
and U16851 (N_16851,N_15205,N_15455);
and U16852 (N_16852,N_15195,N_15469);
nor U16853 (N_16853,N_15305,N_15723);
and U16854 (N_16854,N_15452,N_15228);
and U16855 (N_16855,N_15789,N_15836);
xor U16856 (N_16856,N_15716,N_15400);
nand U16857 (N_16857,N_15438,N_15506);
and U16858 (N_16858,N_15277,N_15644);
nor U16859 (N_16859,N_15269,N_15058);
nor U16860 (N_16860,N_15204,N_15844);
nor U16861 (N_16861,N_15805,N_15883);
nand U16862 (N_16862,N_15341,N_15409);
nand U16863 (N_16863,N_15279,N_15931);
nand U16864 (N_16864,N_15123,N_15356);
nand U16865 (N_16865,N_15763,N_15964);
nor U16866 (N_16866,N_15035,N_15953);
or U16867 (N_16867,N_15928,N_15148);
or U16868 (N_16868,N_15584,N_15484);
xnor U16869 (N_16869,N_15145,N_15128);
nor U16870 (N_16870,N_15659,N_15925);
nor U16871 (N_16871,N_15942,N_15255);
xor U16872 (N_16872,N_15809,N_15642);
and U16873 (N_16873,N_15339,N_15136);
nor U16874 (N_16874,N_15709,N_15760);
nor U16875 (N_16875,N_15429,N_15345);
or U16876 (N_16876,N_15575,N_15445);
or U16877 (N_16877,N_15468,N_15213);
and U16878 (N_16878,N_15301,N_15386);
nand U16879 (N_16879,N_15653,N_15757);
and U16880 (N_16880,N_15674,N_15000);
or U16881 (N_16881,N_15152,N_15613);
nand U16882 (N_16882,N_15355,N_15659);
nor U16883 (N_16883,N_15578,N_15967);
nand U16884 (N_16884,N_15554,N_15836);
nor U16885 (N_16885,N_15385,N_15354);
nand U16886 (N_16886,N_15078,N_15064);
xnor U16887 (N_16887,N_15472,N_15887);
nand U16888 (N_16888,N_15592,N_15860);
nand U16889 (N_16889,N_15460,N_15950);
nor U16890 (N_16890,N_15449,N_15453);
or U16891 (N_16891,N_15047,N_15153);
nand U16892 (N_16892,N_15372,N_15605);
xnor U16893 (N_16893,N_15269,N_15548);
nor U16894 (N_16894,N_15215,N_15722);
or U16895 (N_16895,N_15590,N_15719);
nor U16896 (N_16896,N_15606,N_15953);
nor U16897 (N_16897,N_15018,N_15094);
and U16898 (N_16898,N_15276,N_15392);
xnor U16899 (N_16899,N_15718,N_15293);
xnor U16900 (N_16900,N_15025,N_15713);
xnor U16901 (N_16901,N_15754,N_15353);
and U16902 (N_16902,N_15869,N_15475);
nand U16903 (N_16903,N_15491,N_15142);
or U16904 (N_16904,N_15971,N_15171);
nand U16905 (N_16905,N_15859,N_15012);
nand U16906 (N_16906,N_15145,N_15173);
xor U16907 (N_16907,N_15565,N_15762);
or U16908 (N_16908,N_15864,N_15739);
nand U16909 (N_16909,N_15852,N_15458);
nand U16910 (N_16910,N_15468,N_15036);
nand U16911 (N_16911,N_15125,N_15729);
or U16912 (N_16912,N_15678,N_15895);
or U16913 (N_16913,N_15515,N_15323);
and U16914 (N_16914,N_15369,N_15536);
or U16915 (N_16915,N_15446,N_15631);
nor U16916 (N_16916,N_15430,N_15782);
xor U16917 (N_16917,N_15475,N_15261);
and U16918 (N_16918,N_15271,N_15642);
xnor U16919 (N_16919,N_15089,N_15518);
nand U16920 (N_16920,N_15819,N_15737);
or U16921 (N_16921,N_15807,N_15197);
nand U16922 (N_16922,N_15585,N_15324);
or U16923 (N_16923,N_15213,N_15198);
xor U16924 (N_16924,N_15581,N_15421);
nand U16925 (N_16925,N_15966,N_15084);
or U16926 (N_16926,N_15751,N_15742);
nor U16927 (N_16927,N_15562,N_15640);
xor U16928 (N_16928,N_15934,N_15100);
nand U16929 (N_16929,N_15670,N_15656);
or U16930 (N_16930,N_15069,N_15315);
or U16931 (N_16931,N_15768,N_15882);
nor U16932 (N_16932,N_15176,N_15328);
and U16933 (N_16933,N_15575,N_15292);
or U16934 (N_16934,N_15878,N_15412);
xnor U16935 (N_16935,N_15001,N_15304);
nand U16936 (N_16936,N_15712,N_15463);
nand U16937 (N_16937,N_15274,N_15021);
and U16938 (N_16938,N_15320,N_15849);
and U16939 (N_16939,N_15930,N_15621);
xnor U16940 (N_16940,N_15552,N_15833);
nor U16941 (N_16941,N_15571,N_15390);
nand U16942 (N_16942,N_15722,N_15739);
xnor U16943 (N_16943,N_15102,N_15574);
or U16944 (N_16944,N_15961,N_15152);
nand U16945 (N_16945,N_15931,N_15629);
xnor U16946 (N_16946,N_15962,N_15033);
nand U16947 (N_16947,N_15525,N_15469);
xnor U16948 (N_16948,N_15529,N_15366);
nand U16949 (N_16949,N_15891,N_15422);
nand U16950 (N_16950,N_15859,N_15400);
nor U16951 (N_16951,N_15679,N_15742);
and U16952 (N_16952,N_15639,N_15833);
and U16953 (N_16953,N_15931,N_15226);
or U16954 (N_16954,N_15135,N_15767);
nand U16955 (N_16955,N_15295,N_15873);
xor U16956 (N_16956,N_15190,N_15501);
and U16957 (N_16957,N_15054,N_15996);
xnor U16958 (N_16958,N_15904,N_15825);
and U16959 (N_16959,N_15808,N_15886);
nor U16960 (N_16960,N_15403,N_15384);
xnor U16961 (N_16961,N_15702,N_15074);
nand U16962 (N_16962,N_15117,N_15935);
and U16963 (N_16963,N_15195,N_15684);
nand U16964 (N_16964,N_15683,N_15567);
nor U16965 (N_16965,N_15585,N_15756);
nor U16966 (N_16966,N_15420,N_15027);
and U16967 (N_16967,N_15551,N_15217);
nand U16968 (N_16968,N_15647,N_15444);
or U16969 (N_16969,N_15207,N_15677);
and U16970 (N_16970,N_15296,N_15822);
and U16971 (N_16971,N_15113,N_15374);
xor U16972 (N_16972,N_15985,N_15905);
and U16973 (N_16973,N_15345,N_15237);
nor U16974 (N_16974,N_15119,N_15732);
nand U16975 (N_16975,N_15459,N_15546);
nor U16976 (N_16976,N_15529,N_15454);
or U16977 (N_16977,N_15763,N_15519);
nand U16978 (N_16978,N_15022,N_15188);
xnor U16979 (N_16979,N_15658,N_15707);
nor U16980 (N_16980,N_15981,N_15580);
nand U16981 (N_16981,N_15315,N_15286);
xnor U16982 (N_16982,N_15242,N_15176);
nand U16983 (N_16983,N_15838,N_15777);
xnor U16984 (N_16984,N_15949,N_15029);
xor U16985 (N_16985,N_15298,N_15857);
or U16986 (N_16986,N_15445,N_15374);
nor U16987 (N_16987,N_15355,N_15750);
nor U16988 (N_16988,N_15691,N_15624);
nor U16989 (N_16989,N_15538,N_15793);
nor U16990 (N_16990,N_15914,N_15149);
or U16991 (N_16991,N_15725,N_15767);
nand U16992 (N_16992,N_15493,N_15921);
xor U16993 (N_16993,N_15808,N_15138);
nand U16994 (N_16994,N_15443,N_15299);
nand U16995 (N_16995,N_15458,N_15565);
nor U16996 (N_16996,N_15081,N_15685);
nand U16997 (N_16997,N_15391,N_15925);
nand U16998 (N_16998,N_15372,N_15924);
nor U16999 (N_16999,N_15832,N_15097);
nor U17000 (N_17000,N_16408,N_16134);
nand U17001 (N_17001,N_16426,N_16621);
nand U17002 (N_17002,N_16595,N_16752);
nand U17003 (N_17003,N_16350,N_16416);
or U17004 (N_17004,N_16329,N_16533);
nor U17005 (N_17005,N_16894,N_16254);
xor U17006 (N_17006,N_16530,N_16542);
xor U17007 (N_17007,N_16368,N_16093);
and U17008 (N_17008,N_16005,N_16458);
and U17009 (N_17009,N_16417,N_16104);
nand U17010 (N_17010,N_16502,N_16317);
or U17011 (N_17011,N_16414,N_16880);
or U17012 (N_17012,N_16614,N_16852);
nor U17013 (N_17013,N_16187,N_16831);
xnor U17014 (N_17014,N_16810,N_16069);
nand U17015 (N_17015,N_16722,N_16899);
or U17016 (N_17016,N_16782,N_16150);
nand U17017 (N_17017,N_16320,N_16668);
xnor U17018 (N_17018,N_16029,N_16656);
xor U17019 (N_17019,N_16133,N_16686);
or U17020 (N_17020,N_16296,N_16212);
or U17021 (N_17021,N_16519,N_16356);
or U17022 (N_17022,N_16698,N_16049);
or U17023 (N_17023,N_16809,N_16255);
or U17024 (N_17024,N_16751,N_16805);
xor U17025 (N_17025,N_16312,N_16390);
xnor U17026 (N_17026,N_16919,N_16216);
xor U17027 (N_17027,N_16207,N_16159);
xor U17028 (N_17028,N_16986,N_16323);
nand U17029 (N_17029,N_16827,N_16083);
nand U17030 (N_17030,N_16836,N_16790);
and U17031 (N_17031,N_16404,N_16982);
xnor U17032 (N_17032,N_16513,N_16674);
xnor U17033 (N_17033,N_16916,N_16096);
or U17034 (N_17034,N_16591,N_16094);
nand U17035 (N_17035,N_16436,N_16248);
and U17036 (N_17036,N_16870,N_16945);
nor U17037 (N_17037,N_16279,N_16106);
or U17038 (N_17038,N_16362,N_16817);
and U17039 (N_17039,N_16003,N_16540);
xor U17040 (N_17040,N_16048,N_16963);
or U17041 (N_17041,N_16126,N_16812);
or U17042 (N_17042,N_16731,N_16160);
and U17043 (N_17043,N_16153,N_16068);
and U17044 (N_17044,N_16703,N_16626);
xnor U17045 (N_17045,N_16051,N_16943);
nand U17046 (N_17046,N_16879,N_16842);
and U17047 (N_17047,N_16816,N_16795);
or U17048 (N_17048,N_16167,N_16475);
or U17049 (N_17049,N_16220,N_16324);
and U17050 (N_17050,N_16901,N_16933);
or U17051 (N_17051,N_16654,N_16398);
or U17052 (N_17052,N_16715,N_16344);
and U17053 (N_17053,N_16907,N_16141);
and U17054 (N_17054,N_16859,N_16478);
nand U17055 (N_17055,N_16256,N_16459);
and U17056 (N_17056,N_16864,N_16774);
nor U17057 (N_17057,N_16673,N_16823);
and U17058 (N_17058,N_16689,N_16284);
or U17059 (N_17059,N_16536,N_16738);
nor U17060 (N_17060,N_16578,N_16095);
or U17061 (N_17061,N_16662,N_16843);
or U17062 (N_17062,N_16549,N_16575);
nand U17063 (N_17063,N_16528,N_16599);
and U17064 (N_17064,N_16709,N_16780);
nand U17065 (N_17065,N_16596,N_16940);
or U17066 (N_17066,N_16690,N_16209);
nand U17067 (N_17067,N_16788,N_16609);
and U17068 (N_17068,N_16440,N_16033);
xnor U17069 (N_17069,N_16031,N_16957);
nand U17070 (N_17070,N_16219,N_16878);
and U17071 (N_17071,N_16607,N_16018);
nand U17072 (N_17072,N_16201,N_16156);
xnor U17073 (N_17073,N_16177,N_16973);
and U17074 (N_17074,N_16235,N_16341);
nand U17075 (N_17075,N_16808,N_16789);
xnor U17076 (N_17076,N_16064,N_16286);
or U17077 (N_17077,N_16411,N_16950);
xnor U17078 (N_17078,N_16625,N_16022);
xnor U17079 (N_17079,N_16965,N_16084);
xor U17080 (N_17080,N_16331,N_16639);
nor U17081 (N_17081,N_16643,N_16054);
and U17082 (N_17082,N_16088,N_16939);
nand U17083 (N_17083,N_16234,N_16432);
nor U17084 (N_17084,N_16562,N_16259);
or U17085 (N_17085,N_16613,N_16466);
nor U17086 (N_17086,N_16551,N_16192);
or U17087 (N_17087,N_16053,N_16984);
nand U17088 (N_17088,N_16659,N_16797);
nand U17089 (N_17089,N_16733,N_16061);
nand U17090 (N_17090,N_16764,N_16838);
nand U17091 (N_17091,N_16685,N_16748);
and U17092 (N_17092,N_16392,N_16166);
xnor U17093 (N_17093,N_16503,N_16706);
and U17094 (N_17094,N_16820,N_16474);
and U17095 (N_17095,N_16188,N_16360);
xor U17096 (N_17096,N_16861,N_16687);
and U17097 (N_17097,N_16981,N_16741);
xnor U17098 (N_17098,N_16730,N_16330);
nand U17099 (N_17099,N_16516,N_16967);
nand U17100 (N_17100,N_16071,N_16070);
nand U17101 (N_17101,N_16336,N_16321);
and U17102 (N_17102,N_16688,N_16953);
xor U17103 (N_17103,N_16976,N_16267);
xor U17104 (N_17104,N_16787,N_16338);
or U17105 (N_17105,N_16905,N_16322);
and U17106 (N_17106,N_16245,N_16202);
nor U17107 (N_17107,N_16162,N_16406);
nand U17108 (N_17108,N_16926,N_16629);
or U17109 (N_17109,N_16117,N_16553);
nor U17110 (N_17110,N_16152,N_16196);
nor U17111 (N_17111,N_16052,N_16854);
nand U17112 (N_17112,N_16538,N_16379);
or U17113 (N_17113,N_16098,N_16678);
nand U17114 (N_17114,N_16446,N_16657);
nand U17115 (N_17115,N_16962,N_16924);
nand U17116 (N_17116,N_16251,N_16441);
xnor U17117 (N_17117,N_16734,N_16264);
xnor U17118 (N_17118,N_16079,N_16750);
nor U17119 (N_17119,N_16566,N_16754);
or U17120 (N_17120,N_16995,N_16695);
xor U17121 (N_17121,N_16228,N_16343);
nand U17122 (N_17122,N_16129,N_16349);
and U17123 (N_17123,N_16281,N_16144);
nor U17124 (N_17124,N_16556,N_16498);
nand U17125 (N_17125,N_16840,N_16959);
or U17126 (N_17126,N_16651,N_16884);
xnor U17127 (N_17127,N_16250,N_16479);
xor U17128 (N_17128,N_16922,N_16559);
xnor U17129 (N_17129,N_16139,N_16989);
xnor U17130 (N_17130,N_16047,N_16807);
or U17131 (N_17131,N_16289,N_16565);
and U17132 (N_17132,N_16482,N_16552);
and U17133 (N_17133,N_16198,N_16600);
and U17134 (N_17134,N_16020,N_16765);
nor U17135 (N_17135,N_16298,N_16822);
and U17136 (N_17136,N_16315,N_16158);
nor U17137 (N_17137,N_16929,N_16988);
nor U17138 (N_17138,N_16524,N_16771);
nand U17139 (N_17139,N_16340,N_16646);
and U17140 (N_17140,N_16914,N_16077);
nor U17141 (N_17141,N_16438,N_16714);
or U17142 (N_17142,N_16745,N_16637);
and U17143 (N_17143,N_16735,N_16399);
nor U17144 (N_17144,N_16520,N_16707);
nand U17145 (N_17145,N_16550,N_16142);
and U17146 (N_17146,N_16430,N_16337);
nand U17147 (N_17147,N_16027,N_16736);
nand U17148 (N_17148,N_16623,N_16361);
nand U17149 (N_17149,N_16218,N_16935);
or U17150 (N_17150,N_16044,N_16677);
nor U17151 (N_17151,N_16580,N_16278);
nor U17152 (N_17152,N_16236,N_16389);
nand U17153 (N_17153,N_16036,N_16371);
and U17154 (N_17154,N_16303,N_16608);
nand U17155 (N_17155,N_16647,N_16514);
xnor U17156 (N_17156,N_16941,N_16194);
nand U17157 (N_17157,N_16305,N_16062);
nor U17158 (N_17158,N_16847,N_16848);
and U17159 (N_17159,N_16424,N_16767);
nor U17160 (N_17160,N_16669,N_16785);
nor U17161 (N_17161,N_16841,N_16906);
xnor U17162 (N_17162,N_16171,N_16993);
xnor U17163 (N_17163,N_16143,N_16979);
nand U17164 (N_17164,N_16463,N_16509);
nand U17165 (N_17165,N_16992,N_16369);
and U17166 (N_17166,N_16944,N_16593);
nor U17167 (N_17167,N_16001,N_16856);
nand U17168 (N_17168,N_16043,N_16419);
or U17169 (N_17169,N_16515,N_16108);
or U17170 (N_17170,N_16778,N_16292);
or U17171 (N_17171,N_16727,N_16616);
or U17172 (N_17172,N_16958,N_16874);
or U17173 (N_17173,N_16523,N_16586);
nor U17174 (N_17174,N_16470,N_16759);
xor U17175 (N_17175,N_16109,N_16747);
nand U17176 (N_17176,N_16386,N_16415);
or U17177 (N_17177,N_16762,N_16719);
xnor U17178 (N_17178,N_16472,N_16570);
and U17179 (N_17179,N_16425,N_16006);
xor U17180 (N_17180,N_16431,N_16505);
and U17181 (N_17181,N_16299,N_16381);
and U17182 (N_17182,N_16952,N_16755);
xor U17183 (N_17183,N_16487,N_16757);
nand U17184 (N_17184,N_16547,N_16115);
nor U17185 (N_17185,N_16412,N_16974);
xor U17186 (N_17186,N_16518,N_16866);
or U17187 (N_17187,N_16040,N_16008);
xor U17188 (N_17188,N_16729,N_16232);
and U17189 (N_17189,N_16155,N_16364);
and U17190 (N_17190,N_16781,N_16056);
xor U17191 (N_17191,N_16573,N_16893);
nand U17192 (N_17192,N_16353,N_16978);
or U17193 (N_17193,N_16396,N_16455);
nand U17194 (N_17194,N_16630,N_16877);
or U17195 (N_17195,N_16873,N_16173);
xnor U17196 (N_17196,N_16063,N_16704);
xor U17197 (N_17197,N_16060,N_16791);
and U17198 (N_17198,N_16650,N_16758);
nand U17199 (N_17199,N_16969,N_16110);
xor U17200 (N_17200,N_16041,N_16004);
or U17201 (N_17201,N_16560,N_16494);
nor U17202 (N_17202,N_16761,N_16670);
and U17203 (N_17203,N_16169,N_16086);
and U17204 (N_17204,N_16229,N_16694);
nor U17205 (N_17205,N_16377,N_16249);
xnor U17206 (N_17206,N_16964,N_16042);
or U17207 (N_17207,N_16628,N_16132);
xor U17208 (N_17208,N_16577,N_16226);
nor U17209 (N_17209,N_16871,N_16602);
nor U17210 (N_17210,N_16858,N_16671);
nor U17211 (N_17211,N_16339,N_16495);
nor U17212 (N_17212,N_16499,N_16594);
nor U17213 (N_17213,N_16572,N_16102);
and U17214 (N_17214,N_16853,N_16632);
or U17215 (N_17215,N_16168,N_16749);
nand U17216 (N_17216,N_16358,N_16700);
and U17217 (N_17217,N_16311,N_16009);
xnor U17218 (N_17218,N_16534,N_16994);
or U17219 (N_17219,N_16857,N_16295);
xor U17220 (N_17220,N_16306,N_16302);
nand U17221 (N_17221,N_16434,N_16942);
nor U17222 (N_17222,N_16996,N_16876);
or U17223 (N_17223,N_16113,N_16111);
nor U17224 (N_17224,N_16784,N_16909);
nor U17225 (N_17225,N_16354,N_16511);
and U17226 (N_17226,N_16180,N_16763);
and U17227 (N_17227,N_16429,N_16468);
nor U17228 (N_17228,N_16347,N_16091);
and U17229 (N_17229,N_16409,N_16664);
or U17230 (N_17230,N_16118,N_16696);
nand U17231 (N_17231,N_16391,N_16997);
or U17232 (N_17232,N_16266,N_16260);
nand U17233 (N_17233,N_16057,N_16319);
and U17234 (N_17234,N_16138,N_16839);
or U17235 (N_17235,N_16903,N_16103);
and U17236 (N_17236,N_16442,N_16604);
xor U17237 (N_17237,N_16471,N_16526);
nand U17238 (N_17238,N_16697,N_16225);
xor U17239 (N_17239,N_16372,N_16980);
or U17240 (N_17240,N_16521,N_16172);
nor U17241 (N_17241,N_16313,N_16786);
nor U17242 (N_17242,N_16913,N_16620);
and U17243 (N_17243,N_16375,N_16985);
and U17244 (N_17244,N_16019,N_16039);
xor U17245 (N_17245,N_16793,N_16011);
xor U17246 (N_17246,N_16619,N_16087);
nor U17247 (N_17247,N_16010,N_16247);
and U17248 (N_17248,N_16875,N_16224);
and U17249 (N_17249,N_16612,N_16746);
or U17250 (N_17250,N_16148,N_16720);
nand U17251 (N_17251,N_16378,N_16075);
nor U17252 (N_17252,N_16676,N_16314);
xor U17253 (N_17253,N_16204,N_16448);
xnor U17254 (N_17254,N_16667,N_16923);
or U17255 (N_17255,N_16796,N_16211);
xor U17256 (N_17256,N_16701,N_16915);
xnor U17257 (N_17257,N_16675,N_16119);
and U17258 (N_17258,N_16862,N_16955);
or U17259 (N_17259,N_16035,N_16889);
and U17260 (N_17260,N_16946,N_16558);
and U17261 (N_17261,N_16447,N_16800);
xnor U17262 (N_17262,N_16373,N_16548);
xnor U17263 (N_17263,N_16633,N_16897);
nor U17264 (N_17264,N_16484,N_16554);
or U17265 (N_17265,N_16367,N_16199);
nand U17266 (N_17266,N_16936,N_16265);
xnor U17267 (N_17267,N_16030,N_16253);
or U17268 (N_17268,N_16618,N_16691);
and U17269 (N_17269,N_16660,N_16151);
nand U17270 (N_17270,N_16401,N_16145);
nor U17271 (N_17271,N_16376,N_16481);
xor U17272 (N_17272,N_16522,N_16644);
nor U17273 (N_17273,N_16355,N_16116);
or U17274 (N_17274,N_16131,N_16325);
and U17275 (N_17275,N_16309,N_16833);
nor U17276 (N_17276,N_16579,N_16128);
and U17277 (N_17277,N_16122,N_16301);
nor U17278 (N_17278,N_16863,N_16597);
xor U17279 (N_17279,N_16058,N_16017);
nor U17280 (N_17280,N_16016,N_16428);
nand U17281 (N_17281,N_16539,N_16592);
and U17282 (N_17282,N_16770,N_16140);
and U17283 (N_17283,N_16589,N_16737);
or U17284 (N_17284,N_16335,N_16038);
nand U17285 (N_17285,N_16357,N_16467);
and U17286 (N_17286,N_16825,N_16496);
nor U17287 (N_17287,N_16918,N_16175);
and U17288 (N_17288,N_16273,N_16405);
xnor U17289 (N_17289,N_16887,N_16803);
nand U17290 (N_17290,N_16772,N_16811);
xnor U17291 (N_17291,N_16189,N_16683);
nor U17292 (N_17292,N_16636,N_16990);
or U17293 (N_17293,N_16705,N_16328);
and U17294 (N_17294,N_16123,N_16046);
xor U17295 (N_17295,N_16948,N_16756);
nor U17296 (N_17296,N_16653,N_16182);
and U17297 (N_17297,N_16215,N_16252);
nand U17298 (N_17298,N_16258,N_16025);
nor U17299 (N_17299,N_16032,N_16137);
nor U17300 (N_17300,N_16684,N_16851);
or U17301 (N_17301,N_16222,N_16835);
nand U17302 (N_17302,N_16708,N_16214);
or U17303 (N_17303,N_16457,N_16423);
or U17304 (N_17304,N_16290,N_16233);
or U17305 (N_17305,N_16947,N_16231);
and U17306 (N_17306,N_16930,N_16034);
nand U17307 (N_17307,N_16888,N_16699);
xor U17308 (N_17308,N_16476,N_16184);
xnor U17309 (N_17309,N_16531,N_16555);
nor U17310 (N_17310,N_16462,N_16804);
and U17311 (N_17311,N_16149,N_16200);
nor U17312 (N_17312,N_16393,N_16240);
xnor U17313 (N_17313,N_16512,N_16217);
and U17314 (N_17314,N_16268,N_16297);
and U17315 (N_17315,N_16724,N_16937);
nor U17316 (N_17316,N_16348,N_16504);
nor U17317 (N_17317,N_16775,N_16532);
or U17318 (N_17318,N_16917,N_16576);
and U17319 (N_17319,N_16427,N_16185);
xor U17320 (N_17320,N_16161,N_16453);
nor U17321 (N_17321,N_16635,N_16726);
xor U17322 (N_17322,N_16477,N_16000);
or U17323 (N_17323,N_16725,N_16269);
nand U17324 (N_17324,N_16584,N_16450);
and U17325 (N_17325,N_16304,N_16363);
nand U17326 (N_17326,N_16885,N_16120);
and U17327 (N_17327,N_16065,N_16525);
xor U17328 (N_17328,N_16157,N_16089);
nand U17329 (N_17329,N_16537,N_16318);
nand U17330 (N_17330,N_16452,N_16966);
nor U17331 (N_17331,N_16464,N_16867);
and U17332 (N_17332,N_16615,N_16783);
nand U17333 (N_17333,N_16818,N_16587);
xnor U17334 (N_17334,N_16488,N_16383);
and U17335 (N_17335,N_16227,N_16485);
nand U17336 (N_17336,N_16850,N_16213);
or U17337 (N_17337,N_16346,N_16983);
nor U17338 (N_17338,N_16802,N_16543);
nand U17339 (N_17339,N_16768,N_16545);
nand U17340 (N_17340,N_16385,N_16977);
nand U17341 (N_17341,N_16824,N_16890);
nor U17342 (N_17342,N_16622,N_16590);
or U17343 (N_17343,N_16037,N_16649);
nor U17344 (N_17344,N_16045,N_16640);
nor U17345 (N_17345,N_16583,N_16257);
or U17346 (N_17346,N_16895,N_16420);
nand U17347 (N_17347,N_16483,N_16846);
xnor U17348 (N_17348,N_16099,N_16230);
and U17349 (N_17349,N_16563,N_16603);
nand U17350 (N_17350,N_16300,N_16869);
xnor U17351 (N_17351,N_16456,N_16601);
nor U17352 (N_17352,N_16739,N_16261);
or U17353 (N_17353,N_16239,N_16308);
xnor U17354 (N_17354,N_16627,N_16191);
and U17355 (N_17355,N_16911,N_16624);
nor U17356 (N_17356,N_16611,N_16881);
xnor U17357 (N_17357,N_16275,N_16655);
xnor U17358 (N_17358,N_16742,N_16794);
xnor U17359 (N_17359,N_16740,N_16291);
and U17360 (N_17360,N_16892,N_16316);
xnor U17361 (N_17361,N_16588,N_16801);
nand U17362 (N_17362,N_16345,N_16912);
xnor U17363 (N_17363,N_16101,N_16510);
and U17364 (N_17364,N_16972,N_16910);
nand U17365 (N_17365,N_16693,N_16574);
nand U17366 (N_17366,N_16055,N_16666);
nand U17367 (N_17367,N_16407,N_16598);
or U17368 (N_17368,N_16178,N_16799);
xnor U17369 (N_17369,N_16205,N_16387);
nor U17370 (N_17370,N_16766,N_16883);
nor U17371 (N_17371,N_16285,N_16294);
xnor U17372 (N_17372,N_16561,N_16002);
or U17373 (N_17373,N_16288,N_16527);
nand U17374 (N_17374,N_16114,N_16710);
or U17375 (N_17375,N_16154,N_16821);
nand U17376 (N_17376,N_16568,N_16105);
or U17377 (N_17377,N_16951,N_16949);
and U17378 (N_17378,N_16183,N_16961);
nor U17379 (N_17379,N_16480,N_16461);
nor U17380 (N_17380,N_16310,N_16569);
or U17381 (N_17381,N_16606,N_16059);
nor U17382 (N_17382,N_16680,N_16195);
or U17383 (N_17383,N_16112,N_16679);
or U17384 (N_17384,N_16439,N_16242);
or U17385 (N_17385,N_16370,N_16388);
nand U17386 (N_17386,N_16855,N_16418);
or U17387 (N_17387,N_16433,N_16638);
xor U17388 (N_17388,N_16203,N_16384);
nand U17389 (N_17389,N_16342,N_16050);
nand U17390 (N_17390,N_16090,N_16223);
xor U17391 (N_17391,N_16270,N_16882);
or U17392 (N_17392,N_16723,N_16014);
nand U17393 (N_17393,N_16716,N_16073);
or U17394 (N_17394,N_16074,N_16243);
and U17395 (N_17395,N_16970,N_16938);
and U17396 (N_17396,N_16645,N_16652);
or U17397 (N_17397,N_16272,N_16382);
and U17398 (N_17398,N_16641,N_16712);
xor U17399 (N_17399,N_16374,N_16081);
or U17400 (N_17400,N_16921,N_16642);
xnor U17401 (N_17401,N_16130,N_16956);
xor U17402 (N_17402,N_16682,N_16845);
nor U17403 (N_17403,N_16136,N_16146);
or U17404 (N_17404,N_16263,N_16413);
or U17405 (N_17405,N_16927,N_16648);
or U17406 (N_17406,N_16332,N_16546);
xnor U17407 (N_17407,N_16658,N_16280);
xor U17408 (N_17408,N_16798,N_16181);
and U17409 (N_17409,N_16681,N_16403);
nor U17410 (N_17410,N_16813,N_16422);
and U17411 (N_17411,N_16928,N_16410);
nand U17412 (N_17412,N_16998,N_16991);
and U17413 (N_17413,N_16400,N_16449);
nor U17414 (N_17414,N_16080,N_16366);
nor U17415 (N_17415,N_16097,N_16672);
nor U17416 (N_17416,N_16276,N_16815);
nand U17417 (N_17417,N_16072,N_16830);
nand U17418 (N_17418,N_16634,N_16334);
or U17419 (N_17419,N_16777,N_16773);
and U17420 (N_17420,N_16023,N_16732);
or U17421 (N_17421,N_16564,N_16454);
nand U17422 (N_17422,N_16663,N_16241);
nand U17423 (N_17423,N_16617,N_16501);
or U17424 (N_17424,N_16489,N_16127);
xor U17425 (N_17425,N_16121,N_16896);
and U17426 (N_17426,N_16902,N_16015);
nor U17427 (N_17427,N_16849,N_16506);
xor U17428 (N_17428,N_16007,N_16713);
or U17429 (N_17429,N_16164,N_16262);
nor U17430 (N_17430,N_16326,N_16728);
nand U17431 (N_17431,N_16100,N_16206);
xnor U17432 (N_17432,N_16834,N_16176);
xnor U17433 (N_17433,N_16541,N_16197);
nor U17434 (N_17434,N_16743,N_16582);
nor U17435 (N_17435,N_16567,N_16999);
and U17436 (N_17436,N_16500,N_16237);
xnor U17437 (N_17437,N_16210,N_16987);
nor U17438 (N_17438,N_16492,N_16507);
xnor U17439 (N_17439,N_16085,N_16491);
nor U17440 (N_17440,N_16860,N_16497);
xnor U17441 (N_17441,N_16365,N_16920);
or U17442 (N_17442,N_16179,N_16898);
xor U17443 (N_17443,N_16282,N_16380);
nor U17444 (N_17444,N_16900,N_16473);
nand U17445 (N_17445,N_16975,N_16779);
xnor U17446 (N_17446,N_16493,N_16021);
and U17447 (N_17447,N_16960,N_16610);
xnor U17448 (N_17448,N_16327,N_16544);
nand U17449 (N_17449,N_16868,N_16283);
xnor U17450 (N_17450,N_16165,N_16891);
and U17451 (N_17451,N_16147,N_16517);
nor U17452 (N_17452,N_16934,N_16221);
xor U17453 (N_17453,N_16529,N_16753);
xnor U17454 (N_17454,N_16066,N_16394);
and U17455 (N_17455,N_16333,N_16828);
xor U17456 (N_17456,N_16744,N_16557);
nor U17457 (N_17457,N_16435,N_16012);
or U17458 (N_17458,N_16397,N_16421);
or U17459 (N_17459,N_16631,N_16271);
nand U17460 (N_17460,N_16135,N_16508);
and U17461 (N_17461,N_16490,N_16925);
nor U17462 (N_17462,N_16486,N_16076);
xor U17463 (N_17463,N_16274,N_16776);
or U17464 (N_17464,N_16125,N_16829);
xnor U17465 (N_17465,N_16444,N_16163);
nor U17466 (N_17466,N_16954,N_16814);
and U17467 (N_17467,N_16904,N_16402);
nor U17468 (N_17468,N_16124,N_16826);
and U17469 (N_17469,N_16186,N_16351);
nand U17470 (N_17470,N_16193,N_16692);
nor U17471 (N_17471,N_16605,N_16718);
and U17472 (N_17472,N_16806,N_16661);
and U17473 (N_17473,N_16535,N_16819);
xor U17474 (N_17474,N_16711,N_16792);
nor U17475 (N_17475,N_16443,N_16769);
or U17476 (N_17476,N_16665,N_16352);
nor U17477 (N_17477,N_16865,N_16067);
and U17478 (N_17478,N_16092,N_16013);
nor U17479 (N_17479,N_16445,N_16844);
nand U17480 (N_17480,N_16469,N_16174);
or U17481 (N_17481,N_16832,N_16208);
nand U17482 (N_17482,N_16721,N_16170);
nor U17483 (N_17483,N_16293,N_16024);
or U17484 (N_17484,N_16760,N_16082);
nor U17485 (N_17485,N_16437,N_16244);
nor U17486 (N_17486,N_16465,N_16190);
and U17487 (N_17487,N_16968,N_16837);
nand U17488 (N_17488,N_16872,N_16238);
nor U17489 (N_17489,N_16971,N_16026);
nor U17490 (N_17490,N_16078,N_16460);
and U17491 (N_17491,N_16451,N_16307);
nand U17492 (N_17492,N_16287,N_16908);
or U17493 (N_17493,N_16246,N_16581);
nor U17494 (N_17494,N_16702,N_16028);
nor U17495 (N_17495,N_16277,N_16571);
xor U17496 (N_17496,N_16931,N_16886);
xnor U17497 (N_17497,N_16932,N_16717);
and U17498 (N_17498,N_16585,N_16359);
xor U17499 (N_17499,N_16395,N_16107);
and U17500 (N_17500,N_16515,N_16755);
or U17501 (N_17501,N_16048,N_16975);
or U17502 (N_17502,N_16713,N_16515);
xnor U17503 (N_17503,N_16932,N_16014);
or U17504 (N_17504,N_16269,N_16157);
or U17505 (N_17505,N_16612,N_16957);
nand U17506 (N_17506,N_16959,N_16360);
or U17507 (N_17507,N_16130,N_16330);
and U17508 (N_17508,N_16417,N_16608);
and U17509 (N_17509,N_16858,N_16252);
nor U17510 (N_17510,N_16910,N_16633);
nor U17511 (N_17511,N_16691,N_16179);
and U17512 (N_17512,N_16754,N_16953);
nor U17513 (N_17513,N_16628,N_16714);
and U17514 (N_17514,N_16793,N_16482);
xnor U17515 (N_17515,N_16295,N_16860);
xor U17516 (N_17516,N_16368,N_16687);
or U17517 (N_17517,N_16546,N_16950);
or U17518 (N_17518,N_16172,N_16176);
nor U17519 (N_17519,N_16068,N_16892);
nand U17520 (N_17520,N_16867,N_16362);
nand U17521 (N_17521,N_16175,N_16260);
nand U17522 (N_17522,N_16544,N_16537);
or U17523 (N_17523,N_16731,N_16600);
xnor U17524 (N_17524,N_16396,N_16907);
nand U17525 (N_17525,N_16087,N_16981);
and U17526 (N_17526,N_16103,N_16406);
or U17527 (N_17527,N_16697,N_16860);
nor U17528 (N_17528,N_16364,N_16183);
nand U17529 (N_17529,N_16275,N_16378);
or U17530 (N_17530,N_16435,N_16033);
nor U17531 (N_17531,N_16720,N_16102);
xnor U17532 (N_17532,N_16283,N_16081);
and U17533 (N_17533,N_16929,N_16585);
nand U17534 (N_17534,N_16547,N_16978);
nor U17535 (N_17535,N_16437,N_16436);
or U17536 (N_17536,N_16927,N_16463);
nor U17537 (N_17537,N_16808,N_16550);
nor U17538 (N_17538,N_16235,N_16038);
or U17539 (N_17539,N_16668,N_16428);
or U17540 (N_17540,N_16471,N_16477);
xor U17541 (N_17541,N_16383,N_16011);
nor U17542 (N_17542,N_16263,N_16041);
nor U17543 (N_17543,N_16592,N_16497);
nand U17544 (N_17544,N_16511,N_16198);
or U17545 (N_17545,N_16767,N_16852);
nor U17546 (N_17546,N_16140,N_16214);
nand U17547 (N_17547,N_16693,N_16823);
xnor U17548 (N_17548,N_16268,N_16910);
and U17549 (N_17549,N_16488,N_16904);
and U17550 (N_17550,N_16998,N_16988);
and U17551 (N_17551,N_16485,N_16595);
xor U17552 (N_17552,N_16655,N_16704);
or U17553 (N_17553,N_16383,N_16028);
nor U17554 (N_17554,N_16631,N_16811);
xor U17555 (N_17555,N_16171,N_16652);
xor U17556 (N_17556,N_16137,N_16115);
nand U17557 (N_17557,N_16315,N_16282);
or U17558 (N_17558,N_16411,N_16772);
or U17559 (N_17559,N_16852,N_16178);
nand U17560 (N_17560,N_16156,N_16396);
nor U17561 (N_17561,N_16559,N_16729);
nand U17562 (N_17562,N_16653,N_16342);
and U17563 (N_17563,N_16642,N_16790);
nor U17564 (N_17564,N_16806,N_16452);
and U17565 (N_17565,N_16929,N_16679);
or U17566 (N_17566,N_16651,N_16904);
nor U17567 (N_17567,N_16290,N_16449);
xnor U17568 (N_17568,N_16475,N_16329);
or U17569 (N_17569,N_16070,N_16858);
nor U17570 (N_17570,N_16580,N_16665);
xnor U17571 (N_17571,N_16477,N_16652);
and U17572 (N_17572,N_16199,N_16427);
nor U17573 (N_17573,N_16341,N_16423);
nand U17574 (N_17574,N_16450,N_16375);
nor U17575 (N_17575,N_16596,N_16800);
or U17576 (N_17576,N_16162,N_16703);
xnor U17577 (N_17577,N_16940,N_16007);
xor U17578 (N_17578,N_16859,N_16198);
nand U17579 (N_17579,N_16728,N_16210);
nor U17580 (N_17580,N_16847,N_16075);
nand U17581 (N_17581,N_16018,N_16977);
xor U17582 (N_17582,N_16798,N_16397);
or U17583 (N_17583,N_16296,N_16091);
nand U17584 (N_17584,N_16945,N_16246);
xor U17585 (N_17585,N_16628,N_16266);
nand U17586 (N_17586,N_16950,N_16604);
nand U17587 (N_17587,N_16368,N_16571);
or U17588 (N_17588,N_16340,N_16698);
or U17589 (N_17589,N_16933,N_16957);
nand U17590 (N_17590,N_16155,N_16316);
and U17591 (N_17591,N_16341,N_16441);
nor U17592 (N_17592,N_16965,N_16847);
nand U17593 (N_17593,N_16412,N_16944);
or U17594 (N_17594,N_16482,N_16319);
nor U17595 (N_17595,N_16581,N_16879);
or U17596 (N_17596,N_16893,N_16622);
xnor U17597 (N_17597,N_16439,N_16305);
xor U17598 (N_17598,N_16135,N_16664);
or U17599 (N_17599,N_16371,N_16972);
xor U17600 (N_17600,N_16690,N_16721);
and U17601 (N_17601,N_16680,N_16317);
xnor U17602 (N_17602,N_16440,N_16490);
and U17603 (N_17603,N_16782,N_16768);
xnor U17604 (N_17604,N_16079,N_16589);
and U17605 (N_17605,N_16932,N_16771);
nand U17606 (N_17606,N_16312,N_16046);
and U17607 (N_17607,N_16205,N_16465);
xor U17608 (N_17608,N_16178,N_16797);
nor U17609 (N_17609,N_16588,N_16787);
or U17610 (N_17610,N_16235,N_16403);
nand U17611 (N_17611,N_16502,N_16338);
xnor U17612 (N_17612,N_16021,N_16990);
and U17613 (N_17613,N_16113,N_16460);
and U17614 (N_17614,N_16333,N_16790);
nor U17615 (N_17615,N_16983,N_16509);
or U17616 (N_17616,N_16914,N_16021);
nand U17617 (N_17617,N_16779,N_16792);
xnor U17618 (N_17618,N_16013,N_16915);
nor U17619 (N_17619,N_16429,N_16239);
nand U17620 (N_17620,N_16236,N_16402);
and U17621 (N_17621,N_16239,N_16821);
nor U17622 (N_17622,N_16190,N_16902);
and U17623 (N_17623,N_16688,N_16402);
or U17624 (N_17624,N_16058,N_16725);
or U17625 (N_17625,N_16643,N_16242);
and U17626 (N_17626,N_16863,N_16313);
xor U17627 (N_17627,N_16726,N_16188);
and U17628 (N_17628,N_16417,N_16763);
and U17629 (N_17629,N_16476,N_16435);
nor U17630 (N_17630,N_16294,N_16734);
or U17631 (N_17631,N_16271,N_16133);
xor U17632 (N_17632,N_16169,N_16162);
and U17633 (N_17633,N_16358,N_16417);
xor U17634 (N_17634,N_16326,N_16572);
or U17635 (N_17635,N_16711,N_16768);
nor U17636 (N_17636,N_16555,N_16530);
xor U17637 (N_17637,N_16329,N_16241);
nor U17638 (N_17638,N_16829,N_16435);
nor U17639 (N_17639,N_16138,N_16515);
xor U17640 (N_17640,N_16208,N_16632);
or U17641 (N_17641,N_16347,N_16718);
nor U17642 (N_17642,N_16614,N_16437);
or U17643 (N_17643,N_16791,N_16780);
xnor U17644 (N_17644,N_16620,N_16225);
nor U17645 (N_17645,N_16398,N_16652);
xnor U17646 (N_17646,N_16685,N_16562);
or U17647 (N_17647,N_16386,N_16832);
xor U17648 (N_17648,N_16046,N_16302);
and U17649 (N_17649,N_16790,N_16593);
xnor U17650 (N_17650,N_16713,N_16287);
xor U17651 (N_17651,N_16795,N_16217);
nor U17652 (N_17652,N_16529,N_16958);
nor U17653 (N_17653,N_16659,N_16860);
xor U17654 (N_17654,N_16943,N_16144);
and U17655 (N_17655,N_16421,N_16978);
nor U17656 (N_17656,N_16903,N_16840);
nor U17657 (N_17657,N_16790,N_16200);
nand U17658 (N_17658,N_16291,N_16478);
and U17659 (N_17659,N_16125,N_16857);
or U17660 (N_17660,N_16497,N_16090);
and U17661 (N_17661,N_16910,N_16882);
or U17662 (N_17662,N_16472,N_16258);
and U17663 (N_17663,N_16113,N_16526);
and U17664 (N_17664,N_16653,N_16439);
nand U17665 (N_17665,N_16402,N_16443);
nor U17666 (N_17666,N_16057,N_16199);
nand U17667 (N_17667,N_16325,N_16962);
nand U17668 (N_17668,N_16816,N_16586);
nor U17669 (N_17669,N_16163,N_16923);
and U17670 (N_17670,N_16540,N_16915);
xor U17671 (N_17671,N_16858,N_16090);
and U17672 (N_17672,N_16066,N_16621);
nor U17673 (N_17673,N_16473,N_16408);
nor U17674 (N_17674,N_16931,N_16534);
xor U17675 (N_17675,N_16294,N_16201);
or U17676 (N_17676,N_16756,N_16729);
nand U17677 (N_17677,N_16932,N_16379);
xor U17678 (N_17678,N_16243,N_16936);
and U17679 (N_17679,N_16641,N_16731);
nor U17680 (N_17680,N_16343,N_16141);
xnor U17681 (N_17681,N_16699,N_16658);
and U17682 (N_17682,N_16347,N_16282);
xor U17683 (N_17683,N_16013,N_16819);
xnor U17684 (N_17684,N_16802,N_16868);
and U17685 (N_17685,N_16853,N_16391);
xnor U17686 (N_17686,N_16244,N_16147);
and U17687 (N_17687,N_16633,N_16492);
nor U17688 (N_17688,N_16693,N_16666);
xnor U17689 (N_17689,N_16616,N_16097);
xnor U17690 (N_17690,N_16740,N_16476);
xor U17691 (N_17691,N_16528,N_16425);
or U17692 (N_17692,N_16110,N_16753);
and U17693 (N_17693,N_16060,N_16926);
or U17694 (N_17694,N_16394,N_16180);
or U17695 (N_17695,N_16331,N_16057);
nor U17696 (N_17696,N_16936,N_16927);
xor U17697 (N_17697,N_16662,N_16482);
and U17698 (N_17698,N_16213,N_16322);
nor U17699 (N_17699,N_16852,N_16065);
nor U17700 (N_17700,N_16404,N_16956);
or U17701 (N_17701,N_16412,N_16704);
nand U17702 (N_17702,N_16818,N_16036);
and U17703 (N_17703,N_16890,N_16257);
nand U17704 (N_17704,N_16265,N_16389);
or U17705 (N_17705,N_16805,N_16654);
nor U17706 (N_17706,N_16428,N_16921);
or U17707 (N_17707,N_16339,N_16168);
nand U17708 (N_17708,N_16573,N_16506);
or U17709 (N_17709,N_16539,N_16031);
nand U17710 (N_17710,N_16840,N_16769);
nor U17711 (N_17711,N_16201,N_16455);
xor U17712 (N_17712,N_16161,N_16845);
and U17713 (N_17713,N_16942,N_16921);
xnor U17714 (N_17714,N_16922,N_16997);
and U17715 (N_17715,N_16058,N_16437);
xor U17716 (N_17716,N_16370,N_16239);
or U17717 (N_17717,N_16448,N_16254);
xor U17718 (N_17718,N_16125,N_16395);
and U17719 (N_17719,N_16517,N_16500);
and U17720 (N_17720,N_16012,N_16179);
and U17721 (N_17721,N_16730,N_16935);
and U17722 (N_17722,N_16291,N_16531);
or U17723 (N_17723,N_16009,N_16057);
nand U17724 (N_17724,N_16896,N_16792);
or U17725 (N_17725,N_16892,N_16384);
nand U17726 (N_17726,N_16432,N_16414);
nor U17727 (N_17727,N_16376,N_16498);
xnor U17728 (N_17728,N_16291,N_16682);
nand U17729 (N_17729,N_16773,N_16645);
and U17730 (N_17730,N_16028,N_16281);
xnor U17731 (N_17731,N_16755,N_16593);
nor U17732 (N_17732,N_16927,N_16605);
or U17733 (N_17733,N_16691,N_16011);
nand U17734 (N_17734,N_16474,N_16220);
and U17735 (N_17735,N_16383,N_16553);
xor U17736 (N_17736,N_16345,N_16076);
nand U17737 (N_17737,N_16223,N_16497);
nor U17738 (N_17738,N_16966,N_16060);
or U17739 (N_17739,N_16048,N_16218);
nor U17740 (N_17740,N_16117,N_16046);
and U17741 (N_17741,N_16844,N_16551);
and U17742 (N_17742,N_16140,N_16499);
nand U17743 (N_17743,N_16926,N_16532);
xor U17744 (N_17744,N_16578,N_16440);
or U17745 (N_17745,N_16094,N_16563);
or U17746 (N_17746,N_16113,N_16137);
and U17747 (N_17747,N_16430,N_16413);
or U17748 (N_17748,N_16864,N_16748);
xnor U17749 (N_17749,N_16405,N_16610);
nor U17750 (N_17750,N_16021,N_16090);
nor U17751 (N_17751,N_16169,N_16582);
or U17752 (N_17752,N_16137,N_16165);
and U17753 (N_17753,N_16618,N_16619);
xor U17754 (N_17754,N_16921,N_16071);
and U17755 (N_17755,N_16445,N_16816);
xor U17756 (N_17756,N_16637,N_16127);
nand U17757 (N_17757,N_16689,N_16589);
and U17758 (N_17758,N_16347,N_16566);
xor U17759 (N_17759,N_16553,N_16470);
xor U17760 (N_17760,N_16954,N_16503);
or U17761 (N_17761,N_16429,N_16788);
nor U17762 (N_17762,N_16945,N_16190);
nor U17763 (N_17763,N_16567,N_16089);
and U17764 (N_17764,N_16140,N_16090);
xor U17765 (N_17765,N_16807,N_16315);
nand U17766 (N_17766,N_16093,N_16968);
nor U17767 (N_17767,N_16471,N_16416);
nor U17768 (N_17768,N_16978,N_16947);
nor U17769 (N_17769,N_16182,N_16506);
xor U17770 (N_17770,N_16778,N_16239);
or U17771 (N_17771,N_16362,N_16681);
and U17772 (N_17772,N_16512,N_16651);
or U17773 (N_17773,N_16132,N_16807);
xnor U17774 (N_17774,N_16596,N_16060);
nand U17775 (N_17775,N_16141,N_16563);
and U17776 (N_17776,N_16073,N_16385);
and U17777 (N_17777,N_16838,N_16886);
or U17778 (N_17778,N_16107,N_16218);
or U17779 (N_17779,N_16954,N_16203);
xor U17780 (N_17780,N_16652,N_16384);
nor U17781 (N_17781,N_16339,N_16181);
and U17782 (N_17782,N_16014,N_16971);
and U17783 (N_17783,N_16021,N_16359);
xor U17784 (N_17784,N_16290,N_16769);
and U17785 (N_17785,N_16231,N_16644);
or U17786 (N_17786,N_16322,N_16537);
xor U17787 (N_17787,N_16781,N_16974);
nand U17788 (N_17788,N_16048,N_16478);
or U17789 (N_17789,N_16062,N_16784);
xor U17790 (N_17790,N_16342,N_16228);
and U17791 (N_17791,N_16199,N_16936);
nand U17792 (N_17792,N_16807,N_16712);
nand U17793 (N_17793,N_16917,N_16979);
or U17794 (N_17794,N_16530,N_16273);
xnor U17795 (N_17795,N_16197,N_16012);
xnor U17796 (N_17796,N_16110,N_16019);
xnor U17797 (N_17797,N_16993,N_16554);
nor U17798 (N_17798,N_16758,N_16084);
and U17799 (N_17799,N_16172,N_16151);
xnor U17800 (N_17800,N_16561,N_16765);
nor U17801 (N_17801,N_16939,N_16545);
xnor U17802 (N_17802,N_16810,N_16691);
xnor U17803 (N_17803,N_16505,N_16465);
xnor U17804 (N_17804,N_16689,N_16938);
nor U17805 (N_17805,N_16013,N_16791);
nand U17806 (N_17806,N_16759,N_16420);
xnor U17807 (N_17807,N_16333,N_16959);
nand U17808 (N_17808,N_16560,N_16518);
nor U17809 (N_17809,N_16680,N_16677);
and U17810 (N_17810,N_16296,N_16062);
xnor U17811 (N_17811,N_16797,N_16769);
or U17812 (N_17812,N_16279,N_16625);
and U17813 (N_17813,N_16636,N_16284);
nand U17814 (N_17814,N_16278,N_16326);
nor U17815 (N_17815,N_16432,N_16734);
or U17816 (N_17816,N_16456,N_16877);
nand U17817 (N_17817,N_16018,N_16837);
nor U17818 (N_17818,N_16631,N_16925);
nand U17819 (N_17819,N_16951,N_16395);
and U17820 (N_17820,N_16718,N_16560);
nor U17821 (N_17821,N_16653,N_16661);
xnor U17822 (N_17822,N_16241,N_16937);
or U17823 (N_17823,N_16624,N_16498);
and U17824 (N_17824,N_16340,N_16166);
nand U17825 (N_17825,N_16994,N_16648);
nor U17826 (N_17826,N_16674,N_16488);
or U17827 (N_17827,N_16413,N_16347);
or U17828 (N_17828,N_16691,N_16813);
nor U17829 (N_17829,N_16536,N_16030);
and U17830 (N_17830,N_16191,N_16093);
nand U17831 (N_17831,N_16144,N_16063);
nor U17832 (N_17832,N_16234,N_16447);
xor U17833 (N_17833,N_16609,N_16778);
nand U17834 (N_17834,N_16270,N_16670);
or U17835 (N_17835,N_16420,N_16089);
and U17836 (N_17836,N_16791,N_16149);
xnor U17837 (N_17837,N_16763,N_16316);
nor U17838 (N_17838,N_16076,N_16521);
and U17839 (N_17839,N_16320,N_16486);
and U17840 (N_17840,N_16403,N_16674);
nor U17841 (N_17841,N_16155,N_16038);
and U17842 (N_17842,N_16287,N_16886);
xor U17843 (N_17843,N_16662,N_16555);
or U17844 (N_17844,N_16034,N_16385);
and U17845 (N_17845,N_16144,N_16988);
nor U17846 (N_17846,N_16368,N_16703);
or U17847 (N_17847,N_16757,N_16293);
nor U17848 (N_17848,N_16347,N_16875);
and U17849 (N_17849,N_16176,N_16590);
or U17850 (N_17850,N_16348,N_16851);
nor U17851 (N_17851,N_16347,N_16222);
nor U17852 (N_17852,N_16440,N_16351);
xnor U17853 (N_17853,N_16077,N_16657);
xnor U17854 (N_17854,N_16297,N_16830);
nand U17855 (N_17855,N_16553,N_16371);
or U17856 (N_17856,N_16154,N_16952);
nor U17857 (N_17857,N_16248,N_16714);
xor U17858 (N_17858,N_16243,N_16272);
nand U17859 (N_17859,N_16521,N_16953);
nand U17860 (N_17860,N_16777,N_16453);
and U17861 (N_17861,N_16063,N_16107);
xor U17862 (N_17862,N_16743,N_16789);
and U17863 (N_17863,N_16488,N_16600);
nand U17864 (N_17864,N_16548,N_16594);
xnor U17865 (N_17865,N_16002,N_16493);
xnor U17866 (N_17866,N_16256,N_16336);
nor U17867 (N_17867,N_16140,N_16779);
nor U17868 (N_17868,N_16303,N_16590);
nor U17869 (N_17869,N_16231,N_16868);
xnor U17870 (N_17870,N_16581,N_16631);
nor U17871 (N_17871,N_16913,N_16979);
and U17872 (N_17872,N_16873,N_16421);
xor U17873 (N_17873,N_16036,N_16552);
nor U17874 (N_17874,N_16433,N_16034);
nand U17875 (N_17875,N_16322,N_16524);
or U17876 (N_17876,N_16371,N_16684);
or U17877 (N_17877,N_16392,N_16543);
xor U17878 (N_17878,N_16613,N_16278);
and U17879 (N_17879,N_16048,N_16972);
xnor U17880 (N_17880,N_16067,N_16167);
and U17881 (N_17881,N_16283,N_16344);
or U17882 (N_17882,N_16868,N_16622);
xnor U17883 (N_17883,N_16986,N_16919);
nor U17884 (N_17884,N_16620,N_16813);
nand U17885 (N_17885,N_16148,N_16908);
or U17886 (N_17886,N_16477,N_16790);
or U17887 (N_17887,N_16493,N_16373);
nor U17888 (N_17888,N_16945,N_16516);
nor U17889 (N_17889,N_16643,N_16103);
and U17890 (N_17890,N_16813,N_16146);
and U17891 (N_17891,N_16358,N_16869);
nand U17892 (N_17892,N_16156,N_16525);
and U17893 (N_17893,N_16694,N_16072);
or U17894 (N_17894,N_16060,N_16237);
xnor U17895 (N_17895,N_16966,N_16487);
or U17896 (N_17896,N_16235,N_16845);
xnor U17897 (N_17897,N_16143,N_16471);
or U17898 (N_17898,N_16926,N_16617);
or U17899 (N_17899,N_16292,N_16434);
nor U17900 (N_17900,N_16315,N_16434);
xnor U17901 (N_17901,N_16368,N_16709);
nand U17902 (N_17902,N_16694,N_16270);
nand U17903 (N_17903,N_16630,N_16395);
and U17904 (N_17904,N_16666,N_16023);
xnor U17905 (N_17905,N_16812,N_16462);
or U17906 (N_17906,N_16243,N_16908);
xnor U17907 (N_17907,N_16433,N_16867);
nor U17908 (N_17908,N_16765,N_16260);
nand U17909 (N_17909,N_16722,N_16657);
or U17910 (N_17910,N_16701,N_16061);
xor U17911 (N_17911,N_16453,N_16199);
and U17912 (N_17912,N_16823,N_16010);
xor U17913 (N_17913,N_16072,N_16822);
xor U17914 (N_17914,N_16822,N_16222);
nand U17915 (N_17915,N_16443,N_16118);
xnor U17916 (N_17916,N_16770,N_16146);
nand U17917 (N_17917,N_16022,N_16483);
and U17918 (N_17918,N_16958,N_16642);
xnor U17919 (N_17919,N_16931,N_16887);
nor U17920 (N_17920,N_16686,N_16561);
xnor U17921 (N_17921,N_16397,N_16534);
and U17922 (N_17922,N_16541,N_16985);
xor U17923 (N_17923,N_16955,N_16255);
nand U17924 (N_17924,N_16562,N_16387);
or U17925 (N_17925,N_16472,N_16662);
nor U17926 (N_17926,N_16315,N_16928);
or U17927 (N_17927,N_16468,N_16991);
nor U17928 (N_17928,N_16291,N_16382);
nor U17929 (N_17929,N_16219,N_16229);
or U17930 (N_17930,N_16147,N_16493);
or U17931 (N_17931,N_16466,N_16516);
nand U17932 (N_17932,N_16925,N_16003);
or U17933 (N_17933,N_16189,N_16762);
xnor U17934 (N_17934,N_16265,N_16485);
and U17935 (N_17935,N_16251,N_16788);
xor U17936 (N_17936,N_16150,N_16228);
or U17937 (N_17937,N_16149,N_16007);
and U17938 (N_17938,N_16600,N_16884);
nand U17939 (N_17939,N_16864,N_16962);
and U17940 (N_17940,N_16578,N_16909);
nor U17941 (N_17941,N_16416,N_16999);
nand U17942 (N_17942,N_16696,N_16027);
nor U17943 (N_17943,N_16514,N_16895);
and U17944 (N_17944,N_16677,N_16435);
or U17945 (N_17945,N_16534,N_16277);
and U17946 (N_17946,N_16700,N_16951);
xor U17947 (N_17947,N_16724,N_16008);
and U17948 (N_17948,N_16833,N_16202);
xnor U17949 (N_17949,N_16534,N_16109);
nand U17950 (N_17950,N_16224,N_16751);
nor U17951 (N_17951,N_16802,N_16825);
xor U17952 (N_17952,N_16037,N_16200);
or U17953 (N_17953,N_16750,N_16554);
and U17954 (N_17954,N_16896,N_16318);
nor U17955 (N_17955,N_16721,N_16895);
nand U17956 (N_17956,N_16270,N_16108);
or U17957 (N_17957,N_16062,N_16138);
nor U17958 (N_17958,N_16680,N_16839);
nand U17959 (N_17959,N_16457,N_16652);
or U17960 (N_17960,N_16404,N_16955);
and U17961 (N_17961,N_16137,N_16530);
and U17962 (N_17962,N_16742,N_16044);
nand U17963 (N_17963,N_16440,N_16684);
or U17964 (N_17964,N_16673,N_16920);
nand U17965 (N_17965,N_16534,N_16827);
nand U17966 (N_17966,N_16589,N_16816);
xor U17967 (N_17967,N_16329,N_16337);
and U17968 (N_17968,N_16520,N_16712);
nand U17969 (N_17969,N_16625,N_16724);
or U17970 (N_17970,N_16349,N_16343);
and U17971 (N_17971,N_16582,N_16316);
and U17972 (N_17972,N_16504,N_16608);
or U17973 (N_17973,N_16768,N_16889);
nand U17974 (N_17974,N_16400,N_16204);
or U17975 (N_17975,N_16268,N_16137);
and U17976 (N_17976,N_16399,N_16275);
nor U17977 (N_17977,N_16313,N_16314);
xnor U17978 (N_17978,N_16498,N_16994);
and U17979 (N_17979,N_16158,N_16743);
xnor U17980 (N_17980,N_16723,N_16810);
nand U17981 (N_17981,N_16446,N_16297);
and U17982 (N_17982,N_16118,N_16594);
and U17983 (N_17983,N_16068,N_16694);
nand U17984 (N_17984,N_16277,N_16285);
nand U17985 (N_17985,N_16558,N_16127);
nand U17986 (N_17986,N_16786,N_16264);
xnor U17987 (N_17987,N_16406,N_16301);
or U17988 (N_17988,N_16769,N_16748);
xor U17989 (N_17989,N_16986,N_16856);
and U17990 (N_17990,N_16072,N_16359);
or U17991 (N_17991,N_16982,N_16558);
and U17992 (N_17992,N_16156,N_16630);
nand U17993 (N_17993,N_16404,N_16115);
nor U17994 (N_17994,N_16451,N_16716);
and U17995 (N_17995,N_16169,N_16388);
nor U17996 (N_17996,N_16191,N_16010);
or U17997 (N_17997,N_16371,N_16926);
nor U17998 (N_17998,N_16363,N_16842);
nor U17999 (N_17999,N_16131,N_16552);
xnor U18000 (N_18000,N_17282,N_17513);
nand U18001 (N_18001,N_17512,N_17619);
xnor U18002 (N_18002,N_17386,N_17889);
nor U18003 (N_18003,N_17362,N_17315);
nand U18004 (N_18004,N_17924,N_17859);
or U18005 (N_18005,N_17874,N_17931);
and U18006 (N_18006,N_17661,N_17450);
nand U18007 (N_18007,N_17254,N_17920);
nor U18008 (N_18008,N_17652,N_17674);
and U18009 (N_18009,N_17142,N_17430);
xor U18010 (N_18010,N_17785,N_17480);
and U18011 (N_18011,N_17197,N_17022);
or U18012 (N_18012,N_17606,N_17101);
or U18013 (N_18013,N_17326,N_17981);
nor U18014 (N_18014,N_17568,N_17995);
and U18015 (N_18015,N_17733,N_17983);
xnor U18016 (N_18016,N_17387,N_17530);
and U18017 (N_18017,N_17626,N_17697);
nand U18018 (N_18018,N_17237,N_17737);
or U18019 (N_18019,N_17992,N_17514);
xor U18020 (N_18020,N_17541,N_17989);
xnor U18021 (N_18021,N_17922,N_17336);
or U18022 (N_18022,N_17456,N_17267);
nor U18023 (N_18023,N_17919,N_17018);
nor U18024 (N_18024,N_17609,N_17420);
and U18025 (N_18025,N_17104,N_17993);
xnor U18026 (N_18026,N_17586,N_17975);
nand U18027 (N_18027,N_17719,N_17881);
nand U18028 (N_18028,N_17232,N_17249);
and U18029 (N_18029,N_17896,N_17778);
nand U18030 (N_18030,N_17521,N_17890);
and U18031 (N_18031,N_17219,N_17167);
nand U18032 (N_18032,N_17478,N_17926);
or U18033 (N_18033,N_17903,N_17441);
or U18034 (N_18034,N_17868,N_17509);
nand U18035 (N_18035,N_17062,N_17696);
or U18036 (N_18036,N_17321,N_17493);
nand U18037 (N_18037,N_17687,N_17349);
xnor U18038 (N_18038,N_17694,N_17345);
nor U18039 (N_18039,N_17297,N_17431);
or U18040 (N_18040,N_17375,N_17414);
nor U18041 (N_18041,N_17632,N_17229);
nand U18042 (N_18042,N_17762,N_17986);
xor U18043 (N_18043,N_17793,N_17819);
or U18044 (N_18044,N_17372,N_17141);
or U18045 (N_18045,N_17335,N_17873);
nand U18046 (N_18046,N_17002,N_17777);
xnor U18047 (N_18047,N_17550,N_17089);
xor U18048 (N_18048,N_17436,N_17581);
xnor U18049 (N_18049,N_17798,N_17157);
xnor U18050 (N_18050,N_17394,N_17534);
nand U18051 (N_18051,N_17753,N_17973);
and U18052 (N_18052,N_17474,N_17090);
xor U18053 (N_18053,N_17111,N_17880);
nor U18054 (N_18054,N_17004,N_17502);
xnor U18055 (N_18055,N_17013,N_17154);
or U18056 (N_18056,N_17221,N_17806);
nand U18057 (N_18057,N_17065,N_17875);
and U18058 (N_18058,N_17510,N_17852);
or U18059 (N_18059,N_17392,N_17312);
or U18060 (N_18060,N_17127,N_17564);
and U18061 (N_18061,N_17884,N_17311);
and U18062 (N_18062,N_17941,N_17817);
xor U18063 (N_18063,N_17956,N_17664);
or U18064 (N_18064,N_17938,N_17908);
xnor U18065 (N_18065,N_17342,N_17485);
nor U18066 (N_18066,N_17608,N_17073);
or U18067 (N_18067,N_17505,N_17855);
nor U18068 (N_18068,N_17287,N_17066);
nand U18069 (N_18069,N_17883,N_17932);
and U18070 (N_18070,N_17400,N_17069);
nor U18071 (N_18071,N_17594,N_17252);
xor U18072 (N_18072,N_17088,N_17198);
and U18073 (N_18073,N_17904,N_17113);
nand U18074 (N_18074,N_17792,N_17290);
and U18075 (N_18075,N_17517,N_17729);
xor U18076 (N_18076,N_17028,N_17424);
or U18077 (N_18077,N_17757,N_17155);
nand U18078 (N_18078,N_17508,N_17364);
and U18079 (N_18079,N_17279,N_17166);
xnor U18080 (N_18080,N_17948,N_17208);
or U18081 (N_18081,N_17280,N_17681);
nor U18082 (N_18082,N_17132,N_17548);
nor U18083 (N_18083,N_17196,N_17228);
xor U18084 (N_18084,N_17341,N_17026);
and U18085 (N_18085,N_17363,N_17921);
or U18086 (N_18086,N_17707,N_17476);
nand U18087 (N_18087,N_17909,N_17783);
xor U18088 (N_18088,N_17153,N_17080);
nand U18089 (N_18089,N_17771,N_17620);
or U18090 (N_18090,N_17828,N_17291);
nor U18091 (N_18091,N_17499,N_17987);
xor U18092 (N_18092,N_17751,N_17827);
xor U18093 (N_18093,N_17288,N_17665);
nand U18094 (N_18094,N_17850,N_17683);
xnor U18095 (N_18095,N_17805,N_17218);
nand U18096 (N_18096,N_17329,N_17091);
or U18097 (N_18097,N_17325,N_17555);
xor U18098 (N_18098,N_17255,N_17444);
xnor U18099 (N_18099,N_17865,N_17982);
and U18100 (N_18100,N_17801,N_17671);
xor U18101 (N_18101,N_17901,N_17007);
nor U18102 (N_18102,N_17712,N_17575);
nand U18103 (N_18103,N_17054,N_17577);
or U18104 (N_18104,N_17123,N_17727);
and U18105 (N_18105,N_17624,N_17454);
nand U18106 (N_18106,N_17092,N_17536);
and U18107 (N_18107,N_17409,N_17231);
nor U18108 (N_18108,N_17690,N_17673);
nor U18109 (N_18109,N_17570,N_17885);
or U18110 (N_18110,N_17437,N_17899);
nand U18111 (N_18111,N_17718,N_17782);
or U18112 (N_18112,N_17257,N_17537);
nor U18113 (N_18113,N_17067,N_17892);
nor U18114 (N_18114,N_17945,N_17204);
and U18115 (N_18115,N_17466,N_17274);
and U18116 (N_18116,N_17128,N_17377);
xor U18117 (N_18117,N_17809,N_17121);
nor U18118 (N_18118,N_17452,N_17693);
or U18119 (N_18119,N_17445,N_17724);
xor U18120 (N_18120,N_17049,N_17005);
nand U18121 (N_18121,N_17864,N_17172);
nand U18122 (N_18122,N_17563,N_17650);
nand U18123 (N_18123,N_17600,N_17680);
xor U18124 (N_18124,N_17569,N_17578);
xor U18125 (N_18125,N_17976,N_17937);
or U18126 (N_18126,N_17872,N_17604);
and U18127 (N_18127,N_17455,N_17222);
nor U18128 (N_18128,N_17784,N_17384);
and U18129 (N_18129,N_17776,N_17471);
or U18130 (N_18130,N_17348,N_17126);
nor U18131 (N_18131,N_17567,N_17081);
nor U18132 (N_18132,N_17266,N_17678);
xor U18133 (N_18133,N_17496,N_17915);
nand U18134 (N_18134,N_17191,N_17518);
and U18135 (N_18135,N_17843,N_17971);
or U18136 (N_18136,N_17284,N_17658);
nand U18137 (N_18137,N_17957,N_17648);
nor U18138 (N_18138,N_17482,N_17950);
or U18139 (N_18139,N_17756,N_17882);
xnor U18140 (N_18140,N_17935,N_17415);
nand U18141 (N_18141,N_17391,N_17192);
nor U18142 (N_18142,N_17395,N_17333);
or U18143 (N_18143,N_17133,N_17587);
nand U18144 (N_18144,N_17877,N_17492);
nand U18145 (N_18145,N_17876,N_17645);
nand U18146 (N_18146,N_17692,N_17105);
nor U18147 (N_18147,N_17438,N_17140);
nor U18148 (N_18148,N_17403,N_17497);
nor U18149 (N_18149,N_17490,N_17344);
nor U18150 (N_18150,N_17826,N_17780);
nor U18151 (N_18151,N_17009,N_17070);
or U18152 (N_18152,N_17230,N_17553);
and U18153 (N_18153,N_17754,N_17636);
nor U18154 (N_18154,N_17786,N_17347);
nand U18155 (N_18155,N_17682,N_17309);
nand U18156 (N_18156,N_17177,N_17135);
xor U18157 (N_18157,N_17405,N_17103);
nor U18158 (N_18158,N_17401,N_17353);
or U18159 (N_18159,N_17328,N_17406);
nor U18160 (N_18160,N_17464,N_17565);
or U18161 (N_18161,N_17432,N_17691);
and U18162 (N_18162,N_17745,N_17655);
and U18163 (N_18163,N_17633,N_17708);
and U18164 (N_18164,N_17419,N_17717);
or U18165 (N_18165,N_17841,N_17185);
nor U18166 (N_18166,N_17533,N_17029);
nand U18167 (N_18167,N_17589,N_17246);
or U18168 (N_18168,N_17138,N_17808);
nand U18169 (N_18169,N_17146,N_17357);
and U18170 (N_18170,N_17281,N_17775);
and U18171 (N_18171,N_17366,N_17407);
or U18172 (N_18172,N_17742,N_17412);
or U18173 (N_18173,N_17939,N_17598);
or U18174 (N_18174,N_17295,N_17851);
nor U18175 (N_18175,N_17726,N_17912);
or U18176 (N_18176,N_17358,N_17946);
or U18177 (N_18177,N_17794,N_17529);
and U18178 (N_18178,N_17764,N_17443);
and U18179 (N_18179,N_17878,N_17019);
nand U18180 (N_18180,N_17165,N_17559);
or U18181 (N_18181,N_17467,N_17170);
nand U18182 (N_18182,N_17867,N_17151);
xor U18183 (N_18183,N_17458,N_17902);
nand U18184 (N_18184,N_17593,N_17398);
nand U18185 (N_18185,N_17035,N_17913);
and U18186 (N_18186,N_17831,N_17662);
or U18187 (N_18187,N_17447,N_17037);
nand U18188 (N_18188,N_17666,N_17985);
and U18189 (N_18189,N_17685,N_17887);
nor U18190 (N_18190,N_17747,N_17340);
xor U18191 (N_18191,N_17179,N_17317);
nor U18192 (N_18192,N_17709,N_17959);
xnor U18193 (N_18193,N_17207,N_17334);
or U18194 (N_18194,N_17916,N_17265);
and U18195 (N_18195,N_17905,N_17383);
and U18196 (N_18196,N_17519,N_17316);
nor U18197 (N_18197,N_17917,N_17791);
xnor U18198 (N_18198,N_17053,N_17156);
nand U18199 (N_18199,N_17145,N_17839);
xnor U18200 (N_18200,N_17462,N_17623);
or U18201 (N_18201,N_17094,N_17251);
and U18202 (N_18202,N_17322,N_17356);
or U18203 (N_18203,N_17077,N_17253);
nand U18204 (N_18204,N_17417,N_17974);
nor U18205 (N_18205,N_17642,N_17630);
or U18206 (N_18206,N_17711,N_17927);
and U18207 (N_18207,N_17720,N_17670);
and U18208 (N_18208,N_17731,N_17571);
nor U18209 (N_18209,N_17557,N_17410);
xnor U18210 (N_18210,N_17675,N_17660);
nand U18211 (N_18211,N_17668,N_17484);
nand U18212 (N_18212,N_17591,N_17108);
nor U18213 (N_18213,N_17433,N_17998);
or U18214 (N_18214,N_17829,N_17134);
nor U18215 (N_18215,N_17672,N_17639);
or U18216 (N_18216,N_17629,N_17465);
nor U18217 (N_18217,N_17840,N_17501);
xor U18218 (N_18218,N_17730,N_17136);
or U18219 (N_18219,N_17008,N_17857);
nand U18220 (N_18220,N_17679,N_17379);
or U18221 (N_18221,N_17283,N_17583);
or U18222 (N_18222,N_17725,N_17016);
nand U18223 (N_18223,N_17503,N_17750);
nor U18224 (N_18224,N_17977,N_17178);
xnor U18225 (N_18225,N_17030,N_17821);
or U18226 (N_18226,N_17504,N_17241);
and U18227 (N_18227,N_17343,N_17175);
nor U18228 (N_18228,N_17285,N_17300);
or U18229 (N_18229,N_17886,N_17301);
nand U18230 (N_18230,N_17399,N_17148);
nand U18231 (N_18231,N_17582,N_17338);
xor U18232 (N_18232,N_17050,N_17996);
xnor U18233 (N_18233,N_17802,N_17041);
xor U18234 (N_18234,N_17027,N_17954);
or U18235 (N_18235,N_17273,N_17527);
and U18236 (N_18236,N_17271,N_17525);
nand U18237 (N_18237,N_17614,N_17613);
nand U18238 (N_18238,N_17597,N_17900);
nor U18239 (N_18239,N_17048,N_17327);
nand U18240 (N_18240,N_17728,N_17515);
and U18241 (N_18241,N_17769,N_17421);
xor U18242 (N_18242,N_17923,N_17256);
or U18243 (N_18243,N_17914,N_17483);
nand U18244 (N_18244,N_17098,N_17699);
or U18245 (N_18245,N_17663,N_17084);
or U18246 (N_18246,N_17184,N_17055);
nor U18247 (N_18247,N_17440,N_17314);
nand U18248 (N_18248,N_17735,N_17446);
and U18249 (N_18249,N_17137,N_17930);
xnor U18250 (N_18250,N_17910,N_17180);
nand U18251 (N_18251,N_17816,N_17962);
xnor U18252 (N_18252,N_17213,N_17427);
nand U18253 (N_18253,N_17052,N_17117);
and U18254 (N_18254,N_17031,N_17305);
nor U18255 (N_18255,N_17079,N_17997);
nor U18256 (N_18256,N_17835,N_17631);
nand U18257 (N_18257,N_17804,N_17122);
or U18258 (N_18258,N_17990,N_17226);
nor U18259 (N_18259,N_17324,N_17918);
nand U18260 (N_18260,N_17547,N_17369);
and U18261 (N_18261,N_17741,N_17303);
and U18262 (N_18262,N_17893,N_17261);
nand U18263 (N_18263,N_17595,N_17834);
or U18264 (N_18264,N_17772,N_17763);
nand U18265 (N_18265,N_17698,N_17934);
and U18266 (N_18266,N_17034,N_17715);
or U18267 (N_18267,N_17380,N_17020);
and U18268 (N_18268,N_17500,N_17714);
xor U18269 (N_18269,N_17453,N_17602);
or U18270 (N_18270,N_17516,N_17980);
nor U18271 (N_18271,N_17259,N_17473);
nand U18272 (N_18272,N_17612,N_17109);
and U18273 (N_18273,N_17949,N_17072);
and U18274 (N_18274,N_17195,N_17641);
xnor U18275 (N_18275,N_17649,N_17964);
nand U18276 (N_18276,N_17732,N_17451);
nand U18277 (N_18277,N_17734,N_17790);
and U18278 (N_18278,N_17248,N_17118);
nand U18279 (N_18279,N_17528,N_17460);
nand U18280 (N_18280,N_17965,N_17540);
nor U18281 (N_18281,N_17339,N_17224);
nand U18282 (N_18282,N_17489,N_17546);
xor U18283 (N_18283,N_17056,N_17585);
and U18284 (N_18284,N_17523,N_17599);
or U18285 (N_18285,N_17045,N_17955);
nand U18286 (N_18286,N_17319,N_17183);
or U18287 (N_18287,N_17713,N_17627);
xor U18288 (N_18288,N_17129,N_17243);
and U18289 (N_18289,N_17242,N_17758);
nor U18290 (N_18290,N_17706,N_17220);
xor U18291 (N_18291,N_17173,N_17078);
and U18292 (N_18292,N_17272,N_17535);
xor U18293 (N_18293,N_17097,N_17071);
or U18294 (N_18294,N_17355,N_17833);
nor U18295 (N_18295,N_17238,N_17203);
nor U18296 (N_18296,N_17160,N_17469);
xnor U18297 (N_18297,N_17601,N_17161);
or U18298 (N_18298,N_17488,N_17032);
or U18299 (N_18299,N_17388,N_17023);
and U18300 (N_18300,N_17051,N_17814);
nand U18301 (N_18301,N_17838,N_17187);
or U18302 (N_18302,N_17584,N_17190);
xor U18303 (N_18303,N_17573,N_17869);
nor U18304 (N_18304,N_17677,N_17643);
and U18305 (N_18305,N_17963,N_17233);
nand U18306 (N_18306,N_17799,N_17014);
or U18307 (N_18307,N_17147,N_17795);
nand U18308 (N_18308,N_17653,N_17688);
nand U18309 (N_18309,N_17162,N_17010);
nor U18310 (N_18310,N_17373,N_17657);
or U18311 (N_18311,N_17705,N_17944);
nor U18312 (N_18312,N_17991,N_17907);
nor U18313 (N_18313,N_17359,N_17526);
nand U18314 (N_18314,N_17545,N_17393);
or U18315 (N_18315,N_17367,N_17205);
nand U18316 (N_18316,N_17064,N_17001);
nand U18317 (N_18317,N_17209,N_17025);
and U18318 (N_18318,N_17561,N_17689);
xor U18319 (N_18319,N_17603,N_17552);
and U18320 (N_18320,N_17988,N_17434);
or U18321 (N_18321,N_17310,N_17223);
xnor U18322 (N_18322,N_17644,N_17656);
or U18323 (N_18323,N_17651,N_17235);
and U18324 (N_18324,N_17746,N_17115);
nand U18325 (N_18325,N_17539,N_17163);
or U18326 (N_18326,N_17592,N_17459);
nor U18327 (N_18327,N_17330,N_17667);
and U18328 (N_18328,N_17481,N_17350);
or U18329 (N_18329,N_17858,N_17374);
or U18330 (N_18330,N_17761,N_17871);
and U18331 (N_18331,N_17119,N_17788);
xnor U18332 (N_18332,N_17810,N_17087);
and U18333 (N_18333,N_17580,N_17640);
nor U18334 (N_18334,N_17891,N_17531);
xnor U18335 (N_18335,N_17418,N_17425);
nor U18336 (N_18336,N_17933,N_17862);
nor U18337 (N_18337,N_17498,N_17616);
xnor U18338 (N_18338,N_17625,N_17848);
nand U18339 (N_18339,N_17100,N_17402);
nor U18340 (N_18340,N_17770,N_17506);
nand U18341 (N_18341,N_17863,N_17378);
or U18342 (N_18342,N_17979,N_17302);
or U18343 (N_18343,N_17560,N_17442);
or U18344 (N_18344,N_17749,N_17532);
or U18345 (N_18345,N_17099,N_17385);
or U18346 (N_18346,N_17522,N_17800);
xor U18347 (N_18347,N_17046,N_17320);
nand U18348 (N_18348,N_17576,N_17365);
nor U18349 (N_18349,N_17943,N_17739);
nor U18350 (N_18350,N_17202,N_17174);
xnor U18351 (N_18351,N_17968,N_17461);
nand U18352 (N_18352,N_17086,N_17978);
nor U18353 (N_18353,N_17755,N_17368);
nand U18354 (N_18354,N_17736,N_17060);
nor U18355 (N_18355,N_17716,N_17003);
nand U18356 (N_18356,N_17618,N_17245);
nor U18357 (N_18357,N_17487,N_17429);
xor U18358 (N_18358,N_17928,N_17966);
xor U18359 (N_18359,N_17448,N_17842);
nor U18360 (N_18360,N_17063,N_17947);
xor U18361 (N_18361,N_17354,N_17846);
or U18362 (N_18362,N_17304,N_17370);
nor U18363 (N_18363,N_17176,N_17634);
xnor U18364 (N_18364,N_17646,N_17686);
nand U18365 (N_18365,N_17120,N_17960);
nor U18366 (N_18366,N_17942,N_17507);
nand U18367 (N_18367,N_17139,N_17813);
nor U18368 (N_18368,N_17389,N_17748);
nor U18369 (N_18369,N_17076,N_17044);
nand U18370 (N_18370,N_17796,N_17292);
nand U18371 (N_18371,N_17413,N_17217);
and U18372 (N_18372,N_17164,N_17970);
and U18373 (N_18373,N_17168,N_17404);
and U18374 (N_18374,N_17186,N_17866);
nand U18375 (N_18375,N_17972,N_17820);
nor U18376 (N_18376,N_17171,N_17012);
or U18377 (N_18377,N_17150,N_17566);
nor U18378 (N_18378,N_17210,N_17215);
or U18379 (N_18379,N_17061,N_17216);
and U18380 (N_18380,N_17610,N_17556);
or U18381 (N_18381,N_17611,N_17036);
nand U18382 (N_18382,N_17579,N_17486);
nor U18383 (N_18383,N_17247,N_17759);
nand U18384 (N_18384,N_17654,N_17635);
xnor U18385 (N_18385,N_17895,N_17520);
or U18386 (N_18386,N_17352,N_17953);
nand U18387 (N_18387,N_17894,N_17836);
nand U18388 (N_18388,N_17738,N_17040);
xnor U18389 (N_18389,N_17743,N_17017);
nand U18390 (N_18390,N_17428,N_17837);
xnor U18391 (N_18391,N_17225,N_17999);
nor U18392 (N_18392,N_17695,N_17194);
nand U18393 (N_18393,N_17083,N_17258);
nor U18394 (N_18394,N_17766,N_17371);
nor U18395 (N_18395,N_17189,N_17193);
xor U18396 (N_18396,N_17470,N_17449);
nor U18397 (N_18397,N_17463,N_17262);
xnor U18398 (N_18398,N_17306,N_17549);
or U18399 (N_18399,N_17144,N_17332);
nand U18400 (N_18400,N_17832,N_17308);
nand U18401 (N_18401,N_17472,N_17423);
nor U18402 (N_18402,N_17114,N_17936);
nor U18403 (N_18403,N_17058,N_17765);
nand U18404 (N_18404,N_17822,N_17376);
and U18405 (N_18405,N_17538,N_17110);
nand U18406 (N_18406,N_17382,N_17475);
nand U18407 (N_18407,N_17323,N_17879);
or U18408 (N_18408,N_17811,N_17264);
nand U18409 (N_18409,N_17787,N_17244);
nor U18410 (N_18410,N_17169,N_17059);
nor U18411 (N_18411,N_17477,N_17495);
xnor U18412 (N_18412,N_17422,N_17558);
nand U18413 (N_18413,N_17112,N_17408);
nand U18414 (N_18414,N_17268,N_17637);
and U18415 (N_18415,N_17125,N_17294);
nor U18416 (N_18416,N_17039,N_17085);
or U18417 (N_18417,N_17897,N_17823);
nand U18418 (N_18418,N_17906,N_17723);
nor U18419 (N_18419,N_17543,N_17298);
and U18420 (N_18420,N_17116,N_17607);
nor U18421 (N_18421,N_17011,N_17853);
and U18422 (N_18422,N_17617,N_17925);
or U18423 (N_18423,N_17830,N_17015);
xnor U18424 (N_18424,N_17812,N_17524);
nor U18425 (N_18425,N_17270,N_17337);
and U18426 (N_18426,N_17130,N_17621);
nor U18427 (N_18427,N_17106,N_17647);
xnor U18428 (N_18428,N_17752,N_17068);
or U18429 (N_18429,N_17006,N_17107);
nor U18430 (N_18430,N_17124,N_17701);
or U18431 (N_18431,N_17888,N_17313);
nand U18432 (N_18432,N_17331,N_17911);
nand U18433 (N_18433,N_17898,N_17562);
nor U18434 (N_18434,N_17622,N_17278);
nand U18435 (N_18435,N_17293,N_17596);
nand U18436 (N_18436,N_17958,N_17605);
xnor U18437 (N_18437,N_17703,N_17206);
nand U18438 (N_18438,N_17426,N_17744);
xor U18439 (N_18439,N_17275,N_17768);
xnor U18440 (N_18440,N_17149,N_17361);
xnor U18441 (N_18441,N_17082,N_17479);
or U18442 (N_18442,N_17269,N_17158);
and U18443 (N_18443,N_17860,N_17638);
xnor U18444 (N_18444,N_17074,N_17807);
xnor U18445 (N_18445,N_17773,N_17057);
nor U18446 (N_18446,N_17491,N_17797);
xnor U18447 (N_18447,N_17307,N_17093);
and U18448 (N_18448,N_17844,N_17588);
nor U18449 (N_18449,N_17952,N_17854);
or U18450 (N_18450,N_17435,N_17075);
xor U18451 (N_18451,N_17227,N_17760);
and U18452 (N_18452,N_17381,N_17042);
and U18453 (N_18453,N_17390,N_17200);
nand U18454 (N_18454,N_17286,N_17000);
and U18455 (N_18455,N_17659,N_17590);
nand U18456 (N_18456,N_17722,N_17260);
xor U18457 (N_18457,N_17318,N_17700);
xor U18458 (N_18458,N_17789,N_17416);
or U18459 (N_18459,N_17849,N_17152);
and U18460 (N_18460,N_17212,N_17277);
nor U18461 (N_18461,N_17263,N_17861);
nor U18462 (N_18462,N_17131,N_17803);
nand U18463 (N_18463,N_17940,N_17182);
and U18464 (N_18464,N_17779,N_17572);
nand U18465 (N_18465,N_17188,N_17551);
and U18466 (N_18466,N_17351,N_17439);
or U18467 (N_18467,N_17702,N_17494);
and U18468 (N_18468,N_17199,N_17929);
and U18469 (N_18469,N_17824,N_17669);
nor U18470 (N_18470,N_17774,N_17095);
or U18471 (N_18471,N_17024,N_17214);
and U18472 (N_18472,N_17236,N_17047);
nor U18473 (N_18473,N_17457,N_17994);
xor U18474 (N_18474,N_17289,N_17299);
xnor U18475 (N_18475,N_17961,N_17710);
nand U18476 (N_18476,N_17845,N_17984);
nor U18477 (N_18477,N_17239,N_17511);
nor U18478 (N_18478,N_17969,N_17096);
nor U18479 (N_18479,N_17542,N_17201);
nand U18480 (N_18480,N_17740,N_17276);
nand U18481 (N_18481,N_17767,N_17721);
and U18482 (N_18482,N_17396,N_17951);
or U18483 (N_18483,N_17628,N_17615);
or U18484 (N_18484,N_17967,N_17038);
nor U18485 (N_18485,N_17544,N_17102);
or U18486 (N_18486,N_17856,N_17818);
nor U18487 (N_18487,N_17033,N_17781);
nor U18488 (N_18488,N_17250,N_17021);
nand U18489 (N_18489,N_17043,N_17676);
nand U18490 (N_18490,N_17234,N_17346);
nand U18491 (N_18491,N_17181,N_17360);
xnor U18492 (N_18492,N_17143,N_17468);
and U18493 (N_18493,N_17211,N_17240);
or U18494 (N_18494,N_17397,N_17825);
and U18495 (N_18495,N_17411,N_17554);
or U18496 (N_18496,N_17870,N_17684);
and U18497 (N_18497,N_17847,N_17704);
and U18498 (N_18498,N_17296,N_17574);
nor U18499 (N_18499,N_17159,N_17815);
or U18500 (N_18500,N_17279,N_17659);
and U18501 (N_18501,N_17857,N_17445);
nand U18502 (N_18502,N_17297,N_17883);
nand U18503 (N_18503,N_17879,N_17488);
nand U18504 (N_18504,N_17311,N_17117);
or U18505 (N_18505,N_17719,N_17187);
and U18506 (N_18506,N_17023,N_17529);
xor U18507 (N_18507,N_17049,N_17609);
nor U18508 (N_18508,N_17760,N_17384);
and U18509 (N_18509,N_17885,N_17580);
nor U18510 (N_18510,N_17770,N_17859);
nor U18511 (N_18511,N_17401,N_17691);
nand U18512 (N_18512,N_17193,N_17153);
and U18513 (N_18513,N_17624,N_17424);
and U18514 (N_18514,N_17261,N_17318);
or U18515 (N_18515,N_17653,N_17595);
or U18516 (N_18516,N_17837,N_17534);
nor U18517 (N_18517,N_17178,N_17880);
or U18518 (N_18518,N_17711,N_17978);
xnor U18519 (N_18519,N_17922,N_17237);
or U18520 (N_18520,N_17635,N_17101);
xor U18521 (N_18521,N_17272,N_17440);
xor U18522 (N_18522,N_17983,N_17788);
nor U18523 (N_18523,N_17245,N_17589);
or U18524 (N_18524,N_17997,N_17731);
or U18525 (N_18525,N_17462,N_17994);
xor U18526 (N_18526,N_17030,N_17565);
nand U18527 (N_18527,N_17319,N_17035);
xnor U18528 (N_18528,N_17330,N_17631);
xor U18529 (N_18529,N_17143,N_17356);
and U18530 (N_18530,N_17417,N_17819);
xor U18531 (N_18531,N_17284,N_17509);
nand U18532 (N_18532,N_17461,N_17294);
and U18533 (N_18533,N_17792,N_17140);
nand U18534 (N_18534,N_17405,N_17082);
or U18535 (N_18535,N_17786,N_17046);
or U18536 (N_18536,N_17432,N_17556);
nand U18537 (N_18537,N_17150,N_17121);
and U18538 (N_18538,N_17954,N_17738);
or U18539 (N_18539,N_17341,N_17938);
nor U18540 (N_18540,N_17356,N_17124);
and U18541 (N_18541,N_17289,N_17513);
nor U18542 (N_18542,N_17268,N_17530);
or U18543 (N_18543,N_17106,N_17594);
or U18544 (N_18544,N_17743,N_17953);
nor U18545 (N_18545,N_17265,N_17262);
xnor U18546 (N_18546,N_17086,N_17783);
or U18547 (N_18547,N_17125,N_17067);
xor U18548 (N_18548,N_17504,N_17319);
and U18549 (N_18549,N_17771,N_17416);
and U18550 (N_18550,N_17964,N_17034);
nor U18551 (N_18551,N_17217,N_17208);
nand U18552 (N_18552,N_17104,N_17637);
xnor U18553 (N_18553,N_17249,N_17468);
and U18554 (N_18554,N_17482,N_17648);
nand U18555 (N_18555,N_17837,N_17110);
nand U18556 (N_18556,N_17838,N_17217);
xnor U18557 (N_18557,N_17552,N_17783);
nor U18558 (N_18558,N_17542,N_17285);
or U18559 (N_18559,N_17185,N_17231);
or U18560 (N_18560,N_17418,N_17410);
nand U18561 (N_18561,N_17530,N_17442);
xnor U18562 (N_18562,N_17114,N_17673);
xor U18563 (N_18563,N_17381,N_17096);
xor U18564 (N_18564,N_17304,N_17536);
and U18565 (N_18565,N_17900,N_17867);
nor U18566 (N_18566,N_17310,N_17327);
and U18567 (N_18567,N_17791,N_17630);
xor U18568 (N_18568,N_17381,N_17447);
nand U18569 (N_18569,N_17151,N_17374);
nand U18570 (N_18570,N_17315,N_17548);
nor U18571 (N_18571,N_17341,N_17569);
xor U18572 (N_18572,N_17476,N_17338);
nor U18573 (N_18573,N_17248,N_17672);
nor U18574 (N_18574,N_17265,N_17543);
and U18575 (N_18575,N_17328,N_17226);
nor U18576 (N_18576,N_17043,N_17552);
or U18577 (N_18577,N_17461,N_17449);
nand U18578 (N_18578,N_17463,N_17019);
xnor U18579 (N_18579,N_17709,N_17376);
nand U18580 (N_18580,N_17358,N_17656);
and U18581 (N_18581,N_17444,N_17432);
nand U18582 (N_18582,N_17059,N_17762);
or U18583 (N_18583,N_17825,N_17207);
and U18584 (N_18584,N_17849,N_17202);
xor U18585 (N_18585,N_17138,N_17131);
nand U18586 (N_18586,N_17314,N_17565);
nand U18587 (N_18587,N_17594,N_17993);
and U18588 (N_18588,N_17288,N_17383);
nor U18589 (N_18589,N_17012,N_17435);
and U18590 (N_18590,N_17093,N_17168);
and U18591 (N_18591,N_17313,N_17927);
or U18592 (N_18592,N_17170,N_17050);
nand U18593 (N_18593,N_17426,N_17427);
and U18594 (N_18594,N_17080,N_17411);
or U18595 (N_18595,N_17589,N_17407);
xor U18596 (N_18596,N_17767,N_17193);
nor U18597 (N_18597,N_17091,N_17149);
and U18598 (N_18598,N_17826,N_17865);
or U18599 (N_18599,N_17868,N_17823);
nor U18600 (N_18600,N_17089,N_17980);
and U18601 (N_18601,N_17047,N_17423);
or U18602 (N_18602,N_17349,N_17466);
nor U18603 (N_18603,N_17594,N_17373);
xor U18604 (N_18604,N_17632,N_17218);
and U18605 (N_18605,N_17674,N_17560);
and U18606 (N_18606,N_17084,N_17469);
nor U18607 (N_18607,N_17126,N_17003);
nor U18608 (N_18608,N_17039,N_17452);
and U18609 (N_18609,N_17626,N_17211);
xnor U18610 (N_18610,N_17152,N_17494);
xnor U18611 (N_18611,N_17536,N_17028);
and U18612 (N_18612,N_17655,N_17765);
or U18613 (N_18613,N_17812,N_17979);
nor U18614 (N_18614,N_17684,N_17934);
or U18615 (N_18615,N_17218,N_17020);
xor U18616 (N_18616,N_17926,N_17531);
nand U18617 (N_18617,N_17023,N_17826);
nor U18618 (N_18618,N_17610,N_17945);
or U18619 (N_18619,N_17883,N_17675);
nor U18620 (N_18620,N_17662,N_17326);
xnor U18621 (N_18621,N_17131,N_17712);
or U18622 (N_18622,N_17392,N_17271);
nor U18623 (N_18623,N_17477,N_17912);
nand U18624 (N_18624,N_17324,N_17338);
xnor U18625 (N_18625,N_17384,N_17848);
and U18626 (N_18626,N_17375,N_17919);
and U18627 (N_18627,N_17011,N_17652);
xnor U18628 (N_18628,N_17509,N_17040);
and U18629 (N_18629,N_17873,N_17109);
xnor U18630 (N_18630,N_17010,N_17158);
and U18631 (N_18631,N_17167,N_17513);
and U18632 (N_18632,N_17145,N_17438);
nand U18633 (N_18633,N_17436,N_17360);
nand U18634 (N_18634,N_17011,N_17409);
xor U18635 (N_18635,N_17232,N_17010);
nand U18636 (N_18636,N_17176,N_17808);
or U18637 (N_18637,N_17731,N_17725);
or U18638 (N_18638,N_17800,N_17738);
xnor U18639 (N_18639,N_17244,N_17264);
nor U18640 (N_18640,N_17512,N_17483);
nor U18641 (N_18641,N_17598,N_17249);
and U18642 (N_18642,N_17084,N_17535);
or U18643 (N_18643,N_17799,N_17838);
and U18644 (N_18644,N_17012,N_17771);
or U18645 (N_18645,N_17370,N_17974);
nor U18646 (N_18646,N_17515,N_17652);
nand U18647 (N_18647,N_17592,N_17978);
or U18648 (N_18648,N_17264,N_17304);
or U18649 (N_18649,N_17972,N_17917);
xor U18650 (N_18650,N_17785,N_17302);
nor U18651 (N_18651,N_17723,N_17519);
nor U18652 (N_18652,N_17045,N_17334);
xor U18653 (N_18653,N_17043,N_17594);
nor U18654 (N_18654,N_17505,N_17264);
nand U18655 (N_18655,N_17865,N_17885);
nor U18656 (N_18656,N_17536,N_17544);
and U18657 (N_18657,N_17816,N_17444);
xor U18658 (N_18658,N_17823,N_17118);
nand U18659 (N_18659,N_17437,N_17808);
nor U18660 (N_18660,N_17153,N_17885);
nand U18661 (N_18661,N_17663,N_17673);
nand U18662 (N_18662,N_17433,N_17302);
or U18663 (N_18663,N_17620,N_17734);
or U18664 (N_18664,N_17140,N_17766);
nor U18665 (N_18665,N_17764,N_17105);
nor U18666 (N_18666,N_17342,N_17795);
xor U18667 (N_18667,N_17883,N_17092);
and U18668 (N_18668,N_17106,N_17779);
nor U18669 (N_18669,N_17518,N_17656);
or U18670 (N_18670,N_17832,N_17666);
and U18671 (N_18671,N_17405,N_17257);
nor U18672 (N_18672,N_17046,N_17983);
xor U18673 (N_18673,N_17458,N_17175);
or U18674 (N_18674,N_17398,N_17872);
and U18675 (N_18675,N_17484,N_17726);
xnor U18676 (N_18676,N_17389,N_17601);
or U18677 (N_18677,N_17765,N_17368);
nand U18678 (N_18678,N_17781,N_17388);
or U18679 (N_18679,N_17817,N_17568);
nor U18680 (N_18680,N_17610,N_17584);
xnor U18681 (N_18681,N_17675,N_17713);
xnor U18682 (N_18682,N_17895,N_17370);
xnor U18683 (N_18683,N_17052,N_17937);
xor U18684 (N_18684,N_17043,N_17182);
or U18685 (N_18685,N_17055,N_17166);
or U18686 (N_18686,N_17390,N_17284);
xnor U18687 (N_18687,N_17385,N_17841);
and U18688 (N_18688,N_17291,N_17890);
nor U18689 (N_18689,N_17576,N_17014);
nand U18690 (N_18690,N_17633,N_17826);
nor U18691 (N_18691,N_17956,N_17734);
and U18692 (N_18692,N_17093,N_17808);
or U18693 (N_18693,N_17611,N_17769);
and U18694 (N_18694,N_17000,N_17711);
or U18695 (N_18695,N_17086,N_17536);
nor U18696 (N_18696,N_17500,N_17751);
nand U18697 (N_18697,N_17720,N_17853);
nor U18698 (N_18698,N_17807,N_17189);
xnor U18699 (N_18699,N_17900,N_17866);
nand U18700 (N_18700,N_17363,N_17977);
or U18701 (N_18701,N_17957,N_17790);
or U18702 (N_18702,N_17797,N_17302);
nor U18703 (N_18703,N_17774,N_17236);
nor U18704 (N_18704,N_17843,N_17826);
nor U18705 (N_18705,N_17038,N_17373);
xor U18706 (N_18706,N_17875,N_17159);
nor U18707 (N_18707,N_17033,N_17900);
nor U18708 (N_18708,N_17808,N_17301);
nor U18709 (N_18709,N_17117,N_17977);
xor U18710 (N_18710,N_17844,N_17404);
nand U18711 (N_18711,N_17865,N_17469);
xnor U18712 (N_18712,N_17015,N_17056);
or U18713 (N_18713,N_17028,N_17167);
and U18714 (N_18714,N_17416,N_17930);
nor U18715 (N_18715,N_17152,N_17964);
nand U18716 (N_18716,N_17406,N_17883);
xor U18717 (N_18717,N_17745,N_17567);
and U18718 (N_18718,N_17309,N_17025);
xor U18719 (N_18719,N_17765,N_17557);
nand U18720 (N_18720,N_17431,N_17951);
xor U18721 (N_18721,N_17759,N_17637);
or U18722 (N_18722,N_17718,N_17485);
or U18723 (N_18723,N_17611,N_17122);
nor U18724 (N_18724,N_17954,N_17191);
and U18725 (N_18725,N_17283,N_17033);
and U18726 (N_18726,N_17595,N_17518);
and U18727 (N_18727,N_17454,N_17746);
or U18728 (N_18728,N_17259,N_17059);
xor U18729 (N_18729,N_17720,N_17029);
and U18730 (N_18730,N_17225,N_17707);
nand U18731 (N_18731,N_17363,N_17022);
or U18732 (N_18732,N_17429,N_17519);
nor U18733 (N_18733,N_17089,N_17022);
nor U18734 (N_18734,N_17414,N_17444);
and U18735 (N_18735,N_17368,N_17879);
nor U18736 (N_18736,N_17847,N_17021);
and U18737 (N_18737,N_17922,N_17643);
nor U18738 (N_18738,N_17700,N_17782);
xnor U18739 (N_18739,N_17914,N_17202);
xnor U18740 (N_18740,N_17563,N_17829);
and U18741 (N_18741,N_17520,N_17373);
or U18742 (N_18742,N_17071,N_17333);
and U18743 (N_18743,N_17841,N_17623);
or U18744 (N_18744,N_17090,N_17965);
nor U18745 (N_18745,N_17798,N_17808);
nor U18746 (N_18746,N_17528,N_17690);
nor U18747 (N_18747,N_17491,N_17566);
and U18748 (N_18748,N_17194,N_17433);
nor U18749 (N_18749,N_17282,N_17750);
xor U18750 (N_18750,N_17411,N_17565);
nand U18751 (N_18751,N_17100,N_17439);
xnor U18752 (N_18752,N_17002,N_17402);
nand U18753 (N_18753,N_17987,N_17669);
nor U18754 (N_18754,N_17060,N_17366);
xor U18755 (N_18755,N_17827,N_17134);
xnor U18756 (N_18756,N_17099,N_17499);
nor U18757 (N_18757,N_17512,N_17830);
or U18758 (N_18758,N_17747,N_17896);
and U18759 (N_18759,N_17890,N_17047);
xnor U18760 (N_18760,N_17743,N_17049);
xor U18761 (N_18761,N_17223,N_17504);
nor U18762 (N_18762,N_17151,N_17263);
nor U18763 (N_18763,N_17140,N_17859);
xnor U18764 (N_18764,N_17729,N_17404);
xnor U18765 (N_18765,N_17323,N_17482);
nor U18766 (N_18766,N_17230,N_17805);
xnor U18767 (N_18767,N_17191,N_17147);
or U18768 (N_18768,N_17792,N_17689);
and U18769 (N_18769,N_17029,N_17503);
xor U18770 (N_18770,N_17707,N_17574);
or U18771 (N_18771,N_17292,N_17683);
xor U18772 (N_18772,N_17430,N_17186);
nor U18773 (N_18773,N_17443,N_17860);
xor U18774 (N_18774,N_17087,N_17264);
xor U18775 (N_18775,N_17419,N_17209);
nand U18776 (N_18776,N_17249,N_17402);
nor U18777 (N_18777,N_17092,N_17426);
and U18778 (N_18778,N_17760,N_17592);
xor U18779 (N_18779,N_17251,N_17049);
nor U18780 (N_18780,N_17626,N_17614);
and U18781 (N_18781,N_17840,N_17675);
nand U18782 (N_18782,N_17236,N_17308);
nand U18783 (N_18783,N_17416,N_17629);
nand U18784 (N_18784,N_17731,N_17374);
xnor U18785 (N_18785,N_17767,N_17879);
and U18786 (N_18786,N_17319,N_17071);
xor U18787 (N_18787,N_17852,N_17989);
and U18788 (N_18788,N_17878,N_17641);
nor U18789 (N_18789,N_17938,N_17377);
and U18790 (N_18790,N_17826,N_17100);
or U18791 (N_18791,N_17492,N_17772);
xnor U18792 (N_18792,N_17162,N_17600);
or U18793 (N_18793,N_17670,N_17693);
or U18794 (N_18794,N_17973,N_17924);
and U18795 (N_18795,N_17465,N_17718);
and U18796 (N_18796,N_17014,N_17343);
nand U18797 (N_18797,N_17577,N_17861);
or U18798 (N_18798,N_17945,N_17293);
nand U18799 (N_18799,N_17204,N_17255);
nand U18800 (N_18800,N_17774,N_17607);
and U18801 (N_18801,N_17841,N_17918);
nand U18802 (N_18802,N_17526,N_17933);
nand U18803 (N_18803,N_17077,N_17026);
xor U18804 (N_18804,N_17361,N_17403);
nand U18805 (N_18805,N_17124,N_17010);
nand U18806 (N_18806,N_17595,N_17983);
or U18807 (N_18807,N_17282,N_17071);
nand U18808 (N_18808,N_17154,N_17422);
nand U18809 (N_18809,N_17653,N_17134);
and U18810 (N_18810,N_17684,N_17002);
nor U18811 (N_18811,N_17982,N_17146);
and U18812 (N_18812,N_17411,N_17665);
nor U18813 (N_18813,N_17981,N_17033);
xnor U18814 (N_18814,N_17817,N_17793);
and U18815 (N_18815,N_17957,N_17509);
or U18816 (N_18816,N_17980,N_17177);
xnor U18817 (N_18817,N_17485,N_17092);
nor U18818 (N_18818,N_17440,N_17289);
nor U18819 (N_18819,N_17463,N_17450);
or U18820 (N_18820,N_17822,N_17241);
and U18821 (N_18821,N_17011,N_17884);
nand U18822 (N_18822,N_17766,N_17098);
nand U18823 (N_18823,N_17501,N_17951);
nor U18824 (N_18824,N_17689,N_17592);
nand U18825 (N_18825,N_17640,N_17635);
or U18826 (N_18826,N_17257,N_17324);
nand U18827 (N_18827,N_17687,N_17668);
nor U18828 (N_18828,N_17971,N_17248);
nor U18829 (N_18829,N_17932,N_17029);
nand U18830 (N_18830,N_17807,N_17397);
xor U18831 (N_18831,N_17415,N_17875);
or U18832 (N_18832,N_17625,N_17772);
nor U18833 (N_18833,N_17565,N_17371);
nand U18834 (N_18834,N_17860,N_17484);
xnor U18835 (N_18835,N_17156,N_17854);
and U18836 (N_18836,N_17874,N_17184);
or U18837 (N_18837,N_17673,N_17124);
nand U18838 (N_18838,N_17033,N_17560);
and U18839 (N_18839,N_17601,N_17772);
and U18840 (N_18840,N_17639,N_17432);
nor U18841 (N_18841,N_17361,N_17998);
or U18842 (N_18842,N_17430,N_17676);
nor U18843 (N_18843,N_17595,N_17523);
nand U18844 (N_18844,N_17583,N_17186);
or U18845 (N_18845,N_17568,N_17407);
or U18846 (N_18846,N_17819,N_17788);
or U18847 (N_18847,N_17882,N_17556);
and U18848 (N_18848,N_17403,N_17385);
xor U18849 (N_18849,N_17198,N_17466);
nor U18850 (N_18850,N_17304,N_17986);
and U18851 (N_18851,N_17087,N_17361);
xor U18852 (N_18852,N_17909,N_17574);
nor U18853 (N_18853,N_17380,N_17882);
and U18854 (N_18854,N_17586,N_17010);
or U18855 (N_18855,N_17181,N_17517);
and U18856 (N_18856,N_17882,N_17376);
or U18857 (N_18857,N_17513,N_17895);
xnor U18858 (N_18858,N_17007,N_17436);
nand U18859 (N_18859,N_17155,N_17438);
xor U18860 (N_18860,N_17921,N_17973);
or U18861 (N_18861,N_17246,N_17789);
and U18862 (N_18862,N_17303,N_17154);
and U18863 (N_18863,N_17033,N_17408);
and U18864 (N_18864,N_17958,N_17718);
xor U18865 (N_18865,N_17385,N_17098);
nor U18866 (N_18866,N_17188,N_17928);
and U18867 (N_18867,N_17078,N_17749);
xnor U18868 (N_18868,N_17740,N_17494);
nor U18869 (N_18869,N_17765,N_17555);
or U18870 (N_18870,N_17379,N_17817);
nand U18871 (N_18871,N_17919,N_17981);
nand U18872 (N_18872,N_17608,N_17045);
xnor U18873 (N_18873,N_17082,N_17890);
and U18874 (N_18874,N_17045,N_17349);
xnor U18875 (N_18875,N_17431,N_17259);
nor U18876 (N_18876,N_17366,N_17208);
or U18877 (N_18877,N_17196,N_17778);
or U18878 (N_18878,N_17572,N_17818);
nor U18879 (N_18879,N_17871,N_17439);
or U18880 (N_18880,N_17623,N_17555);
nand U18881 (N_18881,N_17662,N_17267);
xor U18882 (N_18882,N_17985,N_17065);
nor U18883 (N_18883,N_17711,N_17912);
nand U18884 (N_18884,N_17963,N_17452);
nand U18885 (N_18885,N_17317,N_17817);
and U18886 (N_18886,N_17137,N_17792);
or U18887 (N_18887,N_17606,N_17007);
xnor U18888 (N_18888,N_17936,N_17217);
and U18889 (N_18889,N_17687,N_17281);
and U18890 (N_18890,N_17951,N_17201);
and U18891 (N_18891,N_17338,N_17924);
nor U18892 (N_18892,N_17269,N_17434);
or U18893 (N_18893,N_17685,N_17758);
nand U18894 (N_18894,N_17789,N_17908);
nand U18895 (N_18895,N_17404,N_17750);
or U18896 (N_18896,N_17087,N_17759);
nor U18897 (N_18897,N_17342,N_17080);
or U18898 (N_18898,N_17954,N_17830);
nor U18899 (N_18899,N_17703,N_17776);
or U18900 (N_18900,N_17323,N_17185);
nor U18901 (N_18901,N_17981,N_17386);
nand U18902 (N_18902,N_17596,N_17842);
and U18903 (N_18903,N_17250,N_17024);
and U18904 (N_18904,N_17638,N_17974);
nor U18905 (N_18905,N_17127,N_17401);
nand U18906 (N_18906,N_17796,N_17057);
and U18907 (N_18907,N_17791,N_17261);
nand U18908 (N_18908,N_17858,N_17259);
nor U18909 (N_18909,N_17181,N_17578);
and U18910 (N_18910,N_17096,N_17729);
xor U18911 (N_18911,N_17077,N_17243);
nor U18912 (N_18912,N_17988,N_17520);
nor U18913 (N_18913,N_17168,N_17177);
nor U18914 (N_18914,N_17698,N_17225);
nor U18915 (N_18915,N_17255,N_17338);
nand U18916 (N_18916,N_17748,N_17742);
nor U18917 (N_18917,N_17746,N_17945);
nor U18918 (N_18918,N_17649,N_17418);
nand U18919 (N_18919,N_17638,N_17721);
and U18920 (N_18920,N_17822,N_17817);
or U18921 (N_18921,N_17841,N_17624);
nand U18922 (N_18922,N_17206,N_17076);
nor U18923 (N_18923,N_17595,N_17577);
xnor U18924 (N_18924,N_17271,N_17267);
nor U18925 (N_18925,N_17203,N_17629);
xor U18926 (N_18926,N_17055,N_17709);
and U18927 (N_18927,N_17801,N_17104);
and U18928 (N_18928,N_17472,N_17990);
nand U18929 (N_18929,N_17875,N_17145);
and U18930 (N_18930,N_17631,N_17043);
nand U18931 (N_18931,N_17618,N_17483);
or U18932 (N_18932,N_17347,N_17440);
or U18933 (N_18933,N_17936,N_17384);
nor U18934 (N_18934,N_17215,N_17596);
nor U18935 (N_18935,N_17839,N_17834);
and U18936 (N_18936,N_17922,N_17809);
xor U18937 (N_18937,N_17041,N_17192);
nand U18938 (N_18938,N_17958,N_17158);
xnor U18939 (N_18939,N_17769,N_17853);
or U18940 (N_18940,N_17882,N_17363);
xnor U18941 (N_18941,N_17128,N_17451);
nor U18942 (N_18942,N_17116,N_17974);
xor U18943 (N_18943,N_17015,N_17048);
nand U18944 (N_18944,N_17122,N_17084);
or U18945 (N_18945,N_17933,N_17861);
xor U18946 (N_18946,N_17811,N_17390);
nand U18947 (N_18947,N_17457,N_17410);
nand U18948 (N_18948,N_17833,N_17616);
or U18949 (N_18949,N_17291,N_17836);
or U18950 (N_18950,N_17121,N_17378);
nor U18951 (N_18951,N_17898,N_17785);
xnor U18952 (N_18952,N_17061,N_17293);
nor U18953 (N_18953,N_17592,N_17890);
xor U18954 (N_18954,N_17543,N_17633);
xor U18955 (N_18955,N_17565,N_17610);
nor U18956 (N_18956,N_17865,N_17980);
xor U18957 (N_18957,N_17227,N_17572);
and U18958 (N_18958,N_17698,N_17486);
or U18959 (N_18959,N_17763,N_17523);
nand U18960 (N_18960,N_17476,N_17727);
nor U18961 (N_18961,N_17511,N_17969);
nor U18962 (N_18962,N_17963,N_17477);
nand U18963 (N_18963,N_17582,N_17873);
or U18964 (N_18964,N_17040,N_17496);
or U18965 (N_18965,N_17286,N_17829);
nand U18966 (N_18966,N_17509,N_17666);
xnor U18967 (N_18967,N_17009,N_17663);
and U18968 (N_18968,N_17992,N_17195);
nand U18969 (N_18969,N_17249,N_17884);
or U18970 (N_18970,N_17920,N_17991);
nor U18971 (N_18971,N_17286,N_17207);
xor U18972 (N_18972,N_17969,N_17824);
or U18973 (N_18973,N_17237,N_17490);
nand U18974 (N_18974,N_17564,N_17145);
or U18975 (N_18975,N_17664,N_17370);
nor U18976 (N_18976,N_17151,N_17883);
xnor U18977 (N_18977,N_17259,N_17609);
and U18978 (N_18978,N_17283,N_17237);
or U18979 (N_18979,N_17956,N_17683);
and U18980 (N_18980,N_17752,N_17935);
nor U18981 (N_18981,N_17112,N_17553);
xnor U18982 (N_18982,N_17115,N_17271);
xnor U18983 (N_18983,N_17834,N_17901);
xor U18984 (N_18984,N_17124,N_17948);
nand U18985 (N_18985,N_17776,N_17749);
xnor U18986 (N_18986,N_17385,N_17775);
or U18987 (N_18987,N_17029,N_17656);
nor U18988 (N_18988,N_17999,N_17776);
xor U18989 (N_18989,N_17746,N_17270);
nor U18990 (N_18990,N_17936,N_17913);
xor U18991 (N_18991,N_17024,N_17442);
or U18992 (N_18992,N_17383,N_17065);
or U18993 (N_18993,N_17198,N_17452);
and U18994 (N_18994,N_17586,N_17866);
nor U18995 (N_18995,N_17488,N_17271);
or U18996 (N_18996,N_17271,N_17419);
or U18997 (N_18997,N_17341,N_17078);
xor U18998 (N_18998,N_17030,N_17739);
nand U18999 (N_18999,N_17344,N_17646);
nand U19000 (N_19000,N_18299,N_18259);
and U19001 (N_19001,N_18943,N_18755);
and U19002 (N_19002,N_18032,N_18751);
and U19003 (N_19003,N_18489,N_18798);
xor U19004 (N_19004,N_18612,N_18266);
nand U19005 (N_19005,N_18724,N_18823);
nor U19006 (N_19006,N_18397,N_18687);
nor U19007 (N_19007,N_18513,N_18799);
and U19008 (N_19008,N_18664,N_18298);
and U19009 (N_19009,N_18231,N_18522);
and U19010 (N_19010,N_18191,N_18353);
nand U19011 (N_19011,N_18783,N_18909);
xor U19012 (N_19012,N_18127,N_18817);
nand U19013 (N_19013,N_18312,N_18589);
nand U19014 (N_19014,N_18990,N_18016);
or U19015 (N_19015,N_18761,N_18218);
or U19016 (N_19016,N_18381,N_18126);
or U19017 (N_19017,N_18083,N_18949);
and U19018 (N_19018,N_18486,N_18746);
or U19019 (N_19019,N_18902,N_18694);
xnor U19020 (N_19020,N_18084,N_18323);
or U19021 (N_19021,N_18560,N_18056);
and U19022 (N_19022,N_18713,N_18403);
or U19023 (N_19023,N_18594,N_18374);
nand U19024 (N_19024,N_18964,N_18770);
xnor U19025 (N_19025,N_18287,N_18654);
or U19026 (N_19026,N_18430,N_18454);
xor U19027 (N_19027,N_18558,N_18520);
xnor U19028 (N_19028,N_18966,N_18566);
xnor U19029 (N_19029,N_18002,N_18448);
or U19030 (N_19030,N_18340,N_18094);
nor U19031 (N_19031,N_18553,N_18624);
nand U19032 (N_19032,N_18601,N_18791);
nand U19033 (N_19033,N_18866,N_18112);
and U19034 (N_19034,N_18268,N_18618);
nor U19035 (N_19035,N_18756,N_18590);
and U19036 (N_19036,N_18762,N_18147);
or U19037 (N_19037,N_18436,N_18473);
xnor U19038 (N_19038,N_18113,N_18030);
or U19039 (N_19039,N_18675,N_18765);
nand U19040 (N_19040,N_18580,N_18081);
or U19041 (N_19041,N_18103,N_18398);
nand U19042 (N_19042,N_18456,N_18254);
or U19043 (N_19043,N_18918,N_18673);
nor U19044 (N_19044,N_18243,N_18018);
and U19045 (N_19045,N_18452,N_18500);
and U19046 (N_19046,N_18386,N_18945);
nand U19047 (N_19047,N_18021,N_18371);
nand U19048 (N_19048,N_18435,N_18764);
nand U19049 (N_19049,N_18773,N_18038);
xor U19050 (N_19050,N_18503,N_18582);
nor U19051 (N_19051,N_18459,N_18696);
or U19052 (N_19052,N_18297,N_18301);
or U19053 (N_19053,N_18058,N_18959);
and U19054 (N_19054,N_18588,N_18311);
xnor U19055 (N_19055,N_18467,N_18977);
and U19056 (N_19056,N_18292,N_18651);
xor U19057 (N_19057,N_18236,N_18046);
nor U19058 (N_19058,N_18421,N_18223);
or U19059 (N_19059,N_18031,N_18986);
and U19060 (N_19060,N_18289,N_18458);
nand U19061 (N_19061,N_18778,N_18176);
xor U19062 (N_19062,N_18365,N_18822);
nand U19063 (N_19063,N_18348,N_18750);
nor U19064 (N_19064,N_18009,N_18608);
nand U19065 (N_19065,N_18174,N_18416);
xnor U19066 (N_19066,N_18239,N_18211);
or U19067 (N_19067,N_18728,N_18954);
and U19068 (N_19068,N_18335,N_18437);
nor U19069 (N_19069,N_18542,N_18793);
xnor U19070 (N_19070,N_18146,N_18166);
and U19071 (N_19071,N_18149,N_18173);
nor U19072 (N_19072,N_18382,N_18704);
or U19073 (N_19073,N_18116,N_18524);
or U19074 (N_19074,N_18640,N_18702);
nor U19075 (N_19075,N_18646,N_18586);
nor U19076 (N_19076,N_18110,N_18282);
or U19077 (N_19077,N_18787,N_18893);
or U19078 (N_19078,N_18206,N_18306);
and U19079 (N_19079,N_18603,N_18156);
nor U19080 (N_19080,N_18812,N_18376);
nand U19081 (N_19081,N_18622,N_18415);
or U19082 (N_19082,N_18616,N_18923);
nand U19083 (N_19083,N_18499,N_18725);
xnor U19084 (N_19084,N_18737,N_18495);
nor U19085 (N_19085,N_18815,N_18846);
and U19086 (N_19086,N_18853,N_18827);
and U19087 (N_19087,N_18731,N_18802);
xor U19088 (N_19088,N_18875,N_18203);
and U19089 (N_19089,N_18633,N_18248);
or U19090 (N_19090,N_18691,N_18961);
or U19091 (N_19091,N_18001,N_18721);
and U19092 (N_19092,N_18372,N_18670);
nor U19093 (N_19093,N_18479,N_18294);
xnor U19094 (N_19094,N_18035,N_18858);
nor U19095 (N_19095,N_18375,N_18184);
nand U19096 (N_19096,N_18310,N_18327);
nor U19097 (N_19097,N_18790,N_18991);
xnor U19098 (N_19098,N_18530,N_18826);
and U19099 (N_19099,N_18663,N_18965);
nor U19100 (N_19100,N_18881,N_18051);
or U19101 (N_19101,N_18296,N_18552);
or U19102 (N_19102,N_18474,N_18369);
or U19103 (N_19103,N_18220,N_18012);
nor U19104 (N_19104,N_18962,N_18636);
nand U19105 (N_19105,N_18219,N_18641);
or U19106 (N_19106,N_18333,N_18526);
xor U19107 (N_19107,N_18057,N_18272);
nor U19108 (N_19108,N_18786,N_18975);
nand U19109 (N_19109,N_18114,N_18304);
and U19110 (N_19110,N_18736,N_18475);
and U19111 (N_19111,N_18920,N_18477);
and U19112 (N_19112,N_18124,N_18738);
nand U19113 (N_19113,N_18816,N_18532);
nor U19114 (N_19114,N_18652,N_18619);
xor U19115 (N_19115,N_18908,N_18538);
or U19116 (N_19116,N_18614,N_18300);
nor U19117 (N_19117,N_18125,N_18422);
or U19118 (N_19118,N_18133,N_18659);
nor U19119 (N_19119,N_18706,N_18888);
xnor U19120 (N_19120,N_18144,N_18672);
xor U19121 (N_19121,N_18175,N_18722);
and U19122 (N_19122,N_18583,N_18395);
xnor U19123 (N_19123,N_18726,N_18252);
nand U19124 (N_19124,N_18584,N_18662);
or U19125 (N_19125,N_18068,N_18838);
and U19126 (N_19126,N_18941,N_18054);
nand U19127 (N_19127,N_18565,N_18914);
or U19128 (N_19128,N_18278,N_18101);
and U19129 (N_19129,N_18997,N_18181);
nand U19130 (N_19130,N_18086,N_18187);
nor U19131 (N_19131,N_18564,N_18072);
xor U19132 (N_19132,N_18401,N_18285);
nor U19133 (N_19133,N_18082,N_18302);
or U19134 (N_19134,N_18788,N_18984);
and U19135 (N_19135,N_18036,N_18255);
xor U19136 (N_19136,N_18803,N_18411);
nand U19137 (N_19137,N_18154,N_18545);
and U19138 (N_19138,N_18801,N_18992);
nand U19139 (N_19139,N_18698,N_18076);
or U19140 (N_19140,N_18228,N_18221);
xor U19141 (N_19141,N_18469,N_18115);
nand U19142 (N_19142,N_18820,N_18955);
or U19143 (N_19143,N_18025,N_18763);
and U19144 (N_19144,N_18688,N_18198);
or U19145 (N_19145,N_18648,N_18967);
or U19146 (N_19146,N_18158,N_18396);
nor U19147 (N_19147,N_18572,N_18085);
or U19148 (N_19148,N_18892,N_18048);
and U19149 (N_19149,N_18994,N_18981);
xnor U19150 (N_19150,N_18742,N_18050);
xor U19151 (N_19151,N_18857,N_18732);
or U19152 (N_19152,N_18045,N_18825);
or U19153 (N_19153,N_18202,N_18078);
and U19154 (N_19154,N_18719,N_18769);
nand U19155 (N_19155,N_18766,N_18033);
nor U19156 (N_19156,N_18004,N_18693);
or U19157 (N_19157,N_18891,N_18245);
nor U19158 (N_19158,N_18425,N_18399);
nor U19159 (N_19159,N_18919,N_18214);
nand U19160 (N_19160,N_18844,N_18325);
xnor U19161 (N_19161,N_18157,N_18195);
nand U19162 (N_19162,N_18426,N_18490);
nand U19163 (N_19163,N_18972,N_18876);
and U19164 (N_19164,N_18837,N_18217);
xor U19165 (N_19165,N_18208,N_18339);
and U19166 (N_19166,N_18170,N_18808);
or U19167 (N_19167,N_18439,N_18507);
nand U19168 (N_19168,N_18019,N_18433);
xor U19169 (N_19169,N_18451,N_18434);
or U19170 (N_19170,N_18819,N_18143);
xnor U19171 (N_19171,N_18460,N_18098);
or U19172 (N_19172,N_18518,N_18859);
nand U19173 (N_19173,N_18547,N_18227);
or U19174 (N_19174,N_18749,N_18105);
and U19175 (N_19175,N_18406,N_18831);
nor U19176 (N_19176,N_18118,N_18256);
and U19177 (N_19177,N_18833,N_18644);
nand U19178 (N_19178,N_18328,N_18631);
nand U19179 (N_19179,N_18661,N_18655);
xnor U19180 (N_19180,N_18466,N_18167);
nand U19181 (N_19181,N_18043,N_18052);
nor U19182 (N_19182,N_18155,N_18940);
nor U19183 (N_19183,N_18006,N_18079);
nand U19184 (N_19184,N_18315,N_18013);
nor U19185 (N_19185,N_18359,N_18942);
nand U19186 (N_19186,N_18322,N_18948);
and U19187 (N_19187,N_18258,N_18544);
nor U19188 (N_19188,N_18276,N_18805);
nor U19189 (N_19189,N_18226,N_18141);
nor U19190 (N_19190,N_18039,N_18182);
and U19191 (N_19191,N_18017,N_18506);
nor U19192 (N_19192,N_18334,N_18657);
and U19193 (N_19193,N_18213,N_18008);
and U19194 (N_19194,N_18179,N_18476);
and U19195 (N_19195,N_18674,N_18951);
xnor U19196 (N_19196,N_18368,N_18153);
and U19197 (N_19197,N_18678,N_18850);
or U19198 (N_19198,N_18505,N_18090);
xor U19199 (N_19199,N_18634,N_18679);
nor U19200 (N_19200,N_18865,N_18549);
or U19201 (N_19201,N_18165,N_18134);
nor U19202 (N_19202,N_18928,N_18461);
nor U19203 (N_19203,N_18539,N_18864);
or U19204 (N_19204,N_18936,N_18447);
nor U19205 (N_19205,N_18380,N_18117);
or U19206 (N_19206,N_18352,N_18781);
or U19207 (N_19207,N_18595,N_18767);
or U19208 (N_19208,N_18059,N_18625);
nor U19209 (N_19209,N_18491,N_18355);
or U19210 (N_19210,N_18754,N_18324);
nor U19211 (N_19211,N_18349,N_18921);
and U19212 (N_19212,N_18987,N_18326);
nor U19213 (N_19213,N_18024,N_18494);
xor U19214 (N_19214,N_18824,N_18797);
xor U19215 (N_19215,N_18795,N_18207);
nand U19216 (N_19216,N_18164,N_18354);
nand U19217 (N_19217,N_18373,N_18501);
and U19218 (N_19218,N_18630,N_18318);
or U19219 (N_19219,N_18344,N_18370);
nor U19220 (N_19220,N_18834,N_18960);
or U19221 (N_19221,N_18135,N_18502);
xnor U19222 (N_19222,N_18771,N_18671);
xor U19223 (N_19223,N_18201,N_18177);
or U19224 (N_19224,N_18504,N_18172);
nor U19225 (N_19225,N_18600,N_18345);
nand U19226 (N_19226,N_18969,N_18482);
nand U19227 (N_19227,N_18851,N_18700);
and U19228 (N_19228,N_18757,N_18237);
or U19229 (N_19229,N_18944,N_18014);
xor U19230 (N_19230,N_18064,N_18988);
xnor U19231 (N_19231,N_18615,N_18023);
nand U19232 (N_19232,N_18870,N_18468);
and U19233 (N_19233,N_18982,N_18901);
or U19234 (N_19234,N_18896,N_18029);
nand U19235 (N_19235,N_18424,N_18658);
xnor U19236 (N_19236,N_18257,N_18168);
xnor U19237 (N_19237,N_18455,N_18387);
nand U19238 (N_19238,N_18937,N_18493);
and U19239 (N_19239,N_18111,N_18894);
and U19240 (N_19240,N_18515,N_18860);
or U19241 (N_19241,N_18561,N_18250);
or U19242 (N_19242,N_18579,N_18734);
xor U19243 (N_19243,N_18427,N_18604);
nor U19244 (N_19244,N_18958,N_18996);
nand U19245 (N_19245,N_18358,N_18978);
xnor U19246 (N_19246,N_18956,N_18649);
nor U19247 (N_19247,N_18645,N_18899);
or U19248 (N_19248,N_18741,N_18230);
and U19249 (N_19249,N_18449,N_18718);
or U19250 (N_19250,N_18096,N_18613);
or U19251 (N_19251,N_18939,N_18343);
nor U19252 (N_19252,N_18995,N_18492);
and U19253 (N_19253,N_18271,N_18895);
or U19254 (N_19254,N_18209,N_18903);
nor U19255 (N_19255,N_18362,N_18745);
nor U19256 (N_19256,N_18041,N_18137);
nand U19257 (N_19257,N_18022,N_18280);
or U19258 (N_19258,N_18104,N_18440);
nor U19259 (N_19259,N_18238,N_18665);
xor U19260 (N_19260,N_18385,N_18121);
and U19261 (N_19261,N_18015,N_18739);
or U19262 (N_19262,N_18262,N_18119);
xor U19263 (N_19263,N_18980,N_18514);
nor U19264 (N_19264,N_18185,N_18841);
xnor U19265 (N_19265,N_18338,N_18314);
or U19266 (N_19266,N_18383,N_18882);
xor U19267 (N_19267,N_18776,N_18528);
xor U19268 (N_19268,N_18044,N_18308);
nor U19269 (N_19269,N_18316,N_18319);
and U19270 (N_19270,N_18686,N_18329);
xor U19271 (N_19271,N_18963,N_18517);
nor U19272 (N_19272,N_18088,N_18284);
nand U19273 (N_19273,N_18568,N_18171);
xnor U19274 (N_19274,N_18874,N_18419);
xnor U19275 (N_19275,N_18136,N_18178);
xnor U19276 (N_19276,N_18620,N_18818);
xnor U19277 (N_19277,N_18192,N_18389);
and U19278 (N_19278,N_18701,N_18071);
or U19279 (N_19279,N_18905,N_18912);
nand U19280 (N_19280,N_18814,N_18626);
nand U19281 (N_19281,N_18186,N_18950);
xor U19282 (N_19282,N_18091,N_18989);
nand U19283 (N_19283,N_18034,N_18650);
or U19284 (N_19284,N_18346,N_18933);
nor U19285 (N_19285,N_18350,N_18402);
nor U19286 (N_19286,N_18394,N_18683);
or U19287 (N_19287,N_18180,N_18462);
and U19288 (N_19288,N_18132,N_18260);
xnor U19289 (N_19289,N_18692,N_18151);
or U19290 (N_19290,N_18587,N_18813);
nor U19291 (N_19291,N_18360,N_18336);
and U19292 (N_19292,N_18690,N_18444);
or U19293 (N_19293,N_18843,N_18653);
xnor U19294 (N_19294,N_18487,N_18189);
xor U19295 (N_19295,N_18830,N_18593);
nand U19296 (N_19296,N_18069,N_18122);
nor U19297 (N_19297,N_18063,N_18804);
or U19298 (N_19298,N_18077,N_18845);
nor U19299 (N_19299,N_18541,N_18074);
xor U19300 (N_19300,N_18872,N_18796);
nor U19301 (N_19301,N_18277,N_18011);
nand U19302 (N_19302,N_18669,N_18794);
and U19303 (N_19303,N_18481,N_18660);
xnor U19304 (N_19304,N_18829,N_18927);
and U19305 (N_19305,N_18295,N_18720);
and U19306 (N_19306,N_18210,N_18224);
nand U19307 (N_19307,N_18733,N_18414);
nor U19308 (N_19308,N_18540,N_18160);
nor U19309 (N_19309,N_18922,N_18712);
nand U19310 (N_19310,N_18556,N_18723);
nor U19311 (N_19311,N_18635,N_18811);
and U19312 (N_19312,N_18759,N_18525);
and U19313 (N_19313,N_18443,N_18839);
nand U19314 (N_19314,N_18924,N_18357);
nor U19315 (N_19315,N_18596,N_18639);
xor U19316 (N_19316,N_18128,N_18807);
nor U19317 (N_19317,N_18779,N_18607);
and U19318 (N_19318,N_18042,N_18317);
nand U19319 (N_19319,N_18758,N_18247);
or U19320 (N_19320,N_18251,N_18780);
nor U19321 (N_19321,N_18193,N_18511);
or U19322 (N_19322,N_18470,N_18667);
or U19323 (N_19323,N_18800,N_18628);
nor U19324 (N_19324,N_18131,N_18621);
and U19325 (N_19325,N_18777,N_18241);
nor U19326 (N_19326,N_18854,N_18676);
xnor U19327 (N_19327,N_18931,N_18465);
nand U19328 (N_19328,N_18432,N_18785);
and U19329 (N_19329,N_18890,N_18313);
nand U19330 (N_19330,N_18263,N_18848);
and U19331 (N_19331,N_18863,N_18656);
or U19332 (N_19332,N_18431,N_18571);
xnor U19333 (N_19333,N_18407,N_18585);
nor U19334 (N_19334,N_18752,N_18792);
nor U19335 (N_19335,N_18159,N_18567);
and U19336 (N_19336,N_18705,N_18130);
or U19337 (N_19337,N_18410,N_18488);
and U19338 (N_19338,N_18429,N_18789);
nor U19339 (N_19339,N_18569,N_18265);
and U19340 (N_19340,N_18998,N_18708);
nand U19341 (N_19341,N_18573,N_18450);
or U19342 (N_19342,N_18710,N_18087);
nand U19343 (N_19343,N_18000,N_18095);
and U19344 (N_19344,N_18970,N_18772);
nor U19345 (N_19345,N_18108,N_18557);
xnor U19346 (N_19346,N_18760,N_18089);
nand U19347 (N_19347,N_18010,N_18832);
nor U19348 (N_19348,N_18286,N_18536);
xor U19349 (N_19349,N_18379,N_18204);
nand U19350 (N_19350,N_18682,N_18910);
xnor U19351 (N_19351,N_18930,N_18748);
nand U19352 (N_19352,N_18983,N_18264);
nor U19353 (N_19353,N_18123,N_18550);
xor U19354 (N_19354,N_18140,N_18332);
xor U19355 (N_19355,N_18497,N_18246);
or U19356 (N_19356,N_18632,N_18623);
nand U19357 (N_19357,N_18049,N_18856);
nor U19358 (N_19358,N_18129,N_18026);
or U19359 (N_19359,N_18453,N_18152);
nand U19360 (N_19360,N_18485,N_18199);
xor U19361 (N_19361,N_18689,N_18139);
or U19362 (N_19362,N_18885,N_18351);
and U19363 (N_19363,N_18531,N_18161);
or U19364 (N_19364,N_18190,N_18703);
and U19365 (N_19365,N_18979,N_18281);
or U19366 (N_19366,N_18889,N_18364);
and U19367 (N_19367,N_18442,N_18717);
nand U19368 (N_19368,N_18897,N_18535);
xnor U19369 (N_19369,N_18483,N_18099);
and U19370 (N_19370,N_18320,N_18331);
or U19371 (N_19371,N_18784,N_18929);
xnor U19372 (N_19372,N_18602,N_18576);
or U19373 (N_19373,N_18205,N_18559);
and U19374 (N_19374,N_18508,N_18138);
and U19375 (N_19375,N_18575,N_18999);
xnor U19376 (N_19376,N_18020,N_18681);
xor U19377 (N_19377,N_18120,N_18109);
xor U19378 (N_19378,N_18993,N_18642);
and U19379 (N_19379,N_18925,N_18985);
nand U19380 (N_19380,N_18543,N_18408);
or U19381 (N_19381,N_18100,N_18709);
nand U19382 (N_19382,N_18384,N_18598);
or U19383 (N_19383,N_18269,N_18534);
or U19384 (N_19384,N_18347,N_18768);
xor U19385 (N_19385,N_18067,N_18555);
or U19386 (N_19386,N_18685,N_18225);
nor U19387 (N_19387,N_18464,N_18070);
xor U19388 (N_19388,N_18915,N_18968);
nand U19389 (N_19389,N_18877,N_18215);
or U19390 (N_19390,N_18871,N_18445);
and U19391 (N_19391,N_18378,N_18197);
or U19392 (N_19392,N_18926,N_18947);
and U19393 (N_19393,N_18821,N_18546);
and U19394 (N_19394,N_18868,N_18233);
xor U19395 (N_19395,N_18849,N_18194);
nand U19396 (N_19396,N_18869,N_18599);
nor U19397 (N_19397,N_18581,N_18413);
xnor U19398 (N_19398,N_18743,N_18478);
nand U19399 (N_19399,N_18169,N_18911);
nor U19400 (N_19400,N_18341,N_18291);
or U19401 (N_19401,N_18471,N_18684);
xnor U19402 (N_19402,N_18093,N_18303);
nor U19403 (N_19403,N_18847,N_18747);
nand U19404 (N_19404,N_18200,N_18405);
and U19405 (N_19405,N_18973,N_18400);
or U19406 (N_19406,N_18677,N_18570);
and U19407 (N_19407,N_18007,N_18512);
or U19408 (N_19408,N_18412,N_18275);
nor U19409 (N_19409,N_18027,N_18367);
or U19410 (N_19410,N_18420,N_18629);
and U19411 (N_19411,N_18188,N_18509);
nor U19412 (N_19412,N_18609,N_18107);
and U19413 (N_19413,N_18574,N_18836);
xor U19414 (N_19414,N_18235,N_18288);
and U19415 (N_19415,N_18976,N_18971);
or U19416 (N_19416,N_18307,N_18974);
or U19417 (N_19417,N_18073,N_18441);
xnor U19418 (N_19418,N_18907,N_18668);
nor U19419 (N_19419,N_18309,N_18774);
xnor U19420 (N_19420,N_18782,N_18342);
xnor U19421 (N_19421,N_18699,N_18554);
and U19422 (N_19422,N_18055,N_18887);
or U19423 (N_19423,N_18627,N_18716);
or U19424 (N_19424,N_18715,N_18183);
nor U19425 (N_19425,N_18562,N_18253);
nand U19426 (N_19426,N_18080,N_18957);
and U19427 (N_19427,N_18610,N_18953);
nor U19428 (N_19428,N_18938,N_18886);
xnor U19429 (N_19429,N_18906,N_18212);
or U19430 (N_19430,N_18577,N_18409);
nand U19431 (N_19431,N_18643,N_18356);
nor U19432 (N_19432,N_18934,N_18066);
xnor U19433 (N_19433,N_18003,N_18735);
or U19434 (N_19434,N_18521,N_18321);
and U19435 (N_19435,N_18290,N_18878);
and U19436 (N_19436,N_18606,N_18578);
nor U19437 (N_19437,N_18730,N_18862);
nor U19438 (N_19438,N_18196,N_18142);
nand U19439 (N_19439,N_18283,N_18806);
or U19440 (N_19440,N_18463,N_18840);
nand U19441 (N_19441,N_18145,N_18446);
xnor U19442 (N_19442,N_18744,N_18244);
or U19443 (N_19443,N_18711,N_18527);
or U19444 (N_19444,N_18533,N_18842);
xor U19445 (N_19445,N_18714,N_18391);
or U19446 (N_19446,N_18537,N_18232);
xnor U19447 (N_19447,N_18727,N_18516);
nor U19448 (N_19448,N_18740,N_18873);
nand U19449 (N_19449,N_18548,N_18060);
or U19450 (N_19450,N_18330,N_18484);
nor U19451 (N_19451,N_18605,N_18563);
nand U19452 (N_19452,N_18753,N_18075);
or U19453 (N_19453,N_18828,N_18472);
nor U19454 (N_19454,N_18092,N_18065);
nand U19455 (N_19455,N_18273,N_18498);
or U19456 (N_19456,N_18935,N_18880);
nor U19457 (N_19457,N_18597,N_18163);
nor U19458 (N_19458,N_18835,N_18519);
or U19459 (N_19459,N_18611,N_18707);
or U19460 (N_19460,N_18695,N_18249);
xnor U19461 (N_19461,N_18279,N_18270);
and U19462 (N_19462,N_18293,N_18392);
nor U19463 (N_19463,N_18867,N_18393);
nand U19464 (N_19464,N_18457,N_18900);
and U19465 (N_19465,N_18529,N_18377);
and U19466 (N_19466,N_18855,N_18261);
and U19467 (N_19467,N_18390,N_18040);
nand U19468 (N_19468,N_18637,N_18879);
xnor U19469 (N_19469,N_18053,N_18913);
or U19470 (N_19470,N_18062,N_18274);
or U19471 (N_19471,N_18592,N_18697);
or U19472 (N_19472,N_18932,N_18898);
xnor U19473 (N_19473,N_18680,N_18366);
xnor U19474 (N_19474,N_18438,N_18404);
nor U19475 (N_19475,N_18617,N_18666);
and U19476 (N_19476,N_18523,N_18551);
or U19477 (N_19477,N_18423,N_18916);
xnor U19478 (N_19478,N_18240,N_18647);
and U19479 (N_19479,N_18480,N_18884);
nor U19480 (N_19480,N_18005,N_18809);
or U19481 (N_19481,N_18496,N_18150);
nor U19482 (N_19482,N_18234,N_18305);
nor U19483 (N_19483,N_18810,N_18510);
xor U19484 (N_19484,N_18106,N_18097);
or U19485 (N_19485,N_18363,N_18428);
nand U19486 (N_19486,N_18729,N_18102);
and U19487 (N_19487,N_18361,N_18242);
or U19488 (N_19488,N_18028,N_18037);
or U19489 (N_19489,N_18229,N_18591);
and U19490 (N_19490,N_18946,N_18418);
nand U19491 (N_19491,N_18883,N_18638);
nor U19492 (N_19492,N_18267,N_18162);
and U19493 (N_19493,N_18417,N_18047);
and U19494 (N_19494,N_18222,N_18388);
xnor U19495 (N_19495,N_18148,N_18852);
nor U19496 (N_19496,N_18904,N_18775);
nand U19497 (N_19497,N_18061,N_18337);
xor U19498 (N_19498,N_18952,N_18861);
nor U19499 (N_19499,N_18917,N_18216);
nor U19500 (N_19500,N_18138,N_18769);
and U19501 (N_19501,N_18960,N_18094);
nand U19502 (N_19502,N_18688,N_18537);
xnor U19503 (N_19503,N_18751,N_18685);
or U19504 (N_19504,N_18493,N_18957);
nor U19505 (N_19505,N_18667,N_18493);
nand U19506 (N_19506,N_18075,N_18403);
or U19507 (N_19507,N_18244,N_18373);
and U19508 (N_19508,N_18024,N_18571);
and U19509 (N_19509,N_18697,N_18465);
and U19510 (N_19510,N_18669,N_18462);
or U19511 (N_19511,N_18901,N_18232);
and U19512 (N_19512,N_18219,N_18241);
xor U19513 (N_19513,N_18292,N_18843);
xor U19514 (N_19514,N_18915,N_18322);
nor U19515 (N_19515,N_18680,N_18028);
and U19516 (N_19516,N_18787,N_18707);
or U19517 (N_19517,N_18811,N_18015);
or U19518 (N_19518,N_18535,N_18310);
and U19519 (N_19519,N_18749,N_18225);
xor U19520 (N_19520,N_18948,N_18762);
or U19521 (N_19521,N_18768,N_18196);
and U19522 (N_19522,N_18051,N_18356);
or U19523 (N_19523,N_18602,N_18075);
nand U19524 (N_19524,N_18720,N_18670);
or U19525 (N_19525,N_18215,N_18517);
nor U19526 (N_19526,N_18814,N_18507);
nor U19527 (N_19527,N_18687,N_18901);
or U19528 (N_19528,N_18005,N_18650);
and U19529 (N_19529,N_18799,N_18306);
nand U19530 (N_19530,N_18442,N_18525);
xnor U19531 (N_19531,N_18677,N_18726);
and U19532 (N_19532,N_18579,N_18102);
xnor U19533 (N_19533,N_18761,N_18015);
nand U19534 (N_19534,N_18423,N_18041);
xnor U19535 (N_19535,N_18114,N_18214);
and U19536 (N_19536,N_18939,N_18488);
or U19537 (N_19537,N_18272,N_18222);
nor U19538 (N_19538,N_18449,N_18266);
nor U19539 (N_19539,N_18093,N_18512);
nand U19540 (N_19540,N_18832,N_18983);
or U19541 (N_19541,N_18804,N_18111);
and U19542 (N_19542,N_18733,N_18665);
nor U19543 (N_19543,N_18664,N_18542);
or U19544 (N_19544,N_18573,N_18087);
nor U19545 (N_19545,N_18136,N_18651);
and U19546 (N_19546,N_18525,N_18352);
nand U19547 (N_19547,N_18847,N_18666);
xnor U19548 (N_19548,N_18664,N_18716);
xnor U19549 (N_19549,N_18957,N_18763);
and U19550 (N_19550,N_18918,N_18127);
and U19551 (N_19551,N_18883,N_18964);
and U19552 (N_19552,N_18191,N_18886);
xor U19553 (N_19553,N_18687,N_18885);
or U19554 (N_19554,N_18393,N_18113);
or U19555 (N_19555,N_18709,N_18504);
and U19556 (N_19556,N_18162,N_18495);
or U19557 (N_19557,N_18888,N_18204);
nand U19558 (N_19558,N_18980,N_18538);
nand U19559 (N_19559,N_18968,N_18242);
nor U19560 (N_19560,N_18878,N_18704);
or U19561 (N_19561,N_18527,N_18698);
nand U19562 (N_19562,N_18051,N_18461);
nor U19563 (N_19563,N_18912,N_18263);
and U19564 (N_19564,N_18394,N_18567);
xnor U19565 (N_19565,N_18016,N_18756);
nand U19566 (N_19566,N_18015,N_18208);
nor U19567 (N_19567,N_18494,N_18664);
nand U19568 (N_19568,N_18668,N_18245);
nor U19569 (N_19569,N_18298,N_18892);
nor U19570 (N_19570,N_18839,N_18406);
nand U19571 (N_19571,N_18801,N_18840);
nor U19572 (N_19572,N_18521,N_18673);
and U19573 (N_19573,N_18538,N_18813);
or U19574 (N_19574,N_18451,N_18356);
nand U19575 (N_19575,N_18681,N_18078);
nand U19576 (N_19576,N_18765,N_18962);
nand U19577 (N_19577,N_18637,N_18417);
or U19578 (N_19578,N_18236,N_18895);
nor U19579 (N_19579,N_18233,N_18833);
or U19580 (N_19580,N_18022,N_18576);
xnor U19581 (N_19581,N_18060,N_18183);
nand U19582 (N_19582,N_18980,N_18230);
nor U19583 (N_19583,N_18353,N_18016);
nand U19584 (N_19584,N_18415,N_18849);
nor U19585 (N_19585,N_18988,N_18695);
xnor U19586 (N_19586,N_18091,N_18421);
and U19587 (N_19587,N_18185,N_18935);
nor U19588 (N_19588,N_18478,N_18761);
nand U19589 (N_19589,N_18121,N_18288);
nor U19590 (N_19590,N_18217,N_18432);
nor U19591 (N_19591,N_18186,N_18793);
and U19592 (N_19592,N_18172,N_18231);
xor U19593 (N_19593,N_18480,N_18013);
nand U19594 (N_19594,N_18726,N_18273);
nor U19595 (N_19595,N_18675,N_18635);
and U19596 (N_19596,N_18809,N_18169);
nand U19597 (N_19597,N_18480,N_18797);
and U19598 (N_19598,N_18840,N_18464);
nor U19599 (N_19599,N_18452,N_18713);
nor U19600 (N_19600,N_18125,N_18061);
nand U19601 (N_19601,N_18575,N_18747);
nand U19602 (N_19602,N_18314,N_18803);
or U19603 (N_19603,N_18495,N_18190);
or U19604 (N_19604,N_18993,N_18623);
or U19605 (N_19605,N_18124,N_18338);
xor U19606 (N_19606,N_18363,N_18760);
nor U19607 (N_19607,N_18219,N_18775);
or U19608 (N_19608,N_18993,N_18313);
nand U19609 (N_19609,N_18528,N_18765);
and U19610 (N_19610,N_18531,N_18523);
and U19611 (N_19611,N_18849,N_18235);
nand U19612 (N_19612,N_18290,N_18042);
nor U19613 (N_19613,N_18509,N_18816);
nor U19614 (N_19614,N_18512,N_18664);
nor U19615 (N_19615,N_18178,N_18856);
or U19616 (N_19616,N_18416,N_18531);
and U19617 (N_19617,N_18977,N_18253);
and U19618 (N_19618,N_18028,N_18305);
xnor U19619 (N_19619,N_18554,N_18324);
nor U19620 (N_19620,N_18620,N_18055);
and U19621 (N_19621,N_18195,N_18214);
or U19622 (N_19622,N_18918,N_18004);
or U19623 (N_19623,N_18580,N_18402);
or U19624 (N_19624,N_18572,N_18422);
nor U19625 (N_19625,N_18519,N_18718);
or U19626 (N_19626,N_18164,N_18793);
nand U19627 (N_19627,N_18261,N_18401);
nand U19628 (N_19628,N_18665,N_18070);
nor U19629 (N_19629,N_18503,N_18936);
nand U19630 (N_19630,N_18640,N_18588);
nand U19631 (N_19631,N_18832,N_18264);
and U19632 (N_19632,N_18662,N_18171);
xnor U19633 (N_19633,N_18259,N_18707);
nand U19634 (N_19634,N_18232,N_18567);
and U19635 (N_19635,N_18972,N_18464);
nor U19636 (N_19636,N_18449,N_18019);
or U19637 (N_19637,N_18330,N_18441);
xnor U19638 (N_19638,N_18228,N_18338);
nand U19639 (N_19639,N_18513,N_18961);
nor U19640 (N_19640,N_18151,N_18985);
nor U19641 (N_19641,N_18759,N_18064);
nor U19642 (N_19642,N_18114,N_18098);
and U19643 (N_19643,N_18690,N_18283);
nand U19644 (N_19644,N_18744,N_18752);
or U19645 (N_19645,N_18066,N_18414);
nor U19646 (N_19646,N_18962,N_18900);
or U19647 (N_19647,N_18927,N_18157);
nand U19648 (N_19648,N_18482,N_18613);
xor U19649 (N_19649,N_18368,N_18424);
and U19650 (N_19650,N_18384,N_18940);
xnor U19651 (N_19651,N_18632,N_18627);
or U19652 (N_19652,N_18632,N_18662);
nor U19653 (N_19653,N_18783,N_18090);
nor U19654 (N_19654,N_18106,N_18120);
nor U19655 (N_19655,N_18618,N_18977);
nand U19656 (N_19656,N_18080,N_18370);
and U19657 (N_19657,N_18907,N_18892);
and U19658 (N_19658,N_18433,N_18331);
and U19659 (N_19659,N_18528,N_18896);
or U19660 (N_19660,N_18868,N_18033);
nand U19661 (N_19661,N_18426,N_18260);
xnor U19662 (N_19662,N_18639,N_18608);
nand U19663 (N_19663,N_18250,N_18020);
nor U19664 (N_19664,N_18669,N_18158);
or U19665 (N_19665,N_18702,N_18173);
or U19666 (N_19666,N_18677,N_18081);
nor U19667 (N_19667,N_18737,N_18293);
and U19668 (N_19668,N_18407,N_18574);
xor U19669 (N_19669,N_18772,N_18083);
xor U19670 (N_19670,N_18357,N_18719);
or U19671 (N_19671,N_18426,N_18731);
or U19672 (N_19672,N_18187,N_18105);
nor U19673 (N_19673,N_18019,N_18762);
nor U19674 (N_19674,N_18675,N_18209);
nand U19675 (N_19675,N_18378,N_18640);
or U19676 (N_19676,N_18022,N_18774);
or U19677 (N_19677,N_18143,N_18672);
or U19678 (N_19678,N_18411,N_18414);
nor U19679 (N_19679,N_18022,N_18021);
xnor U19680 (N_19680,N_18743,N_18252);
or U19681 (N_19681,N_18624,N_18185);
and U19682 (N_19682,N_18202,N_18372);
nor U19683 (N_19683,N_18653,N_18183);
and U19684 (N_19684,N_18739,N_18501);
and U19685 (N_19685,N_18985,N_18178);
nor U19686 (N_19686,N_18774,N_18427);
xor U19687 (N_19687,N_18245,N_18903);
or U19688 (N_19688,N_18571,N_18973);
and U19689 (N_19689,N_18264,N_18110);
or U19690 (N_19690,N_18961,N_18001);
or U19691 (N_19691,N_18386,N_18764);
xnor U19692 (N_19692,N_18039,N_18680);
or U19693 (N_19693,N_18091,N_18669);
or U19694 (N_19694,N_18110,N_18549);
nor U19695 (N_19695,N_18857,N_18426);
nor U19696 (N_19696,N_18129,N_18877);
and U19697 (N_19697,N_18709,N_18011);
nand U19698 (N_19698,N_18072,N_18600);
nor U19699 (N_19699,N_18690,N_18608);
nand U19700 (N_19700,N_18190,N_18771);
nand U19701 (N_19701,N_18364,N_18538);
or U19702 (N_19702,N_18692,N_18675);
nor U19703 (N_19703,N_18452,N_18695);
nor U19704 (N_19704,N_18776,N_18803);
or U19705 (N_19705,N_18496,N_18324);
xor U19706 (N_19706,N_18623,N_18895);
or U19707 (N_19707,N_18835,N_18179);
or U19708 (N_19708,N_18873,N_18600);
xnor U19709 (N_19709,N_18241,N_18592);
nor U19710 (N_19710,N_18195,N_18403);
xor U19711 (N_19711,N_18512,N_18687);
nand U19712 (N_19712,N_18714,N_18354);
xor U19713 (N_19713,N_18174,N_18854);
or U19714 (N_19714,N_18972,N_18456);
nand U19715 (N_19715,N_18978,N_18572);
xnor U19716 (N_19716,N_18981,N_18924);
nand U19717 (N_19717,N_18277,N_18351);
or U19718 (N_19718,N_18473,N_18421);
and U19719 (N_19719,N_18575,N_18908);
or U19720 (N_19720,N_18878,N_18177);
nand U19721 (N_19721,N_18487,N_18001);
and U19722 (N_19722,N_18983,N_18160);
nand U19723 (N_19723,N_18805,N_18818);
xnor U19724 (N_19724,N_18312,N_18835);
nor U19725 (N_19725,N_18369,N_18166);
and U19726 (N_19726,N_18149,N_18892);
or U19727 (N_19727,N_18034,N_18525);
and U19728 (N_19728,N_18575,N_18238);
or U19729 (N_19729,N_18839,N_18662);
and U19730 (N_19730,N_18703,N_18970);
nand U19731 (N_19731,N_18218,N_18341);
nand U19732 (N_19732,N_18977,N_18809);
xor U19733 (N_19733,N_18958,N_18102);
nor U19734 (N_19734,N_18970,N_18250);
and U19735 (N_19735,N_18912,N_18829);
nor U19736 (N_19736,N_18983,N_18138);
nand U19737 (N_19737,N_18533,N_18250);
nand U19738 (N_19738,N_18945,N_18148);
nor U19739 (N_19739,N_18459,N_18184);
nor U19740 (N_19740,N_18806,N_18278);
nor U19741 (N_19741,N_18302,N_18820);
nand U19742 (N_19742,N_18385,N_18799);
or U19743 (N_19743,N_18353,N_18012);
xor U19744 (N_19744,N_18035,N_18194);
xnor U19745 (N_19745,N_18539,N_18899);
nor U19746 (N_19746,N_18181,N_18782);
or U19747 (N_19747,N_18106,N_18045);
or U19748 (N_19748,N_18035,N_18004);
nand U19749 (N_19749,N_18314,N_18262);
nor U19750 (N_19750,N_18073,N_18046);
xor U19751 (N_19751,N_18691,N_18184);
and U19752 (N_19752,N_18749,N_18238);
nand U19753 (N_19753,N_18580,N_18278);
nor U19754 (N_19754,N_18696,N_18395);
nor U19755 (N_19755,N_18282,N_18296);
xnor U19756 (N_19756,N_18512,N_18692);
and U19757 (N_19757,N_18718,N_18813);
and U19758 (N_19758,N_18221,N_18923);
or U19759 (N_19759,N_18838,N_18232);
nand U19760 (N_19760,N_18083,N_18210);
xnor U19761 (N_19761,N_18202,N_18723);
nor U19762 (N_19762,N_18362,N_18475);
nand U19763 (N_19763,N_18628,N_18506);
and U19764 (N_19764,N_18559,N_18944);
nand U19765 (N_19765,N_18894,N_18897);
xnor U19766 (N_19766,N_18799,N_18874);
nor U19767 (N_19767,N_18775,N_18985);
and U19768 (N_19768,N_18220,N_18240);
xnor U19769 (N_19769,N_18543,N_18537);
and U19770 (N_19770,N_18312,N_18229);
nor U19771 (N_19771,N_18579,N_18256);
nand U19772 (N_19772,N_18998,N_18421);
or U19773 (N_19773,N_18649,N_18851);
nand U19774 (N_19774,N_18073,N_18568);
or U19775 (N_19775,N_18129,N_18303);
or U19776 (N_19776,N_18309,N_18758);
xor U19777 (N_19777,N_18071,N_18153);
xnor U19778 (N_19778,N_18396,N_18782);
and U19779 (N_19779,N_18391,N_18276);
or U19780 (N_19780,N_18544,N_18073);
nand U19781 (N_19781,N_18169,N_18552);
nand U19782 (N_19782,N_18044,N_18974);
xor U19783 (N_19783,N_18631,N_18955);
nor U19784 (N_19784,N_18943,N_18150);
and U19785 (N_19785,N_18408,N_18382);
nand U19786 (N_19786,N_18136,N_18366);
nand U19787 (N_19787,N_18888,N_18189);
nand U19788 (N_19788,N_18431,N_18126);
and U19789 (N_19789,N_18240,N_18751);
or U19790 (N_19790,N_18972,N_18428);
nor U19791 (N_19791,N_18008,N_18140);
xor U19792 (N_19792,N_18992,N_18068);
nor U19793 (N_19793,N_18347,N_18130);
nand U19794 (N_19794,N_18460,N_18694);
xnor U19795 (N_19795,N_18246,N_18342);
xor U19796 (N_19796,N_18751,N_18680);
or U19797 (N_19797,N_18206,N_18387);
nor U19798 (N_19798,N_18514,N_18011);
nand U19799 (N_19799,N_18325,N_18832);
nor U19800 (N_19800,N_18935,N_18103);
nand U19801 (N_19801,N_18856,N_18559);
or U19802 (N_19802,N_18788,N_18548);
or U19803 (N_19803,N_18075,N_18154);
xnor U19804 (N_19804,N_18427,N_18406);
xor U19805 (N_19805,N_18177,N_18780);
xor U19806 (N_19806,N_18619,N_18070);
xor U19807 (N_19807,N_18094,N_18690);
or U19808 (N_19808,N_18288,N_18299);
and U19809 (N_19809,N_18340,N_18985);
and U19810 (N_19810,N_18541,N_18918);
or U19811 (N_19811,N_18508,N_18535);
and U19812 (N_19812,N_18185,N_18747);
nand U19813 (N_19813,N_18266,N_18569);
nor U19814 (N_19814,N_18127,N_18961);
or U19815 (N_19815,N_18206,N_18584);
nor U19816 (N_19816,N_18983,N_18065);
or U19817 (N_19817,N_18457,N_18201);
and U19818 (N_19818,N_18200,N_18551);
nand U19819 (N_19819,N_18791,N_18894);
or U19820 (N_19820,N_18211,N_18325);
nand U19821 (N_19821,N_18509,N_18675);
or U19822 (N_19822,N_18076,N_18106);
and U19823 (N_19823,N_18104,N_18002);
xnor U19824 (N_19824,N_18142,N_18187);
xor U19825 (N_19825,N_18097,N_18349);
nor U19826 (N_19826,N_18139,N_18384);
nand U19827 (N_19827,N_18483,N_18686);
nand U19828 (N_19828,N_18197,N_18417);
and U19829 (N_19829,N_18101,N_18808);
or U19830 (N_19830,N_18308,N_18830);
or U19831 (N_19831,N_18059,N_18479);
nand U19832 (N_19832,N_18452,N_18532);
nor U19833 (N_19833,N_18019,N_18583);
or U19834 (N_19834,N_18525,N_18330);
nand U19835 (N_19835,N_18911,N_18335);
and U19836 (N_19836,N_18714,N_18720);
and U19837 (N_19837,N_18881,N_18834);
nand U19838 (N_19838,N_18359,N_18657);
nor U19839 (N_19839,N_18902,N_18607);
and U19840 (N_19840,N_18817,N_18139);
xor U19841 (N_19841,N_18226,N_18691);
or U19842 (N_19842,N_18049,N_18522);
xnor U19843 (N_19843,N_18418,N_18649);
xor U19844 (N_19844,N_18119,N_18770);
or U19845 (N_19845,N_18253,N_18622);
xnor U19846 (N_19846,N_18489,N_18913);
xnor U19847 (N_19847,N_18596,N_18696);
xnor U19848 (N_19848,N_18139,N_18924);
xnor U19849 (N_19849,N_18251,N_18400);
nor U19850 (N_19850,N_18955,N_18907);
nor U19851 (N_19851,N_18899,N_18507);
nor U19852 (N_19852,N_18948,N_18889);
and U19853 (N_19853,N_18492,N_18535);
nor U19854 (N_19854,N_18488,N_18917);
xor U19855 (N_19855,N_18172,N_18155);
xor U19856 (N_19856,N_18514,N_18584);
or U19857 (N_19857,N_18884,N_18036);
or U19858 (N_19858,N_18484,N_18639);
or U19859 (N_19859,N_18376,N_18341);
nor U19860 (N_19860,N_18123,N_18395);
or U19861 (N_19861,N_18615,N_18992);
nor U19862 (N_19862,N_18457,N_18608);
nor U19863 (N_19863,N_18955,N_18784);
nand U19864 (N_19864,N_18161,N_18790);
nand U19865 (N_19865,N_18422,N_18244);
xnor U19866 (N_19866,N_18767,N_18194);
and U19867 (N_19867,N_18960,N_18030);
or U19868 (N_19868,N_18224,N_18496);
nand U19869 (N_19869,N_18882,N_18827);
and U19870 (N_19870,N_18519,N_18177);
nor U19871 (N_19871,N_18807,N_18245);
xor U19872 (N_19872,N_18184,N_18061);
or U19873 (N_19873,N_18851,N_18537);
and U19874 (N_19874,N_18704,N_18369);
or U19875 (N_19875,N_18358,N_18115);
nand U19876 (N_19876,N_18709,N_18151);
nand U19877 (N_19877,N_18494,N_18957);
nor U19878 (N_19878,N_18678,N_18908);
nand U19879 (N_19879,N_18315,N_18457);
or U19880 (N_19880,N_18035,N_18601);
nand U19881 (N_19881,N_18156,N_18747);
nor U19882 (N_19882,N_18973,N_18612);
or U19883 (N_19883,N_18127,N_18159);
or U19884 (N_19884,N_18988,N_18275);
nand U19885 (N_19885,N_18818,N_18568);
nand U19886 (N_19886,N_18794,N_18391);
or U19887 (N_19887,N_18358,N_18399);
and U19888 (N_19888,N_18597,N_18349);
or U19889 (N_19889,N_18228,N_18042);
nor U19890 (N_19890,N_18347,N_18840);
nor U19891 (N_19891,N_18248,N_18360);
or U19892 (N_19892,N_18860,N_18220);
and U19893 (N_19893,N_18142,N_18067);
or U19894 (N_19894,N_18023,N_18301);
or U19895 (N_19895,N_18618,N_18275);
nor U19896 (N_19896,N_18780,N_18345);
xnor U19897 (N_19897,N_18463,N_18560);
and U19898 (N_19898,N_18398,N_18976);
nand U19899 (N_19899,N_18551,N_18405);
and U19900 (N_19900,N_18254,N_18287);
or U19901 (N_19901,N_18487,N_18745);
nor U19902 (N_19902,N_18867,N_18756);
nand U19903 (N_19903,N_18541,N_18596);
or U19904 (N_19904,N_18525,N_18538);
nor U19905 (N_19905,N_18276,N_18833);
and U19906 (N_19906,N_18922,N_18123);
xor U19907 (N_19907,N_18979,N_18557);
and U19908 (N_19908,N_18165,N_18185);
or U19909 (N_19909,N_18458,N_18384);
nor U19910 (N_19910,N_18103,N_18514);
xnor U19911 (N_19911,N_18362,N_18277);
nor U19912 (N_19912,N_18141,N_18453);
nand U19913 (N_19913,N_18664,N_18826);
xor U19914 (N_19914,N_18513,N_18912);
nor U19915 (N_19915,N_18655,N_18642);
xor U19916 (N_19916,N_18745,N_18452);
nand U19917 (N_19917,N_18928,N_18559);
and U19918 (N_19918,N_18486,N_18788);
nand U19919 (N_19919,N_18814,N_18136);
nand U19920 (N_19920,N_18465,N_18071);
nand U19921 (N_19921,N_18892,N_18608);
nand U19922 (N_19922,N_18034,N_18550);
and U19923 (N_19923,N_18270,N_18592);
nor U19924 (N_19924,N_18021,N_18188);
or U19925 (N_19925,N_18123,N_18629);
xor U19926 (N_19926,N_18059,N_18884);
xor U19927 (N_19927,N_18491,N_18401);
and U19928 (N_19928,N_18912,N_18262);
and U19929 (N_19929,N_18158,N_18449);
nor U19930 (N_19930,N_18927,N_18689);
nand U19931 (N_19931,N_18475,N_18366);
xor U19932 (N_19932,N_18244,N_18148);
or U19933 (N_19933,N_18360,N_18070);
nor U19934 (N_19934,N_18356,N_18000);
and U19935 (N_19935,N_18172,N_18118);
xor U19936 (N_19936,N_18775,N_18403);
or U19937 (N_19937,N_18063,N_18903);
or U19938 (N_19938,N_18351,N_18912);
or U19939 (N_19939,N_18310,N_18214);
nor U19940 (N_19940,N_18971,N_18058);
xnor U19941 (N_19941,N_18850,N_18549);
nor U19942 (N_19942,N_18649,N_18023);
xor U19943 (N_19943,N_18365,N_18367);
nor U19944 (N_19944,N_18792,N_18270);
nor U19945 (N_19945,N_18409,N_18857);
or U19946 (N_19946,N_18113,N_18292);
nor U19947 (N_19947,N_18526,N_18235);
xnor U19948 (N_19948,N_18893,N_18729);
nor U19949 (N_19949,N_18918,N_18036);
nand U19950 (N_19950,N_18571,N_18007);
xnor U19951 (N_19951,N_18545,N_18800);
or U19952 (N_19952,N_18597,N_18710);
nor U19953 (N_19953,N_18961,N_18360);
or U19954 (N_19954,N_18123,N_18722);
nor U19955 (N_19955,N_18429,N_18630);
or U19956 (N_19956,N_18559,N_18942);
nand U19957 (N_19957,N_18687,N_18372);
nand U19958 (N_19958,N_18471,N_18626);
or U19959 (N_19959,N_18625,N_18261);
nand U19960 (N_19960,N_18939,N_18145);
and U19961 (N_19961,N_18903,N_18206);
nand U19962 (N_19962,N_18880,N_18207);
nand U19963 (N_19963,N_18679,N_18064);
xor U19964 (N_19964,N_18144,N_18042);
and U19965 (N_19965,N_18033,N_18671);
and U19966 (N_19966,N_18167,N_18384);
nand U19967 (N_19967,N_18135,N_18515);
or U19968 (N_19968,N_18273,N_18000);
nor U19969 (N_19969,N_18922,N_18515);
and U19970 (N_19970,N_18203,N_18065);
xnor U19971 (N_19971,N_18412,N_18938);
nand U19972 (N_19972,N_18505,N_18572);
or U19973 (N_19973,N_18613,N_18634);
xnor U19974 (N_19974,N_18759,N_18485);
nor U19975 (N_19975,N_18625,N_18108);
nor U19976 (N_19976,N_18078,N_18852);
or U19977 (N_19977,N_18047,N_18138);
nand U19978 (N_19978,N_18631,N_18614);
or U19979 (N_19979,N_18573,N_18263);
xor U19980 (N_19980,N_18011,N_18289);
nor U19981 (N_19981,N_18745,N_18031);
and U19982 (N_19982,N_18861,N_18869);
nor U19983 (N_19983,N_18345,N_18929);
nand U19984 (N_19984,N_18544,N_18185);
xor U19985 (N_19985,N_18096,N_18445);
nand U19986 (N_19986,N_18465,N_18291);
nor U19987 (N_19987,N_18613,N_18918);
and U19988 (N_19988,N_18159,N_18193);
nor U19989 (N_19989,N_18720,N_18291);
nor U19990 (N_19990,N_18197,N_18914);
and U19991 (N_19991,N_18647,N_18773);
xnor U19992 (N_19992,N_18034,N_18669);
or U19993 (N_19993,N_18834,N_18529);
xor U19994 (N_19994,N_18935,N_18170);
xnor U19995 (N_19995,N_18100,N_18553);
nor U19996 (N_19996,N_18395,N_18739);
or U19997 (N_19997,N_18103,N_18599);
or U19998 (N_19998,N_18873,N_18690);
and U19999 (N_19999,N_18660,N_18724);
nand U20000 (N_20000,N_19893,N_19560);
nand U20001 (N_20001,N_19946,N_19666);
nand U20002 (N_20002,N_19591,N_19119);
nand U20003 (N_20003,N_19207,N_19442);
and U20004 (N_20004,N_19278,N_19901);
xnor U20005 (N_20005,N_19972,N_19269);
nand U20006 (N_20006,N_19483,N_19837);
or U20007 (N_20007,N_19768,N_19225);
or U20008 (N_20008,N_19685,N_19998);
and U20009 (N_20009,N_19538,N_19910);
xor U20010 (N_20010,N_19782,N_19062);
or U20011 (N_20011,N_19005,N_19715);
nand U20012 (N_20012,N_19969,N_19667);
or U20013 (N_20013,N_19510,N_19388);
and U20014 (N_20014,N_19630,N_19822);
or U20015 (N_20015,N_19522,N_19279);
nor U20016 (N_20016,N_19475,N_19897);
or U20017 (N_20017,N_19034,N_19178);
and U20018 (N_20018,N_19230,N_19850);
nor U20019 (N_20019,N_19356,N_19835);
or U20020 (N_20020,N_19843,N_19481);
xor U20021 (N_20021,N_19504,N_19749);
and U20022 (N_20022,N_19792,N_19721);
xnor U20023 (N_20023,N_19010,N_19929);
nand U20024 (N_20024,N_19271,N_19675);
or U20025 (N_20025,N_19760,N_19750);
or U20026 (N_20026,N_19620,N_19347);
or U20027 (N_20027,N_19416,N_19970);
nand U20028 (N_20028,N_19135,N_19680);
nor U20029 (N_20029,N_19171,N_19950);
and U20030 (N_20030,N_19267,N_19864);
or U20031 (N_20031,N_19447,N_19916);
nand U20032 (N_20032,N_19917,N_19148);
nor U20033 (N_20033,N_19352,N_19439);
nor U20034 (N_20034,N_19490,N_19928);
xnor U20035 (N_20035,N_19016,N_19369);
nand U20036 (N_20036,N_19121,N_19213);
nand U20037 (N_20037,N_19492,N_19624);
nand U20038 (N_20038,N_19714,N_19634);
nor U20039 (N_20039,N_19006,N_19384);
nor U20040 (N_20040,N_19628,N_19737);
or U20041 (N_20041,N_19240,N_19825);
nand U20042 (N_20042,N_19488,N_19453);
or U20043 (N_20043,N_19875,N_19988);
nand U20044 (N_20044,N_19736,N_19373);
or U20045 (N_20045,N_19498,N_19295);
or U20046 (N_20046,N_19212,N_19017);
and U20047 (N_20047,N_19274,N_19090);
xnor U20048 (N_20048,N_19283,N_19505);
nor U20049 (N_20049,N_19124,N_19434);
nand U20050 (N_20050,N_19186,N_19469);
and U20051 (N_20051,N_19448,N_19131);
nand U20052 (N_20052,N_19605,N_19994);
and U20053 (N_20053,N_19661,N_19256);
nor U20054 (N_20054,N_19912,N_19487);
nand U20055 (N_20055,N_19933,N_19085);
nand U20056 (N_20056,N_19165,N_19080);
xor U20057 (N_20057,N_19349,N_19519);
or U20058 (N_20058,N_19745,N_19470);
nand U20059 (N_20059,N_19321,N_19486);
xnor U20060 (N_20060,N_19293,N_19451);
and U20061 (N_20061,N_19799,N_19597);
or U20062 (N_20062,N_19140,N_19095);
nor U20063 (N_20063,N_19485,N_19502);
nor U20064 (N_20064,N_19073,N_19342);
xnor U20065 (N_20065,N_19662,N_19518);
or U20066 (N_20066,N_19294,N_19019);
nor U20067 (N_20067,N_19888,N_19215);
and U20068 (N_20068,N_19959,N_19691);
nor U20069 (N_20069,N_19590,N_19372);
or U20070 (N_20070,N_19652,N_19687);
nand U20071 (N_20071,N_19922,N_19094);
or U20072 (N_20072,N_19371,N_19291);
and U20073 (N_20073,N_19851,N_19249);
and U20074 (N_20074,N_19194,N_19462);
nor U20075 (N_20075,N_19930,N_19823);
or U20076 (N_20076,N_19325,N_19552);
xnor U20077 (N_20077,N_19397,N_19414);
or U20078 (N_20078,N_19264,N_19364);
and U20079 (N_20079,N_19335,N_19855);
nor U20080 (N_20080,N_19104,N_19746);
or U20081 (N_20081,N_19698,N_19508);
nor U20082 (N_20082,N_19586,N_19748);
and U20083 (N_20083,N_19198,N_19100);
nor U20084 (N_20084,N_19362,N_19753);
nand U20085 (N_20085,N_19789,N_19257);
and U20086 (N_20086,N_19568,N_19758);
nand U20087 (N_20087,N_19684,N_19730);
and U20088 (N_20088,N_19322,N_19220);
or U20089 (N_20089,N_19868,N_19067);
xnor U20090 (N_20090,N_19682,N_19467);
xnor U20091 (N_20091,N_19553,N_19353);
xnor U20092 (N_20092,N_19169,N_19339);
or U20093 (N_20093,N_19044,N_19253);
and U20094 (N_20094,N_19204,N_19642);
nor U20095 (N_20095,N_19881,N_19379);
nor U20096 (N_20096,N_19791,N_19811);
nor U20097 (N_20097,N_19132,N_19513);
nand U20098 (N_20098,N_19557,N_19027);
xor U20099 (N_20099,N_19996,N_19232);
xnor U20100 (N_20100,N_19457,N_19593);
nor U20101 (N_20101,N_19966,N_19587);
or U20102 (N_20102,N_19637,N_19218);
and U20103 (N_20103,N_19292,N_19944);
or U20104 (N_20104,N_19656,N_19188);
or U20105 (N_20105,N_19496,N_19381);
or U20106 (N_20106,N_19138,N_19201);
nand U20107 (N_20107,N_19111,N_19474);
nor U20108 (N_20108,N_19221,N_19506);
nand U20109 (N_20109,N_19683,N_19906);
xor U20110 (N_20110,N_19535,N_19246);
nand U20111 (N_20111,N_19521,N_19625);
or U20112 (N_20112,N_19156,N_19526);
xnor U20113 (N_20113,N_19826,N_19890);
xor U20114 (N_20114,N_19979,N_19742);
or U20115 (N_20115,N_19733,N_19978);
or U20116 (N_20116,N_19524,N_19954);
nor U20117 (N_20117,N_19144,N_19117);
and U20118 (N_20118,N_19626,N_19007);
xnor U20119 (N_20119,N_19167,N_19895);
nor U20120 (N_20120,N_19407,N_19761);
xor U20121 (N_20121,N_19842,N_19960);
xor U20122 (N_20122,N_19456,N_19082);
xor U20123 (N_20123,N_19290,N_19306);
nand U20124 (N_20124,N_19341,N_19641);
xnor U20125 (N_20125,N_19635,N_19987);
xnor U20126 (N_20126,N_19192,N_19468);
nand U20127 (N_20127,N_19412,N_19766);
nand U20128 (N_20128,N_19941,N_19147);
nand U20129 (N_20129,N_19162,N_19939);
xnor U20130 (N_20130,N_19125,N_19182);
or U20131 (N_20131,N_19801,N_19904);
nand U20132 (N_20132,N_19350,N_19810);
nand U20133 (N_20133,N_19075,N_19337);
and U20134 (N_20134,N_19907,N_19478);
nor U20135 (N_20135,N_19055,N_19976);
and U20136 (N_20136,N_19619,N_19032);
xor U20137 (N_20137,N_19920,N_19458);
nor U20138 (N_20138,N_19298,N_19035);
and U20139 (N_20139,N_19814,N_19716);
nor U20140 (N_20140,N_19613,N_19255);
nand U20141 (N_20141,N_19284,N_19563);
nor U20142 (N_20142,N_19719,N_19103);
or U20143 (N_20143,N_19202,N_19426);
or U20144 (N_20144,N_19049,N_19289);
xnor U20145 (N_20145,N_19849,N_19217);
or U20146 (N_20146,N_19479,N_19168);
and U20147 (N_20147,N_19455,N_19759);
xor U20148 (N_20148,N_19551,N_19208);
nor U20149 (N_20149,N_19564,N_19919);
xor U20150 (N_20150,N_19744,N_19064);
or U20151 (N_20151,N_19640,N_19435);
nor U20152 (N_20152,N_19909,N_19270);
and U20153 (N_20153,N_19884,N_19541);
or U20154 (N_20154,N_19161,N_19530);
xnor U20155 (N_20155,N_19495,N_19664);
xnor U20156 (N_20156,N_19203,N_19892);
nor U20157 (N_20157,N_19422,N_19237);
or U20158 (N_20158,N_19376,N_19860);
and U20159 (N_20159,N_19818,N_19989);
or U20160 (N_20160,N_19913,N_19367);
and U20161 (N_20161,N_19784,N_19967);
or U20162 (N_20162,N_19644,N_19840);
xor U20163 (N_20163,N_19011,N_19210);
nand U20164 (N_20164,N_19172,N_19785);
xnor U20165 (N_20165,N_19804,N_19392);
and U20166 (N_20166,N_19594,N_19238);
nor U20167 (N_20167,N_19588,N_19399);
and U20168 (N_20168,N_19874,N_19977);
or U20169 (N_20169,N_19756,N_19421);
or U20170 (N_20170,N_19394,N_19424);
nand U20171 (N_20171,N_19889,N_19400);
xor U20172 (N_20172,N_19183,N_19561);
and U20173 (N_20173,N_19657,N_19710);
xor U20174 (N_20174,N_19779,N_19562);
xor U20175 (N_20175,N_19187,N_19627);
xnor U20176 (N_20176,N_19107,N_19465);
or U20177 (N_20177,N_19673,N_19190);
or U20178 (N_20178,N_19176,N_19146);
xor U20179 (N_20179,N_19450,N_19320);
and U20180 (N_20180,N_19038,N_19956);
xnor U20181 (N_20181,N_19351,N_19741);
xnor U20182 (N_20182,N_19821,N_19209);
and U20183 (N_20183,N_19357,N_19360);
nor U20184 (N_20184,N_19806,N_19589);
xor U20185 (N_20185,N_19409,N_19430);
nor U20186 (N_20186,N_19155,N_19793);
nand U20187 (N_20187,N_19558,N_19420);
and U20188 (N_20188,N_19765,N_19332);
nor U20189 (N_20189,N_19654,N_19219);
nor U20190 (N_20190,N_19815,N_19918);
nor U20191 (N_20191,N_19728,N_19948);
nor U20192 (N_20192,N_19199,N_19983);
nor U20193 (N_20193,N_19297,N_19261);
xor U20194 (N_20194,N_19859,N_19711);
and U20195 (N_20195,N_19343,N_19771);
and U20196 (N_20196,N_19705,N_19757);
nand U20197 (N_20197,N_19239,N_19299);
nor U20198 (N_20198,N_19031,N_19039);
or U20199 (N_20199,N_19145,N_19370);
nand U20200 (N_20200,N_19277,N_19309);
and U20201 (N_20201,N_19947,N_19528);
or U20202 (N_20202,N_19489,N_19908);
nand U20203 (N_20203,N_19731,N_19681);
or U20204 (N_20204,N_19798,N_19633);
or U20205 (N_20205,N_19401,N_19962);
xnor U20206 (N_20206,N_19428,N_19051);
and U20207 (N_20207,N_19417,N_19263);
nand U20208 (N_20208,N_19053,N_19047);
xor U20209 (N_20209,N_19778,N_19054);
and U20210 (N_20210,N_19612,N_19911);
and U20211 (N_20211,N_19014,N_19026);
or U20212 (N_20212,N_19328,N_19709);
xor U20213 (N_20213,N_19025,N_19653);
nor U20214 (N_20214,N_19878,N_19595);
and U20215 (N_20215,N_19216,N_19582);
or U20216 (N_20216,N_19195,N_19565);
or U20217 (N_20217,N_19554,N_19830);
and U20218 (N_20218,N_19173,N_19068);
or U20219 (N_20219,N_19762,N_19340);
xnor U20220 (N_20220,N_19385,N_19958);
nand U20221 (N_20221,N_19752,N_19266);
nand U20222 (N_20222,N_19797,N_19193);
nor U20223 (N_20223,N_19235,N_19317);
nand U20224 (N_20224,N_19775,N_19265);
or U20225 (N_20225,N_19807,N_19050);
nor U20226 (N_20226,N_19460,N_19608);
xor U20227 (N_20227,N_19514,N_19833);
and U20228 (N_20228,N_19924,N_19272);
nand U20229 (N_20229,N_19985,N_19346);
and U20230 (N_20230,N_19431,N_19720);
nor U20231 (N_20231,N_19233,N_19938);
xor U20232 (N_20232,N_19993,N_19990);
nand U20233 (N_20233,N_19477,N_19886);
or U20234 (N_20234,N_19268,N_19312);
xnor U20235 (N_20235,N_19527,N_19729);
or U20236 (N_20236,N_19764,N_19609);
nor U20237 (N_20237,N_19882,N_19816);
nand U20238 (N_20238,N_19348,N_19022);
or U20239 (N_20239,N_19197,N_19905);
or U20240 (N_20240,N_19338,N_19493);
nand U20241 (N_20241,N_19639,N_19224);
or U20242 (N_20242,N_19048,N_19914);
and U20243 (N_20243,N_19160,N_19543);
and U20244 (N_20244,N_19122,N_19252);
and U20245 (N_20245,N_19607,N_19699);
xnor U20246 (N_20246,N_19743,N_19577);
nor U20247 (N_20247,N_19559,N_19157);
or U20248 (N_20248,N_19942,N_19516);
or U20249 (N_20249,N_19894,N_19196);
nor U20250 (N_20250,N_19056,N_19177);
nor U20251 (N_20251,N_19275,N_19689);
and U20252 (N_20252,N_19316,N_19432);
or U20253 (N_20253,N_19857,N_19033);
or U20254 (N_20254,N_19110,N_19688);
nor U20255 (N_20255,N_19181,N_19602);
and U20256 (N_20256,N_19128,N_19581);
and U20257 (N_20257,N_19126,N_19647);
nand U20258 (N_20258,N_19902,N_19393);
nand U20259 (N_20259,N_19174,N_19674);
and U20260 (N_20260,N_19623,N_19229);
or U20261 (N_20261,N_19735,N_19898);
or U20262 (N_20262,N_19153,N_19961);
or U20263 (N_20263,N_19867,N_19858);
xor U20264 (N_20264,N_19361,N_19540);
nor U20265 (N_20265,N_19621,N_19088);
nand U20266 (N_20266,N_19323,N_19517);
nor U20267 (N_20267,N_19002,N_19824);
xnor U20268 (N_20268,N_19755,N_19576);
nor U20269 (N_20269,N_19787,N_19276);
nand U20270 (N_20270,N_19081,N_19191);
nand U20271 (N_20271,N_19604,N_19115);
nand U20272 (N_20272,N_19651,N_19872);
and U20273 (N_20273,N_19045,N_19658);
and U20274 (N_20274,N_19141,N_19550);
or U20275 (N_20275,N_19795,N_19041);
xor U20276 (N_20276,N_19114,N_19314);
nand U20277 (N_20277,N_19231,N_19001);
and U20278 (N_20278,N_19973,N_19794);
xnor U20279 (N_20279,N_19767,N_19387);
xnor U20280 (N_20280,N_19763,N_19102);
xnor U20281 (N_20281,N_19015,N_19503);
nand U20282 (N_20282,N_19712,N_19777);
and U20283 (N_20283,N_19109,N_19163);
nand U20284 (N_20284,N_19573,N_19004);
nand U20285 (N_20285,N_19703,N_19258);
xnor U20286 (N_20286,N_19288,N_19052);
or U20287 (N_20287,N_19812,N_19441);
and U20288 (N_20288,N_19411,N_19499);
or U20289 (N_20289,N_19515,N_19836);
and U20290 (N_20290,N_19286,N_19772);
nand U20291 (N_20291,N_19433,N_19984);
nand U20292 (N_20292,N_19395,N_19690);
and U20293 (N_20293,N_19139,N_19774);
and U20294 (N_20294,N_19834,N_19964);
nor U20295 (N_20295,N_19154,N_19861);
nand U20296 (N_20296,N_19000,N_19180);
nor U20297 (N_20297,N_19136,N_19925);
nand U20298 (N_20298,N_19243,N_19606);
and U20299 (N_20299,N_19869,N_19366);
xnor U20300 (N_20300,N_19358,N_19065);
or U20301 (N_20301,N_19324,N_19018);
xnor U20302 (N_20302,N_19086,N_19643);
nand U20303 (N_20303,N_19660,N_19547);
and U20304 (N_20304,N_19596,N_19273);
and U20305 (N_20305,N_19009,N_19622);
and U20306 (N_20306,N_19648,N_19028);
xnor U20307 (N_20307,N_19404,N_19423);
xnor U20308 (N_20308,N_19319,N_19368);
nor U20309 (N_20309,N_19365,N_19092);
nor U20310 (N_20310,N_19382,N_19649);
xor U20311 (N_20311,N_19251,N_19659);
nor U20312 (N_20312,N_19981,N_19436);
or U20313 (N_20313,N_19112,N_19301);
and U20314 (N_20314,N_19900,N_19935);
nand U20315 (N_20315,N_19402,N_19310);
or U20316 (N_20316,N_19079,N_19800);
xnor U20317 (N_20317,N_19677,N_19438);
xnor U20318 (N_20318,N_19214,N_19072);
and U20319 (N_20319,N_19694,N_19780);
xnor U20320 (N_20320,N_19975,N_19704);
or U20321 (N_20321,N_19727,N_19440);
xor U20322 (N_20322,N_19548,N_19040);
or U20323 (N_20323,N_19702,N_19802);
and U20324 (N_20324,N_19571,N_19839);
nand U20325 (N_20325,N_19334,N_19724);
nand U20326 (N_20326,N_19511,N_19300);
or U20327 (N_20327,N_19537,N_19512);
nand U20328 (N_20328,N_19500,N_19472);
and U20329 (N_20329,N_19856,N_19739);
or U20330 (N_20330,N_19446,N_19578);
nand U20331 (N_20331,N_19087,N_19783);
or U20332 (N_20332,N_19646,N_19676);
xnor U20333 (N_20333,N_19575,N_19096);
and U20334 (N_20334,N_19244,N_19280);
or U20335 (N_20335,N_19476,N_19302);
or U20336 (N_20336,N_19665,N_19200);
or U20337 (N_20337,N_19406,N_19378);
and U20338 (N_20338,N_19380,N_19971);
or U20339 (N_20339,N_19584,N_19844);
nand U20340 (N_20340,N_19819,N_19020);
xnor U20341 (N_20341,N_19569,N_19965);
xor U20342 (N_20342,N_19042,N_19151);
xnor U20343 (N_20343,N_19003,N_19951);
and U20344 (N_20344,N_19106,N_19873);
nor U20345 (N_20345,N_19980,N_19722);
nand U20346 (N_20346,N_19123,N_19354);
nor U20347 (N_20347,N_19159,N_19287);
xnor U20348 (N_20348,N_19556,N_19482);
nor U20349 (N_20349,N_19847,N_19854);
or U20350 (N_20350,N_19304,N_19326);
xnor U20351 (N_20351,N_19754,N_19507);
or U20352 (N_20352,N_19281,N_19118);
nor U20353 (N_20353,N_19036,N_19738);
xor U20354 (N_20354,N_19669,N_19845);
and U20355 (N_20355,N_19828,N_19061);
xor U20356 (N_20356,N_19863,N_19282);
and U20357 (N_20357,N_19668,N_19059);
or U20358 (N_20358,N_19459,N_19037);
xnor U20359 (N_20359,N_19262,N_19166);
and U20360 (N_20360,N_19531,N_19883);
xnor U20361 (N_20361,N_19137,N_19853);
nor U20362 (N_20362,N_19846,N_19494);
and U20363 (N_20363,N_19127,N_19078);
nand U20364 (N_20364,N_19170,N_19831);
nor U20365 (N_20365,N_19211,N_19509);
nand U20366 (N_20366,N_19701,N_19091);
xor U20367 (N_20367,N_19296,N_19327);
or U20368 (N_20368,N_19158,N_19580);
nand U20369 (N_20369,N_19534,N_19877);
xnor U20370 (N_20370,N_19259,N_19254);
or U20371 (N_20371,N_19069,N_19615);
nor U20372 (N_20372,N_19986,N_19043);
or U20373 (N_20373,N_19717,N_19449);
xnor U20374 (N_20374,N_19315,N_19813);
nor U20375 (N_20375,N_19023,N_19134);
xor U20376 (N_20376,N_19097,N_19331);
or U20377 (N_20377,N_19601,N_19773);
nand U20378 (N_20378,N_19077,N_19344);
or U20379 (N_20379,N_19308,N_19501);
nor U20380 (N_20380,N_19497,N_19670);
nor U20381 (N_20381,N_19632,N_19903);
or U20382 (N_20382,N_19391,N_19247);
or U20383 (N_20383,N_19063,N_19599);
or U20384 (N_20384,N_19585,N_19943);
nor U20385 (N_20385,N_19150,N_19887);
or U20386 (N_20386,N_19718,N_19101);
xnor U20387 (N_20387,N_19781,N_19880);
and U20388 (N_20388,N_19057,N_19133);
and U20389 (N_20389,N_19143,N_19463);
nor U20390 (N_20390,N_19437,N_19953);
nor U20391 (N_20391,N_19999,N_19454);
and U20392 (N_20392,N_19829,N_19809);
xor U20393 (N_20393,N_19862,N_19957);
and U20394 (N_20394,N_19723,N_19876);
or U20395 (N_20395,N_19024,N_19841);
or U20396 (N_20396,N_19084,N_19241);
or U20397 (N_20397,N_19374,N_19260);
and U20398 (N_20398,N_19429,N_19923);
or U20399 (N_20399,N_19245,N_19600);
xnor U20400 (N_20400,N_19732,N_19525);
nor U20401 (N_20401,N_19466,N_19021);
nor U20402 (N_20402,N_19936,N_19222);
nor U20403 (N_20403,N_19539,N_19997);
nor U20404 (N_20404,N_19931,N_19076);
nor U20405 (N_20405,N_19650,N_19142);
xor U20406 (N_20406,N_19189,N_19226);
xor U20407 (N_20407,N_19410,N_19671);
and U20408 (N_20408,N_19228,N_19796);
nor U20409 (N_20409,N_19940,N_19242);
or U20410 (N_20410,N_19066,N_19227);
nor U20411 (N_20411,N_19566,N_19663);
nor U20412 (N_20412,N_19915,N_19205);
and U20413 (N_20413,N_19390,N_19926);
xor U20414 (N_20414,N_19152,N_19932);
xnor U20415 (N_20415,N_19471,N_19945);
nand U20416 (N_20416,N_19769,N_19734);
xnor U20417 (N_20417,N_19473,N_19896);
nand U20418 (N_20418,N_19484,N_19788);
xnor U20419 (N_20419,N_19598,N_19248);
nand U20420 (N_20420,N_19817,N_19113);
and U20421 (N_20421,N_19415,N_19164);
or U20422 (N_20422,N_19700,N_19707);
nand U20423 (N_20423,N_19389,N_19638);
nand U20424 (N_20424,N_19046,N_19129);
or U20425 (N_20425,N_19398,N_19206);
nand U20426 (N_20426,N_19567,N_19546);
xnor U20427 (N_20427,N_19464,N_19848);
and U20428 (N_20428,N_19870,N_19236);
or U20429 (N_20429,N_19099,N_19803);
xnor U20430 (N_20430,N_19747,N_19305);
and U20431 (N_20431,N_19832,N_19333);
and U20432 (N_20432,N_19927,N_19570);
nand U20433 (N_20433,N_19359,N_19452);
nor U20434 (N_20434,N_19377,N_19645);
xnor U20435 (N_20435,N_19545,N_19313);
nor U20436 (N_20436,N_19695,N_19529);
nor U20437 (N_20437,N_19770,N_19852);
nand U20438 (N_20438,N_19899,N_19583);
xor U20439 (N_20439,N_19523,N_19318);
nor U20440 (N_20440,N_19184,N_19403);
or U20441 (N_20441,N_19405,N_19030);
and U20442 (N_20442,N_19692,N_19461);
nand U20443 (N_20443,N_19175,N_19108);
or U20444 (N_20444,N_19532,N_19013);
xor U20445 (N_20445,N_19616,N_19083);
and U20446 (N_20446,N_19311,N_19934);
xnor U20447 (N_20447,N_19549,N_19250);
xnor U20448 (N_20448,N_19678,N_19443);
or U20449 (N_20449,N_19413,N_19375);
xnor U20450 (N_20450,N_19693,N_19995);
nor U20451 (N_20451,N_19592,N_19579);
nand U20452 (N_20452,N_19491,N_19130);
and U20453 (N_20453,N_19725,N_19070);
or U20454 (N_20454,N_19885,N_19149);
nor U20455 (N_20455,N_19603,N_19303);
nor U20456 (N_20456,N_19329,N_19805);
or U20457 (N_20457,N_19074,N_19629);
or U20458 (N_20458,N_19610,N_19879);
nand U20459 (N_20459,N_19330,N_19533);
or U20460 (N_20460,N_19336,N_19921);
and U20461 (N_20461,N_19974,N_19968);
xor U20462 (N_20462,N_19786,N_19937);
nor U20463 (N_20463,N_19574,N_19105);
nand U20464 (N_20464,N_19383,N_19120);
nor U20465 (N_20465,N_19542,N_19408);
and U20466 (N_20466,N_19618,N_19982);
or U20467 (N_20467,N_19955,N_19093);
xnor U20468 (N_20468,N_19991,N_19672);
nand U20469 (N_20469,N_19345,N_19726);
nand U20470 (N_20470,N_19655,N_19679);
nand U20471 (N_20471,N_19572,N_19427);
nor U20472 (N_20472,N_19234,N_19445);
nor U20473 (N_20473,N_19686,N_19713);
and U20474 (N_20474,N_19116,N_19706);
xnor U20475 (N_20475,N_19617,N_19963);
nor U20476 (N_20476,N_19611,N_19614);
nor U20477 (N_20477,N_19865,N_19952);
nor U20478 (N_20478,N_19520,N_19058);
and U20479 (N_20479,N_19992,N_19871);
xnor U20480 (N_20480,N_19636,N_19790);
or U20481 (N_20481,N_19820,N_19089);
or U20482 (N_20482,N_19555,N_19029);
nand U20483 (N_20483,N_19223,N_19363);
nor U20484 (N_20484,N_19285,N_19708);
nand U20485 (N_20485,N_19419,N_19536);
nand U20486 (N_20486,N_19631,N_19396);
and U20487 (N_20487,N_19425,N_19386);
or U20488 (N_20488,N_19480,N_19418);
xor U20489 (N_20489,N_19866,N_19696);
xnor U20490 (N_20490,N_19355,N_19891);
xnor U20491 (N_20491,N_19307,N_19185);
nor U20492 (N_20492,N_19444,N_19060);
xnor U20493 (N_20493,N_19776,N_19838);
or U20494 (N_20494,N_19740,N_19179);
xor U20495 (N_20495,N_19012,N_19808);
xor U20496 (N_20496,N_19697,N_19008);
nor U20497 (N_20497,N_19098,N_19071);
xnor U20498 (N_20498,N_19949,N_19544);
xnor U20499 (N_20499,N_19751,N_19827);
xor U20500 (N_20500,N_19395,N_19725);
xor U20501 (N_20501,N_19917,N_19691);
xnor U20502 (N_20502,N_19063,N_19898);
xnor U20503 (N_20503,N_19993,N_19429);
or U20504 (N_20504,N_19285,N_19566);
xnor U20505 (N_20505,N_19968,N_19988);
or U20506 (N_20506,N_19584,N_19518);
xnor U20507 (N_20507,N_19343,N_19062);
nand U20508 (N_20508,N_19561,N_19163);
nor U20509 (N_20509,N_19583,N_19033);
nand U20510 (N_20510,N_19605,N_19062);
nor U20511 (N_20511,N_19404,N_19719);
and U20512 (N_20512,N_19134,N_19773);
xor U20513 (N_20513,N_19756,N_19560);
xor U20514 (N_20514,N_19945,N_19135);
or U20515 (N_20515,N_19054,N_19803);
or U20516 (N_20516,N_19074,N_19767);
or U20517 (N_20517,N_19542,N_19535);
nor U20518 (N_20518,N_19625,N_19693);
nand U20519 (N_20519,N_19379,N_19859);
nand U20520 (N_20520,N_19960,N_19614);
or U20521 (N_20521,N_19886,N_19312);
nand U20522 (N_20522,N_19172,N_19823);
and U20523 (N_20523,N_19685,N_19745);
nor U20524 (N_20524,N_19319,N_19053);
or U20525 (N_20525,N_19530,N_19069);
and U20526 (N_20526,N_19671,N_19234);
xor U20527 (N_20527,N_19710,N_19636);
nor U20528 (N_20528,N_19293,N_19816);
nand U20529 (N_20529,N_19806,N_19132);
nor U20530 (N_20530,N_19836,N_19322);
xor U20531 (N_20531,N_19276,N_19769);
or U20532 (N_20532,N_19245,N_19909);
and U20533 (N_20533,N_19862,N_19863);
nand U20534 (N_20534,N_19988,N_19637);
xor U20535 (N_20535,N_19667,N_19095);
nor U20536 (N_20536,N_19877,N_19661);
and U20537 (N_20537,N_19266,N_19943);
or U20538 (N_20538,N_19270,N_19091);
nand U20539 (N_20539,N_19359,N_19614);
nor U20540 (N_20540,N_19327,N_19627);
nor U20541 (N_20541,N_19798,N_19973);
nand U20542 (N_20542,N_19011,N_19878);
nand U20543 (N_20543,N_19340,N_19639);
and U20544 (N_20544,N_19972,N_19766);
xnor U20545 (N_20545,N_19742,N_19676);
and U20546 (N_20546,N_19454,N_19401);
nand U20547 (N_20547,N_19089,N_19699);
nand U20548 (N_20548,N_19432,N_19262);
nand U20549 (N_20549,N_19881,N_19507);
nor U20550 (N_20550,N_19678,N_19354);
or U20551 (N_20551,N_19231,N_19850);
and U20552 (N_20552,N_19126,N_19963);
nand U20553 (N_20553,N_19552,N_19666);
or U20554 (N_20554,N_19797,N_19217);
xnor U20555 (N_20555,N_19996,N_19936);
nand U20556 (N_20556,N_19465,N_19959);
or U20557 (N_20557,N_19632,N_19997);
nor U20558 (N_20558,N_19309,N_19501);
and U20559 (N_20559,N_19244,N_19521);
and U20560 (N_20560,N_19492,N_19190);
nand U20561 (N_20561,N_19948,N_19752);
nor U20562 (N_20562,N_19159,N_19611);
nor U20563 (N_20563,N_19536,N_19556);
nand U20564 (N_20564,N_19237,N_19332);
or U20565 (N_20565,N_19406,N_19404);
xnor U20566 (N_20566,N_19583,N_19260);
and U20567 (N_20567,N_19176,N_19780);
xor U20568 (N_20568,N_19138,N_19380);
nor U20569 (N_20569,N_19081,N_19966);
nand U20570 (N_20570,N_19864,N_19374);
or U20571 (N_20571,N_19004,N_19386);
nor U20572 (N_20572,N_19091,N_19372);
nand U20573 (N_20573,N_19168,N_19028);
and U20574 (N_20574,N_19286,N_19664);
and U20575 (N_20575,N_19845,N_19835);
or U20576 (N_20576,N_19008,N_19742);
and U20577 (N_20577,N_19884,N_19098);
and U20578 (N_20578,N_19200,N_19524);
and U20579 (N_20579,N_19886,N_19313);
or U20580 (N_20580,N_19887,N_19394);
and U20581 (N_20581,N_19448,N_19046);
nand U20582 (N_20582,N_19212,N_19882);
and U20583 (N_20583,N_19318,N_19639);
and U20584 (N_20584,N_19405,N_19393);
or U20585 (N_20585,N_19235,N_19930);
and U20586 (N_20586,N_19319,N_19370);
nand U20587 (N_20587,N_19657,N_19139);
xor U20588 (N_20588,N_19444,N_19951);
nand U20589 (N_20589,N_19322,N_19488);
nand U20590 (N_20590,N_19016,N_19217);
xnor U20591 (N_20591,N_19531,N_19740);
nor U20592 (N_20592,N_19167,N_19816);
or U20593 (N_20593,N_19802,N_19852);
nor U20594 (N_20594,N_19308,N_19332);
xor U20595 (N_20595,N_19370,N_19354);
xor U20596 (N_20596,N_19441,N_19214);
xor U20597 (N_20597,N_19881,N_19620);
nand U20598 (N_20598,N_19590,N_19626);
and U20599 (N_20599,N_19102,N_19765);
nand U20600 (N_20600,N_19148,N_19208);
xnor U20601 (N_20601,N_19487,N_19611);
nor U20602 (N_20602,N_19517,N_19881);
nand U20603 (N_20603,N_19945,N_19487);
nor U20604 (N_20604,N_19662,N_19442);
nor U20605 (N_20605,N_19731,N_19930);
or U20606 (N_20606,N_19104,N_19365);
nor U20607 (N_20607,N_19441,N_19174);
or U20608 (N_20608,N_19094,N_19521);
xor U20609 (N_20609,N_19339,N_19597);
nand U20610 (N_20610,N_19675,N_19230);
or U20611 (N_20611,N_19862,N_19092);
nand U20612 (N_20612,N_19937,N_19797);
nand U20613 (N_20613,N_19375,N_19182);
nand U20614 (N_20614,N_19045,N_19668);
xor U20615 (N_20615,N_19789,N_19488);
nand U20616 (N_20616,N_19700,N_19144);
or U20617 (N_20617,N_19778,N_19908);
xnor U20618 (N_20618,N_19795,N_19567);
nor U20619 (N_20619,N_19240,N_19505);
or U20620 (N_20620,N_19145,N_19051);
or U20621 (N_20621,N_19128,N_19988);
nand U20622 (N_20622,N_19254,N_19560);
nor U20623 (N_20623,N_19412,N_19722);
and U20624 (N_20624,N_19262,N_19317);
or U20625 (N_20625,N_19795,N_19375);
nand U20626 (N_20626,N_19257,N_19178);
nand U20627 (N_20627,N_19590,N_19210);
or U20628 (N_20628,N_19188,N_19951);
nor U20629 (N_20629,N_19185,N_19790);
and U20630 (N_20630,N_19487,N_19485);
xor U20631 (N_20631,N_19522,N_19487);
or U20632 (N_20632,N_19530,N_19846);
xor U20633 (N_20633,N_19838,N_19258);
and U20634 (N_20634,N_19772,N_19887);
xor U20635 (N_20635,N_19079,N_19891);
xor U20636 (N_20636,N_19085,N_19350);
nor U20637 (N_20637,N_19477,N_19142);
nor U20638 (N_20638,N_19127,N_19295);
and U20639 (N_20639,N_19198,N_19256);
or U20640 (N_20640,N_19449,N_19461);
and U20641 (N_20641,N_19377,N_19259);
or U20642 (N_20642,N_19194,N_19760);
and U20643 (N_20643,N_19426,N_19402);
and U20644 (N_20644,N_19187,N_19160);
nor U20645 (N_20645,N_19493,N_19376);
and U20646 (N_20646,N_19232,N_19726);
or U20647 (N_20647,N_19896,N_19518);
and U20648 (N_20648,N_19190,N_19711);
and U20649 (N_20649,N_19962,N_19159);
nor U20650 (N_20650,N_19351,N_19706);
nor U20651 (N_20651,N_19966,N_19472);
xor U20652 (N_20652,N_19276,N_19337);
nand U20653 (N_20653,N_19937,N_19884);
xor U20654 (N_20654,N_19724,N_19923);
xor U20655 (N_20655,N_19350,N_19376);
and U20656 (N_20656,N_19967,N_19683);
and U20657 (N_20657,N_19413,N_19400);
xnor U20658 (N_20658,N_19867,N_19007);
nand U20659 (N_20659,N_19383,N_19333);
nor U20660 (N_20660,N_19865,N_19403);
and U20661 (N_20661,N_19846,N_19275);
or U20662 (N_20662,N_19564,N_19210);
or U20663 (N_20663,N_19446,N_19361);
or U20664 (N_20664,N_19988,N_19104);
xnor U20665 (N_20665,N_19723,N_19051);
nor U20666 (N_20666,N_19262,N_19679);
xor U20667 (N_20667,N_19388,N_19356);
nor U20668 (N_20668,N_19773,N_19690);
and U20669 (N_20669,N_19019,N_19436);
xor U20670 (N_20670,N_19658,N_19900);
or U20671 (N_20671,N_19065,N_19554);
and U20672 (N_20672,N_19955,N_19192);
nand U20673 (N_20673,N_19524,N_19612);
and U20674 (N_20674,N_19365,N_19391);
and U20675 (N_20675,N_19031,N_19891);
nor U20676 (N_20676,N_19269,N_19875);
nor U20677 (N_20677,N_19181,N_19120);
and U20678 (N_20678,N_19238,N_19404);
nor U20679 (N_20679,N_19103,N_19867);
nor U20680 (N_20680,N_19337,N_19694);
nor U20681 (N_20681,N_19888,N_19746);
xor U20682 (N_20682,N_19076,N_19933);
nor U20683 (N_20683,N_19543,N_19030);
nor U20684 (N_20684,N_19321,N_19649);
and U20685 (N_20685,N_19995,N_19575);
nand U20686 (N_20686,N_19397,N_19452);
xor U20687 (N_20687,N_19095,N_19251);
and U20688 (N_20688,N_19660,N_19700);
nand U20689 (N_20689,N_19061,N_19016);
nor U20690 (N_20690,N_19205,N_19792);
and U20691 (N_20691,N_19954,N_19591);
and U20692 (N_20692,N_19292,N_19541);
xnor U20693 (N_20693,N_19772,N_19055);
or U20694 (N_20694,N_19652,N_19699);
nand U20695 (N_20695,N_19734,N_19757);
nand U20696 (N_20696,N_19275,N_19479);
xnor U20697 (N_20697,N_19329,N_19966);
nand U20698 (N_20698,N_19118,N_19168);
and U20699 (N_20699,N_19274,N_19943);
xnor U20700 (N_20700,N_19761,N_19579);
and U20701 (N_20701,N_19579,N_19593);
nor U20702 (N_20702,N_19426,N_19310);
xnor U20703 (N_20703,N_19420,N_19662);
or U20704 (N_20704,N_19175,N_19478);
nor U20705 (N_20705,N_19299,N_19911);
nand U20706 (N_20706,N_19689,N_19967);
or U20707 (N_20707,N_19658,N_19742);
or U20708 (N_20708,N_19688,N_19313);
nor U20709 (N_20709,N_19777,N_19491);
nor U20710 (N_20710,N_19764,N_19207);
nand U20711 (N_20711,N_19280,N_19611);
nand U20712 (N_20712,N_19870,N_19559);
and U20713 (N_20713,N_19378,N_19673);
and U20714 (N_20714,N_19131,N_19926);
and U20715 (N_20715,N_19557,N_19717);
or U20716 (N_20716,N_19775,N_19931);
xnor U20717 (N_20717,N_19313,N_19887);
or U20718 (N_20718,N_19086,N_19167);
nand U20719 (N_20719,N_19898,N_19500);
nand U20720 (N_20720,N_19231,N_19530);
or U20721 (N_20721,N_19599,N_19640);
nor U20722 (N_20722,N_19511,N_19913);
nand U20723 (N_20723,N_19238,N_19555);
nor U20724 (N_20724,N_19469,N_19349);
nand U20725 (N_20725,N_19274,N_19537);
nor U20726 (N_20726,N_19416,N_19998);
and U20727 (N_20727,N_19646,N_19776);
nand U20728 (N_20728,N_19214,N_19413);
nor U20729 (N_20729,N_19547,N_19512);
nand U20730 (N_20730,N_19362,N_19940);
or U20731 (N_20731,N_19049,N_19689);
nand U20732 (N_20732,N_19453,N_19199);
nor U20733 (N_20733,N_19336,N_19316);
xor U20734 (N_20734,N_19148,N_19032);
or U20735 (N_20735,N_19283,N_19328);
and U20736 (N_20736,N_19204,N_19855);
nor U20737 (N_20737,N_19955,N_19892);
nor U20738 (N_20738,N_19370,N_19489);
nand U20739 (N_20739,N_19208,N_19296);
and U20740 (N_20740,N_19692,N_19407);
or U20741 (N_20741,N_19715,N_19104);
or U20742 (N_20742,N_19243,N_19474);
nand U20743 (N_20743,N_19897,N_19959);
nand U20744 (N_20744,N_19958,N_19088);
or U20745 (N_20745,N_19787,N_19126);
nor U20746 (N_20746,N_19377,N_19814);
and U20747 (N_20747,N_19862,N_19547);
nor U20748 (N_20748,N_19711,N_19035);
xor U20749 (N_20749,N_19944,N_19039);
xnor U20750 (N_20750,N_19741,N_19577);
xnor U20751 (N_20751,N_19509,N_19612);
nor U20752 (N_20752,N_19496,N_19270);
xor U20753 (N_20753,N_19839,N_19699);
or U20754 (N_20754,N_19239,N_19691);
or U20755 (N_20755,N_19142,N_19015);
nand U20756 (N_20756,N_19372,N_19968);
xor U20757 (N_20757,N_19575,N_19275);
or U20758 (N_20758,N_19426,N_19791);
or U20759 (N_20759,N_19747,N_19344);
nor U20760 (N_20760,N_19297,N_19896);
nor U20761 (N_20761,N_19674,N_19185);
nor U20762 (N_20762,N_19703,N_19303);
xnor U20763 (N_20763,N_19817,N_19627);
nand U20764 (N_20764,N_19232,N_19932);
and U20765 (N_20765,N_19027,N_19500);
xnor U20766 (N_20766,N_19454,N_19131);
and U20767 (N_20767,N_19722,N_19656);
nand U20768 (N_20768,N_19321,N_19188);
nand U20769 (N_20769,N_19429,N_19724);
nor U20770 (N_20770,N_19486,N_19609);
and U20771 (N_20771,N_19624,N_19890);
or U20772 (N_20772,N_19499,N_19084);
nor U20773 (N_20773,N_19563,N_19344);
xor U20774 (N_20774,N_19396,N_19208);
or U20775 (N_20775,N_19601,N_19452);
and U20776 (N_20776,N_19070,N_19480);
and U20777 (N_20777,N_19789,N_19871);
and U20778 (N_20778,N_19825,N_19414);
and U20779 (N_20779,N_19624,N_19974);
nand U20780 (N_20780,N_19882,N_19002);
or U20781 (N_20781,N_19358,N_19199);
and U20782 (N_20782,N_19618,N_19599);
nand U20783 (N_20783,N_19477,N_19605);
nand U20784 (N_20784,N_19908,N_19162);
xnor U20785 (N_20785,N_19649,N_19048);
or U20786 (N_20786,N_19093,N_19942);
xor U20787 (N_20787,N_19788,N_19722);
or U20788 (N_20788,N_19608,N_19328);
and U20789 (N_20789,N_19235,N_19981);
nor U20790 (N_20790,N_19145,N_19182);
or U20791 (N_20791,N_19882,N_19447);
nor U20792 (N_20792,N_19270,N_19884);
or U20793 (N_20793,N_19758,N_19745);
xnor U20794 (N_20794,N_19442,N_19973);
and U20795 (N_20795,N_19813,N_19730);
nor U20796 (N_20796,N_19209,N_19051);
or U20797 (N_20797,N_19022,N_19089);
xor U20798 (N_20798,N_19420,N_19517);
nand U20799 (N_20799,N_19058,N_19801);
xnor U20800 (N_20800,N_19758,N_19150);
nand U20801 (N_20801,N_19526,N_19892);
and U20802 (N_20802,N_19238,N_19284);
nand U20803 (N_20803,N_19285,N_19189);
nand U20804 (N_20804,N_19042,N_19345);
and U20805 (N_20805,N_19726,N_19439);
or U20806 (N_20806,N_19162,N_19783);
and U20807 (N_20807,N_19881,N_19700);
nand U20808 (N_20808,N_19162,N_19350);
nand U20809 (N_20809,N_19826,N_19267);
xnor U20810 (N_20810,N_19008,N_19956);
or U20811 (N_20811,N_19047,N_19778);
or U20812 (N_20812,N_19782,N_19889);
and U20813 (N_20813,N_19309,N_19490);
nand U20814 (N_20814,N_19039,N_19720);
nand U20815 (N_20815,N_19662,N_19130);
xnor U20816 (N_20816,N_19844,N_19482);
nand U20817 (N_20817,N_19894,N_19053);
or U20818 (N_20818,N_19416,N_19658);
or U20819 (N_20819,N_19239,N_19929);
nor U20820 (N_20820,N_19243,N_19994);
nor U20821 (N_20821,N_19224,N_19569);
or U20822 (N_20822,N_19339,N_19086);
xnor U20823 (N_20823,N_19333,N_19502);
xnor U20824 (N_20824,N_19302,N_19879);
nor U20825 (N_20825,N_19474,N_19595);
xnor U20826 (N_20826,N_19502,N_19398);
nor U20827 (N_20827,N_19725,N_19066);
or U20828 (N_20828,N_19430,N_19792);
xnor U20829 (N_20829,N_19239,N_19627);
xnor U20830 (N_20830,N_19713,N_19408);
nor U20831 (N_20831,N_19026,N_19341);
nand U20832 (N_20832,N_19641,N_19700);
nand U20833 (N_20833,N_19762,N_19637);
or U20834 (N_20834,N_19485,N_19176);
xor U20835 (N_20835,N_19406,N_19256);
or U20836 (N_20836,N_19208,N_19964);
nand U20837 (N_20837,N_19131,N_19677);
nor U20838 (N_20838,N_19229,N_19118);
nor U20839 (N_20839,N_19786,N_19169);
nor U20840 (N_20840,N_19885,N_19808);
nand U20841 (N_20841,N_19310,N_19716);
and U20842 (N_20842,N_19043,N_19635);
nand U20843 (N_20843,N_19057,N_19606);
or U20844 (N_20844,N_19150,N_19090);
xnor U20845 (N_20845,N_19545,N_19860);
nand U20846 (N_20846,N_19312,N_19099);
nor U20847 (N_20847,N_19039,N_19375);
or U20848 (N_20848,N_19529,N_19604);
nor U20849 (N_20849,N_19956,N_19259);
xnor U20850 (N_20850,N_19023,N_19153);
and U20851 (N_20851,N_19022,N_19379);
and U20852 (N_20852,N_19525,N_19235);
nand U20853 (N_20853,N_19564,N_19134);
nand U20854 (N_20854,N_19180,N_19286);
or U20855 (N_20855,N_19910,N_19506);
xnor U20856 (N_20856,N_19267,N_19202);
xor U20857 (N_20857,N_19973,N_19250);
xnor U20858 (N_20858,N_19911,N_19744);
xnor U20859 (N_20859,N_19921,N_19050);
xor U20860 (N_20860,N_19779,N_19802);
nor U20861 (N_20861,N_19200,N_19890);
xor U20862 (N_20862,N_19123,N_19672);
nand U20863 (N_20863,N_19877,N_19225);
nor U20864 (N_20864,N_19159,N_19815);
xnor U20865 (N_20865,N_19577,N_19928);
and U20866 (N_20866,N_19525,N_19002);
or U20867 (N_20867,N_19947,N_19661);
xor U20868 (N_20868,N_19044,N_19171);
xnor U20869 (N_20869,N_19045,N_19043);
nand U20870 (N_20870,N_19553,N_19210);
nor U20871 (N_20871,N_19159,N_19426);
xnor U20872 (N_20872,N_19577,N_19626);
or U20873 (N_20873,N_19129,N_19043);
nand U20874 (N_20874,N_19816,N_19032);
nor U20875 (N_20875,N_19212,N_19922);
or U20876 (N_20876,N_19652,N_19733);
and U20877 (N_20877,N_19247,N_19999);
and U20878 (N_20878,N_19158,N_19387);
nand U20879 (N_20879,N_19603,N_19597);
nor U20880 (N_20880,N_19680,N_19362);
xor U20881 (N_20881,N_19766,N_19164);
nand U20882 (N_20882,N_19398,N_19807);
or U20883 (N_20883,N_19585,N_19962);
and U20884 (N_20884,N_19446,N_19187);
xor U20885 (N_20885,N_19766,N_19613);
nor U20886 (N_20886,N_19125,N_19617);
or U20887 (N_20887,N_19089,N_19362);
and U20888 (N_20888,N_19807,N_19933);
or U20889 (N_20889,N_19947,N_19641);
nor U20890 (N_20890,N_19546,N_19797);
and U20891 (N_20891,N_19297,N_19237);
nand U20892 (N_20892,N_19802,N_19135);
nand U20893 (N_20893,N_19792,N_19811);
and U20894 (N_20894,N_19867,N_19288);
xor U20895 (N_20895,N_19980,N_19075);
and U20896 (N_20896,N_19615,N_19925);
nand U20897 (N_20897,N_19051,N_19822);
or U20898 (N_20898,N_19325,N_19416);
xnor U20899 (N_20899,N_19996,N_19316);
nand U20900 (N_20900,N_19544,N_19189);
and U20901 (N_20901,N_19075,N_19448);
and U20902 (N_20902,N_19562,N_19332);
and U20903 (N_20903,N_19894,N_19145);
nand U20904 (N_20904,N_19691,N_19766);
and U20905 (N_20905,N_19776,N_19131);
nor U20906 (N_20906,N_19454,N_19888);
nor U20907 (N_20907,N_19936,N_19061);
nand U20908 (N_20908,N_19340,N_19427);
and U20909 (N_20909,N_19422,N_19199);
nor U20910 (N_20910,N_19193,N_19220);
and U20911 (N_20911,N_19150,N_19072);
nand U20912 (N_20912,N_19519,N_19366);
or U20913 (N_20913,N_19612,N_19282);
xnor U20914 (N_20914,N_19205,N_19267);
nand U20915 (N_20915,N_19100,N_19025);
and U20916 (N_20916,N_19558,N_19102);
and U20917 (N_20917,N_19259,N_19917);
and U20918 (N_20918,N_19590,N_19939);
and U20919 (N_20919,N_19084,N_19928);
nor U20920 (N_20920,N_19394,N_19692);
or U20921 (N_20921,N_19685,N_19516);
xor U20922 (N_20922,N_19624,N_19884);
and U20923 (N_20923,N_19994,N_19932);
or U20924 (N_20924,N_19662,N_19032);
nand U20925 (N_20925,N_19481,N_19355);
and U20926 (N_20926,N_19479,N_19470);
xor U20927 (N_20927,N_19272,N_19099);
or U20928 (N_20928,N_19092,N_19210);
nor U20929 (N_20929,N_19143,N_19479);
nand U20930 (N_20930,N_19332,N_19388);
nor U20931 (N_20931,N_19578,N_19251);
and U20932 (N_20932,N_19963,N_19809);
and U20933 (N_20933,N_19111,N_19326);
xor U20934 (N_20934,N_19051,N_19817);
and U20935 (N_20935,N_19186,N_19574);
nand U20936 (N_20936,N_19862,N_19235);
nand U20937 (N_20937,N_19698,N_19358);
or U20938 (N_20938,N_19657,N_19368);
nor U20939 (N_20939,N_19036,N_19296);
or U20940 (N_20940,N_19511,N_19759);
nor U20941 (N_20941,N_19319,N_19062);
xor U20942 (N_20942,N_19534,N_19055);
nor U20943 (N_20943,N_19448,N_19313);
xor U20944 (N_20944,N_19697,N_19810);
nand U20945 (N_20945,N_19641,N_19694);
xnor U20946 (N_20946,N_19788,N_19250);
or U20947 (N_20947,N_19812,N_19204);
or U20948 (N_20948,N_19734,N_19929);
or U20949 (N_20949,N_19352,N_19327);
nor U20950 (N_20950,N_19843,N_19642);
xor U20951 (N_20951,N_19106,N_19383);
xnor U20952 (N_20952,N_19223,N_19206);
or U20953 (N_20953,N_19566,N_19894);
nand U20954 (N_20954,N_19127,N_19916);
nand U20955 (N_20955,N_19516,N_19249);
or U20956 (N_20956,N_19036,N_19429);
nor U20957 (N_20957,N_19811,N_19635);
nand U20958 (N_20958,N_19464,N_19430);
and U20959 (N_20959,N_19459,N_19669);
and U20960 (N_20960,N_19338,N_19578);
xor U20961 (N_20961,N_19246,N_19563);
nor U20962 (N_20962,N_19196,N_19703);
and U20963 (N_20963,N_19916,N_19497);
and U20964 (N_20964,N_19532,N_19172);
xnor U20965 (N_20965,N_19796,N_19011);
xnor U20966 (N_20966,N_19628,N_19559);
nor U20967 (N_20967,N_19318,N_19890);
xnor U20968 (N_20968,N_19076,N_19669);
nor U20969 (N_20969,N_19831,N_19983);
nand U20970 (N_20970,N_19525,N_19114);
and U20971 (N_20971,N_19529,N_19721);
xor U20972 (N_20972,N_19559,N_19337);
nand U20973 (N_20973,N_19944,N_19131);
or U20974 (N_20974,N_19874,N_19484);
or U20975 (N_20975,N_19744,N_19586);
or U20976 (N_20976,N_19049,N_19640);
nand U20977 (N_20977,N_19998,N_19578);
nand U20978 (N_20978,N_19317,N_19015);
nor U20979 (N_20979,N_19703,N_19601);
nand U20980 (N_20980,N_19395,N_19089);
xor U20981 (N_20981,N_19378,N_19576);
and U20982 (N_20982,N_19402,N_19131);
xnor U20983 (N_20983,N_19589,N_19213);
nand U20984 (N_20984,N_19430,N_19345);
and U20985 (N_20985,N_19612,N_19872);
and U20986 (N_20986,N_19574,N_19745);
nand U20987 (N_20987,N_19196,N_19388);
or U20988 (N_20988,N_19905,N_19285);
nor U20989 (N_20989,N_19631,N_19205);
nand U20990 (N_20990,N_19138,N_19947);
nor U20991 (N_20991,N_19616,N_19261);
nor U20992 (N_20992,N_19642,N_19276);
nor U20993 (N_20993,N_19542,N_19118);
nor U20994 (N_20994,N_19800,N_19096);
and U20995 (N_20995,N_19135,N_19445);
nand U20996 (N_20996,N_19929,N_19361);
xnor U20997 (N_20997,N_19301,N_19969);
nor U20998 (N_20998,N_19162,N_19116);
or U20999 (N_20999,N_19867,N_19514);
xnor U21000 (N_21000,N_20926,N_20737);
nand U21001 (N_21001,N_20488,N_20710);
and U21002 (N_21002,N_20694,N_20681);
xnor U21003 (N_21003,N_20650,N_20670);
xnor U21004 (N_21004,N_20143,N_20350);
nand U21005 (N_21005,N_20547,N_20351);
nand U21006 (N_21006,N_20044,N_20025);
xnor U21007 (N_21007,N_20930,N_20882);
nand U21008 (N_21008,N_20968,N_20908);
and U21009 (N_21009,N_20022,N_20580);
and U21010 (N_21010,N_20951,N_20712);
and U21011 (N_21011,N_20303,N_20080);
xnor U21012 (N_21012,N_20414,N_20395);
nor U21013 (N_21013,N_20765,N_20452);
nor U21014 (N_21014,N_20188,N_20886);
xnor U21015 (N_21015,N_20029,N_20090);
xor U21016 (N_21016,N_20625,N_20128);
and U21017 (N_21017,N_20788,N_20995);
and U21018 (N_21018,N_20654,N_20286);
xor U21019 (N_21019,N_20552,N_20457);
and U21020 (N_21020,N_20219,N_20170);
or U21021 (N_21021,N_20049,N_20535);
nand U21022 (N_21022,N_20876,N_20508);
or U21023 (N_21023,N_20119,N_20083);
xnor U21024 (N_21024,N_20730,N_20655);
nand U21025 (N_21025,N_20904,N_20549);
nor U21026 (N_21026,N_20568,N_20370);
nor U21027 (N_21027,N_20852,N_20036);
nand U21028 (N_21028,N_20894,N_20880);
nor U21029 (N_21029,N_20829,N_20111);
nand U21030 (N_21030,N_20726,N_20125);
xor U21031 (N_21031,N_20622,N_20074);
or U21032 (N_21032,N_20872,N_20653);
xor U21033 (N_21033,N_20828,N_20636);
or U21034 (N_21034,N_20548,N_20984);
nor U21035 (N_21035,N_20129,N_20330);
nor U21036 (N_21036,N_20838,N_20861);
nand U21037 (N_21037,N_20084,N_20259);
xor U21038 (N_21038,N_20200,N_20898);
or U21039 (N_21039,N_20952,N_20152);
nand U21040 (N_21040,N_20742,N_20344);
xor U21041 (N_21041,N_20629,N_20062);
and U21042 (N_21042,N_20624,N_20678);
or U21043 (N_21043,N_20999,N_20638);
or U21044 (N_21044,N_20393,N_20224);
nand U21045 (N_21045,N_20635,N_20486);
nor U21046 (N_21046,N_20236,N_20179);
xor U21047 (N_21047,N_20379,N_20656);
and U21048 (N_21048,N_20682,N_20177);
or U21049 (N_21049,N_20273,N_20251);
nor U21050 (N_21050,N_20100,N_20498);
nand U21051 (N_21051,N_20600,N_20927);
and U21052 (N_21052,N_20359,N_20247);
xnor U21053 (N_21053,N_20896,N_20182);
nor U21054 (N_21054,N_20348,N_20504);
xnor U21055 (N_21055,N_20139,N_20309);
nand U21056 (N_21056,N_20711,N_20147);
and U21057 (N_21057,N_20342,N_20963);
nand U21058 (N_21058,N_20263,N_20523);
and U21059 (N_21059,N_20881,N_20832);
nor U21060 (N_21060,N_20464,N_20287);
xor U21061 (N_21061,N_20162,N_20870);
nor U21062 (N_21062,N_20060,N_20643);
nor U21063 (N_21063,N_20284,N_20437);
and U21064 (N_21064,N_20094,N_20248);
nor U21065 (N_21065,N_20764,N_20198);
xnor U21066 (N_21066,N_20133,N_20028);
nand U21067 (N_21067,N_20264,N_20441);
nand U21068 (N_21068,N_20567,N_20992);
xnor U21069 (N_21069,N_20993,N_20631);
or U21070 (N_21070,N_20146,N_20641);
nand U21071 (N_21071,N_20132,N_20740);
nor U21072 (N_21072,N_20315,N_20061);
nand U21073 (N_21073,N_20810,N_20722);
or U21074 (N_21074,N_20959,N_20749);
xnor U21075 (N_21075,N_20483,N_20990);
nand U21076 (N_21076,N_20561,N_20860);
and U21077 (N_21077,N_20250,N_20554);
nand U21078 (N_21078,N_20845,N_20501);
nor U21079 (N_21079,N_20478,N_20557);
or U21080 (N_21080,N_20467,N_20418);
xor U21081 (N_21081,N_20759,N_20801);
and U21082 (N_21082,N_20958,N_20203);
nor U21083 (N_21083,N_20704,N_20648);
xor U21084 (N_21084,N_20897,N_20607);
nand U21085 (N_21085,N_20169,N_20277);
nand U21086 (N_21086,N_20874,N_20098);
and U21087 (N_21087,N_20687,N_20447);
xnor U21088 (N_21088,N_20269,N_20782);
nand U21089 (N_21089,N_20888,N_20695);
xor U21090 (N_21090,N_20307,N_20043);
and U21091 (N_21091,N_20421,N_20879);
nand U21092 (N_21092,N_20525,N_20242);
nand U21093 (N_21093,N_20649,N_20619);
or U21094 (N_21094,N_20366,N_20374);
or U21095 (N_21095,N_20050,N_20774);
and U21096 (N_21096,N_20652,N_20675);
nand U21097 (N_21097,N_20538,N_20118);
xnor U21098 (N_21098,N_20982,N_20308);
and U21099 (N_21099,N_20956,N_20067);
or U21100 (N_21100,N_20101,N_20015);
or U21101 (N_21101,N_20750,N_20208);
xnor U21102 (N_21102,N_20240,N_20667);
or U21103 (N_21103,N_20239,N_20728);
and U21104 (N_21104,N_20425,N_20037);
and U21105 (N_21105,N_20617,N_20697);
xor U21106 (N_21106,N_20637,N_20787);
xor U21107 (N_21107,N_20230,N_20592);
and U21108 (N_21108,N_20856,N_20474);
nand U21109 (N_21109,N_20327,N_20966);
nor U21110 (N_21110,N_20804,N_20326);
or U21111 (N_21111,N_20705,N_20046);
or U21112 (N_21112,N_20954,N_20955);
and U21113 (N_21113,N_20201,N_20252);
and U21114 (N_21114,N_20127,N_20521);
and U21115 (N_21115,N_20850,N_20791);
nand U21116 (N_21116,N_20254,N_20701);
or U21117 (N_21117,N_20500,N_20371);
nand U21118 (N_21118,N_20068,N_20871);
xnor U21119 (N_21119,N_20581,N_20003);
xnor U21120 (N_21120,N_20092,N_20495);
nand U21121 (N_21121,N_20276,N_20988);
xor U21122 (N_21122,N_20399,N_20794);
xnor U21123 (N_21123,N_20925,N_20082);
nor U21124 (N_21124,N_20628,N_20411);
and U21125 (N_21125,N_20356,N_20962);
and U21126 (N_21126,N_20391,N_20205);
or U21127 (N_21127,N_20964,N_20477);
nand U21128 (N_21128,N_20747,N_20070);
xor U21129 (N_21129,N_20633,N_20442);
nor U21130 (N_21130,N_20940,N_20081);
or U21131 (N_21131,N_20427,N_20559);
nand U21132 (N_21132,N_20974,N_20479);
xor U21133 (N_21133,N_20555,N_20134);
xor U21134 (N_21134,N_20151,N_20258);
nand U21135 (N_21135,N_20748,N_20931);
nand U21136 (N_21136,N_20953,N_20338);
or U21137 (N_21137,N_20302,N_20145);
and U21138 (N_21138,N_20822,N_20154);
or U21139 (N_21139,N_20382,N_20294);
and U21140 (N_21140,N_20187,N_20432);
and U21141 (N_21141,N_20531,N_20126);
nand U21142 (N_21142,N_20965,N_20657);
xnor U21143 (N_21143,N_20980,N_20784);
or U21144 (N_21144,N_20497,N_20144);
xor U21145 (N_21145,N_20325,N_20833);
or U21146 (N_21146,N_20196,N_20367);
or U21147 (N_21147,N_20117,N_20602);
nand U21148 (N_21148,N_20830,N_20720);
xor U21149 (N_21149,N_20715,N_20175);
nand U21150 (N_21150,N_20570,N_20862);
or U21151 (N_21151,N_20934,N_20013);
and U21152 (N_21152,N_20033,N_20916);
xnor U21153 (N_21153,N_20550,N_20413);
xnor U21154 (N_21154,N_20642,N_20016);
xor U21155 (N_21155,N_20257,N_20770);
nor U21156 (N_21156,N_20085,N_20903);
or U21157 (N_21157,N_20292,N_20053);
and U21158 (N_21158,N_20313,N_20481);
and U21159 (N_21159,N_20579,N_20466);
and U21160 (N_21160,N_20725,N_20912);
or U21161 (N_21161,N_20422,N_20582);
or U21162 (N_21162,N_20390,N_20223);
xnor U21163 (N_21163,N_20340,N_20910);
or U21164 (N_21164,N_20578,N_20972);
or U21165 (N_21165,N_20676,N_20855);
xor U21166 (N_21166,N_20210,N_20989);
and U21167 (N_21167,N_20458,N_20091);
nand U21168 (N_21168,N_20847,N_20797);
or U21169 (N_21169,N_20489,N_20807);
and U21170 (N_21170,N_20666,N_20598);
and U21171 (N_21171,N_20394,N_20562);
and U21172 (N_21172,N_20777,N_20361);
xnor U21173 (N_21173,N_20064,N_20795);
or U21174 (N_21174,N_20480,N_20517);
nand U21175 (N_21175,N_20433,N_20499);
nand U21176 (N_21176,N_20723,N_20270);
xor U21177 (N_21177,N_20793,N_20563);
nand U21178 (N_21178,N_20194,N_20757);
xnor U21179 (N_21179,N_20155,N_20335);
and U21180 (N_21180,N_20047,N_20751);
nand U21181 (N_21181,N_20265,N_20076);
or U21182 (N_21182,N_20560,N_20368);
nand U21183 (N_21183,N_20096,N_20227);
or U21184 (N_21184,N_20789,N_20255);
xnor U21185 (N_21185,N_20435,N_20410);
and U21186 (N_21186,N_20280,N_20848);
xnor U21187 (N_21187,N_20506,N_20456);
nor U21188 (N_21188,N_20213,N_20799);
or U21189 (N_21189,N_20986,N_20817);
nand U21190 (N_21190,N_20352,N_20305);
and U21191 (N_21191,N_20544,N_20796);
xnor U21192 (N_21192,N_20978,N_20174);
nand U21193 (N_21193,N_20802,N_20123);
and U21194 (N_21194,N_20431,N_20674);
or U21195 (N_21195,N_20272,N_20420);
nor U21196 (N_21196,N_20450,N_20318);
or U21197 (N_21197,N_20815,N_20661);
nand U21198 (N_21198,N_20983,N_20868);
or U21199 (N_21199,N_20032,N_20780);
nor U21200 (N_21200,N_20097,N_20785);
or U21201 (N_21201,N_20839,N_20148);
and U21202 (N_21202,N_20482,N_20189);
nand U21203 (N_21203,N_20403,N_20779);
xor U21204 (N_21204,N_20851,N_20513);
xor U21205 (N_21205,N_20824,N_20333);
nor U21206 (N_21206,N_20245,N_20002);
xnor U21207 (N_21207,N_20130,N_20599);
xnor U21208 (N_21208,N_20472,N_20436);
nand U21209 (N_21209,N_20669,N_20295);
nand U21210 (N_21210,N_20753,N_20553);
nand U21211 (N_21211,N_20238,N_20372);
xor U21212 (N_21212,N_20569,N_20768);
nand U21213 (N_21213,N_20416,N_20970);
nand U21214 (N_21214,N_20496,N_20719);
and U21215 (N_21215,N_20843,N_20734);
xor U21216 (N_21216,N_20319,N_20444);
nand U21217 (N_21217,N_20124,N_20938);
or U21218 (N_21218,N_20677,N_20645);
nor U21219 (N_21219,N_20296,N_20979);
nor U21220 (N_21220,N_20322,N_20994);
xnor U21221 (N_21221,N_20533,N_20102);
or U21222 (N_21222,N_20088,N_20738);
nand U21223 (N_21223,N_20866,N_20854);
xor U21224 (N_21224,N_20618,N_20805);
or U21225 (N_21225,N_20933,N_20221);
nor U21226 (N_21226,N_20271,N_20171);
nor U21227 (N_21227,N_20369,N_20688);
nor U21228 (N_21228,N_20543,N_20353);
and U21229 (N_21229,N_20329,N_20680);
nand U21230 (N_21230,N_20893,N_20355);
nor U21231 (N_21231,N_20626,N_20586);
nor U21232 (N_21232,N_20758,N_20150);
nor U21233 (N_21233,N_20929,N_20917);
nor U21234 (N_21234,N_20298,N_20463);
nand U21235 (N_21235,N_20505,N_20214);
xor U21236 (N_21236,N_20253,N_20228);
and U21237 (N_21237,N_20919,N_20998);
nand U21238 (N_21238,N_20494,N_20072);
and U21239 (N_21239,N_20363,N_20594);
and U21240 (N_21240,N_20991,N_20875);
xor U21241 (N_21241,N_20647,N_20587);
nor U21242 (N_21242,N_20008,N_20935);
nand U21243 (N_21243,N_20243,N_20591);
or U21244 (N_21244,N_20375,N_20840);
xor U21245 (N_21245,N_20961,N_20052);
and U21246 (N_21246,N_20942,N_20975);
and U21247 (N_21247,N_20244,N_20608);
nor U21248 (N_21248,N_20603,N_20469);
nor U21249 (N_21249,N_20138,N_20288);
nor U21250 (N_21250,N_20589,N_20057);
or U21251 (N_21251,N_20944,N_20609);
or U21252 (N_21252,N_20686,N_20529);
and U21253 (N_21253,N_20345,N_20160);
and U21254 (N_21254,N_20142,N_20923);
or U21255 (N_21255,N_20571,N_20341);
and U21256 (N_21256,N_20229,N_20588);
or U21257 (N_21257,N_20110,N_20009);
xnor U21258 (N_21258,N_20030,N_20261);
and U21259 (N_21259,N_20502,N_20842);
or U21260 (N_21260,N_20664,N_20527);
nor U21261 (N_21261,N_20167,N_20987);
xor U21262 (N_21262,N_20834,N_20107);
or U21263 (N_21263,N_20672,N_20443);
xnor U21264 (N_21264,N_20197,N_20109);
or U21265 (N_21265,N_20460,N_20721);
nor U21266 (N_21266,N_20180,N_20211);
nor U21267 (N_21267,N_20398,N_20204);
or U21268 (N_21268,N_20772,N_20545);
xnor U21269 (N_21269,N_20172,N_20823);
or U21270 (N_21270,N_20116,N_20163);
nand U21271 (N_21271,N_20706,N_20744);
nand U21272 (N_21272,N_20763,N_20428);
and U21273 (N_21273,N_20583,N_20684);
xnor U21274 (N_21274,N_20386,N_20274);
and U21275 (N_21275,N_20023,N_20515);
xor U21276 (N_21276,N_20606,N_20887);
xnor U21277 (N_21277,N_20818,N_20509);
or U21278 (N_21278,N_20546,N_20365);
xor U21279 (N_21279,N_20262,N_20424);
xnor U21280 (N_21280,N_20183,N_20027);
xor U21281 (N_21281,N_20114,N_20218);
and U21282 (N_21282,N_20536,N_20140);
or U21283 (N_21283,N_20756,N_20743);
nor U21284 (N_21284,N_20724,N_20440);
xor U21285 (N_21285,N_20007,N_20439);
nor U21286 (N_21286,N_20892,N_20191);
xnor U21287 (N_21287,N_20106,N_20212);
xor U21288 (N_21288,N_20312,N_20853);
nand U21289 (N_21289,N_20806,N_20453);
and U21290 (N_21290,N_20973,N_20528);
xnor U21291 (N_21291,N_20108,N_20291);
xnor U21292 (N_21292,N_20918,N_20066);
xnor U21293 (N_21293,N_20071,N_20914);
nor U21294 (N_21294,N_20937,N_20639);
nor U21295 (N_21295,N_20864,N_20299);
and U21296 (N_21296,N_20634,N_20304);
nor U21297 (N_21297,N_20819,N_20899);
xor U21298 (N_21298,N_20006,N_20976);
and U21299 (N_21299,N_20522,N_20005);
xnor U21300 (N_21300,N_20800,N_20051);
nand U21301 (N_21301,N_20401,N_20895);
nor U21302 (N_21302,N_20977,N_20836);
or U21303 (N_21303,N_20408,N_20089);
xor U21304 (N_21304,N_20769,N_20825);
and U21305 (N_21305,N_20232,N_20217);
or U21306 (N_21306,N_20156,N_20475);
nor U21307 (N_21307,N_20890,N_20889);
nand U21308 (N_21308,N_20275,N_20630);
xnor U21309 (N_21309,N_20660,N_20266);
xor U21310 (N_21310,N_20445,N_20698);
xnor U21311 (N_21311,N_20857,N_20803);
or U21312 (N_21312,N_20293,N_20473);
nand U21313 (N_21313,N_20426,N_20249);
nor U21314 (N_21314,N_20065,N_20692);
and U21315 (N_21315,N_20202,N_20377);
or U21316 (N_21316,N_20024,N_20115);
and U21317 (N_21317,N_20658,N_20120);
or U21318 (N_21318,N_20564,N_20397);
nand U21319 (N_21319,N_20613,N_20595);
nor U21320 (N_21320,N_20928,N_20610);
nor U21321 (N_21321,N_20075,N_20811);
xor U21322 (N_21322,N_20462,N_20031);
and U21323 (N_21323,N_20615,N_20392);
and U21324 (N_21324,N_20320,N_20373);
or U21325 (N_21325,N_20997,N_20943);
nand U21326 (N_21326,N_20507,N_20913);
nand U21327 (N_21327,N_20735,N_20297);
xor U21328 (N_21328,N_20181,N_20640);
or U21329 (N_21329,N_20485,N_20948);
nand U21330 (N_21330,N_20446,N_20883);
nand U21331 (N_21331,N_20026,N_20235);
nand U21332 (N_21332,N_20404,N_20158);
or U21333 (N_21333,N_20808,N_20331);
or U21334 (N_21334,N_20891,N_20354);
and U21335 (N_21335,N_20969,N_20662);
and U21336 (N_21336,N_20821,N_20841);
nor U21337 (N_21337,N_20901,N_20596);
or U21338 (N_21338,N_20381,N_20849);
or U21339 (N_21339,N_20741,N_20063);
nand U21340 (N_21340,N_20572,N_20632);
and U21341 (N_21341,N_20590,N_20947);
xnor U21342 (N_21342,N_20192,N_20718);
or U21343 (N_21343,N_20945,N_20691);
and U21344 (N_21344,N_20783,N_20512);
and U21345 (N_21345,N_20716,N_20683);
nand U21346 (N_21346,N_20186,N_20471);
or U21347 (N_21347,N_20511,N_20941);
nor U21348 (N_21348,N_20798,N_20449);
nor U21349 (N_21349,N_20316,N_20957);
or U21350 (N_21350,N_20907,N_20310);
and U21351 (N_21351,N_20717,N_20004);
and U21352 (N_21352,N_20470,N_20328);
nand U21353 (N_21353,N_20099,N_20778);
and U21354 (N_21354,N_20360,N_20566);
or U21355 (N_21355,N_20209,N_20378);
nand U21356 (N_21356,N_20537,N_20745);
or U21357 (N_21357,N_20279,N_20018);
nand U21358 (N_21358,N_20539,N_20415);
nor U21359 (N_21359,N_20056,N_20323);
xnor U21360 (N_21360,N_20905,N_20317);
and U21361 (N_21361,N_20376,N_20017);
and U21362 (N_21362,N_20290,N_20178);
nor U21363 (N_21363,N_20021,N_20349);
and U21364 (N_21364,N_20216,N_20001);
xnor U21365 (N_21365,N_20461,N_20534);
xor U21366 (N_21366,N_20434,N_20014);
or U21367 (N_21367,N_20222,N_20161);
and U21368 (N_21368,N_20733,N_20679);
and U21369 (N_21369,N_20574,N_20707);
xor U21370 (N_21370,N_20520,N_20644);
nand U21371 (N_21371,N_20651,N_20809);
xor U21372 (N_21372,N_20324,N_20524);
xor U21373 (N_21373,N_20936,N_20225);
or U21374 (N_21374,N_20492,N_20556);
xnor U21375 (N_21375,N_20752,N_20766);
nand U21376 (N_21376,N_20455,N_20605);
or U21377 (N_21377,N_20476,N_20487);
or U21378 (N_21378,N_20920,N_20226);
or U21379 (N_21379,N_20321,N_20585);
or U21380 (N_21380,N_20362,N_20405);
or U21381 (N_21381,N_20300,N_20690);
nand U21382 (N_21382,N_20911,N_20604);
xor U21383 (N_21383,N_20621,N_20220);
nor U21384 (N_21384,N_20967,N_20059);
and U21385 (N_21385,N_20438,N_20924);
and U21386 (N_21386,N_20576,N_20584);
nor U21387 (N_21387,N_20575,N_20010);
nor U21388 (N_21388,N_20996,N_20429);
or U21389 (N_21389,N_20078,N_20448);
and U21390 (N_21390,N_20157,N_20268);
nand U21391 (N_21391,N_20776,N_20858);
xor U21392 (N_21392,N_20755,N_20754);
xnor U21393 (N_21393,N_20159,N_20673);
nand U21394 (N_21394,N_20900,N_20086);
nor U21395 (N_21395,N_20419,N_20551);
nor U21396 (N_21396,N_20185,N_20034);
nand U21397 (N_21397,N_20339,N_20732);
nor U21398 (N_21398,N_20558,N_20484);
nor U21399 (N_21399,N_20454,N_20199);
or U21400 (N_21400,N_20387,N_20077);
nor U21401 (N_21401,N_20812,N_20234);
nand U21402 (N_21402,N_20260,N_20491);
or U21403 (N_21403,N_20385,N_20985);
nand U21404 (N_21404,N_20950,N_20058);
nand U21405 (N_21405,N_20863,N_20038);
nor U21406 (N_21406,N_20135,N_20000);
nor U21407 (N_21407,N_20614,N_20241);
or U21408 (N_21408,N_20423,N_20702);
nand U21409 (N_21409,N_20493,N_20337);
or U21410 (N_21410,N_20468,N_20055);
and U21411 (N_21411,N_20530,N_20859);
xor U21412 (N_21412,N_20542,N_20939);
nand U21413 (N_21413,N_20095,N_20087);
or U21414 (N_21414,N_20069,N_20693);
nor U21415 (N_21415,N_20915,N_20659);
xnor U21416 (N_21416,N_20761,N_20946);
and U21417 (N_21417,N_20627,N_20790);
nand U21418 (N_21418,N_20665,N_20771);
xnor U21419 (N_21419,N_20465,N_20623);
and U21420 (N_21420,N_20282,N_20922);
nor U21421 (N_21421,N_20184,N_20909);
nor U21422 (N_21422,N_20792,N_20714);
nor U21423 (N_21423,N_20519,N_20827);
nor U21424 (N_21424,N_20612,N_20760);
and U21425 (N_21425,N_20565,N_20451);
xor U21426 (N_21426,N_20949,N_20869);
xor U21427 (N_21427,N_20577,N_20400);
xor U21428 (N_21428,N_20193,N_20762);
and U21429 (N_21429,N_20816,N_20835);
or U21430 (N_21430,N_20906,N_20685);
nor U21431 (N_21431,N_20113,N_20048);
nor U21432 (N_21432,N_20173,N_20019);
and U21433 (N_21433,N_20620,N_20103);
and U21434 (N_21434,N_20514,N_20921);
nand U21435 (N_21435,N_20884,N_20593);
nand U21436 (N_21436,N_20767,N_20409);
or U21437 (N_21437,N_20164,N_20831);
nand U21438 (N_21438,N_20826,N_20166);
and U21439 (N_21439,N_20700,N_20301);
nor U21440 (N_21440,N_20336,N_20865);
nor U21441 (N_21441,N_20079,N_20844);
nor U21442 (N_21442,N_20380,N_20786);
or U21443 (N_21443,N_20781,N_20960);
and U21444 (N_21444,N_20877,N_20713);
nor U21445 (N_21445,N_20773,N_20703);
or U21446 (N_21446,N_20289,N_20122);
nor U21447 (N_21447,N_20054,N_20541);
and U21448 (N_21448,N_20417,N_20278);
or U21449 (N_21449,N_20503,N_20837);
xor U21450 (N_21450,N_20813,N_20215);
and U21451 (N_21451,N_20041,N_20346);
and U21452 (N_21452,N_20739,N_20190);
nor U21453 (N_21453,N_20121,N_20104);
and U21454 (N_21454,N_20490,N_20035);
nand U21455 (N_21455,N_20153,N_20207);
nand U21456 (N_21456,N_20873,N_20042);
nor U21457 (N_21457,N_20141,N_20256);
nor U21458 (N_21458,N_20699,N_20540);
and U21459 (N_21459,N_20729,N_20073);
xor U21460 (N_21460,N_20932,N_20136);
and U21461 (N_21461,N_20510,N_20389);
or U21462 (N_21462,N_20045,N_20663);
or U21463 (N_21463,N_20709,N_20396);
or U21464 (N_21464,N_20233,N_20708);
xor U21465 (N_21465,N_20820,N_20285);
and U21466 (N_21466,N_20343,N_20412);
or U21467 (N_21467,N_20011,N_20358);
or U21468 (N_21468,N_20518,N_20696);
and U21469 (N_21469,N_20149,N_20131);
and U21470 (N_21470,N_20039,N_20383);
nor U21471 (N_21471,N_20306,N_20689);
and U21472 (N_21472,N_20206,N_20736);
nor U21473 (N_21473,N_20246,N_20601);
and U21474 (N_21474,N_20281,N_20459);
or U21475 (N_21475,N_20971,N_20867);
xnor U21476 (N_21476,N_20616,N_20668);
and U21477 (N_21477,N_20195,N_20012);
nor U21478 (N_21478,N_20112,N_20814);
or U21479 (N_21479,N_20532,N_20407);
xor U21480 (N_21480,N_20402,N_20311);
nand U21481 (N_21481,N_20176,N_20573);
and U21482 (N_21482,N_20746,N_20597);
nor U21483 (N_21483,N_20364,N_20671);
xnor U21484 (N_21484,N_20878,N_20332);
xor U21485 (N_21485,N_20093,N_20040);
and U21486 (N_21486,N_20516,N_20731);
xor U21487 (N_21487,N_20388,N_20611);
xor U21488 (N_21488,N_20020,N_20283);
xor U21489 (N_21489,N_20646,N_20168);
nand U21490 (N_21490,N_20237,N_20105);
nor U21491 (N_21491,N_20775,N_20981);
and U21492 (N_21492,N_20526,N_20231);
or U21493 (N_21493,N_20727,N_20137);
or U21494 (N_21494,N_20357,N_20347);
and U21495 (N_21495,N_20406,N_20846);
and U21496 (N_21496,N_20384,N_20165);
nor U21497 (N_21497,N_20885,N_20314);
or U21498 (N_21498,N_20430,N_20334);
and U21499 (N_21499,N_20267,N_20902);
nor U21500 (N_21500,N_20897,N_20495);
and U21501 (N_21501,N_20850,N_20132);
nor U21502 (N_21502,N_20234,N_20380);
and U21503 (N_21503,N_20601,N_20564);
xnor U21504 (N_21504,N_20739,N_20935);
or U21505 (N_21505,N_20798,N_20486);
xor U21506 (N_21506,N_20980,N_20714);
nor U21507 (N_21507,N_20118,N_20518);
xnor U21508 (N_21508,N_20446,N_20936);
nand U21509 (N_21509,N_20546,N_20010);
and U21510 (N_21510,N_20084,N_20662);
xor U21511 (N_21511,N_20216,N_20899);
nand U21512 (N_21512,N_20705,N_20346);
nand U21513 (N_21513,N_20047,N_20756);
xor U21514 (N_21514,N_20770,N_20383);
or U21515 (N_21515,N_20556,N_20970);
or U21516 (N_21516,N_20106,N_20316);
xor U21517 (N_21517,N_20854,N_20234);
or U21518 (N_21518,N_20907,N_20008);
xnor U21519 (N_21519,N_20062,N_20565);
nand U21520 (N_21520,N_20059,N_20891);
nand U21521 (N_21521,N_20050,N_20395);
nand U21522 (N_21522,N_20313,N_20979);
and U21523 (N_21523,N_20276,N_20883);
xor U21524 (N_21524,N_20860,N_20047);
and U21525 (N_21525,N_20008,N_20150);
or U21526 (N_21526,N_20888,N_20765);
nor U21527 (N_21527,N_20133,N_20462);
xor U21528 (N_21528,N_20443,N_20774);
and U21529 (N_21529,N_20352,N_20546);
and U21530 (N_21530,N_20943,N_20178);
or U21531 (N_21531,N_20660,N_20557);
and U21532 (N_21532,N_20669,N_20229);
nand U21533 (N_21533,N_20833,N_20201);
nor U21534 (N_21534,N_20010,N_20767);
or U21535 (N_21535,N_20084,N_20123);
xor U21536 (N_21536,N_20196,N_20694);
xor U21537 (N_21537,N_20094,N_20095);
nor U21538 (N_21538,N_20341,N_20418);
and U21539 (N_21539,N_20538,N_20408);
nand U21540 (N_21540,N_20252,N_20050);
nand U21541 (N_21541,N_20547,N_20829);
or U21542 (N_21542,N_20660,N_20911);
or U21543 (N_21543,N_20660,N_20933);
nand U21544 (N_21544,N_20213,N_20116);
xor U21545 (N_21545,N_20401,N_20665);
and U21546 (N_21546,N_20113,N_20013);
nand U21547 (N_21547,N_20877,N_20962);
nor U21548 (N_21548,N_20305,N_20903);
or U21549 (N_21549,N_20071,N_20474);
nor U21550 (N_21550,N_20656,N_20900);
nor U21551 (N_21551,N_20755,N_20933);
or U21552 (N_21552,N_20244,N_20951);
and U21553 (N_21553,N_20091,N_20538);
nand U21554 (N_21554,N_20289,N_20713);
xor U21555 (N_21555,N_20390,N_20104);
and U21556 (N_21556,N_20506,N_20377);
and U21557 (N_21557,N_20882,N_20793);
nand U21558 (N_21558,N_20538,N_20502);
xnor U21559 (N_21559,N_20435,N_20172);
nor U21560 (N_21560,N_20659,N_20862);
nand U21561 (N_21561,N_20421,N_20586);
or U21562 (N_21562,N_20421,N_20279);
and U21563 (N_21563,N_20124,N_20345);
nor U21564 (N_21564,N_20588,N_20408);
xor U21565 (N_21565,N_20709,N_20028);
nand U21566 (N_21566,N_20000,N_20761);
nor U21567 (N_21567,N_20237,N_20987);
and U21568 (N_21568,N_20394,N_20359);
or U21569 (N_21569,N_20973,N_20722);
xor U21570 (N_21570,N_20050,N_20825);
or U21571 (N_21571,N_20887,N_20526);
and U21572 (N_21572,N_20628,N_20895);
xor U21573 (N_21573,N_20757,N_20061);
nand U21574 (N_21574,N_20610,N_20924);
nand U21575 (N_21575,N_20244,N_20179);
xnor U21576 (N_21576,N_20662,N_20005);
nand U21577 (N_21577,N_20143,N_20516);
nand U21578 (N_21578,N_20853,N_20213);
nor U21579 (N_21579,N_20282,N_20250);
nor U21580 (N_21580,N_20285,N_20338);
and U21581 (N_21581,N_20015,N_20586);
or U21582 (N_21582,N_20714,N_20662);
nand U21583 (N_21583,N_20185,N_20886);
or U21584 (N_21584,N_20328,N_20019);
nor U21585 (N_21585,N_20414,N_20346);
and U21586 (N_21586,N_20458,N_20482);
nor U21587 (N_21587,N_20201,N_20477);
or U21588 (N_21588,N_20567,N_20735);
xnor U21589 (N_21589,N_20805,N_20770);
and U21590 (N_21590,N_20555,N_20358);
xor U21591 (N_21591,N_20132,N_20822);
and U21592 (N_21592,N_20485,N_20880);
or U21593 (N_21593,N_20957,N_20135);
nand U21594 (N_21594,N_20581,N_20923);
nand U21595 (N_21595,N_20080,N_20161);
or U21596 (N_21596,N_20206,N_20780);
or U21597 (N_21597,N_20110,N_20260);
nor U21598 (N_21598,N_20717,N_20034);
or U21599 (N_21599,N_20655,N_20292);
nand U21600 (N_21600,N_20313,N_20267);
or U21601 (N_21601,N_20481,N_20080);
nor U21602 (N_21602,N_20241,N_20820);
or U21603 (N_21603,N_20402,N_20902);
xnor U21604 (N_21604,N_20877,N_20986);
xnor U21605 (N_21605,N_20149,N_20010);
and U21606 (N_21606,N_20486,N_20481);
or U21607 (N_21607,N_20687,N_20093);
or U21608 (N_21608,N_20070,N_20972);
nand U21609 (N_21609,N_20081,N_20994);
and U21610 (N_21610,N_20228,N_20715);
and U21611 (N_21611,N_20437,N_20019);
nor U21612 (N_21612,N_20089,N_20057);
nor U21613 (N_21613,N_20377,N_20010);
nand U21614 (N_21614,N_20458,N_20999);
nor U21615 (N_21615,N_20775,N_20400);
nand U21616 (N_21616,N_20674,N_20019);
nor U21617 (N_21617,N_20955,N_20497);
nor U21618 (N_21618,N_20044,N_20327);
nand U21619 (N_21619,N_20712,N_20583);
nand U21620 (N_21620,N_20862,N_20026);
nor U21621 (N_21621,N_20623,N_20055);
nand U21622 (N_21622,N_20151,N_20501);
nand U21623 (N_21623,N_20893,N_20453);
nand U21624 (N_21624,N_20258,N_20684);
or U21625 (N_21625,N_20130,N_20469);
and U21626 (N_21626,N_20606,N_20745);
nor U21627 (N_21627,N_20141,N_20026);
nor U21628 (N_21628,N_20823,N_20059);
and U21629 (N_21629,N_20877,N_20887);
and U21630 (N_21630,N_20628,N_20386);
or U21631 (N_21631,N_20096,N_20859);
and U21632 (N_21632,N_20534,N_20920);
xnor U21633 (N_21633,N_20813,N_20740);
or U21634 (N_21634,N_20544,N_20969);
or U21635 (N_21635,N_20586,N_20972);
and U21636 (N_21636,N_20455,N_20864);
or U21637 (N_21637,N_20408,N_20173);
xor U21638 (N_21638,N_20466,N_20483);
nor U21639 (N_21639,N_20704,N_20213);
nand U21640 (N_21640,N_20049,N_20421);
or U21641 (N_21641,N_20610,N_20794);
or U21642 (N_21642,N_20650,N_20700);
and U21643 (N_21643,N_20393,N_20496);
or U21644 (N_21644,N_20803,N_20578);
xor U21645 (N_21645,N_20073,N_20632);
or U21646 (N_21646,N_20522,N_20238);
nor U21647 (N_21647,N_20914,N_20029);
or U21648 (N_21648,N_20588,N_20506);
nor U21649 (N_21649,N_20040,N_20031);
and U21650 (N_21650,N_20355,N_20143);
xor U21651 (N_21651,N_20134,N_20452);
xnor U21652 (N_21652,N_20511,N_20575);
nand U21653 (N_21653,N_20344,N_20832);
xor U21654 (N_21654,N_20677,N_20801);
xor U21655 (N_21655,N_20672,N_20083);
or U21656 (N_21656,N_20155,N_20805);
and U21657 (N_21657,N_20949,N_20901);
xor U21658 (N_21658,N_20215,N_20552);
xor U21659 (N_21659,N_20010,N_20185);
or U21660 (N_21660,N_20579,N_20293);
or U21661 (N_21661,N_20164,N_20070);
xnor U21662 (N_21662,N_20588,N_20333);
nand U21663 (N_21663,N_20106,N_20589);
xnor U21664 (N_21664,N_20470,N_20987);
nand U21665 (N_21665,N_20916,N_20375);
and U21666 (N_21666,N_20765,N_20517);
and U21667 (N_21667,N_20527,N_20903);
nand U21668 (N_21668,N_20132,N_20529);
nand U21669 (N_21669,N_20441,N_20976);
nor U21670 (N_21670,N_20792,N_20837);
nor U21671 (N_21671,N_20034,N_20514);
nand U21672 (N_21672,N_20507,N_20447);
nand U21673 (N_21673,N_20801,N_20713);
nor U21674 (N_21674,N_20689,N_20212);
xor U21675 (N_21675,N_20588,N_20021);
nand U21676 (N_21676,N_20217,N_20113);
and U21677 (N_21677,N_20487,N_20438);
nand U21678 (N_21678,N_20224,N_20166);
nor U21679 (N_21679,N_20884,N_20887);
nand U21680 (N_21680,N_20468,N_20880);
nor U21681 (N_21681,N_20852,N_20455);
or U21682 (N_21682,N_20931,N_20792);
nor U21683 (N_21683,N_20728,N_20648);
or U21684 (N_21684,N_20180,N_20896);
xnor U21685 (N_21685,N_20053,N_20345);
and U21686 (N_21686,N_20926,N_20465);
or U21687 (N_21687,N_20874,N_20544);
or U21688 (N_21688,N_20370,N_20063);
nand U21689 (N_21689,N_20901,N_20135);
xor U21690 (N_21690,N_20390,N_20629);
and U21691 (N_21691,N_20456,N_20174);
nand U21692 (N_21692,N_20635,N_20288);
xnor U21693 (N_21693,N_20330,N_20261);
xor U21694 (N_21694,N_20635,N_20445);
xor U21695 (N_21695,N_20606,N_20237);
nor U21696 (N_21696,N_20409,N_20093);
nand U21697 (N_21697,N_20080,N_20331);
or U21698 (N_21698,N_20982,N_20630);
and U21699 (N_21699,N_20342,N_20754);
and U21700 (N_21700,N_20097,N_20017);
xor U21701 (N_21701,N_20478,N_20074);
and U21702 (N_21702,N_20839,N_20100);
nand U21703 (N_21703,N_20342,N_20372);
xor U21704 (N_21704,N_20742,N_20382);
and U21705 (N_21705,N_20537,N_20269);
and U21706 (N_21706,N_20336,N_20080);
nor U21707 (N_21707,N_20737,N_20194);
or U21708 (N_21708,N_20258,N_20221);
or U21709 (N_21709,N_20759,N_20571);
nor U21710 (N_21710,N_20190,N_20728);
nand U21711 (N_21711,N_20518,N_20626);
and U21712 (N_21712,N_20976,N_20793);
nand U21713 (N_21713,N_20112,N_20430);
and U21714 (N_21714,N_20506,N_20472);
nor U21715 (N_21715,N_20351,N_20365);
xor U21716 (N_21716,N_20955,N_20546);
and U21717 (N_21717,N_20531,N_20704);
xnor U21718 (N_21718,N_20050,N_20424);
nand U21719 (N_21719,N_20530,N_20614);
nor U21720 (N_21720,N_20306,N_20020);
and U21721 (N_21721,N_20166,N_20684);
nand U21722 (N_21722,N_20581,N_20203);
or U21723 (N_21723,N_20449,N_20299);
nand U21724 (N_21724,N_20648,N_20577);
and U21725 (N_21725,N_20240,N_20425);
nand U21726 (N_21726,N_20657,N_20457);
xnor U21727 (N_21727,N_20788,N_20799);
and U21728 (N_21728,N_20780,N_20858);
and U21729 (N_21729,N_20851,N_20352);
nand U21730 (N_21730,N_20456,N_20486);
and U21731 (N_21731,N_20659,N_20324);
nand U21732 (N_21732,N_20122,N_20052);
or U21733 (N_21733,N_20049,N_20843);
xor U21734 (N_21734,N_20851,N_20608);
nand U21735 (N_21735,N_20883,N_20155);
or U21736 (N_21736,N_20815,N_20120);
nor U21737 (N_21737,N_20816,N_20754);
xnor U21738 (N_21738,N_20912,N_20663);
nor U21739 (N_21739,N_20456,N_20199);
and U21740 (N_21740,N_20078,N_20157);
nand U21741 (N_21741,N_20841,N_20508);
and U21742 (N_21742,N_20807,N_20299);
nand U21743 (N_21743,N_20761,N_20223);
or U21744 (N_21744,N_20519,N_20890);
nor U21745 (N_21745,N_20654,N_20252);
nand U21746 (N_21746,N_20806,N_20776);
or U21747 (N_21747,N_20973,N_20977);
and U21748 (N_21748,N_20247,N_20740);
and U21749 (N_21749,N_20727,N_20976);
and U21750 (N_21750,N_20456,N_20529);
or U21751 (N_21751,N_20942,N_20374);
and U21752 (N_21752,N_20033,N_20182);
and U21753 (N_21753,N_20547,N_20118);
xor U21754 (N_21754,N_20612,N_20191);
nand U21755 (N_21755,N_20709,N_20877);
nor U21756 (N_21756,N_20310,N_20862);
and U21757 (N_21757,N_20291,N_20603);
nor U21758 (N_21758,N_20502,N_20525);
and U21759 (N_21759,N_20850,N_20996);
or U21760 (N_21760,N_20233,N_20447);
nor U21761 (N_21761,N_20307,N_20841);
nand U21762 (N_21762,N_20770,N_20162);
nor U21763 (N_21763,N_20286,N_20524);
and U21764 (N_21764,N_20083,N_20000);
or U21765 (N_21765,N_20002,N_20551);
nor U21766 (N_21766,N_20332,N_20726);
or U21767 (N_21767,N_20982,N_20852);
and U21768 (N_21768,N_20054,N_20315);
nor U21769 (N_21769,N_20082,N_20134);
or U21770 (N_21770,N_20433,N_20109);
and U21771 (N_21771,N_20833,N_20077);
nor U21772 (N_21772,N_20353,N_20657);
xor U21773 (N_21773,N_20707,N_20112);
nor U21774 (N_21774,N_20769,N_20529);
nor U21775 (N_21775,N_20887,N_20012);
nand U21776 (N_21776,N_20870,N_20643);
nand U21777 (N_21777,N_20902,N_20952);
xnor U21778 (N_21778,N_20138,N_20971);
nand U21779 (N_21779,N_20448,N_20681);
nor U21780 (N_21780,N_20544,N_20230);
xnor U21781 (N_21781,N_20715,N_20200);
or U21782 (N_21782,N_20600,N_20360);
nand U21783 (N_21783,N_20308,N_20580);
nand U21784 (N_21784,N_20505,N_20700);
or U21785 (N_21785,N_20023,N_20052);
or U21786 (N_21786,N_20270,N_20809);
nand U21787 (N_21787,N_20545,N_20225);
and U21788 (N_21788,N_20163,N_20676);
or U21789 (N_21789,N_20954,N_20884);
xor U21790 (N_21790,N_20395,N_20133);
xnor U21791 (N_21791,N_20634,N_20257);
xor U21792 (N_21792,N_20638,N_20808);
xor U21793 (N_21793,N_20433,N_20543);
and U21794 (N_21794,N_20466,N_20334);
and U21795 (N_21795,N_20134,N_20841);
nand U21796 (N_21796,N_20558,N_20318);
and U21797 (N_21797,N_20602,N_20586);
nand U21798 (N_21798,N_20921,N_20395);
xor U21799 (N_21799,N_20670,N_20516);
nand U21800 (N_21800,N_20900,N_20416);
or U21801 (N_21801,N_20523,N_20899);
or U21802 (N_21802,N_20977,N_20940);
xor U21803 (N_21803,N_20911,N_20126);
nor U21804 (N_21804,N_20971,N_20623);
xor U21805 (N_21805,N_20202,N_20428);
xnor U21806 (N_21806,N_20941,N_20926);
and U21807 (N_21807,N_20661,N_20894);
or U21808 (N_21808,N_20978,N_20781);
or U21809 (N_21809,N_20216,N_20438);
or U21810 (N_21810,N_20128,N_20601);
nor U21811 (N_21811,N_20072,N_20968);
xor U21812 (N_21812,N_20533,N_20000);
nand U21813 (N_21813,N_20925,N_20516);
and U21814 (N_21814,N_20636,N_20445);
xnor U21815 (N_21815,N_20422,N_20936);
xnor U21816 (N_21816,N_20358,N_20463);
xor U21817 (N_21817,N_20348,N_20252);
nor U21818 (N_21818,N_20035,N_20507);
or U21819 (N_21819,N_20259,N_20057);
nand U21820 (N_21820,N_20612,N_20808);
or U21821 (N_21821,N_20266,N_20403);
or U21822 (N_21822,N_20570,N_20424);
nor U21823 (N_21823,N_20611,N_20634);
xor U21824 (N_21824,N_20198,N_20908);
nor U21825 (N_21825,N_20482,N_20616);
nor U21826 (N_21826,N_20708,N_20490);
and U21827 (N_21827,N_20189,N_20469);
nand U21828 (N_21828,N_20962,N_20731);
nor U21829 (N_21829,N_20529,N_20477);
nor U21830 (N_21830,N_20507,N_20472);
nor U21831 (N_21831,N_20036,N_20524);
and U21832 (N_21832,N_20916,N_20942);
nor U21833 (N_21833,N_20790,N_20523);
nand U21834 (N_21834,N_20717,N_20705);
xnor U21835 (N_21835,N_20189,N_20105);
nor U21836 (N_21836,N_20866,N_20777);
or U21837 (N_21837,N_20140,N_20439);
xnor U21838 (N_21838,N_20562,N_20845);
xor U21839 (N_21839,N_20029,N_20700);
and U21840 (N_21840,N_20785,N_20850);
xor U21841 (N_21841,N_20375,N_20246);
nand U21842 (N_21842,N_20244,N_20528);
nor U21843 (N_21843,N_20488,N_20914);
nor U21844 (N_21844,N_20360,N_20293);
and U21845 (N_21845,N_20325,N_20645);
nor U21846 (N_21846,N_20946,N_20594);
or U21847 (N_21847,N_20184,N_20133);
nor U21848 (N_21848,N_20411,N_20453);
nand U21849 (N_21849,N_20089,N_20515);
nand U21850 (N_21850,N_20843,N_20202);
xor U21851 (N_21851,N_20049,N_20138);
xnor U21852 (N_21852,N_20206,N_20396);
xor U21853 (N_21853,N_20957,N_20715);
nor U21854 (N_21854,N_20942,N_20674);
xnor U21855 (N_21855,N_20254,N_20772);
or U21856 (N_21856,N_20424,N_20684);
xor U21857 (N_21857,N_20711,N_20471);
nor U21858 (N_21858,N_20458,N_20235);
xnor U21859 (N_21859,N_20962,N_20716);
nor U21860 (N_21860,N_20215,N_20517);
xnor U21861 (N_21861,N_20845,N_20611);
nand U21862 (N_21862,N_20292,N_20092);
or U21863 (N_21863,N_20463,N_20667);
xnor U21864 (N_21864,N_20286,N_20288);
xor U21865 (N_21865,N_20864,N_20000);
or U21866 (N_21866,N_20855,N_20294);
and U21867 (N_21867,N_20744,N_20406);
nand U21868 (N_21868,N_20617,N_20616);
xnor U21869 (N_21869,N_20951,N_20232);
nor U21870 (N_21870,N_20408,N_20910);
xnor U21871 (N_21871,N_20444,N_20295);
nor U21872 (N_21872,N_20072,N_20937);
xnor U21873 (N_21873,N_20353,N_20057);
and U21874 (N_21874,N_20535,N_20657);
and U21875 (N_21875,N_20028,N_20002);
nand U21876 (N_21876,N_20423,N_20428);
nand U21877 (N_21877,N_20201,N_20249);
nand U21878 (N_21878,N_20089,N_20782);
and U21879 (N_21879,N_20754,N_20153);
nand U21880 (N_21880,N_20341,N_20737);
nor U21881 (N_21881,N_20435,N_20795);
nor U21882 (N_21882,N_20820,N_20977);
or U21883 (N_21883,N_20907,N_20615);
and U21884 (N_21884,N_20534,N_20342);
nor U21885 (N_21885,N_20769,N_20554);
nor U21886 (N_21886,N_20267,N_20438);
and U21887 (N_21887,N_20859,N_20863);
xor U21888 (N_21888,N_20170,N_20998);
nor U21889 (N_21889,N_20337,N_20314);
nand U21890 (N_21890,N_20216,N_20054);
nor U21891 (N_21891,N_20103,N_20789);
xor U21892 (N_21892,N_20237,N_20527);
xnor U21893 (N_21893,N_20025,N_20831);
nor U21894 (N_21894,N_20167,N_20847);
xor U21895 (N_21895,N_20111,N_20886);
or U21896 (N_21896,N_20155,N_20041);
nor U21897 (N_21897,N_20288,N_20700);
nor U21898 (N_21898,N_20144,N_20282);
or U21899 (N_21899,N_20317,N_20121);
and U21900 (N_21900,N_20816,N_20246);
or U21901 (N_21901,N_20704,N_20600);
and U21902 (N_21902,N_20338,N_20077);
or U21903 (N_21903,N_20062,N_20856);
nand U21904 (N_21904,N_20541,N_20342);
or U21905 (N_21905,N_20882,N_20695);
nor U21906 (N_21906,N_20588,N_20001);
or U21907 (N_21907,N_20322,N_20588);
nand U21908 (N_21908,N_20485,N_20723);
nand U21909 (N_21909,N_20380,N_20919);
or U21910 (N_21910,N_20860,N_20256);
or U21911 (N_21911,N_20695,N_20132);
nand U21912 (N_21912,N_20087,N_20023);
nand U21913 (N_21913,N_20167,N_20746);
and U21914 (N_21914,N_20090,N_20186);
or U21915 (N_21915,N_20138,N_20871);
xor U21916 (N_21916,N_20430,N_20833);
nand U21917 (N_21917,N_20513,N_20807);
and U21918 (N_21918,N_20139,N_20193);
xor U21919 (N_21919,N_20427,N_20179);
xnor U21920 (N_21920,N_20673,N_20761);
or U21921 (N_21921,N_20977,N_20193);
or U21922 (N_21922,N_20011,N_20881);
nand U21923 (N_21923,N_20324,N_20664);
xor U21924 (N_21924,N_20413,N_20830);
nor U21925 (N_21925,N_20593,N_20296);
and U21926 (N_21926,N_20517,N_20749);
nand U21927 (N_21927,N_20956,N_20434);
nor U21928 (N_21928,N_20718,N_20544);
nor U21929 (N_21929,N_20412,N_20730);
nand U21930 (N_21930,N_20976,N_20292);
xnor U21931 (N_21931,N_20683,N_20143);
nor U21932 (N_21932,N_20078,N_20854);
nand U21933 (N_21933,N_20607,N_20509);
xor U21934 (N_21934,N_20050,N_20852);
and U21935 (N_21935,N_20047,N_20463);
or U21936 (N_21936,N_20039,N_20479);
and U21937 (N_21937,N_20307,N_20889);
and U21938 (N_21938,N_20438,N_20253);
and U21939 (N_21939,N_20415,N_20253);
and U21940 (N_21940,N_20605,N_20931);
nor U21941 (N_21941,N_20394,N_20393);
and U21942 (N_21942,N_20794,N_20263);
nand U21943 (N_21943,N_20755,N_20141);
nor U21944 (N_21944,N_20924,N_20175);
xor U21945 (N_21945,N_20481,N_20536);
nand U21946 (N_21946,N_20532,N_20438);
nand U21947 (N_21947,N_20217,N_20026);
nor U21948 (N_21948,N_20046,N_20249);
and U21949 (N_21949,N_20496,N_20910);
nand U21950 (N_21950,N_20644,N_20107);
nand U21951 (N_21951,N_20257,N_20395);
xor U21952 (N_21952,N_20610,N_20857);
xor U21953 (N_21953,N_20907,N_20217);
nand U21954 (N_21954,N_20826,N_20607);
nand U21955 (N_21955,N_20616,N_20449);
nand U21956 (N_21956,N_20447,N_20071);
nor U21957 (N_21957,N_20348,N_20076);
or U21958 (N_21958,N_20337,N_20467);
and U21959 (N_21959,N_20264,N_20064);
and U21960 (N_21960,N_20178,N_20993);
nand U21961 (N_21961,N_20861,N_20413);
nor U21962 (N_21962,N_20278,N_20693);
or U21963 (N_21963,N_20612,N_20618);
nor U21964 (N_21964,N_20960,N_20396);
or U21965 (N_21965,N_20834,N_20179);
or U21966 (N_21966,N_20662,N_20508);
and U21967 (N_21967,N_20010,N_20593);
and U21968 (N_21968,N_20708,N_20032);
and U21969 (N_21969,N_20051,N_20844);
and U21970 (N_21970,N_20506,N_20871);
nand U21971 (N_21971,N_20006,N_20749);
or U21972 (N_21972,N_20441,N_20664);
nor U21973 (N_21973,N_20055,N_20783);
or U21974 (N_21974,N_20232,N_20205);
xor U21975 (N_21975,N_20160,N_20220);
nor U21976 (N_21976,N_20018,N_20605);
xor U21977 (N_21977,N_20578,N_20478);
nand U21978 (N_21978,N_20831,N_20883);
and U21979 (N_21979,N_20484,N_20337);
nor U21980 (N_21980,N_20494,N_20813);
or U21981 (N_21981,N_20465,N_20657);
nand U21982 (N_21982,N_20228,N_20699);
or U21983 (N_21983,N_20363,N_20203);
nand U21984 (N_21984,N_20048,N_20122);
nor U21985 (N_21985,N_20366,N_20277);
nand U21986 (N_21986,N_20723,N_20053);
nor U21987 (N_21987,N_20207,N_20053);
xor U21988 (N_21988,N_20524,N_20149);
and U21989 (N_21989,N_20216,N_20524);
and U21990 (N_21990,N_20559,N_20068);
xnor U21991 (N_21991,N_20754,N_20395);
nor U21992 (N_21992,N_20871,N_20246);
or U21993 (N_21993,N_20607,N_20577);
or U21994 (N_21994,N_20063,N_20747);
or U21995 (N_21995,N_20739,N_20731);
nor U21996 (N_21996,N_20140,N_20820);
nand U21997 (N_21997,N_20003,N_20551);
and U21998 (N_21998,N_20813,N_20219);
and U21999 (N_21999,N_20021,N_20373);
xnor U22000 (N_22000,N_21908,N_21921);
and U22001 (N_22001,N_21078,N_21521);
and U22002 (N_22002,N_21211,N_21034);
nand U22003 (N_22003,N_21097,N_21631);
nand U22004 (N_22004,N_21165,N_21744);
and U22005 (N_22005,N_21766,N_21138);
or U22006 (N_22006,N_21153,N_21300);
xnor U22007 (N_22007,N_21751,N_21713);
and U22008 (N_22008,N_21230,N_21120);
nor U22009 (N_22009,N_21103,N_21293);
xor U22010 (N_22010,N_21564,N_21819);
and U22011 (N_22011,N_21607,N_21099);
nor U22012 (N_22012,N_21167,N_21304);
and U22013 (N_22013,N_21722,N_21694);
xnor U22014 (N_22014,N_21926,N_21410);
nor U22015 (N_22015,N_21669,N_21439);
xor U22016 (N_22016,N_21937,N_21644);
xor U22017 (N_22017,N_21731,N_21295);
nor U22018 (N_22018,N_21770,N_21507);
and U22019 (N_22019,N_21922,N_21584);
xor U22020 (N_22020,N_21656,N_21436);
xnor U22021 (N_22021,N_21031,N_21058);
xnor U22022 (N_22022,N_21091,N_21540);
and U22023 (N_22023,N_21784,N_21449);
and U22024 (N_22024,N_21259,N_21973);
xor U22025 (N_22025,N_21458,N_21805);
xnor U22026 (N_22026,N_21646,N_21387);
nor U22027 (N_22027,N_21615,N_21579);
xnor U22028 (N_22028,N_21358,N_21945);
or U22029 (N_22029,N_21068,N_21581);
nand U22030 (N_22030,N_21965,N_21528);
nand U22031 (N_22031,N_21026,N_21501);
nand U22032 (N_22032,N_21613,N_21611);
and U22033 (N_22033,N_21009,N_21585);
nand U22034 (N_22034,N_21201,N_21318);
nor U22035 (N_22035,N_21172,N_21002);
nand U22036 (N_22036,N_21089,N_21244);
nand U22037 (N_22037,N_21620,N_21196);
and U22038 (N_22038,N_21070,N_21075);
and U22039 (N_22039,N_21468,N_21351);
nor U22040 (N_22040,N_21241,N_21000);
nand U22041 (N_22041,N_21375,N_21434);
and U22042 (N_22042,N_21727,N_21326);
or U22043 (N_22043,N_21189,N_21148);
or U22044 (N_22044,N_21866,N_21511);
or U22045 (N_22045,N_21319,N_21264);
and U22046 (N_22046,N_21905,N_21638);
or U22047 (N_22047,N_21182,N_21232);
and U22048 (N_22048,N_21724,N_21983);
nand U22049 (N_22049,N_21812,N_21831);
nand U22050 (N_22050,N_21255,N_21723);
or U22051 (N_22051,N_21537,N_21231);
xor U22052 (N_22052,N_21701,N_21526);
or U22053 (N_22053,N_21160,N_21597);
nor U22054 (N_22054,N_21726,N_21538);
nor U22055 (N_22055,N_21683,N_21257);
and U22056 (N_22056,N_21207,N_21296);
xnor U22057 (N_22057,N_21833,N_21475);
xor U22058 (N_22058,N_21136,N_21778);
xnor U22059 (N_22059,N_21588,N_21466);
nand U22060 (N_22060,N_21963,N_21117);
and U22061 (N_22061,N_21742,N_21942);
and U22062 (N_22062,N_21903,N_21420);
or U22063 (N_22063,N_21048,N_21333);
or U22064 (N_22064,N_21912,N_21532);
xor U22065 (N_22065,N_21177,N_21971);
and U22066 (N_22066,N_21576,N_21847);
nand U22067 (N_22067,N_21039,N_21567);
xnor U22068 (N_22068,N_21658,N_21663);
and U22069 (N_22069,N_21886,N_21443);
nand U22070 (N_22070,N_21206,N_21561);
or U22071 (N_22071,N_21106,N_21856);
nand U22072 (N_22072,N_21703,N_21592);
nor U22073 (N_22073,N_21515,N_21513);
nand U22074 (N_22074,N_21686,N_21174);
or U22075 (N_22075,N_21964,N_21226);
xor U22076 (N_22076,N_21841,N_21682);
nand U22077 (N_22077,N_21881,N_21634);
nand U22078 (N_22078,N_21479,N_21815);
and U22079 (N_22079,N_21141,N_21888);
nand U22080 (N_22080,N_21630,N_21010);
and U22081 (N_22081,N_21720,N_21889);
nor U22082 (N_22082,N_21876,N_21762);
or U22083 (N_22083,N_21559,N_21090);
nand U22084 (N_22084,N_21645,N_21178);
and U22085 (N_22085,N_21793,N_21494);
and U22086 (N_22086,N_21809,N_21426);
and U22087 (N_22087,N_21523,N_21763);
and U22088 (N_22088,N_21913,N_21556);
xor U22089 (N_22089,N_21531,N_21957);
nand U22090 (N_22090,N_21250,N_21400);
xor U22091 (N_22091,N_21252,N_21814);
nor U22092 (N_22092,N_21782,N_21041);
nand U22093 (N_22093,N_21418,N_21144);
and U22094 (N_22094,N_21168,N_21134);
xnor U22095 (N_22095,N_21381,N_21665);
xnor U22096 (N_22096,N_21279,N_21807);
nor U22097 (N_22097,N_21543,N_21469);
nand U22098 (N_22098,N_21786,N_21935);
or U22099 (N_22099,N_21691,N_21367);
nor U22100 (N_22100,N_21743,N_21525);
nor U22101 (N_22101,N_21083,N_21647);
xnor U22102 (N_22102,N_21895,N_21535);
or U22103 (N_22103,N_21715,N_21643);
or U22104 (N_22104,N_21882,N_21332);
or U22105 (N_22105,N_21376,N_21791);
or U22106 (N_22106,N_21697,N_21917);
nor U22107 (N_22107,N_21877,N_21612);
nor U22108 (N_22108,N_21518,N_21461);
or U22109 (N_22109,N_21008,N_21336);
nand U22110 (N_22110,N_21549,N_21865);
nor U22111 (N_22111,N_21191,N_21920);
and U22112 (N_22112,N_21517,N_21169);
nand U22113 (N_22113,N_21383,N_21896);
or U22114 (N_22114,N_21234,N_21872);
or U22115 (N_22115,N_21648,N_21176);
or U22116 (N_22116,N_21672,N_21498);
xnor U22117 (N_22117,N_21562,N_21893);
nor U22118 (N_22118,N_21308,N_21098);
or U22119 (N_22119,N_21804,N_21578);
and U22120 (N_22120,N_21988,N_21664);
nand U22121 (N_22121,N_21551,N_21080);
nand U22122 (N_22122,N_21282,N_21218);
xnor U22123 (N_22123,N_21455,N_21229);
nor U22124 (N_22124,N_21452,N_21133);
or U22125 (N_22125,N_21087,N_21539);
nor U22126 (N_22126,N_21321,N_21698);
nor U22127 (N_22127,N_21073,N_21056);
nand U22128 (N_22128,N_21021,N_21649);
or U22129 (N_22129,N_21810,N_21057);
xor U22130 (N_22130,N_21030,N_21309);
nand U22131 (N_22131,N_21454,N_21830);
or U22132 (N_22132,N_21844,N_21994);
nor U22133 (N_22133,N_21186,N_21050);
xnor U22134 (N_22134,N_21156,N_21341);
xor U22135 (N_22135,N_21352,N_21173);
and U22136 (N_22136,N_21685,N_21316);
and U22137 (N_22137,N_21977,N_21108);
nor U22138 (N_22138,N_21104,N_21571);
xor U22139 (N_22139,N_21959,N_21604);
or U22140 (N_22140,N_21962,N_21750);
nor U22141 (N_22141,N_21943,N_21142);
xnor U22142 (N_22142,N_21371,N_21480);
nor U22143 (N_22143,N_21553,N_21955);
nand U22144 (N_22144,N_21931,N_21628);
nor U22145 (N_22145,N_21736,N_21402);
nor U22146 (N_22146,N_21981,N_21310);
xor U22147 (N_22147,N_21848,N_21051);
xnor U22148 (N_22148,N_21361,N_21278);
nor U22149 (N_22149,N_21450,N_21359);
or U22150 (N_22150,N_21923,N_21711);
nand U22151 (N_22151,N_21674,N_21222);
or U22152 (N_22152,N_21799,N_21929);
xnor U22153 (N_22153,N_21440,N_21126);
or U22154 (N_22154,N_21933,N_21473);
nand U22155 (N_22155,N_21033,N_21406);
and U22156 (N_22156,N_21353,N_21424);
or U22157 (N_22157,N_21808,N_21155);
and U22158 (N_22158,N_21569,N_21852);
nor U22159 (N_22159,N_21224,N_21357);
nor U22160 (N_22160,N_21772,N_21769);
xnor U22161 (N_22161,N_21476,N_21199);
and U22162 (N_22162,N_21777,N_21552);
xor U22163 (N_22163,N_21688,N_21055);
nand U22164 (N_22164,N_21131,N_21997);
nor U22165 (N_22165,N_21349,N_21835);
or U22166 (N_22166,N_21629,N_21448);
nand U22167 (N_22167,N_21395,N_21392);
and U22168 (N_22168,N_21123,N_21114);
nor U22169 (N_22169,N_21437,N_21188);
and U22170 (N_22170,N_21880,N_21028);
and U22171 (N_22171,N_21758,N_21502);
nor U22172 (N_22172,N_21529,N_21781);
nor U22173 (N_22173,N_21335,N_21006);
nand U22174 (N_22174,N_21785,N_21286);
and U22175 (N_22175,N_21348,N_21737);
xor U22176 (N_22176,N_21487,N_21885);
xnor U22177 (N_22177,N_21347,N_21490);
nor U22178 (N_22178,N_21509,N_21826);
and U22179 (N_22179,N_21415,N_21776);
nand U22180 (N_22180,N_21065,N_21307);
nor U22181 (N_22181,N_21753,N_21143);
nor U22182 (N_22182,N_21012,N_21128);
and U22183 (N_22183,N_21297,N_21795);
or U22184 (N_22184,N_21015,N_21838);
xor U22185 (N_22185,N_21818,N_21305);
and U22186 (N_22186,N_21632,N_21911);
nand U22187 (N_22187,N_21898,N_21356);
nor U22188 (N_22188,N_21122,N_21716);
nor U22189 (N_22189,N_21857,N_21601);
and U22190 (N_22190,N_21100,N_21868);
or U22191 (N_22191,N_21076,N_21240);
nor U22192 (N_22192,N_21702,N_21851);
and U22193 (N_22193,N_21331,N_21024);
and U22194 (N_22194,N_21394,N_21811);
or U22195 (N_22195,N_21657,N_21175);
or U22196 (N_22196,N_21453,N_21695);
nand U22197 (N_22197,N_21652,N_21640);
nor U22198 (N_22198,N_21580,N_21023);
xnor U22199 (N_22199,N_21754,N_21897);
and U22200 (N_22200,N_21533,N_21269);
and U22201 (N_22201,N_21582,N_21520);
nand U22202 (N_22202,N_21684,N_21813);
nor U22203 (N_22203,N_21823,N_21590);
and U22204 (N_22204,N_21329,N_21111);
and U22205 (N_22205,N_21205,N_21314);
or U22206 (N_22206,N_21465,N_21978);
xnor U22207 (N_22207,N_21047,N_21832);
or U22208 (N_22208,N_21270,N_21760);
xnor U22209 (N_22209,N_21970,N_21574);
nand U22210 (N_22210,N_21292,N_21680);
nand U22211 (N_22211,N_21639,N_21478);
or U22212 (N_22212,N_21982,N_21339);
xor U22213 (N_22213,N_21281,N_21239);
xnor U22214 (N_22214,N_21334,N_21779);
nand U22215 (N_22215,N_21547,N_21679);
xnor U22216 (N_22216,N_21867,N_21855);
nand U22217 (N_22217,N_21161,N_21029);
and U22218 (N_22218,N_21514,N_21102);
nand U22219 (N_22219,N_21958,N_21276);
and U22220 (N_22220,N_21527,N_21946);
or U22221 (N_22221,N_21904,N_21414);
nand U22222 (N_22222,N_21049,N_21976);
and U22223 (N_22223,N_21510,N_21005);
nand U22224 (N_22224,N_21875,N_21116);
nor U22225 (N_22225,N_21197,N_21858);
nand U22226 (N_22226,N_21398,N_21642);
nand U22227 (N_22227,N_21947,N_21162);
and U22228 (N_22228,N_21140,N_21074);
nor U22229 (N_22229,N_21360,N_21560);
nand U22230 (N_22230,N_21043,N_21902);
and U22231 (N_22231,N_21052,N_21824);
or U22232 (N_22232,N_21204,N_21302);
and U22233 (N_22233,N_21350,N_21442);
nor U22234 (N_22234,N_21317,N_21625);
or U22235 (N_22235,N_21253,N_21745);
and U22236 (N_22236,N_21312,N_21194);
nand U22237 (N_22237,N_21566,N_21067);
and U22238 (N_22238,N_21616,N_21635);
or U22239 (N_22239,N_21470,N_21079);
and U22240 (N_22240,N_21214,N_21659);
or U22241 (N_22241,N_21198,N_21725);
and U22242 (N_22242,N_21765,N_21405);
or U22243 (N_22243,N_21409,N_21287);
nand U22244 (N_22244,N_21949,N_21825);
xnor U22245 (N_22245,N_21227,N_21545);
nor U22246 (N_22246,N_21863,N_21018);
and U22247 (N_22247,N_21488,N_21671);
and U22248 (N_22248,N_21456,N_21666);
and U22249 (N_22249,N_21121,N_21907);
or U22250 (N_22250,N_21481,N_21673);
nor U22251 (N_22251,N_21365,N_21457);
xnor U22252 (N_22252,N_21071,N_21274);
and U22253 (N_22253,N_21342,N_21396);
nand U22254 (N_22254,N_21602,N_21085);
nor U22255 (N_22255,N_21710,N_21203);
xnor U22256 (N_22256,N_21894,N_21508);
xor U22257 (N_22257,N_21283,N_21215);
and U22258 (N_22258,N_21718,N_21413);
nand U22259 (N_22259,N_21389,N_21570);
or U22260 (N_22260,N_21132,N_21368);
and U22261 (N_22261,N_21555,N_21344);
or U22262 (N_22262,N_21020,N_21064);
and U22263 (N_22263,N_21046,N_21884);
or U22264 (N_22264,N_21924,N_21438);
and U22265 (N_22265,N_21219,N_21447);
nor U22266 (N_22266,N_21054,N_21789);
nor U22267 (N_22267,N_21265,N_21506);
or U22268 (N_22268,N_21407,N_21572);
nor U22269 (N_22269,N_21990,N_21397);
and U22270 (N_22270,N_21843,N_21914);
and U22271 (N_22271,N_21719,N_21157);
and U22272 (N_22272,N_21734,N_21446);
xor U22273 (N_22273,N_21417,N_21113);
or U22274 (N_22274,N_21610,N_21284);
nand U22275 (N_22275,N_21154,N_21032);
nor U22276 (N_22276,N_21275,N_21596);
or U22277 (N_22277,N_21699,N_21130);
or U22278 (N_22278,N_21993,N_21557);
nor U22279 (N_22279,N_21267,N_21906);
and U22280 (N_22280,N_21842,N_21707);
and U22281 (N_22281,N_21337,N_21489);
nand U22282 (N_22282,N_21119,N_21954);
or U22283 (N_22283,N_21803,N_21228);
nand U22284 (N_22284,N_21084,N_21554);
or U22285 (N_22285,N_21996,N_21878);
or U22286 (N_22286,N_21193,N_21313);
nor U22287 (N_22287,N_21441,N_21870);
or U22288 (N_22288,N_21503,N_21916);
and U22289 (N_22289,N_21245,N_21401);
or U22290 (N_22290,N_21693,N_21081);
or U22291 (N_22291,N_21593,N_21624);
or U22292 (N_22292,N_21806,N_21516);
xnor U22293 (N_22293,N_21919,N_21474);
or U22294 (N_22294,N_21505,N_21427);
nor U22295 (N_22295,N_21834,N_21676);
xnor U22296 (N_22296,N_21213,N_21190);
and U22297 (N_22297,N_21027,N_21661);
or U22298 (N_22298,N_21237,N_21690);
and U22299 (N_22299,N_21692,N_21208);
and U22300 (N_22300,N_21626,N_21989);
or U22301 (N_22301,N_21273,N_21416);
or U22302 (N_22302,N_21233,N_21740);
or U22303 (N_22303,N_21938,N_21235);
nor U22304 (N_22304,N_21411,N_21256);
nand U22305 (N_22305,N_21836,N_21845);
nand U22306 (N_22306,N_21217,N_21179);
xor U22307 (N_22307,N_21192,N_21599);
nand U22308 (N_22308,N_21355,N_21678);
nor U22309 (N_22309,N_21864,N_21247);
nor U22310 (N_22310,N_21166,N_21901);
or U22311 (N_22311,N_21974,N_21594);
nand U22312 (N_22312,N_21362,N_21464);
nand U22313 (N_22313,N_21223,N_21550);
and U22314 (N_22314,N_21790,N_21088);
nor U22315 (N_22315,N_21794,N_21595);
nand U22316 (N_22316,N_21650,N_21747);
nand U22317 (N_22317,N_21950,N_21377);
nand U22318 (N_22318,N_21721,N_21925);
nand U22319 (N_22319,N_21484,N_21756);
or U22320 (N_22320,N_21042,N_21568);
and U22321 (N_22321,N_21374,N_21839);
xnor U22322 (N_22322,N_21254,N_21600);
nand U22323 (N_22323,N_21732,N_21757);
or U22324 (N_22324,N_21986,N_21952);
nand U22325 (N_22325,N_21563,N_21059);
or U22326 (N_22326,N_21268,N_21340);
nand U22327 (N_22327,N_21654,N_21522);
and U22328 (N_22328,N_21800,N_21712);
and U22329 (N_22329,N_21496,N_21534);
and U22330 (N_22330,N_21759,N_21618);
nand U22331 (N_22331,N_21202,N_21180);
nor U22332 (N_22332,N_21112,N_21101);
nand U22333 (N_22333,N_21500,N_21783);
xor U22334 (N_22334,N_21565,N_21311);
nor U22335 (N_22335,N_21771,N_21787);
and U22336 (N_22336,N_21798,N_21729);
nor U22337 (N_22337,N_21419,N_21003);
or U22338 (N_22338,N_21934,N_21338);
or U22339 (N_22339,N_21491,N_21236);
nand U22340 (N_22340,N_21939,N_21960);
or U22341 (N_22341,N_21086,N_21967);
nor U22342 (N_22342,N_21752,N_21109);
xor U22343 (N_22343,N_21472,N_21306);
nand U22344 (N_22344,N_21622,N_21975);
nor U22345 (N_22345,N_21343,N_21135);
xnor U22346 (N_22346,N_21951,N_21512);
nand U22347 (N_22347,N_21322,N_21445);
and U22348 (N_22348,N_21382,N_21820);
or U22349 (N_22349,N_21433,N_21956);
nor U22350 (N_22350,N_21151,N_21060);
nand U22351 (N_22351,N_21460,N_21748);
or U22352 (N_22352,N_21431,N_21738);
nand U22353 (N_22353,N_21542,N_21242);
and U22354 (N_22354,N_21899,N_21670);
nor U22355 (N_22355,N_21984,N_21587);
xor U22356 (N_22356,N_21216,N_21277);
xor U22357 (N_22357,N_21181,N_21195);
and U22358 (N_22358,N_21299,N_21854);
nor U22359 (N_22359,N_21164,N_21862);
nor U22360 (N_22360,N_21909,N_21152);
or U22361 (N_22361,N_21828,N_21849);
xor U22362 (N_22362,N_21346,N_21733);
or U22363 (N_22363,N_21384,N_21948);
or U22364 (N_22364,N_21301,N_21764);
xnor U22365 (N_22365,N_21094,N_21797);
and U22366 (N_22366,N_21159,N_21775);
or U22367 (N_22367,N_21115,N_21017);
nor U22368 (N_22368,N_21363,N_21037);
and U22369 (N_22369,N_21541,N_21910);
or U22370 (N_22370,N_21072,N_21873);
and U22371 (N_22371,N_21887,N_21524);
and U22372 (N_22372,N_21290,N_21591);
nor U22373 (N_22373,N_21183,N_21714);
nand U22374 (N_22374,N_21007,N_21036);
or U22375 (N_22375,N_21932,N_21260);
or U22376 (N_22376,N_21822,N_21040);
or U22377 (N_22377,N_21105,N_21477);
xor U22378 (N_22378,N_21651,N_21266);
nand U22379 (N_22379,N_21330,N_21969);
nand U22380 (N_22380,N_21493,N_21598);
and U22381 (N_22381,N_21077,N_21871);
or U22382 (N_22382,N_21621,N_21294);
nor U22383 (N_22383,N_21927,N_21062);
nand U22384 (N_22384,N_21315,N_21749);
nand U22385 (N_22385,N_21767,N_21280);
and U22386 (N_22386,N_21485,N_21589);
or U22387 (N_22387,N_21373,N_21016);
and U22388 (N_22388,N_21422,N_21482);
nor U22389 (N_22389,N_21243,N_21463);
or U22390 (N_22390,N_21019,N_21263);
nand U22391 (N_22391,N_21861,N_21998);
or U22392 (N_22392,N_21660,N_21096);
nor U22393 (N_22393,N_21495,N_21892);
or U22394 (N_22394,N_21044,N_21704);
xnor U22395 (N_22395,N_21385,N_21092);
xor U22396 (N_22396,N_21788,N_21827);
or U22397 (N_22397,N_21430,N_21558);
nand U22398 (N_22398,N_21125,N_21379);
nand U22399 (N_22399,N_21735,N_21623);
and U22400 (N_22400,N_21486,N_21082);
xor U22401 (N_22401,N_21936,N_21380);
or U22402 (N_22402,N_21289,N_21200);
or U22403 (N_22403,N_21700,N_21303);
and U22404 (N_22404,N_21614,N_21435);
nor U22405 (N_22405,N_21246,N_21999);
nor U22406 (N_22406,N_21467,N_21428);
and U22407 (N_22407,N_21390,N_21364);
nor U22408 (N_22408,N_21404,N_21345);
nor U22409 (N_22409,N_21966,N_21953);
nor U22410 (N_22410,N_21608,N_21874);
xor U22411 (N_22411,N_21627,N_21483);
nand U22412 (N_22412,N_21548,N_21220);
nand U22413 (N_22413,N_21066,N_21504);
and U22414 (N_22414,N_21991,N_21829);
xor U22415 (N_22415,N_21285,N_21022);
or U22416 (N_22416,N_21796,N_21158);
nand U22417 (N_22417,N_21163,N_21425);
nor U22418 (N_22418,N_21251,N_21928);
xnor U22419 (N_22419,N_21792,N_21147);
xor U22420 (N_22420,N_21837,N_21900);
or U22421 (N_22421,N_21107,N_21972);
nor U22422 (N_22422,N_21497,N_21378);
or U22423 (N_22423,N_21408,N_21212);
and U22424 (N_22424,N_21961,N_21846);
nand U22425 (N_22425,N_21850,N_21768);
nand U22426 (N_22426,N_21677,N_21746);
nor U22427 (N_22427,N_21451,N_21209);
nand U22428 (N_22428,N_21323,N_21110);
xnor U22429 (N_22429,N_21655,N_21603);
nor U22430 (N_22430,N_21124,N_21586);
nor U22431 (N_22431,N_21980,N_21968);
or U22432 (N_22432,N_21262,N_21883);
xor U22433 (N_22433,N_21930,N_21817);
nand U22434 (N_22434,N_21370,N_21577);
xor U22435 (N_22435,N_21272,N_21429);
nand U22436 (N_22436,N_21421,N_21221);
nand U22437 (N_22437,N_21717,N_21462);
xor U22438 (N_22438,N_21755,N_21860);
nor U22439 (N_22439,N_21609,N_21519);
and U22440 (N_22440,N_21859,N_21891);
and U22441 (N_22441,N_21249,N_21399);
and U22442 (N_22442,N_21146,N_21271);
nor U22443 (N_22443,N_21992,N_21014);
nor U22444 (N_22444,N_21816,N_21004);
nand U22445 (N_22445,N_21139,N_21773);
or U22446 (N_22446,N_21170,N_21011);
and U22447 (N_22447,N_21320,N_21328);
nand U22448 (N_22448,N_21530,N_21979);
nand U22449 (N_22449,N_21915,N_21187);
and U22450 (N_22450,N_21633,N_21354);
xnor U22451 (N_22451,N_21403,N_21471);
or U22452 (N_22452,N_21730,N_21492);
xor U22453 (N_22453,N_21637,N_21689);
and U22454 (N_22454,N_21093,N_21137);
xnor U22455 (N_22455,N_21583,N_21261);
and U22456 (N_22456,N_21127,N_21780);
or U22457 (N_22457,N_21879,N_21298);
and U22458 (N_22458,N_21705,N_21940);
or U22459 (N_22459,N_21063,N_21369);
nor U22460 (N_22460,N_21069,N_21821);
or U22461 (N_22461,N_21184,N_21739);
nor U22462 (N_22462,N_21606,N_21653);
and U22463 (N_22463,N_21225,N_21444);
and U22464 (N_22464,N_21546,N_21995);
nor U22465 (N_22465,N_21459,N_21741);
or U22466 (N_22466,N_21210,N_21118);
nand U22467 (N_22467,N_21709,N_21918);
or U22468 (N_22468,N_21696,N_21366);
nand U22469 (N_22469,N_21761,N_21944);
nor U22470 (N_22470,N_21985,N_21619);
xor U22471 (N_22471,N_21038,N_21432);
xnor U22472 (N_22472,N_21890,N_21372);
nor U22473 (N_22473,N_21045,N_21061);
nor U22474 (N_22474,N_21393,N_21288);
xnor U22475 (N_22475,N_21801,N_21013);
nor U22476 (N_22476,N_21291,N_21573);
nor U22477 (N_22477,N_21544,N_21145);
and U22478 (N_22478,N_21238,N_21941);
nand U22479 (N_22479,N_21687,N_21681);
and U22480 (N_22480,N_21706,N_21386);
and U22481 (N_22481,N_21171,N_21575);
and U22482 (N_22482,N_21150,N_21391);
nand U22483 (N_22483,N_21605,N_21325);
and U22484 (N_22484,N_21840,N_21675);
nand U22485 (N_22485,N_21708,N_21774);
or U22486 (N_22486,N_21667,N_21869);
xnor U22487 (N_22487,N_21035,N_21258);
nor U22488 (N_22488,N_21668,N_21248);
or U22489 (N_22489,N_21499,N_21025);
or U22490 (N_22490,N_21853,N_21327);
and U22491 (N_22491,N_21129,N_21001);
nor U22492 (N_22492,N_21388,N_21095);
and U22493 (N_22493,N_21987,N_21423);
or U22494 (N_22494,N_21185,N_21324);
and U22495 (N_22495,N_21617,N_21802);
xnor U22496 (N_22496,N_21536,N_21636);
and U22497 (N_22497,N_21053,N_21641);
nand U22498 (N_22498,N_21412,N_21662);
and U22499 (N_22499,N_21149,N_21728);
and U22500 (N_22500,N_21001,N_21246);
nand U22501 (N_22501,N_21048,N_21491);
nand U22502 (N_22502,N_21770,N_21256);
or U22503 (N_22503,N_21100,N_21140);
xor U22504 (N_22504,N_21246,N_21071);
nand U22505 (N_22505,N_21535,N_21143);
or U22506 (N_22506,N_21658,N_21501);
or U22507 (N_22507,N_21106,N_21019);
or U22508 (N_22508,N_21010,N_21889);
nor U22509 (N_22509,N_21701,N_21566);
xor U22510 (N_22510,N_21524,N_21265);
xnor U22511 (N_22511,N_21003,N_21994);
nor U22512 (N_22512,N_21290,N_21358);
or U22513 (N_22513,N_21716,N_21617);
nor U22514 (N_22514,N_21762,N_21228);
and U22515 (N_22515,N_21247,N_21399);
or U22516 (N_22516,N_21838,N_21635);
or U22517 (N_22517,N_21845,N_21576);
nor U22518 (N_22518,N_21645,N_21037);
and U22519 (N_22519,N_21620,N_21377);
nand U22520 (N_22520,N_21263,N_21347);
nor U22521 (N_22521,N_21177,N_21556);
and U22522 (N_22522,N_21596,N_21563);
xnor U22523 (N_22523,N_21185,N_21067);
xor U22524 (N_22524,N_21751,N_21645);
xnor U22525 (N_22525,N_21122,N_21801);
nor U22526 (N_22526,N_21626,N_21722);
nor U22527 (N_22527,N_21411,N_21068);
and U22528 (N_22528,N_21505,N_21035);
nor U22529 (N_22529,N_21604,N_21563);
or U22530 (N_22530,N_21203,N_21612);
xor U22531 (N_22531,N_21331,N_21650);
nor U22532 (N_22532,N_21786,N_21447);
xnor U22533 (N_22533,N_21006,N_21597);
nor U22534 (N_22534,N_21887,N_21427);
nor U22535 (N_22535,N_21326,N_21534);
or U22536 (N_22536,N_21800,N_21043);
and U22537 (N_22537,N_21280,N_21030);
or U22538 (N_22538,N_21900,N_21206);
or U22539 (N_22539,N_21612,N_21417);
nand U22540 (N_22540,N_21102,N_21982);
nand U22541 (N_22541,N_21140,N_21646);
xor U22542 (N_22542,N_21008,N_21035);
or U22543 (N_22543,N_21771,N_21274);
or U22544 (N_22544,N_21316,N_21143);
nand U22545 (N_22545,N_21894,N_21845);
and U22546 (N_22546,N_21603,N_21808);
or U22547 (N_22547,N_21220,N_21182);
and U22548 (N_22548,N_21423,N_21997);
or U22549 (N_22549,N_21596,N_21081);
and U22550 (N_22550,N_21149,N_21716);
xnor U22551 (N_22551,N_21428,N_21388);
or U22552 (N_22552,N_21276,N_21176);
nand U22553 (N_22553,N_21228,N_21650);
nor U22554 (N_22554,N_21092,N_21695);
nor U22555 (N_22555,N_21698,N_21707);
or U22556 (N_22556,N_21764,N_21569);
nor U22557 (N_22557,N_21893,N_21956);
nand U22558 (N_22558,N_21500,N_21107);
nand U22559 (N_22559,N_21362,N_21577);
nor U22560 (N_22560,N_21969,N_21520);
xor U22561 (N_22561,N_21289,N_21853);
or U22562 (N_22562,N_21056,N_21447);
nand U22563 (N_22563,N_21431,N_21727);
or U22564 (N_22564,N_21399,N_21463);
and U22565 (N_22565,N_21695,N_21145);
nor U22566 (N_22566,N_21066,N_21041);
or U22567 (N_22567,N_21540,N_21649);
and U22568 (N_22568,N_21118,N_21281);
or U22569 (N_22569,N_21934,N_21175);
xnor U22570 (N_22570,N_21947,N_21743);
nand U22571 (N_22571,N_21484,N_21374);
nor U22572 (N_22572,N_21560,N_21302);
xor U22573 (N_22573,N_21555,N_21629);
nand U22574 (N_22574,N_21243,N_21445);
nand U22575 (N_22575,N_21496,N_21432);
or U22576 (N_22576,N_21110,N_21273);
or U22577 (N_22577,N_21901,N_21448);
xnor U22578 (N_22578,N_21526,N_21649);
nor U22579 (N_22579,N_21240,N_21402);
nor U22580 (N_22580,N_21667,N_21223);
xor U22581 (N_22581,N_21298,N_21816);
xnor U22582 (N_22582,N_21962,N_21218);
and U22583 (N_22583,N_21040,N_21646);
and U22584 (N_22584,N_21710,N_21237);
nor U22585 (N_22585,N_21914,N_21602);
or U22586 (N_22586,N_21015,N_21950);
nand U22587 (N_22587,N_21098,N_21337);
or U22588 (N_22588,N_21414,N_21720);
nand U22589 (N_22589,N_21428,N_21524);
and U22590 (N_22590,N_21955,N_21956);
nor U22591 (N_22591,N_21331,N_21820);
nand U22592 (N_22592,N_21380,N_21982);
nor U22593 (N_22593,N_21007,N_21440);
nand U22594 (N_22594,N_21542,N_21344);
nor U22595 (N_22595,N_21489,N_21947);
nor U22596 (N_22596,N_21352,N_21738);
or U22597 (N_22597,N_21601,N_21109);
nand U22598 (N_22598,N_21516,N_21529);
and U22599 (N_22599,N_21849,N_21163);
nor U22600 (N_22600,N_21277,N_21015);
or U22601 (N_22601,N_21458,N_21879);
nor U22602 (N_22602,N_21164,N_21220);
nor U22603 (N_22603,N_21813,N_21093);
nand U22604 (N_22604,N_21448,N_21421);
nor U22605 (N_22605,N_21965,N_21885);
nor U22606 (N_22606,N_21264,N_21763);
nor U22607 (N_22607,N_21408,N_21619);
nand U22608 (N_22608,N_21026,N_21032);
and U22609 (N_22609,N_21169,N_21848);
or U22610 (N_22610,N_21420,N_21700);
and U22611 (N_22611,N_21562,N_21250);
or U22612 (N_22612,N_21334,N_21981);
xor U22613 (N_22613,N_21860,N_21055);
nor U22614 (N_22614,N_21066,N_21242);
or U22615 (N_22615,N_21700,N_21182);
and U22616 (N_22616,N_21088,N_21093);
or U22617 (N_22617,N_21771,N_21081);
and U22618 (N_22618,N_21435,N_21891);
xor U22619 (N_22619,N_21523,N_21280);
nand U22620 (N_22620,N_21257,N_21030);
and U22621 (N_22621,N_21102,N_21672);
xor U22622 (N_22622,N_21321,N_21014);
xor U22623 (N_22623,N_21457,N_21330);
nand U22624 (N_22624,N_21576,N_21757);
xor U22625 (N_22625,N_21674,N_21472);
xnor U22626 (N_22626,N_21582,N_21719);
or U22627 (N_22627,N_21806,N_21967);
xnor U22628 (N_22628,N_21093,N_21250);
xnor U22629 (N_22629,N_21477,N_21889);
or U22630 (N_22630,N_21096,N_21970);
xor U22631 (N_22631,N_21508,N_21831);
nor U22632 (N_22632,N_21224,N_21240);
nand U22633 (N_22633,N_21682,N_21922);
and U22634 (N_22634,N_21341,N_21843);
nand U22635 (N_22635,N_21094,N_21493);
nand U22636 (N_22636,N_21897,N_21483);
xnor U22637 (N_22637,N_21222,N_21635);
or U22638 (N_22638,N_21944,N_21888);
xnor U22639 (N_22639,N_21594,N_21148);
nand U22640 (N_22640,N_21018,N_21313);
nand U22641 (N_22641,N_21630,N_21172);
xor U22642 (N_22642,N_21746,N_21730);
nand U22643 (N_22643,N_21524,N_21630);
nor U22644 (N_22644,N_21316,N_21313);
or U22645 (N_22645,N_21031,N_21605);
or U22646 (N_22646,N_21061,N_21238);
nand U22647 (N_22647,N_21055,N_21656);
or U22648 (N_22648,N_21191,N_21771);
and U22649 (N_22649,N_21605,N_21693);
nand U22650 (N_22650,N_21364,N_21573);
xnor U22651 (N_22651,N_21589,N_21632);
nor U22652 (N_22652,N_21474,N_21983);
nand U22653 (N_22653,N_21464,N_21840);
nand U22654 (N_22654,N_21659,N_21733);
or U22655 (N_22655,N_21259,N_21494);
and U22656 (N_22656,N_21337,N_21532);
or U22657 (N_22657,N_21466,N_21847);
and U22658 (N_22658,N_21298,N_21593);
and U22659 (N_22659,N_21220,N_21363);
nor U22660 (N_22660,N_21210,N_21972);
or U22661 (N_22661,N_21887,N_21145);
nor U22662 (N_22662,N_21042,N_21855);
or U22663 (N_22663,N_21985,N_21258);
xnor U22664 (N_22664,N_21615,N_21790);
nand U22665 (N_22665,N_21011,N_21270);
xnor U22666 (N_22666,N_21417,N_21086);
or U22667 (N_22667,N_21162,N_21895);
xor U22668 (N_22668,N_21343,N_21884);
xor U22669 (N_22669,N_21905,N_21899);
xor U22670 (N_22670,N_21166,N_21609);
and U22671 (N_22671,N_21797,N_21633);
xor U22672 (N_22672,N_21738,N_21199);
nor U22673 (N_22673,N_21563,N_21087);
and U22674 (N_22674,N_21942,N_21109);
nand U22675 (N_22675,N_21901,N_21943);
or U22676 (N_22676,N_21144,N_21103);
xor U22677 (N_22677,N_21232,N_21398);
or U22678 (N_22678,N_21803,N_21393);
nor U22679 (N_22679,N_21866,N_21249);
and U22680 (N_22680,N_21375,N_21450);
and U22681 (N_22681,N_21811,N_21562);
or U22682 (N_22682,N_21353,N_21196);
or U22683 (N_22683,N_21523,N_21773);
and U22684 (N_22684,N_21295,N_21590);
or U22685 (N_22685,N_21708,N_21066);
or U22686 (N_22686,N_21934,N_21686);
xor U22687 (N_22687,N_21503,N_21172);
or U22688 (N_22688,N_21393,N_21796);
nor U22689 (N_22689,N_21143,N_21641);
or U22690 (N_22690,N_21642,N_21052);
nor U22691 (N_22691,N_21455,N_21553);
nor U22692 (N_22692,N_21046,N_21465);
nand U22693 (N_22693,N_21018,N_21380);
nand U22694 (N_22694,N_21980,N_21249);
nand U22695 (N_22695,N_21449,N_21470);
or U22696 (N_22696,N_21895,N_21723);
and U22697 (N_22697,N_21290,N_21070);
xor U22698 (N_22698,N_21642,N_21604);
and U22699 (N_22699,N_21747,N_21873);
nor U22700 (N_22700,N_21236,N_21250);
nor U22701 (N_22701,N_21972,N_21583);
nor U22702 (N_22702,N_21867,N_21529);
nor U22703 (N_22703,N_21542,N_21522);
or U22704 (N_22704,N_21667,N_21445);
and U22705 (N_22705,N_21380,N_21279);
and U22706 (N_22706,N_21784,N_21876);
xnor U22707 (N_22707,N_21626,N_21495);
xor U22708 (N_22708,N_21527,N_21824);
and U22709 (N_22709,N_21659,N_21009);
nand U22710 (N_22710,N_21885,N_21989);
nand U22711 (N_22711,N_21243,N_21456);
and U22712 (N_22712,N_21941,N_21436);
nand U22713 (N_22713,N_21149,N_21271);
nand U22714 (N_22714,N_21901,N_21629);
nand U22715 (N_22715,N_21634,N_21289);
nand U22716 (N_22716,N_21032,N_21257);
and U22717 (N_22717,N_21728,N_21433);
nor U22718 (N_22718,N_21813,N_21585);
nor U22719 (N_22719,N_21150,N_21450);
nand U22720 (N_22720,N_21132,N_21565);
xnor U22721 (N_22721,N_21033,N_21883);
or U22722 (N_22722,N_21103,N_21816);
nor U22723 (N_22723,N_21488,N_21068);
nand U22724 (N_22724,N_21904,N_21893);
nor U22725 (N_22725,N_21698,N_21985);
or U22726 (N_22726,N_21125,N_21713);
or U22727 (N_22727,N_21242,N_21452);
xor U22728 (N_22728,N_21495,N_21788);
nor U22729 (N_22729,N_21418,N_21292);
nand U22730 (N_22730,N_21864,N_21298);
and U22731 (N_22731,N_21587,N_21453);
or U22732 (N_22732,N_21507,N_21401);
xor U22733 (N_22733,N_21775,N_21779);
and U22734 (N_22734,N_21245,N_21617);
nor U22735 (N_22735,N_21799,N_21479);
or U22736 (N_22736,N_21444,N_21719);
nand U22737 (N_22737,N_21795,N_21497);
nor U22738 (N_22738,N_21662,N_21337);
or U22739 (N_22739,N_21882,N_21719);
and U22740 (N_22740,N_21866,N_21779);
nor U22741 (N_22741,N_21399,N_21875);
nor U22742 (N_22742,N_21444,N_21945);
nor U22743 (N_22743,N_21173,N_21667);
nor U22744 (N_22744,N_21132,N_21626);
xnor U22745 (N_22745,N_21799,N_21302);
nor U22746 (N_22746,N_21750,N_21739);
nor U22747 (N_22747,N_21199,N_21898);
and U22748 (N_22748,N_21598,N_21419);
nor U22749 (N_22749,N_21070,N_21393);
nand U22750 (N_22750,N_21438,N_21281);
and U22751 (N_22751,N_21054,N_21486);
and U22752 (N_22752,N_21252,N_21177);
or U22753 (N_22753,N_21829,N_21186);
xor U22754 (N_22754,N_21532,N_21816);
nor U22755 (N_22755,N_21460,N_21179);
and U22756 (N_22756,N_21745,N_21725);
nand U22757 (N_22757,N_21854,N_21290);
or U22758 (N_22758,N_21323,N_21754);
nand U22759 (N_22759,N_21178,N_21931);
nand U22760 (N_22760,N_21279,N_21123);
and U22761 (N_22761,N_21594,N_21991);
nand U22762 (N_22762,N_21571,N_21454);
and U22763 (N_22763,N_21542,N_21173);
and U22764 (N_22764,N_21259,N_21418);
nand U22765 (N_22765,N_21866,N_21440);
nand U22766 (N_22766,N_21887,N_21694);
xor U22767 (N_22767,N_21524,N_21307);
xor U22768 (N_22768,N_21172,N_21304);
and U22769 (N_22769,N_21531,N_21071);
and U22770 (N_22770,N_21088,N_21109);
nand U22771 (N_22771,N_21994,N_21857);
nand U22772 (N_22772,N_21294,N_21507);
and U22773 (N_22773,N_21335,N_21613);
and U22774 (N_22774,N_21749,N_21051);
nand U22775 (N_22775,N_21327,N_21291);
and U22776 (N_22776,N_21015,N_21082);
and U22777 (N_22777,N_21563,N_21639);
or U22778 (N_22778,N_21974,N_21907);
nand U22779 (N_22779,N_21384,N_21780);
and U22780 (N_22780,N_21159,N_21295);
nand U22781 (N_22781,N_21733,N_21078);
xor U22782 (N_22782,N_21967,N_21938);
xnor U22783 (N_22783,N_21501,N_21583);
and U22784 (N_22784,N_21434,N_21008);
and U22785 (N_22785,N_21672,N_21958);
or U22786 (N_22786,N_21463,N_21209);
xnor U22787 (N_22787,N_21023,N_21455);
nor U22788 (N_22788,N_21941,N_21815);
nor U22789 (N_22789,N_21270,N_21881);
nor U22790 (N_22790,N_21397,N_21289);
nand U22791 (N_22791,N_21137,N_21275);
nand U22792 (N_22792,N_21727,N_21163);
nor U22793 (N_22793,N_21263,N_21552);
nand U22794 (N_22794,N_21618,N_21424);
and U22795 (N_22795,N_21706,N_21110);
nand U22796 (N_22796,N_21853,N_21207);
nand U22797 (N_22797,N_21224,N_21968);
xor U22798 (N_22798,N_21501,N_21886);
or U22799 (N_22799,N_21874,N_21213);
or U22800 (N_22800,N_21642,N_21246);
or U22801 (N_22801,N_21825,N_21999);
or U22802 (N_22802,N_21931,N_21915);
xnor U22803 (N_22803,N_21262,N_21861);
or U22804 (N_22804,N_21244,N_21516);
or U22805 (N_22805,N_21223,N_21647);
nand U22806 (N_22806,N_21519,N_21820);
nor U22807 (N_22807,N_21051,N_21170);
or U22808 (N_22808,N_21679,N_21005);
and U22809 (N_22809,N_21540,N_21045);
xnor U22810 (N_22810,N_21217,N_21451);
nor U22811 (N_22811,N_21828,N_21430);
nand U22812 (N_22812,N_21561,N_21699);
xnor U22813 (N_22813,N_21451,N_21136);
nor U22814 (N_22814,N_21083,N_21112);
nor U22815 (N_22815,N_21498,N_21154);
nand U22816 (N_22816,N_21506,N_21868);
xor U22817 (N_22817,N_21051,N_21396);
nand U22818 (N_22818,N_21585,N_21559);
and U22819 (N_22819,N_21873,N_21315);
nor U22820 (N_22820,N_21925,N_21053);
xnor U22821 (N_22821,N_21162,N_21500);
xor U22822 (N_22822,N_21710,N_21090);
nand U22823 (N_22823,N_21257,N_21546);
and U22824 (N_22824,N_21074,N_21327);
nand U22825 (N_22825,N_21989,N_21300);
or U22826 (N_22826,N_21322,N_21300);
and U22827 (N_22827,N_21755,N_21175);
nor U22828 (N_22828,N_21977,N_21197);
or U22829 (N_22829,N_21758,N_21969);
or U22830 (N_22830,N_21629,N_21820);
and U22831 (N_22831,N_21694,N_21321);
nor U22832 (N_22832,N_21176,N_21094);
nand U22833 (N_22833,N_21422,N_21654);
and U22834 (N_22834,N_21187,N_21373);
and U22835 (N_22835,N_21101,N_21025);
nand U22836 (N_22836,N_21477,N_21906);
and U22837 (N_22837,N_21880,N_21670);
nand U22838 (N_22838,N_21257,N_21893);
nor U22839 (N_22839,N_21383,N_21404);
xnor U22840 (N_22840,N_21259,N_21537);
nand U22841 (N_22841,N_21782,N_21189);
xor U22842 (N_22842,N_21775,N_21141);
and U22843 (N_22843,N_21665,N_21964);
xnor U22844 (N_22844,N_21337,N_21504);
or U22845 (N_22845,N_21292,N_21987);
and U22846 (N_22846,N_21874,N_21357);
nand U22847 (N_22847,N_21912,N_21179);
nor U22848 (N_22848,N_21385,N_21676);
nor U22849 (N_22849,N_21005,N_21408);
nor U22850 (N_22850,N_21083,N_21509);
nor U22851 (N_22851,N_21883,N_21759);
or U22852 (N_22852,N_21736,N_21279);
nand U22853 (N_22853,N_21743,N_21584);
nor U22854 (N_22854,N_21477,N_21324);
xor U22855 (N_22855,N_21566,N_21789);
and U22856 (N_22856,N_21550,N_21153);
or U22857 (N_22857,N_21268,N_21402);
xor U22858 (N_22858,N_21468,N_21141);
and U22859 (N_22859,N_21959,N_21283);
or U22860 (N_22860,N_21067,N_21631);
nand U22861 (N_22861,N_21673,N_21824);
nor U22862 (N_22862,N_21354,N_21945);
or U22863 (N_22863,N_21439,N_21180);
nand U22864 (N_22864,N_21803,N_21414);
nand U22865 (N_22865,N_21972,N_21560);
nor U22866 (N_22866,N_21114,N_21074);
nor U22867 (N_22867,N_21564,N_21858);
nand U22868 (N_22868,N_21649,N_21220);
xnor U22869 (N_22869,N_21569,N_21512);
nand U22870 (N_22870,N_21536,N_21589);
nor U22871 (N_22871,N_21591,N_21302);
or U22872 (N_22872,N_21391,N_21889);
and U22873 (N_22873,N_21662,N_21605);
nand U22874 (N_22874,N_21215,N_21819);
xnor U22875 (N_22875,N_21036,N_21625);
nor U22876 (N_22876,N_21173,N_21102);
or U22877 (N_22877,N_21062,N_21648);
nand U22878 (N_22878,N_21510,N_21903);
nor U22879 (N_22879,N_21848,N_21428);
or U22880 (N_22880,N_21519,N_21403);
nor U22881 (N_22881,N_21951,N_21341);
nor U22882 (N_22882,N_21089,N_21975);
nor U22883 (N_22883,N_21988,N_21205);
or U22884 (N_22884,N_21751,N_21347);
nand U22885 (N_22885,N_21993,N_21561);
nor U22886 (N_22886,N_21904,N_21619);
or U22887 (N_22887,N_21405,N_21093);
and U22888 (N_22888,N_21475,N_21668);
and U22889 (N_22889,N_21333,N_21863);
nand U22890 (N_22890,N_21811,N_21425);
nor U22891 (N_22891,N_21325,N_21338);
xor U22892 (N_22892,N_21548,N_21370);
and U22893 (N_22893,N_21186,N_21469);
or U22894 (N_22894,N_21591,N_21228);
and U22895 (N_22895,N_21697,N_21132);
and U22896 (N_22896,N_21863,N_21364);
nor U22897 (N_22897,N_21729,N_21854);
xnor U22898 (N_22898,N_21269,N_21601);
and U22899 (N_22899,N_21380,N_21722);
or U22900 (N_22900,N_21576,N_21325);
or U22901 (N_22901,N_21972,N_21465);
or U22902 (N_22902,N_21577,N_21771);
xnor U22903 (N_22903,N_21131,N_21463);
nor U22904 (N_22904,N_21161,N_21205);
nand U22905 (N_22905,N_21755,N_21773);
nand U22906 (N_22906,N_21754,N_21356);
or U22907 (N_22907,N_21404,N_21053);
nand U22908 (N_22908,N_21674,N_21812);
and U22909 (N_22909,N_21156,N_21119);
and U22910 (N_22910,N_21761,N_21783);
or U22911 (N_22911,N_21909,N_21197);
xnor U22912 (N_22912,N_21975,N_21550);
xnor U22913 (N_22913,N_21536,N_21801);
xor U22914 (N_22914,N_21020,N_21166);
nor U22915 (N_22915,N_21619,N_21616);
or U22916 (N_22916,N_21428,N_21345);
nor U22917 (N_22917,N_21457,N_21200);
xnor U22918 (N_22918,N_21227,N_21261);
xnor U22919 (N_22919,N_21717,N_21342);
or U22920 (N_22920,N_21086,N_21659);
nor U22921 (N_22921,N_21480,N_21169);
and U22922 (N_22922,N_21150,N_21547);
or U22923 (N_22923,N_21808,N_21261);
or U22924 (N_22924,N_21416,N_21620);
or U22925 (N_22925,N_21367,N_21960);
nand U22926 (N_22926,N_21319,N_21178);
nand U22927 (N_22927,N_21124,N_21808);
nand U22928 (N_22928,N_21873,N_21135);
xnor U22929 (N_22929,N_21120,N_21910);
and U22930 (N_22930,N_21012,N_21256);
or U22931 (N_22931,N_21656,N_21955);
or U22932 (N_22932,N_21674,N_21087);
xor U22933 (N_22933,N_21701,N_21391);
nor U22934 (N_22934,N_21085,N_21848);
and U22935 (N_22935,N_21410,N_21209);
or U22936 (N_22936,N_21682,N_21708);
xnor U22937 (N_22937,N_21953,N_21882);
nand U22938 (N_22938,N_21329,N_21281);
nor U22939 (N_22939,N_21689,N_21792);
or U22940 (N_22940,N_21055,N_21947);
xor U22941 (N_22941,N_21745,N_21013);
and U22942 (N_22942,N_21937,N_21184);
and U22943 (N_22943,N_21673,N_21981);
nor U22944 (N_22944,N_21057,N_21583);
and U22945 (N_22945,N_21008,N_21409);
and U22946 (N_22946,N_21050,N_21283);
nand U22947 (N_22947,N_21906,N_21788);
and U22948 (N_22948,N_21546,N_21161);
nor U22949 (N_22949,N_21383,N_21708);
nand U22950 (N_22950,N_21174,N_21911);
xnor U22951 (N_22951,N_21012,N_21572);
nand U22952 (N_22952,N_21343,N_21594);
xnor U22953 (N_22953,N_21656,N_21326);
nor U22954 (N_22954,N_21650,N_21446);
xnor U22955 (N_22955,N_21323,N_21984);
nand U22956 (N_22956,N_21901,N_21087);
xnor U22957 (N_22957,N_21596,N_21191);
xnor U22958 (N_22958,N_21826,N_21175);
nor U22959 (N_22959,N_21447,N_21260);
or U22960 (N_22960,N_21772,N_21845);
nand U22961 (N_22961,N_21708,N_21853);
or U22962 (N_22962,N_21037,N_21936);
nor U22963 (N_22963,N_21220,N_21553);
nor U22964 (N_22964,N_21097,N_21128);
nand U22965 (N_22965,N_21211,N_21888);
nor U22966 (N_22966,N_21994,N_21612);
xnor U22967 (N_22967,N_21594,N_21521);
or U22968 (N_22968,N_21668,N_21742);
or U22969 (N_22969,N_21527,N_21167);
and U22970 (N_22970,N_21825,N_21099);
or U22971 (N_22971,N_21244,N_21366);
nor U22972 (N_22972,N_21132,N_21455);
xor U22973 (N_22973,N_21446,N_21123);
and U22974 (N_22974,N_21783,N_21781);
nand U22975 (N_22975,N_21123,N_21792);
xor U22976 (N_22976,N_21993,N_21847);
xor U22977 (N_22977,N_21380,N_21752);
xnor U22978 (N_22978,N_21810,N_21001);
nor U22979 (N_22979,N_21794,N_21702);
or U22980 (N_22980,N_21439,N_21204);
or U22981 (N_22981,N_21598,N_21480);
or U22982 (N_22982,N_21204,N_21349);
nand U22983 (N_22983,N_21448,N_21461);
nor U22984 (N_22984,N_21040,N_21081);
xnor U22985 (N_22985,N_21768,N_21310);
and U22986 (N_22986,N_21617,N_21826);
xor U22987 (N_22987,N_21208,N_21516);
and U22988 (N_22988,N_21611,N_21394);
nand U22989 (N_22989,N_21159,N_21307);
nand U22990 (N_22990,N_21357,N_21200);
or U22991 (N_22991,N_21110,N_21996);
xnor U22992 (N_22992,N_21961,N_21482);
nand U22993 (N_22993,N_21184,N_21140);
nand U22994 (N_22994,N_21445,N_21489);
nand U22995 (N_22995,N_21153,N_21361);
nor U22996 (N_22996,N_21276,N_21493);
and U22997 (N_22997,N_21588,N_21763);
nand U22998 (N_22998,N_21339,N_21132);
nand U22999 (N_22999,N_21844,N_21329);
and U23000 (N_23000,N_22648,N_22961);
and U23001 (N_23001,N_22720,N_22899);
nand U23002 (N_23002,N_22384,N_22099);
nor U23003 (N_23003,N_22054,N_22319);
nand U23004 (N_23004,N_22653,N_22784);
or U23005 (N_23005,N_22218,N_22615);
xnor U23006 (N_23006,N_22925,N_22018);
nand U23007 (N_23007,N_22423,N_22242);
xnor U23008 (N_23008,N_22581,N_22589);
xnor U23009 (N_23009,N_22462,N_22832);
xor U23010 (N_23010,N_22947,N_22592);
nor U23011 (N_23011,N_22564,N_22826);
nor U23012 (N_23012,N_22183,N_22714);
nor U23013 (N_23013,N_22883,N_22862);
and U23014 (N_23014,N_22773,N_22821);
xor U23015 (N_23015,N_22071,N_22058);
xnor U23016 (N_23016,N_22020,N_22776);
nand U23017 (N_23017,N_22701,N_22199);
or U23018 (N_23018,N_22602,N_22876);
nor U23019 (N_23019,N_22979,N_22737);
xnor U23020 (N_23020,N_22822,N_22417);
xnor U23021 (N_23021,N_22493,N_22142);
or U23022 (N_23022,N_22852,N_22053);
or U23023 (N_23023,N_22579,N_22075);
xor U23024 (N_23024,N_22982,N_22061);
and U23025 (N_23025,N_22831,N_22757);
xnor U23026 (N_23026,N_22125,N_22512);
and U23027 (N_23027,N_22835,N_22953);
nor U23028 (N_23028,N_22471,N_22972);
nand U23029 (N_23029,N_22594,N_22572);
nand U23030 (N_23030,N_22435,N_22496);
nor U23031 (N_23031,N_22401,N_22238);
nand U23032 (N_23032,N_22524,N_22041);
and U23033 (N_23033,N_22726,N_22452);
or U23034 (N_23034,N_22654,N_22409);
nand U23035 (N_23035,N_22710,N_22711);
nor U23036 (N_23036,N_22984,N_22474);
nor U23037 (N_23037,N_22366,N_22480);
nor U23038 (N_23038,N_22059,N_22767);
or U23039 (N_23039,N_22208,N_22554);
nor U23040 (N_23040,N_22387,N_22671);
nor U23041 (N_23041,N_22576,N_22818);
and U23042 (N_23042,N_22312,N_22944);
or U23043 (N_23043,N_22004,N_22523);
and U23044 (N_23044,N_22731,N_22655);
nand U23045 (N_23045,N_22901,N_22519);
or U23046 (N_23046,N_22008,N_22211);
nand U23047 (N_23047,N_22151,N_22836);
xor U23048 (N_23048,N_22015,N_22611);
nand U23049 (N_23049,N_22413,N_22282);
nor U23050 (N_23050,N_22880,N_22067);
or U23051 (N_23051,N_22200,N_22422);
and U23052 (N_23052,N_22191,N_22500);
xor U23053 (N_23053,N_22190,N_22149);
or U23054 (N_23054,N_22318,N_22233);
xor U23055 (N_23055,N_22243,N_22516);
xor U23056 (N_23056,N_22341,N_22373);
xnor U23057 (N_23057,N_22303,N_22716);
or U23058 (N_23058,N_22324,N_22336);
and U23059 (N_23059,N_22884,N_22133);
and U23060 (N_23060,N_22703,N_22178);
and U23061 (N_23061,N_22839,N_22891);
and U23062 (N_23062,N_22717,N_22315);
and U23063 (N_23063,N_22355,N_22508);
and U23064 (N_23064,N_22206,N_22875);
xnor U23065 (N_23065,N_22582,N_22706);
or U23066 (N_23066,N_22718,N_22721);
or U23067 (N_23067,N_22170,N_22035);
or U23068 (N_23068,N_22158,N_22912);
nor U23069 (N_23069,N_22863,N_22106);
nor U23070 (N_23070,N_22325,N_22472);
nand U23071 (N_23071,N_22503,N_22097);
nand U23072 (N_23072,N_22692,N_22492);
nor U23073 (N_23073,N_22056,N_22269);
and U23074 (N_23074,N_22250,N_22560);
nand U23075 (N_23075,N_22381,N_22437);
and U23076 (N_23076,N_22505,N_22403);
or U23077 (N_23077,N_22569,N_22977);
nor U23078 (N_23078,N_22389,N_22956);
nand U23079 (N_23079,N_22749,N_22604);
nand U23080 (N_23080,N_22487,N_22690);
nor U23081 (N_23081,N_22394,N_22935);
nand U23082 (N_23082,N_22552,N_22301);
or U23083 (N_23083,N_22856,N_22857);
nor U23084 (N_23084,N_22478,N_22495);
and U23085 (N_23085,N_22320,N_22098);
xnor U23086 (N_23086,N_22544,N_22688);
xnor U23087 (N_23087,N_22814,N_22180);
nand U23088 (N_23088,N_22745,N_22501);
or U23089 (N_23089,N_22526,N_22625);
nor U23090 (N_23090,N_22981,N_22380);
xnor U23091 (N_23091,N_22144,N_22878);
nor U23092 (N_23092,N_22732,N_22750);
and U23093 (N_23093,N_22874,N_22386);
nor U23094 (N_23094,N_22351,N_22088);
xnor U23095 (N_23095,N_22135,N_22210);
xor U23096 (N_23096,N_22967,N_22877);
nand U23097 (N_23097,N_22370,N_22385);
nor U23098 (N_23098,N_22800,N_22825);
or U23099 (N_23099,N_22739,N_22440);
and U23100 (N_23100,N_22938,N_22165);
nor U23101 (N_23101,N_22651,N_22697);
or U23102 (N_23102,N_22795,N_22057);
nor U23103 (N_23103,N_22873,N_22477);
xnor U23104 (N_23104,N_22425,N_22382);
nor U23105 (N_23105,N_22793,N_22332);
nor U23106 (N_23106,N_22637,N_22568);
nor U23107 (N_23107,N_22963,N_22511);
nor U23108 (N_23108,N_22689,N_22545);
nor U23109 (N_23109,N_22404,N_22159);
nor U23110 (N_23110,N_22696,N_22904);
nor U23111 (N_23111,N_22127,N_22867);
xor U23112 (N_23112,N_22713,N_22284);
or U23113 (N_23113,N_22743,N_22712);
or U23114 (N_23114,N_22675,N_22755);
and U23115 (N_23115,N_22618,N_22473);
xor U23116 (N_23116,N_22194,N_22702);
nor U23117 (N_23117,N_22136,N_22920);
nor U23118 (N_23118,N_22065,N_22890);
nor U23119 (N_23119,N_22960,N_22796);
nor U23120 (N_23120,N_22761,N_22283);
nor U23121 (N_23121,N_22104,N_22217);
or U23122 (N_23122,N_22343,N_22350);
nand U23123 (N_23123,N_22114,N_22410);
nor U23124 (N_23124,N_22570,N_22286);
xnor U23125 (N_23125,N_22590,N_22486);
xnor U23126 (N_23126,N_22276,N_22682);
nand U23127 (N_23127,N_22605,N_22102);
xnor U23128 (N_23128,N_22415,N_22305);
nor U23129 (N_23129,N_22879,N_22215);
or U23130 (N_23130,N_22117,N_22887);
nand U23131 (N_23131,N_22823,N_22946);
nand U23132 (N_23132,N_22778,N_22416);
or U23133 (N_23133,N_22663,N_22804);
nor U23134 (N_23134,N_22620,N_22518);
nor U23135 (N_23135,N_22640,N_22976);
xor U23136 (N_23136,N_22771,N_22265);
xnor U23137 (N_23137,N_22608,N_22715);
nor U23138 (N_23138,N_22521,N_22596);
nand U23139 (N_23139,N_22274,N_22816);
nand U23140 (N_23140,N_22288,N_22006);
xor U23141 (N_23141,N_22230,N_22817);
nor U23142 (N_23142,N_22859,N_22534);
nor U23143 (N_23143,N_22695,N_22528);
and U23144 (N_23144,N_22644,N_22687);
or U23145 (N_23145,N_22583,N_22834);
and U23146 (N_23146,N_22353,N_22331);
nand U23147 (N_23147,N_22824,N_22709);
and U23148 (N_23148,N_22820,N_22073);
nor U23149 (N_23149,N_22334,N_22786);
or U23150 (N_23150,N_22672,N_22851);
nor U23151 (N_23151,N_22257,N_22803);
xnor U23152 (N_23152,N_22236,N_22293);
xor U23153 (N_23153,N_22089,N_22270);
xor U23154 (N_23154,N_22727,N_22011);
or U23155 (N_23155,N_22064,N_22335);
xor U23156 (N_23156,N_22617,N_22326);
or U23157 (N_23157,N_22221,N_22549);
nand U23158 (N_23158,N_22141,N_22992);
nor U23159 (N_23159,N_22337,N_22461);
and U23160 (N_23160,N_22012,N_22705);
or U23161 (N_23161,N_22321,N_22153);
or U23162 (N_23162,N_22076,N_22150);
or U23163 (N_23163,N_22950,N_22077);
nor U23164 (N_23164,N_22886,N_22971);
nor U23165 (N_23165,N_22533,N_22551);
and U23166 (N_23166,N_22974,N_22201);
and U23167 (N_23167,N_22844,N_22996);
xnor U23168 (N_23168,N_22694,N_22391);
nor U23169 (N_23169,N_22154,N_22498);
nor U23170 (N_23170,N_22264,N_22550);
nand U23171 (N_23171,N_22898,N_22223);
nor U23172 (N_23172,N_22686,N_22476);
or U23173 (N_23173,N_22155,N_22978);
nor U23174 (N_23174,N_22148,N_22542);
nor U23175 (N_23175,N_22787,N_22484);
xnor U23176 (N_23176,N_22197,N_22724);
or U23177 (N_23177,N_22402,N_22042);
or U23178 (N_23178,N_22556,N_22966);
or U23179 (N_23179,N_22225,N_22311);
nand U23180 (N_23180,N_22063,N_22198);
or U23181 (N_23181,N_22989,N_22371);
xnor U23182 (N_23182,N_22555,N_22735);
nor U23183 (N_23183,N_22628,N_22419);
nand U23184 (N_23184,N_22802,N_22289);
xnor U23185 (N_23185,N_22147,N_22575);
nand U23186 (N_23186,N_22050,N_22850);
and U23187 (N_23187,N_22455,N_22490);
xor U23188 (N_23188,N_22454,N_22219);
or U23189 (N_23189,N_22685,N_22189);
nor U23190 (N_23190,N_22203,N_22424);
nor U23191 (N_23191,N_22509,N_22108);
xor U23192 (N_23192,N_22143,N_22708);
xnor U23193 (N_23193,N_22662,N_22788);
or U23194 (N_23194,N_22954,N_22226);
or U23195 (N_23195,N_22139,N_22295);
or U23196 (N_23196,N_22300,N_22122);
xnor U23197 (N_23197,N_22043,N_22801);
nand U23198 (N_23198,N_22600,N_22782);
nor U23199 (N_23199,N_22434,N_22532);
and U23200 (N_23200,N_22306,N_22613);
and U23201 (N_23201,N_22182,N_22680);
and U23202 (N_23202,N_22999,N_22845);
or U23203 (N_23203,N_22634,N_22864);
xnor U23204 (N_23204,N_22038,N_22291);
and U23205 (N_23205,N_22016,N_22779);
or U23206 (N_23206,N_22007,N_22441);
xnor U23207 (N_23207,N_22917,N_22399);
xnor U23208 (N_23208,N_22345,N_22955);
nand U23209 (N_23209,N_22362,N_22895);
or U23210 (N_23210,N_22936,N_22196);
or U23211 (N_23211,N_22458,N_22900);
xnor U23212 (N_23212,N_22748,N_22268);
and U23213 (N_23213,N_22297,N_22805);
nand U23214 (N_23214,N_22445,N_22888);
nor U23215 (N_23215,N_22418,N_22964);
nand U23216 (N_23216,N_22517,N_22892);
nand U23217 (N_23217,N_22298,N_22681);
nor U23218 (N_23218,N_22798,N_22623);
xnor U23219 (N_23219,N_22031,N_22673);
xor U23220 (N_23220,N_22930,N_22024);
and U23221 (N_23221,N_22991,N_22388);
nand U23222 (N_23222,N_22941,N_22429);
xnor U23223 (N_23223,N_22442,N_22376);
xnor U23224 (N_23224,N_22645,N_22624);
nor U23225 (N_23225,N_22780,N_22965);
xnor U23226 (N_23226,N_22395,N_22292);
xor U23227 (N_23227,N_22329,N_22111);
or U23228 (N_23228,N_22338,N_22535);
and U23229 (N_23229,N_22513,N_22040);
or U23230 (N_23230,N_22195,N_22421);
or U23231 (N_23231,N_22449,N_22174);
and U23232 (N_23232,N_22833,N_22010);
and U23233 (N_23233,N_22907,N_22157);
and U23234 (N_23234,N_22095,N_22668);
or U23235 (N_23235,N_22456,N_22033);
nand U23236 (N_23236,N_22094,N_22485);
or U23237 (N_23237,N_22760,N_22475);
nand U23238 (N_23238,N_22746,N_22083);
or U23239 (N_23239,N_22842,N_22866);
xor U23240 (N_23240,N_22765,N_22164);
or U23241 (N_23241,N_22599,N_22598);
xnor U23242 (N_23242,N_22168,N_22248);
xor U23243 (N_23243,N_22910,N_22553);
and U23244 (N_23244,N_22664,N_22631);
or U23245 (N_23245,N_22251,N_22412);
or U23246 (N_23246,N_22121,N_22667);
nor U23247 (N_23247,N_22356,N_22893);
or U23248 (N_23248,N_22214,N_22392);
nand U23249 (N_23249,N_22614,N_22633);
or U23250 (N_23250,N_22060,N_22903);
nor U23251 (N_23251,N_22940,N_22411);
and U23252 (N_23252,N_22129,N_22497);
xor U23253 (N_23253,N_22138,N_22548);
nor U23254 (N_23254,N_22536,N_22530);
nor U23255 (N_23255,N_22220,N_22632);
nand U23256 (N_23256,N_22998,N_22584);
nand U23257 (N_23257,N_22252,N_22034);
or U23258 (N_23258,N_22278,N_22086);
nor U23259 (N_23259,N_22256,N_22557);
nand U23260 (N_23260,N_22656,N_22647);
and U23261 (N_23261,N_22665,N_22162);
and U23262 (N_23262,N_22048,N_22047);
nand U23263 (N_23263,N_22641,N_22578);
nand U23264 (N_23264,N_22995,N_22489);
nor U23265 (N_23265,N_22819,N_22408);
nand U23266 (N_23266,N_22453,N_22317);
nand U23267 (N_23267,N_22116,N_22464);
or U23268 (N_23268,N_22729,N_22593);
nor U23269 (N_23269,N_22541,N_22650);
and U23270 (N_23270,N_22467,N_22302);
nor U23271 (N_23271,N_22091,N_22255);
xnor U23272 (N_23272,N_22860,N_22450);
and U23273 (N_23273,N_22934,N_22830);
xor U23274 (N_23274,N_22032,N_22333);
nor U23275 (N_23275,N_22186,N_22433);
nand U23276 (N_23276,N_22277,N_22175);
and U23277 (N_23277,N_22968,N_22307);
and U23278 (N_23278,N_22591,N_22567);
nand U23279 (N_23279,N_22393,N_22885);
nand U23280 (N_23280,N_22342,N_22296);
nand U23281 (N_23281,N_22751,N_22023);
nor U23282 (N_23282,N_22101,N_22027);
nand U23283 (N_23283,N_22082,N_22759);
xor U23284 (N_23284,N_22428,N_22616);
nor U23285 (N_23285,N_22908,N_22267);
nor U23286 (N_23286,N_22357,N_22962);
or U23287 (N_23287,N_22514,N_22213);
xnor U23288 (N_23288,N_22110,N_22853);
and U23289 (N_23289,N_22595,N_22398);
nor U23290 (N_23290,N_22112,N_22290);
nor U23291 (N_23291,N_22679,N_22074);
xor U23292 (N_23292,N_22897,N_22085);
nor U23293 (N_23293,N_22754,N_22407);
or U23294 (N_23294,N_22205,N_22889);
or U23295 (N_23295,N_22610,N_22843);
xor U23296 (N_23296,N_22466,N_22084);
or U23297 (N_23297,N_22271,N_22914);
or U23298 (N_23298,N_22093,N_22369);
xnor U23299 (N_23299,N_22520,N_22014);
nand U23300 (N_23300,N_22119,N_22942);
xnor U23301 (N_23301,N_22451,N_22118);
nor U23302 (N_23302,N_22738,N_22444);
or U23303 (N_23303,N_22367,N_22601);
nor U23304 (N_23304,N_22540,N_22349);
xnor U23305 (N_23305,N_22799,N_22192);
xor U23306 (N_23306,N_22021,N_22529);
nand U23307 (N_23307,N_22609,N_22522);
nand U23308 (N_23308,N_22330,N_22510);
nand U23309 (N_23309,N_22565,N_22896);
and U23310 (N_23310,N_22022,N_22868);
or U23311 (N_23311,N_22629,N_22163);
xor U23312 (N_23312,N_22177,N_22109);
or U23313 (N_23313,N_22988,N_22502);
or U23314 (N_23314,N_22669,N_22588);
xor U23315 (N_23315,N_22068,N_22612);
xor U23316 (N_23316,N_22725,N_22400);
nor U23317 (N_23317,N_22100,N_22239);
nor U23318 (N_23318,N_22137,N_22287);
or U23319 (N_23319,N_22915,N_22927);
nand U23320 (N_23320,N_22003,N_22132);
nand U23321 (N_23321,N_22310,N_22921);
nand U23322 (N_23322,N_22660,N_22911);
or U23323 (N_23323,N_22052,N_22986);
xnor U23324 (N_23324,N_22092,N_22728);
or U23325 (N_23325,N_22865,N_22531);
and U23326 (N_23326,N_22483,N_22987);
and U23327 (N_23327,N_22202,N_22126);
nor U23328 (N_23328,N_22081,N_22849);
xnor U23329 (N_23329,N_22753,N_22546);
xor U23330 (N_23330,N_22676,N_22090);
xnor U23331 (N_23331,N_22146,N_22113);
xor U23332 (N_23332,N_22973,N_22432);
or U23333 (N_23333,N_22263,N_22002);
nand U23334 (N_23334,N_22327,N_22062);
or U23335 (N_23335,N_22229,N_22249);
and U23336 (N_23336,N_22469,N_22313);
or U23337 (N_23337,N_22247,N_22375);
nor U23338 (N_23338,N_22235,N_22993);
or U23339 (N_23339,N_22231,N_22772);
nor U23340 (N_23340,N_22871,N_22430);
nor U23341 (N_23341,N_22752,N_22919);
and U23342 (N_23342,N_22931,N_22698);
nor U23343 (N_23343,N_22161,N_22639);
nor U23344 (N_23344,N_22756,N_22131);
and U23345 (N_23345,N_22515,N_22358);
nor U23346 (N_23346,N_22029,N_22273);
nand U23347 (N_23347,N_22619,N_22758);
nand U23348 (N_23348,N_22446,N_22246);
xor U23349 (N_23349,N_22783,N_22363);
or U23350 (N_23350,N_22436,N_22630);
xor U23351 (N_23351,N_22080,N_22806);
nand U23352 (N_23352,N_22294,N_22079);
nor U23353 (N_23353,N_22228,N_22790);
nand U23354 (N_23354,N_22019,N_22847);
xor U23355 (N_23355,N_22348,N_22427);
nor U23356 (N_23356,N_22580,N_22809);
nor U23357 (N_23357,N_22187,N_22506);
nor U23358 (N_23358,N_22468,N_22747);
nand U23359 (N_23359,N_22244,N_22176);
or U23360 (N_23360,N_22722,N_22670);
and U23361 (N_23361,N_22744,N_22969);
xnor U23362 (N_23362,N_22789,N_22443);
xor U23363 (N_23363,N_22115,N_22431);
nand U23364 (N_23364,N_22959,N_22426);
nand U23365 (N_23365,N_22078,N_22636);
or U23366 (N_23366,N_22145,N_22087);
and U23367 (N_23367,N_22571,N_22627);
and U23368 (N_23368,N_22559,N_22241);
and U23369 (N_23369,N_22561,N_22837);
nor U23370 (N_23370,N_22922,N_22339);
and U23371 (N_23371,N_22212,N_22028);
and U23372 (N_23372,N_22237,N_22488);
xor U23373 (N_23373,N_22543,N_22829);
and U23374 (N_23374,N_22813,N_22128);
nor U23375 (N_23375,N_22621,N_22704);
or U23376 (N_23376,N_22828,N_22794);
and U23377 (N_23377,N_22952,N_22691);
or U23378 (N_23378,N_22929,N_22460);
nor U23379 (N_23379,N_22649,N_22396);
nor U23380 (N_23380,N_22207,N_22909);
nand U23381 (N_23381,N_22674,N_22957);
or U23382 (N_23382,N_22323,N_22933);
nor U23383 (N_23383,N_22005,N_22360);
and U23384 (N_23384,N_22626,N_22245);
nor U23385 (N_23385,N_22308,N_22285);
nand U23386 (N_23386,N_22768,N_22659);
nor U23387 (N_23387,N_22525,N_22894);
nor U23388 (N_23388,N_22538,N_22377);
and U23389 (N_23389,N_22924,N_22763);
nor U23390 (N_23390,N_22167,N_22368);
xor U23391 (N_23391,N_22438,N_22181);
or U23392 (N_23392,N_22587,N_22171);
nand U23393 (N_23393,N_22766,N_22209);
xor U23394 (N_23394,N_22140,N_22983);
or U23395 (N_23395,N_22039,N_22643);
nand U23396 (N_23396,N_22470,N_22791);
and U23397 (N_23397,N_22906,N_22072);
or U23398 (N_23398,N_22103,N_22328);
and U23399 (N_23399,N_22945,N_22025);
or U23400 (N_23400,N_22785,N_22741);
and U23401 (N_23401,N_22719,N_22642);
xnor U23402 (N_23402,N_22390,N_22537);
or U23403 (N_23403,N_22951,N_22266);
and U23404 (N_23404,N_22352,N_22797);
or U23405 (N_23405,N_22262,N_22902);
nand U23406 (N_23406,N_22232,N_22044);
and U23407 (N_23407,N_22562,N_22359);
nand U23408 (N_23408,N_22405,N_22185);
or U23409 (N_23409,N_22397,N_22037);
nand U23410 (N_23410,N_22808,N_22734);
nor U23411 (N_23411,N_22566,N_22279);
nor U23412 (N_23412,N_22275,N_22361);
or U23413 (N_23413,N_22603,N_22046);
and U23414 (N_23414,N_22272,N_22260);
xnor U23415 (N_23415,N_22928,N_22193);
xor U23416 (N_23416,N_22499,N_22000);
and U23417 (N_23417,N_22507,N_22130);
and U23418 (N_23418,N_22573,N_22120);
xnor U23419 (N_23419,N_22314,N_22638);
or U23420 (N_23420,N_22563,N_22253);
and U23421 (N_23421,N_22216,N_22346);
xnor U23422 (N_23422,N_22558,N_22848);
and U23423 (N_23423,N_22762,N_22775);
nor U23424 (N_23424,N_22070,N_22152);
or U23425 (N_23425,N_22457,N_22280);
nand U23426 (N_23426,N_22678,N_22134);
or U23427 (N_23427,N_22322,N_22657);
xor U23428 (N_23428,N_22465,N_22838);
nor U23429 (N_23429,N_22870,N_22365);
and U23430 (N_23430,N_22036,N_22166);
and U23431 (N_23431,N_22316,N_22420);
nor U23432 (N_23432,N_22309,N_22693);
xor U23433 (N_23433,N_22869,N_22736);
nor U23434 (N_23434,N_22013,N_22069);
nor U23435 (N_23435,N_22622,N_22840);
or U23436 (N_23436,N_22658,N_22700);
and U23437 (N_23437,N_22970,N_22652);
nand U23438 (N_23438,N_22855,N_22009);
and U23439 (N_23439,N_22261,N_22607);
nor U23440 (N_23440,N_22049,N_22354);
nand U23441 (N_23441,N_22224,N_22222);
or U23442 (N_23442,N_22574,N_22939);
nor U23443 (N_23443,N_22406,N_22344);
or U23444 (N_23444,N_22447,N_22740);
or U23445 (N_23445,N_22188,N_22124);
and U23446 (N_23446,N_22846,N_22539);
or U23447 (N_23447,N_22764,N_22107);
xnor U23448 (N_23448,N_22494,N_22123);
xor U23449 (N_23449,N_22975,N_22932);
or U23450 (N_23450,N_22372,N_22913);
nand U23451 (N_23451,N_22234,N_22527);
nand U23452 (N_23452,N_22586,N_22807);
xnor U23453 (N_23453,N_22730,N_22105);
and U23454 (N_23454,N_22707,N_22227);
and U23455 (N_23455,N_22666,N_22949);
and U23456 (N_23456,N_22854,N_22479);
nand U23457 (N_23457,N_22364,N_22918);
and U23458 (N_23458,N_22179,N_22905);
and U23459 (N_23459,N_22769,N_22547);
and U23460 (N_23460,N_22204,N_22299);
or U23461 (N_23461,N_22872,N_22439);
nand U23462 (N_23462,N_22184,N_22781);
xor U23463 (N_23463,N_22777,N_22937);
nand U23464 (N_23464,N_22684,N_22017);
and U23465 (N_23465,N_22943,N_22926);
or U23466 (N_23466,N_22774,N_22051);
and U23467 (N_23467,N_22001,N_22378);
and U23468 (N_23468,N_22683,N_22414);
nand U23469 (N_23469,N_22096,N_22958);
nor U23470 (N_23470,N_22948,N_22045);
nand U23471 (N_23471,N_22448,N_22585);
xor U23472 (N_23472,N_22459,N_22923);
nor U23473 (N_23473,N_22026,N_22858);
nand U23474 (N_23474,N_22985,N_22066);
xor U23475 (N_23475,N_22173,N_22916);
xnor U23476 (N_23476,N_22463,N_22990);
nand U23477 (N_23477,N_22172,N_22481);
and U23478 (N_23478,N_22994,N_22254);
xnor U23479 (N_23479,N_22258,N_22055);
and U23480 (N_23480,N_22030,N_22881);
nor U23481 (N_23481,N_22792,N_22661);
nand U23482 (N_23482,N_22733,N_22160);
and U23483 (N_23483,N_22304,N_22340);
nor U23484 (N_23484,N_22504,N_22882);
or U23485 (N_23485,N_22723,N_22812);
or U23486 (N_23486,N_22374,N_22379);
or U23487 (N_23487,N_22677,N_22347);
nand U23488 (N_23488,N_22597,N_22699);
or U23489 (N_23489,N_22577,N_22240);
and U23490 (N_23490,N_22770,N_22281);
or U23491 (N_23491,N_22742,N_22482);
or U23492 (N_23492,N_22491,N_22827);
xor U23493 (N_23493,N_22861,N_22169);
nor U23494 (N_23494,N_22811,N_22646);
and U23495 (N_23495,N_22606,N_22841);
and U23496 (N_23496,N_22383,N_22997);
and U23497 (N_23497,N_22635,N_22156);
or U23498 (N_23498,N_22815,N_22980);
and U23499 (N_23499,N_22259,N_22810);
or U23500 (N_23500,N_22510,N_22278);
or U23501 (N_23501,N_22663,N_22682);
nand U23502 (N_23502,N_22412,N_22047);
or U23503 (N_23503,N_22481,N_22318);
and U23504 (N_23504,N_22040,N_22151);
and U23505 (N_23505,N_22801,N_22387);
and U23506 (N_23506,N_22691,N_22228);
nand U23507 (N_23507,N_22622,N_22432);
xor U23508 (N_23508,N_22593,N_22856);
nand U23509 (N_23509,N_22713,N_22441);
xor U23510 (N_23510,N_22008,N_22350);
nand U23511 (N_23511,N_22255,N_22655);
or U23512 (N_23512,N_22458,N_22141);
xnor U23513 (N_23513,N_22051,N_22684);
xnor U23514 (N_23514,N_22237,N_22592);
nand U23515 (N_23515,N_22025,N_22163);
and U23516 (N_23516,N_22945,N_22055);
and U23517 (N_23517,N_22179,N_22205);
and U23518 (N_23518,N_22616,N_22264);
and U23519 (N_23519,N_22360,N_22114);
and U23520 (N_23520,N_22275,N_22405);
xor U23521 (N_23521,N_22025,N_22606);
or U23522 (N_23522,N_22357,N_22778);
or U23523 (N_23523,N_22814,N_22941);
xnor U23524 (N_23524,N_22344,N_22519);
or U23525 (N_23525,N_22632,N_22022);
xnor U23526 (N_23526,N_22710,N_22495);
and U23527 (N_23527,N_22104,N_22558);
or U23528 (N_23528,N_22239,N_22498);
xor U23529 (N_23529,N_22550,N_22565);
and U23530 (N_23530,N_22031,N_22685);
nand U23531 (N_23531,N_22241,N_22986);
nor U23532 (N_23532,N_22561,N_22915);
or U23533 (N_23533,N_22587,N_22548);
and U23534 (N_23534,N_22046,N_22751);
or U23535 (N_23535,N_22757,N_22217);
nor U23536 (N_23536,N_22431,N_22585);
nand U23537 (N_23537,N_22824,N_22999);
nand U23538 (N_23538,N_22511,N_22952);
or U23539 (N_23539,N_22321,N_22885);
xnor U23540 (N_23540,N_22397,N_22875);
nand U23541 (N_23541,N_22790,N_22627);
or U23542 (N_23542,N_22989,N_22141);
nor U23543 (N_23543,N_22315,N_22959);
nor U23544 (N_23544,N_22782,N_22613);
nor U23545 (N_23545,N_22152,N_22892);
and U23546 (N_23546,N_22752,N_22990);
and U23547 (N_23547,N_22724,N_22441);
nand U23548 (N_23548,N_22417,N_22280);
xnor U23549 (N_23549,N_22698,N_22279);
nand U23550 (N_23550,N_22183,N_22965);
and U23551 (N_23551,N_22505,N_22467);
nor U23552 (N_23552,N_22193,N_22237);
or U23553 (N_23553,N_22240,N_22068);
or U23554 (N_23554,N_22682,N_22900);
or U23555 (N_23555,N_22719,N_22196);
nor U23556 (N_23556,N_22623,N_22168);
xor U23557 (N_23557,N_22500,N_22092);
xor U23558 (N_23558,N_22617,N_22478);
nor U23559 (N_23559,N_22304,N_22245);
and U23560 (N_23560,N_22758,N_22197);
nor U23561 (N_23561,N_22528,N_22198);
xor U23562 (N_23562,N_22465,N_22549);
and U23563 (N_23563,N_22059,N_22324);
nor U23564 (N_23564,N_22690,N_22175);
xor U23565 (N_23565,N_22481,N_22577);
xnor U23566 (N_23566,N_22522,N_22566);
nor U23567 (N_23567,N_22181,N_22602);
xor U23568 (N_23568,N_22749,N_22011);
and U23569 (N_23569,N_22435,N_22672);
and U23570 (N_23570,N_22089,N_22623);
or U23571 (N_23571,N_22409,N_22397);
or U23572 (N_23572,N_22956,N_22115);
or U23573 (N_23573,N_22807,N_22637);
nor U23574 (N_23574,N_22709,N_22129);
and U23575 (N_23575,N_22717,N_22761);
xnor U23576 (N_23576,N_22752,N_22518);
and U23577 (N_23577,N_22266,N_22528);
nand U23578 (N_23578,N_22558,N_22766);
xor U23579 (N_23579,N_22715,N_22197);
and U23580 (N_23580,N_22270,N_22423);
xor U23581 (N_23581,N_22021,N_22245);
nor U23582 (N_23582,N_22570,N_22750);
nor U23583 (N_23583,N_22594,N_22344);
nand U23584 (N_23584,N_22858,N_22541);
nand U23585 (N_23585,N_22163,N_22031);
and U23586 (N_23586,N_22811,N_22203);
nand U23587 (N_23587,N_22456,N_22107);
xor U23588 (N_23588,N_22450,N_22624);
nand U23589 (N_23589,N_22673,N_22772);
or U23590 (N_23590,N_22568,N_22866);
nand U23591 (N_23591,N_22369,N_22774);
xor U23592 (N_23592,N_22523,N_22768);
xor U23593 (N_23593,N_22443,N_22418);
nand U23594 (N_23594,N_22752,N_22390);
nor U23595 (N_23595,N_22895,N_22405);
nor U23596 (N_23596,N_22149,N_22440);
or U23597 (N_23597,N_22808,N_22242);
xnor U23598 (N_23598,N_22286,N_22644);
and U23599 (N_23599,N_22499,N_22821);
nand U23600 (N_23600,N_22199,N_22848);
nor U23601 (N_23601,N_22413,N_22757);
xnor U23602 (N_23602,N_22328,N_22360);
nand U23603 (N_23603,N_22563,N_22665);
nor U23604 (N_23604,N_22341,N_22627);
or U23605 (N_23605,N_22264,N_22305);
nor U23606 (N_23606,N_22072,N_22372);
or U23607 (N_23607,N_22949,N_22288);
or U23608 (N_23608,N_22545,N_22343);
xnor U23609 (N_23609,N_22693,N_22715);
and U23610 (N_23610,N_22771,N_22531);
nor U23611 (N_23611,N_22890,N_22465);
and U23612 (N_23612,N_22161,N_22972);
or U23613 (N_23613,N_22755,N_22825);
xor U23614 (N_23614,N_22106,N_22455);
or U23615 (N_23615,N_22055,N_22124);
and U23616 (N_23616,N_22964,N_22745);
or U23617 (N_23617,N_22572,N_22524);
nand U23618 (N_23618,N_22359,N_22535);
or U23619 (N_23619,N_22464,N_22033);
nand U23620 (N_23620,N_22079,N_22839);
or U23621 (N_23621,N_22366,N_22774);
or U23622 (N_23622,N_22800,N_22158);
or U23623 (N_23623,N_22587,N_22432);
xnor U23624 (N_23624,N_22485,N_22959);
nand U23625 (N_23625,N_22881,N_22814);
nand U23626 (N_23626,N_22937,N_22541);
nand U23627 (N_23627,N_22859,N_22212);
nand U23628 (N_23628,N_22724,N_22696);
nor U23629 (N_23629,N_22573,N_22726);
and U23630 (N_23630,N_22118,N_22008);
nand U23631 (N_23631,N_22083,N_22143);
nand U23632 (N_23632,N_22040,N_22246);
nand U23633 (N_23633,N_22975,N_22567);
or U23634 (N_23634,N_22728,N_22077);
nor U23635 (N_23635,N_22861,N_22176);
and U23636 (N_23636,N_22172,N_22342);
or U23637 (N_23637,N_22866,N_22659);
and U23638 (N_23638,N_22672,N_22612);
or U23639 (N_23639,N_22645,N_22965);
and U23640 (N_23640,N_22314,N_22137);
nand U23641 (N_23641,N_22742,N_22036);
and U23642 (N_23642,N_22487,N_22434);
or U23643 (N_23643,N_22866,N_22367);
nor U23644 (N_23644,N_22065,N_22456);
or U23645 (N_23645,N_22730,N_22815);
nand U23646 (N_23646,N_22238,N_22767);
nand U23647 (N_23647,N_22921,N_22822);
nand U23648 (N_23648,N_22972,N_22879);
nor U23649 (N_23649,N_22748,N_22314);
or U23650 (N_23650,N_22723,N_22151);
nor U23651 (N_23651,N_22522,N_22423);
nor U23652 (N_23652,N_22773,N_22115);
xor U23653 (N_23653,N_22031,N_22232);
and U23654 (N_23654,N_22629,N_22613);
nand U23655 (N_23655,N_22817,N_22711);
xnor U23656 (N_23656,N_22569,N_22660);
xnor U23657 (N_23657,N_22053,N_22986);
and U23658 (N_23658,N_22864,N_22356);
xnor U23659 (N_23659,N_22623,N_22165);
xor U23660 (N_23660,N_22566,N_22153);
and U23661 (N_23661,N_22654,N_22250);
and U23662 (N_23662,N_22625,N_22995);
nor U23663 (N_23663,N_22619,N_22865);
nor U23664 (N_23664,N_22718,N_22892);
or U23665 (N_23665,N_22408,N_22315);
or U23666 (N_23666,N_22131,N_22527);
nor U23667 (N_23667,N_22829,N_22715);
or U23668 (N_23668,N_22816,N_22723);
nand U23669 (N_23669,N_22456,N_22022);
or U23670 (N_23670,N_22653,N_22676);
xor U23671 (N_23671,N_22885,N_22774);
xnor U23672 (N_23672,N_22642,N_22061);
nand U23673 (N_23673,N_22112,N_22123);
xor U23674 (N_23674,N_22198,N_22303);
or U23675 (N_23675,N_22100,N_22492);
and U23676 (N_23676,N_22034,N_22045);
or U23677 (N_23677,N_22350,N_22726);
and U23678 (N_23678,N_22382,N_22771);
xnor U23679 (N_23679,N_22157,N_22068);
or U23680 (N_23680,N_22541,N_22605);
xor U23681 (N_23681,N_22222,N_22034);
and U23682 (N_23682,N_22547,N_22652);
or U23683 (N_23683,N_22860,N_22572);
and U23684 (N_23684,N_22716,N_22126);
nor U23685 (N_23685,N_22450,N_22811);
or U23686 (N_23686,N_22407,N_22507);
and U23687 (N_23687,N_22743,N_22884);
and U23688 (N_23688,N_22877,N_22240);
xor U23689 (N_23689,N_22347,N_22228);
xnor U23690 (N_23690,N_22792,N_22691);
and U23691 (N_23691,N_22128,N_22213);
nand U23692 (N_23692,N_22785,N_22773);
nor U23693 (N_23693,N_22699,N_22817);
xor U23694 (N_23694,N_22162,N_22999);
nand U23695 (N_23695,N_22278,N_22499);
and U23696 (N_23696,N_22618,N_22954);
or U23697 (N_23697,N_22534,N_22466);
xnor U23698 (N_23698,N_22203,N_22282);
or U23699 (N_23699,N_22005,N_22461);
nor U23700 (N_23700,N_22218,N_22465);
nand U23701 (N_23701,N_22894,N_22418);
nor U23702 (N_23702,N_22884,N_22536);
and U23703 (N_23703,N_22602,N_22281);
or U23704 (N_23704,N_22794,N_22281);
and U23705 (N_23705,N_22210,N_22266);
and U23706 (N_23706,N_22659,N_22951);
xor U23707 (N_23707,N_22826,N_22513);
xnor U23708 (N_23708,N_22626,N_22653);
nand U23709 (N_23709,N_22967,N_22243);
and U23710 (N_23710,N_22729,N_22330);
and U23711 (N_23711,N_22644,N_22248);
and U23712 (N_23712,N_22679,N_22503);
nand U23713 (N_23713,N_22351,N_22791);
nor U23714 (N_23714,N_22488,N_22509);
nor U23715 (N_23715,N_22605,N_22997);
nand U23716 (N_23716,N_22495,N_22648);
and U23717 (N_23717,N_22511,N_22793);
nand U23718 (N_23718,N_22632,N_22703);
xnor U23719 (N_23719,N_22097,N_22861);
nand U23720 (N_23720,N_22138,N_22850);
or U23721 (N_23721,N_22909,N_22728);
nand U23722 (N_23722,N_22102,N_22528);
xor U23723 (N_23723,N_22845,N_22504);
xor U23724 (N_23724,N_22333,N_22231);
nand U23725 (N_23725,N_22109,N_22758);
nor U23726 (N_23726,N_22862,N_22296);
xor U23727 (N_23727,N_22769,N_22244);
xor U23728 (N_23728,N_22957,N_22350);
or U23729 (N_23729,N_22440,N_22172);
nand U23730 (N_23730,N_22014,N_22595);
nor U23731 (N_23731,N_22814,N_22409);
and U23732 (N_23732,N_22744,N_22196);
or U23733 (N_23733,N_22744,N_22909);
nor U23734 (N_23734,N_22080,N_22437);
and U23735 (N_23735,N_22765,N_22283);
nor U23736 (N_23736,N_22108,N_22435);
and U23737 (N_23737,N_22513,N_22554);
nor U23738 (N_23738,N_22553,N_22545);
nor U23739 (N_23739,N_22421,N_22068);
and U23740 (N_23740,N_22392,N_22029);
nand U23741 (N_23741,N_22742,N_22707);
xor U23742 (N_23742,N_22669,N_22534);
or U23743 (N_23743,N_22922,N_22031);
nand U23744 (N_23744,N_22681,N_22225);
or U23745 (N_23745,N_22808,N_22601);
or U23746 (N_23746,N_22184,N_22014);
or U23747 (N_23747,N_22144,N_22526);
nand U23748 (N_23748,N_22211,N_22751);
nand U23749 (N_23749,N_22869,N_22753);
nand U23750 (N_23750,N_22039,N_22260);
xnor U23751 (N_23751,N_22303,N_22644);
or U23752 (N_23752,N_22458,N_22658);
xnor U23753 (N_23753,N_22149,N_22051);
and U23754 (N_23754,N_22559,N_22868);
and U23755 (N_23755,N_22178,N_22368);
xor U23756 (N_23756,N_22667,N_22107);
xnor U23757 (N_23757,N_22941,N_22527);
or U23758 (N_23758,N_22676,N_22791);
nor U23759 (N_23759,N_22682,N_22547);
nand U23760 (N_23760,N_22780,N_22210);
xor U23761 (N_23761,N_22457,N_22843);
or U23762 (N_23762,N_22966,N_22691);
nand U23763 (N_23763,N_22057,N_22120);
nor U23764 (N_23764,N_22263,N_22059);
and U23765 (N_23765,N_22487,N_22152);
xnor U23766 (N_23766,N_22467,N_22927);
xnor U23767 (N_23767,N_22243,N_22019);
and U23768 (N_23768,N_22613,N_22670);
nor U23769 (N_23769,N_22363,N_22444);
nor U23770 (N_23770,N_22467,N_22596);
nor U23771 (N_23771,N_22650,N_22885);
nand U23772 (N_23772,N_22620,N_22393);
xor U23773 (N_23773,N_22880,N_22591);
and U23774 (N_23774,N_22649,N_22492);
or U23775 (N_23775,N_22859,N_22402);
xnor U23776 (N_23776,N_22666,N_22503);
nand U23777 (N_23777,N_22711,N_22473);
xnor U23778 (N_23778,N_22584,N_22241);
and U23779 (N_23779,N_22025,N_22736);
xor U23780 (N_23780,N_22094,N_22351);
nand U23781 (N_23781,N_22872,N_22783);
and U23782 (N_23782,N_22092,N_22042);
or U23783 (N_23783,N_22517,N_22607);
nand U23784 (N_23784,N_22473,N_22534);
xnor U23785 (N_23785,N_22819,N_22822);
nor U23786 (N_23786,N_22109,N_22820);
and U23787 (N_23787,N_22849,N_22728);
xor U23788 (N_23788,N_22052,N_22560);
and U23789 (N_23789,N_22093,N_22763);
and U23790 (N_23790,N_22024,N_22373);
or U23791 (N_23791,N_22096,N_22550);
nand U23792 (N_23792,N_22600,N_22125);
nor U23793 (N_23793,N_22815,N_22473);
or U23794 (N_23794,N_22712,N_22463);
or U23795 (N_23795,N_22502,N_22737);
xnor U23796 (N_23796,N_22801,N_22465);
or U23797 (N_23797,N_22657,N_22748);
and U23798 (N_23798,N_22004,N_22613);
nand U23799 (N_23799,N_22363,N_22011);
nand U23800 (N_23800,N_22746,N_22706);
or U23801 (N_23801,N_22255,N_22230);
xnor U23802 (N_23802,N_22672,N_22998);
and U23803 (N_23803,N_22523,N_22295);
nor U23804 (N_23804,N_22113,N_22852);
or U23805 (N_23805,N_22896,N_22169);
nand U23806 (N_23806,N_22970,N_22137);
and U23807 (N_23807,N_22128,N_22169);
nor U23808 (N_23808,N_22038,N_22220);
nor U23809 (N_23809,N_22164,N_22701);
and U23810 (N_23810,N_22119,N_22142);
nor U23811 (N_23811,N_22528,N_22225);
and U23812 (N_23812,N_22150,N_22390);
or U23813 (N_23813,N_22665,N_22411);
and U23814 (N_23814,N_22464,N_22958);
nand U23815 (N_23815,N_22035,N_22875);
nor U23816 (N_23816,N_22148,N_22192);
and U23817 (N_23817,N_22069,N_22554);
nor U23818 (N_23818,N_22871,N_22197);
or U23819 (N_23819,N_22181,N_22244);
xor U23820 (N_23820,N_22106,N_22655);
nand U23821 (N_23821,N_22069,N_22185);
or U23822 (N_23822,N_22608,N_22260);
or U23823 (N_23823,N_22081,N_22268);
nor U23824 (N_23824,N_22197,N_22055);
nor U23825 (N_23825,N_22385,N_22681);
or U23826 (N_23826,N_22129,N_22402);
nor U23827 (N_23827,N_22900,N_22504);
and U23828 (N_23828,N_22793,N_22958);
or U23829 (N_23829,N_22811,N_22137);
xnor U23830 (N_23830,N_22075,N_22710);
nand U23831 (N_23831,N_22248,N_22193);
nor U23832 (N_23832,N_22409,N_22884);
or U23833 (N_23833,N_22696,N_22757);
or U23834 (N_23834,N_22144,N_22466);
nand U23835 (N_23835,N_22609,N_22632);
nor U23836 (N_23836,N_22397,N_22953);
nor U23837 (N_23837,N_22060,N_22367);
nor U23838 (N_23838,N_22334,N_22881);
and U23839 (N_23839,N_22694,N_22056);
or U23840 (N_23840,N_22760,N_22481);
nand U23841 (N_23841,N_22739,N_22564);
and U23842 (N_23842,N_22442,N_22891);
and U23843 (N_23843,N_22167,N_22259);
xor U23844 (N_23844,N_22668,N_22771);
or U23845 (N_23845,N_22248,N_22917);
nor U23846 (N_23846,N_22802,N_22649);
nand U23847 (N_23847,N_22705,N_22474);
or U23848 (N_23848,N_22002,N_22016);
xnor U23849 (N_23849,N_22482,N_22693);
nand U23850 (N_23850,N_22989,N_22075);
xor U23851 (N_23851,N_22513,N_22745);
xor U23852 (N_23852,N_22675,N_22420);
xnor U23853 (N_23853,N_22285,N_22469);
and U23854 (N_23854,N_22387,N_22783);
or U23855 (N_23855,N_22792,N_22893);
or U23856 (N_23856,N_22115,N_22411);
or U23857 (N_23857,N_22413,N_22895);
or U23858 (N_23858,N_22431,N_22780);
nand U23859 (N_23859,N_22097,N_22410);
nand U23860 (N_23860,N_22049,N_22526);
and U23861 (N_23861,N_22359,N_22820);
xnor U23862 (N_23862,N_22242,N_22249);
nor U23863 (N_23863,N_22927,N_22067);
or U23864 (N_23864,N_22939,N_22866);
and U23865 (N_23865,N_22804,N_22944);
xnor U23866 (N_23866,N_22101,N_22451);
and U23867 (N_23867,N_22921,N_22062);
and U23868 (N_23868,N_22540,N_22247);
and U23869 (N_23869,N_22817,N_22710);
or U23870 (N_23870,N_22359,N_22637);
nor U23871 (N_23871,N_22689,N_22766);
nand U23872 (N_23872,N_22833,N_22426);
nor U23873 (N_23873,N_22261,N_22654);
nor U23874 (N_23874,N_22797,N_22602);
nand U23875 (N_23875,N_22751,N_22189);
and U23876 (N_23876,N_22767,N_22902);
nor U23877 (N_23877,N_22892,N_22058);
or U23878 (N_23878,N_22230,N_22067);
nor U23879 (N_23879,N_22360,N_22704);
nor U23880 (N_23880,N_22170,N_22423);
and U23881 (N_23881,N_22046,N_22233);
xor U23882 (N_23882,N_22621,N_22999);
nand U23883 (N_23883,N_22339,N_22940);
xor U23884 (N_23884,N_22317,N_22217);
or U23885 (N_23885,N_22568,N_22779);
or U23886 (N_23886,N_22866,N_22031);
and U23887 (N_23887,N_22041,N_22517);
nand U23888 (N_23888,N_22131,N_22279);
and U23889 (N_23889,N_22711,N_22232);
or U23890 (N_23890,N_22051,N_22664);
nand U23891 (N_23891,N_22690,N_22439);
nand U23892 (N_23892,N_22634,N_22471);
or U23893 (N_23893,N_22745,N_22684);
nor U23894 (N_23894,N_22156,N_22412);
nand U23895 (N_23895,N_22818,N_22746);
and U23896 (N_23896,N_22297,N_22690);
or U23897 (N_23897,N_22917,N_22573);
nor U23898 (N_23898,N_22553,N_22685);
xor U23899 (N_23899,N_22458,N_22574);
and U23900 (N_23900,N_22188,N_22612);
nor U23901 (N_23901,N_22697,N_22639);
xnor U23902 (N_23902,N_22108,N_22467);
nor U23903 (N_23903,N_22046,N_22366);
or U23904 (N_23904,N_22083,N_22813);
nand U23905 (N_23905,N_22039,N_22512);
xnor U23906 (N_23906,N_22438,N_22706);
xnor U23907 (N_23907,N_22829,N_22124);
nand U23908 (N_23908,N_22256,N_22075);
and U23909 (N_23909,N_22278,N_22660);
xor U23910 (N_23910,N_22655,N_22947);
nor U23911 (N_23911,N_22471,N_22259);
and U23912 (N_23912,N_22049,N_22870);
or U23913 (N_23913,N_22010,N_22669);
nor U23914 (N_23914,N_22601,N_22745);
or U23915 (N_23915,N_22270,N_22345);
xor U23916 (N_23916,N_22196,N_22674);
nand U23917 (N_23917,N_22472,N_22781);
and U23918 (N_23918,N_22411,N_22099);
nand U23919 (N_23919,N_22800,N_22264);
or U23920 (N_23920,N_22889,N_22739);
and U23921 (N_23921,N_22070,N_22147);
xor U23922 (N_23922,N_22668,N_22988);
xnor U23923 (N_23923,N_22935,N_22363);
nand U23924 (N_23924,N_22456,N_22444);
and U23925 (N_23925,N_22984,N_22766);
nor U23926 (N_23926,N_22996,N_22836);
xnor U23927 (N_23927,N_22821,N_22789);
or U23928 (N_23928,N_22969,N_22869);
nor U23929 (N_23929,N_22736,N_22462);
or U23930 (N_23930,N_22064,N_22657);
or U23931 (N_23931,N_22042,N_22990);
and U23932 (N_23932,N_22660,N_22756);
nor U23933 (N_23933,N_22935,N_22388);
nand U23934 (N_23934,N_22969,N_22110);
nor U23935 (N_23935,N_22669,N_22223);
nand U23936 (N_23936,N_22745,N_22699);
and U23937 (N_23937,N_22265,N_22636);
and U23938 (N_23938,N_22334,N_22944);
nor U23939 (N_23939,N_22393,N_22618);
nand U23940 (N_23940,N_22526,N_22275);
xnor U23941 (N_23941,N_22364,N_22475);
xnor U23942 (N_23942,N_22910,N_22174);
and U23943 (N_23943,N_22498,N_22483);
nand U23944 (N_23944,N_22388,N_22546);
nor U23945 (N_23945,N_22361,N_22935);
nor U23946 (N_23946,N_22403,N_22078);
nor U23947 (N_23947,N_22205,N_22089);
nand U23948 (N_23948,N_22873,N_22670);
and U23949 (N_23949,N_22575,N_22305);
nor U23950 (N_23950,N_22570,N_22192);
nand U23951 (N_23951,N_22746,N_22416);
or U23952 (N_23952,N_22839,N_22720);
xnor U23953 (N_23953,N_22038,N_22792);
nand U23954 (N_23954,N_22719,N_22044);
nor U23955 (N_23955,N_22343,N_22914);
nand U23956 (N_23956,N_22391,N_22803);
xor U23957 (N_23957,N_22584,N_22966);
and U23958 (N_23958,N_22373,N_22823);
nand U23959 (N_23959,N_22059,N_22322);
xor U23960 (N_23960,N_22327,N_22790);
nor U23961 (N_23961,N_22983,N_22114);
and U23962 (N_23962,N_22144,N_22980);
nand U23963 (N_23963,N_22591,N_22500);
and U23964 (N_23964,N_22738,N_22552);
or U23965 (N_23965,N_22716,N_22032);
xnor U23966 (N_23966,N_22096,N_22034);
and U23967 (N_23967,N_22782,N_22083);
nand U23968 (N_23968,N_22875,N_22171);
xor U23969 (N_23969,N_22667,N_22044);
nor U23970 (N_23970,N_22448,N_22136);
xor U23971 (N_23971,N_22208,N_22818);
and U23972 (N_23972,N_22369,N_22066);
nand U23973 (N_23973,N_22264,N_22176);
nand U23974 (N_23974,N_22244,N_22874);
or U23975 (N_23975,N_22019,N_22931);
nor U23976 (N_23976,N_22401,N_22338);
nand U23977 (N_23977,N_22990,N_22195);
and U23978 (N_23978,N_22958,N_22651);
nand U23979 (N_23979,N_22562,N_22957);
xor U23980 (N_23980,N_22876,N_22625);
xnor U23981 (N_23981,N_22434,N_22881);
and U23982 (N_23982,N_22266,N_22351);
and U23983 (N_23983,N_22916,N_22761);
and U23984 (N_23984,N_22458,N_22686);
or U23985 (N_23985,N_22747,N_22011);
nor U23986 (N_23986,N_22497,N_22959);
or U23987 (N_23987,N_22563,N_22629);
nand U23988 (N_23988,N_22404,N_22019);
nor U23989 (N_23989,N_22510,N_22849);
or U23990 (N_23990,N_22316,N_22966);
nor U23991 (N_23991,N_22835,N_22171);
xnor U23992 (N_23992,N_22222,N_22822);
and U23993 (N_23993,N_22043,N_22908);
nor U23994 (N_23994,N_22578,N_22717);
nor U23995 (N_23995,N_22755,N_22230);
or U23996 (N_23996,N_22138,N_22885);
nor U23997 (N_23997,N_22550,N_22300);
xnor U23998 (N_23998,N_22923,N_22493);
xnor U23999 (N_23999,N_22952,N_22659);
and U24000 (N_24000,N_23138,N_23219);
nor U24001 (N_24001,N_23664,N_23245);
nor U24002 (N_24002,N_23801,N_23575);
nand U24003 (N_24003,N_23679,N_23904);
and U24004 (N_24004,N_23702,N_23080);
xor U24005 (N_24005,N_23683,N_23215);
and U24006 (N_24006,N_23480,N_23186);
nor U24007 (N_24007,N_23891,N_23564);
xnor U24008 (N_24008,N_23563,N_23546);
nor U24009 (N_24009,N_23284,N_23743);
xnor U24010 (N_24010,N_23662,N_23759);
nor U24011 (N_24011,N_23440,N_23741);
nor U24012 (N_24012,N_23039,N_23503);
xnor U24013 (N_24013,N_23557,N_23568);
or U24014 (N_24014,N_23740,N_23250);
and U24015 (N_24015,N_23578,N_23548);
xor U24016 (N_24016,N_23691,N_23017);
xnor U24017 (N_24017,N_23948,N_23920);
nand U24018 (N_24018,N_23968,N_23814);
and U24019 (N_24019,N_23765,N_23853);
or U24020 (N_24020,N_23828,N_23234);
or U24021 (N_24021,N_23705,N_23323);
xnor U24022 (N_24022,N_23133,N_23012);
or U24023 (N_24023,N_23704,N_23657);
nand U24024 (N_24024,N_23602,N_23656);
and U24025 (N_24025,N_23352,N_23504);
nand U24026 (N_24026,N_23509,N_23607);
xor U24027 (N_24027,N_23579,N_23388);
nand U24028 (N_24028,N_23744,N_23241);
nor U24029 (N_24029,N_23748,N_23682);
nor U24030 (N_24030,N_23979,N_23906);
xor U24031 (N_24031,N_23175,N_23959);
xnor U24032 (N_24032,N_23417,N_23180);
xor U24033 (N_24033,N_23093,N_23128);
xor U24034 (N_24034,N_23430,N_23488);
nand U24035 (N_24035,N_23451,N_23608);
and U24036 (N_24036,N_23701,N_23519);
and U24037 (N_24037,N_23994,N_23925);
nor U24038 (N_24038,N_23350,N_23767);
nand U24039 (N_24039,N_23224,N_23206);
nand U24040 (N_24040,N_23811,N_23552);
or U24041 (N_24041,N_23275,N_23877);
and U24042 (N_24042,N_23130,N_23021);
nand U24043 (N_24043,N_23867,N_23263);
or U24044 (N_24044,N_23949,N_23745);
and U24045 (N_24045,N_23884,N_23062);
xor U24046 (N_24046,N_23232,N_23373);
nor U24047 (N_24047,N_23048,N_23567);
xnor U24048 (N_24048,N_23084,N_23518);
xnor U24049 (N_24049,N_23190,N_23908);
nand U24050 (N_24050,N_23760,N_23221);
nor U24051 (N_24051,N_23537,N_23136);
or U24052 (N_24052,N_23145,N_23897);
nand U24053 (N_24053,N_23095,N_23817);
nor U24054 (N_24054,N_23609,N_23363);
and U24055 (N_24055,N_23663,N_23225);
xor U24056 (N_24056,N_23650,N_23617);
xnor U24057 (N_24057,N_23902,N_23002);
nor U24058 (N_24058,N_23590,N_23634);
nor U24059 (N_24059,N_23766,N_23613);
and U24060 (N_24060,N_23629,N_23622);
or U24061 (N_24061,N_23696,N_23140);
nor U24062 (N_24062,N_23846,N_23969);
nor U24063 (N_24063,N_23070,N_23202);
and U24064 (N_24064,N_23954,N_23854);
and U24065 (N_24065,N_23318,N_23468);
xnor U24066 (N_24066,N_23097,N_23424);
nand U24067 (N_24067,N_23860,N_23573);
xor U24068 (N_24068,N_23534,N_23732);
or U24069 (N_24069,N_23758,N_23840);
xnor U24070 (N_24070,N_23924,N_23781);
or U24071 (N_24071,N_23049,N_23463);
and U24072 (N_24072,N_23928,N_23916);
xnor U24073 (N_24073,N_23266,N_23269);
nor U24074 (N_24074,N_23614,N_23479);
nor U24075 (N_24075,N_23319,N_23396);
xor U24076 (N_24076,N_23460,N_23076);
xor U24077 (N_24077,N_23303,N_23692);
and U24078 (N_24078,N_23471,N_23653);
and U24079 (N_24079,N_23217,N_23777);
nand U24080 (N_24080,N_23796,N_23977);
xor U24081 (N_24081,N_23357,N_23187);
xor U24082 (N_24082,N_23718,N_23652);
xor U24083 (N_24083,N_23423,N_23061);
and U24084 (N_24084,N_23272,N_23978);
nor U24085 (N_24085,N_23866,N_23072);
nor U24086 (N_24086,N_23645,N_23207);
nor U24087 (N_24087,N_23171,N_23922);
nor U24088 (N_24088,N_23859,N_23820);
or U24089 (N_24089,N_23943,N_23379);
or U24090 (N_24090,N_23527,N_23085);
nor U24091 (N_24091,N_23163,N_23415);
nor U24092 (N_24092,N_23485,N_23688);
nand U24093 (N_24093,N_23746,N_23950);
xor U24094 (N_24094,N_23115,N_23574);
nor U24095 (N_24095,N_23299,N_23341);
or U24096 (N_24096,N_23235,N_23627);
nor U24097 (N_24097,N_23214,N_23999);
or U24098 (N_24098,N_23389,N_23862);
or U24099 (N_24099,N_23001,N_23756);
nand U24100 (N_24100,N_23466,N_23886);
or U24101 (N_24101,N_23510,N_23813);
and U24102 (N_24102,N_23330,N_23201);
nor U24103 (N_24103,N_23459,N_23022);
and U24104 (N_24104,N_23780,N_23894);
xnor U24105 (N_24105,N_23386,N_23099);
xor U24106 (N_24106,N_23774,N_23166);
nor U24107 (N_24107,N_23285,N_23462);
or U24108 (N_24108,N_23831,N_23015);
nand U24109 (N_24109,N_23031,N_23581);
nor U24110 (N_24110,N_23324,N_23342);
and U24111 (N_24111,N_23339,N_23051);
nor U24112 (N_24112,N_23254,N_23251);
or U24113 (N_24113,N_23678,N_23794);
and U24114 (N_24114,N_23942,N_23901);
or U24115 (N_24115,N_23110,N_23249);
and U24116 (N_24116,N_23298,N_23848);
nand U24117 (N_24117,N_23461,N_23077);
nor U24118 (N_24118,N_23496,N_23806);
nor U24119 (N_24119,N_23108,N_23422);
or U24120 (N_24120,N_23804,N_23727);
or U24121 (N_24121,N_23346,N_23103);
nand U24122 (N_24122,N_23872,N_23812);
nor U24123 (N_24123,N_23952,N_23029);
xnor U24124 (N_24124,N_23577,N_23000);
or U24125 (N_24125,N_23554,N_23047);
nor U24126 (N_24126,N_23403,N_23020);
and U24127 (N_24127,N_23671,N_23040);
nor U24128 (N_24128,N_23591,N_23535);
or U24129 (N_24129,N_23231,N_23680);
nand U24130 (N_24130,N_23927,N_23615);
and U24131 (N_24131,N_23402,N_23880);
nand U24132 (N_24132,N_23238,N_23864);
xor U24133 (N_24133,N_23540,N_23827);
nor U24134 (N_24134,N_23934,N_23932);
and U24135 (N_24135,N_23371,N_23304);
and U24136 (N_24136,N_23027,N_23405);
and U24137 (N_24137,N_23420,N_23165);
nor U24138 (N_24138,N_23797,N_23320);
and U24139 (N_24139,N_23962,N_23625);
or U24140 (N_24140,N_23809,N_23054);
xnor U24141 (N_24141,N_23729,N_23909);
nand U24142 (N_24142,N_23689,N_23270);
nand U24143 (N_24143,N_23871,N_23967);
or U24144 (N_24144,N_23648,N_23869);
and U24145 (N_24145,N_23915,N_23690);
nand U24146 (N_24146,N_23944,N_23694);
or U24147 (N_24147,N_23294,N_23153);
or U24148 (N_24148,N_23695,N_23161);
and U24149 (N_24149,N_23003,N_23951);
xor U24150 (N_24150,N_23899,N_23127);
nor U24151 (N_24151,N_23257,N_23368);
nand U24152 (N_24152,N_23068,N_23287);
nand U24153 (N_24153,N_23725,N_23052);
or U24154 (N_24154,N_23595,N_23588);
nor U24155 (N_24155,N_23268,N_23053);
or U24156 (N_24156,N_23734,N_23632);
or U24157 (N_24157,N_23078,N_23787);
nor U24158 (N_24158,N_23436,N_23309);
and U24159 (N_24159,N_23026,N_23086);
or U24160 (N_24160,N_23511,N_23390);
xor U24161 (N_24161,N_23983,N_23283);
and U24162 (N_24162,N_23401,N_23385);
or U24163 (N_24163,N_23965,N_23300);
and U24164 (N_24164,N_23685,N_23911);
and U24165 (N_24165,N_23432,N_23660);
nor U24166 (N_24166,N_23322,N_23314);
nand U24167 (N_24167,N_23895,N_23446);
or U24168 (N_24168,N_23148,N_23450);
nand U24169 (N_24169,N_23870,N_23146);
xnor U24170 (N_24170,N_23857,N_23096);
nor U24171 (N_24171,N_23142,N_23297);
xnor U24172 (N_24172,N_23639,N_23223);
nand U24173 (N_24173,N_23400,N_23089);
nor U24174 (N_24174,N_23984,N_23628);
xnor U24175 (N_24175,N_23155,N_23264);
nor U24176 (N_24176,N_23467,N_23365);
nor U24177 (N_24177,N_23056,N_23456);
nor U24178 (N_24178,N_23836,N_23106);
nand U24179 (N_24179,N_23789,N_23776);
nand U24180 (N_24180,N_23624,N_23307);
or U24181 (N_24181,N_23976,N_23454);
and U24182 (N_24182,N_23913,N_23315);
and U24183 (N_24183,N_23798,N_23094);
and U24184 (N_24184,N_23344,N_23733);
or U24185 (N_24185,N_23542,N_23404);
nor U24186 (N_24186,N_23075,N_23289);
nor U24187 (N_24187,N_23550,N_23633);
nor U24188 (N_24188,N_23649,N_23749);
nand U24189 (N_24189,N_23807,N_23670);
xor U24190 (N_24190,N_23113,N_23247);
xor U24191 (N_24191,N_23757,N_23448);
xnor U24192 (N_24192,N_23525,N_23541);
nand U24193 (N_24193,N_23229,N_23659);
or U24194 (N_24194,N_23929,N_23167);
or U24195 (N_24195,N_23008,N_23675);
nand U24196 (N_24196,N_23367,N_23998);
or U24197 (N_24197,N_23406,N_23487);
nand U24198 (N_24198,N_23100,N_23018);
nor U24199 (N_24199,N_23782,N_23159);
or U24200 (N_24200,N_23035,N_23770);
xnor U24201 (N_24201,N_23865,N_23712);
and U24202 (N_24202,N_23343,N_23412);
nor U24203 (N_24203,N_23521,N_23042);
and U24204 (N_24204,N_23612,N_23316);
or U24205 (N_24205,N_23286,N_23174);
xnor U24206 (N_24206,N_23011,N_23987);
nand U24207 (N_24207,N_23843,N_23391);
or U24208 (N_24208,N_23839,N_23885);
and U24209 (N_24209,N_23879,N_23311);
nor U24210 (N_24210,N_23618,N_23707);
nor U24211 (N_24211,N_23980,N_23939);
and U24212 (N_24212,N_23930,N_23296);
nor U24213 (N_24213,N_23730,N_23667);
and U24214 (N_24214,N_23105,N_23646);
nor U24215 (N_24215,N_23007,N_23710);
nand U24216 (N_24216,N_23255,N_23935);
or U24217 (N_24217,N_23005,N_23507);
nand U24218 (N_24218,N_23045,N_23668);
and U24219 (N_24219,N_23055,N_23555);
xor U24220 (N_24220,N_23384,N_23855);
nor U24221 (N_24221,N_23416,N_23244);
xnor U24222 (N_24222,N_23262,N_23370);
nand U24223 (N_24223,N_23355,N_23754);
or U24224 (N_24224,N_23562,N_23775);
and U24225 (N_24225,N_23476,N_23261);
and U24226 (N_24226,N_23973,N_23566);
and U24227 (N_24227,N_23763,N_23558);
nand U24228 (N_24228,N_23141,N_23783);
and U24229 (N_24229,N_23892,N_23842);
and U24230 (N_24230,N_23687,N_23785);
nand U24231 (N_24231,N_23861,N_23449);
nor U24232 (N_24232,N_23570,N_23116);
xor U24233 (N_24233,N_23119,N_23966);
nand U24234 (N_24234,N_23889,N_23800);
nand U24235 (N_24235,N_23313,N_23635);
or U24236 (N_24236,N_23046,N_23372);
nor U24237 (N_24237,N_23220,N_23387);
nor U24238 (N_24238,N_23458,N_23610);
and U24239 (N_24239,N_23538,N_23997);
nand U24240 (N_24240,N_23936,N_23677);
nand U24241 (N_24241,N_23144,N_23524);
or U24242 (N_24242,N_23457,N_23178);
xor U24243 (N_24243,N_23536,N_23023);
and U24244 (N_24244,N_23723,N_23673);
or U24245 (N_24245,N_23258,N_23443);
nor U24246 (N_24246,N_23874,N_23724);
nor U24247 (N_24247,N_23583,N_23619);
nand U24248 (N_24248,N_23267,N_23064);
nand U24249 (N_24249,N_23835,N_23398);
and U24250 (N_24250,N_23523,N_23762);
nor U24251 (N_24251,N_23325,N_23706);
nor U24252 (N_24252,N_23397,N_23547);
nand U24253 (N_24253,N_23408,N_23970);
or U24254 (N_24254,N_23698,N_23009);
or U24255 (N_24255,N_23502,N_23394);
and U24256 (N_24256,N_23837,N_23681);
xnor U24257 (N_24257,N_23111,N_23700);
nand U24258 (N_24258,N_23465,N_23883);
and U24259 (N_24259,N_23213,N_23572);
nand U24260 (N_24260,N_23152,N_23469);
or U24261 (N_24261,N_23829,N_23844);
nand U24262 (N_24262,N_23981,N_23990);
nor U24263 (N_24263,N_23516,N_23963);
nor U24264 (N_24264,N_23553,N_23338);
nand U24265 (N_24265,N_23728,N_23816);
xnor U24266 (N_24266,N_23358,N_23335);
nand U24267 (N_24267,N_23222,N_23114);
xnor U24268 (N_24268,N_23382,N_23074);
nor U24269 (N_24269,N_23209,N_23079);
nand U24270 (N_24270,N_23090,N_23198);
nand U24271 (N_24271,N_23526,N_23147);
or U24272 (N_24272,N_23317,N_23065);
or U24273 (N_24273,N_23362,N_23279);
or U24274 (N_24274,N_23135,N_23060);
nand U24275 (N_24275,N_23717,N_23273);
nor U24276 (N_24276,N_23203,N_23772);
or U24277 (N_24277,N_23123,N_23810);
nand U24278 (N_24278,N_23571,N_23508);
nand U24279 (N_24279,N_23193,N_23742);
xor U24280 (N_24280,N_23421,N_23228);
xnor U24281 (N_24281,N_23109,N_23520);
or U24282 (N_24282,N_23237,N_23900);
or U24283 (N_24283,N_23600,N_23960);
xnor U24284 (N_24284,N_23822,N_23082);
nand U24285 (N_24285,N_23442,N_23996);
nand U24286 (N_24286,N_23019,N_23851);
and U24287 (N_24287,N_23938,N_23071);
and U24288 (N_24288,N_23910,N_23713);
or U24289 (N_24289,N_23993,N_23280);
or U24290 (N_24290,N_23143,N_23971);
nand U24291 (N_24291,N_23102,N_23189);
or U24292 (N_24292,N_23905,N_23149);
xor U24293 (N_24293,N_23066,N_23834);
nor U24294 (N_24294,N_23150,N_23196);
or U24295 (N_24295,N_23771,N_23183);
or U24296 (N_24296,N_23033,N_23374);
nand U24297 (N_24297,N_23711,N_23778);
nor U24298 (N_24298,N_23098,N_23043);
and U24299 (N_24299,N_23821,N_23332);
nand U24300 (N_24300,N_23719,N_23531);
or U24301 (N_24301,N_23972,N_23192);
xnor U24302 (N_24302,N_23088,N_23751);
or U24303 (N_24303,N_23277,N_23293);
nor U24304 (N_24304,N_23212,N_23755);
nand U24305 (N_24305,N_23032,N_23118);
xor U24306 (N_24306,N_23559,N_23252);
nor U24307 (N_24307,N_23014,N_23992);
or U24308 (N_24308,N_23549,N_23647);
or U24309 (N_24309,N_23592,N_23483);
and U24310 (N_24310,N_23274,N_23931);
nand U24311 (N_24311,N_23326,N_23940);
nor U24312 (N_24312,N_23517,N_23383);
or U24313 (N_24313,N_23515,N_23427);
and U24314 (N_24314,N_23359,N_23425);
nor U24315 (N_24315,N_23117,N_23565);
nand U24316 (N_24316,N_23982,N_23151);
nand U24317 (N_24317,N_23893,N_23561);
nor U24318 (N_24318,N_23124,N_23411);
and U24319 (N_24319,N_23773,N_23271);
nor U24320 (N_24320,N_23482,N_23708);
or U24321 (N_24321,N_23455,N_23529);
or U24322 (N_24322,N_23907,N_23500);
xnor U24323 (N_24323,N_23069,N_23447);
and U24324 (N_24324,N_23958,N_23532);
xnor U24325 (N_24325,N_23666,N_23464);
nand U24326 (N_24326,N_23351,N_23321);
xor U24327 (N_24327,N_23988,N_23709);
nand U24328 (N_24328,N_23059,N_23890);
nand U24329 (N_24329,N_23941,N_23158);
xor U24330 (N_24330,N_23896,N_23506);
and U24331 (N_24331,N_23216,N_23197);
xnor U24332 (N_24332,N_23490,N_23306);
nand U24333 (N_24333,N_23703,N_23256);
and U24334 (N_24334,N_23495,N_23038);
xnor U24335 (N_24335,N_23331,N_23686);
or U24336 (N_24336,N_23218,N_23620);
or U24337 (N_24337,N_23030,N_23587);
or U24338 (N_24338,N_23499,N_23194);
and U24339 (N_24339,N_23131,N_23605);
nand U24340 (N_24340,N_23651,N_23439);
nand U24341 (N_24341,N_23208,N_23641);
xnor U24342 (N_24342,N_23819,N_23137);
nand U24343 (N_24343,N_23584,N_23528);
or U24344 (N_24344,N_23361,N_23750);
nand U24345 (N_24345,N_23621,N_23434);
and U24346 (N_24346,N_23986,N_23768);
nand U24347 (N_24347,N_23716,N_23539);
or U24348 (N_24348,N_23302,N_23409);
nand U24349 (N_24349,N_23168,N_23779);
xor U24350 (N_24350,N_23291,N_23199);
and U24351 (N_24351,N_23429,N_23661);
nor U24352 (N_24352,N_23946,N_23057);
xor U24353 (N_24353,N_23024,N_23281);
xnor U24354 (N_24354,N_23926,N_23337);
xor U24355 (N_24355,N_23191,N_23636);
xor U24356 (N_24356,N_23125,N_23841);
nand U24357 (N_24357,N_23964,N_23881);
nand U24358 (N_24358,N_23081,N_23852);
xor U24359 (N_24359,N_23543,N_23722);
and U24360 (N_24360,N_23898,N_23050);
and U24361 (N_24361,N_23699,N_23808);
or U24362 (N_24362,N_23156,N_23989);
nor U24363 (N_24363,N_23594,N_23248);
nor U24364 (N_24364,N_23107,N_23580);
or U24365 (N_24365,N_23340,N_23377);
and U24366 (N_24366,N_23016,N_23672);
nor U24367 (N_24367,N_23334,N_23917);
nand U24368 (N_24368,N_23603,N_23230);
nor U24369 (N_24369,N_23172,N_23582);
nor U24370 (N_24370,N_23784,N_23470);
nand U24371 (N_24371,N_23576,N_23721);
xor U24372 (N_24372,N_23551,N_23112);
nor U24373 (N_24373,N_23288,N_23164);
and U24374 (N_24374,N_23444,N_23010);
and U24375 (N_24375,N_23497,N_23157);
xnor U24376 (N_24376,N_23182,N_23364);
and U24377 (N_24377,N_23642,N_23282);
or U24378 (N_24378,N_23513,N_23715);
or U24379 (N_24379,N_23239,N_23995);
nand U24380 (N_24380,N_23393,N_23025);
xnor U24381 (N_24381,N_23903,N_23735);
or U24382 (N_24382,N_23947,N_23638);
nor U24383 (N_24383,N_23292,N_23975);
and U24384 (N_24384,N_23037,N_23747);
nor U24385 (N_24385,N_23791,N_23833);
or U24386 (N_24386,N_23586,N_23345);
or U24387 (N_24387,N_23176,N_23790);
and U24388 (N_24388,N_23290,N_23850);
nor U24389 (N_24389,N_23188,N_23753);
nor U24390 (N_24390,N_23593,N_23626);
xnor U24391 (N_24391,N_23585,N_23769);
xnor U24392 (N_24392,N_23227,N_23825);
xnor U24393 (N_24393,N_23631,N_23505);
nor U24394 (N_24394,N_23083,N_23604);
nand U24395 (N_24395,N_23623,N_23184);
or U24396 (N_24396,N_23985,N_23328);
xnor U24397 (N_24397,N_23013,N_23478);
xnor U24398 (N_24398,N_23265,N_23132);
and U24399 (N_24399,N_23956,N_23381);
and U24400 (N_24400,N_23498,N_23376);
or U24401 (N_24401,N_23676,N_23738);
xor U24402 (N_24402,N_23752,N_23139);
xor U24403 (N_24403,N_23134,N_23826);
xor U24404 (N_24404,N_23173,N_23243);
or U24405 (N_24405,N_23177,N_23353);
nand U24406 (N_24406,N_23640,N_23418);
and U24407 (N_24407,N_23034,N_23426);
nor U24408 (N_24408,N_23560,N_23305);
or U24409 (N_24409,N_23492,N_23354);
xor U24410 (N_24410,N_23347,N_23569);
nand U24411 (N_24411,N_23803,N_23475);
nand U24412 (N_24412,N_23545,N_23611);
nand U24413 (N_24413,N_23530,N_23210);
or U24414 (N_24414,N_23438,N_23974);
nor U24415 (N_24415,N_23616,N_23799);
nand U24416 (N_24416,N_23805,N_23832);
and U24417 (N_24417,N_23445,N_23493);
or U24418 (N_24418,N_23697,N_23204);
or U24419 (N_24419,N_23731,N_23858);
and U24420 (N_24420,N_23349,N_23477);
xnor U24421 (N_24421,N_23308,N_23606);
xor U24422 (N_24422,N_23036,N_23253);
and U24423 (N_24423,N_23126,N_23120);
or U24424 (N_24424,N_23399,N_23882);
and U24425 (N_24425,N_23643,N_23875);
and U24426 (N_24426,N_23484,N_23669);
nand U24427 (N_24427,N_23453,N_23195);
and U24428 (N_24428,N_23788,N_23792);
or U24429 (N_24429,N_23336,N_23955);
nand U24430 (N_24430,N_23665,N_23856);
and U24431 (N_24431,N_23838,N_23878);
and U24432 (N_24432,N_23491,N_23044);
and U24433 (N_24433,N_23556,N_23953);
or U24434 (N_24434,N_23474,N_23067);
nor U24435 (N_24435,N_23849,N_23333);
nand U24436 (N_24436,N_23658,N_23181);
nor U24437 (N_24437,N_23830,N_23823);
nand U24438 (N_24438,N_23887,N_23433);
and U24439 (N_24439,N_23414,N_23654);
nor U24440 (N_24440,N_23795,N_23514);
and U24441 (N_24441,N_23121,N_23957);
and U24442 (N_24442,N_23589,N_23876);
nor U24443 (N_24443,N_23522,N_23092);
nor U24444 (N_24444,N_23378,N_23041);
and U24445 (N_24445,N_23533,N_23598);
and U24446 (N_24446,N_23726,N_23937);
xor U24447 (N_24447,N_23129,N_23091);
nand U24448 (N_24448,N_23063,N_23233);
and U24449 (N_24449,N_23240,N_23260);
or U24450 (N_24450,N_23205,N_23162);
nand U24451 (N_24451,N_23441,N_23737);
nor U24452 (N_24452,N_23597,N_23918);
xnor U24453 (N_24453,N_23786,N_23369);
or U24454 (N_24454,N_23793,N_23278);
or U24455 (N_24455,N_23185,N_23888);
nor U24456 (N_24456,N_23226,N_23912);
nor U24457 (N_24457,N_23923,N_23246);
xor U24458 (N_24458,N_23329,N_23637);
and U24459 (N_24459,N_23655,N_23544);
xnor U24460 (N_24460,N_23473,N_23961);
nor U24461 (N_24461,N_23242,N_23170);
or U24462 (N_24462,N_23481,N_23366);
and U24463 (N_24463,N_23058,N_23863);
nor U24464 (N_24464,N_23847,N_23601);
and U24465 (N_24465,N_23360,N_23684);
nor U24466 (N_24466,N_23348,N_23375);
or U24467 (N_24467,N_23945,N_23452);
and U24468 (N_24468,N_23407,N_23736);
or U24469 (N_24469,N_23489,N_23073);
and U24470 (N_24470,N_23824,N_23104);
and U24471 (N_24471,N_23310,N_23428);
xnor U24472 (N_24472,N_23087,N_23739);
nand U24473 (N_24473,N_23714,N_23921);
xor U24474 (N_24474,N_23380,N_23818);
or U24475 (N_24475,N_23200,N_23327);
and U24476 (N_24476,N_23435,N_23764);
nor U24477 (N_24477,N_23501,N_23720);
and U24478 (N_24478,N_23596,N_23160);
and U24479 (N_24479,N_23410,N_23295);
nor U24480 (N_24480,N_23512,N_23914);
or U24481 (N_24481,N_23919,N_23644);
nor U24482 (N_24482,N_23494,N_23154);
xnor U24483 (N_24483,N_23276,N_23169);
xnor U24484 (N_24484,N_23395,N_23437);
xor U24485 (N_24485,N_23122,N_23599);
nor U24486 (N_24486,N_23259,N_23211);
nor U24487 (N_24487,N_23802,N_23356);
nor U24488 (N_24488,N_23004,N_23236);
or U24489 (N_24489,N_23419,N_23761);
xor U24490 (N_24490,N_23312,N_23028);
nor U24491 (N_24491,N_23472,N_23991);
xnor U24492 (N_24492,N_23486,N_23693);
and U24493 (N_24493,N_23674,N_23101);
nor U24494 (N_24494,N_23431,N_23845);
xnor U24495 (N_24495,N_23392,N_23815);
nor U24496 (N_24496,N_23873,N_23868);
nand U24497 (N_24497,N_23006,N_23933);
xnor U24498 (N_24498,N_23413,N_23301);
nor U24499 (N_24499,N_23179,N_23630);
and U24500 (N_24500,N_23866,N_23932);
nor U24501 (N_24501,N_23258,N_23698);
nand U24502 (N_24502,N_23371,N_23367);
nor U24503 (N_24503,N_23553,N_23877);
nand U24504 (N_24504,N_23950,N_23723);
and U24505 (N_24505,N_23429,N_23046);
or U24506 (N_24506,N_23072,N_23750);
nor U24507 (N_24507,N_23663,N_23425);
and U24508 (N_24508,N_23641,N_23838);
and U24509 (N_24509,N_23578,N_23066);
xnor U24510 (N_24510,N_23157,N_23578);
nor U24511 (N_24511,N_23679,N_23404);
nand U24512 (N_24512,N_23942,N_23882);
nand U24513 (N_24513,N_23607,N_23096);
xnor U24514 (N_24514,N_23054,N_23452);
nand U24515 (N_24515,N_23522,N_23608);
and U24516 (N_24516,N_23736,N_23181);
nor U24517 (N_24517,N_23104,N_23262);
and U24518 (N_24518,N_23235,N_23714);
nor U24519 (N_24519,N_23287,N_23437);
nand U24520 (N_24520,N_23678,N_23519);
nand U24521 (N_24521,N_23389,N_23484);
xnor U24522 (N_24522,N_23759,N_23612);
nand U24523 (N_24523,N_23408,N_23127);
and U24524 (N_24524,N_23873,N_23991);
and U24525 (N_24525,N_23108,N_23678);
nand U24526 (N_24526,N_23101,N_23891);
nor U24527 (N_24527,N_23087,N_23283);
xor U24528 (N_24528,N_23859,N_23197);
or U24529 (N_24529,N_23460,N_23896);
and U24530 (N_24530,N_23548,N_23458);
xor U24531 (N_24531,N_23587,N_23938);
and U24532 (N_24532,N_23407,N_23570);
or U24533 (N_24533,N_23567,N_23401);
and U24534 (N_24534,N_23436,N_23198);
and U24535 (N_24535,N_23585,N_23827);
nor U24536 (N_24536,N_23468,N_23713);
or U24537 (N_24537,N_23811,N_23681);
xnor U24538 (N_24538,N_23197,N_23337);
nand U24539 (N_24539,N_23664,N_23636);
or U24540 (N_24540,N_23710,N_23078);
xor U24541 (N_24541,N_23430,N_23320);
nand U24542 (N_24542,N_23625,N_23815);
nor U24543 (N_24543,N_23060,N_23764);
and U24544 (N_24544,N_23547,N_23707);
and U24545 (N_24545,N_23285,N_23486);
xnor U24546 (N_24546,N_23888,N_23824);
and U24547 (N_24547,N_23329,N_23222);
nor U24548 (N_24548,N_23537,N_23014);
and U24549 (N_24549,N_23274,N_23839);
xor U24550 (N_24550,N_23887,N_23502);
nand U24551 (N_24551,N_23560,N_23868);
or U24552 (N_24552,N_23476,N_23263);
nor U24553 (N_24553,N_23945,N_23349);
xor U24554 (N_24554,N_23925,N_23610);
and U24555 (N_24555,N_23993,N_23812);
nand U24556 (N_24556,N_23106,N_23549);
xor U24557 (N_24557,N_23883,N_23521);
xor U24558 (N_24558,N_23182,N_23708);
nor U24559 (N_24559,N_23418,N_23655);
and U24560 (N_24560,N_23675,N_23866);
and U24561 (N_24561,N_23164,N_23780);
xor U24562 (N_24562,N_23064,N_23537);
or U24563 (N_24563,N_23752,N_23393);
and U24564 (N_24564,N_23710,N_23063);
and U24565 (N_24565,N_23964,N_23551);
or U24566 (N_24566,N_23180,N_23701);
and U24567 (N_24567,N_23031,N_23530);
or U24568 (N_24568,N_23001,N_23123);
nor U24569 (N_24569,N_23817,N_23807);
or U24570 (N_24570,N_23647,N_23418);
and U24571 (N_24571,N_23550,N_23122);
nor U24572 (N_24572,N_23573,N_23477);
nand U24573 (N_24573,N_23983,N_23613);
and U24574 (N_24574,N_23360,N_23736);
or U24575 (N_24575,N_23481,N_23293);
and U24576 (N_24576,N_23129,N_23892);
nor U24577 (N_24577,N_23186,N_23563);
xor U24578 (N_24578,N_23555,N_23755);
or U24579 (N_24579,N_23314,N_23625);
and U24580 (N_24580,N_23982,N_23752);
nor U24581 (N_24581,N_23484,N_23214);
xor U24582 (N_24582,N_23636,N_23042);
or U24583 (N_24583,N_23436,N_23093);
nand U24584 (N_24584,N_23837,N_23096);
or U24585 (N_24585,N_23696,N_23011);
and U24586 (N_24586,N_23043,N_23897);
nand U24587 (N_24587,N_23117,N_23388);
or U24588 (N_24588,N_23157,N_23179);
nand U24589 (N_24589,N_23729,N_23100);
or U24590 (N_24590,N_23782,N_23501);
nor U24591 (N_24591,N_23133,N_23250);
nor U24592 (N_24592,N_23498,N_23779);
xnor U24593 (N_24593,N_23186,N_23879);
nor U24594 (N_24594,N_23376,N_23819);
nor U24595 (N_24595,N_23732,N_23609);
nor U24596 (N_24596,N_23115,N_23915);
xnor U24597 (N_24597,N_23841,N_23780);
or U24598 (N_24598,N_23521,N_23364);
nand U24599 (N_24599,N_23498,N_23226);
nand U24600 (N_24600,N_23018,N_23324);
or U24601 (N_24601,N_23662,N_23346);
or U24602 (N_24602,N_23642,N_23533);
nand U24603 (N_24603,N_23690,N_23792);
xnor U24604 (N_24604,N_23480,N_23355);
nand U24605 (N_24605,N_23932,N_23107);
nor U24606 (N_24606,N_23069,N_23628);
nor U24607 (N_24607,N_23069,N_23826);
or U24608 (N_24608,N_23334,N_23429);
xor U24609 (N_24609,N_23519,N_23603);
and U24610 (N_24610,N_23959,N_23295);
nand U24611 (N_24611,N_23593,N_23933);
nor U24612 (N_24612,N_23172,N_23585);
nand U24613 (N_24613,N_23251,N_23093);
and U24614 (N_24614,N_23879,N_23443);
or U24615 (N_24615,N_23529,N_23068);
nor U24616 (N_24616,N_23370,N_23324);
nor U24617 (N_24617,N_23656,N_23301);
nor U24618 (N_24618,N_23266,N_23657);
or U24619 (N_24619,N_23685,N_23984);
nand U24620 (N_24620,N_23571,N_23939);
nand U24621 (N_24621,N_23116,N_23244);
and U24622 (N_24622,N_23421,N_23894);
nor U24623 (N_24623,N_23028,N_23094);
nand U24624 (N_24624,N_23185,N_23076);
and U24625 (N_24625,N_23195,N_23029);
and U24626 (N_24626,N_23438,N_23456);
nand U24627 (N_24627,N_23141,N_23715);
nand U24628 (N_24628,N_23231,N_23948);
nand U24629 (N_24629,N_23837,N_23894);
or U24630 (N_24630,N_23670,N_23012);
or U24631 (N_24631,N_23274,N_23558);
nor U24632 (N_24632,N_23603,N_23430);
nor U24633 (N_24633,N_23703,N_23793);
xor U24634 (N_24634,N_23240,N_23707);
and U24635 (N_24635,N_23207,N_23132);
and U24636 (N_24636,N_23399,N_23603);
nand U24637 (N_24637,N_23046,N_23056);
xnor U24638 (N_24638,N_23717,N_23714);
nand U24639 (N_24639,N_23275,N_23871);
nor U24640 (N_24640,N_23359,N_23705);
and U24641 (N_24641,N_23812,N_23436);
nand U24642 (N_24642,N_23552,N_23805);
xor U24643 (N_24643,N_23193,N_23383);
xor U24644 (N_24644,N_23690,N_23248);
xor U24645 (N_24645,N_23174,N_23287);
or U24646 (N_24646,N_23029,N_23956);
or U24647 (N_24647,N_23335,N_23460);
nand U24648 (N_24648,N_23867,N_23532);
xor U24649 (N_24649,N_23730,N_23504);
xor U24650 (N_24650,N_23078,N_23654);
nor U24651 (N_24651,N_23319,N_23107);
or U24652 (N_24652,N_23524,N_23243);
and U24653 (N_24653,N_23013,N_23626);
xnor U24654 (N_24654,N_23743,N_23571);
nor U24655 (N_24655,N_23607,N_23540);
nor U24656 (N_24656,N_23783,N_23778);
or U24657 (N_24657,N_23718,N_23664);
or U24658 (N_24658,N_23782,N_23609);
or U24659 (N_24659,N_23184,N_23652);
nor U24660 (N_24660,N_23010,N_23575);
nand U24661 (N_24661,N_23731,N_23732);
and U24662 (N_24662,N_23133,N_23172);
and U24663 (N_24663,N_23570,N_23985);
and U24664 (N_24664,N_23566,N_23436);
nand U24665 (N_24665,N_23569,N_23467);
and U24666 (N_24666,N_23731,N_23805);
or U24667 (N_24667,N_23823,N_23467);
nor U24668 (N_24668,N_23487,N_23079);
nand U24669 (N_24669,N_23055,N_23457);
nor U24670 (N_24670,N_23161,N_23049);
nor U24671 (N_24671,N_23879,N_23106);
nand U24672 (N_24672,N_23042,N_23357);
nand U24673 (N_24673,N_23802,N_23108);
xnor U24674 (N_24674,N_23887,N_23593);
nand U24675 (N_24675,N_23556,N_23812);
nor U24676 (N_24676,N_23138,N_23786);
nand U24677 (N_24677,N_23983,N_23399);
nor U24678 (N_24678,N_23694,N_23616);
nand U24679 (N_24679,N_23512,N_23514);
xnor U24680 (N_24680,N_23015,N_23174);
or U24681 (N_24681,N_23993,N_23554);
xor U24682 (N_24682,N_23365,N_23664);
or U24683 (N_24683,N_23006,N_23376);
xor U24684 (N_24684,N_23114,N_23397);
nand U24685 (N_24685,N_23330,N_23750);
or U24686 (N_24686,N_23077,N_23165);
nor U24687 (N_24687,N_23099,N_23150);
nand U24688 (N_24688,N_23252,N_23620);
xnor U24689 (N_24689,N_23159,N_23335);
nand U24690 (N_24690,N_23891,N_23866);
xor U24691 (N_24691,N_23852,N_23222);
and U24692 (N_24692,N_23280,N_23697);
xnor U24693 (N_24693,N_23474,N_23261);
and U24694 (N_24694,N_23345,N_23599);
or U24695 (N_24695,N_23871,N_23844);
nor U24696 (N_24696,N_23149,N_23667);
or U24697 (N_24697,N_23370,N_23552);
nor U24698 (N_24698,N_23988,N_23320);
nand U24699 (N_24699,N_23103,N_23294);
nor U24700 (N_24700,N_23463,N_23259);
nor U24701 (N_24701,N_23435,N_23662);
nor U24702 (N_24702,N_23450,N_23535);
or U24703 (N_24703,N_23286,N_23265);
xnor U24704 (N_24704,N_23688,N_23350);
nor U24705 (N_24705,N_23692,N_23184);
nand U24706 (N_24706,N_23216,N_23920);
nor U24707 (N_24707,N_23167,N_23503);
xor U24708 (N_24708,N_23376,N_23695);
nand U24709 (N_24709,N_23342,N_23608);
xnor U24710 (N_24710,N_23368,N_23327);
and U24711 (N_24711,N_23671,N_23368);
nor U24712 (N_24712,N_23722,N_23051);
xor U24713 (N_24713,N_23061,N_23549);
or U24714 (N_24714,N_23872,N_23393);
and U24715 (N_24715,N_23280,N_23304);
or U24716 (N_24716,N_23985,N_23534);
xor U24717 (N_24717,N_23180,N_23852);
and U24718 (N_24718,N_23527,N_23936);
nand U24719 (N_24719,N_23612,N_23965);
or U24720 (N_24720,N_23726,N_23256);
nor U24721 (N_24721,N_23968,N_23054);
xnor U24722 (N_24722,N_23128,N_23671);
nand U24723 (N_24723,N_23754,N_23731);
and U24724 (N_24724,N_23217,N_23937);
xnor U24725 (N_24725,N_23196,N_23355);
or U24726 (N_24726,N_23316,N_23208);
or U24727 (N_24727,N_23830,N_23952);
or U24728 (N_24728,N_23316,N_23392);
and U24729 (N_24729,N_23904,N_23460);
xor U24730 (N_24730,N_23353,N_23858);
nor U24731 (N_24731,N_23882,N_23435);
and U24732 (N_24732,N_23263,N_23354);
or U24733 (N_24733,N_23525,N_23463);
or U24734 (N_24734,N_23394,N_23127);
or U24735 (N_24735,N_23333,N_23748);
xnor U24736 (N_24736,N_23597,N_23838);
nand U24737 (N_24737,N_23775,N_23307);
nand U24738 (N_24738,N_23349,N_23858);
or U24739 (N_24739,N_23929,N_23838);
nor U24740 (N_24740,N_23609,N_23018);
and U24741 (N_24741,N_23735,N_23141);
xor U24742 (N_24742,N_23016,N_23507);
nand U24743 (N_24743,N_23481,N_23544);
nand U24744 (N_24744,N_23657,N_23595);
xnor U24745 (N_24745,N_23675,N_23959);
and U24746 (N_24746,N_23745,N_23599);
nor U24747 (N_24747,N_23744,N_23072);
xor U24748 (N_24748,N_23216,N_23035);
nand U24749 (N_24749,N_23900,N_23310);
or U24750 (N_24750,N_23380,N_23071);
or U24751 (N_24751,N_23389,N_23503);
and U24752 (N_24752,N_23025,N_23455);
and U24753 (N_24753,N_23180,N_23497);
nor U24754 (N_24754,N_23869,N_23554);
nor U24755 (N_24755,N_23173,N_23682);
nand U24756 (N_24756,N_23855,N_23313);
nand U24757 (N_24757,N_23073,N_23879);
xnor U24758 (N_24758,N_23455,N_23158);
nor U24759 (N_24759,N_23709,N_23056);
or U24760 (N_24760,N_23939,N_23291);
nand U24761 (N_24761,N_23373,N_23404);
nand U24762 (N_24762,N_23670,N_23372);
xor U24763 (N_24763,N_23103,N_23892);
nand U24764 (N_24764,N_23948,N_23331);
or U24765 (N_24765,N_23422,N_23153);
and U24766 (N_24766,N_23059,N_23341);
xor U24767 (N_24767,N_23656,N_23765);
nor U24768 (N_24768,N_23758,N_23918);
nand U24769 (N_24769,N_23607,N_23309);
or U24770 (N_24770,N_23836,N_23667);
xor U24771 (N_24771,N_23166,N_23115);
or U24772 (N_24772,N_23451,N_23206);
or U24773 (N_24773,N_23178,N_23337);
or U24774 (N_24774,N_23385,N_23695);
nor U24775 (N_24775,N_23599,N_23612);
nand U24776 (N_24776,N_23611,N_23373);
or U24777 (N_24777,N_23029,N_23097);
xor U24778 (N_24778,N_23993,N_23633);
xor U24779 (N_24779,N_23682,N_23262);
or U24780 (N_24780,N_23526,N_23730);
nand U24781 (N_24781,N_23218,N_23206);
xor U24782 (N_24782,N_23923,N_23483);
xor U24783 (N_24783,N_23928,N_23781);
or U24784 (N_24784,N_23931,N_23902);
and U24785 (N_24785,N_23466,N_23846);
xor U24786 (N_24786,N_23171,N_23691);
or U24787 (N_24787,N_23436,N_23629);
or U24788 (N_24788,N_23415,N_23178);
nor U24789 (N_24789,N_23199,N_23303);
xnor U24790 (N_24790,N_23057,N_23777);
and U24791 (N_24791,N_23959,N_23180);
nor U24792 (N_24792,N_23340,N_23537);
and U24793 (N_24793,N_23796,N_23806);
and U24794 (N_24794,N_23109,N_23443);
or U24795 (N_24795,N_23446,N_23999);
or U24796 (N_24796,N_23859,N_23129);
nand U24797 (N_24797,N_23436,N_23709);
or U24798 (N_24798,N_23948,N_23823);
or U24799 (N_24799,N_23113,N_23892);
or U24800 (N_24800,N_23517,N_23553);
or U24801 (N_24801,N_23812,N_23921);
xor U24802 (N_24802,N_23508,N_23482);
nor U24803 (N_24803,N_23211,N_23868);
and U24804 (N_24804,N_23984,N_23933);
xnor U24805 (N_24805,N_23870,N_23587);
nand U24806 (N_24806,N_23509,N_23132);
or U24807 (N_24807,N_23197,N_23051);
nand U24808 (N_24808,N_23646,N_23892);
nor U24809 (N_24809,N_23283,N_23026);
or U24810 (N_24810,N_23327,N_23293);
xor U24811 (N_24811,N_23021,N_23937);
nand U24812 (N_24812,N_23064,N_23045);
and U24813 (N_24813,N_23734,N_23236);
or U24814 (N_24814,N_23048,N_23015);
nand U24815 (N_24815,N_23200,N_23009);
nand U24816 (N_24816,N_23042,N_23251);
nand U24817 (N_24817,N_23773,N_23991);
xnor U24818 (N_24818,N_23457,N_23524);
xor U24819 (N_24819,N_23738,N_23794);
nor U24820 (N_24820,N_23666,N_23785);
nand U24821 (N_24821,N_23251,N_23720);
xor U24822 (N_24822,N_23376,N_23190);
nor U24823 (N_24823,N_23777,N_23613);
nor U24824 (N_24824,N_23975,N_23379);
xor U24825 (N_24825,N_23343,N_23403);
nor U24826 (N_24826,N_23244,N_23045);
nand U24827 (N_24827,N_23280,N_23070);
and U24828 (N_24828,N_23002,N_23191);
xor U24829 (N_24829,N_23058,N_23132);
or U24830 (N_24830,N_23961,N_23765);
nand U24831 (N_24831,N_23782,N_23707);
xnor U24832 (N_24832,N_23019,N_23364);
nand U24833 (N_24833,N_23839,N_23794);
and U24834 (N_24834,N_23904,N_23663);
and U24835 (N_24835,N_23049,N_23885);
nand U24836 (N_24836,N_23913,N_23580);
xnor U24837 (N_24837,N_23810,N_23887);
or U24838 (N_24838,N_23814,N_23565);
xor U24839 (N_24839,N_23376,N_23615);
or U24840 (N_24840,N_23794,N_23782);
and U24841 (N_24841,N_23699,N_23597);
nor U24842 (N_24842,N_23106,N_23536);
nand U24843 (N_24843,N_23986,N_23658);
xnor U24844 (N_24844,N_23945,N_23082);
nand U24845 (N_24845,N_23183,N_23012);
and U24846 (N_24846,N_23205,N_23146);
xnor U24847 (N_24847,N_23063,N_23832);
xnor U24848 (N_24848,N_23311,N_23847);
xor U24849 (N_24849,N_23794,N_23757);
nand U24850 (N_24850,N_23530,N_23508);
and U24851 (N_24851,N_23323,N_23395);
xor U24852 (N_24852,N_23851,N_23832);
xnor U24853 (N_24853,N_23701,N_23860);
nand U24854 (N_24854,N_23178,N_23139);
xnor U24855 (N_24855,N_23945,N_23246);
xor U24856 (N_24856,N_23347,N_23239);
and U24857 (N_24857,N_23600,N_23930);
and U24858 (N_24858,N_23800,N_23774);
and U24859 (N_24859,N_23541,N_23380);
and U24860 (N_24860,N_23183,N_23112);
nand U24861 (N_24861,N_23092,N_23049);
nor U24862 (N_24862,N_23324,N_23264);
nor U24863 (N_24863,N_23920,N_23788);
and U24864 (N_24864,N_23302,N_23414);
nor U24865 (N_24865,N_23669,N_23069);
nor U24866 (N_24866,N_23603,N_23576);
and U24867 (N_24867,N_23079,N_23301);
nor U24868 (N_24868,N_23258,N_23551);
or U24869 (N_24869,N_23515,N_23546);
xor U24870 (N_24870,N_23629,N_23343);
or U24871 (N_24871,N_23952,N_23655);
and U24872 (N_24872,N_23667,N_23835);
or U24873 (N_24873,N_23031,N_23135);
or U24874 (N_24874,N_23824,N_23951);
and U24875 (N_24875,N_23119,N_23657);
or U24876 (N_24876,N_23042,N_23767);
and U24877 (N_24877,N_23148,N_23508);
nand U24878 (N_24878,N_23185,N_23353);
nor U24879 (N_24879,N_23717,N_23550);
xor U24880 (N_24880,N_23521,N_23933);
or U24881 (N_24881,N_23268,N_23530);
xor U24882 (N_24882,N_23956,N_23203);
and U24883 (N_24883,N_23320,N_23313);
or U24884 (N_24884,N_23302,N_23793);
nor U24885 (N_24885,N_23288,N_23128);
or U24886 (N_24886,N_23639,N_23957);
or U24887 (N_24887,N_23995,N_23491);
nand U24888 (N_24888,N_23722,N_23793);
or U24889 (N_24889,N_23701,N_23375);
nor U24890 (N_24890,N_23557,N_23904);
nand U24891 (N_24891,N_23265,N_23274);
nand U24892 (N_24892,N_23490,N_23855);
nand U24893 (N_24893,N_23072,N_23599);
xnor U24894 (N_24894,N_23093,N_23880);
and U24895 (N_24895,N_23283,N_23883);
xor U24896 (N_24896,N_23557,N_23032);
and U24897 (N_24897,N_23808,N_23374);
or U24898 (N_24898,N_23049,N_23794);
nor U24899 (N_24899,N_23708,N_23933);
or U24900 (N_24900,N_23453,N_23370);
nand U24901 (N_24901,N_23772,N_23873);
and U24902 (N_24902,N_23263,N_23820);
or U24903 (N_24903,N_23920,N_23449);
or U24904 (N_24904,N_23671,N_23866);
or U24905 (N_24905,N_23507,N_23527);
nand U24906 (N_24906,N_23759,N_23015);
nor U24907 (N_24907,N_23697,N_23441);
nor U24908 (N_24908,N_23620,N_23672);
or U24909 (N_24909,N_23175,N_23052);
and U24910 (N_24910,N_23261,N_23008);
or U24911 (N_24911,N_23477,N_23169);
nor U24912 (N_24912,N_23228,N_23509);
nand U24913 (N_24913,N_23686,N_23774);
nand U24914 (N_24914,N_23375,N_23933);
and U24915 (N_24915,N_23271,N_23063);
nand U24916 (N_24916,N_23264,N_23074);
or U24917 (N_24917,N_23670,N_23184);
nand U24918 (N_24918,N_23165,N_23968);
or U24919 (N_24919,N_23635,N_23750);
or U24920 (N_24920,N_23637,N_23204);
nor U24921 (N_24921,N_23023,N_23706);
and U24922 (N_24922,N_23998,N_23899);
or U24923 (N_24923,N_23015,N_23503);
xnor U24924 (N_24924,N_23176,N_23375);
nor U24925 (N_24925,N_23105,N_23468);
nor U24926 (N_24926,N_23175,N_23028);
or U24927 (N_24927,N_23472,N_23714);
nand U24928 (N_24928,N_23229,N_23757);
xor U24929 (N_24929,N_23378,N_23148);
nor U24930 (N_24930,N_23459,N_23918);
or U24931 (N_24931,N_23265,N_23320);
nor U24932 (N_24932,N_23812,N_23087);
nand U24933 (N_24933,N_23219,N_23153);
and U24934 (N_24934,N_23819,N_23893);
nor U24935 (N_24935,N_23997,N_23778);
nand U24936 (N_24936,N_23801,N_23051);
nand U24937 (N_24937,N_23610,N_23725);
xnor U24938 (N_24938,N_23244,N_23784);
and U24939 (N_24939,N_23711,N_23092);
and U24940 (N_24940,N_23520,N_23842);
xor U24941 (N_24941,N_23401,N_23587);
nor U24942 (N_24942,N_23950,N_23894);
xor U24943 (N_24943,N_23451,N_23502);
and U24944 (N_24944,N_23086,N_23338);
or U24945 (N_24945,N_23236,N_23547);
and U24946 (N_24946,N_23888,N_23102);
and U24947 (N_24947,N_23895,N_23728);
nand U24948 (N_24948,N_23609,N_23034);
nor U24949 (N_24949,N_23829,N_23993);
and U24950 (N_24950,N_23326,N_23685);
or U24951 (N_24951,N_23576,N_23596);
nand U24952 (N_24952,N_23165,N_23212);
nor U24953 (N_24953,N_23245,N_23092);
xnor U24954 (N_24954,N_23427,N_23211);
nand U24955 (N_24955,N_23872,N_23847);
xnor U24956 (N_24956,N_23313,N_23551);
and U24957 (N_24957,N_23481,N_23579);
xnor U24958 (N_24958,N_23864,N_23472);
or U24959 (N_24959,N_23183,N_23356);
nand U24960 (N_24960,N_23873,N_23479);
and U24961 (N_24961,N_23405,N_23770);
and U24962 (N_24962,N_23991,N_23128);
and U24963 (N_24963,N_23522,N_23625);
and U24964 (N_24964,N_23848,N_23663);
and U24965 (N_24965,N_23815,N_23584);
nand U24966 (N_24966,N_23453,N_23288);
nor U24967 (N_24967,N_23952,N_23164);
nor U24968 (N_24968,N_23675,N_23963);
and U24969 (N_24969,N_23125,N_23818);
nand U24970 (N_24970,N_23979,N_23709);
nor U24971 (N_24971,N_23425,N_23433);
or U24972 (N_24972,N_23597,N_23151);
or U24973 (N_24973,N_23178,N_23821);
xor U24974 (N_24974,N_23795,N_23059);
nor U24975 (N_24975,N_23316,N_23722);
and U24976 (N_24976,N_23616,N_23416);
and U24977 (N_24977,N_23980,N_23741);
nor U24978 (N_24978,N_23769,N_23323);
xor U24979 (N_24979,N_23376,N_23692);
nand U24980 (N_24980,N_23489,N_23627);
or U24981 (N_24981,N_23968,N_23807);
and U24982 (N_24982,N_23030,N_23772);
and U24983 (N_24983,N_23674,N_23592);
nor U24984 (N_24984,N_23685,N_23954);
and U24985 (N_24985,N_23175,N_23192);
and U24986 (N_24986,N_23120,N_23456);
nor U24987 (N_24987,N_23336,N_23410);
nor U24988 (N_24988,N_23851,N_23277);
nor U24989 (N_24989,N_23698,N_23438);
nand U24990 (N_24990,N_23858,N_23895);
nand U24991 (N_24991,N_23375,N_23897);
nand U24992 (N_24992,N_23106,N_23712);
xor U24993 (N_24993,N_23248,N_23619);
and U24994 (N_24994,N_23268,N_23835);
nand U24995 (N_24995,N_23015,N_23257);
nor U24996 (N_24996,N_23528,N_23706);
nand U24997 (N_24997,N_23102,N_23850);
nor U24998 (N_24998,N_23554,N_23010);
xnor U24999 (N_24999,N_23235,N_23028);
nor U25000 (N_25000,N_24246,N_24055);
xnor U25001 (N_25001,N_24577,N_24301);
and U25002 (N_25002,N_24544,N_24439);
nand U25003 (N_25003,N_24894,N_24421);
nor U25004 (N_25004,N_24718,N_24463);
or U25005 (N_25005,N_24760,N_24183);
xnor U25006 (N_25006,N_24061,N_24001);
xor U25007 (N_25007,N_24304,N_24141);
xnor U25008 (N_25008,N_24923,N_24038);
nand U25009 (N_25009,N_24773,N_24405);
nor U25010 (N_25010,N_24298,N_24532);
nand U25011 (N_25011,N_24845,N_24646);
nand U25012 (N_25012,N_24391,N_24390);
nor U25013 (N_25013,N_24919,N_24170);
nor U25014 (N_25014,N_24582,N_24809);
nand U25015 (N_25015,N_24967,N_24163);
xnor U25016 (N_25016,N_24393,N_24545);
nor U25017 (N_25017,N_24455,N_24802);
nand U25018 (N_25018,N_24557,N_24999);
nand U25019 (N_25019,N_24364,N_24279);
nand U25020 (N_25020,N_24536,N_24131);
xnor U25021 (N_25021,N_24824,N_24106);
nand U25022 (N_25022,N_24674,N_24158);
or U25023 (N_25023,N_24093,N_24974);
and U25024 (N_25024,N_24542,N_24041);
or U25025 (N_25025,N_24196,N_24933);
xnor U25026 (N_25026,N_24202,N_24368);
or U25027 (N_25027,N_24901,N_24278);
nor U25028 (N_25028,N_24663,N_24852);
and U25029 (N_25029,N_24988,N_24083);
and U25030 (N_25030,N_24281,N_24793);
or U25031 (N_25031,N_24791,N_24282);
and U25032 (N_25032,N_24199,N_24173);
or U25033 (N_25033,N_24494,N_24177);
xor U25034 (N_25034,N_24691,N_24273);
and U25035 (N_25035,N_24152,N_24261);
xor U25036 (N_25036,N_24518,N_24925);
nor U25037 (N_25037,N_24960,N_24594);
or U25038 (N_25038,N_24440,N_24831);
and U25039 (N_25039,N_24539,N_24314);
nor U25040 (N_25040,N_24896,N_24351);
xnor U25041 (N_25041,N_24406,N_24175);
and U25042 (N_25042,N_24937,N_24921);
nand U25043 (N_25043,N_24576,N_24374);
nor U25044 (N_25044,N_24387,N_24514);
nand U25045 (N_25045,N_24699,N_24307);
and U25046 (N_25046,N_24072,N_24251);
nor U25047 (N_25047,N_24610,N_24469);
or U25048 (N_25048,N_24616,N_24157);
nor U25049 (N_25049,N_24633,N_24159);
nand U25050 (N_25050,N_24321,N_24819);
or U25051 (N_25051,N_24748,N_24954);
and U25052 (N_25052,N_24034,N_24741);
and U25053 (N_25053,N_24336,N_24531);
and U25054 (N_25054,N_24655,N_24503);
nand U25055 (N_25055,N_24541,N_24825);
nand U25056 (N_25056,N_24027,N_24111);
xnor U25057 (N_25057,N_24924,N_24909);
or U25058 (N_25058,N_24313,N_24692);
nor U25059 (N_25059,N_24957,N_24046);
nand U25060 (N_25060,N_24964,N_24778);
nand U25061 (N_25061,N_24140,N_24130);
nand U25062 (N_25062,N_24520,N_24452);
nor U25063 (N_25063,N_24795,N_24537);
xnor U25064 (N_25064,N_24398,N_24883);
and U25065 (N_25065,N_24029,N_24839);
and U25066 (N_25066,N_24114,N_24227);
nor U25067 (N_25067,N_24358,N_24898);
xnor U25068 (N_25068,N_24299,N_24436);
nor U25069 (N_25069,N_24165,N_24709);
and U25070 (N_25070,N_24833,N_24977);
nand U25071 (N_25071,N_24206,N_24289);
xnor U25072 (N_25072,N_24458,N_24088);
or U25073 (N_25073,N_24205,N_24681);
xor U25074 (N_25074,N_24510,N_24752);
and U25075 (N_25075,N_24184,N_24640);
nor U25076 (N_25076,N_24983,N_24069);
or U25077 (N_25077,N_24653,N_24203);
nand U25078 (N_25078,N_24892,N_24353);
or U25079 (N_25079,N_24738,N_24065);
or U25080 (N_25080,N_24447,N_24099);
nand U25081 (N_25081,N_24756,N_24888);
nor U25082 (N_25082,N_24036,N_24618);
nand U25083 (N_25083,N_24565,N_24734);
nor U25084 (N_25084,N_24235,N_24932);
nor U25085 (N_25085,N_24776,N_24103);
nand U25086 (N_25086,N_24249,N_24116);
and U25087 (N_25087,N_24325,N_24590);
and U25088 (N_25088,N_24643,N_24993);
xor U25089 (N_25089,N_24252,N_24587);
nor U25090 (N_25090,N_24712,N_24108);
and U25091 (N_25091,N_24953,N_24497);
or U25092 (N_25092,N_24451,N_24425);
nand U25093 (N_25093,N_24651,N_24051);
nor U25094 (N_25094,N_24700,N_24063);
nand U25095 (N_25095,N_24929,N_24850);
xor U25096 (N_25096,N_24904,N_24614);
nand U25097 (N_25097,N_24736,N_24560);
nand U25098 (N_25098,N_24021,N_24223);
or U25099 (N_25099,N_24288,N_24426);
or U25100 (N_25100,N_24349,N_24037);
or U25101 (N_25101,N_24178,N_24475);
nor U25102 (N_25102,N_24829,N_24443);
and U25103 (N_25103,N_24724,N_24574);
and U25104 (N_25104,N_24492,N_24930);
or U25105 (N_25105,N_24630,N_24373);
or U25106 (N_25106,N_24955,N_24613);
or U25107 (N_25107,N_24423,N_24491);
nand U25108 (N_25108,N_24369,N_24316);
or U25109 (N_25109,N_24759,N_24385);
and U25110 (N_25110,N_24271,N_24232);
and U25111 (N_25111,N_24101,N_24876);
and U25112 (N_25112,N_24730,N_24478);
and U25113 (N_25113,N_24354,N_24982);
nor U25114 (N_25114,N_24528,N_24684);
nand U25115 (N_25115,N_24474,N_24127);
or U25116 (N_25116,N_24379,N_24874);
xnor U25117 (N_25117,N_24976,N_24024);
xor U25118 (N_25118,N_24865,N_24145);
nor U25119 (N_25119,N_24318,N_24376);
or U25120 (N_25120,N_24987,N_24556);
nand U25121 (N_25121,N_24326,N_24952);
xnor U25122 (N_25122,N_24840,N_24908);
or U25123 (N_25123,N_24890,N_24333);
or U25124 (N_25124,N_24416,N_24290);
nand U25125 (N_25125,N_24787,N_24637);
or U25126 (N_25126,N_24669,N_24625);
or U25127 (N_25127,N_24507,N_24673);
xor U25128 (N_25128,N_24262,N_24899);
and U25129 (N_25129,N_24464,N_24264);
nand U25130 (N_25130,N_24155,N_24725);
nor U25131 (N_25131,N_24688,N_24062);
xor U25132 (N_25132,N_24784,N_24335);
xnor U25133 (N_25133,N_24240,N_24167);
or U25134 (N_25134,N_24303,N_24608);
nand U25135 (N_25135,N_24465,N_24632);
or U25136 (N_25136,N_24553,N_24000);
xor U25137 (N_25137,N_24025,N_24331);
xnor U25138 (N_25138,N_24562,N_24220);
or U25139 (N_25139,N_24035,N_24149);
and U25140 (N_25140,N_24221,N_24212);
and U25141 (N_25141,N_24498,N_24356);
or U25142 (N_25142,N_24311,N_24509);
xor U25143 (N_25143,N_24887,N_24783);
nor U25144 (N_25144,N_24181,N_24346);
xor U25145 (N_25145,N_24732,N_24030);
and U25146 (N_25146,N_24371,N_24294);
nand U25147 (N_25147,N_24234,N_24182);
nand U25148 (N_25148,N_24857,N_24818);
nor U25149 (N_25149,N_24889,N_24685);
nand U25150 (N_25150,N_24459,N_24715);
nand U25151 (N_25151,N_24073,N_24104);
nor U25152 (N_25152,N_24885,N_24868);
and U25153 (N_25153,N_24767,N_24645);
or U25154 (N_25154,N_24529,N_24779);
and U25155 (N_25155,N_24543,N_24519);
nor U25156 (N_25156,N_24766,N_24702);
nand U25157 (N_25157,N_24657,N_24151);
and U25158 (N_25158,N_24798,N_24597);
nand U25159 (N_25159,N_24838,N_24365);
nand U25160 (N_25160,N_24757,N_24462);
nand U25161 (N_25161,N_24711,N_24812);
nor U25162 (N_25162,N_24785,N_24366);
nand U25163 (N_25163,N_24445,N_24744);
and U25164 (N_25164,N_24635,N_24284);
and U25165 (N_25165,N_24777,N_24926);
and U25166 (N_25166,N_24579,N_24248);
nor U25167 (N_25167,N_24631,N_24031);
xnor U25168 (N_25168,N_24360,N_24012);
or U25169 (N_25169,N_24124,N_24603);
nand U25170 (N_25170,N_24017,N_24677);
nand U25171 (N_25171,N_24676,N_24198);
xor U25172 (N_25172,N_24096,N_24226);
nor U25173 (N_25173,N_24836,N_24753);
nand U25174 (N_25174,N_24241,N_24255);
or U25175 (N_25175,N_24132,N_24270);
nand U25176 (N_25176,N_24694,N_24350);
nand U25177 (N_25177,N_24059,N_24296);
nor U25178 (N_25178,N_24580,N_24142);
or U25179 (N_25179,N_24022,N_24701);
nor U25180 (N_25180,N_24266,N_24547);
or U25181 (N_25181,N_24068,N_24705);
xor U25182 (N_25182,N_24678,N_24512);
and U25183 (N_25183,N_24575,N_24397);
and U25184 (N_25184,N_24292,N_24312);
xnor U25185 (N_25185,N_24230,N_24814);
and U25186 (N_25186,N_24070,N_24972);
nor U25187 (N_25187,N_24995,N_24847);
nor U25188 (N_25188,N_24011,N_24747);
xnor U25189 (N_25189,N_24675,N_24555);
and U25190 (N_25190,N_24432,N_24714);
or U25191 (N_25191,N_24731,N_24665);
and U25192 (N_25192,N_24109,N_24352);
nand U25193 (N_25193,N_24570,N_24242);
or U25194 (N_25194,N_24066,N_24704);
or U25195 (N_25195,N_24985,N_24961);
nor U25196 (N_25196,N_24233,N_24293);
and U25197 (N_25197,N_24064,N_24128);
or U25198 (N_25198,N_24413,N_24723);
nand U25199 (N_25199,N_24189,N_24843);
xor U25200 (N_25200,N_24117,N_24048);
nand U25201 (N_25201,N_24039,N_24735);
xnor U25202 (N_25202,N_24218,N_24323);
or U25203 (N_25203,N_24297,N_24944);
or U25204 (N_25204,N_24375,N_24115);
and U25205 (N_25205,N_24265,N_24895);
nand U25206 (N_25206,N_24834,N_24485);
and U25207 (N_25207,N_24661,N_24045);
xor U25208 (N_25208,N_24214,N_24156);
or U25209 (N_25209,N_24951,N_24092);
nand U25210 (N_25210,N_24496,N_24441);
nand U25211 (N_25211,N_24309,N_24564);
and U25212 (N_25212,N_24229,N_24329);
xor U25213 (N_25213,N_24342,N_24437);
nand U25214 (N_25214,N_24144,N_24384);
or U25215 (N_25215,N_24482,N_24609);
nand U25216 (N_25216,N_24433,N_24372);
or U25217 (N_25217,N_24860,N_24648);
nand U25218 (N_25218,N_24668,N_24863);
nor U25219 (N_25219,N_24906,N_24219);
and U25220 (N_25220,N_24672,N_24363);
nand U25221 (N_25221,N_24774,N_24569);
and U25222 (N_25222,N_24826,N_24522);
and U25223 (N_25223,N_24858,N_24453);
nor U25224 (N_25224,N_24624,N_24081);
and U25225 (N_25225,N_24125,N_24571);
and U25226 (N_25226,N_24018,N_24984);
nor U25227 (N_25227,N_24043,N_24658);
nand U25228 (N_25228,N_24412,N_24135);
or U25229 (N_25229,N_24341,N_24168);
nand U25230 (N_25230,N_24171,N_24193);
xor U25231 (N_25231,N_24471,N_24136);
and U25232 (N_25232,N_24780,N_24508);
nand U25233 (N_25233,N_24044,N_24419);
xor U25234 (N_25234,N_24277,N_24480);
or U25235 (N_25235,N_24728,N_24770);
nor U25236 (N_25236,N_24344,N_24884);
nand U25237 (N_25237,N_24224,N_24495);
xor U25238 (N_25238,N_24717,N_24195);
nor U25239 (N_25239,N_24411,N_24745);
nor U25240 (N_25240,N_24666,N_24856);
nor U25241 (N_25241,N_24291,N_24877);
and U25242 (N_25242,N_24418,N_24882);
and U25243 (N_25243,N_24454,N_24500);
xor U25244 (N_25244,N_24654,N_24566);
and U25245 (N_25245,N_24763,N_24286);
and U25246 (N_25246,N_24094,N_24499);
xnor U25247 (N_25247,N_24164,N_24743);
xnor U25248 (N_25248,N_24615,N_24690);
xor U25249 (N_25249,N_24956,N_24057);
nor U25250 (N_25250,N_24516,N_24968);
or U25251 (N_25251,N_24697,N_24939);
and U25252 (N_25252,N_24370,N_24147);
xnor U25253 (N_25253,N_24862,N_24191);
or U25254 (N_25254,N_24864,N_24851);
and U25255 (N_25255,N_24942,N_24698);
xor U25256 (N_25256,N_24636,N_24805);
or U25257 (N_25257,N_24260,N_24513);
xor U25258 (N_25258,N_24523,N_24917);
or U25259 (N_25259,N_24832,N_24788);
xor U25260 (N_25260,N_24662,N_24197);
xnor U25261 (N_25261,N_24134,N_24584);
nand U25262 (N_25262,N_24589,N_24559);
nand U25263 (N_25263,N_24486,N_24721);
nor U25264 (N_25264,N_24750,N_24345);
nand U25265 (N_25265,N_24970,N_24020);
nor U25266 (N_25266,N_24505,N_24100);
nor U25267 (N_25267,N_24003,N_24595);
and U25268 (N_25268,N_24472,N_24327);
or U25269 (N_25269,N_24764,N_24275);
nand U25270 (N_25270,N_24530,N_24903);
xnor U25271 (N_25271,N_24285,N_24915);
nor U25272 (N_25272,N_24816,N_24386);
and U25273 (N_25273,N_24550,N_24707);
nand U25274 (N_25274,N_24253,N_24225);
xnor U25275 (N_25275,N_24799,N_24879);
nor U25276 (N_25276,N_24841,N_24400);
or U25277 (N_25277,N_24897,N_24607);
and U25278 (N_25278,N_24187,N_24074);
xor U25279 (N_25279,N_24087,N_24913);
or U25280 (N_25280,N_24077,N_24938);
or U25281 (N_25281,N_24755,N_24295);
or U25282 (N_25282,N_24696,N_24593);
and U25283 (N_25283,N_24450,N_24120);
xor U25284 (N_25284,N_24650,N_24981);
nand U25285 (N_25285,N_24190,N_24310);
nand U25286 (N_25286,N_24849,N_24414);
xnor U25287 (N_25287,N_24213,N_24588);
xor U25288 (N_25288,N_24775,N_24146);
xnor U25289 (N_25289,N_24180,N_24986);
and U25290 (N_25290,N_24493,N_24483);
nor U25291 (N_25291,N_24751,N_24830);
or U25292 (N_25292,N_24647,N_24687);
nor U25293 (N_25293,N_24382,N_24706);
nor U25294 (N_25294,N_24016,N_24807);
or U25295 (N_25295,N_24713,N_24431);
xor U25296 (N_25296,N_24058,N_24209);
or U25297 (N_25297,N_24786,N_24664);
nand U25298 (N_25298,N_24754,N_24082);
and U25299 (N_25299,N_24815,N_24238);
nand U25300 (N_25300,N_24546,N_24361);
nor U25301 (N_25301,N_24269,N_24680);
and U25302 (N_25302,N_24481,N_24434);
nand U25303 (N_25303,N_24797,N_24328);
nor U25304 (N_25304,N_24935,N_24800);
nor U25305 (N_25305,N_24533,N_24160);
nand U25306 (N_25306,N_24727,N_24920);
nor U25307 (N_25307,N_24620,N_24015);
nand U25308 (N_25308,N_24438,N_24075);
nor U25309 (N_25309,N_24028,N_24875);
xor U25310 (N_25310,N_24842,N_24444);
nor U25311 (N_25311,N_24283,N_24410);
nor U25312 (N_25312,N_24272,N_24817);
or U25313 (N_25313,N_24552,N_24716);
xor U25314 (N_25314,N_24873,N_24859);
nor U25315 (N_25315,N_24102,N_24097);
xor U25316 (N_25316,N_24322,N_24504);
nor U25317 (N_25317,N_24473,N_24487);
xnor U25318 (N_25318,N_24758,N_24837);
nor U25319 (N_25319,N_24243,N_24112);
xnor U25320 (N_25320,N_24005,N_24404);
and U25321 (N_25321,N_24600,N_24010);
or U25322 (N_25322,N_24257,N_24835);
and U25323 (N_25323,N_24287,N_24040);
nor U25324 (N_25324,N_24804,N_24634);
xor U25325 (N_25325,N_24940,N_24945);
or U25326 (N_25326,N_24330,N_24506);
and U25327 (N_25327,N_24245,N_24305);
xnor U25328 (N_25328,N_24216,N_24162);
nor U25329 (N_25329,N_24172,N_24823);
nor U25330 (N_25330,N_24975,N_24320);
or U25331 (N_25331,N_24334,N_24586);
nor U25332 (N_25332,N_24317,N_24617);
or U25333 (N_25333,N_24084,N_24827);
xor U25334 (N_25334,N_24086,N_24639);
nor U25335 (N_25335,N_24395,N_24470);
xnor U25336 (N_25336,N_24644,N_24948);
nor U25337 (N_25337,N_24378,N_24893);
or U25338 (N_25338,N_24551,N_24820);
nand U25339 (N_25339,N_24477,N_24319);
and U25340 (N_25340,N_24535,N_24971);
xnor U25341 (N_25341,N_24679,N_24990);
nand U25342 (N_25342,N_24403,N_24409);
xnor U25343 (N_25343,N_24392,N_24121);
or U25344 (N_25344,N_24581,N_24340);
and U25345 (N_25345,N_24790,N_24200);
nor U25346 (N_25346,N_24222,N_24592);
and U25347 (N_25347,N_24489,N_24561);
xor U25348 (N_25348,N_24050,N_24407);
nand U25349 (N_25349,N_24768,N_24007);
and U25350 (N_25350,N_24660,N_24091);
nand U25351 (N_25351,N_24947,N_24324);
and U25352 (N_25352,N_24997,N_24710);
or U25353 (N_25353,N_24239,N_24122);
and U25354 (N_25354,N_24578,N_24796);
xnor U25355 (N_25355,N_24527,N_24315);
nand U25356 (N_25356,N_24558,N_24442);
nand U25357 (N_25357,N_24649,N_24720);
xor U25358 (N_25358,N_24258,N_24377);
or U25359 (N_25359,N_24396,N_24060);
nand U25360 (N_25360,N_24231,N_24502);
and U25361 (N_25361,N_24525,N_24907);
nand U25362 (N_25362,N_24962,N_24308);
or U25363 (N_25363,N_24129,N_24813);
nor U25364 (N_25364,N_24501,N_24280);
nand U25365 (N_25365,N_24174,N_24602);
or U25366 (N_25366,N_24612,N_24186);
and U25367 (N_25367,N_24428,N_24009);
or U25368 (N_25368,N_24927,N_24772);
or U25369 (N_25369,N_24161,N_24761);
nor U25370 (N_25370,N_24192,N_24789);
nand U25371 (N_25371,N_24380,N_24049);
xor U25372 (N_25372,N_24166,N_24148);
nand U25373 (N_25373,N_24762,N_24207);
nand U25374 (N_25374,N_24337,N_24362);
or U25375 (N_25375,N_24596,N_24468);
nor U25376 (N_25376,N_24922,N_24682);
nor U25377 (N_25377,N_24461,N_24821);
nor U25378 (N_25378,N_24629,N_24965);
and U25379 (N_25379,N_24019,N_24769);
or U25380 (N_25380,N_24719,N_24381);
nor U25381 (N_25381,N_24306,N_24598);
and U25382 (N_25382,N_24236,N_24123);
or U25383 (N_25383,N_24693,N_24746);
nand U25384 (N_25384,N_24521,N_24388);
or U25385 (N_25385,N_24338,N_24343);
xor U25386 (N_25386,N_24994,N_24568);
or U25387 (N_25387,N_24708,N_24359);
nor U25388 (N_25388,N_24878,N_24765);
or U25389 (N_25389,N_24902,N_24268);
nand U25390 (N_25390,N_24476,N_24729);
xnor U25391 (N_25391,N_24515,N_24417);
nand U25392 (N_25392,N_24511,N_24429);
xnor U25393 (N_25393,N_24274,N_24628);
nor U25394 (N_25394,N_24228,N_24347);
nand U25395 (N_25395,N_24583,N_24861);
and U25396 (N_25396,N_24042,N_24934);
xnor U25397 (N_25397,N_24866,N_24008);
xnor U25398 (N_25398,N_24722,N_24573);
or U25399 (N_25399,N_24169,N_24667);
or U25400 (N_25400,N_24949,N_24211);
or U25401 (N_25401,N_24911,N_24959);
and U25402 (N_25402,N_24803,N_24969);
and U25403 (N_25403,N_24811,N_24958);
xnor U25404 (N_25404,N_24854,N_24150);
nand U25405 (N_25405,N_24383,N_24740);
nor U25406 (N_25406,N_24534,N_24980);
or U25407 (N_25407,N_24399,N_24259);
and U25408 (N_25408,N_24071,N_24963);
nand U25409 (N_25409,N_24052,N_24026);
xnor U25410 (N_25410,N_24076,N_24998);
xor U25411 (N_25411,N_24880,N_24686);
or U25412 (N_25412,N_24659,N_24641);
or U25413 (N_25413,N_24599,N_24139);
nand U25414 (N_25414,N_24742,N_24891);
and U25415 (N_25415,N_24006,N_24126);
and U25416 (N_25416,N_24806,N_24703);
or U25417 (N_25417,N_24201,N_24430);
xnor U25418 (N_25418,N_24867,N_24912);
nor U25419 (N_25419,N_24053,N_24105);
or U25420 (N_25420,N_24871,N_24110);
xnor U25421 (N_25421,N_24881,N_24910);
xnor U25422 (N_25422,N_24978,N_24517);
or U25423 (N_25423,N_24627,N_24916);
xor U25424 (N_25424,N_24733,N_24078);
xor U25425 (N_25425,N_24143,N_24604);
nand U25426 (N_25426,N_24782,N_24946);
xor U25427 (N_25427,N_24449,N_24979);
or U25428 (N_25428,N_24540,N_24348);
nand U25429 (N_25429,N_24210,N_24217);
or U25430 (N_25430,N_24047,N_24781);
nand U25431 (N_25431,N_24176,N_24966);
nor U25432 (N_25432,N_24726,N_24606);
nand U25433 (N_25433,N_24848,N_24204);
xnor U25434 (N_25434,N_24080,N_24456);
or U25435 (N_25435,N_24402,N_24671);
xor U25436 (N_25436,N_24918,N_24991);
nand U25437 (N_25437,N_24822,N_24931);
or U25438 (N_25438,N_24623,N_24208);
xor U25439 (N_25439,N_24992,N_24095);
and U25440 (N_25440,N_24808,N_24810);
and U25441 (N_25441,N_24855,N_24332);
nand U25442 (N_25442,N_24828,N_24973);
xor U25443 (N_25443,N_24113,N_24941);
xor U25444 (N_25444,N_24185,N_24089);
xnor U25445 (N_25445,N_24107,N_24137);
nand U25446 (N_25446,N_24263,N_24119);
xnor U25447 (N_25447,N_24526,N_24611);
or U25448 (N_25448,N_24215,N_24572);
xnor U25449 (N_25449,N_24652,N_24626);
and U25450 (N_25450,N_24401,N_24154);
and U25451 (N_25451,N_24355,N_24032);
nand U25452 (N_25452,N_24567,N_24886);
nand U25453 (N_25453,N_24642,N_24563);
nor U25454 (N_25454,N_24622,N_24300);
nor U25455 (N_25455,N_24928,N_24548);
xnor U25456 (N_25456,N_24339,N_24002);
or U25457 (N_25457,N_24749,N_24394);
xnor U25458 (N_25458,N_24133,N_24118);
nor U25459 (N_25459,N_24689,N_24254);
xor U25460 (N_25460,N_24524,N_24794);
or U25461 (N_25461,N_24415,N_24554);
and U25462 (N_25462,N_24638,N_24585);
nand U25463 (N_25463,N_24619,N_24737);
or U25464 (N_25464,N_24844,N_24389);
xor U25465 (N_25465,N_24367,N_24256);
nor U25466 (N_25466,N_24601,N_24943);
or U25467 (N_25467,N_24188,N_24422);
or U25468 (N_25468,N_24448,N_24179);
or U25469 (N_25469,N_24138,N_24357);
or U25470 (N_25470,N_24023,N_24670);
xnor U25471 (N_25471,N_24079,N_24989);
or U25472 (N_25472,N_24090,N_24739);
xnor U25473 (N_25473,N_24853,N_24771);
xnor U25474 (N_25474,N_24460,N_24244);
and U25475 (N_25475,N_24408,N_24950);
and U25476 (N_25476,N_24914,N_24695);
xor U25477 (N_25477,N_24484,N_24549);
or U25478 (N_25478,N_24420,N_24056);
nor U25479 (N_25479,N_24247,N_24591);
nand U25480 (N_25480,N_24446,N_24457);
xnor U25481 (N_25481,N_24656,N_24900);
and U25482 (N_25482,N_24792,N_24237);
or U25483 (N_25483,N_24435,N_24067);
or U25484 (N_25484,N_24466,N_24872);
or U25485 (N_25485,N_24870,N_24427);
xnor U25486 (N_25486,N_24479,N_24004);
xor U25487 (N_25487,N_24801,N_24424);
xnor U25488 (N_25488,N_24538,N_24467);
or U25489 (N_25489,N_24153,N_24054);
or U25490 (N_25490,N_24302,N_24846);
and U25491 (N_25491,N_24267,N_24033);
and U25492 (N_25492,N_24276,N_24488);
and U25493 (N_25493,N_24683,N_24605);
nor U25494 (N_25494,N_24085,N_24869);
or U25495 (N_25495,N_24905,N_24194);
nand U25496 (N_25496,N_24936,N_24250);
and U25497 (N_25497,N_24621,N_24013);
xor U25498 (N_25498,N_24014,N_24490);
or U25499 (N_25499,N_24098,N_24996);
and U25500 (N_25500,N_24510,N_24139);
nand U25501 (N_25501,N_24811,N_24286);
xor U25502 (N_25502,N_24489,N_24864);
nand U25503 (N_25503,N_24048,N_24598);
nor U25504 (N_25504,N_24512,N_24861);
nor U25505 (N_25505,N_24262,N_24002);
and U25506 (N_25506,N_24734,N_24602);
or U25507 (N_25507,N_24153,N_24727);
and U25508 (N_25508,N_24362,N_24751);
and U25509 (N_25509,N_24546,N_24454);
nor U25510 (N_25510,N_24254,N_24579);
or U25511 (N_25511,N_24928,N_24565);
or U25512 (N_25512,N_24085,N_24801);
nand U25513 (N_25513,N_24833,N_24064);
nor U25514 (N_25514,N_24891,N_24078);
or U25515 (N_25515,N_24184,N_24946);
or U25516 (N_25516,N_24463,N_24065);
nor U25517 (N_25517,N_24674,N_24080);
and U25518 (N_25518,N_24730,N_24843);
nor U25519 (N_25519,N_24644,N_24405);
nor U25520 (N_25520,N_24453,N_24010);
nand U25521 (N_25521,N_24355,N_24588);
or U25522 (N_25522,N_24974,N_24655);
or U25523 (N_25523,N_24192,N_24854);
xor U25524 (N_25524,N_24112,N_24696);
and U25525 (N_25525,N_24511,N_24132);
nor U25526 (N_25526,N_24413,N_24110);
nor U25527 (N_25527,N_24709,N_24588);
xnor U25528 (N_25528,N_24974,N_24969);
or U25529 (N_25529,N_24485,N_24060);
nand U25530 (N_25530,N_24384,N_24288);
and U25531 (N_25531,N_24035,N_24019);
xnor U25532 (N_25532,N_24687,N_24416);
xnor U25533 (N_25533,N_24798,N_24982);
xor U25534 (N_25534,N_24499,N_24852);
or U25535 (N_25535,N_24627,N_24084);
and U25536 (N_25536,N_24546,N_24497);
nor U25537 (N_25537,N_24272,N_24026);
nor U25538 (N_25538,N_24311,N_24577);
and U25539 (N_25539,N_24261,N_24182);
or U25540 (N_25540,N_24492,N_24553);
or U25541 (N_25541,N_24043,N_24996);
or U25542 (N_25542,N_24408,N_24399);
and U25543 (N_25543,N_24176,N_24637);
or U25544 (N_25544,N_24015,N_24616);
or U25545 (N_25545,N_24749,N_24231);
xor U25546 (N_25546,N_24221,N_24935);
xor U25547 (N_25547,N_24078,N_24552);
xnor U25548 (N_25548,N_24974,N_24983);
nand U25549 (N_25549,N_24056,N_24537);
nor U25550 (N_25550,N_24260,N_24826);
and U25551 (N_25551,N_24964,N_24351);
xor U25552 (N_25552,N_24948,N_24742);
or U25553 (N_25553,N_24738,N_24651);
nor U25554 (N_25554,N_24650,N_24398);
nor U25555 (N_25555,N_24468,N_24514);
and U25556 (N_25556,N_24913,N_24872);
or U25557 (N_25557,N_24117,N_24533);
or U25558 (N_25558,N_24770,N_24396);
nor U25559 (N_25559,N_24836,N_24031);
and U25560 (N_25560,N_24719,N_24555);
xnor U25561 (N_25561,N_24787,N_24960);
xor U25562 (N_25562,N_24457,N_24392);
nor U25563 (N_25563,N_24460,N_24227);
and U25564 (N_25564,N_24670,N_24270);
and U25565 (N_25565,N_24751,N_24814);
nor U25566 (N_25566,N_24476,N_24009);
xnor U25567 (N_25567,N_24305,N_24237);
nor U25568 (N_25568,N_24809,N_24613);
nand U25569 (N_25569,N_24675,N_24128);
xnor U25570 (N_25570,N_24246,N_24244);
nor U25571 (N_25571,N_24121,N_24298);
nand U25572 (N_25572,N_24414,N_24367);
nand U25573 (N_25573,N_24009,N_24726);
or U25574 (N_25574,N_24522,N_24825);
and U25575 (N_25575,N_24144,N_24556);
nand U25576 (N_25576,N_24569,N_24138);
xnor U25577 (N_25577,N_24013,N_24896);
nor U25578 (N_25578,N_24554,N_24661);
or U25579 (N_25579,N_24286,N_24301);
or U25580 (N_25580,N_24606,N_24824);
nor U25581 (N_25581,N_24998,N_24891);
nand U25582 (N_25582,N_24792,N_24115);
nor U25583 (N_25583,N_24800,N_24631);
or U25584 (N_25584,N_24110,N_24341);
and U25585 (N_25585,N_24073,N_24163);
nor U25586 (N_25586,N_24901,N_24720);
nor U25587 (N_25587,N_24915,N_24214);
or U25588 (N_25588,N_24250,N_24493);
xnor U25589 (N_25589,N_24065,N_24491);
nand U25590 (N_25590,N_24831,N_24713);
nand U25591 (N_25591,N_24863,N_24694);
nand U25592 (N_25592,N_24899,N_24032);
nand U25593 (N_25593,N_24012,N_24067);
and U25594 (N_25594,N_24964,N_24233);
or U25595 (N_25595,N_24232,N_24972);
or U25596 (N_25596,N_24751,N_24714);
xnor U25597 (N_25597,N_24183,N_24771);
xnor U25598 (N_25598,N_24606,N_24267);
nand U25599 (N_25599,N_24406,N_24383);
and U25600 (N_25600,N_24402,N_24571);
xor U25601 (N_25601,N_24192,N_24015);
or U25602 (N_25602,N_24352,N_24532);
xor U25603 (N_25603,N_24150,N_24222);
nand U25604 (N_25604,N_24058,N_24998);
nor U25605 (N_25605,N_24900,N_24770);
xnor U25606 (N_25606,N_24548,N_24625);
nor U25607 (N_25607,N_24217,N_24047);
nor U25608 (N_25608,N_24235,N_24234);
nand U25609 (N_25609,N_24540,N_24743);
xnor U25610 (N_25610,N_24674,N_24467);
and U25611 (N_25611,N_24182,N_24310);
nand U25612 (N_25612,N_24711,N_24800);
nand U25613 (N_25613,N_24440,N_24780);
or U25614 (N_25614,N_24513,N_24163);
xnor U25615 (N_25615,N_24471,N_24181);
xnor U25616 (N_25616,N_24565,N_24275);
and U25617 (N_25617,N_24136,N_24113);
xnor U25618 (N_25618,N_24692,N_24596);
nand U25619 (N_25619,N_24785,N_24658);
nand U25620 (N_25620,N_24091,N_24407);
nand U25621 (N_25621,N_24210,N_24412);
and U25622 (N_25622,N_24565,N_24477);
or U25623 (N_25623,N_24897,N_24950);
and U25624 (N_25624,N_24797,N_24418);
or U25625 (N_25625,N_24124,N_24759);
and U25626 (N_25626,N_24134,N_24346);
xnor U25627 (N_25627,N_24051,N_24819);
xnor U25628 (N_25628,N_24716,N_24833);
nand U25629 (N_25629,N_24048,N_24290);
nor U25630 (N_25630,N_24217,N_24952);
or U25631 (N_25631,N_24477,N_24963);
and U25632 (N_25632,N_24904,N_24114);
or U25633 (N_25633,N_24305,N_24508);
nand U25634 (N_25634,N_24302,N_24370);
xnor U25635 (N_25635,N_24558,N_24415);
and U25636 (N_25636,N_24077,N_24788);
or U25637 (N_25637,N_24345,N_24642);
xnor U25638 (N_25638,N_24072,N_24938);
and U25639 (N_25639,N_24289,N_24437);
nand U25640 (N_25640,N_24513,N_24994);
or U25641 (N_25641,N_24480,N_24018);
and U25642 (N_25642,N_24815,N_24701);
nand U25643 (N_25643,N_24560,N_24851);
nor U25644 (N_25644,N_24287,N_24592);
nor U25645 (N_25645,N_24591,N_24148);
nor U25646 (N_25646,N_24487,N_24102);
nor U25647 (N_25647,N_24622,N_24437);
or U25648 (N_25648,N_24154,N_24869);
nand U25649 (N_25649,N_24994,N_24879);
nand U25650 (N_25650,N_24099,N_24305);
nor U25651 (N_25651,N_24963,N_24578);
xor U25652 (N_25652,N_24146,N_24429);
nor U25653 (N_25653,N_24585,N_24672);
or U25654 (N_25654,N_24840,N_24195);
nor U25655 (N_25655,N_24106,N_24873);
nor U25656 (N_25656,N_24313,N_24033);
nor U25657 (N_25657,N_24970,N_24088);
xnor U25658 (N_25658,N_24578,N_24576);
nor U25659 (N_25659,N_24824,N_24244);
nand U25660 (N_25660,N_24785,N_24825);
xor U25661 (N_25661,N_24825,N_24169);
or U25662 (N_25662,N_24311,N_24591);
nor U25663 (N_25663,N_24233,N_24193);
xnor U25664 (N_25664,N_24687,N_24592);
nand U25665 (N_25665,N_24761,N_24872);
or U25666 (N_25666,N_24008,N_24980);
nor U25667 (N_25667,N_24294,N_24022);
or U25668 (N_25668,N_24685,N_24438);
nor U25669 (N_25669,N_24058,N_24856);
and U25670 (N_25670,N_24926,N_24153);
nand U25671 (N_25671,N_24643,N_24663);
xor U25672 (N_25672,N_24192,N_24048);
nor U25673 (N_25673,N_24690,N_24523);
nor U25674 (N_25674,N_24208,N_24070);
nand U25675 (N_25675,N_24649,N_24293);
nor U25676 (N_25676,N_24617,N_24147);
and U25677 (N_25677,N_24476,N_24306);
nor U25678 (N_25678,N_24076,N_24139);
nand U25679 (N_25679,N_24204,N_24712);
or U25680 (N_25680,N_24567,N_24773);
or U25681 (N_25681,N_24908,N_24391);
nand U25682 (N_25682,N_24698,N_24195);
and U25683 (N_25683,N_24949,N_24697);
nor U25684 (N_25684,N_24988,N_24034);
nor U25685 (N_25685,N_24813,N_24594);
nand U25686 (N_25686,N_24128,N_24120);
nand U25687 (N_25687,N_24743,N_24112);
or U25688 (N_25688,N_24234,N_24328);
nand U25689 (N_25689,N_24335,N_24410);
and U25690 (N_25690,N_24589,N_24762);
nand U25691 (N_25691,N_24563,N_24961);
or U25692 (N_25692,N_24048,N_24835);
nand U25693 (N_25693,N_24493,N_24910);
and U25694 (N_25694,N_24472,N_24072);
xnor U25695 (N_25695,N_24895,N_24033);
and U25696 (N_25696,N_24489,N_24979);
or U25697 (N_25697,N_24775,N_24405);
and U25698 (N_25698,N_24561,N_24316);
or U25699 (N_25699,N_24117,N_24023);
or U25700 (N_25700,N_24397,N_24645);
nor U25701 (N_25701,N_24478,N_24036);
or U25702 (N_25702,N_24724,N_24008);
nor U25703 (N_25703,N_24234,N_24726);
or U25704 (N_25704,N_24257,N_24657);
or U25705 (N_25705,N_24236,N_24179);
nand U25706 (N_25706,N_24282,N_24412);
and U25707 (N_25707,N_24087,N_24290);
and U25708 (N_25708,N_24243,N_24478);
or U25709 (N_25709,N_24488,N_24251);
nor U25710 (N_25710,N_24678,N_24919);
nand U25711 (N_25711,N_24043,N_24964);
nand U25712 (N_25712,N_24388,N_24924);
nand U25713 (N_25713,N_24724,N_24444);
nand U25714 (N_25714,N_24038,N_24962);
nand U25715 (N_25715,N_24147,N_24143);
nand U25716 (N_25716,N_24725,N_24679);
nor U25717 (N_25717,N_24800,N_24017);
nand U25718 (N_25718,N_24331,N_24732);
or U25719 (N_25719,N_24747,N_24956);
nand U25720 (N_25720,N_24180,N_24734);
xnor U25721 (N_25721,N_24940,N_24835);
nand U25722 (N_25722,N_24510,N_24422);
nand U25723 (N_25723,N_24322,N_24025);
nor U25724 (N_25724,N_24680,N_24282);
nor U25725 (N_25725,N_24797,N_24298);
or U25726 (N_25726,N_24376,N_24916);
xor U25727 (N_25727,N_24258,N_24133);
nand U25728 (N_25728,N_24245,N_24458);
and U25729 (N_25729,N_24817,N_24224);
or U25730 (N_25730,N_24473,N_24898);
and U25731 (N_25731,N_24257,N_24033);
nor U25732 (N_25732,N_24388,N_24503);
nor U25733 (N_25733,N_24472,N_24107);
or U25734 (N_25734,N_24049,N_24415);
nand U25735 (N_25735,N_24053,N_24747);
or U25736 (N_25736,N_24950,N_24225);
and U25737 (N_25737,N_24193,N_24982);
or U25738 (N_25738,N_24360,N_24837);
or U25739 (N_25739,N_24788,N_24253);
or U25740 (N_25740,N_24209,N_24272);
nand U25741 (N_25741,N_24225,N_24679);
nor U25742 (N_25742,N_24205,N_24842);
and U25743 (N_25743,N_24782,N_24315);
xor U25744 (N_25744,N_24123,N_24441);
nor U25745 (N_25745,N_24383,N_24673);
xor U25746 (N_25746,N_24170,N_24477);
nor U25747 (N_25747,N_24748,N_24512);
nand U25748 (N_25748,N_24935,N_24516);
or U25749 (N_25749,N_24001,N_24867);
and U25750 (N_25750,N_24025,N_24006);
and U25751 (N_25751,N_24578,N_24311);
nand U25752 (N_25752,N_24012,N_24721);
or U25753 (N_25753,N_24434,N_24876);
nand U25754 (N_25754,N_24732,N_24583);
xor U25755 (N_25755,N_24896,N_24073);
or U25756 (N_25756,N_24018,N_24926);
xor U25757 (N_25757,N_24099,N_24333);
and U25758 (N_25758,N_24286,N_24271);
or U25759 (N_25759,N_24282,N_24684);
and U25760 (N_25760,N_24023,N_24736);
or U25761 (N_25761,N_24525,N_24474);
xor U25762 (N_25762,N_24402,N_24468);
nor U25763 (N_25763,N_24786,N_24298);
and U25764 (N_25764,N_24180,N_24082);
or U25765 (N_25765,N_24568,N_24186);
nand U25766 (N_25766,N_24793,N_24536);
nor U25767 (N_25767,N_24136,N_24672);
and U25768 (N_25768,N_24580,N_24335);
or U25769 (N_25769,N_24549,N_24620);
nand U25770 (N_25770,N_24192,N_24300);
nand U25771 (N_25771,N_24554,N_24644);
nor U25772 (N_25772,N_24244,N_24357);
and U25773 (N_25773,N_24993,N_24960);
or U25774 (N_25774,N_24594,N_24358);
and U25775 (N_25775,N_24017,N_24647);
and U25776 (N_25776,N_24006,N_24852);
nor U25777 (N_25777,N_24219,N_24192);
nand U25778 (N_25778,N_24113,N_24256);
and U25779 (N_25779,N_24405,N_24736);
nand U25780 (N_25780,N_24772,N_24637);
nand U25781 (N_25781,N_24619,N_24300);
nand U25782 (N_25782,N_24449,N_24289);
and U25783 (N_25783,N_24018,N_24618);
nand U25784 (N_25784,N_24203,N_24564);
nand U25785 (N_25785,N_24963,N_24708);
and U25786 (N_25786,N_24868,N_24027);
nor U25787 (N_25787,N_24600,N_24634);
or U25788 (N_25788,N_24342,N_24970);
and U25789 (N_25789,N_24712,N_24576);
nor U25790 (N_25790,N_24559,N_24701);
nor U25791 (N_25791,N_24787,N_24941);
nand U25792 (N_25792,N_24426,N_24676);
xor U25793 (N_25793,N_24350,N_24496);
and U25794 (N_25794,N_24550,N_24790);
xnor U25795 (N_25795,N_24924,N_24404);
xnor U25796 (N_25796,N_24419,N_24155);
xnor U25797 (N_25797,N_24569,N_24393);
nor U25798 (N_25798,N_24807,N_24331);
nor U25799 (N_25799,N_24109,N_24227);
and U25800 (N_25800,N_24497,N_24588);
and U25801 (N_25801,N_24111,N_24669);
xor U25802 (N_25802,N_24516,N_24863);
xnor U25803 (N_25803,N_24087,N_24552);
nand U25804 (N_25804,N_24420,N_24235);
xnor U25805 (N_25805,N_24011,N_24394);
and U25806 (N_25806,N_24689,N_24544);
or U25807 (N_25807,N_24689,N_24271);
nor U25808 (N_25808,N_24919,N_24892);
nor U25809 (N_25809,N_24222,N_24016);
nor U25810 (N_25810,N_24261,N_24922);
xnor U25811 (N_25811,N_24320,N_24877);
or U25812 (N_25812,N_24893,N_24736);
or U25813 (N_25813,N_24780,N_24854);
nand U25814 (N_25814,N_24537,N_24417);
and U25815 (N_25815,N_24643,N_24931);
xnor U25816 (N_25816,N_24136,N_24523);
or U25817 (N_25817,N_24065,N_24693);
and U25818 (N_25818,N_24401,N_24357);
xnor U25819 (N_25819,N_24989,N_24256);
nand U25820 (N_25820,N_24437,N_24725);
or U25821 (N_25821,N_24427,N_24655);
or U25822 (N_25822,N_24072,N_24841);
or U25823 (N_25823,N_24021,N_24465);
or U25824 (N_25824,N_24918,N_24568);
nand U25825 (N_25825,N_24298,N_24858);
and U25826 (N_25826,N_24649,N_24794);
nor U25827 (N_25827,N_24860,N_24322);
nor U25828 (N_25828,N_24389,N_24993);
nand U25829 (N_25829,N_24431,N_24030);
nor U25830 (N_25830,N_24075,N_24558);
nand U25831 (N_25831,N_24313,N_24511);
or U25832 (N_25832,N_24570,N_24354);
and U25833 (N_25833,N_24546,N_24903);
nor U25834 (N_25834,N_24643,N_24586);
or U25835 (N_25835,N_24220,N_24061);
and U25836 (N_25836,N_24341,N_24623);
or U25837 (N_25837,N_24053,N_24378);
nor U25838 (N_25838,N_24654,N_24082);
xnor U25839 (N_25839,N_24101,N_24882);
xor U25840 (N_25840,N_24731,N_24500);
xnor U25841 (N_25841,N_24226,N_24388);
and U25842 (N_25842,N_24572,N_24635);
xor U25843 (N_25843,N_24424,N_24359);
nor U25844 (N_25844,N_24519,N_24247);
or U25845 (N_25845,N_24875,N_24591);
and U25846 (N_25846,N_24931,N_24958);
xnor U25847 (N_25847,N_24961,N_24436);
nor U25848 (N_25848,N_24313,N_24233);
or U25849 (N_25849,N_24392,N_24174);
nor U25850 (N_25850,N_24700,N_24783);
and U25851 (N_25851,N_24896,N_24141);
xor U25852 (N_25852,N_24752,N_24945);
nor U25853 (N_25853,N_24015,N_24764);
and U25854 (N_25854,N_24013,N_24948);
and U25855 (N_25855,N_24440,N_24827);
nand U25856 (N_25856,N_24526,N_24615);
xor U25857 (N_25857,N_24667,N_24427);
or U25858 (N_25858,N_24009,N_24782);
nand U25859 (N_25859,N_24035,N_24625);
and U25860 (N_25860,N_24536,N_24826);
xnor U25861 (N_25861,N_24397,N_24596);
nand U25862 (N_25862,N_24482,N_24231);
or U25863 (N_25863,N_24921,N_24594);
xnor U25864 (N_25864,N_24543,N_24294);
nor U25865 (N_25865,N_24427,N_24867);
nand U25866 (N_25866,N_24392,N_24823);
and U25867 (N_25867,N_24020,N_24115);
nor U25868 (N_25868,N_24450,N_24890);
xnor U25869 (N_25869,N_24491,N_24218);
xnor U25870 (N_25870,N_24040,N_24609);
xnor U25871 (N_25871,N_24753,N_24090);
nor U25872 (N_25872,N_24933,N_24721);
and U25873 (N_25873,N_24929,N_24493);
nor U25874 (N_25874,N_24071,N_24824);
nand U25875 (N_25875,N_24972,N_24186);
and U25876 (N_25876,N_24813,N_24629);
or U25877 (N_25877,N_24244,N_24050);
xnor U25878 (N_25878,N_24704,N_24777);
nand U25879 (N_25879,N_24301,N_24182);
nand U25880 (N_25880,N_24428,N_24120);
xnor U25881 (N_25881,N_24835,N_24845);
or U25882 (N_25882,N_24255,N_24153);
nor U25883 (N_25883,N_24418,N_24144);
or U25884 (N_25884,N_24290,N_24567);
or U25885 (N_25885,N_24485,N_24128);
or U25886 (N_25886,N_24067,N_24945);
xor U25887 (N_25887,N_24161,N_24648);
and U25888 (N_25888,N_24018,N_24864);
xor U25889 (N_25889,N_24161,N_24995);
or U25890 (N_25890,N_24762,N_24855);
nor U25891 (N_25891,N_24299,N_24964);
xor U25892 (N_25892,N_24840,N_24637);
xor U25893 (N_25893,N_24753,N_24594);
xor U25894 (N_25894,N_24850,N_24528);
nor U25895 (N_25895,N_24212,N_24369);
xnor U25896 (N_25896,N_24638,N_24652);
or U25897 (N_25897,N_24545,N_24475);
nor U25898 (N_25898,N_24059,N_24820);
nor U25899 (N_25899,N_24451,N_24236);
and U25900 (N_25900,N_24069,N_24385);
or U25901 (N_25901,N_24625,N_24758);
xnor U25902 (N_25902,N_24582,N_24715);
or U25903 (N_25903,N_24288,N_24909);
and U25904 (N_25904,N_24883,N_24539);
nor U25905 (N_25905,N_24955,N_24780);
or U25906 (N_25906,N_24779,N_24060);
xnor U25907 (N_25907,N_24425,N_24992);
nor U25908 (N_25908,N_24265,N_24733);
nor U25909 (N_25909,N_24013,N_24589);
nor U25910 (N_25910,N_24464,N_24938);
or U25911 (N_25911,N_24189,N_24131);
and U25912 (N_25912,N_24922,N_24140);
nor U25913 (N_25913,N_24713,N_24226);
or U25914 (N_25914,N_24218,N_24877);
nor U25915 (N_25915,N_24743,N_24571);
nand U25916 (N_25916,N_24258,N_24810);
and U25917 (N_25917,N_24216,N_24923);
nor U25918 (N_25918,N_24366,N_24632);
nor U25919 (N_25919,N_24815,N_24443);
and U25920 (N_25920,N_24069,N_24042);
xor U25921 (N_25921,N_24209,N_24732);
nand U25922 (N_25922,N_24946,N_24450);
nand U25923 (N_25923,N_24764,N_24841);
or U25924 (N_25924,N_24107,N_24911);
nand U25925 (N_25925,N_24930,N_24095);
nand U25926 (N_25926,N_24804,N_24780);
nor U25927 (N_25927,N_24600,N_24839);
xor U25928 (N_25928,N_24369,N_24474);
nor U25929 (N_25929,N_24001,N_24505);
and U25930 (N_25930,N_24591,N_24979);
or U25931 (N_25931,N_24213,N_24404);
nor U25932 (N_25932,N_24381,N_24687);
nand U25933 (N_25933,N_24115,N_24516);
xnor U25934 (N_25934,N_24308,N_24293);
or U25935 (N_25935,N_24617,N_24677);
and U25936 (N_25936,N_24513,N_24199);
nand U25937 (N_25937,N_24438,N_24453);
xnor U25938 (N_25938,N_24738,N_24247);
xnor U25939 (N_25939,N_24596,N_24617);
xor U25940 (N_25940,N_24842,N_24034);
xor U25941 (N_25941,N_24985,N_24340);
and U25942 (N_25942,N_24840,N_24507);
nor U25943 (N_25943,N_24073,N_24666);
and U25944 (N_25944,N_24115,N_24143);
nand U25945 (N_25945,N_24509,N_24303);
xor U25946 (N_25946,N_24737,N_24572);
xnor U25947 (N_25947,N_24380,N_24098);
and U25948 (N_25948,N_24278,N_24510);
nand U25949 (N_25949,N_24570,N_24791);
nand U25950 (N_25950,N_24600,N_24309);
and U25951 (N_25951,N_24099,N_24560);
and U25952 (N_25952,N_24756,N_24674);
and U25953 (N_25953,N_24464,N_24125);
or U25954 (N_25954,N_24461,N_24655);
xor U25955 (N_25955,N_24347,N_24191);
xnor U25956 (N_25956,N_24090,N_24028);
or U25957 (N_25957,N_24739,N_24427);
xor U25958 (N_25958,N_24400,N_24794);
or U25959 (N_25959,N_24282,N_24447);
xor U25960 (N_25960,N_24084,N_24726);
nand U25961 (N_25961,N_24137,N_24129);
xor U25962 (N_25962,N_24524,N_24925);
or U25963 (N_25963,N_24922,N_24601);
nand U25964 (N_25964,N_24015,N_24605);
and U25965 (N_25965,N_24109,N_24219);
or U25966 (N_25966,N_24567,N_24979);
nand U25967 (N_25967,N_24258,N_24279);
xor U25968 (N_25968,N_24372,N_24148);
or U25969 (N_25969,N_24174,N_24896);
or U25970 (N_25970,N_24838,N_24310);
or U25971 (N_25971,N_24436,N_24409);
or U25972 (N_25972,N_24208,N_24304);
and U25973 (N_25973,N_24996,N_24312);
and U25974 (N_25974,N_24266,N_24372);
nor U25975 (N_25975,N_24897,N_24719);
xor U25976 (N_25976,N_24569,N_24444);
nor U25977 (N_25977,N_24976,N_24420);
nand U25978 (N_25978,N_24675,N_24394);
nor U25979 (N_25979,N_24727,N_24669);
nor U25980 (N_25980,N_24955,N_24337);
xnor U25981 (N_25981,N_24912,N_24194);
and U25982 (N_25982,N_24394,N_24537);
xor U25983 (N_25983,N_24385,N_24311);
nor U25984 (N_25984,N_24397,N_24200);
nor U25985 (N_25985,N_24230,N_24023);
or U25986 (N_25986,N_24403,N_24184);
nor U25987 (N_25987,N_24792,N_24461);
and U25988 (N_25988,N_24379,N_24836);
xor U25989 (N_25989,N_24255,N_24370);
nor U25990 (N_25990,N_24918,N_24851);
and U25991 (N_25991,N_24471,N_24925);
or U25992 (N_25992,N_24271,N_24729);
nand U25993 (N_25993,N_24047,N_24258);
nor U25994 (N_25994,N_24000,N_24213);
or U25995 (N_25995,N_24541,N_24684);
and U25996 (N_25996,N_24838,N_24421);
and U25997 (N_25997,N_24758,N_24528);
and U25998 (N_25998,N_24986,N_24731);
nor U25999 (N_25999,N_24369,N_24002);
and U26000 (N_26000,N_25256,N_25948);
nand U26001 (N_26001,N_25670,N_25831);
xor U26002 (N_26002,N_25559,N_25403);
nand U26003 (N_26003,N_25995,N_25111);
or U26004 (N_26004,N_25088,N_25378);
or U26005 (N_26005,N_25449,N_25472);
and U26006 (N_26006,N_25060,N_25025);
nand U26007 (N_26007,N_25090,N_25194);
nand U26008 (N_26008,N_25187,N_25599);
nor U26009 (N_26009,N_25035,N_25476);
or U26010 (N_26010,N_25807,N_25844);
nand U26011 (N_26011,N_25118,N_25855);
nand U26012 (N_26012,N_25487,N_25655);
and U26013 (N_26013,N_25873,N_25737);
or U26014 (N_26014,N_25624,N_25836);
and U26015 (N_26015,N_25799,N_25208);
or U26016 (N_26016,N_25997,N_25993);
nand U26017 (N_26017,N_25897,N_25164);
xnor U26018 (N_26018,N_25261,N_25656);
and U26019 (N_26019,N_25399,N_25311);
nor U26020 (N_26020,N_25486,N_25499);
or U26021 (N_26021,N_25241,N_25113);
nand U26022 (N_26022,N_25019,N_25856);
nand U26023 (N_26023,N_25646,N_25020);
nand U26024 (N_26024,N_25409,N_25264);
or U26025 (N_26025,N_25772,N_25752);
nand U26026 (N_26026,N_25453,N_25785);
xnor U26027 (N_26027,N_25732,N_25602);
and U26028 (N_26028,N_25571,N_25673);
nand U26029 (N_26029,N_25628,N_25106);
and U26030 (N_26030,N_25105,N_25136);
xnor U26031 (N_26031,N_25726,N_25991);
or U26032 (N_26032,N_25258,N_25355);
xnor U26033 (N_26033,N_25994,N_25288);
nand U26034 (N_26034,N_25653,N_25826);
and U26035 (N_26035,N_25488,N_25870);
and U26036 (N_26036,N_25346,N_25260);
and U26037 (N_26037,N_25824,N_25102);
nand U26038 (N_26038,N_25617,N_25362);
or U26039 (N_26039,N_25871,N_25689);
and U26040 (N_26040,N_25473,N_25648);
nor U26041 (N_26041,N_25928,N_25998);
xor U26042 (N_26042,N_25698,N_25846);
and U26043 (N_26043,N_25370,N_25611);
xnor U26044 (N_26044,N_25489,N_25352);
and U26045 (N_26045,N_25857,N_25275);
nor U26046 (N_26046,N_25251,N_25757);
and U26047 (N_26047,N_25454,N_25960);
xor U26048 (N_26048,N_25334,N_25533);
and U26049 (N_26049,N_25684,N_25467);
and U26050 (N_26050,N_25003,N_25971);
or U26051 (N_26051,N_25371,N_25812);
and U26052 (N_26052,N_25427,N_25988);
xnor U26053 (N_26053,N_25581,N_25043);
or U26054 (N_26054,N_25140,N_25188);
and U26055 (N_26055,N_25420,N_25890);
xnor U26056 (N_26056,N_25722,N_25556);
nand U26057 (N_26057,N_25085,N_25555);
nand U26058 (N_26058,N_25958,N_25468);
nor U26059 (N_26059,N_25970,N_25451);
and U26060 (N_26060,N_25766,N_25823);
and U26061 (N_26061,N_25250,N_25665);
nand U26062 (N_26062,N_25037,N_25137);
and U26063 (N_26063,N_25558,N_25784);
xnor U26064 (N_26064,N_25416,N_25961);
xor U26065 (N_26065,N_25906,N_25778);
nand U26066 (N_26066,N_25601,N_25234);
and U26067 (N_26067,N_25567,N_25398);
and U26068 (N_26068,N_25606,N_25696);
or U26069 (N_26069,N_25820,N_25987);
nand U26070 (N_26070,N_25797,N_25641);
nand U26071 (N_26071,N_25830,N_25701);
xor U26072 (N_26072,N_25806,N_25072);
and U26073 (N_26073,N_25032,N_25298);
and U26074 (N_26074,N_25130,N_25864);
nand U26075 (N_26075,N_25540,N_25097);
and U26076 (N_26076,N_25674,N_25619);
nor U26077 (N_26077,N_25691,N_25680);
nand U26078 (N_26078,N_25947,N_25123);
nor U26079 (N_26079,N_25969,N_25055);
xor U26080 (N_26080,N_25210,N_25514);
and U26081 (N_26081,N_25139,N_25613);
xnor U26082 (N_26082,N_25711,N_25186);
nor U26083 (N_26083,N_25790,N_25980);
nand U26084 (N_26084,N_25209,N_25719);
or U26085 (N_26085,N_25979,N_25084);
and U26086 (N_26086,N_25788,N_25171);
xor U26087 (N_26087,N_25340,N_25973);
nand U26088 (N_26088,N_25480,N_25972);
and U26089 (N_26089,N_25916,N_25984);
and U26090 (N_26090,N_25804,N_25433);
xnor U26091 (N_26091,N_25900,N_25821);
and U26092 (N_26092,N_25153,N_25432);
nand U26093 (N_26093,N_25326,N_25749);
nand U26094 (N_26094,N_25093,N_25783);
and U26095 (N_26095,N_25206,N_25460);
and U26096 (N_26096,N_25396,N_25905);
xnor U26097 (N_26097,N_25443,N_25932);
nor U26098 (N_26098,N_25714,N_25437);
nor U26099 (N_26099,N_25729,N_25623);
or U26100 (N_26100,N_25029,N_25796);
nand U26101 (N_26101,N_25394,N_25964);
nand U26102 (N_26102,N_25798,N_25730);
xor U26103 (N_26103,N_25047,N_25716);
and U26104 (N_26104,N_25103,N_25678);
nand U26105 (N_26105,N_25828,N_25270);
nand U26106 (N_26106,N_25951,N_25535);
nor U26107 (N_26107,N_25228,N_25803);
nor U26108 (N_26108,N_25541,N_25509);
xnor U26109 (N_26109,N_25813,N_25944);
xor U26110 (N_26110,N_25070,N_25384);
or U26111 (N_26111,N_25095,N_25837);
xor U26112 (N_26112,N_25195,N_25452);
xnor U26113 (N_26113,N_25727,N_25201);
nor U26114 (N_26114,N_25814,N_25491);
nor U26115 (N_26115,N_25762,N_25710);
or U26116 (N_26116,N_25238,N_25505);
nor U26117 (N_26117,N_25955,N_25832);
or U26118 (N_26118,N_25200,N_25156);
or U26119 (N_26119,N_25386,N_25498);
nand U26120 (N_26120,N_25351,N_25078);
nand U26121 (N_26121,N_25404,N_25204);
xnor U26122 (N_26122,N_25073,N_25747);
nor U26123 (N_26123,N_25397,N_25708);
nand U26124 (N_26124,N_25912,N_25527);
or U26125 (N_26125,N_25743,N_25733);
nand U26126 (N_26126,N_25728,N_25579);
nor U26127 (N_26127,N_25317,N_25364);
nand U26128 (N_26128,N_25939,N_25190);
or U26129 (N_26129,N_25380,N_25212);
nand U26130 (N_26130,N_25848,N_25005);
or U26131 (N_26131,N_25021,N_25440);
nand U26132 (N_26132,N_25224,N_25240);
nand U26133 (N_26133,N_25996,N_25931);
nor U26134 (N_26134,N_25339,N_25297);
nor U26135 (N_26135,N_25356,N_25030);
nor U26136 (N_26136,N_25415,N_25622);
or U26137 (N_26137,N_25408,N_25328);
and U26138 (N_26138,N_25750,N_25576);
nand U26139 (N_26139,N_25127,N_25582);
nand U26140 (N_26140,N_25385,N_25512);
xnor U26141 (N_26141,N_25649,N_25162);
xor U26142 (N_26142,N_25508,N_25539);
nor U26143 (N_26143,N_25921,N_25954);
nand U26144 (N_26144,N_25281,N_25896);
and U26145 (N_26145,N_25941,N_25700);
and U26146 (N_26146,N_25161,N_25822);
xor U26147 (N_26147,N_25827,N_25523);
or U26148 (N_26148,N_25406,N_25736);
or U26149 (N_26149,N_25902,N_25319);
or U26150 (N_26150,N_25718,N_25235);
xnor U26151 (N_26151,N_25926,N_25911);
nand U26152 (N_26152,N_25052,N_25259);
or U26153 (N_26153,N_25782,N_25192);
nor U26154 (N_26154,N_25838,N_25843);
nand U26155 (N_26155,N_25273,N_25348);
xor U26156 (N_26156,N_25688,N_25354);
nand U26157 (N_26157,N_25746,N_25325);
xor U26158 (N_26158,N_25287,N_25564);
nor U26159 (N_26159,N_25868,N_25017);
nor U26160 (N_26160,N_25545,N_25342);
nand U26161 (N_26161,N_25963,N_25125);
xor U26162 (N_26162,N_25640,N_25484);
xor U26163 (N_26163,N_25652,N_25651);
xor U26164 (N_26164,N_25933,N_25436);
nor U26165 (N_26165,N_25575,N_25891);
and U26166 (N_26166,N_25143,N_25647);
xnor U26167 (N_26167,N_25537,N_25522);
nor U26168 (N_26168,N_25202,N_25760);
xnor U26169 (N_26169,N_25272,N_25934);
xnor U26170 (N_26170,N_25849,N_25293);
and U26171 (N_26171,N_25840,N_25337);
nor U26172 (N_26172,N_25618,N_25424);
or U26173 (N_26173,N_25310,N_25874);
and U26174 (N_26174,N_25280,N_25059);
xor U26175 (N_26175,N_25586,N_25096);
xor U26176 (N_26176,N_25182,N_25080);
nand U26177 (N_26177,N_25616,N_25442);
nand U26178 (N_26178,N_25949,N_25879);
or U26179 (N_26179,N_25341,N_25359);
or U26180 (N_26180,N_25758,N_25529);
nand U26181 (N_26181,N_25063,N_25568);
nand U26182 (N_26182,N_25101,N_25637);
nand U26183 (N_26183,N_25759,N_25115);
xnor U26184 (N_26184,N_25006,N_25283);
nor U26185 (N_26185,N_25501,N_25146);
xnor U26186 (N_26186,N_25267,N_25448);
nand U26187 (N_26187,N_25867,N_25455);
nand U26188 (N_26188,N_25603,N_25662);
xnor U26189 (N_26189,N_25860,N_25069);
nor U26190 (N_26190,N_25461,N_25439);
nor U26191 (N_26191,N_25819,N_25605);
and U26192 (N_26192,N_25071,N_25196);
nand U26193 (N_26193,N_25626,N_25299);
nor U26194 (N_26194,N_25612,N_25062);
and U26195 (N_26195,N_25692,N_25044);
and U26196 (N_26196,N_25253,N_25744);
or U26197 (N_26197,N_25686,N_25227);
nor U26198 (N_26198,N_25098,N_25671);
and U26199 (N_26199,N_25742,N_25707);
xor U26200 (N_26200,N_25308,N_25469);
xor U26201 (N_26201,N_25922,N_25051);
xor U26202 (N_26202,N_25390,N_25347);
nor U26203 (N_26203,N_25572,N_25165);
nor U26204 (N_26204,N_25459,N_25191);
and U26205 (N_26205,N_25229,N_25914);
and U26206 (N_26206,N_25734,N_25316);
nand U26207 (N_26207,N_25596,N_25144);
nor U26208 (N_26208,N_25061,N_25343);
or U26209 (N_26209,N_25669,N_25366);
or U26210 (N_26210,N_25952,N_25119);
nor U26211 (N_26211,N_25252,N_25774);
xor U26212 (N_26212,N_25549,N_25092);
nor U26213 (N_26213,N_25754,N_25738);
or U26214 (N_26214,N_25511,N_25330);
nand U26215 (N_26215,N_25001,N_25172);
nor U26216 (N_26216,N_25243,N_25014);
or U26217 (N_26217,N_25135,N_25079);
and U26218 (N_26218,N_25026,N_25391);
xnor U26219 (N_26219,N_25482,N_25740);
xor U26220 (N_26220,N_25181,N_25040);
and U26221 (N_26221,N_25008,N_25672);
and U26222 (N_26222,N_25777,N_25429);
xor U26223 (N_26223,N_25199,N_25271);
nand U26224 (N_26224,N_25887,N_25091);
nor U26225 (N_26225,N_25050,N_25817);
nand U26226 (N_26226,N_25205,N_25081);
nand U26227 (N_26227,N_25574,N_25120);
nor U26228 (N_26228,N_25490,N_25776);
xnor U26229 (N_26229,N_25417,N_25917);
and U26230 (N_26230,N_25910,N_25479);
and U26231 (N_26231,N_25739,N_25519);
xnor U26232 (N_26232,N_25741,N_25155);
xnor U26233 (N_26233,N_25290,N_25681);
nand U26234 (N_26234,N_25590,N_25054);
or U26235 (N_26235,N_25907,N_25076);
xor U26236 (N_26236,N_25862,N_25411);
xnor U26237 (N_26237,N_25634,N_25923);
xnor U26238 (N_26238,N_25633,N_25002);
and U26239 (N_26239,N_25465,N_25918);
nor U26240 (N_26240,N_25876,N_25151);
nor U26241 (N_26241,N_25336,N_25869);
nand U26242 (N_26242,N_25977,N_25363);
nor U26243 (N_26243,N_25222,N_25913);
nor U26244 (N_26244,N_25690,N_25481);
and U26245 (N_26245,N_25213,N_25134);
nor U26246 (N_26246,N_25068,N_25811);
or U26247 (N_26247,N_25245,N_25056);
or U26248 (N_26248,N_25112,N_25329);
nand U26249 (N_26249,N_25495,N_25793);
nand U26250 (N_26250,N_25886,N_25013);
xnor U26251 (N_26251,N_25983,N_25632);
nand U26252 (N_26252,N_25183,N_25769);
nor U26253 (N_26253,N_25654,N_25882);
nand U26254 (N_26254,N_25500,N_25520);
and U26255 (N_26255,N_25808,N_25990);
xnor U26256 (N_26256,N_25421,N_25561);
and U26257 (N_26257,N_25395,N_25239);
nor U26258 (N_26258,N_25735,N_25975);
or U26259 (N_26259,N_25219,N_25792);
and U26260 (N_26260,N_25577,N_25851);
xor U26261 (N_26261,N_25075,N_25262);
or U26262 (N_26262,N_25434,N_25554);
xor U26263 (N_26263,N_25198,N_25620);
nand U26264 (N_26264,N_25189,N_25945);
or U26265 (N_26265,N_25254,N_25528);
xor U26266 (N_26266,N_25349,N_25493);
nor U26267 (N_26267,N_25464,N_25012);
and U26268 (N_26268,N_25940,N_25318);
nor U26269 (N_26269,N_25203,N_25682);
nor U26270 (N_26270,N_25230,N_25908);
or U26271 (N_26271,N_25033,N_25425);
or U26272 (N_26272,N_25122,N_25375);
nor U26273 (N_26273,N_25478,N_25129);
xor U26274 (N_26274,N_25751,N_25124);
nor U26275 (N_26275,N_25038,N_25638);
or U26276 (N_26276,N_25810,N_25631);
or U26277 (N_26277,N_25463,N_25284);
nand U26278 (N_26278,N_25957,N_25242);
nand U26279 (N_26279,N_25041,N_25789);
nor U26280 (N_26280,N_25657,N_25315);
and U26281 (N_26281,N_25748,N_25534);
and U26282 (N_26282,N_25609,N_25358);
xnor U26283 (N_26283,N_25116,N_25389);
and U26284 (N_26284,N_25000,N_25953);
xnor U26285 (N_26285,N_25833,N_25407);
nand U26286 (N_26286,N_25114,N_25946);
nor U26287 (N_26287,N_25158,N_25683);
or U26288 (N_26288,N_25121,N_25303);
nand U26289 (N_26289,N_25901,N_25510);
and U26290 (N_26290,N_25180,N_25627);
nor U26291 (N_26291,N_25430,N_25850);
nand U26292 (N_26292,N_25989,N_25834);
and U26293 (N_26293,N_25015,N_25768);
or U26294 (N_26294,N_25207,N_25445);
nand U26295 (N_26295,N_25694,N_25536);
nand U26296 (N_26296,N_25755,N_25550);
nand U26297 (N_26297,N_25392,N_25009);
nand U26298 (N_26298,N_25110,N_25592);
or U26299 (N_26299,N_25246,N_25723);
or U26300 (N_26300,N_25898,N_25553);
nand U26301 (N_26301,N_25884,N_25625);
and U26302 (N_26302,N_25094,N_25233);
xnor U26303 (N_26303,N_25285,N_25878);
or U26304 (N_26304,N_25438,N_25526);
xor U26305 (N_26305,N_25909,N_25402);
nand U26306 (N_26306,N_25082,N_25053);
or U26307 (N_26307,N_25257,N_25530);
or U26308 (N_26308,N_25466,N_25525);
xor U26309 (N_26309,N_25327,N_25816);
nand U26310 (N_26310,N_25598,N_25724);
and U26311 (N_26311,N_25551,N_25147);
or U26312 (N_26312,N_25138,N_25695);
nor U26313 (N_26313,N_25089,N_25064);
or U26314 (N_26314,N_25100,N_25169);
xor U26315 (N_26315,N_25773,N_25565);
and U26316 (N_26316,N_25801,N_25036);
or U26317 (N_26317,N_25899,N_25313);
nor U26318 (N_26318,N_25865,N_25231);
xnor U26319 (N_26319,N_25462,N_25458);
xnor U26320 (N_26320,N_25184,N_25516);
or U26321 (N_26321,N_25639,N_25142);
nor U26322 (N_26322,N_25381,N_25604);
and U26323 (N_26323,N_25978,N_25943);
and U26324 (N_26324,N_25787,N_25185);
xnor U26325 (N_26325,N_25761,N_25950);
or U26326 (N_26326,N_25393,N_25109);
xor U26327 (N_26327,N_25721,N_25515);
nand U26328 (N_26328,N_25175,N_25705);
nor U26329 (N_26329,N_25046,N_25875);
nand U26330 (N_26330,N_25217,N_25497);
and U26331 (N_26331,N_25767,N_25966);
nand U26332 (N_26332,N_25117,N_25145);
nand U26333 (N_26333,N_25457,N_25818);
and U26334 (N_26334,N_25852,N_25058);
nand U26335 (N_26335,N_25765,N_25935);
xnor U26336 (N_26336,N_25300,N_25331);
nand U26337 (N_26337,N_25992,N_25277);
and U26338 (N_26338,N_25544,N_25794);
and U26339 (N_26339,N_25675,N_25644);
and U26340 (N_26340,N_25924,N_25566);
xor U26341 (N_26341,N_25382,N_25255);
and U26342 (N_26342,N_25004,N_25413);
or U26343 (N_26343,N_25706,N_25635);
and U26344 (N_26344,N_25133,N_25306);
nor U26345 (N_26345,N_25858,N_25915);
or U26346 (N_26346,N_25154,N_25636);
and U26347 (N_26347,N_25888,N_25108);
and U26348 (N_26348,N_25338,N_25236);
xor U26349 (N_26349,N_25016,N_25597);
or U26350 (N_26350,N_25712,N_25226);
or U26351 (N_26351,N_25225,N_25563);
nand U26352 (N_26352,N_25494,N_25745);
nand U26353 (N_26353,N_25981,N_25320);
and U26354 (N_26354,N_25074,N_25506);
xnor U26355 (N_26355,N_25295,N_25401);
xnor U26356 (N_26356,N_25786,N_25894);
nor U26357 (N_26357,N_25679,N_25099);
or U26358 (N_26358,N_25148,N_25086);
or U26359 (N_26359,N_25713,N_25795);
nor U26360 (N_26360,N_25919,N_25126);
and U26361 (N_26361,N_25580,N_25502);
or U26362 (N_26362,N_25815,N_25274);
or U26363 (N_26363,N_25412,N_25847);
or U26364 (N_26364,N_25621,N_25067);
nor U26365 (N_26365,N_25368,N_25211);
nor U26366 (N_26366,N_25825,N_25292);
xor U26367 (N_26367,N_25756,N_25560);
nand U26368 (N_26368,N_25312,N_25282);
or U26369 (N_26369,N_25664,N_25193);
xor U26370 (N_26370,N_25007,N_25335);
or U26371 (N_26371,N_25278,N_25607);
nand U26372 (N_26372,N_25309,N_25893);
nor U26373 (N_26373,N_25057,N_25324);
and U26374 (N_26374,N_25507,N_25699);
or U26375 (N_26375,N_25296,N_25314);
and U26376 (N_26376,N_25781,N_25150);
nand U26377 (N_26377,N_25426,N_25853);
nand U26378 (N_26378,N_25697,N_25223);
nand U26379 (N_26379,N_25503,N_25232);
and U26380 (N_26380,N_25885,N_25387);
nor U26381 (N_26381,N_25800,N_25141);
nand U26382 (N_26382,N_25023,N_25702);
or U26383 (N_26383,N_25400,N_25925);
nor U26384 (N_26384,N_25999,N_25608);
xor U26385 (N_26385,N_25881,N_25132);
and U26386 (N_26386,N_25471,N_25521);
and U26387 (N_26387,N_25357,N_25027);
and U26388 (N_26388,N_25446,N_25546);
xor U26389 (N_26389,N_25492,N_25174);
and U26390 (N_26390,N_25304,N_25302);
nor U26391 (N_26391,N_25360,N_25163);
nand U26392 (N_26392,N_25709,N_25976);
xor U26393 (N_26393,N_25031,N_25286);
xnor U26394 (N_26394,N_25345,N_25863);
or U26395 (N_26395,N_25584,N_25011);
or U26396 (N_26396,N_25562,N_25383);
and U26397 (N_26397,N_25570,N_25373);
nand U26398 (N_26398,N_25483,N_25965);
xnor U26399 (N_26399,N_25221,N_25895);
xnor U26400 (N_26400,N_25920,N_25414);
or U26401 (N_26401,N_25247,N_25967);
and U26402 (N_26402,N_25159,N_25379);
and U26403 (N_26403,N_25104,N_25845);
nor U26404 (N_26404,N_25720,N_25369);
nor U26405 (N_26405,N_25176,N_25450);
nor U26406 (N_26406,N_25410,N_25477);
xnor U26407 (N_26407,N_25587,N_25128);
nand U26408 (N_26408,N_25431,N_25422);
xor U26409 (N_26409,N_25024,N_25531);
and U26410 (N_26410,N_25615,N_25666);
nand U26411 (N_26411,N_25441,N_25048);
nand U26412 (N_26412,N_25805,N_25214);
nand U26413 (N_26413,N_25841,N_25880);
xor U26414 (N_26414,N_25872,N_25107);
nor U26415 (N_26415,N_25197,N_25367);
or U26416 (N_26416,N_25861,N_25157);
and U26417 (N_26417,N_25645,N_25168);
xor U26418 (N_26418,N_25517,N_25218);
or U26419 (N_26419,N_25668,N_25532);
or U26420 (N_26420,N_25543,N_25959);
nor U26421 (N_26421,N_25986,N_25780);
xor U26422 (N_26422,N_25065,N_25301);
nand U26423 (N_26423,N_25170,N_25083);
and U26424 (N_26424,N_25591,N_25937);
or U26425 (N_26425,N_25661,N_25475);
xnor U26426 (N_26426,N_25276,N_25474);
xnor U26427 (N_26427,N_25859,N_25929);
nand U26428 (N_26428,N_25405,N_25548);
or U26429 (N_26429,N_25269,N_25660);
and U26430 (N_26430,N_25216,N_25593);
and U26431 (N_26431,N_25444,N_25585);
and U26432 (N_26432,N_25763,N_25496);
xnor U26433 (N_26433,N_25985,N_25249);
xnor U26434 (N_26434,N_25677,N_25693);
and U26435 (N_26435,N_25418,N_25854);
or U26436 (N_26436,N_25152,N_25703);
nand U26437 (N_26437,N_25323,N_25764);
or U26438 (N_26438,N_25809,N_25903);
xnor U26439 (N_26439,N_25687,N_25419);
xor U26440 (N_26440,N_25968,N_25049);
and U26441 (N_26441,N_25962,N_25866);
nor U26442 (N_26442,N_25717,N_25350);
and U26443 (N_26443,N_25629,N_25485);
and U26444 (N_26444,N_25279,N_25077);
nand U26445 (N_26445,N_25839,N_25538);
or U26446 (N_26446,N_25956,N_25294);
or U26447 (N_26447,N_25435,N_25039);
or U26448 (N_26448,N_25028,N_25265);
xor U26449 (N_26449,N_25753,N_25388);
nor U26450 (N_26450,N_25927,N_25428);
nand U26451 (N_26451,N_25160,N_25547);
or U26452 (N_26452,N_25889,N_25374);
nor U26453 (N_26453,N_25569,N_25042);
xor U26454 (N_26454,N_25087,N_25600);
or U26455 (N_26455,N_25344,N_25307);
nor U26456 (N_26456,N_25361,N_25470);
nand U26457 (N_26457,N_25372,N_25589);
nand U26458 (N_26458,N_25578,N_25725);
xnor U26459 (N_26459,N_25237,N_25731);
xnor U26460 (N_26460,N_25173,N_25595);
or U26461 (N_26461,N_25676,N_25685);
nor U26462 (N_26462,N_25883,N_25456);
and U26463 (N_26463,N_25936,N_25010);
and U26464 (N_26464,N_25610,N_25557);
xor U26465 (N_26465,N_25663,N_25877);
xnor U26466 (N_26466,N_25715,N_25542);
nand U26467 (N_26467,N_25513,N_25377);
xnor U26468 (N_26468,N_25775,N_25321);
or U26469 (N_26469,N_25588,N_25791);
nor U26470 (N_26470,N_25518,N_25289);
nor U26471 (N_26471,N_25177,N_25667);
nor U26472 (N_26472,N_25447,N_25376);
or U26473 (N_26473,N_25802,N_25835);
and U26474 (N_26474,N_25322,N_25594);
or U26475 (N_26475,N_25504,N_25149);
or U26476 (N_26476,N_25248,N_25018);
xor U26477 (N_26477,N_25305,N_25583);
nand U26478 (N_26478,N_25982,N_25938);
nand U26479 (N_26479,N_25365,N_25892);
or U26480 (N_26480,N_25167,N_25263);
or U26481 (N_26481,N_25904,N_25179);
or U26482 (N_26482,N_25333,N_25332);
or U26483 (N_26483,N_25650,N_25704);
nor U26484 (N_26484,N_25034,N_25842);
nor U26485 (N_26485,N_25930,N_25268);
and U26486 (N_26486,N_25658,N_25244);
xnor U26487 (N_26487,N_25770,N_25045);
nand U26488 (N_26488,N_25614,N_25353);
xnor U26489 (N_26489,N_25166,N_25291);
nand U26490 (N_26490,N_25573,N_25829);
nand U26491 (N_26491,N_25266,N_25643);
or U26492 (N_26492,N_25215,N_25524);
nand U26493 (N_26493,N_25552,N_25659);
nand U26494 (N_26494,N_25423,N_25642);
or U26495 (N_26495,N_25131,N_25630);
xor U26496 (N_26496,N_25022,N_25942);
and U26497 (N_26497,N_25178,N_25771);
and U26498 (N_26498,N_25220,N_25066);
or U26499 (N_26499,N_25779,N_25974);
nand U26500 (N_26500,N_25890,N_25435);
xor U26501 (N_26501,N_25513,N_25168);
nor U26502 (N_26502,N_25219,N_25273);
or U26503 (N_26503,N_25059,N_25796);
nand U26504 (N_26504,N_25994,N_25078);
nor U26505 (N_26505,N_25142,N_25274);
or U26506 (N_26506,N_25858,N_25402);
xor U26507 (N_26507,N_25034,N_25399);
and U26508 (N_26508,N_25562,N_25584);
and U26509 (N_26509,N_25977,N_25259);
and U26510 (N_26510,N_25325,N_25639);
or U26511 (N_26511,N_25242,N_25758);
xnor U26512 (N_26512,N_25156,N_25491);
nand U26513 (N_26513,N_25165,N_25521);
nand U26514 (N_26514,N_25568,N_25624);
xnor U26515 (N_26515,N_25029,N_25825);
nor U26516 (N_26516,N_25570,N_25316);
xnor U26517 (N_26517,N_25905,N_25260);
xor U26518 (N_26518,N_25833,N_25351);
or U26519 (N_26519,N_25090,N_25118);
nand U26520 (N_26520,N_25307,N_25406);
or U26521 (N_26521,N_25154,N_25025);
and U26522 (N_26522,N_25081,N_25678);
nor U26523 (N_26523,N_25858,N_25772);
and U26524 (N_26524,N_25875,N_25424);
nand U26525 (N_26525,N_25913,N_25168);
and U26526 (N_26526,N_25281,N_25892);
nor U26527 (N_26527,N_25078,N_25108);
and U26528 (N_26528,N_25692,N_25728);
nor U26529 (N_26529,N_25165,N_25890);
nor U26530 (N_26530,N_25462,N_25656);
or U26531 (N_26531,N_25984,N_25636);
nand U26532 (N_26532,N_25804,N_25979);
xnor U26533 (N_26533,N_25476,N_25257);
nand U26534 (N_26534,N_25427,N_25425);
xnor U26535 (N_26535,N_25110,N_25779);
and U26536 (N_26536,N_25278,N_25526);
or U26537 (N_26537,N_25010,N_25793);
nand U26538 (N_26538,N_25724,N_25291);
and U26539 (N_26539,N_25943,N_25204);
nor U26540 (N_26540,N_25655,N_25641);
nor U26541 (N_26541,N_25225,N_25024);
and U26542 (N_26542,N_25250,N_25402);
and U26543 (N_26543,N_25774,N_25983);
or U26544 (N_26544,N_25251,N_25387);
nand U26545 (N_26545,N_25269,N_25697);
nand U26546 (N_26546,N_25777,N_25768);
nor U26547 (N_26547,N_25211,N_25407);
xnor U26548 (N_26548,N_25114,N_25453);
nand U26549 (N_26549,N_25396,N_25716);
xor U26550 (N_26550,N_25357,N_25005);
xnor U26551 (N_26551,N_25813,N_25014);
nor U26552 (N_26552,N_25262,N_25404);
nor U26553 (N_26553,N_25047,N_25066);
or U26554 (N_26554,N_25205,N_25794);
nand U26555 (N_26555,N_25486,N_25085);
or U26556 (N_26556,N_25829,N_25878);
xnor U26557 (N_26557,N_25756,N_25022);
xor U26558 (N_26558,N_25124,N_25075);
or U26559 (N_26559,N_25364,N_25188);
nand U26560 (N_26560,N_25681,N_25871);
nand U26561 (N_26561,N_25450,N_25546);
nand U26562 (N_26562,N_25071,N_25645);
nor U26563 (N_26563,N_25182,N_25308);
and U26564 (N_26564,N_25186,N_25405);
xnor U26565 (N_26565,N_25750,N_25948);
nor U26566 (N_26566,N_25292,N_25817);
nor U26567 (N_26567,N_25860,N_25663);
or U26568 (N_26568,N_25755,N_25713);
xnor U26569 (N_26569,N_25775,N_25066);
and U26570 (N_26570,N_25891,N_25144);
and U26571 (N_26571,N_25038,N_25560);
and U26572 (N_26572,N_25908,N_25319);
xor U26573 (N_26573,N_25620,N_25594);
or U26574 (N_26574,N_25462,N_25366);
and U26575 (N_26575,N_25267,N_25069);
and U26576 (N_26576,N_25318,N_25210);
or U26577 (N_26577,N_25877,N_25519);
nand U26578 (N_26578,N_25762,N_25883);
xnor U26579 (N_26579,N_25266,N_25619);
xnor U26580 (N_26580,N_25376,N_25081);
and U26581 (N_26581,N_25481,N_25156);
xor U26582 (N_26582,N_25191,N_25171);
xnor U26583 (N_26583,N_25224,N_25730);
nor U26584 (N_26584,N_25339,N_25456);
nor U26585 (N_26585,N_25711,N_25648);
nor U26586 (N_26586,N_25313,N_25871);
xnor U26587 (N_26587,N_25107,N_25992);
nand U26588 (N_26588,N_25895,N_25328);
and U26589 (N_26589,N_25475,N_25285);
or U26590 (N_26590,N_25427,N_25517);
xnor U26591 (N_26591,N_25774,N_25919);
and U26592 (N_26592,N_25266,N_25091);
and U26593 (N_26593,N_25182,N_25913);
or U26594 (N_26594,N_25328,N_25392);
or U26595 (N_26595,N_25759,N_25510);
and U26596 (N_26596,N_25227,N_25013);
nor U26597 (N_26597,N_25836,N_25534);
xnor U26598 (N_26598,N_25715,N_25485);
nor U26599 (N_26599,N_25193,N_25454);
nand U26600 (N_26600,N_25768,N_25614);
nand U26601 (N_26601,N_25485,N_25875);
xnor U26602 (N_26602,N_25972,N_25299);
nand U26603 (N_26603,N_25065,N_25189);
nor U26604 (N_26604,N_25932,N_25507);
nand U26605 (N_26605,N_25524,N_25171);
nor U26606 (N_26606,N_25044,N_25637);
xnor U26607 (N_26607,N_25352,N_25865);
or U26608 (N_26608,N_25149,N_25691);
nor U26609 (N_26609,N_25265,N_25799);
nor U26610 (N_26610,N_25723,N_25227);
or U26611 (N_26611,N_25927,N_25338);
nor U26612 (N_26612,N_25086,N_25760);
or U26613 (N_26613,N_25910,N_25723);
xor U26614 (N_26614,N_25069,N_25993);
and U26615 (N_26615,N_25265,N_25001);
and U26616 (N_26616,N_25750,N_25419);
xor U26617 (N_26617,N_25384,N_25036);
nor U26618 (N_26618,N_25084,N_25082);
or U26619 (N_26619,N_25166,N_25036);
xor U26620 (N_26620,N_25730,N_25029);
and U26621 (N_26621,N_25080,N_25676);
and U26622 (N_26622,N_25734,N_25003);
nor U26623 (N_26623,N_25020,N_25449);
nor U26624 (N_26624,N_25526,N_25643);
nand U26625 (N_26625,N_25756,N_25459);
nand U26626 (N_26626,N_25036,N_25463);
or U26627 (N_26627,N_25730,N_25067);
nor U26628 (N_26628,N_25338,N_25300);
and U26629 (N_26629,N_25859,N_25954);
nor U26630 (N_26630,N_25450,N_25772);
and U26631 (N_26631,N_25186,N_25037);
nor U26632 (N_26632,N_25769,N_25531);
xnor U26633 (N_26633,N_25821,N_25954);
nand U26634 (N_26634,N_25685,N_25119);
and U26635 (N_26635,N_25740,N_25874);
nand U26636 (N_26636,N_25024,N_25572);
nand U26637 (N_26637,N_25945,N_25808);
nand U26638 (N_26638,N_25872,N_25704);
nor U26639 (N_26639,N_25808,N_25166);
nand U26640 (N_26640,N_25444,N_25753);
nor U26641 (N_26641,N_25425,N_25113);
nor U26642 (N_26642,N_25343,N_25008);
or U26643 (N_26643,N_25905,N_25156);
xor U26644 (N_26644,N_25264,N_25818);
nand U26645 (N_26645,N_25092,N_25969);
xnor U26646 (N_26646,N_25519,N_25032);
xnor U26647 (N_26647,N_25633,N_25532);
xnor U26648 (N_26648,N_25937,N_25916);
and U26649 (N_26649,N_25718,N_25593);
and U26650 (N_26650,N_25646,N_25948);
and U26651 (N_26651,N_25219,N_25649);
or U26652 (N_26652,N_25607,N_25605);
and U26653 (N_26653,N_25686,N_25655);
and U26654 (N_26654,N_25995,N_25842);
xor U26655 (N_26655,N_25931,N_25025);
nand U26656 (N_26656,N_25257,N_25693);
or U26657 (N_26657,N_25841,N_25426);
xor U26658 (N_26658,N_25600,N_25730);
or U26659 (N_26659,N_25705,N_25634);
nand U26660 (N_26660,N_25506,N_25185);
xnor U26661 (N_26661,N_25654,N_25573);
nand U26662 (N_26662,N_25305,N_25174);
nor U26663 (N_26663,N_25300,N_25998);
nor U26664 (N_26664,N_25995,N_25282);
nand U26665 (N_26665,N_25424,N_25953);
nor U26666 (N_26666,N_25571,N_25671);
and U26667 (N_26667,N_25059,N_25585);
xor U26668 (N_26668,N_25301,N_25764);
nand U26669 (N_26669,N_25349,N_25045);
nor U26670 (N_26670,N_25747,N_25244);
nor U26671 (N_26671,N_25000,N_25758);
or U26672 (N_26672,N_25526,N_25749);
xor U26673 (N_26673,N_25067,N_25483);
nand U26674 (N_26674,N_25406,N_25035);
and U26675 (N_26675,N_25453,N_25004);
xor U26676 (N_26676,N_25827,N_25595);
xnor U26677 (N_26677,N_25055,N_25160);
and U26678 (N_26678,N_25956,N_25753);
or U26679 (N_26679,N_25007,N_25495);
xnor U26680 (N_26680,N_25951,N_25660);
nor U26681 (N_26681,N_25533,N_25627);
or U26682 (N_26682,N_25943,N_25564);
or U26683 (N_26683,N_25561,N_25743);
or U26684 (N_26684,N_25589,N_25744);
or U26685 (N_26685,N_25880,N_25095);
or U26686 (N_26686,N_25777,N_25174);
xor U26687 (N_26687,N_25143,N_25495);
and U26688 (N_26688,N_25634,N_25322);
and U26689 (N_26689,N_25030,N_25170);
nand U26690 (N_26690,N_25860,N_25697);
nor U26691 (N_26691,N_25305,N_25587);
and U26692 (N_26692,N_25943,N_25961);
and U26693 (N_26693,N_25584,N_25811);
nand U26694 (N_26694,N_25281,N_25584);
nand U26695 (N_26695,N_25503,N_25239);
and U26696 (N_26696,N_25304,N_25312);
or U26697 (N_26697,N_25586,N_25015);
xnor U26698 (N_26698,N_25727,N_25827);
or U26699 (N_26699,N_25256,N_25898);
nand U26700 (N_26700,N_25652,N_25083);
and U26701 (N_26701,N_25072,N_25103);
and U26702 (N_26702,N_25558,N_25246);
nor U26703 (N_26703,N_25289,N_25186);
nor U26704 (N_26704,N_25007,N_25546);
nand U26705 (N_26705,N_25121,N_25068);
xor U26706 (N_26706,N_25394,N_25004);
nor U26707 (N_26707,N_25778,N_25556);
or U26708 (N_26708,N_25460,N_25287);
xor U26709 (N_26709,N_25681,N_25845);
xor U26710 (N_26710,N_25570,N_25597);
xor U26711 (N_26711,N_25177,N_25734);
xor U26712 (N_26712,N_25485,N_25577);
and U26713 (N_26713,N_25238,N_25069);
xor U26714 (N_26714,N_25741,N_25989);
and U26715 (N_26715,N_25738,N_25911);
or U26716 (N_26716,N_25167,N_25885);
nand U26717 (N_26717,N_25430,N_25481);
nor U26718 (N_26718,N_25393,N_25223);
nor U26719 (N_26719,N_25419,N_25417);
nand U26720 (N_26720,N_25906,N_25612);
or U26721 (N_26721,N_25064,N_25402);
and U26722 (N_26722,N_25140,N_25297);
nand U26723 (N_26723,N_25073,N_25754);
nor U26724 (N_26724,N_25688,N_25314);
nor U26725 (N_26725,N_25240,N_25472);
nand U26726 (N_26726,N_25544,N_25784);
nand U26727 (N_26727,N_25530,N_25623);
and U26728 (N_26728,N_25971,N_25582);
and U26729 (N_26729,N_25978,N_25885);
nor U26730 (N_26730,N_25044,N_25985);
or U26731 (N_26731,N_25067,N_25512);
nand U26732 (N_26732,N_25865,N_25322);
xnor U26733 (N_26733,N_25585,N_25662);
xor U26734 (N_26734,N_25657,N_25408);
and U26735 (N_26735,N_25281,N_25009);
or U26736 (N_26736,N_25698,N_25821);
nand U26737 (N_26737,N_25994,N_25868);
or U26738 (N_26738,N_25891,N_25285);
nor U26739 (N_26739,N_25015,N_25648);
nor U26740 (N_26740,N_25494,N_25245);
xor U26741 (N_26741,N_25465,N_25291);
nor U26742 (N_26742,N_25437,N_25039);
nand U26743 (N_26743,N_25226,N_25429);
and U26744 (N_26744,N_25315,N_25463);
xor U26745 (N_26745,N_25415,N_25859);
xor U26746 (N_26746,N_25629,N_25800);
and U26747 (N_26747,N_25146,N_25268);
nand U26748 (N_26748,N_25847,N_25086);
nand U26749 (N_26749,N_25382,N_25005);
nor U26750 (N_26750,N_25532,N_25183);
xnor U26751 (N_26751,N_25025,N_25279);
or U26752 (N_26752,N_25037,N_25232);
nor U26753 (N_26753,N_25243,N_25090);
nand U26754 (N_26754,N_25850,N_25213);
xor U26755 (N_26755,N_25509,N_25815);
nand U26756 (N_26756,N_25644,N_25685);
xnor U26757 (N_26757,N_25005,N_25441);
and U26758 (N_26758,N_25445,N_25972);
and U26759 (N_26759,N_25510,N_25429);
or U26760 (N_26760,N_25489,N_25066);
nand U26761 (N_26761,N_25911,N_25045);
nand U26762 (N_26762,N_25656,N_25393);
nand U26763 (N_26763,N_25384,N_25637);
nand U26764 (N_26764,N_25140,N_25776);
nand U26765 (N_26765,N_25927,N_25166);
xor U26766 (N_26766,N_25399,N_25141);
nor U26767 (N_26767,N_25108,N_25291);
xnor U26768 (N_26768,N_25206,N_25911);
and U26769 (N_26769,N_25887,N_25950);
nor U26770 (N_26770,N_25941,N_25699);
xor U26771 (N_26771,N_25128,N_25847);
nand U26772 (N_26772,N_25441,N_25841);
nor U26773 (N_26773,N_25014,N_25239);
or U26774 (N_26774,N_25704,N_25253);
xnor U26775 (N_26775,N_25787,N_25356);
or U26776 (N_26776,N_25223,N_25899);
and U26777 (N_26777,N_25104,N_25656);
nor U26778 (N_26778,N_25401,N_25797);
and U26779 (N_26779,N_25025,N_25656);
xnor U26780 (N_26780,N_25825,N_25524);
or U26781 (N_26781,N_25143,N_25081);
nor U26782 (N_26782,N_25342,N_25478);
and U26783 (N_26783,N_25369,N_25479);
xor U26784 (N_26784,N_25923,N_25813);
or U26785 (N_26785,N_25957,N_25692);
xor U26786 (N_26786,N_25943,N_25703);
or U26787 (N_26787,N_25538,N_25558);
or U26788 (N_26788,N_25567,N_25634);
nor U26789 (N_26789,N_25103,N_25183);
nand U26790 (N_26790,N_25369,N_25970);
or U26791 (N_26791,N_25336,N_25875);
nand U26792 (N_26792,N_25309,N_25714);
or U26793 (N_26793,N_25042,N_25618);
nand U26794 (N_26794,N_25664,N_25061);
nor U26795 (N_26795,N_25658,N_25380);
nand U26796 (N_26796,N_25098,N_25174);
or U26797 (N_26797,N_25976,N_25544);
nand U26798 (N_26798,N_25099,N_25900);
and U26799 (N_26799,N_25550,N_25385);
nand U26800 (N_26800,N_25650,N_25713);
and U26801 (N_26801,N_25726,N_25139);
nand U26802 (N_26802,N_25558,N_25103);
or U26803 (N_26803,N_25615,N_25940);
or U26804 (N_26804,N_25610,N_25533);
nor U26805 (N_26805,N_25212,N_25459);
and U26806 (N_26806,N_25719,N_25612);
and U26807 (N_26807,N_25146,N_25656);
or U26808 (N_26808,N_25200,N_25865);
nand U26809 (N_26809,N_25811,N_25850);
nor U26810 (N_26810,N_25092,N_25519);
nand U26811 (N_26811,N_25543,N_25292);
xnor U26812 (N_26812,N_25966,N_25304);
nor U26813 (N_26813,N_25932,N_25577);
or U26814 (N_26814,N_25694,N_25268);
xor U26815 (N_26815,N_25253,N_25798);
and U26816 (N_26816,N_25501,N_25099);
nand U26817 (N_26817,N_25974,N_25245);
nand U26818 (N_26818,N_25917,N_25790);
xnor U26819 (N_26819,N_25487,N_25918);
or U26820 (N_26820,N_25343,N_25266);
and U26821 (N_26821,N_25223,N_25865);
or U26822 (N_26822,N_25189,N_25807);
or U26823 (N_26823,N_25785,N_25715);
and U26824 (N_26824,N_25364,N_25146);
or U26825 (N_26825,N_25135,N_25049);
nand U26826 (N_26826,N_25625,N_25190);
xor U26827 (N_26827,N_25682,N_25772);
and U26828 (N_26828,N_25183,N_25881);
nor U26829 (N_26829,N_25642,N_25867);
nand U26830 (N_26830,N_25906,N_25551);
nand U26831 (N_26831,N_25257,N_25826);
or U26832 (N_26832,N_25544,N_25021);
or U26833 (N_26833,N_25922,N_25936);
nand U26834 (N_26834,N_25147,N_25293);
xor U26835 (N_26835,N_25773,N_25697);
xnor U26836 (N_26836,N_25701,N_25906);
xnor U26837 (N_26837,N_25270,N_25383);
nor U26838 (N_26838,N_25809,N_25981);
or U26839 (N_26839,N_25627,N_25045);
or U26840 (N_26840,N_25249,N_25566);
nand U26841 (N_26841,N_25570,N_25351);
and U26842 (N_26842,N_25953,N_25786);
or U26843 (N_26843,N_25525,N_25247);
nand U26844 (N_26844,N_25621,N_25962);
xnor U26845 (N_26845,N_25989,N_25413);
nor U26846 (N_26846,N_25845,N_25742);
xnor U26847 (N_26847,N_25737,N_25535);
nor U26848 (N_26848,N_25389,N_25081);
and U26849 (N_26849,N_25998,N_25004);
or U26850 (N_26850,N_25575,N_25385);
and U26851 (N_26851,N_25624,N_25665);
nand U26852 (N_26852,N_25967,N_25172);
nor U26853 (N_26853,N_25504,N_25775);
nor U26854 (N_26854,N_25717,N_25979);
nor U26855 (N_26855,N_25553,N_25832);
nand U26856 (N_26856,N_25616,N_25262);
nand U26857 (N_26857,N_25500,N_25827);
xor U26858 (N_26858,N_25173,N_25351);
or U26859 (N_26859,N_25760,N_25479);
and U26860 (N_26860,N_25853,N_25111);
and U26861 (N_26861,N_25634,N_25280);
nor U26862 (N_26862,N_25997,N_25505);
xnor U26863 (N_26863,N_25817,N_25760);
and U26864 (N_26864,N_25941,N_25819);
nand U26865 (N_26865,N_25990,N_25838);
and U26866 (N_26866,N_25414,N_25694);
nor U26867 (N_26867,N_25193,N_25387);
nor U26868 (N_26868,N_25456,N_25057);
or U26869 (N_26869,N_25871,N_25480);
nand U26870 (N_26870,N_25320,N_25592);
nor U26871 (N_26871,N_25980,N_25865);
and U26872 (N_26872,N_25557,N_25924);
nor U26873 (N_26873,N_25144,N_25491);
or U26874 (N_26874,N_25801,N_25642);
nor U26875 (N_26875,N_25876,N_25291);
or U26876 (N_26876,N_25201,N_25465);
or U26877 (N_26877,N_25555,N_25407);
nor U26878 (N_26878,N_25011,N_25269);
xnor U26879 (N_26879,N_25222,N_25870);
and U26880 (N_26880,N_25105,N_25735);
or U26881 (N_26881,N_25773,N_25568);
nand U26882 (N_26882,N_25771,N_25828);
or U26883 (N_26883,N_25680,N_25233);
nand U26884 (N_26884,N_25357,N_25935);
or U26885 (N_26885,N_25311,N_25718);
xnor U26886 (N_26886,N_25808,N_25660);
nand U26887 (N_26887,N_25173,N_25271);
or U26888 (N_26888,N_25875,N_25719);
nand U26889 (N_26889,N_25623,N_25815);
or U26890 (N_26890,N_25360,N_25025);
or U26891 (N_26891,N_25029,N_25126);
xnor U26892 (N_26892,N_25711,N_25856);
nor U26893 (N_26893,N_25156,N_25612);
and U26894 (N_26894,N_25779,N_25058);
nand U26895 (N_26895,N_25969,N_25576);
xor U26896 (N_26896,N_25953,N_25883);
nor U26897 (N_26897,N_25468,N_25894);
nand U26898 (N_26898,N_25960,N_25041);
xnor U26899 (N_26899,N_25754,N_25839);
nand U26900 (N_26900,N_25173,N_25533);
nand U26901 (N_26901,N_25200,N_25716);
and U26902 (N_26902,N_25145,N_25072);
nor U26903 (N_26903,N_25738,N_25747);
xnor U26904 (N_26904,N_25381,N_25013);
and U26905 (N_26905,N_25862,N_25703);
nand U26906 (N_26906,N_25880,N_25795);
xor U26907 (N_26907,N_25321,N_25647);
xnor U26908 (N_26908,N_25966,N_25811);
nand U26909 (N_26909,N_25640,N_25741);
and U26910 (N_26910,N_25393,N_25697);
nand U26911 (N_26911,N_25897,N_25216);
xor U26912 (N_26912,N_25915,N_25873);
xnor U26913 (N_26913,N_25020,N_25510);
xnor U26914 (N_26914,N_25189,N_25719);
nand U26915 (N_26915,N_25918,N_25759);
xor U26916 (N_26916,N_25688,N_25507);
xor U26917 (N_26917,N_25959,N_25350);
and U26918 (N_26918,N_25846,N_25697);
and U26919 (N_26919,N_25091,N_25115);
or U26920 (N_26920,N_25397,N_25973);
and U26921 (N_26921,N_25941,N_25076);
nor U26922 (N_26922,N_25126,N_25156);
or U26923 (N_26923,N_25269,N_25938);
and U26924 (N_26924,N_25881,N_25485);
or U26925 (N_26925,N_25592,N_25647);
nor U26926 (N_26926,N_25226,N_25936);
xnor U26927 (N_26927,N_25428,N_25996);
or U26928 (N_26928,N_25765,N_25062);
xor U26929 (N_26929,N_25886,N_25772);
xor U26930 (N_26930,N_25296,N_25143);
nand U26931 (N_26931,N_25352,N_25311);
nor U26932 (N_26932,N_25928,N_25560);
or U26933 (N_26933,N_25536,N_25388);
xnor U26934 (N_26934,N_25921,N_25438);
nand U26935 (N_26935,N_25590,N_25211);
nor U26936 (N_26936,N_25750,N_25231);
nand U26937 (N_26937,N_25401,N_25081);
or U26938 (N_26938,N_25714,N_25203);
xnor U26939 (N_26939,N_25365,N_25233);
and U26940 (N_26940,N_25126,N_25271);
nor U26941 (N_26941,N_25912,N_25992);
nor U26942 (N_26942,N_25872,N_25284);
nor U26943 (N_26943,N_25923,N_25394);
and U26944 (N_26944,N_25029,N_25015);
or U26945 (N_26945,N_25025,N_25161);
xor U26946 (N_26946,N_25484,N_25473);
and U26947 (N_26947,N_25064,N_25855);
and U26948 (N_26948,N_25834,N_25502);
and U26949 (N_26949,N_25447,N_25750);
nor U26950 (N_26950,N_25945,N_25052);
xor U26951 (N_26951,N_25069,N_25823);
nand U26952 (N_26952,N_25002,N_25799);
xor U26953 (N_26953,N_25697,N_25214);
nand U26954 (N_26954,N_25689,N_25791);
and U26955 (N_26955,N_25619,N_25611);
or U26956 (N_26956,N_25089,N_25220);
xor U26957 (N_26957,N_25566,N_25938);
nor U26958 (N_26958,N_25100,N_25843);
or U26959 (N_26959,N_25672,N_25907);
nand U26960 (N_26960,N_25006,N_25735);
nor U26961 (N_26961,N_25011,N_25814);
nand U26962 (N_26962,N_25748,N_25792);
nor U26963 (N_26963,N_25468,N_25218);
xnor U26964 (N_26964,N_25280,N_25515);
and U26965 (N_26965,N_25253,N_25950);
nor U26966 (N_26966,N_25104,N_25542);
nor U26967 (N_26967,N_25001,N_25204);
or U26968 (N_26968,N_25385,N_25208);
and U26969 (N_26969,N_25698,N_25283);
xor U26970 (N_26970,N_25970,N_25868);
nor U26971 (N_26971,N_25647,N_25253);
nor U26972 (N_26972,N_25059,N_25518);
nand U26973 (N_26973,N_25195,N_25495);
xor U26974 (N_26974,N_25192,N_25138);
or U26975 (N_26975,N_25249,N_25707);
and U26976 (N_26976,N_25566,N_25808);
nor U26977 (N_26977,N_25465,N_25819);
nor U26978 (N_26978,N_25518,N_25756);
nor U26979 (N_26979,N_25263,N_25273);
xnor U26980 (N_26980,N_25546,N_25685);
nand U26981 (N_26981,N_25558,N_25147);
nand U26982 (N_26982,N_25196,N_25144);
nand U26983 (N_26983,N_25188,N_25525);
nand U26984 (N_26984,N_25274,N_25015);
or U26985 (N_26985,N_25273,N_25333);
or U26986 (N_26986,N_25840,N_25203);
or U26987 (N_26987,N_25147,N_25223);
xnor U26988 (N_26988,N_25772,N_25129);
nand U26989 (N_26989,N_25179,N_25572);
or U26990 (N_26990,N_25660,N_25988);
xor U26991 (N_26991,N_25615,N_25143);
and U26992 (N_26992,N_25599,N_25190);
xnor U26993 (N_26993,N_25992,N_25253);
nand U26994 (N_26994,N_25528,N_25411);
or U26995 (N_26995,N_25543,N_25592);
nor U26996 (N_26996,N_25084,N_25861);
xor U26997 (N_26997,N_25368,N_25655);
nand U26998 (N_26998,N_25330,N_25219);
or U26999 (N_26999,N_25663,N_25300);
and U27000 (N_27000,N_26058,N_26815);
nor U27001 (N_27001,N_26189,N_26575);
nand U27002 (N_27002,N_26187,N_26136);
and U27003 (N_27003,N_26203,N_26447);
nand U27004 (N_27004,N_26593,N_26452);
xnor U27005 (N_27005,N_26248,N_26569);
nand U27006 (N_27006,N_26534,N_26637);
or U27007 (N_27007,N_26926,N_26797);
nand U27008 (N_27008,N_26829,N_26555);
xor U27009 (N_27009,N_26836,N_26530);
nand U27010 (N_27010,N_26657,N_26953);
and U27011 (N_27011,N_26751,N_26473);
nor U27012 (N_27012,N_26289,N_26433);
or U27013 (N_27013,N_26604,N_26415);
nand U27014 (N_27014,N_26246,N_26319);
and U27015 (N_27015,N_26454,N_26388);
nor U27016 (N_27016,N_26052,N_26260);
nand U27017 (N_27017,N_26622,N_26726);
nand U27018 (N_27018,N_26700,N_26019);
nor U27019 (N_27019,N_26079,N_26191);
xor U27020 (N_27020,N_26123,N_26764);
nor U27021 (N_27021,N_26455,N_26412);
xor U27022 (N_27022,N_26725,N_26151);
or U27023 (N_27023,N_26065,N_26170);
or U27024 (N_27024,N_26262,N_26074);
or U27025 (N_27025,N_26892,N_26563);
xor U27026 (N_27026,N_26028,N_26711);
or U27027 (N_27027,N_26982,N_26313);
nand U27028 (N_27028,N_26630,N_26648);
and U27029 (N_27029,N_26460,N_26004);
nand U27030 (N_27030,N_26684,N_26862);
xnor U27031 (N_27031,N_26023,N_26215);
and U27032 (N_27032,N_26337,N_26472);
or U27033 (N_27033,N_26015,N_26972);
xor U27034 (N_27034,N_26933,N_26020);
or U27035 (N_27035,N_26470,N_26955);
and U27036 (N_27036,N_26961,N_26212);
nand U27037 (N_27037,N_26492,N_26226);
nor U27038 (N_27038,N_26837,N_26238);
nor U27039 (N_27039,N_26060,N_26995);
or U27040 (N_27040,N_26763,N_26293);
and U27041 (N_27041,N_26394,N_26169);
nor U27042 (N_27042,N_26744,N_26545);
xor U27043 (N_27043,N_26301,N_26948);
xor U27044 (N_27044,N_26649,N_26882);
xnor U27045 (N_27045,N_26780,N_26939);
xor U27046 (N_27046,N_26807,N_26574);
and U27047 (N_27047,N_26218,N_26273);
or U27048 (N_27048,N_26716,N_26167);
nand U27049 (N_27049,N_26639,N_26588);
xnor U27050 (N_27050,N_26309,N_26267);
and U27051 (N_27051,N_26853,N_26325);
xor U27052 (N_27052,N_26626,N_26214);
xor U27053 (N_27053,N_26655,N_26042);
and U27054 (N_27054,N_26731,N_26000);
xor U27055 (N_27055,N_26149,N_26565);
or U27056 (N_27056,N_26066,N_26476);
and U27057 (N_27057,N_26242,N_26265);
or U27058 (N_27058,N_26614,N_26976);
or U27059 (N_27059,N_26366,N_26934);
nor U27060 (N_27060,N_26664,N_26329);
or U27061 (N_27061,N_26101,N_26888);
xnor U27062 (N_27062,N_26268,N_26677);
nor U27063 (N_27063,N_26160,N_26596);
xor U27064 (N_27064,N_26606,N_26792);
nor U27065 (N_27065,N_26501,N_26782);
nand U27066 (N_27066,N_26498,N_26244);
and U27067 (N_27067,N_26016,N_26465);
or U27068 (N_27068,N_26463,N_26977);
nor U27069 (N_27069,N_26854,N_26391);
xor U27070 (N_27070,N_26735,N_26958);
xnor U27071 (N_27071,N_26537,N_26785);
xor U27072 (N_27072,N_26334,N_26485);
xnor U27073 (N_27073,N_26354,N_26222);
xnor U27074 (N_27074,N_26445,N_26627);
nand U27075 (N_27075,N_26789,N_26119);
nand U27076 (N_27076,N_26640,N_26316);
and U27077 (N_27077,N_26761,N_26475);
nor U27078 (N_27078,N_26283,N_26271);
and U27079 (N_27079,N_26063,N_26442);
nand U27080 (N_27080,N_26724,N_26570);
nand U27081 (N_27081,N_26287,N_26103);
xor U27082 (N_27082,N_26757,N_26154);
or U27083 (N_27083,N_26860,N_26227);
xor U27084 (N_27084,N_26512,N_26839);
and U27085 (N_27085,N_26910,N_26559);
nand U27086 (N_27086,N_26249,N_26487);
nor U27087 (N_27087,N_26183,N_26859);
nor U27088 (N_27088,N_26276,N_26033);
xor U27089 (N_27089,N_26440,N_26471);
nand U27090 (N_27090,N_26798,N_26762);
and U27091 (N_27091,N_26610,N_26687);
or U27092 (N_27092,N_26819,N_26461);
or U27093 (N_27093,N_26235,N_26903);
xor U27094 (N_27094,N_26421,N_26924);
nor U27095 (N_27095,N_26297,N_26175);
nand U27096 (N_27096,N_26011,N_26755);
nand U27097 (N_27097,N_26371,N_26038);
xor U27098 (N_27098,N_26355,N_26723);
and U27099 (N_27099,N_26230,N_26634);
nor U27100 (N_27100,N_26210,N_26091);
nor U27101 (N_27101,N_26304,N_26543);
and U27102 (N_27102,N_26095,N_26332);
or U27103 (N_27103,N_26223,N_26457);
nand U27104 (N_27104,N_26201,N_26007);
and U27105 (N_27105,N_26362,N_26040);
nor U27106 (N_27106,N_26318,N_26776);
and U27107 (N_27107,N_26282,N_26618);
and U27108 (N_27108,N_26696,N_26823);
and U27109 (N_27109,N_26324,N_26148);
nor U27110 (N_27110,N_26247,N_26450);
nor U27111 (N_27111,N_26535,N_26635);
nor U27112 (N_27112,N_26213,N_26712);
nand U27113 (N_27113,N_26335,N_26360);
and U27114 (N_27114,N_26959,N_26017);
nand U27115 (N_27115,N_26505,N_26872);
nor U27116 (N_27116,N_26707,N_26086);
nor U27117 (N_27117,N_26130,N_26740);
nand U27118 (N_27118,N_26057,N_26541);
and U27119 (N_27119,N_26024,N_26279);
nor U27120 (N_27120,N_26399,N_26269);
or U27121 (N_27121,N_26422,N_26044);
and U27122 (N_27122,N_26600,N_26526);
nand U27123 (N_27123,N_26437,N_26509);
or U27124 (N_27124,N_26685,N_26147);
xnor U27125 (N_27125,N_26581,N_26306);
nor U27126 (N_27126,N_26291,N_26479);
xnor U27127 (N_27127,N_26893,N_26107);
and U27128 (N_27128,N_26869,N_26796);
or U27129 (N_27129,N_26441,N_26427);
xnor U27130 (N_27130,N_26523,N_26220);
nor U27131 (N_27131,N_26376,N_26571);
or U27132 (N_27132,N_26930,N_26952);
and U27133 (N_27133,N_26504,N_26368);
and U27134 (N_27134,N_26389,N_26568);
and U27135 (N_27135,N_26878,N_26204);
nand U27136 (N_27136,N_26928,N_26145);
xnor U27137 (N_27137,N_26184,N_26483);
and U27138 (N_27138,N_26721,N_26840);
nand U27139 (N_27139,N_26733,N_26308);
or U27140 (N_27140,N_26979,N_26030);
and U27141 (N_27141,N_26353,N_26732);
xor U27142 (N_27142,N_26345,N_26385);
nand U27143 (N_27143,N_26692,N_26288);
or U27144 (N_27144,N_26361,N_26499);
xor U27145 (N_27145,N_26734,N_26825);
or U27146 (N_27146,N_26480,N_26722);
xor U27147 (N_27147,N_26991,N_26331);
xnor U27148 (N_27148,N_26401,N_26949);
nor U27149 (N_27149,N_26690,N_26866);
and U27150 (N_27150,N_26122,N_26981);
or U27151 (N_27151,N_26599,N_26968);
and U27152 (N_27152,N_26665,N_26849);
or U27153 (N_27153,N_26987,N_26402);
xnor U27154 (N_27154,N_26742,N_26397);
nand U27155 (N_27155,N_26378,N_26848);
nor U27156 (N_27156,N_26644,N_26580);
nand U27157 (N_27157,N_26521,N_26039);
and U27158 (N_27158,N_26026,N_26425);
or U27159 (N_27159,N_26506,N_26805);
nand U27160 (N_27160,N_26899,N_26993);
nand U27161 (N_27161,N_26578,N_26536);
nor U27162 (N_27162,N_26947,N_26609);
nand U27163 (N_27163,N_26654,N_26126);
and U27164 (N_27164,N_26211,N_26179);
or U27165 (N_27165,N_26396,N_26980);
nand U27166 (N_27166,N_26810,N_26253);
nor U27167 (N_27167,N_26611,N_26954);
nand U27168 (N_27168,N_26263,N_26984);
or U27169 (N_27169,N_26115,N_26592);
or U27170 (N_27170,N_26072,N_26489);
nor U27171 (N_27171,N_26909,N_26340);
nor U27172 (N_27172,N_26264,N_26229);
xor U27173 (N_27173,N_26748,N_26165);
nor U27174 (N_27174,N_26701,N_26290);
nor U27175 (N_27175,N_26962,N_26199);
and U27176 (N_27176,N_26156,N_26817);
or U27177 (N_27177,N_26804,N_26105);
xnor U27178 (N_27178,N_26747,N_26628);
nor U27179 (N_27179,N_26311,N_26082);
nor U27180 (N_27180,N_26957,N_26841);
and U27181 (N_27181,N_26668,N_26901);
nand U27182 (N_27182,N_26788,N_26795);
nor U27183 (N_27183,N_26743,N_26106);
nor U27184 (N_27184,N_26240,N_26305);
or U27185 (N_27185,N_26193,N_26464);
and U27186 (N_27186,N_26736,N_26889);
xnor U27187 (N_27187,N_26945,N_26851);
nand U27188 (N_27188,N_26390,N_26081);
and U27189 (N_27189,N_26746,N_26653);
nand U27190 (N_27190,N_26927,N_26894);
or U27191 (N_27191,N_26128,N_26012);
nor U27192 (N_27192,N_26254,N_26041);
nand U27193 (N_27193,N_26363,N_26969);
or U27194 (N_27194,N_26937,N_26902);
or U27195 (N_27195,N_26320,N_26978);
nor U27196 (N_27196,N_26558,N_26886);
and U27197 (N_27197,N_26842,N_26132);
nor U27198 (N_27198,N_26908,N_26787);
or U27199 (N_27199,N_26585,N_26863);
xor U27200 (N_27200,N_26688,N_26777);
xor U27201 (N_27201,N_26356,N_26589);
nand U27202 (N_27202,N_26416,N_26525);
nand U27203 (N_27203,N_26047,N_26032);
nand U27204 (N_27204,N_26251,N_26705);
xnor U27205 (N_27205,N_26140,N_26241);
or U27206 (N_27206,N_26673,N_26920);
or U27207 (N_27207,N_26974,N_26414);
nor U27208 (N_27208,N_26392,N_26284);
or U27209 (N_27209,N_26429,N_26679);
and U27210 (N_27210,N_26326,N_26781);
or U27211 (N_27211,N_26410,N_26681);
or U27212 (N_27212,N_26775,N_26307);
xor U27213 (N_27213,N_26216,N_26691);
and U27214 (N_27214,N_26876,N_26508);
nand U27215 (N_27215,N_26921,N_26045);
or U27216 (N_27216,N_26960,N_26704);
and U27217 (N_27217,N_26430,N_26111);
and U27218 (N_27218,N_26900,N_26486);
or U27219 (N_27219,N_26633,N_26820);
nor U27220 (N_27220,N_26084,N_26752);
and U27221 (N_27221,N_26730,N_26186);
nor U27222 (N_27222,N_26034,N_26439);
nand U27223 (N_27223,N_26477,N_26312);
or U27224 (N_27224,N_26598,N_26963);
or U27225 (N_27225,N_26966,N_26617);
xnor U27226 (N_27226,N_26426,N_26760);
xnor U27227 (N_27227,N_26144,N_26135);
xor U27228 (N_27228,N_26689,N_26406);
nor U27229 (N_27229,N_26080,N_26587);
xnor U27230 (N_27230,N_26434,N_26323);
or U27231 (N_27231,N_26884,N_26873);
or U27232 (N_27232,N_26338,N_26502);
or U27233 (N_27233,N_26089,N_26161);
nor U27234 (N_27234,N_26087,N_26322);
or U27235 (N_27235,N_26468,N_26906);
nor U27236 (N_27236,N_26341,N_26001);
or U27237 (N_27237,N_26564,N_26778);
xnor U27238 (N_27238,N_26803,N_26432);
or U27239 (N_27239,N_26163,N_26207);
and U27240 (N_27240,N_26765,N_26720);
nor U27241 (N_27241,N_26623,N_26821);
nor U27242 (N_27242,N_26758,N_26890);
or U27243 (N_27243,N_26374,N_26619);
or U27244 (N_27244,N_26350,N_26484);
nand U27245 (N_27245,N_26615,N_26624);
and U27246 (N_27246,N_26674,N_26714);
or U27247 (N_27247,N_26377,N_26444);
nor U27248 (N_27248,N_26988,N_26613);
or U27249 (N_27249,N_26870,N_26493);
xor U27250 (N_27250,N_26522,N_26155);
or U27251 (N_27251,N_26608,N_26467);
or U27252 (N_27252,N_26274,N_26768);
nand U27253 (N_27253,N_26802,N_26294);
nor U27254 (N_27254,N_26936,N_26395);
xnor U27255 (N_27255,N_26846,N_26102);
xnor U27256 (N_27256,N_26456,N_26076);
nor U27257 (N_27257,N_26050,N_26258);
or U27258 (N_27258,N_26232,N_26027);
and U27259 (N_27259,N_26594,N_26693);
and U27260 (N_27260,N_26970,N_26343);
or U27261 (N_27261,N_26137,N_26794);
xnor U27262 (N_27262,N_26110,N_26844);
and U27263 (N_27263,N_26466,N_26992);
and U27264 (N_27264,N_26647,N_26330);
and U27265 (N_27265,N_26055,N_26698);
nand U27266 (N_27266,N_26557,N_26584);
nor U27267 (N_27267,N_26496,N_26310);
nand U27268 (N_27268,N_26883,N_26579);
nand U27269 (N_27269,N_26531,N_26022);
nand U27270 (N_27270,N_26741,N_26625);
xnor U27271 (N_27271,N_26381,N_26013);
and U27272 (N_27272,N_26127,N_26228);
and U27273 (N_27273,N_26236,N_26510);
nand U27274 (N_27274,N_26099,N_26713);
or U27275 (N_27275,N_26256,N_26998);
or U27276 (N_27276,N_26061,N_26139);
nand U27277 (N_27277,N_26753,N_26864);
nand U27278 (N_27278,N_26738,N_26660);
and U27279 (N_27279,N_26339,N_26046);
nand U27280 (N_27280,N_26922,N_26178);
nor U27281 (N_27281,N_26188,N_26176);
nor U27282 (N_27282,N_26129,N_26152);
or U27283 (N_27283,N_26138,N_26830);
nand U27284 (N_27284,N_26703,N_26358);
xor U27285 (N_27285,N_26818,N_26114);
nand U27286 (N_27286,N_26520,N_26407);
xnor U27287 (N_27287,N_26601,N_26806);
nand U27288 (N_27288,N_26018,N_26113);
xor U27289 (N_27289,N_26275,N_26605);
xor U27290 (N_27290,N_26540,N_26384);
xnor U27291 (N_27291,N_26507,N_26234);
nand U27292 (N_27292,N_26814,N_26519);
and U27293 (N_27293,N_26719,N_26697);
nand U27294 (N_27294,N_26164,N_26759);
and U27295 (N_27295,N_26659,N_26942);
nor U27296 (N_27296,N_26056,N_26117);
and U27297 (N_27297,N_26462,N_26093);
xnor U27298 (N_27298,N_26875,N_26067);
and U27299 (N_27299,N_26783,N_26121);
or U27300 (N_27300,N_26098,N_26811);
or U27301 (N_27301,N_26562,N_26880);
nand U27302 (N_27302,N_26459,N_26669);
and U27303 (N_27303,N_26347,N_26517);
xnor U27304 (N_27304,N_26272,N_26651);
nand U27305 (N_27305,N_26770,N_26597);
xor U27306 (N_27306,N_26295,N_26062);
and U27307 (N_27307,N_26666,N_26420);
and U27308 (N_27308,N_26255,N_26300);
nor U27309 (N_27309,N_26865,N_26200);
or U27310 (N_27310,N_26885,N_26143);
or U27311 (N_27311,N_26469,N_26233);
or U27312 (N_27312,N_26985,N_26418);
or U27313 (N_27313,N_26708,N_26874);
nor U27314 (N_27314,N_26646,N_26159);
nand U27315 (N_27315,N_26513,N_26816);
nor U27316 (N_27316,N_26146,N_26196);
xor U27317 (N_27317,N_26729,N_26727);
or U27318 (N_27318,N_26198,N_26446);
and U27319 (N_27319,N_26166,N_26983);
xnor U27320 (N_27320,N_26094,N_26270);
xnor U27321 (N_27321,N_26458,N_26299);
and U27322 (N_27322,N_26408,N_26495);
and U27323 (N_27323,N_26009,N_26344);
nand U27324 (N_27324,N_26488,N_26277);
and U27325 (N_27325,N_26941,N_26359);
and U27326 (N_27326,N_26551,N_26352);
xnor U27327 (N_27327,N_26582,N_26838);
and U27328 (N_27328,N_26097,N_26409);
and U27329 (N_27329,N_26686,N_26375);
nand U27330 (N_27330,N_26967,N_26386);
xnor U27331 (N_27331,N_26676,N_26544);
xor U27332 (N_27332,N_26750,N_26561);
and U27333 (N_27333,N_26898,N_26956);
xnor U27334 (N_27334,N_26503,N_26208);
and U27335 (N_27335,N_26500,N_26868);
nand U27336 (N_27336,N_26090,N_26049);
nand U27337 (N_27337,N_26852,N_26671);
or U27338 (N_27338,N_26773,N_26907);
nand U27339 (N_27339,N_26717,N_26709);
nand U27340 (N_27340,N_26769,N_26718);
nor U27341 (N_27341,N_26438,N_26950);
or U27342 (N_27342,N_26813,N_26372);
nor U27343 (N_27343,N_26478,N_26048);
and U27344 (N_27344,N_26393,N_26826);
and U27345 (N_27345,N_26031,N_26528);
or U27346 (N_27346,N_26190,N_26560);
xor U27347 (N_27347,N_26423,N_26328);
xnor U27348 (N_27348,N_26857,N_26567);
and U27349 (N_27349,N_26497,N_26250);
nand U27350 (N_27350,N_26351,N_26824);
or U27351 (N_27351,N_26539,N_26918);
nor U27352 (N_27352,N_26784,N_26929);
nor U27353 (N_27353,N_26621,N_26706);
xnor U27354 (N_27354,N_26083,N_26036);
xnor U27355 (N_27355,N_26005,N_26566);
or U27356 (N_27356,N_26965,N_26827);
nand U27357 (N_27357,N_26120,N_26916);
and U27358 (N_27358,N_26096,N_26845);
nand U27359 (N_27359,N_26224,N_26532);
nor U27360 (N_27360,N_26917,N_26638);
xor U27361 (N_27361,N_26382,N_26643);
and U27362 (N_27362,N_26182,N_26315);
and U27363 (N_27363,N_26298,N_26357);
or U27364 (N_27364,N_26014,N_26346);
xnor U27365 (N_27365,N_26524,N_26364);
or U27366 (N_27366,N_26629,N_26153);
nand U27367 (N_27367,N_26202,N_26075);
nor U27368 (N_27368,N_26367,N_26116);
or U27369 (N_27369,N_26749,N_26793);
and U27370 (N_27370,N_26209,N_26411);
nand U27371 (N_27371,N_26702,N_26964);
nor U27372 (N_27372,N_26296,N_26181);
and U27373 (N_27373,N_26943,N_26383);
or U27374 (N_27374,N_26715,N_26975);
nor U27375 (N_27375,N_26006,N_26879);
nor U27376 (N_27376,N_26158,N_26550);
and U27377 (N_27377,N_26131,N_26002);
nand U27378 (N_27378,N_26141,N_26616);
nand U27379 (N_27379,N_26073,N_26088);
or U27380 (N_27380,N_26314,N_26847);
xnor U27381 (N_27381,N_26549,N_26881);
xnor U27382 (N_27382,N_26940,N_26745);
and U27383 (N_27383,N_26990,N_26877);
xor U27384 (N_27384,N_26887,N_26185);
nor U27385 (N_27385,N_26699,N_26333);
and U27386 (N_27386,N_26398,N_26180);
nor U27387 (N_27387,N_26370,N_26077);
and U27388 (N_27388,N_26443,N_26373);
nor U27389 (N_27389,N_26754,N_26070);
xnor U27390 (N_27390,N_26417,N_26054);
nand U27391 (N_27391,N_26195,N_26641);
nand U27392 (N_27392,N_26667,N_26590);
xnor U27393 (N_27393,N_26612,N_26923);
nand U27394 (N_27394,N_26053,N_26835);
xnor U27395 (N_27395,N_26791,N_26553);
and U27396 (N_27396,N_26650,N_26008);
nand U27397 (N_27397,N_26932,N_26085);
xnor U27398 (N_27398,N_26850,N_26833);
or U27399 (N_27399,N_26670,N_26552);
and U27400 (N_27400,N_26944,N_26252);
nor U27401 (N_27401,N_26043,N_26380);
nand U27402 (N_27402,N_26812,N_26678);
and U27403 (N_27403,N_26515,N_26168);
nand U27404 (N_27404,N_26710,N_26904);
nand U27405 (N_27405,N_26799,N_26172);
or U27406 (N_27406,N_26935,N_26680);
and U27407 (N_27407,N_26652,N_26029);
nand U27408 (N_27408,N_26327,N_26092);
xor U27409 (N_27409,N_26453,N_26257);
nand U27410 (N_27410,N_26219,N_26999);
or U27411 (N_27411,N_26349,N_26133);
nand U27412 (N_27412,N_26766,N_26451);
or U27413 (N_27413,N_26834,N_26379);
xor U27414 (N_27414,N_26527,N_26419);
or U27415 (N_27415,N_26591,N_26663);
xnor U27416 (N_27416,N_26772,N_26973);
nor U27417 (N_27417,N_26831,N_26682);
xnor U27418 (N_27418,N_26259,N_26069);
nor U27419 (N_27419,N_26100,N_26786);
or U27420 (N_27420,N_26078,N_26636);
nand U27421 (N_27421,N_26266,N_26336);
nor U27422 (N_27422,N_26951,N_26595);
nand U27423 (N_27423,N_26529,N_26905);
nand U27424 (N_27424,N_26051,N_26620);
nand U27425 (N_27425,N_26728,N_26059);
and U27426 (N_27426,N_26239,N_26342);
and U27427 (N_27427,N_26997,N_26662);
nand U27428 (N_27428,N_26737,N_26603);
xnor U27429 (N_27429,N_26986,N_26808);
nor U27430 (N_27430,N_26809,N_26546);
xor U27431 (N_27431,N_26192,N_26919);
and U27432 (N_27432,N_26683,N_26895);
or U27433 (N_27433,N_26109,N_26642);
nand U27434 (N_27434,N_26832,N_26694);
and U27435 (N_27435,N_26572,N_26573);
xor U27436 (N_27436,N_26661,N_26217);
or U27437 (N_27437,N_26285,N_26404);
and U27438 (N_27438,N_26171,N_26672);
nor U27439 (N_27439,N_26302,N_26861);
nor U27440 (N_27440,N_26645,N_26387);
and U27441 (N_27441,N_26494,N_26779);
or U27442 (N_27442,N_26112,N_26431);
or U27443 (N_27443,N_26896,N_26281);
nand U27444 (N_27444,N_26607,N_26206);
and U27445 (N_27445,N_26435,N_26518);
xnor U27446 (N_27446,N_26424,N_26413);
and U27447 (N_27447,N_26071,N_26245);
nor U27448 (N_27448,N_26292,N_26118);
nand U27449 (N_27449,N_26996,N_26037);
xnor U27450 (N_27450,N_26150,N_26914);
nand U27451 (N_27451,N_26482,N_26449);
and U27452 (N_27452,N_26912,N_26286);
nor U27453 (N_27453,N_26771,N_26790);
xnor U27454 (N_27454,N_26891,N_26602);
nand U27455 (N_27455,N_26280,N_26010);
xor U27456 (N_27456,N_26162,N_26576);
or U27457 (N_27457,N_26871,N_26405);
or U27458 (N_27458,N_26261,N_26533);
xnor U27459 (N_27459,N_26205,N_26915);
and U27460 (N_27460,N_26035,N_26237);
nand U27461 (N_27461,N_26946,N_26317);
nor U27462 (N_27462,N_26490,N_26174);
nand U27463 (N_27463,N_26554,N_26003);
and U27464 (N_27464,N_26867,N_26157);
nor U27465 (N_27465,N_26474,N_26538);
nand U27466 (N_27466,N_26194,N_26774);
or U27467 (N_27467,N_26403,N_26491);
nand U27468 (N_27468,N_26516,N_26971);
nor U27469 (N_27469,N_26556,N_26225);
and U27470 (N_27470,N_26695,N_26586);
xnor U27471 (N_27471,N_26656,N_26756);
or U27472 (N_27472,N_26448,N_26369);
and U27473 (N_27473,N_26911,N_26365);
xor U27474 (N_27474,N_26675,N_26436);
nor U27475 (N_27475,N_26025,N_26481);
or U27476 (N_27476,N_26931,N_26925);
and U27477 (N_27477,N_26124,N_26400);
nand U27478 (N_27478,N_26064,N_26177);
xor U27479 (N_27479,N_26104,N_26303);
xnor U27480 (N_27480,N_26583,N_26514);
and U27481 (N_27481,N_26801,N_26542);
nor U27482 (N_27482,N_26631,N_26243);
nand U27483 (N_27483,N_26221,N_26632);
xnor U27484 (N_27484,N_26068,N_26142);
nor U27485 (N_27485,N_26856,N_26800);
or U27486 (N_27486,N_26739,N_26547);
xor U27487 (N_27487,N_26855,N_26938);
nor U27488 (N_27488,N_26173,N_26231);
xnor U27489 (N_27489,N_26321,N_26843);
and U27490 (N_27490,N_26348,N_26767);
and U27491 (N_27491,N_26278,N_26989);
xnor U27492 (N_27492,N_26125,N_26428);
and U27493 (N_27493,N_26548,N_26511);
nand U27494 (N_27494,N_26858,N_26994);
xnor U27495 (N_27495,N_26913,N_26108);
nand U27496 (N_27496,N_26577,N_26021);
or U27497 (N_27497,N_26197,N_26828);
and U27498 (N_27498,N_26897,N_26134);
nand U27499 (N_27499,N_26658,N_26822);
nor U27500 (N_27500,N_26294,N_26379);
or U27501 (N_27501,N_26728,N_26687);
xnor U27502 (N_27502,N_26182,N_26991);
or U27503 (N_27503,N_26271,N_26339);
or U27504 (N_27504,N_26006,N_26801);
and U27505 (N_27505,N_26654,N_26195);
nor U27506 (N_27506,N_26045,N_26528);
xnor U27507 (N_27507,N_26639,N_26670);
xor U27508 (N_27508,N_26582,N_26914);
nor U27509 (N_27509,N_26740,N_26290);
nor U27510 (N_27510,N_26291,N_26677);
nand U27511 (N_27511,N_26753,N_26909);
and U27512 (N_27512,N_26256,N_26720);
or U27513 (N_27513,N_26542,N_26422);
or U27514 (N_27514,N_26798,N_26854);
and U27515 (N_27515,N_26051,N_26442);
nand U27516 (N_27516,N_26039,N_26167);
and U27517 (N_27517,N_26505,N_26230);
nor U27518 (N_27518,N_26573,N_26707);
xor U27519 (N_27519,N_26096,N_26780);
xnor U27520 (N_27520,N_26402,N_26217);
or U27521 (N_27521,N_26486,N_26378);
nor U27522 (N_27522,N_26901,N_26356);
nor U27523 (N_27523,N_26771,N_26895);
nand U27524 (N_27524,N_26392,N_26160);
xnor U27525 (N_27525,N_26741,N_26482);
nand U27526 (N_27526,N_26399,N_26598);
and U27527 (N_27527,N_26534,N_26329);
and U27528 (N_27528,N_26823,N_26396);
and U27529 (N_27529,N_26968,N_26557);
nand U27530 (N_27530,N_26665,N_26501);
nor U27531 (N_27531,N_26805,N_26226);
nor U27532 (N_27532,N_26305,N_26484);
nor U27533 (N_27533,N_26841,N_26426);
or U27534 (N_27534,N_26166,N_26748);
nor U27535 (N_27535,N_26957,N_26986);
and U27536 (N_27536,N_26756,N_26169);
nor U27537 (N_27537,N_26900,N_26149);
xor U27538 (N_27538,N_26519,N_26066);
nor U27539 (N_27539,N_26348,N_26885);
or U27540 (N_27540,N_26912,N_26718);
or U27541 (N_27541,N_26821,N_26290);
or U27542 (N_27542,N_26178,N_26798);
nand U27543 (N_27543,N_26405,N_26203);
nand U27544 (N_27544,N_26681,N_26106);
xnor U27545 (N_27545,N_26286,N_26595);
nand U27546 (N_27546,N_26855,N_26954);
nor U27547 (N_27547,N_26390,N_26972);
nor U27548 (N_27548,N_26342,N_26955);
xor U27549 (N_27549,N_26201,N_26722);
and U27550 (N_27550,N_26840,N_26285);
or U27551 (N_27551,N_26779,N_26769);
xnor U27552 (N_27552,N_26452,N_26157);
nor U27553 (N_27553,N_26925,N_26654);
nand U27554 (N_27554,N_26477,N_26747);
nand U27555 (N_27555,N_26981,N_26627);
nor U27556 (N_27556,N_26112,N_26032);
xor U27557 (N_27557,N_26384,N_26493);
nor U27558 (N_27558,N_26771,N_26702);
nor U27559 (N_27559,N_26375,N_26599);
nor U27560 (N_27560,N_26385,N_26133);
nand U27561 (N_27561,N_26186,N_26602);
nand U27562 (N_27562,N_26488,N_26471);
and U27563 (N_27563,N_26445,N_26326);
and U27564 (N_27564,N_26009,N_26796);
or U27565 (N_27565,N_26470,N_26953);
or U27566 (N_27566,N_26723,N_26655);
nand U27567 (N_27567,N_26304,N_26381);
or U27568 (N_27568,N_26233,N_26036);
xnor U27569 (N_27569,N_26256,N_26920);
or U27570 (N_27570,N_26682,N_26396);
nor U27571 (N_27571,N_26809,N_26321);
or U27572 (N_27572,N_26832,N_26392);
xnor U27573 (N_27573,N_26449,N_26924);
or U27574 (N_27574,N_26107,N_26890);
or U27575 (N_27575,N_26239,N_26876);
or U27576 (N_27576,N_26329,N_26669);
nand U27577 (N_27577,N_26099,N_26541);
and U27578 (N_27578,N_26654,N_26627);
xor U27579 (N_27579,N_26122,N_26196);
nor U27580 (N_27580,N_26868,N_26388);
and U27581 (N_27581,N_26629,N_26611);
and U27582 (N_27582,N_26704,N_26256);
nor U27583 (N_27583,N_26424,N_26886);
nand U27584 (N_27584,N_26962,N_26651);
and U27585 (N_27585,N_26613,N_26842);
or U27586 (N_27586,N_26015,N_26430);
xnor U27587 (N_27587,N_26165,N_26800);
and U27588 (N_27588,N_26101,N_26673);
and U27589 (N_27589,N_26503,N_26870);
and U27590 (N_27590,N_26929,N_26157);
xor U27591 (N_27591,N_26550,N_26002);
nand U27592 (N_27592,N_26057,N_26146);
xor U27593 (N_27593,N_26894,N_26924);
nor U27594 (N_27594,N_26268,N_26788);
nand U27595 (N_27595,N_26234,N_26168);
or U27596 (N_27596,N_26902,N_26788);
nor U27597 (N_27597,N_26547,N_26116);
nand U27598 (N_27598,N_26194,N_26707);
or U27599 (N_27599,N_26409,N_26206);
nand U27600 (N_27600,N_26469,N_26952);
or U27601 (N_27601,N_26867,N_26510);
and U27602 (N_27602,N_26259,N_26993);
nand U27603 (N_27603,N_26218,N_26402);
nor U27604 (N_27604,N_26749,N_26207);
nand U27605 (N_27605,N_26543,N_26748);
or U27606 (N_27606,N_26660,N_26814);
nor U27607 (N_27607,N_26244,N_26401);
or U27608 (N_27608,N_26029,N_26505);
nor U27609 (N_27609,N_26114,N_26314);
nor U27610 (N_27610,N_26912,N_26625);
or U27611 (N_27611,N_26928,N_26371);
and U27612 (N_27612,N_26500,N_26849);
or U27613 (N_27613,N_26032,N_26147);
or U27614 (N_27614,N_26910,N_26929);
or U27615 (N_27615,N_26118,N_26285);
nand U27616 (N_27616,N_26500,N_26643);
nor U27617 (N_27617,N_26382,N_26461);
nand U27618 (N_27618,N_26237,N_26967);
nor U27619 (N_27619,N_26146,N_26136);
nand U27620 (N_27620,N_26409,N_26120);
nor U27621 (N_27621,N_26619,N_26417);
nand U27622 (N_27622,N_26144,N_26914);
and U27623 (N_27623,N_26053,N_26916);
or U27624 (N_27624,N_26618,N_26491);
xnor U27625 (N_27625,N_26725,N_26190);
and U27626 (N_27626,N_26857,N_26318);
and U27627 (N_27627,N_26981,N_26198);
and U27628 (N_27628,N_26503,N_26467);
nand U27629 (N_27629,N_26628,N_26584);
or U27630 (N_27630,N_26188,N_26620);
nor U27631 (N_27631,N_26449,N_26559);
or U27632 (N_27632,N_26621,N_26652);
or U27633 (N_27633,N_26720,N_26984);
nand U27634 (N_27634,N_26562,N_26723);
nand U27635 (N_27635,N_26662,N_26806);
nor U27636 (N_27636,N_26823,N_26904);
nand U27637 (N_27637,N_26761,N_26898);
nand U27638 (N_27638,N_26711,N_26940);
xnor U27639 (N_27639,N_26639,N_26945);
or U27640 (N_27640,N_26595,N_26201);
or U27641 (N_27641,N_26429,N_26237);
nor U27642 (N_27642,N_26323,N_26874);
and U27643 (N_27643,N_26988,N_26996);
nor U27644 (N_27644,N_26183,N_26627);
and U27645 (N_27645,N_26968,N_26463);
xor U27646 (N_27646,N_26049,N_26258);
nand U27647 (N_27647,N_26123,N_26929);
xor U27648 (N_27648,N_26735,N_26759);
or U27649 (N_27649,N_26097,N_26873);
nand U27650 (N_27650,N_26406,N_26527);
and U27651 (N_27651,N_26151,N_26474);
or U27652 (N_27652,N_26215,N_26008);
xor U27653 (N_27653,N_26571,N_26406);
nor U27654 (N_27654,N_26018,N_26693);
xnor U27655 (N_27655,N_26624,N_26794);
xor U27656 (N_27656,N_26767,N_26980);
xor U27657 (N_27657,N_26172,N_26228);
and U27658 (N_27658,N_26223,N_26420);
nor U27659 (N_27659,N_26071,N_26073);
and U27660 (N_27660,N_26678,N_26956);
or U27661 (N_27661,N_26912,N_26095);
xor U27662 (N_27662,N_26622,N_26250);
nor U27663 (N_27663,N_26068,N_26627);
nor U27664 (N_27664,N_26270,N_26449);
nor U27665 (N_27665,N_26993,N_26610);
nand U27666 (N_27666,N_26441,N_26453);
nor U27667 (N_27667,N_26248,N_26442);
nand U27668 (N_27668,N_26456,N_26688);
or U27669 (N_27669,N_26415,N_26646);
nor U27670 (N_27670,N_26127,N_26993);
xor U27671 (N_27671,N_26258,N_26468);
xor U27672 (N_27672,N_26039,N_26782);
nand U27673 (N_27673,N_26926,N_26886);
or U27674 (N_27674,N_26747,N_26454);
xor U27675 (N_27675,N_26656,N_26420);
nand U27676 (N_27676,N_26320,N_26724);
or U27677 (N_27677,N_26260,N_26044);
nor U27678 (N_27678,N_26652,N_26312);
or U27679 (N_27679,N_26880,N_26876);
nor U27680 (N_27680,N_26288,N_26479);
or U27681 (N_27681,N_26430,N_26989);
nor U27682 (N_27682,N_26903,N_26927);
nor U27683 (N_27683,N_26551,N_26520);
or U27684 (N_27684,N_26373,N_26764);
and U27685 (N_27685,N_26084,N_26607);
or U27686 (N_27686,N_26900,N_26607);
nand U27687 (N_27687,N_26747,N_26725);
and U27688 (N_27688,N_26379,N_26345);
and U27689 (N_27689,N_26016,N_26551);
nand U27690 (N_27690,N_26091,N_26808);
nor U27691 (N_27691,N_26517,N_26275);
xor U27692 (N_27692,N_26136,N_26262);
nor U27693 (N_27693,N_26959,N_26330);
or U27694 (N_27694,N_26753,N_26274);
nand U27695 (N_27695,N_26982,N_26032);
xor U27696 (N_27696,N_26252,N_26041);
nand U27697 (N_27697,N_26720,N_26897);
xnor U27698 (N_27698,N_26763,N_26623);
or U27699 (N_27699,N_26093,N_26882);
nand U27700 (N_27700,N_26914,N_26761);
or U27701 (N_27701,N_26086,N_26945);
and U27702 (N_27702,N_26645,N_26486);
or U27703 (N_27703,N_26840,N_26902);
and U27704 (N_27704,N_26306,N_26835);
and U27705 (N_27705,N_26957,N_26179);
nor U27706 (N_27706,N_26639,N_26664);
nand U27707 (N_27707,N_26410,N_26424);
nor U27708 (N_27708,N_26720,N_26289);
or U27709 (N_27709,N_26706,N_26728);
or U27710 (N_27710,N_26794,N_26049);
nand U27711 (N_27711,N_26589,N_26892);
or U27712 (N_27712,N_26080,N_26445);
and U27713 (N_27713,N_26534,N_26621);
and U27714 (N_27714,N_26414,N_26620);
xor U27715 (N_27715,N_26107,N_26123);
nor U27716 (N_27716,N_26679,N_26936);
or U27717 (N_27717,N_26524,N_26885);
xor U27718 (N_27718,N_26227,N_26363);
nor U27719 (N_27719,N_26681,N_26552);
or U27720 (N_27720,N_26814,N_26171);
nand U27721 (N_27721,N_26254,N_26308);
or U27722 (N_27722,N_26991,N_26658);
and U27723 (N_27723,N_26386,N_26496);
or U27724 (N_27724,N_26040,N_26849);
and U27725 (N_27725,N_26176,N_26351);
or U27726 (N_27726,N_26513,N_26867);
and U27727 (N_27727,N_26842,N_26542);
nor U27728 (N_27728,N_26252,N_26393);
or U27729 (N_27729,N_26446,N_26217);
nand U27730 (N_27730,N_26268,N_26462);
xor U27731 (N_27731,N_26978,N_26987);
nor U27732 (N_27732,N_26797,N_26090);
nor U27733 (N_27733,N_26696,N_26879);
nand U27734 (N_27734,N_26514,N_26580);
and U27735 (N_27735,N_26511,N_26744);
xor U27736 (N_27736,N_26999,N_26232);
or U27737 (N_27737,N_26270,N_26608);
nor U27738 (N_27738,N_26211,N_26904);
or U27739 (N_27739,N_26866,N_26064);
nand U27740 (N_27740,N_26250,N_26096);
nand U27741 (N_27741,N_26209,N_26833);
xor U27742 (N_27742,N_26512,N_26014);
and U27743 (N_27743,N_26394,N_26112);
nor U27744 (N_27744,N_26430,N_26171);
nand U27745 (N_27745,N_26869,N_26471);
and U27746 (N_27746,N_26460,N_26384);
xnor U27747 (N_27747,N_26041,N_26977);
xor U27748 (N_27748,N_26819,N_26985);
or U27749 (N_27749,N_26583,N_26222);
or U27750 (N_27750,N_26356,N_26023);
xnor U27751 (N_27751,N_26499,N_26891);
nand U27752 (N_27752,N_26222,N_26872);
nand U27753 (N_27753,N_26633,N_26594);
xor U27754 (N_27754,N_26787,N_26111);
and U27755 (N_27755,N_26826,N_26282);
nor U27756 (N_27756,N_26971,N_26166);
nand U27757 (N_27757,N_26003,N_26858);
nand U27758 (N_27758,N_26796,N_26593);
xnor U27759 (N_27759,N_26159,N_26853);
nor U27760 (N_27760,N_26976,N_26127);
nor U27761 (N_27761,N_26039,N_26939);
xor U27762 (N_27762,N_26564,N_26933);
xnor U27763 (N_27763,N_26086,N_26095);
and U27764 (N_27764,N_26186,N_26742);
and U27765 (N_27765,N_26918,N_26573);
xnor U27766 (N_27766,N_26509,N_26143);
nand U27767 (N_27767,N_26789,N_26585);
nand U27768 (N_27768,N_26903,N_26069);
or U27769 (N_27769,N_26185,N_26236);
nand U27770 (N_27770,N_26919,N_26373);
xnor U27771 (N_27771,N_26230,N_26020);
or U27772 (N_27772,N_26896,N_26519);
xor U27773 (N_27773,N_26351,N_26338);
nand U27774 (N_27774,N_26768,N_26921);
and U27775 (N_27775,N_26600,N_26760);
xor U27776 (N_27776,N_26474,N_26404);
and U27777 (N_27777,N_26500,N_26197);
nand U27778 (N_27778,N_26417,N_26304);
nand U27779 (N_27779,N_26371,N_26933);
nor U27780 (N_27780,N_26553,N_26426);
nor U27781 (N_27781,N_26860,N_26795);
or U27782 (N_27782,N_26246,N_26130);
or U27783 (N_27783,N_26981,N_26888);
and U27784 (N_27784,N_26275,N_26485);
nor U27785 (N_27785,N_26148,N_26693);
xor U27786 (N_27786,N_26301,N_26466);
xor U27787 (N_27787,N_26620,N_26128);
or U27788 (N_27788,N_26290,N_26427);
or U27789 (N_27789,N_26169,N_26185);
or U27790 (N_27790,N_26121,N_26671);
nand U27791 (N_27791,N_26584,N_26408);
nand U27792 (N_27792,N_26704,N_26606);
or U27793 (N_27793,N_26010,N_26094);
and U27794 (N_27794,N_26562,N_26924);
xnor U27795 (N_27795,N_26254,N_26100);
nor U27796 (N_27796,N_26828,N_26799);
nand U27797 (N_27797,N_26224,N_26926);
xnor U27798 (N_27798,N_26676,N_26839);
or U27799 (N_27799,N_26594,N_26118);
nor U27800 (N_27800,N_26386,N_26334);
xnor U27801 (N_27801,N_26423,N_26532);
nor U27802 (N_27802,N_26034,N_26369);
or U27803 (N_27803,N_26120,N_26826);
nor U27804 (N_27804,N_26226,N_26107);
nor U27805 (N_27805,N_26968,N_26299);
nor U27806 (N_27806,N_26872,N_26174);
xor U27807 (N_27807,N_26041,N_26553);
xnor U27808 (N_27808,N_26560,N_26262);
xor U27809 (N_27809,N_26213,N_26109);
xnor U27810 (N_27810,N_26806,N_26280);
and U27811 (N_27811,N_26243,N_26987);
nand U27812 (N_27812,N_26139,N_26886);
xnor U27813 (N_27813,N_26547,N_26062);
or U27814 (N_27814,N_26088,N_26459);
nand U27815 (N_27815,N_26443,N_26329);
nor U27816 (N_27816,N_26261,N_26724);
or U27817 (N_27817,N_26154,N_26164);
and U27818 (N_27818,N_26352,N_26154);
and U27819 (N_27819,N_26604,N_26564);
nand U27820 (N_27820,N_26733,N_26712);
and U27821 (N_27821,N_26242,N_26782);
or U27822 (N_27822,N_26444,N_26810);
nor U27823 (N_27823,N_26561,N_26485);
nor U27824 (N_27824,N_26215,N_26626);
and U27825 (N_27825,N_26905,N_26490);
nand U27826 (N_27826,N_26539,N_26074);
nand U27827 (N_27827,N_26627,N_26143);
xnor U27828 (N_27828,N_26057,N_26888);
and U27829 (N_27829,N_26558,N_26860);
and U27830 (N_27830,N_26965,N_26541);
or U27831 (N_27831,N_26496,N_26805);
and U27832 (N_27832,N_26271,N_26090);
nand U27833 (N_27833,N_26252,N_26401);
xor U27834 (N_27834,N_26184,N_26662);
and U27835 (N_27835,N_26523,N_26367);
xnor U27836 (N_27836,N_26599,N_26296);
or U27837 (N_27837,N_26301,N_26886);
xnor U27838 (N_27838,N_26279,N_26523);
xnor U27839 (N_27839,N_26989,N_26210);
nor U27840 (N_27840,N_26250,N_26680);
nand U27841 (N_27841,N_26108,N_26894);
nor U27842 (N_27842,N_26336,N_26634);
xnor U27843 (N_27843,N_26529,N_26301);
nor U27844 (N_27844,N_26418,N_26171);
xnor U27845 (N_27845,N_26304,N_26057);
nor U27846 (N_27846,N_26440,N_26310);
xor U27847 (N_27847,N_26805,N_26995);
and U27848 (N_27848,N_26872,N_26572);
xor U27849 (N_27849,N_26806,N_26813);
or U27850 (N_27850,N_26250,N_26970);
xor U27851 (N_27851,N_26299,N_26675);
nand U27852 (N_27852,N_26977,N_26485);
nand U27853 (N_27853,N_26096,N_26025);
xor U27854 (N_27854,N_26134,N_26430);
nand U27855 (N_27855,N_26526,N_26585);
or U27856 (N_27856,N_26229,N_26280);
or U27857 (N_27857,N_26787,N_26494);
xnor U27858 (N_27858,N_26092,N_26522);
and U27859 (N_27859,N_26133,N_26931);
nand U27860 (N_27860,N_26502,N_26664);
or U27861 (N_27861,N_26299,N_26321);
and U27862 (N_27862,N_26842,N_26641);
xor U27863 (N_27863,N_26464,N_26924);
or U27864 (N_27864,N_26560,N_26853);
or U27865 (N_27865,N_26620,N_26309);
nand U27866 (N_27866,N_26018,N_26014);
nor U27867 (N_27867,N_26593,N_26787);
and U27868 (N_27868,N_26769,N_26495);
or U27869 (N_27869,N_26893,N_26182);
nand U27870 (N_27870,N_26893,N_26812);
nand U27871 (N_27871,N_26825,N_26983);
and U27872 (N_27872,N_26049,N_26693);
or U27873 (N_27873,N_26693,N_26857);
and U27874 (N_27874,N_26481,N_26102);
nand U27875 (N_27875,N_26364,N_26712);
xor U27876 (N_27876,N_26721,N_26925);
xor U27877 (N_27877,N_26739,N_26482);
xor U27878 (N_27878,N_26038,N_26259);
nand U27879 (N_27879,N_26739,N_26267);
nor U27880 (N_27880,N_26412,N_26024);
or U27881 (N_27881,N_26586,N_26913);
and U27882 (N_27882,N_26671,N_26196);
or U27883 (N_27883,N_26237,N_26596);
and U27884 (N_27884,N_26244,N_26927);
and U27885 (N_27885,N_26265,N_26145);
xor U27886 (N_27886,N_26508,N_26789);
xnor U27887 (N_27887,N_26890,N_26522);
nand U27888 (N_27888,N_26653,N_26090);
and U27889 (N_27889,N_26260,N_26972);
nand U27890 (N_27890,N_26589,N_26914);
and U27891 (N_27891,N_26185,N_26925);
nand U27892 (N_27892,N_26212,N_26072);
xnor U27893 (N_27893,N_26071,N_26510);
xnor U27894 (N_27894,N_26650,N_26320);
nor U27895 (N_27895,N_26684,N_26161);
xnor U27896 (N_27896,N_26061,N_26728);
and U27897 (N_27897,N_26244,N_26321);
or U27898 (N_27898,N_26861,N_26415);
or U27899 (N_27899,N_26970,N_26857);
or U27900 (N_27900,N_26470,N_26141);
nor U27901 (N_27901,N_26629,N_26276);
xnor U27902 (N_27902,N_26320,N_26907);
and U27903 (N_27903,N_26245,N_26320);
nand U27904 (N_27904,N_26556,N_26315);
and U27905 (N_27905,N_26640,N_26096);
xor U27906 (N_27906,N_26168,N_26146);
xor U27907 (N_27907,N_26244,N_26923);
nor U27908 (N_27908,N_26374,N_26665);
nand U27909 (N_27909,N_26636,N_26894);
nand U27910 (N_27910,N_26722,N_26694);
nand U27911 (N_27911,N_26800,N_26592);
and U27912 (N_27912,N_26904,N_26667);
nor U27913 (N_27913,N_26867,N_26421);
xor U27914 (N_27914,N_26795,N_26887);
nand U27915 (N_27915,N_26492,N_26005);
nand U27916 (N_27916,N_26533,N_26014);
xnor U27917 (N_27917,N_26428,N_26311);
or U27918 (N_27918,N_26113,N_26326);
and U27919 (N_27919,N_26527,N_26567);
nor U27920 (N_27920,N_26410,N_26778);
nor U27921 (N_27921,N_26817,N_26814);
xnor U27922 (N_27922,N_26773,N_26414);
xnor U27923 (N_27923,N_26744,N_26781);
and U27924 (N_27924,N_26654,N_26149);
xnor U27925 (N_27925,N_26753,N_26060);
or U27926 (N_27926,N_26497,N_26114);
or U27927 (N_27927,N_26460,N_26255);
nand U27928 (N_27928,N_26256,N_26203);
and U27929 (N_27929,N_26339,N_26294);
nor U27930 (N_27930,N_26304,N_26903);
or U27931 (N_27931,N_26377,N_26266);
nand U27932 (N_27932,N_26016,N_26380);
or U27933 (N_27933,N_26202,N_26055);
nand U27934 (N_27934,N_26123,N_26449);
nor U27935 (N_27935,N_26088,N_26675);
nor U27936 (N_27936,N_26846,N_26751);
nand U27937 (N_27937,N_26561,N_26364);
xor U27938 (N_27938,N_26006,N_26473);
nand U27939 (N_27939,N_26192,N_26943);
or U27940 (N_27940,N_26400,N_26278);
nand U27941 (N_27941,N_26245,N_26476);
and U27942 (N_27942,N_26442,N_26685);
or U27943 (N_27943,N_26338,N_26227);
and U27944 (N_27944,N_26646,N_26248);
nand U27945 (N_27945,N_26958,N_26027);
or U27946 (N_27946,N_26364,N_26426);
nand U27947 (N_27947,N_26798,N_26873);
and U27948 (N_27948,N_26093,N_26104);
xnor U27949 (N_27949,N_26425,N_26210);
nor U27950 (N_27950,N_26451,N_26298);
nor U27951 (N_27951,N_26820,N_26428);
and U27952 (N_27952,N_26401,N_26668);
nor U27953 (N_27953,N_26284,N_26958);
or U27954 (N_27954,N_26241,N_26416);
or U27955 (N_27955,N_26476,N_26075);
and U27956 (N_27956,N_26487,N_26212);
xor U27957 (N_27957,N_26110,N_26252);
and U27958 (N_27958,N_26215,N_26553);
nor U27959 (N_27959,N_26850,N_26385);
nand U27960 (N_27960,N_26949,N_26976);
xor U27961 (N_27961,N_26105,N_26600);
xor U27962 (N_27962,N_26422,N_26160);
xor U27963 (N_27963,N_26172,N_26346);
and U27964 (N_27964,N_26551,N_26635);
xnor U27965 (N_27965,N_26740,N_26169);
xnor U27966 (N_27966,N_26591,N_26962);
or U27967 (N_27967,N_26416,N_26625);
and U27968 (N_27968,N_26693,N_26434);
xnor U27969 (N_27969,N_26724,N_26544);
nor U27970 (N_27970,N_26867,N_26333);
and U27971 (N_27971,N_26971,N_26635);
and U27972 (N_27972,N_26841,N_26972);
nor U27973 (N_27973,N_26710,N_26651);
nand U27974 (N_27974,N_26219,N_26054);
and U27975 (N_27975,N_26121,N_26970);
nor U27976 (N_27976,N_26841,N_26772);
nor U27977 (N_27977,N_26516,N_26157);
nand U27978 (N_27978,N_26033,N_26498);
or U27979 (N_27979,N_26903,N_26747);
nor U27980 (N_27980,N_26078,N_26556);
or U27981 (N_27981,N_26936,N_26000);
or U27982 (N_27982,N_26576,N_26554);
xnor U27983 (N_27983,N_26849,N_26538);
nand U27984 (N_27984,N_26387,N_26297);
xor U27985 (N_27985,N_26379,N_26469);
xnor U27986 (N_27986,N_26097,N_26844);
xor U27987 (N_27987,N_26582,N_26228);
xnor U27988 (N_27988,N_26130,N_26791);
xor U27989 (N_27989,N_26106,N_26766);
xnor U27990 (N_27990,N_26628,N_26132);
or U27991 (N_27991,N_26270,N_26181);
or U27992 (N_27992,N_26259,N_26216);
nand U27993 (N_27993,N_26751,N_26867);
or U27994 (N_27994,N_26555,N_26777);
and U27995 (N_27995,N_26319,N_26348);
xnor U27996 (N_27996,N_26633,N_26220);
xor U27997 (N_27997,N_26576,N_26698);
nor U27998 (N_27998,N_26119,N_26596);
xor U27999 (N_27999,N_26403,N_26236);
nand U28000 (N_28000,N_27025,N_27711);
xor U28001 (N_28001,N_27879,N_27475);
xnor U28002 (N_28002,N_27418,N_27786);
and U28003 (N_28003,N_27087,N_27054);
nand U28004 (N_28004,N_27616,N_27365);
and U28005 (N_28005,N_27202,N_27580);
xor U28006 (N_28006,N_27305,N_27849);
or U28007 (N_28007,N_27122,N_27628);
xnor U28008 (N_28008,N_27390,N_27785);
xnor U28009 (N_28009,N_27234,N_27922);
xor U28010 (N_28010,N_27892,N_27139);
and U28011 (N_28011,N_27039,N_27593);
nor U28012 (N_28012,N_27421,N_27230);
and U28013 (N_28013,N_27167,N_27319);
nand U28014 (N_28014,N_27448,N_27348);
nor U28015 (N_28015,N_27683,N_27840);
nor U28016 (N_28016,N_27138,N_27859);
and U28017 (N_28017,N_27053,N_27597);
nor U28018 (N_28018,N_27187,N_27267);
nand U28019 (N_28019,N_27431,N_27153);
and U28020 (N_28020,N_27451,N_27841);
and U28021 (N_28021,N_27759,N_27293);
nand U28022 (N_28022,N_27211,N_27097);
xor U28023 (N_28023,N_27046,N_27066);
or U28024 (N_28024,N_27984,N_27930);
xnor U28025 (N_28025,N_27265,N_27399);
nor U28026 (N_28026,N_27615,N_27261);
nor U28027 (N_28027,N_27180,N_27354);
or U28028 (N_28028,N_27441,N_27817);
xor U28029 (N_28029,N_27359,N_27538);
xnor U28030 (N_28030,N_27907,N_27585);
xor U28031 (N_28031,N_27413,N_27326);
xnor U28032 (N_28032,N_27452,N_27308);
nor U28033 (N_28033,N_27581,N_27869);
and U28034 (N_28034,N_27101,N_27292);
nor U28035 (N_28035,N_27419,N_27182);
nor U28036 (N_28036,N_27081,N_27734);
xor U28037 (N_28037,N_27106,N_27056);
nor U28038 (N_28038,N_27744,N_27015);
nand U28039 (N_28039,N_27515,N_27221);
xnor U28040 (N_28040,N_27532,N_27216);
and U28041 (N_28041,N_27979,N_27266);
and U28042 (N_28042,N_27284,N_27188);
xnor U28043 (N_28043,N_27660,N_27014);
xor U28044 (N_28044,N_27131,N_27067);
nand U28045 (N_28045,N_27416,N_27932);
nand U28046 (N_28046,N_27889,N_27980);
and U28047 (N_28047,N_27177,N_27254);
nand U28048 (N_28048,N_27763,N_27070);
nand U28049 (N_28049,N_27232,N_27829);
xnor U28050 (N_28050,N_27862,N_27988);
xnor U28051 (N_28051,N_27827,N_27123);
nand U28052 (N_28052,N_27555,N_27022);
nand U28053 (N_28053,N_27483,N_27601);
nor U28054 (N_28054,N_27779,N_27787);
or U28055 (N_28055,N_27052,N_27834);
and U28056 (N_28056,N_27957,N_27074);
xor U28057 (N_28057,N_27549,N_27968);
xnor U28058 (N_28058,N_27595,N_27249);
xor U28059 (N_28059,N_27026,N_27871);
nor U28060 (N_28060,N_27161,N_27088);
nand U28061 (N_28061,N_27274,N_27237);
or U28062 (N_28062,N_27964,N_27965);
or U28063 (N_28063,N_27329,N_27507);
or U28064 (N_28064,N_27537,N_27133);
or U28065 (N_28065,N_27000,N_27598);
nor U28066 (N_28066,N_27058,N_27923);
nor U28067 (N_28067,N_27774,N_27065);
xor U28068 (N_28068,N_27076,N_27424);
xor U28069 (N_28069,N_27328,N_27544);
and U28070 (N_28070,N_27935,N_27158);
nor U28071 (N_28071,N_27134,N_27749);
nor U28072 (N_28072,N_27878,N_27140);
nand U28073 (N_28073,N_27479,N_27083);
and U28074 (N_28074,N_27799,N_27987);
and U28075 (N_28075,N_27658,N_27034);
xor U28076 (N_28076,N_27875,N_27371);
xor U28077 (N_28077,N_27588,N_27333);
nor U28078 (N_28078,N_27169,N_27652);
or U28079 (N_28079,N_27982,N_27407);
or U28080 (N_28080,N_27462,N_27969);
or U28081 (N_28081,N_27127,N_27038);
nor U28082 (N_28082,N_27440,N_27466);
and U28083 (N_28083,N_27801,N_27813);
or U28084 (N_28084,N_27704,N_27313);
nand U28085 (N_28085,N_27300,N_27499);
nand U28086 (N_28086,N_27807,N_27460);
or U28087 (N_28087,N_27746,N_27794);
or U28088 (N_28088,N_27602,N_27162);
nand U28089 (N_28089,N_27344,N_27568);
and U28090 (N_28090,N_27497,N_27379);
nor U28091 (N_28091,N_27903,N_27500);
or U28092 (N_28092,N_27524,N_27516);
nor U28093 (N_28093,N_27080,N_27008);
or U28094 (N_28094,N_27788,N_27393);
or U28095 (N_28095,N_27341,N_27989);
and U28096 (N_28096,N_27051,N_27727);
xor U28097 (N_28097,N_27558,N_27488);
nand U28098 (N_28098,N_27405,N_27285);
xnor U28099 (N_28099,N_27567,N_27013);
or U28100 (N_28100,N_27583,N_27011);
xor U28101 (N_28101,N_27619,N_27437);
and U28102 (N_28102,N_27600,N_27906);
xor U28103 (N_28103,N_27346,N_27942);
and U28104 (N_28104,N_27573,N_27887);
xnor U28105 (N_28105,N_27403,N_27719);
xnor U28106 (N_28106,N_27103,N_27603);
nand U28107 (N_28107,N_27385,N_27217);
xnor U28108 (N_28108,N_27425,N_27283);
xor U28109 (N_28109,N_27931,N_27156);
nor U28110 (N_28110,N_27229,N_27977);
nand U28111 (N_28111,N_27467,N_27946);
and U28112 (N_28112,N_27814,N_27837);
nand U28113 (N_28113,N_27018,N_27301);
or U28114 (N_28114,N_27246,N_27556);
nand U28115 (N_28115,N_27993,N_27494);
or U28116 (N_28116,N_27891,N_27082);
nor U28117 (N_28117,N_27157,N_27009);
nor U28118 (N_28118,N_27402,N_27427);
or U28119 (N_28119,N_27996,N_27325);
xor U28120 (N_28120,N_27173,N_27874);
nand U28121 (N_28121,N_27294,N_27536);
nand U28122 (N_28122,N_27272,N_27673);
nand U28123 (N_28123,N_27384,N_27322);
xor U28124 (N_28124,N_27278,N_27766);
nand U28125 (N_28125,N_27680,N_27414);
xor U28126 (N_28126,N_27443,N_27238);
xnor U28127 (N_28127,N_27706,N_27688);
or U28128 (N_28128,N_27643,N_27709);
and U28129 (N_28129,N_27925,N_27646);
xor U28130 (N_28130,N_27883,N_27004);
nand U28131 (N_28131,N_27350,N_27526);
or U28132 (N_28132,N_27960,N_27227);
and U28133 (N_28133,N_27468,N_27741);
xnor U28134 (N_28134,N_27019,N_27624);
or U28135 (N_28135,N_27258,N_27132);
and U28136 (N_28136,N_27391,N_27697);
nand U28137 (N_28137,N_27521,N_27193);
xnor U28138 (N_28138,N_27286,N_27802);
or U28139 (N_28139,N_27803,N_27320);
xnor U28140 (N_28140,N_27553,N_27509);
and U28141 (N_28141,N_27148,N_27487);
xnor U28142 (N_28142,N_27165,N_27796);
xnor U28143 (N_28143,N_27708,N_27447);
xnor U28144 (N_28144,N_27810,N_27454);
or U28145 (N_28145,N_27655,N_27474);
or U28146 (N_28146,N_27327,N_27059);
nand U28147 (N_28147,N_27843,N_27458);
nor U28148 (N_28148,N_27712,N_27342);
nand U28149 (N_28149,N_27533,N_27776);
nor U28150 (N_28150,N_27816,N_27369);
and U28151 (N_28151,N_27446,N_27453);
nand U28152 (N_28152,N_27522,N_27061);
nand U28153 (N_28153,N_27951,N_27679);
nand U28154 (N_28154,N_27075,N_27682);
xnor U28155 (N_28155,N_27044,N_27607);
and U28156 (N_28156,N_27715,N_27469);
nand U28157 (N_28157,N_27240,N_27141);
or U28158 (N_28158,N_27504,N_27528);
or U28159 (N_28159,N_27846,N_27164);
xnor U28160 (N_28160,N_27444,N_27137);
nor U28161 (N_28161,N_27896,N_27858);
and U28162 (N_28162,N_27560,N_27853);
and U28163 (N_28163,N_27557,N_27480);
xor U28164 (N_28164,N_27692,N_27842);
nand U28165 (N_28165,N_27364,N_27231);
and U28166 (N_28166,N_27999,N_27698);
nor U28167 (N_28167,N_27376,N_27085);
nand U28168 (N_28168,N_27702,N_27861);
xnor U28169 (N_28169,N_27339,N_27545);
and U28170 (N_28170,N_27733,N_27257);
and U28171 (N_28171,N_27663,N_27060);
nand U28172 (N_28172,N_27863,N_27765);
and U28173 (N_28173,N_27579,N_27491);
nand U28174 (N_28174,N_27184,N_27831);
or U28175 (N_28175,N_27933,N_27811);
nor U28176 (N_28176,N_27909,N_27430);
and U28177 (N_28177,N_27894,N_27501);
or U28178 (N_28178,N_27210,N_27714);
or U28179 (N_28179,N_27605,N_27695);
or U28180 (N_28180,N_27954,N_27147);
xnor U28181 (N_28181,N_27872,N_27481);
or U28182 (N_28182,N_27970,N_27561);
nand U28183 (N_28183,N_27798,N_27484);
xor U28184 (N_28184,N_27535,N_27126);
xnor U28185 (N_28185,N_27928,N_27244);
and U28186 (N_28186,N_27084,N_27685);
or U28187 (N_28187,N_27113,N_27546);
nand U28188 (N_28188,N_27415,N_27657);
or U28189 (N_28189,N_27125,N_27160);
nor U28190 (N_28190,N_27269,N_27168);
or U28191 (N_28191,N_27592,N_27195);
or U28192 (N_28192,N_27299,N_27529);
or U28193 (N_28193,N_27310,N_27335);
xor U28194 (N_28194,N_27422,N_27915);
nor U28195 (N_28195,N_27985,N_27574);
and U28196 (N_28196,N_27362,N_27128);
xor U28197 (N_28197,N_27382,N_27830);
and U28198 (N_28198,N_27208,N_27108);
and U28199 (N_28199,N_27893,N_27949);
xnor U28200 (N_28200,N_27490,N_27028);
xnor U28201 (N_28201,N_27207,N_27476);
nand U28202 (N_28202,N_27352,N_27495);
xor U28203 (N_28203,N_27198,N_27815);
xnor U28204 (N_28204,N_27963,N_27392);
and U28205 (N_28205,N_27865,N_27275);
nor U28206 (N_28206,N_27724,N_27215);
or U28207 (N_28207,N_27099,N_27644);
or U28208 (N_28208,N_27465,N_27656);
and U28209 (N_28209,N_27036,N_27884);
and U28210 (N_28210,N_27040,N_27604);
and U28211 (N_28211,N_27357,N_27701);
xnor U28212 (N_28212,N_27191,N_27944);
and U28213 (N_28213,N_27921,N_27057);
nor U28214 (N_28214,N_27434,N_27591);
and U28215 (N_28215,N_27317,N_27590);
and U28216 (N_28216,N_27255,N_27677);
nor U28217 (N_28217,N_27825,N_27594);
nor U28218 (N_28218,N_27855,N_27091);
and U28219 (N_28219,N_27042,N_27678);
nand U28220 (N_28220,N_27408,N_27653);
nor U28221 (N_28221,N_27378,N_27205);
nand U28222 (N_28222,N_27629,N_27666);
nand U28223 (N_28223,N_27832,N_27991);
and U28224 (N_28224,N_27705,N_27681);
and U28225 (N_28225,N_27927,N_27069);
or U28226 (N_28226,N_27661,N_27966);
or U28227 (N_28227,N_27398,N_27690);
and U28228 (N_28228,N_27730,N_27924);
nand U28229 (N_28229,N_27645,N_27394);
and U28230 (N_28230,N_27718,N_27631);
nor U28231 (N_28231,N_27745,N_27107);
or U28232 (N_28232,N_27135,N_27948);
nor U28233 (N_28233,N_27845,N_27092);
and U28234 (N_28234,N_27510,N_27667);
xor U28235 (N_28235,N_27630,N_27659);
or U28236 (N_28236,N_27256,N_27450);
nor U28237 (N_28237,N_27212,N_27247);
or U28238 (N_28238,N_27050,N_27228);
and U28239 (N_28239,N_27241,N_27296);
nor U28240 (N_28240,N_27569,N_27353);
nor U28241 (N_28241,N_27513,N_27596);
or U28242 (N_28242,N_27613,N_27401);
nor U28243 (N_28243,N_27962,N_27078);
nand U28244 (N_28244,N_27121,N_27116);
xnor U28245 (N_28245,N_27260,N_27445);
nand U28246 (N_28246,N_27197,N_27530);
xnor U28247 (N_28247,N_27821,N_27505);
or U28248 (N_28248,N_27642,N_27145);
or U28249 (N_28249,N_27349,N_27587);
or U28250 (N_28250,N_27477,N_27967);
nand U28251 (N_28251,N_27668,N_27564);
xnor U28252 (N_28252,N_27485,N_27115);
nand U28253 (N_28253,N_27992,N_27201);
and U28254 (N_28254,N_27375,N_27901);
and U28255 (N_28255,N_27971,N_27020);
xnor U28256 (N_28256,N_27559,N_27769);
or U28257 (N_28257,N_27836,N_27850);
or U28258 (N_28258,N_27396,N_27732);
nand U28259 (N_28259,N_27321,N_27174);
or U28260 (N_28260,N_27753,N_27584);
and U28261 (N_28261,N_27760,N_27098);
or U28262 (N_28262,N_27771,N_27742);
and U28263 (N_28263,N_27372,N_27775);
or U28264 (N_28264,N_27345,N_27264);
xor U28265 (N_28265,N_27994,N_27442);
or U28266 (N_28266,N_27072,N_27102);
nand U28267 (N_28267,N_27439,N_27527);
or U28268 (N_28268,N_27886,N_27649);
nor U28269 (N_28269,N_27792,N_27242);
nor U28270 (N_28270,N_27938,N_27897);
nand U28271 (N_28271,N_27151,N_27035);
xor U28272 (N_28272,N_27428,N_27047);
nor U28273 (N_28273,N_27055,N_27270);
xnor U28274 (N_28274,N_27824,N_27772);
xnor U28275 (N_28275,N_27833,N_27793);
xnor U28276 (N_28276,N_27459,N_27016);
or U28277 (N_28277,N_27110,N_27936);
nand U28278 (N_28278,N_27885,N_27611);
or U28279 (N_28279,N_27117,N_27323);
nor U28280 (N_28280,N_27634,N_27370);
nor U28281 (N_28281,N_27178,N_27130);
xnor U28282 (N_28282,N_27812,N_27699);
nor U28283 (N_28283,N_27502,N_27064);
and U28284 (N_28284,N_27343,N_27282);
nand U28285 (N_28285,N_27571,N_27280);
nor U28286 (N_28286,N_27626,N_27163);
xor U28287 (N_28287,N_27956,N_27086);
xnor U28288 (N_28288,N_27472,N_27981);
or U28289 (N_28289,N_27806,N_27176);
or U28290 (N_28290,N_27623,N_27033);
or U28291 (N_28291,N_27728,N_27435);
nand U28292 (N_28292,N_27318,N_27650);
or U28293 (N_28293,N_27412,N_27664);
nand U28294 (N_28294,N_27464,N_27752);
xnor U28295 (N_28295,N_27703,N_27498);
and U28296 (N_28296,N_27622,N_27031);
nor U28297 (N_28297,N_27236,N_27676);
xnor U28298 (N_28298,N_27330,N_27291);
and U28299 (N_28299,N_27143,N_27917);
xnor U28300 (N_28300,N_27795,N_27461);
nor U28301 (N_28301,N_27181,N_27610);
nor U28302 (N_28302,N_27554,N_27154);
and U28303 (N_28303,N_27916,N_27271);
xor U28304 (N_28304,N_27332,N_27689);
nor U28305 (N_28305,N_27614,N_27226);
nor U28306 (N_28306,N_27190,N_27974);
nor U28307 (N_28307,N_27214,N_27914);
or U28308 (N_28308,N_27782,N_27144);
nor U28309 (N_28309,N_27905,N_27170);
nand U28310 (N_28310,N_27700,N_27512);
and U28311 (N_28311,N_27627,N_27941);
xnor U28312 (N_28312,N_27438,N_27279);
nor U28313 (N_28313,N_27492,N_27095);
xor U28314 (N_28314,N_27868,N_27606);
nor U28315 (N_28315,N_27707,N_27518);
nand U28316 (N_28316,N_27609,N_27789);
nand U28317 (N_28317,N_27882,N_27926);
nand U28318 (N_28318,N_27851,N_27783);
nor U28319 (N_28319,N_27196,N_27640);
or U28320 (N_28320,N_27961,N_27496);
xor U28321 (N_28321,N_27423,N_27192);
xnor U28322 (N_28322,N_27118,N_27089);
or U28323 (N_28323,N_27639,N_27073);
xor U28324 (N_28324,N_27189,N_27550);
and U28325 (N_28325,N_27005,N_27404);
and U28326 (N_28326,N_27976,N_27338);
xor U28327 (N_28327,N_27111,N_27790);
xor U28328 (N_28328,N_27312,N_27542);
nand U28329 (N_28329,N_27826,N_27919);
nand U28330 (N_28330,N_27721,N_27710);
and U28331 (N_28331,N_27847,N_27959);
nand U28332 (N_28332,N_27289,N_27360);
xnor U28333 (N_28333,N_27213,N_27621);
nand U28334 (N_28334,N_27514,N_27809);
xor U28335 (N_28335,N_27436,N_27331);
or U28336 (N_28336,N_27315,N_27366);
nor U28337 (N_28337,N_27898,N_27804);
or U28338 (N_28338,N_27090,N_27368);
nand U28339 (N_28339,N_27911,N_27204);
xor U28340 (N_28340,N_27943,N_27854);
xor U28341 (N_28341,N_27367,N_27647);
nor U28342 (N_28342,N_27043,N_27648);
or U28343 (N_28343,N_27222,N_27395);
and U28344 (N_28344,N_27781,N_27671);
or U28345 (N_28345,N_27870,N_27290);
nand U28346 (N_28346,N_27761,N_27735);
nor U28347 (N_28347,N_27867,N_27021);
and U28348 (N_28348,N_27041,N_27929);
xnor U28349 (N_28349,N_27547,N_27400);
xor U28350 (N_28350,N_27314,N_27818);
nand U28351 (N_28351,N_27209,N_27503);
or U28352 (N_28352,N_27027,N_27149);
xor U28353 (N_28353,N_27767,N_27262);
nand U28354 (N_28354,N_27852,N_27159);
and U28355 (N_28355,N_27540,N_27218);
or U28356 (N_28356,N_27429,N_27152);
nor U28357 (N_28357,N_27720,N_27633);
xor U28358 (N_28358,N_27958,N_27309);
xnor U28359 (N_28359,N_27100,N_27150);
xor U28360 (N_28360,N_27662,N_27203);
nand U28361 (N_28361,N_27737,N_27062);
nor U28362 (N_28362,N_27520,N_27912);
nor U28363 (N_28363,N_27273,N_27904);
and U28364 (N_28364,N_27361,N_27881);
or U28365 (N_28365,N_27839,N_27751);
and U28366 (N_28366,N_27420,N_27096);
nor U28367 (N_28367,N_27934,N_27142);
nand U28368 (N_28368,N_27417,N_27489);
or U28369 (N_28369,N_27486,N_27037);
xnor U28370 (N_28370,N_27819,N_27030);
and U28371 (N_28371,N_27835,N_27541);
xnor U28372 (N_28372,N_27800,N_27525);
nand U28373 (N_28373,N_27316,N_27243);
nor U28374 (N_28374,N_27635,N_27572);
xor U28375 (N_28375,N_27860,N_27743);
nand U28376 (N_28376,N_27873,N_27433);
nor U28377 (N_28377,N_27995,N_27768);
and U28378 (N_28378,N_27828,N_27808);
nand U28379 (N_28379,N_27551,N_27687);
nor U28380 (N_28380,N_27939,N_27780);
nand U28381 (N_28381,N_27511,N_27302);
nor U28382 (N_28382,N_27473,N_27007);
and U28383 (N_28383,N_27531,N_27023);
nand U28384 (N_28384,N_27347,N_27471);
nand U28385 (N_28385,N_27277,N_27674);
nor U28386 (N_28386,N_27747,N_27166);
nor U28387 (N_28387,N_27336,N_27268);
xor U28388 (N_28388,N_27713,N_27857);
nor U28389 (N_28389,N_27194,N_27478);
nand U28390 (N_28390,N_27770,N_27844);
nor U28391 (N_28391,N_27206,N_27548);
xnor U28392 (N_28392,N_27750,N_27311);
and U28393 (N_28393,N_27612,N_27432);
and U28394 (N_28394,N_27983,N_27672);
and U28395 (N_28395,N_27045,N_27577);
or U28396 (N_28396,N_27129,N_27112);
nor U28397 (N_28397,N_27575,N_27665);
nor U28398 (N_28398,N_27124,N_27063);
nor U28399 (N_28399,N_27387,N_27017);
nor U28400 (N_28400,N_27457,N_27716);
xor U28401 (N_28401,N_27986,N_27455);
nor U28402 (N_28402,N_27298,N_27777);
or U28403 (N_28403,N_27534,N_27406);
nor U28404 (N_28404,N_27729,N_27397);
xnor U28405 (N_28405,N_27670,N_27470);
and U28406 (N_28406,N_27306,N_27071);
and U28407 (N_28407,N_27105,N_27723);
xor U28408 (N_28408,N_27224,N_27002);
nand U28409 (N_28409,N_27864,N_27651);
or U28410 (N_28410,N_27155,N_27411);
or U28411 (N_28411,N_27654,N_27562);
and U28412 (N_28412,N_27386,N_27848);
and U28413 (N_28413,N_27784,N_27748);
and U28414 (N_28414,N_27493,N_27304);
and U28415 (N_28415,N_27764,N_27726);
xor U28416 (N_28416,N_27625,N_27250);
and U28417 (N_28417,N_27093,N_27693);
nor U28418 (N_28418,N_27109,N_27997);
or U28419 (N_28419,N_27937,N_27281);
xor U28420 (N_28420,N_27186,N_27219);
or U28421 (N_28421,N_27363,N_27620);
and U28422 (N_28422,N_27079,N_27355);
nor U28423 (N_28423,N_27990,N_27029);
xnor U28424 (N_28424,N_27900,N_27945);
nor U28425 (N_28425,N_27136,N_27899);
or U28426 (N_28426,N_27920,N_27589);
nor U28427 (N_28427,N_27972,N_27918);
xor U28428 (N_28428,N_27582,N_27172);
xor U28429 (N_28429,N_27245,N_27175);
or U28430 (N_28430,N_27722,N_27199);
or U28431 (N_28431,N_27998,N_27565);
xor U28432 (N_28432,N_27276,N_27637);
or U28433 (N_28433,N_27003,N_27773);
xnor U28434 (N_28434,N_27248,N_27955);
xnor U28435 (N_28435,N_27739,N_27641);
nand U28436 (N_28436,N_27902,N_27736);
nor U28437 (N_28437,N_27104,N_27295);
xor U28438 (N_28438,N_27694,N_27225);
nor U28439 (N_28439,N_27077,N_27684);
nand U28440 (N_28440,N_27686,N_27910);
nor U28441 (N_28441,N_27940,N_27757);
nand U28442 (N_28442,N_27740,N_27953);
and U28443 (N_28443,N_27303,N_27094);
and U28444 (N_28444,N_27973,N_27717);
and U28445 (N_28445,N_27895,N_27791);
or U28446 (N_28446,N_27381,N_27263);
xor U28447 (N_28447,N_27608,N_27638);
nor U28448 (N_28448,N_27820,N_27552);
nand U28449 (N_28449,N_27755,N_27388);
nor U28450 (N_28450,N_27952,N_27463);
and U28451 (N_28451,N_27950,N_27006);
or U28452 (N_28452,N_27340,N_27337);
nand U28453 (N_28453,N_27183,N_27012);
or U28454 (N_28454,N_27235,N_27506);
nor U28455 (N_28455,N_27576,N_27389);
nand U28456 (N_28456,N_27517,N_27866);
and U28457 (N_28457,N_27888,N_27508);
and U28458 (N_28458,N_27778,N_27179);
nor U28459 (N_28459,N_27599,N_27324);
xor U28460 (N_28460,N_27913,N_27856);
xor U28461 (N_28461,N_27185,N_27171);
nand U28462 (N_28462,N_27975,N_27307);
and U28463 (N_28463,N_27696,N_27120);
nand U28464 (N_28464,N_27632,N_27049);
nor U28465 (N_28465,N_27409,N_27252);
nor U28466 (N_28466,N_27200,N_27618);
xor U28467 (N_28467,N_27410,N_27288);
nor U28468 (N_28468,N_27877,N_27010);
and U28469 (N_28469,N_27797,N_27449);
or U28470 (N_28470,N_27566,N_27543);
or U28471 (N_28471,N_27563,N_27358);
and U28472 (N_28472,N_27758,N_27253);
nor U28473 (N_28473,N_27669,N_27377);
nand U28474 (N_28474,N_27119,N_27146);
nor U28475 (N_28475,N_27876,N_27114);
and U28476 (N_28476,N_27001,N_27351);
nand U28477 (N_28477,N_27426,N_27617);
nor U28478 (N_28478,N_27373,N_27032);
xor U28479 (N_28479,N_27251,N_27725);
nand U28480 (N_28480,N_27880,N_27805);
xor U28481 (N_28481,N_27239,N_27890);
nand U28482 (N_28482,N_27838,N_27523);
xnor U28483 (N_28483,N_27068,N_27978);
nand U28484 (N_28484,N_27287,N_27823);
nor U28485 (N_28485,N_27456,N_27383);
or U28486 (N_28486,N_27586,N_27570);
or U28487 (N_28487,N_27738,N_27636);
xnor U28488 (N_28488,N_27947,N_27233);
xnor U28489 (N_28489,N_27762,N_27334);
or U28490 (N_28490,N_27024,N_27519);
nand U28491 (N_28491,N_27731,N_27374);
nand U28492 (N_28492,N_27297,N_27539);
nor U28493 (N_28493,N_27482,N_27754);
nor U28494 (N_28494,N_27220,N_27356);
nand U28495 (N_28495,N_27223,N_27691);
and U28496 (N_28496,N_27675,N_27756);
xnor U28497 (N_28497,N_27380,N_27259);
nand U28498 (N_28498,N_27578,N_27908);
nand U28499 (N_28499,N_27822,N_27048);
or U28500 (N_28500,N_27106,N_27375);
xor U28501 (N_28501,N_27935,N_27971);
nand U28502 (N_28502,N_27820,N_27891);
xnor U28503 (N_28503,N_27719,N_27769);
nand U28504 (N_28504,N_27419,N_27237);
nor U28505 (N_28505,N_27477,N_27262);
nand U28506 (N_28506,N_27562,N_27418);
or U28507 (N_28507,N_27080,N_27040);
or U28508 (N_28508,N_27685,N_27588);
or U28509 (N_28509,N_27780,N_27147);
nand U28510 (N_28510,N_27366,N_27633);
nor U28511 (N_28511,N_27359,N_27070);
nand U28512 (N_28512,N_27225,N_27830);
and U28513 (N_28513,N_27339,N_27792);
and U28514 (N_28514,N_27234,N_27581);
and U28515 (N_28515,N_27492,N_27949);
nand U28516 (N_28516,N_27640,N_27773);
xor U28517 (N_28517,N_27471,N_27532);
nand U28518 (N_28518,N_27179,N_27358);
nor U28519 (N_28519,N_27148,N_27519);
or U28520 (N_28520,N_27451,N_27271);
or U28521 (N_28521,N_27314,N_27123);
and U28522 (N_28522,N_27866,N_27911);
nand U28523 (N_28523,N_27894,N_27042);
nand U28524 (N_28524,N_27675,N_27366);
nor U28525 (N_28525,N_27375,N_27402);
nand U28526 (N_28526,N_27538,N_27189);
and U28527 (N_28527,N_27092,N_27053);
xor U28528 (N_28528,N_27053,N_27406);
nand U28529 (N_28529,N_27782,N_27527);
xor U28530 (N_28530,N_27916,N_27395);
nand U28531 (N_28531,N_27121,N_27806);
nand U28532 (N_28532,N_27857,N_27246);
nand U28533 (N_28533,N_27135,N_27422);
nor U28534 (N_28534,N_27599,N_27229);
or U28535 (N_28535,N_27828,N_27140);
and U28536 (N_28536,N_27344,N_27461);
or U28537 (N_28537,N_27199,N_27917);
and U28538 (N_28538,N_27456,N_27227);
xnor U28539 (N_28539,N_27285,N_27881);
nand U28540 (N_28540,N_27776,N_27325);
nor U28541 (N_28541,N_27037,N_27177);
and U28542 (N_28542,N_27358,N_27222);
nor U28543 (N_28543,N_27795,N_27530);
xor U28544 (N_28544,N_27892,N_27560);
or U28545 (N_28545,N_27776,N_27724);
xor U28546 (N_28546,N_27947,N_27405);
or U28547 (N_28547,N_27448,N_27402);
xor U28548 (N_28548,N_27266,N_27479);
xnor U28549 (N_28549,N_27368,N_27096);
nor U28550 (N_28550,N_27706,N_27489);
or U28551 (N_28551,N_27190,N_27992);
xnor U28552 (N_28552,N_27887,N_27645);
nor U28553 (N_28553,N_27660,N_27118);
xnor U28554 (N_28554,N_27272,N_27561);
nand U28555 (N_28555,N_27012,N_27157);
xnor U28556 (N_28556,N_27854,N_27346);
or U28557 (N_28557,N_27293,N_27312);
or U28558 (N_28558,N_27927,N_27564);
and U28559 (N_28559,N_27194,N_27102);
or U28560 (N_28560,N_27915,N_27543);
or U28561 (N_28561,N_27321,N_27269);
or U28562 (N_28562,N_27353,N_27866);
xnor U28563 (N_28563,N_27919,N_27710);
nand U28564 (N_28564,N_27359,N_27605);
nand U28565 (N_28565,N_27147,N_27505);
xor U28566 (N_28566,N_27292,N_27727);
nor U28567 (N_28567,N_27583,N_27331);
and U28568 (N_28568,N_27206,N_27159);
or U28569 (N_28569,N_27651,N_27066);
nand U28570 (N_28570,N_27893,N_27738);
nor U28571 (N_28571,N_27662,N_27446);
nand U28572 (N_28572,N_27126,N_27989);
nor U28573 (N_28573,N_27285,N_27548);
nand U28574 (N_28574,N_27017,N_27955);
or U28575 (N_28575,N_27891,N_27575);
nor U28576 (N_28576,N_27263,N_27167);
or U28577 (N_28577,N_27863,N_27736);
nand U28578 (N_28578,N_27659,N_27906);
xnor U28579 (N_28579,N_27585,N_27161);
xnor U28580 (N_28580,N_27425,N_27948);
nand U28581 (N_28581,N_27298,N_27140);
or U28582 (N_28582,N_27380,N_27796);
nor U28583 (N_28583,N_27683,N_27114);
and U28584 (N_28584,N_27034,N_27608);
nand U28585 (N_28585,N_27667,N_27096);
nand U28586 (N_28586,N_27383,N_27175);
xor U28587 (N_28587,N_27631,N_27939);
nand U28588 (N_28588,N_27075,N_27927);
and U28589 (N_28589,N_27105,N_27586);
xnor U28590 (N_28590,N_27115,N_27042);
nand U28591 (N_28591,N_27328,N_27640);
nor U28592 (N_28592,N_27585,N_27214);
and U28593 (N_28593,N_27930,N_27902);
or U28594 (N_28594,N_27629,N_27523);
nor U28595 (N_28595,N_27966,N_27794);
xor U28596 (N_28596,N_27208,N_27817);
or U28597 (N_28597,N_27835,N_27960);
xor U28598 (N_28598,N_27357,N_27027);
nand U28599 (N_28599,N_27670,N_27983);
nand U28600 (N_28600,N_27904,N_27149);
nor U28601 (N_28601,N_27094,N_27021);
nor U28602 (N_28602,N_27266,N_27660);
or U28603 (N_28603,N_27659,N_27897);
xnor U28604 (N_28604,N_27455,N_27364);
or U28605 (N_28605,N_27033,N_27172);
or U28606 (N_28606,N_27710,N_27201);
xnor U28607 (N_28607,N_27039,N_27675);
xnor U28608 (N_28608,N_27898,N_27230);
and U28609 (N_28609,N_27349,N_27049);
nor U28610 (N_28610,N_27856,N_27433);
and U28611 (N_28611,N_27666,N_27131);
or U28612 (N_28612,N_27330,N_27068);
nand U28613 (N_28613,N_27305,N_27072);
and U28614 (N_28614,N_27552,N_27016);
nor U28615 (N_28615,N_27201,N_27809);
nand U28616 (N_28616,N_27171,N_27422);
or U28617 (N_28617,N_27676,N_27237);
or U28618 (N_28618,N_27099,N_27215);
nor U28619 (N_28619,N_27349,N_27095);
or U28620 (N_28620,N_27132,N_27248);
and U28621 (N_28621,N_27770,N_27984);
and U28622 (N_28622,N_27812,N_27266);
nand U28623 (N_28623,N_27403,N_27439);
or U28624 (N_28624,N_27882,N_27179);
and U28625 (N_28625,N_27460,N_27829);
or U28626 (N_28626,N_27920,N_27381);
and U28627 (N_28627,N_27755,N_27408);
or U28628 (N_28628,N_27779,N_27369);
or U28629 (N_28629,N_27982,N_27630);
xor U28630 (N_28630,N_27111,N_27568);
nor U28631 (N_28631,N_27057,N_27833);
nor U28632 (N_28632,N_27212,N_27022);
xor U28633 (N_28633,N_27332,N_27948);
nor U28634 (N_28634,N_27056,N_27310);
nor U28635 (N_28635,N_27828,N_27254);
nand U28636 (N_28636,N_27938,N_27044);
nand U28637 (N_28637,N_27314,N_27479);
xnor U28638 (N_28638,N_27088,N_27110);
or U28639 (N_28639,N_27399,N_27185);
xnor U28640 (N_28640,N_27646,N_27830);
xor U28641 (N_28641,N_27655,N_27105);
and U28642 (N_28642,N_27681,N_27857);
and U28643 (N_28643,N_27464,N_27868);
and U28644 (N_28644,N_27387,N_27379);
nand U28645 (N_28645,N_27443,N_27245);
or U28646 (N_28646,N_27734,N_27812);
or U28647 (N_28647,N_27894,N_27430);
nand U28648 (N_28648,N_27807,N_27450);
and U28649 (N_28649,N_27485,N_27138);
nor U28650 (N_28650,N_27172,N_27089);
nand U28651 (N_28651,N_27394,N_27446);
or U28652 (N_28652,N_27094,N_27378);
nor U28653 (N_28653,N_27312,N_27687);
nor U28654 (N_28654,N_27820,N_27443);
and U28655 (N_28655,N_27821,N_27340);
or U28656 (N_28656,N_27787,N_27698);
nand U28657 (N_28657,N_27517,N_27275);
and U28658 (N_28658,N_27232,N_27047);
or U28659 (N_28659,N_27706,N_27644);
nor U28660 (N_28660,N_27930,N_27852);
nand U28661 (N_28661,N_27249,N_27480);
xnor U28662 (N_28662,N_27431,N_27184);
nor U28663 (N_28663,N_27584,N_27441);
nand U28664 (N_28664,N_27004,N_27133);
xor U28665 (N_28665,N_27249,N_27422);
nand U28666 (N_28666,N_27839,N_27566);
xnor U28667 (N_28667,N_27324,N_27177);
xor U28668 (N_28668,N_27550,N_27361);
nor U28669 (N_28669,N_27498,N_27105);
xor U28670 (N_28670,N_27674,N_27713);
or U28671 (N_28671,N_27744,N_27553);
nor U28672 (N_28672,N_27360,N_27195);
nor U28673 (N_28673,N_27641,N_27625);
xor U28674 (N_28674,N_27722,N_27839);
and U28675 (N_28675,N_27244,N_27336);
nand U28676 (N_28676,N_27284,N_27663);
xnor U28677 (N_28677,N_27497,N_27494);
nand U28678 (N_28678,N_27339,N_27888);
nand U28679 (N_28679,N_27386,N_27477);
nor U28680 (N_28680,N_27177,N_27649);
nor U28681 (N_28681,N_27306,N_27641);
xor U28682 (N_28682,N_27652,N_27580);
nor U28683 (N_28683,N_27216,N_27726);
xor U28684 (N_28684,N_27038,N_27165);
nor U28685 (N_28685,N_27209,N_27879);
nor U28686 (N_28686,N_27147,N_27395);
and U28687 (N_28687,N_27225,N_27281);
and U28688 (N_28688,N_27449,N_27081);
or U28689 (N_28689,N_27019,N_27621);
or U28690 (N_28690,N_27959,N_27698);
nor U28691 (N_28691,N_27625,N_27390);
or U28692 (N_28692,N_27688,N_27811);
or U28693 (N_28693,N_27574,N_27229);
xor U28694 (N_28694,N_27451,N_27981);
or U28695 (N_28695,N_27545,N_27604);
nand U28696 (N_28696,N_27082,N_27936);
and U28697 (N_28697,N_27943,N_27914);
nor U28698 (N_28698,N_27946,N_27666);
nor U28699 (N_28699,N_27142,N_27568);
and U28700 (N_28700,N_27596,N_27661);
xnor U28701 (N_28701,N_27819,N_27884);
and U28702 (N_28702,N_27519,N_27923);
nand U28703 (N_28703,N_27784,N_27440);
nand U28704 (N_28704,N_27707,N_27863);
xor U28705 (N_28705,N_27894,N_27647);
nor U28706 (N_28706,N_27518,N_27254);
and U28707 (N_28707,N_27727,N_27805);
and U28708 (N_28708,N_27653,N_27577);
or U28709 (N_28709,N_27991,N_27040);
xnor U28710 (N_28710,N_27019,N_27103);
xnor U28711 (N_28711,N_27972,N_27521);
and U28712 (N_28712,N_27102,N_27190);
xnor U28713 (N_28713,N_27872,N_27115);
or U28714 (N_28714,N_27776,N_27334);
or U28715 (N_28715,N_27955,N_27444);
nor U28716 (N_28716,N_27034,N_27497);
nand U28717 (N_28717,N_27716,N_27468);
nand U28718 (N_28718,N_27029,N_27055);
or U28719 (N_28719,N_27823,N_27056);
nor U28720 (N_28720,N_27707,N_27859);
and U28721 (N_28721,N_27912,N_27749);
and U28722 (N_28722,N_27715,N_27693);
nand U28723 (N_28723,N_27242,N_27720);
nand U28724 (N_28724,N_27702,N_27200);
and U28725 (N_28725,N_27397,N_27115);
xor U28726 (N_28726,N_27372,N_27968);
and U28727 (N_28727,N_27335,N_27346);
xnor U28728 (N_28728,N_27703,N_27522);
and U28729 (N_28729,N_27796,N_27608);
or U28730 (N_28730,N_27851,N_27564);
nand U28731 (N_28731,N_27038,N_27142);
or U28732 (N_28732,N_27177,N_27265);
nand U28733 (N_28733,N_27840,N_27171);
xor U28734 (N_28734,N_27584,N_27037);
nor U28735 (N_28735,N_27737,N_27994);
nand U28736 (N_28736,N_27156,N_27778);
xnor U28737 (N_28737,N_27536,N_27540);
xor U28738 (N_28738,N_27112,N_27259);
nor U28739 (N_28739,N_27516,N_27602);
nor U28740 (N_28740,N_27404,N_27518);
nor U28741 (N_28741,N_27358,N_27029);
xor U28742 (N_28742,N_27619,N_27600);
and U28743 (N_28743,N_27376,N_27135);
and U28744 (N_28744,N_27261,N_27493);
or U28745 (N_28745,N_27014,N_27978);
or U28746 (N_28746,N_27058,N_27387);
and U28747 (N_28747,N_27988,N_27232);
nand U28748 (N_28748,N_27861,N_27661);
nand U28749 (N_28749,N_27882,N_27729);
xor U28750 (N_28750,N_27434,N_27065);
or U28751 (N_28751,N_27912,N_27785);
nor U28752 (N_28752,N_27394,N_27109);
xor U28753 (N_28753,N_27754,N_27257);
nor U28754 (N_28754,N_27241,N_27395);
and U28755 (N_28755,N_27405,N_27929);
xor U28756 (N_28756,N_27164,N_27439);
and U28757 (N_28757,N_27691,N_27372);
or U28758 (N_28758,N_27654,N_27308);
and U28759 (N_28759,N_27774,N_27152);
nand U28760 (N_28760,N_27301,N_27676);
nand U28761 (N_28761,N_27861,N_27253);
and U28762 (N_28762,N_27698,N_27100);
and U28763 (N_28763,N_27124,N_27233);
nand U28764 (N_28764,N_27644,N_27161);
xor U28765 (N_28765,N_27650,N_27192);
nand U28766 (N_28766,N_27444,N_27714);
nor U28767 (N_28767,N_27292,N_27757);
or U28768 (N_28768,N_27040,N_27306);
xnor U28769 (N_28769,N_27616,N_27202);
nor U28770 (N_28770,N_27070,N_27290);
and U28771 (N_28771,N_27847,N_27277);
nor U28772 (N_28772,N_27417,N_27700);
and U28773 (N_28773,N_27903,N_27078);
and U28774 (N_28774,N_27698,N_27132);
and U28775 (N_28775,N_27862,N_27059);
or U28776 (N_28776,N_27334,N_27023);
xnor U28777 (N_28777,N_27179,N_27688);
nor U28778 (N_28778,N_27294,N_27170);
xnor U28779 (N_28779,N_27690,N_27739);
and U28780 (N_28780,N_27225,N_27231);
xor U28781 (N_28781,N_27305,N_27634);
or U28782 (N_28782,N_27832,N_27743);
xnor U28783 (N_28783,N_27114,N_27689);
or U28784 (N_28784,N_27740,N_27924);
or U28785 (N_28785,N_27430,N_27148);
and U28786 (N_28786,N_27939,N_27411);
or U28787 (N_28787,N_27413,N_27581);
nor U28788 (N_28788,N_27302,N_27619);
nor U28789 (N_28789,N_27342,N_27503);
or U28790 (N_28790,N_27459,N_27654);
xnor U28791 (N_28791,N_27846,N_27689);
nor U28792 (N_28792,N_27692,N_27511);
nor U28793 (N_28793,N_27918,N_27133);
nor U28794 (N_28794,N_27425,N_27951);
or U28795 (N_28795,N_27803,N_27297);
or U28796 (N_28796,N_27429,N_27807);
nor U28797 (N_28797,N_27017,N_27415);
or U28798 (N_28798,N_27635,N_27406);
nand U28799 (N_28799,N_27697,N_27628);
and U28800 (N_28800,N_27690,N_27447);
xnor U28801 (N_28801,N_27496,N_27023);
and U28802 (N_28802,N_27456,N_27183);
or U28803 (N_28803,N_27408,N_27367);
and U28804 (N_28804,N_27875,N_27198);
or U28805 (N_28805,N_27279,N_27378);
and U28806 (N_28806,N_27520,N_27132);
or U28807 (N_28807,N_27170,N_27648);
nand U28808 (N_28808,N_27896,N_27079);
nor U28809 (N_28809,N_27987,N_27019);
nor U28810 (N_28810,N_27198,N_27138);
nor U28811 (N_28811,N_27857,N_27677);
or U28812 (N_28812,N_27620,N_27292);
and U28813 (N_28813,N_27998,N_27085);
nor U28814 (N_28814,N_27992,N_27215);
or U28815 (N_28815,N_27726,N_27859);
nor U28816 (N_28816,N_27483,N_27021);
and U28817 (N_28817,N_27597,N_27816);
and U28818 (N_28818,N_27647,N_27480);
xor U28819 (N_28819,N_27150,N_27238);
nor U28820 (N_28820,N_27217,N_27508);
nand U28821 (N_28821,N_27164,N_27380);
xor U28822 (N_28822,N_27985,N_27101);
xor U28823 (N_28823,N_27232,N_27527);
nand U28824 (N_28824,N_27894,N_27997);
nor U28825 (N_28825,N_27146,N_27982);
and U28826 (N_28826,N_27839,N_27256);
and U28827 (N_28827,N_27628,N_27864);
nor U28828 (N_28828,N_27813,N_27202);
or U28829 (N_28829,N_27094,N_27641);
or U28830 (N_28830,N_27442,N_27494);
or U28831 (N_28831,N_27640,N_27690);
and U28832 (N_28832,N_27938,N_27315);
nand U28833 (N_28833,N_27423,N_27243);
or U28834 (N_28834,N_27557,N_27917);
xnor U28835 (N_28835,N_27463,N_27373);
nand U28836 (N_28836,N_27667,N_27851);
nand U28837 (N_28837,N_27745,N_27861);
nand U28838 (N_28838,N_27862,N_27633);
nand U28839 (N_28839,N_27481,N_27550);
nand U28840 (N_28840,N_27529,N_27009);
nand U28841 (N_28841,N_27583,N_27629);
nand U28842 (N_28842,N_27806,N_27335);
xnor U28843 (N_28843,N_27988,N_27895);
and U28844 (N_28844,N_27918,N_27635);
nand U28845 (N_28845,N_27268,N_27085);
nand U28846 (N_28846,N_27792,N_27756);
xnor U28847 (N_28847,N_27239,N_27410);
xnor U28848 (N_28848,N_27777,N_27349);
or U28849 (N_28849,N_27876,N_27964);
xnor U28850 (N_28850,N_27383,N_27468);
and U28851 (N_28851,N_27113,N_27008);
nor U28852 (N_28852,N_27496,N_27210);
nor U28853 (N_28853,N_27323,N_27113);
xor U28854 (N_28854,N_27911,N_27517);
or U28855 (N_28855,N_27791,N_27309);
nand U28856 (N_28856,N_27114,N_27602);
xor U28857 (N_28857,N_27263,N_27845);
and U28858 (N_28858,N_27070,N_27158);
nand U28859 (N_28859,N_27556,N_27633);
nor U28860 (N_28860,N_27638,N_27292);
or U28861 (N_28861,N_27644,N_27360);
nand U28862 (N_28862,N_27699,N_27382);
or U28863 (N_28863,N_27924,N_27827);
nor U28864 (N_28864,N_27469,N_27362);
and U28865 (N_28865,N_27024,N_27527);
nand U28866 (N_28866,N_27540,N_27064);
nand U28867 (N_28867,N_27857,N_27445);
or U28868 (N_28868,N_27358,N_27002);
or U28869 (N_28869,N_27407,N_27353);
xnor U28870 (N_28870,N_27205,N_27922);
nand U28871 (N_28871,N_27318,N_27975);
xor U28872 (N_28872,N_27170,N_27834);
nor U28873 (N_28873,N_27899,N_27920);
nor U28874 (N_28874,N_27315,N_27963);
xor U28875 (N_28875,N_27039,N_27528);
nor U28876 (N_28876,N_27726,N_27929);
nand U28877 (N_28877,N_27768,N_27272);
or U28878 (N_28878,N_27422,N_27126);
or U28879 (N_28879,N_27675,N_27302);
nor U28880 (N_28880,N_27273,N_27440);
nand U28881 (N_28881,N_27544,N_27252);
nand U28882 (N_28882,N_27030,N_27124);
nor U28883 (N_28883,N_27205,N_27832);
nor U28884 (N_28884,N_27609,N_27897);
and U28885 (N_28885,N_27427,N_27841);
nand U28886 (N_28886,N_27794,N_27735);
or U28887 (N_28887,N_27498,N_27989);
nor U28888 (N_28888,N_27402,N_27765);
xor U28889 (N_28889,N_27681,N_27964);
nor U28890 (N_28890,N_27066,N_27910);
and U28891 (N_28891,N_27738,N_27891);
and U28892 (N_28892,N_27325,N_27820);
and U28893 (N_28893,N_27766,N_27887);
and U28894 (N_28894,N_27583,N_27788);
or U28895 (N_28895,N_27166,N_27725);
or U28896 (N_28896,N_27807,N_27350);
xor U28897 (N_28897,N_27488,N_27968);
nand U28898 (N_28898,N_27277,N_27944);
or U28899 (N_28899,N_27500,N_27776);
nor U28900 (N_28900,N_27066,N_27024);
xor U28901 (N_28901,N_27350,N_27864);
nor U28902 (N_28902,N_27263,N_27970);
xor U28903 (N_28903,N_27315,N_27539);
and U28904 (N_28904,N_27719,N_27575);
xnor U28905 (N_28905,N_27464,N_27555);
and U28906 (N_28906,N_27334,N_27382);
nor U28907 (N_28907,N_27352,N_27634);
nand U28908 (N_28908,N_27111,N_27055);
xnor U28909 (N_28909,N_27545,N_27896);
or U28910 (N_28910,N_27179,N_27894);
nand U28911 (N_28911,N_27548,N_27057);
and U28912 (N_28912,N_27218,N_27844);
xnor U28913 (N_28913,N_27790,N_27107);
nand U28914 (N_28914,N_27064,N_27827);
and U28915 (N_28915,N_27962,N_27172);
xnor U28916 (N_28916,N_27784,N_27453);
and U28917 (N_28917,N_27127,N_27223);
xnor U28918 (N_28918,N_27820,N_27119);
xnor U28919 (N_28919,N_27208,N_27105);
nor U28920 (N_28920,N_27477,N_27577);
xnor U28921 (N_28921,N_27997,N_27791);
nor U28922 (N_28922,N_27306,N_27923);
or U28923 (N_28923,N_27256,N_27825);
nor U28924 (N_28924,N_27893,N_27455);
xnor U28925 (N_28925,N_27865,N_27210);
xnor U28926 (N_28926,N_27606,N_27709);
xor U28927 (N_28927,N_27376,N_27104);
nand U28928 (N_28928,N_27876,N_27927);
or U28929 (N_28929,N_27320,N_27628);
nor U28930 (N_28930,N_27292,N_27664);
and U28931 (N_28931,N_27428,N_27832);
or U28932 (N_28932,N_27484,N_27264);
xnor U28933 (N_28933,N_27466,N_27989);
xnor U28934 (N_28934,N_27176,N_27633);
or U28935 (N_28935,N_27869,N_27236);
nand U28936 (N_28936,N_27479,N_27343);
or U28937 (N_28937,N_27028,N_27708);
and U28938 (N_28938,N_27536,N_27756);
and U28939 (N_28939,N_27904,N_27863);
xor U28940 (N_28940,N_27889,N_27547);
nand U28941 (N_28941,N_27421,N_27994);
xor U28942 (N_28942,N_27615,N_27225);
or U28943 (N_28943,N_27512,N_27550);
nand U28944 (N_28944,N_27133,N_27653);
nand U28945 (N_28945,N_27659,N_27060);
and U28946 (N_28946,N_27873,N_27047);
nand U28947 (N_28947,N_27692,N_27085);
nand U28948 (N_28948,N_27827,N_27651);
nand U28949 (N_28949,N_27835,N_27659);
nand U28950 (N_28950,N_27366,N_27874);
and U28951 (N_28951,N_27066,N_27085);
nor U28952 (N_28952,N_27188,N_27493);
nand U28953 (N_28953,N_27389,N_27263);
and U28954 (N_28954,N_27962,N_27210);
nor U28955 (N_28955,N_27618,N_27387);
and U28956 (N_28956,N_27833,N_27946);
xor U28957 (N_28957,N_27476,N_27172);
nand U28958 (N_28958,N_27857,N_27524);
xnor U28959 (N_28959,N_27727,N_27434);
nand U28960 (N_28960,N_27685,N_27516);
nor U28961 (N_28961,N_27226,N_27370);
and U28962 (N_28962,N_27848,N_27050);
nor U28963 (N_28963,N_27408,N_27558);
or U28964 (N_28964,N_27373,N_27700);
nand U28965 (N_28965,N_27125,N_27306);
and U28966 (N_28966,N_27263,N_27867);
nand U28967 (N_28967,N_27112,N_27353);
xnor U28968 (N_28968,N_27303,N_27994);
xnor U28969 (N_28969,N_27452,N_27636);
nor U28970 (N_28970,N_27099,N_27130);
nand U28971 (N_28971,N_27367,N_27303);
nand U28972 (N_28972,N_27007,N_27542);
and U28973 (N_28973,N_27811,N_27995);
xnor U28974 (N_28974,N_27048,N_27123);
nor U28975 (N_28975,N_27066,N_27564);
and U28976 (N_28976,N_27982,N_27465);
or U28977 (N_28977,N_27071,N_27982);
nand U28978 (N_28978,N_27924,N_27297);
xnor U28979 (N_28979,N_27388,N_27597);
and U28980 (N_28980,N_27775,N_27499);
or U28981 (N_28981,N_27286,N_27427);
or U28982 (N_28982,N_27323,N_27563);
xnor U28983 (N_28983,N_27039,N_27610);
and U28984 (N_28984,N_27094,N_27726);
and U28985 (N_28985,N_27085,N_27749);
xnor U28986 (N_28986,N_27248,N_27462);
and U28987 (N_28987,N_27251,N_27472);
nor U28988 (N_28988,N_27535,N_27976);
nor U28989 (N_28989,N_27321,N_27141);
nand U28990 (N_28990,N_27099,N_27728);
and U28991 (N_28991,N_27021,N_27583);
xnor U28992 (N_28992,N_27840,N_27492);
nand U28993 (N_28993,N_27731,N_27704);
and U28994 (N_28994,N_27652,N_27045);
and U28995 (N_28995,N_27801,N_27848);
or U28996 (N_28996,N_27742,N_27631);
nand U28997 (N_28997,N_27996,N_27745);
xor U28998 (N_28998,N_27642,N_27616);
xor U28999 (N_28999,N_27541,N_27844);
nand U29000 (N_29000,N_28449,N_28306);
xnor U29001 (N_29001,N_28122,N_28187);
nor U29002 (N_29002,N_28905,N_28647);
nor U29003 (N_29003,N_28917,N_28171);
or U29004 (N_29004,N_28781,N_28175);
nor U29005 (N_29005,N_28988,N_28915);
xor U29006 (N_29006,N_28046,N_28337);
or U29007 (N_29007,N_28383,N_28278);
xor U29008 (N_29008,N_28394,N_28293);
nand U29009 (N_29009,N_28238,N_28498);
nor U29010 (N_29010,N_28880,N_28902);
and U29011 (N_29011,N_28554,N_28019);
xnor U29012 (N_29012,N_28897,N_28058);
nand U29013 (N_29013,N_28166,N_28150);
xor U29014 (N_29014,N_28822,N_28323);
and U29015 (N_29015,N_28389,N_28937);
and U29016 (N_29016,N_28939,N_28797);
and U29017 (N_29017,N_28065,N_28120);
nand U29018 (N_29018,N_28220,N_28300);
or U29019 (N_29019,N_28553,N_28655);
nor U29020 (N_29020,N_28645,N_28342);
or U29021 (N_29021,N_28552,N_28452);
nand U29022 (N_29022,N_28321,N_28089);
or U29023 (N_29023,N_28987,N_28505);
nor U29024 (N_29024,N_28989,N_28431);
nand U29025 (N_29025,N_28198,N_28798);
and U29026 (N_29026,N_28954,N_28486);
xor U29027 (N_29027,N_28341,N_28748);
xnor U29028 (N_29028,N_28820,N_28966);
or U29029 (N_29029,N_28304,N_28203);
or U29030 (N_29030,N_28489,N_28417);
and U29031 (N_29031,N_28681,N_28995);
or U29032 (N_29032,N_28158,N_28901);
or U29033 (N_29033,N_28826,N_28453);
nor U29034 (N_29034,N_28879,N_28492);
nor U29035 (N_29035,N_28032,N_28547);
or U29036 (N_29036,N_28701,N_28882);
xor U29037 (N_29037,N_28087,N_28210);
nor U29038 (N_29038,N_28983,N_28715);
and U29039 (N_29039,N_28971,N_28626);
xnor U29040 (N_29040,N_28549,N_28025);
and U29041 (N_29041,N_28181,N_28139);
nand U29042 (N_29042,N_28275,N_28478);
xor U29043 (N_29043,N_28925,N_28422);
and U29044 (N_29044,N_28115,N_28455);
and U29045 (N_29045,N_28199,N_28081);
xnor U29046 (N_29046,N_28972,N_28885);
and U29047 (N_29047,N_28608,N_28672);
nand U29048 (N_29048,N_28393,N_28031);
nor U29049 (N_29049,N_28616,N_28804);
xor U29050 (N_29050,N_28690,N_28410);
xnor U29051 (N_29051,N_28338,N_28918);
nand U29052 (N_29052,N_28962,N_28042);
and U29053 (N_29053,N_28507,N_28644);
and U29054 (N_29054,N_28118,N_28803);
and U29055 (N_29055,N_28841,N_28322);
and U29056 (N_29056,N_28968,N_28783);
nor U29057 (N_29057,N_28869,N_28048);
nand U29058 (N_29058,N_28270,N_28045);
nand U29059 (N_29059,N_28908,N_28805);
nand U29060 (N_29060,N_28105,N_28794);
xnor U29061 (N_29061,N_28572,N_28251);
xor U29062 (N_29062,N_28702,N_28907);
xor U29063 (N_29063,N_28320,N_28381);
or U29064 (N_29064,N_28460,N_28793);
or U29065 (N_29065,N_28358,N_28131);
nand U29066 (N_29066,N_28629,N_28754);
or U29067 (N_29067,N_28414,N_28283);
nand U29068 (N_29068,N_28188,N_28319);
nand U29069 (N_29069,N_28531,N_28176);
nand U29070 (N_29070,N_28134,N_28887);
and U29071 (N_29071,N_28532,N_28237);
nand U29072 (N_29072,N_28407,N_28377);
or U29073 (N_29073,N_28740,N_28288);
nand U29074 (N_29074,N_28438,N_28566);
nand U29075 (N_29075,N_28536,N_28509);
and U29076 (N_29076,N_28420,N_28316);
or U29077 (N_29077,N_28018,N_28504);
nand U29078 (N_29078,N_28662,N_28934);
nor U29079 (N_29079,N_28511,N_28575);
and U29080 (N_29080,N_28390,N_28718);
xor U29081 (N_29081,N_28790,N_28625);
or U29082 (N_29082,N_28858,N_28415);
nand U29083 (N_29083,N_28162,N_28840);
xor U29084 (N_29084,N_28313,N_28052);
nor U29085 (N_29085,N_28580,N_28303);
xor U29086 (N_29086,N_28984,N_28236);
nand U29087 (N_29087,N_28722,N_28611);
or U29088 (N_29088,N_28109,N_28830);
nor U29089 (N_29089,N_28856,N_28761);
nand U29090 (N_29090,N_28838,N_28624);
or U29091 (N_29091,N_28765,N_28368);
or U29092 (N_29092,N_28101,N_28750);
nand U29093 (N_29093,N_28163,N_28221);
xnor U29094 (N_29094,N_28501,N_28851);
nor U29095 (N_29095,N_28396,N_28811);
nand U29096 (N_29096,N_28520,N_28408);
xnor U29097 (N_29097,N_28404,N_28670);
and U29098 (N_29098,N_28073,N_28848);
or U29099 (N_29099,N_28542,N_28627);
nor U29100 (N_29100,N_28413,N_28956);
xnor U29101 (N_29101,N_28529,N_28123);
nor U29102 (N_29102,N_28938,N_28815);
or U29103 (N_29103,N_28759,N_28014);
and U29104 (N_29104,N_28208,N_28117);
xnor U29105 (N_29105,N_28953,N_28684);
or U29106 (N_29106,N_28680,N_28853);
or U29107 (N_29107,N_28898,N_28654);
and U29108 (N_29108,N_28112,N_28516);
nand U29109 (N_29109,N_28430,N_28768);
or U29110 (N_29110,N_28332,N_28865);
or U29111 (N_29111,N_28242,N_28821);
or U29112 (N_29112,N_28854,N_28370);
or U29113 (N_29113,N_28806,N_28193);
nor U29114 (N_29114,N_28660,N_28714);
nor U29115 (N_29115,N_28427,N_28711);
or U29116 (N_29116,N_28209,N_28047);
nor U29117 (N_29117,N_28274,N_28556);
and U29118 (N_29118,N_28445,N_28379);
and U29119 (N_29119,N_28571,N_28291);
nor U29120 (N_29120,N_28965,N_28178);
or U29121 (N_29121,N_28265,N_28344);
nor U29122 (N_29122,N_28072,N_28997);
and U29123 (N_29123,N_28458,N_28307);
nor U29124 (N_29124,N_28837,N_28259);
nor U29125 (N_29125,N_28843,N_28472);
or U29126 (N_29126,N_28563,N_28214);
nand U29127 (N_29127,N_28710,N_28663);
and U29128 (N_29128,N_28948,N_28565);
xor U29129 (N_29129,N_28712,N_28059);
nor U29130 (N_29130,N_28677,N_28355);
nor U29131 (N_29131,N_28021,N_28305);
nand U29132 (N_29132,N_28870,N_28145);
xor U29133 (N_29133,N_28679,N_28814);
or U29134 (N_29134,N_28152,N_28037);
nand U29135 (N_29135,N_28651,N_28129);
or U29136 (N_29136,N_28530,N_28374);
xnor U29137 (N_29137,N_28574,N_28599);
nor U29138 (N_29138,N_28353,N_28577);
nor U29139 (N_29139,N_28622,N_28057);
and U29140 (N_29140,N_28528,N_28756);
nand U29141 (N_29141,N_28034,N_28619);
xor U29142 (N_29142,N_28771,N_28709);
nor U29143 (N_29143,N_28450,N_28088);
xnor U29144 (N_29144,N_28833,N_28085);
nand U29145 (N_29145,N_28212,N_28588);
and U29146 (N_29146,N_28280,N_28919);
xor U29147 (N_29147,N_28391,N_28700);
nor U29148 (N_29148,N_28312,N_28425);
and U29149 (N_29149,N_28373,N_28125);
nand U29150 (N_29150,N_28770,N_28113);
nor U29151 (N_29151,N_28979,N_28148);
nor U29152 (N_29152,N_28403,N_28914);
or U29153 (N_29153,N_28949,N_28816);
or U29154 (N_29154,N_28239,N_28384);
and U29155 (N_29155,N_28874,N_28285);
nand U29156 (N_29156,N_28156,N_28667);
nor U29157 (N_29157,N_28260,N_28524);
xnor U29158 (N_29158,N_28891,N_28920);
nor U29159 (N_29159,N_28096,N_28481);
nand U29160 (N_29160,N_28235,N_28000);
nor U29161 (N_29161,N_28931,N_28365);
and U29162 (N_29162,N_28564,N_28659);
nand U29163 (N_29163,N_28868,N_28197);
nand U29164 (N_29164,N_28196,N_28432);
xor U29165 (N_29165,N_28697,N_28475);
nor U29166 (N_29166,N_28884,N_28069);
nor U29167 (N_29167,N_28910,N_28423);
and U29168 (N_29168,N_28479,N_28185);
nor U29169 (N_29169,N_28512,N_28268);
nand U29170 (N_29170,N_28409,N_28245);
and U29171 (N_29171,N_28380,N_28468);
nand U29172 (N_29172,N_28476,N_28190);
or U29173 (N_29173,N_28114,N_28098);
or U29174 (N_29174,N_28053,N_28721);
nor U29175 (N_29175,N_28108,N_28436);
or U29176 (N_29176,N_28543,N_28827);
xor U29177 (N_29177,N_28986,N_28640);
nor U29178 (N_29178,N_28439,N_28272);
or U29179 (N_29179,N_28001,N_28596);
nor U29180 (N_29180,N_28978,N_28720);
nor U29181 (N_29181,N_28944,N_28585);
and U29182 (N_29182,N_28441,N_28782);
nand U29183 (N_29183,N_28298,N_28729);
and U29184 (N_29184,N_28240,N_28888);
or U29185 (N_29185,N_28703,N_28064);
or U29186 (N_29186,N_28977,N_28766);
nand U29187 (N_29187,N_28023,N_28998);
nor U29188 (N_29188,N_28142,N_28241);
or U29189 (N_29189,N_28991,N_28493);
or U29190 (N_29190,N_28459,N_28339);
nand U29191 (N_29191,N_28202,N_28578);
or U29192 (N_29192,N_28829,N_28138);
and U29193 (N_29193,N_28689,N_28008);
or U29194 (N_29194,N_28287,N_28082);
nor U29195 (N_29195,N_28996,N_28947);
nand U29196 (N_29196,N_28447,N_28533);
nand U29197 (N_29197,N_28839,N_28787);
nand U29198 (N_29198,N_28597,N_28252);
and U29199 (N_29199,N_28961,N_28642);
and U29200 (N_29200,N_28525,N_28144);
or U29201 (N_29201,N_28964,N_28485);
nand U29202 (N_29202,N_28876,N_28435);
or U29203 (N_29203,N_28835,N_28297);
nor U29204 (N_29204,N_28738,N_28006);
nor U29205 (N_29205,N_28906,N_28860);
and U29206 (N_29206,N_28605,N_28846);
xor U29207 (N_29207,N_28174,N_28755);
or U29208 (N_29208,N_28267,N_28067);
nor U29209 (N_29209,N_28567,N_28842);
or U29210 (N_29210,N_28107,N_28933);
nand U29211 (N_29211,N_28086,N_28687);
xor U29212 (N_29212,N_28716,N_28140);
nand U29213 (N_29213,N_28615,N_28799);
nor U29214 (N_29214,N_28426,N_28551);
xnor U29215 (N_29215,N_28537,N_28612);
and U29216 (N_29216,N_28364,N_28369);
and U29217 (N_29217,N_28154,N_28788);
and U29218 (N_29218,N_28650,N_28100);
nor U29219 (N_29219,N_28290,N_28637);
xor U29220 (N_29220,N_28730,N_28168);
nor U29221 (N_29221,N_28593,N_28442);
xnor U29222 (N_29222,N_28490,N_28121);
nand U29223 (N_29223,N_28179,N_28499);
nor U29224 (N_29224,N_28011,N_28315);
nand U29225 (N_29225,N_28469,N_28402);
nor U29226 (N_29226,N_28074,N_28598);
nor U29227 (N_29227,N_28473,N_28433);
nor U29228 (N_29228,N_28124,N_28013);
nand U29229 (N_29229,N_28392,N_28434);
nor U29230 (N_29230,N_28111,N_28292);
or U29231 (N_29231,N_28981,N_28881);
nand U29232 (N_29232,N_28155,N_28692);
or U29233 (N_29233,N_28457,N_28926);
xor U29234 (N_29234,N_28372,N_28103);
or U29235 (N_29235,N_28904,N_28062);
and U29236 (N_29236,N_28982,N_28657);
nand U29237 (N_29237,N_28590,N_28639);
nor U29238 (N_29238,N_28796,N_28040);
nor U29239 (N_29239,N_28527,N_28638);
nand U29240 (N_29240,N_28852,N_28277);
nor U29241 (N_29241,N_28661,N_28912);
and U29242 (N_29242,N_28429,N_28317);
or U29243 (N_29243,N_28694,N_28772);
nor U29244 (N_29244,N_28510,N_28517);
nand U29245 (N_29245,N_28182,N_28078);
nand U29246 (N_29246,N_28041,N_28487);
nand U29247 (N_29247,N_28800,N_28266);
nor U29248 (N_29248,N_28050,N_28515);
or U29249 (N_29249,N_28610,N_28892);
or U29250 (N_29250,N_28061,N_28688);
nor U29251 (N_29251,N_28500,N_28271);
nand U29252 (N_29252,N_28205,N_28620);
nor U29253 (N_29253,N_28932,N_28581);
xnor U29254 (N_29254,N_28132,N_28345);
xnor U29255 (N_29255,N_28204,N_28308);
nor U29256 (N_29256,N_28217,N_28818);
nand U29257 (N_29257,N_28147,N_28896);
xor U29258 (N_29258,N_28502,N_28877);
and U29259 (N_29259,N_28560,N_28617);
or U29260 (N_29260,N_28973,N_28792);
or U29261 (N_29261,N_28160,N_28232);
and U29262 (N_29262,N_28231,N_28159);
nand U29263 (N_29263,N_28301,N_28348);
and U29264 (N_29264,N_28728,N_28351);
nor U29265 (N_29265,N_28388,N_28299);
xnor U29266 (N_29266,N_28828,N_28464);
or U29267 (N_29267,N_28243,N_28136);
or U29268 (N_29268,N_28602,N_28462);
xor U29269 (N_29269,N_28791,N_28745);
or U29270 (N_29270,N_28540,N_28969);
nand U29271 (N_29271,N_28732,N_28227);
or U29272 (N_29272,N_28418,N_28030);
or U29273 (N_29273,N_28051,N_28234);
nand U29274 (N_29274,N_28583,N_28652);
nor U29275 (N_29275,N_28325,N_28673);
xor U29276 (N_29276,N_28678,N_28005);
xor U29277 (N_29277,N_28448,N_28463);
xnor U29278 (N_29278,N_28609,N_28975);
xor U29279 (N_29279,N_28491,N_28106);
or U29280 (N_29280,N_28009,N_28039);
and U29281 (N_29281,N_28928,N_28443);
or U29282 (N_29282,N_28002,N_28823);
nand U29283 (N_29283,N_28352,N_28371);
or U29284 (N_29284,N_28802,N_28866);
or U29285 (N_29285,N_28366,N_28862);
or U29286 (N_29286,N_28929,N_28437);
and U29287 (N_29287,N_28579,N_28324);
nand U29288 (N_29288,N_28923,N_28825);
or U29289 (N_29289,N_28080,N_28411);
and U29290 (N_29290,N_28676,N_28628);
xnor U29291 (N_29291,N_28614,N_28261);
nand U29292 (N_29292,N_28713,N_28257);
and U29293 (N_29293,N_28546,N_28603);
nand U29294 (N_29294,N_28878,N_28777);
nand U29295 (N_29295,N_28810,N_28893);
and U29296 (N_29296,N_28146,N_28993);
nor U29297 (N_29297,N_28035,N_28778);
and U29298 (N_29298,N_28350,N_28165);
nor U29299 (N_29299,N_28256,N_28223);
nor U29300 (N_29300,N_28774,N_28863);
nand U29301 (N_29301,N_28656,N_28269);
nor U29302 (N_29302,N_28727,N_28400);
nand U29303 (N_29303,N_28017,N_28959);
or U29304 (N_29304,N_28386,N_28361);
nand U29305 (N_29305,N_28309,N_28924);
or U29306 (N_29306,N_28043,N_28927);
xnor U29307 (N_29307,N_28587,N_28294);
nor U29308 (N_29308,N_28607,N_28936);
and U29309 (N_29309,N_28328,N_28719);
nand U29310 (N_29310,N_28398,N_28173);
and U29311 (N_29311,N_28763,N_28539);
or U29312 (N_29312,N_28570,N_28725);
xor U29313 (N_29313,N_28584,N_28871);
nor U29314 (N_29314,N_28586,N_28643);
nor U29315 (N_29315,N_28895,N_28942);
nand U29316 (N_29316,N_28250,N_28582);
nor U29317 (N_29317,N_28762,N_28191);
or U29318 (N_29318,N_28521,N_28974);
nand U29319 (N_29319,N_28784,N_28026);
nand U29320 (N_29320,N_28296,N_28758);
nor U29321 (N_29321,N_28378,N_28985);
and U29322 (N_29322,N_28387,N_28864);
and U29323 (N_29323,N_28248,N_28224);
and U29324 (N_29324,N_28094,N_28801);
nand U29325 (N_29325,N_28480,N_28164);
xnor U29326 (N_29326,N_28844,N_28743);
xor U29327 (N_29327,N_28861,N_28569);
or U29328 (N_29328,N_28749,N_28723);
nor U29329 (N_29329,N_28326,N_28015);
and U29330 (N_29330,N_28066,N_28595);
or U29331 (N_29331,N_28336,N_28594);
xnor U29332 (N_29332,N_28471,N_28883);
nand U29333 (N_29333,N_28376,N_28935);
nor U29334 (N_29334,N_28960,N_28060);
xnor U29335 (N_29335,N_28746,N_28696);
or U29336 (N_29336,N_28812,N_28141);
xnor U29337 (N_29337,N_28859,N_28029);
xor U29338 (N_29338,N_28076,N_28263);
nand U29339 (N_29339,N_28466,N_28254);
nand U29340 (N_29340,N_28211,N_28289);
nand U29341 (N_29341,N_28207,N_28228);
nor U29342 (N_29342,N_28990,N_28340);
nor U29343 (N_29343,N_28813,N_28128);
nand U29344 (N_29344,N_28465,N_28623);
xor U29345 (N_29345,N_28523,N_28786);
and U29346 (N_29346,N_28195,N_28653);
and U29347 (N_29347,N_28091,N_28601);
and U29348 (N_29348,N_28632,N_28922);
nor U29349 (N_29349,N_28226,N_28967);
nor U29350 (N_29350,N_28295,N_28012);
and U29351 (N_29351,N_28641,N_28909);
or U29352 (N_29352,N_28218,N_28110);
xnor U29353 (N_29353,N_28343,N_28752);
nand U29354 (N_29354,N_28286,N_28683);
nand U29355 (N_29355,N_28216,N_28127);
xnor U29356 (N_29356,N_28079,N_28671);
nand U29357 (N_29357,N_28606,N_28170);
or U29358 (N_29358,N_28695,N_28318);
nand U29359 (N_29359,N_28514,N_28461);
or U29360 (N_29360,N_28375,N_28200);
xor U29361 (N_29361,N_28613,N_28310);
or U29362 (N_29362,N_28757,N_28724);
xnor U29363 (N_29363,N_28576,N_28055);
nand U29364 (N_29364,N_28399,N_28706);
and U29365 (N_29365,N_28262,N_28246);
nor U29366 (N_29366,N_28604,N_28284);
and U29367 (N_29367,N_28071,N_28767);
or U29368 (N_29368,N_28192,N_28832);
xnor U29369 (N_29369,N_28872,N_28664);
or U29370 (N_29370,N_28022,N_28359);
and U29371 (N_29371,N_28495,N_28685);
nor U29372 (N_29372,N_28809,N_28589);
or U29373 (N_29373,N_28137,N_28247);
nor U29374 (N_29374,N_28726,N_28161);
and U29375 (N_29375,N_28130,N_28665);
nor U29376 (N_29376,N_28135,N_28704);
nor U29377 (N_29377,N_28327,N_28559);
and U29378 (N_29378,N_28126,N_28484);
and U29379 (N_29379,N_28253,N_28646);
xnor U29380 (N_29380,N_28102,N_28682);
or U29381 (N_29381,N_28099,N_28780);
and U29382 (N_29382,N_28686,N_28033);
nor U29383 (N_29383,N_28016,N_28775);
xnor U29384 (N_29384,N_28807,N_28385);
xor U29385 (N_29385,N_28741,N_28092);
nor U29386 (N_29386,N_28496,N_28751);
xnor U29387 (N_29387,N_28649,N_28474);
nand U29388 (N_29388,N_28302,N_28666);
or U29389 (N_29389,N_28333,N_28093);
and U29390 (N_29390,N_28538,N_28428);
xnor U29391 (N_29391,N_28331,N_28279);
nand U29392 (N_29392,N_28970,N_28488);
nor U29393 (N_29393,N_28873,N_28027);
nor U29394 (N_29394,N_28360,N_28951);
nand U29395 (N_29395,N_28503,N_28769);
and U29396 (N_29396,N_28349,N_28063);
nand U29397 (N_29397,N_28674,N_28519);
nand U29398 (N_29398,N_28518,N_28056);
and U29399 (N_29399,N_28186,N_28255);
or U29400 (N_29400,N_28742,N_28899);
and U29401 (N_29401,N_28941,N_28104);
and U29402 (N_29402,N_28180,N_28698);
xor U29403 (N_29403,N_28133,N_28857);
nand U29404 (N_29404,N_28747,N_28177);
nand U29405 (N_29405,N_28036,N_28444);
or U29406 (N_29406,N_28003,N_28467);
and U29407 (N_29407,N_28889,N_28075);
nand U29408 (N_29408,N_28779,N_28733);
nand U29409 (N_29409,N_28054,N_28867);
nand U29410 (N_29410,N_28215,N_28206);
xnor U29411 (N_29411,N_28847,N_28946);
or U29412 (N_29412,N_28446,N_28795);
and U29413 (N_29413,N_28849,N_28070);
nor U29414 (N_29414,N_28172,N_28648);
nor U29415 (N_29415,N_28739,N_28264);
or U29416 (N_29416,N_28213,N_28201);
nor U29417 (N_29417,N_28419,N_28943);
nand U29418 (N_29418,N_28167,N_28382);
or U29419 (N_29419,N_28557,N_28886);
xor U29420 (N_29420,N_28194,N_28470);
and U29421 (N_29421,N_28699,N_28335);
and U29422 (N_29422,N_28367,N_28049);
and U29423 (N_29423,N_28945,N_28169);
and U29424 (N_29424,N_28921,N_28817);
and U29425 (N_29425,N_28785,N_28330);
xor U29426 (N_29426,N_28401,N_28834);
nor U29427 (N_29427,N_28153,N_28958);
nor U29428 (N_29428,N_28508,N_28183);
or U29429 (N_29429,N_28900,N_28184);
and U29430 (N_29430,N_28592,N_28545);
nand U29431 (N_29431,N_28281,N_28913);
and U29432 (N_29432,N_28621,N_28618);
or U29433 (N_29433,N_28405,N_28845);
nand U29434 (N_29434,N_28855,N_28705);
or U29435 (N_29435,N_28535,N_28992);
xor U29436 (N_29436,N_28555,N_28736);
nand U29437 (N_29437,N_28635,N_28451);
or U29438 (N_29438,N_28038,N_28189);
nand U29439 (N_29439,N_28116,N_28095);
nor U29440 (N_29440,N_28083,N_28406);
nor U29441 (N_29441,N_28010,N_28276);
xnor U29442 (N_29442,N_28994,N_28416);
and U29443 (N_29443,N_28824,N_28329);
and U29444 (N_29444,N_28494,N_28282);
nor U29445 (N_29445,N_28258,N_28412);
or U29446 (N_29446,N_28955,N_28753);
and U29447 (N_29447,N_28634,N_28357);
nor U29448 (N_29448,N_28691,N_28522);
or U29449 (N_29449,N_28477,N_28911);
nand U29450 (N_29450,N_28482,N_28143);
nor U29451 (N_29451,N_28244,N_28819);
xnor U29452 (N_29452,N_28249,N_28963);
nand U29453 (N_29453,N_28957,N_28668);
nand U29454 (N_29454,N_28311,N_28773);
and U29455 (N_29455,N_28831,N_28020);
nor U29456 (N_29456,N_28980,N_28562);
xor U29457 (N_29457,N_28764,N_28356);
xor U29458 (N_29458,N_28534,N_28483);
nand U29459 (N_29459,N_28068,N_28497);
xor U29460 (N_29460,N_28273,N_28084);
or U29461 (N_29461,N_28568,N_28894);
nor U29462 (N_29462,N_28930,N_28836);
nand U29463 (N_29463,N_28776,N_28151);
and U29464 (N_29464,N_28346,N_28541);
nand U29465 (N_29465,N_28573,N_28631);
and U29466 (N_29466,N_28149,N_28421);
nand U29467 (N_29467,N_28440,N_28558);
and U29468 (N_29468,N_28636,N_28334);
xor U29469 (N_29469,N_28875,N_28456);
or U29470 (N_29470,N_28395,N_28004);
or U29471 (N_29471,N_28550,N_28735);
xor U29472 (N_29472,N_28077,N_28693);
nand U29473 (N_29473,N_28808,N_28976);
nand U29474 (N_29474,N_28314,N_28708);
nand U29475 (N_29475,N_28561,N_28760);
nor U29476 (N_29476,N_28669,N_28219);
and U29477 (N_29477,N_28225,N_28454);
nand U29478 (N_29478,N_28675,N_28548);
xor U29479 (N_29479,N_28097,N_28424);
or U29480 (N_29480,N_28090,N_28397);
xnor U29481 (N_29481,N_28940,N_28890);
and U29482 (N_29482,N_28707,N_28526);
or U29483 (N_29483,N_28744,N_28999);
nor U29484 (N_29484,N_28734,N_28157);
and U29485 (N_29485,N_28633,N_28717);
xnor U29486 (N_29486,N_28007,N_28513);
and U29487 (N_29487,N_28229,N_28916);
or U29488 (N_29488,N_28354,N_28024);
nor U29489 (N_29489,N_28347,N_28230);
and U29490 (N_29490,N_28850,N_28952);
nor U29491 (N_29491,N_28506,N_28363);
nand U29492 (N_29492,N_28789,N_28044);
xnor U29493 (N_29493,N_28233,N_28658);
or U29494 (N_29494,N_28222,N_28737);
and U29495 (N_29495,N_28950,N_28362);
nor U29496 (N_29496,N_28028,N_28731);
xor U29497 (N_29497,N_28600,N_28630);
nand U29498 (N_29498,N_28544,N_28591);
nand U29499 (N_29499,N_28119,N_28903);
xor U29500 (N_29500,N_28480,N_28750);
nor U29501 (N_29501,N_28429,N_28542);
nor U29502 (N_29502,N_28671,N_28838);
nor U29503 (N_29503,N_28892,N_28946);
xor U29504 (N_29504,N_28594,N_28212);
or U29505 (N_29505,N_28890,N_28685);
or U29506 (N_29506,N_28911,N_28589);
xnor U29507 (N_29507,N_28956,N_28458);
xnor U29508 (N_29508,N_28145,N_28442);
and U29509 (N_29509,N_28246,N_28311);
xor U29510 (N_29510,N_28265,N_28477);
and U29511 (N_29511,N_28112,N_28771);
nand U29512 (N_29512,N_28677,N_28653);
and U29513 (N_29513,N_28883,N_28840);
and U29514 (N_29514,N_28404,N_28556);
or U29515 (N_29515,N_28936,N_28352);
or U29516 (N_29516,N_28368,N_28299);
and U29517 (N_29517,N_28583,N_28844);
and U29518 (N_29518,N_28671,N_28827);
nand U29519 (N_29519,N_28702,N_28460);
nand U29520 (N_29520,N_28646,N_28748);
xor U29521 (N_29521,N_28873,N_28115);
xnor U29522 (N_29522,N_28638,N_28110);
or U29523 (N_29523,N_28391,N_28317);
nand U29524 (N_29524,N_28753,N_28399);
xnor U29525 (N_29525,N_28141,N_28765);
nand U29526 (N_29526,N_28182,N_28381);
nand U29527 (N_29527,N_28321,N_28872);
nor U29528 (N_29528,N_28661,N_28508);
xnor U29529 (N_29529,N_28975,N_28121);
or U29530 (N_29530,N_28350,N_28041);
nand U29531 (N_29531,N_28260,N_28226);
nor U29532 (N_29532,N_28603,N_28071);
and U29533 (N_29533,N_28692,N_28542);
nor U29534 (N_29534,N_28042,N_28159);
nand U29535 (N_29535,N_28658,N_28758);
and U29536 (N_29536,N_28593,N_28179);
xnor U29537 (N_29537,N_28013,N_28662);
xor U29538 (N_29538,N_28053,N_28847);
xor U29539 (N_29539,N_28634,N_28005);
nor U29540 (N_29540,N_28246,N_28039);
or U29541 (N_29541,N_28957,N_28615);
nand U29542 (N_29542,N_28086,N_28774);
and U29543 (N_29543,N_28534,N_28790);
or U29544 (N_29544,N_28165,N_28392);
nand U29545 (N_29545,N_28458,N_28856);
nor U29546 (N_29546,N_28003,N_28363);
nand U29547 (N_29547,N_28716,N_28074);
and U29548 (N_29548,N_28423,N_28233);
xnor U29549 (N_29549,N_28263,N_28281);
and U29550 (N_29550,N_28476,N_28502);
nand U29551 (N_29551,N_28437,N_28906);
nor U29552 (N_29552,N_28302,N_28931);
and U29553 (N_29553,N_28590,N_28866);
nand U29554 (N_29554,N_28366,N_28474);
or U29555 (N_29555,N_28420,N_28932);
xnor U29556 (N_29556,N_28003,N_28021);
and U29557 (N_29557,N_28077,N_28639);
nor U29558 (N_29558,N_28887,N_28318);
nor U29559 (N_29559,N_28086,N_28165);
or U29560 (N_29560,N_28023,N_28071);
nor U29561 (N_29561,N_28716,N_28824);
xor U29562 (N_29562,N_28770,N_28570);
nor U29563 (N_29563,N_28180,N_28399);
nand U29564 (N_29564,N_28536,N_28458);
xor U29565 (N_29565,N_28739,N_28827);
xnor U29566 (N_29566,N_28425,N_28644);
or U29567 (N_29567,N_28426,N_28060);
and U29568 (N_29568,N_28337,N_28449);
xor U29569 (N_29569,N_28134,N_28827);
nor U29570 (N_29570,N_28463,N_28745);
nor U29571 (N_29571,N_28570,N_28698);
xor U29572 (N_29572,N_28516,N_28970);
or U29573 (N_29573,N_28453,N_28892);
or U29574 (N_29574,N_28483,N_28498);
xor U29575 (N_29575,N_28593,N_28394);
and U29576 (N_29576,N_28977,N_28404);
and U29577 (N_29577,N_28413,N_28132);
xnor U29578 (N_29578,N_28810,N_28497);
xor U29579 (N_29579,N_28789,N_28549);
and U29580 (N_29580,N_28789,N_28839);
xor U29581 (N_29581,N_28554,N_28213);
nand U29582 (N_29582,N_28996,N_28630);
xor U29583 (N_29583,N_28596,N_28325);
and U29584 (N_29584,N_28291,N_28506);
xor U29585 (N_29585,N_28533,N_28191);
xor U29586 (N_29586,N_28680,N_28052);
xnor U29587 (N_29587,N_28728,N_28919);
or U29588 (N_29588,N_28478,N_28798);
or U29589 (N_29589,N_28580,N_28570);
xnor U29590 (N_29590,N_28155,N_28105);
xnor U29591 (N_29591,N_28054,N_28298);
nand U29592 (N_29592,N_28045,N_28617);
or U29593 (N_29593,N_28542,N_28972);
nand U29594 (N_29594,N_28881,N_28161);
nor U29595 (N_29595,N_28652,N_28284);
xnor U29596 (N_29596,N_28121,N_28510);
xor U29597 (N_29597,N_28821,N_28880);
or U29598 (N_29598,N_28393,N_28167);
or U29599 (N_29599,N_28867,N_28153);
xnor U29600 (N_29600,N_28684,N_28695);
or U29601 (N_29601,N_28220,N_28638);
nand U29602 (N_29602,N_28805,N_28315);
nor U29603 (N_29603,N_28753,N_28165);
and U29604 (N_29604,N_28978,N_28245);
nand U29605 (N_29605,N_28390,N_28689);
xor U29606 (N_29606,N_28862,N_28992);
or U29607 (N_29607,N_28726,N_28942);
nor U29608 (N_29608,N_28696,N_28567);
xor U29609 (N_29609,N_28505,N_28400);
and U29610 (N_29610,N_28220,N_28065);
and U29611 (N_29611,N_28569,N_28926);
nor U29612 (N_29612,N_28421,N_28697);
or U29613 (N_29613,N_28292,N_28795);
xnor U29614 (N_29614,N_28795,N_28876);
and U29615 (N_29615,N_28721,N_28015);
xor U29616 (N_29616,N_28893,N_28204);
nor U29617 (N_29617,N_28939,N_28648);
xnor U29618 (N_29618,N_28693,N_28469);
xnor U29619 (N_29619,N_28198,N_28751);
or U29620 (N_29620,N_28487,N_28610);
or U29621 (N_29621,N_28275,N_28096);
and U29622 (N_29622,N_28192,N_28264);
xnor U29623 (N_29623,N_28491,N_28319);
nand U29624 (N_29624,N_28807,N_28084);
nor U29625 (N_29625,N_28647,N_28333);
xnor U29626 (N_29626,N_28103,N_28230);
xnor U29627 (N_29627,N_28701,N_28120);
nand U29628 (N_29628,N_28504,N_28811);
or U29629 (N_29629,N_28551,N_28948);
or U29630 (N_29630,N_28452,N_28397);
nand U29631 (N_29631,N_28397,N_28189);
nor U29632 (N_29632,N_28629,N_28861);
and U29633 (N_29633,N_28267,N_28964);
nor U29634 (N_29634,N_28670,N_28206);
nand U29635 (N_29635,N_28000,N_28073);
nor U29636 (N_29636,N_28514,N_28664);
xnor U29637 (N_29637,N_28188,N_28554);
or U29638 (N_29638,N_28710,N_28757);
xor U29639 (N_29639,N_28222,N_28949);
xnor U29640 (N_29640,N_28854,N_28621);
nor U29641 (N_29641,N_28598,N_28087);
xor U29642 (N_29642,N_28815,N_28406);
and U29643 (N_29643,N_28676,N_28340);
xor U29644 (N_29644,N_28787,N_28093);
nor U29645 (N_29645,N_28816,N_28567);
nand U29646 (N_29646,N_28577,N_28745);
xor U29647 (N_29647,N_28977,N_28097);
nor U29648 (N_29648,N_28792,N_28482);
nand U29649 (N_29649,N_28710,N_28803);
or U29650 (N_29650,N_28832,N_28699);
or U29651 (N_29651,N_28615,N_28238);
xnor U29652 (N_29652,N_28583,N_28969);
and U29653 (N_29653,N_28563,N_28674);
nor U29654 (N_29654,N_28640,N_28509);
nand U29655 (N_29655,N_28101,N_28357);
nor U29656 (N_29656,N_28496,N_28670);
nand U29657 (N_29657,N_28738,N_28640);
xor U29658 (N_29658,N_28574,N_28771);
xnor U29659 (N_29659,N_28721,N_28616);
and U29660 (N_29660,N_28096,N_28601);
xnor U29661 (N_29661,N_28333,N_28659);
xor U29662 (N_29662,N_28487,N_28449);
and U29663 (N_29663,N_28426,N_28748);
nor U29664 (N_29664,N_28772,N_28193);
nand U29665 (N_29665,N_28906,N_28715);
or U29666 (N_29666,N_28448,N_28291);
xor U29667 (N_29667,N_28933,N_28028);
or U29668 (N_29668,N_28559,N_28226);
or U29669 (N_29669,N_28633,N_28454);
xor U29670 (N_29670,N_28441,N_28215);
or U29671 (N_29671,N_28653,N_28358);
nand U29672 (N_29672,N_28462,N_28726);
and U29673 (N_29673,N_28480,N_28583);
and U29674 (N_29674,N_28348,N_28516);
nor U29675 (N_29675,N_28034,N_28447);
xnor U29676 (N_29676,N_28276,N_28945);
nand U29677 (N_29677,N_28193,N_28879);
nor U29678 (N_29678,N_28404,N_28107);
and U29679 (N_29679,N_28165,N_28035);
and U29680 (N_29680,N_28704,N_28747);
and U29681 (N_29681,N_28025,N_28270);
xnor U29682 (N_29682,N_28754,N_28350);
nor U29683 (N_29683,N_28148,N_28569);
and U29684 (N_29684,N_28797,N_28694);
nand U29685 (N_29685,N_28882,N_28224);
and U29686 (N_29686,N_28017,N_28123);
or U29687 (N_29687,N_28712,N_28721);
xor U29688 (N_29688,N_28554,N_28079);
and U29689 (N_29689,N_28807,N_28487);
xor U29690 (N_29690,N_28210,N_28109);
nor U29691 (N_29691,N_28377,N_28359);
xnor U29692 (N_29692,N_28319,N_28266);
and U29693 (N_29693,N_28768,N_28038);
or U29694 (N_29694,N_28621,N_28797);
xor U29695 (N_29695,N_28293,N_28594);
and U29696 (N_29696,N_28373,N_28101);
xnor U29697 (N_29697,N_28465,N_28092);
or U29698 (N_29698,N_28442,N_28781);
xnor U29699 (N_29699,N_28351,N_28323);
or U29700 (N_29700,N_28743,N_28726);
and U29701 (N_29701,N_28177,N_28106);
xnor U29702 (N_29702,N_28431,N_28715);
nand U29703 (N_29703,N_28235,N_28527);
nor U29704 (N_29704,N_28515,N_28032);
xnor U29705 (N_29705,N_28688,N_28116);
or U29706 (N_29706,N_28555,N_28696);
nand U29707 (N_29707,N_28309,N_28427);
nand U29708 (N_29708,N_28010,N_28579);
or U29709 (N_29709,N_28830,N_28584);
or U29710 (N_29710,N_28812,N_28923);
nand U29711 (N_29711,N_28603,N_28340);
xor U29712 (N_29712,N_28246,N_28959);
nand U29713 (N_29713,N_28027,N_28522);
xor U29714 (N_29714,N_28255,N_28924);
or U29715 (N_29715,N_28238,N_28953);
and U29716 (N_29716,N_28465,N_28299);
nor U29717 (N_29717,N_28293,N_28454);
nor U29718 (N_29718,N_28114,N_28155);
and U29719 (N_29719,N_28377,N_28861);
nor U29720 (N_29720,N_28088,N_28337);
and U29721 (N_29721,N_28778,N_28542);
xor U29722 (N_29722,N_28153,N_28616);
nor U29723 (N_29723,N_28845,N_28523);
nand U29724 (N_29724,N_28646,N_28875);
xnor U29725 (N_29725,N_28304,N_28206);
xnor U29726 (N_29726,N_28854,N_28532);
and U29727 (N_29727,N_28501,N_28751);
and U29728 (N_29728,N_28903,N_28136);
nor U29729 (N_29729,N_28713,N_28533);
nor U29730 (N_29730,N_28889,N_28723);
or U29731 (N_29731,N_28942,N_28826);
and U29732 (N_29732,N_28622,N_28387);
and U29733 (N_29733,N_28636,N_28009);
nor U29734 (N_29734,N_28421,N_28453);
or U29735 (N_29735,N_28846,N_28981);
nand U29736 (N_29736,N_28796,N_28526);
nand U29737 (N_29737,N_28762,N_28857);
and U29738 (N_29738,N_28510,N_28981);
nor U29739 (N_29739,N_28482,N_28287);
nor U29740 (N_29740,N_28552,N_28021);
or U29741 (N_29741,N_28421,N_28816);
and U29742 (N_29742,N_28535,N_28362);
and U29743 (N_29743,N_28315,N_28561);
and U29744 (N_29744,N_28145,N_28794);
nand U29745 (N_29745,N_28442,N_28494);
nand U29746 (N_29746,N_28221,N_28758);
and U29747 (N_29747,N_28817,N_28449);
or U29748 (N_29748,N_28938,N_28304);
or U29749 (N_29749,N_28007,N_28987);
xor U29750 (N_29750,N_28772,N_28426);
nand U29751 (N_29751,N_28934,N_28292);
nor U29752 (N_29752,N_28645,N_28427);
xor U29753 (N_29753,N_28264,N_28141);
or U29754 (N_29754,N_28070,N_28280);
or U29755 (N_29755,N_28254,N_28686);
nand U29756 (N_29756,N_28949,N_28725);
nor U29757 (N_29757,N_28410,N_28465);
and U29758 (N_29758,N_28046,N_28755);
xor U29759 (N_29759,N_28982,N_28100);
or U29760 (N_29760,N_28484,N_28339);
or U29761 (N_29761,N_28787,N_28538);
nand U29762 (N_29762,N_28843,N_28146);
nand U29763 (N_29763,N_28622,N_28495);
xnor U29764 (N_29764,N_28295,N_28527);
and U29765 (N_29765,N_28872,N_28216);
xnor U29766 (N_29766,N_28078,N_28558);
xnor U29767 (N_29767,N_28309,N_28200);
nor U29768 (N_29768,N_28013,N_28343);
and U29769 (N_29769,N_28432,N_28565);
nor U29770 (N_29770,N_28941,N_28244);
and U29771 (N_29771,N_28946,N_28820);
nor U29772 (N_29772,N_28124,N_28563);
xor U29773 (N_29773,N_28917,N_28079);
nand U29774 (N_29774,N_28194,N_28031);
nand U29775 (N_29775,N_28704,N_28972);
nand U29776 (N_29776,N_28513,N_28036);
nand U29777 (N_29777,N_28404,N_28602);
or U29778 (N_29778,N_28219,N_28003);
nand U29779 (N_29779,N_28624,N_28410);
and U29780 (N_29780,N_28079,N_28022);
nor U29781 (N_29781,N_28848,N_28176);
nor U29782 (N_29782,N_28152,N_28077);
and U29783 (N_29783,N_28999,N_28926);
xor U29784 (N_29784,N_28724,N_28424);
nand U29785 (N_29785,N_28461,N_28909);
or U29786 (N_29786,N_28621,N_28693);
nand U29787 (N_29787,N_28975,N_28057);
nor U29788 (N_29788,N_28570,N_28344);
and U29789 (N_29789,N_28267,N_28330);
nand U29790 (N_29790,N_28890,N_28561);
xor U29791 (N_29791,N_28571,N_28244);
and U29792 (N_29792,N_28901,N_28836);
nor U29793 (N_29793,N_28263,N_28536);
xor U29794 (N_29794,N_28589,N_28064);
or U29795 (N_29795,N_28257,N_28443);
or U29796 (N_29796,N_28151,N_28407);
nand U29797 (N_29797,N_28084,N_28523);
and U29798 (N_29798,N_28798,N_28519);
nand U29799 (N_29799,N_28438,N_28726);
and U29800 (N_29800,N_28122,N_28979);
nor U29801 (N_29801,N_28538,N_28166);
xor U29802 (N_29802,N_28827,N_28500);
and U29803 (N_29803,N_28052,N_28345);
or U29804 (N_29804,N_28971,N_28291);
xnor U29805 (N_29805,N_28681,N_28278);
and U29806 (N_29806,N_28891,N_28896);
and U29807 (N_29807,N_28923,N_28481);
or U29808 (N_29808,N_28749,N_28060);
and U29809 (N_29809,N_28271,N_28911);
nand U29810 (N_29810,N_28679,N_28481);
xnor U29811 (N_29811,N_28293,N_28829);
xnor U29812 (N_29812,N_28184,N_28252);
nor U29813 (N_29813,N_28056,N_28226);
nand U29814 (N_29814,N_28435,N_28456);
xnor U29815 (N_29815,N_28705,N_28716);
or U29816 (N_29816,N_28517,N_28443);
and U29817 (N_29817,N_28110,N_28697);
and U29818 (N_29818,N_28139,N_28961);
or U29819 (N_29819,N_28833,N_28074);
xnor U29820 (N_29820,N_28528,N_28350);
or U29821 (N_29821,N_28558,N_28377);
nor U29822 (N_29822,N_28676,N_28493);
or U29823 (N_29823,N_28679,N_28274);
or U29824 (N_29824,N_28255,N_28028);
or U29825 (N_29825,N_28725,N_28921);
xnor U29826 (N_29826,N_28246,N_28965);
nand U29827 (N_29827,N_28629,N_28029);
xor U29828 (N_29828,N_28186,N_28789);
nand U29829 (N_29829,N_28448,N_28662);
xnor U29830 (N_29830,N_28876,N_28787);
or U29831 (N_29831,N_28840,N_28408);
or U29832 (N_29832,N_28692,N_28002);
or U29833 (N_29833,N_28304,N_28411);
or U29834 (N_29834,N_28828,N_28312);
and U29835 (N_29835,N_28146,N_28072);
nor U29836 (N_29836,N_28269,N_28377);
or U29837 (N_29837,N_28747,N_28732);
nor U29838 (N_29838,N_28964,N_28647);
nand U29839 (N_29839,N_28371,N_28874);
or U29840 (N_29840,N_28758,N_28472);
xor U29841 (N_29841,N_28624,N_28376);
nor U29842 (N_29842,N_28747,N_28491);
nor U29843 (N_29843,N_28242,N_28179);
nor U29844 (N_29844,N_28757,N_28883);
and U29845 (N_29845,N_28007,N_28907);
or U29846 (N_29846,N_28269,N_28327);
nand U29847 (N_29847,N_28735,N_28905);
nand U29848 (N_29848,N_28628,N_28456);
and U29849 (N_29849,N_28932,N_28794);
nand U29850 (N_29850,N_28382,N_28159);
and U29851 (N_29851,N_28204,N_28116);
nand U29852 (N_29852,N_28611,N_28568);
or U29853 (N_29853,N_28339,N_28734);
nor U29854 (N_29854,N_28231,N_28368);
nand U29855 (N_29855,N_28654,N_28792);
nand U29856 (N_29856,N_28137,N_28650);
xnor U29857 (N_29857,N_28975,N_28474);
xor U29858 (N_29858,N_28264,N_28786);
nor U29859 (N_29859,N_28853,N_28288);
nand U29860 (N_29860,N_28896,N_28139);
nand U29861 (N_29861,N_28694,N_28002);
nand U29862 (N_29862,N_28293,N_28984);
xor U29863 (N_29863,N_28021,N_28329);
and U29864 (N_29864,N_28707,N_28778);
xor U29865 (N_29865,N_28210,N_28182);
and U29866 (N_29866,N_28706,N_28123);
xnor U29867 (N_29867,N_28415,N_28493);
nand U29868 (N_29868,N_28754,N_28676);
nor U29869 (N_29869,N_28043,N_28229);
nand U29870 (N_29870,N_28889,N_28090);
and U29871 (N_29871,N_28034,N_28535);
nor U29872 (N_29872,N_28350,N_28914);
and U29873 (N_29873,N_28979,N_28085);
nor U29874 (N_29874,N_28226,N_28981);
xor U29875 (N_29875,N_28983,N_28210);
or U29876 (N_29876,N_28366,N_28391);
nand U29877 (N_29877,N_28331,N_28465);
or U29878 (N_29878,N_28227,N_28391);
and U29879 (N_29879,N_28164,N_28525);
nor U29880 (N_29880,N_28498,N_28249);
or U29881 (N_29881,N_28319,N_28540);
or U29882 (N_29882,N_28931,N_28848);
or U29883 (N_29883,N_28125,N_28713);
xor U29884 (N_29884,N_28609,N_28591);
nor U29885 (N_29885,N_28574,N_28036);
xnor U29886 (N_29886,N_28582,N_28893);
nand U29887 (N_29887,N_28167,N_28724);
and U29888 (N_29888,N_28412,N_28937);
xor U29889 (N_29889,N_28226,N_28854);
nand U29890 (N_29890,N_28945,N_28413);
nor U29891 (N_29891,N_28369,N_28393);
or U29892 (N_29892,N_28137,N_28951);
or U29893 (N_29893,N_28094,N_28519);
nor U29894 (N_29894,N_28002,N_28656);
nand U29895 (N_29895,N_28361,N_28595);
and U29896 (N_29896,N_28046,N_28214);
xnor U29897 (N_29897,N_28717,N_28349);
or U29898 (N_29898,N_28485,N_28628);
nand U29899 (N_29899,N_28585,N_28241);
and U29900 (N_29900,N_28913,N_28310);
nor U29901 (N_29901,N_28106,N_28303);
nor U29902 (N_29902,N_28697,N_28160);
xnor U29903 (N_29903,N_28017,N_28121);
and U29904 (N_29904,N_28625,N_28407);
or U29905 (N_29905,N_28598,N_28060);
or U29906 (N_29906,N_28931,N_28542);
or U29907 (N_29907,N_28456,N_28198);
or U29908 (N_29908,N_28323,N_28009);
nor U29909 (N_29909,N_28184,N_28587);
and U29910 (N_29910,N_28082,N_28040);
nor U29911 (N_29911,N_28613,N_28210);
or U29912 (N_29912,N_28133,N_28936);
or U29913 (N_29913,N_28849,N_28152);
xnor U29914 (N_29914,N_28113,N_28813);
xnor U29915 (N_29915,N_28926,N_28618);
nor U29916 (N_29916,N_28856,N_28813);
nor U29917 (N_29917,N_28155,N_28273);
nand U29918 (N_29918,N_28661,N_28705);
and U29919 (N_29919,N_28553,N_28353);
or U29920 (N_29920,N_28690,N_28480);
xor U29921 (N_29921,N_28860,N_28831);
and U29922 (N_29922,N_28642,N_28922);
or U29923 (N_29923,N_28212,N_28630);
nor U29924 (N_29924,N_28128,N_28924);
nand U29925 (N_29925,N_28242,N_28607);
nand U29926 (N_29926,N_28842,N_28340);
nand U29927 (N_29927,N_28714,N_28584);
nand U29928 (N_29928,N_28364,N_28156);
nor U29929 (N_29929,N_28751,N_28459);
and U29930 (N_29930,N_28260,N_28210);
nor U29931 (N_29931,N_28281,N_28559);
xnor U29932 (N_29932,N_28904,N_28209);
nor U29933 (N_29933,N_28688,N_28702);
xor U29934 (N_29934,N_28021,N_28082);
or U29935 (N_29935,N_28936,N_28802);
xor U29936 (N_29936,N_28949,N_28900);
nand U29937 (N_29937,N_28085,N_28186);
or U29938 (N_29938,N_28681,N_28422);
xor U29939 (N_29939,N_28531,N_28302);
nor U29940 (N_29940,N_28954,N_28204);
or U29941 (N_29941,N_28392,N_28267);
or U29942 (N_29942,N_28545,N_28429);
and U29943 (N_29943,N_28356,N_28671);
and U29944 (N_29944,N_28436,N_28764);
or U29945 (N_29945,N_28229,N_28226);
nor U29946 (N_29946,N_28551,N_28621);
or U29947 (N_29947,N_28361,N_28039);
or U29948 (N_29948,N_28997,N_28699);
nor U29949 (N_29949,N_28444,N_28372);
nand U29950 (N_29950,N_28204,N_28498);
and U29951 (N_29951,N_28184,N_28632);
and U29952 (N_29952,N_28771,N_28597);
nand U29953 (N_29953,N_28166,N_28438);
nand U29954 (N_29954,N_28715,N_28515);
and U29955 (N_29955,N_28741,N_28147);
xnor U29956 (N_29956,N_28126,N_28826);
xor U29957 (N_29957,N_28232,N_28979);
and U29958 (N_29958,N_28079,N_28318);
and U29959 (N_29959,N_28875,N_28823);
nand U29960 (N_29960,N_28659,N_28174);
or U29961 (N_29961,N_28802,N_28856);
or U29962 (N_29962,N_28673,N_28049);
nor U29963 (N_29963,N_28867,N_28443);
and U29964 (N_29964,N_28411,N_28316);
nand U29965 (N_29965,N_28839,N_28123);
and U29966 (N_29966,N_28127,N_28457);
nand U29967 (N_29967,N_28365,N_28505);
xor U29968 (N_29968,N_28148,N_28826);
xor U29969 (N_29969,N_28175,N_28989);
nor U29970 (N_29970,N_28848,N_28578);
nor U29971 (N_29971,N_28873,N_28270);
xor U29972 (N_29972,N_28946,N_28721);
or U29973 (N_29973,N_28127,N_28979);
and U29974 (N_29974,N_28503,N_28757);
and U29975 (N_29975,N_28374,N_28286);
or U29976 (N_29976,N_28653,N_28009);
xnor U29977 (N_29977,N_28325,N_28984);
or U29978 (N_29978,N_28472,N_28298);
and U29979 (N_29979,N_28723,N_28126);
and U29980 (N_29980,N_28129,N_28843);
xor U29981 (N_29981,N_28734,N_28992);
nand U29982 (N_29982,N_28355,N_28699);
xor U29983 (N_29983,N_28024,N_28475);
nand U29984 (N_29984,N_28458,N_28684);
or U29985 (N_29985,N_28211,N_28007);
and U29986 (N_29986,N_28481,N_28695);
or U29987 (N_29987,N_28498,N_28312);
nand U29988 (N_29988,N_28904,N_28470);
nand U29989 (N_29989,N_28082,N_28117);
and U29990 (N_29990,N_28869,N_28828);
nand U29991 (N_29991,N_28426,N_28170);
nand U29992 (N_29992,N_28171,N_28935);
and U29993 (N_29993,N_28335,N_28269);
nor U29994 (N_29994,N_28781,N_28212);
and U29995 (N_29995,N_28772,N_28655);
and U29996 (N_29996,N_28274,N_28527);
nand U29997 (N_29997,N_28484,N_28819);
xor U29998 (N_29998,N_28011,N_28398);
nor U29999 (N_29999,N_28167,N_28715);
and UO_0 (O_0,N_29751,N_29336);
nor UO_1 (O_1,N_29040,N_29168);
and UO_2 (O_2,N_29414,N_29601);
nand UO_3 (O_3,N_29779,N_29837);
nor UO_4 (O_4,N_29771,N_29720);
xor UO_5 (O_5,N_29370,N_29120);
xnor UO_6 (O_6,N_29464,N_29936);
nor UO_7 (O_7,N_29470,N_29243);
or UO_8 (O_8,N_29229,N_29160);
xor UO_9 (O_9,N_29701,N_29942);
xor UO_10 (O_10,N_29842,N_29116);
xor UO_11 (O_11,N_29871,N_29466);
nand UO_12 (O_12,N_29235,N_29798);
xor UO_13 (O_13,N_29367,N_29115);
xnor UO_14 (O_14,N_29118,N_29662);
nor UO_15 (O_15,N_29063,N_29208);
or UO_16 (O_16,N_29631,N_29223);
and UO_17 (O_17,N_29585,N_29467);
or UO_18 (O_18,N_29158,N_29179);
and UO_19 (O_19,N_29970,N_29571);
xor UO_20 (O_20,N_29524,N_29050);
and UO_21 (O_21,N_29540,N_29981);
xnor UO_22 (O_22,N_29390,N_29596);
or UO_23 (O_23,N_29422,N_29277);
nor UO_24 (O_24,N_29833,N_29226);
nor UO_25 (O_25,N_29248,N_29916);
nor UO_26 (O_26,N_29282,N_29512);
nor UO_27 (O_27,N_29971,N_29032);
or UO_28 (O_28,N_29977,N_29018);
and UO_29 (O_29,N_29508,N_29621);
or UO_30 (O_30,N_29998,N_29857);
and UO_31 (O_31,N_29748,N_29001);
or UO_32 (O_32,N_29677,N_29581);
and UO_33 (O_33,N_29537,N_29444);
nand UO_34 (O_34,N_29084,N_29093);
or UO_35 (O_35,N_29366,N_29108);
or UO_36 (O_36,N_29900,N_29325);
or UO_37 (O_37,N_29768,N_29230);
nand UO_38 (O_38,N_29427,N_29424);
nand UO_39 (O_39,N_29551,N_29385);
nand UO_40 (O_40,N_29532,N_29197);
and UO_41 (O_41,N_29559,N_29724);
nor UO_42 (O_42,N_29838,N_29345);
and UO_43 (O_43,N_29250,N_29595);
and UO_44 (O_44,N_29920,N_29496);
nor UO_45 (O_45,N_29213,N_29693);
or UO_46 (O_46,N_29755,N_29142);
xor UO_47 (O_47,N_29324,N_29156);
xnor UO_48 (O_48,N_29877,N_29059);
xor UO_49 (O_49,N_29257,N_29404);
xnor UO_50 (O_50,N_29687,N_29099);
and UO_51 (O_51,N_29828,N_29445);
nor UO_52 (O_52,N_29173,N_29354);
and UO_53 (O_53,N_29679,N_29371);
or UO_54 (O_54,N_29881,N_29456);
nand UO_55 (O_55,N_29839,N_29207);
nor UO_56 (O_56,N_29786,N_29594);
or UO_57 (O_57,N_29454,N_29525);
or UO_58 (O_58,N_29020,N_29908);
nor UO_59 (O_59,N_29265,N_29162);
or UO_60 (O_60,N_29847,N_29823);
or UO_61 (O_61,N_29752,N_29502);
or UO_62 (O_62,N_29211,N_29256);
or UO_63 (O_63,N_29038,N_29686);
xnor UO_64 (O_64,N_29025,N_29364);
nor UO_65 (O_65,N_29304,N_29562);
xor UO_66 (O_66,N_29441,N_29391);
and UO_67 (O_67,N_29004,N_29110);
xor UO_68 (O_68,N_29029,N_29107);
xnor UO_69 (O_69,N_29906,N_29696);
nor UO_70 (O_70,N_29067,N_29246);
xnor UO_71 (O_71,N_29943,N_29225);
xnor UO_72 (O_72,N_29355,N_29535);
and UO_73 (O_73,N_29474,N_29669);
nor UO_74 (O_74,N_29984,N_29937);
and UO_75 (O_75,N_29397,N_29046);
and UO_76 (O_76,N_29522,N_29593);
xor UO_77 (O_77,N_29151,N_29547);
xnor UO_78 (O_78,N_29599,N_29268);
nand UO_79 (O_79,N_29732,N_29861);
nor UO_80 (O_80,N_29335,N_29453);
nand UO_81 (O_81,N_29836,N_29255);
nand UO_82 (O_82,N_29053,N_29242);
xor UO_83 (O_83,N_29545,N_29733);
nor UO_84 (O_84,N_29281,N_29529);
nor UO_85 (O_85,N_29079,N_29017);
nor UO_86 (O_86,N_29910,N_29258);
xnor UO_87 (O_87,N_29612,N_29347);
or UO_88 (O_88,N_29015,N_29893);
nor UO_89 (O_89,N_29781,N_29448);
nor UO_90 (O_90,N_29388,N_29215);
nand UO_91 (O_91,N_29715,N_29418);
or UO_92 (O_92,N_29864,N_29756);
and UO_93 (O_93,N_29379,N_29503);
nand UO_94 (O_94,N_29539,N_29446);
nand UO_95 (O_95,N_29866,N_29629);
nand UO_96 (O_96,N_29209,N_29917);
or UO_97 (O_97,N_29430,N_29090);
nand UO_98 (O_98,N_29723,N_29420);
nor UO_99 (O_99,N_29963,N_29718);
and UO_100 (O_100,N_29504,N_29203);
xor UO_101 (O_101,N_29815,N_29238);
xnor UO_102 (O_102,N_29363,N_29523);
or UO_103 (O_103,N_29184,N_29763);
or UO_104 (O_104,N_29583,N_29003);
nor UO_105 (O_105,N_29794,N_29848);
and UO_106 (O_106,N_29966,N_29811);
and UO_107 (O_107,N_29616,N_29261);
nor UO_108 (O_108,N_29219,N_29071);
xnor UO_109 (O_109,N_29618,N_29021);
or UO_110 (O_110,N_29816,N_29873);
nor UO_111 (O_111,N_29403,N_29054);
or UO_112 (O_112,N_29055,N_29617);
nand UO_113 (O_113,N_29176,N_29514);
nor UO_114 (O_114,N_29558,N_29495);
and UO_115 (O_115,N_29125,N_29736);
nand UO_116 (O_116,N_29997,N_29401);
or UO_117 (O_117,N_29452,N_29615);
and UO_118 (O_118,N_29664,N_29267);
nand UO_119 (O_119,N_29949,N_29827);
and UO_120 (O_120,N_29510,N_29276);
xnor UO_121 (O_121,N_29309,N_29232);
xnor UO_122 (O_122,N_29331,N_29096);
and UO_123 (O_123,N_29538,N_29793);
and UO_124 (O_124,N_29518,N_29123);
and UO_125 (O_125,N_29024,N_29465);
nand UO_126 (O_126,N_29516,N_29384);
and UO_127 (O_127,N_29244,N_29252);
and UO_128 (O_128,N_29132,N_29240);
or UO_129 (O_129,N_29023,N_29249);
or UO_130 (O_130,N_29759,N_29577);
xor UO_131 (O_131,N_29925,N_29329);
nor UO_132 (O_132,N_29435,N_29515);
and UO_133 (O_133,N_29704,N_29328);
nand UO_134 (O_134,N_29402,N_29645);
xnor UO_135 (O_135,N_29620,N_29098);
nand UO_136 (O_136,N_29580,N_29554);
xor UO_137 (O_137,N_29210,N_29350);
and UO_138 (O_138,N_29883,N_29859);
or UO_139 (O_139,N_29691,N_29239);
and UO_140 (O_140,N_29819,N_29578);
and UO_141 (O_141,N_29939,N_29273);
nand UO_142 (O_142,N_29862,N_29953);
nor UO_143 (O_143,N_29305,N_29590);
and UO_144 (O_144,N_29012,N_29684);
and UO_145 (O_145,N_29668,N_29341);
or UO_146 (O_146,N_29138,N_29216);
nor UO_147 (O_147,N_29117,N_29463);
xor UO_148 (O_148,N_29542,N_29741);
nor UO_149 (O_149,N_29573,N_29202);
nor UO_150 (O_150,N_29803,N_29566);
or UO_151 (O_151,N_29043,N_29929);
xnor UO_152 (O_152,N_29564,N_29778);
nor UO_153 (O_153,N_29316,N_29673);
and UO_154 (O_154,N_29530,N_29841);
or UO_155 (O_155,N_29697,N_29365);
xor UO_156 (O_156,N_29106,N_29960);
nand UO_157 (O_157,N_29802,N_29852);
and UO_158 (O_158,N_29431,N_29163);
xnor UO_159 (O_159,N_29185,N_29392);
nor UO_160 (O_160,N_29344,N_29996);
xor UO_161 (O_161,N_29576,N_29911);
or UO_162 (O_162,N_29849,N_29806);
nor UO_163 (O_163,N_29659,N_29716);
nand UO_164 (O_164,N_29995,N_29476);
and UO_165 (O_165,N_29228,N_29818);
nor UO_166 (O_166,N_29134,N_29126);
nand UO_167 (O_167,N_29764,N_29436);
nor UO_168 (O_168,N_29956,N_29865);
and UO_169 (O_169,N_29633,N_29485);
or UO_170 (O_170,N_29245,N_29086);
nor UO_171 (O_171,N_29507,N_29892);
nand UO_172 (O_172,N_29342,N_29622);
nand UO_173 (O_173,N_29195,N_29274);
nand UO_174 (O_174,N_29993,N_29382);
and UO_175 (O_175,N_29582,N_29835);
nand UO_176 (O_176,N_29983,N_29747);
xnor UO_177 (O_177,N_29780,N_29170);
xnor UO_178 (O_178,N_29766,N_29473);
or UO_179 (O_179,N_29772,N_29863);
nor UO_180 (O_180,N_29812,N_29681);
xnor UO_181 (O_181,N_29380,N_29484);
and UO_182 (O_182,N_29076,N_29776);
nor UO_183 (O_183,N_29061,N_29520);
xor UO_184 (O_184,N_29725,N_29870);
or UO_185 (O_185,N_29413,N_29611);
xnor UO_186 (O_186,N_29307,N_29152);
nand UO_187 (O_187,N_29565,N_29682);
and UO_188 (O_188,N_29475,N_29932);
and UO_189 (O_189,N_29398,N_29019);
xnor UO_190 (O_190,N_29519,N_29703);
nand UO_191 (O_191,N_29979,N_29898);
and UO_192 (O_192,N_29005,N_29461);
nand UO_193 (O_193,N_29855,N_29770);
nand UO_194 (O_194,N_29869,N_29039);
nand UO_195 (O_195,N_29491,N_29721);
xor UO_196 (O_196,N_29395,N_29657);
and UO_197 (O_197,N_29699,N_29785);
nor UO_198 (O_198,N_29127,N_29415);
and UO_199 (O_199,N_29455,N_29320);
xnor UO_200 (O_200,N_29783,N_29407);
nand UO_201 (O_201,N_29787,N_29080);
xor UO_202 (O_202,N_29951,N_29556);
nor UO_203 (O_203,N_29130,N_29894);
nand UO_204 (O_204,N_29016,N_29899);
nand UO_205 (O_205,N_29233,N_29598);
nor UO_206 (O_206,N_29886,N_29319);
and UO_207 (O_207,N_29490,N_29136);
nand UO_208 (O_208,N_29757,N_29817);
nand UO_209 (O_209,N_29416,N_29685);
nand UO_210 (O_210,N_29891,N_29405);
xor UO_211 (O_211,N_29034,N_29710);
and UO_212 (O_212,N_29945,N_29746);
xnor UO_213 (O_213,N_29044,N_29434);
nand UO_214 (O_214,N_29178,N_29634);
and UO_215 (O_215,N_29087,N_29149);
or UO_216 (O_216,N_29042,N_29333);
and UO_217 (O_217,N_29650,N_29393);
nand UO_218 (O_218,N_29990,N_29978);
and UO_219 (O_219,N_29543,N_29030);
or UO_220 (O_220,N_29670,N_29935);
xnor UO_221 (O_221,N_29317,N_29613);
xor UO_222 (O_222,N_29112,N_29605);
xnor UO_223 (O_223,N_29026,N_29991);
or UO_224 (O_224,N_29440,N_29394);
or UO_225 (O_225,N_29745,N_29555);
nor UO_226 (O_226,N_29789,N_29154);
nand UO_227 (O_227,N_29389,N_29161);
and UO_228 (O_228,N_29468,N_29419);
and UO_229 (O_229,N_29070,N_29109);
nand UO_230 (O_230,N_29089,N_29726);
nor UO_231 (O_231,N_29264,N_29694);
nor UO_232 (O_232,N_29560,N_29509);
nor UO_233 (O_233,N_29101,N_29065);
nand UO_234 (O_234,N_29150,N_29334);
and UO_235 (O_235,N_29909,N_29280);
nor UO_236 (O_236,N_29078,N_29073);
nor UO_237 (O_237,N_29628,N_29064);
and UO_238 (O_238,N_29805,N_29832);
xor UO_239 (O_239,N_29563,N_29744);
or UO_240 (O_240,N_29879,N_29296);
xnor UO_241 (O_241,N_29698,N_29471);
or UO_242 (O_242,N_29712,N_29714);
and UO_243 (O_243,N_29671,N_29135);
or UO_244 (O_244,N_29036,N_29443);
and UO_245 (O_245,N_29619,N_29840);
nand UO_246 (O_246,N_29874,N_29777);
xnor UO_247 (O_247,N_29813,N_29626);
nand UO_248 (O_248,N_29591,N_29623);
or UO_249 (O_249,N_29561,N_29340);
nor UO_250 (O_250,N_29856,N_29128);
xor UO_251 (O_251,N_29878,N_29675);
xor UO_252 (O_252,N_29536,N_29360);
nor UO_253 (O_253,N_29103,N_29579);
nand UO_254 (O_254,N_29646,N_29915);
or UO_255 (O_255,N_29638,N_29498);
nor UO_256 (O_256,N_29905,N_29541);
and UO_257 (O_257,N_29986,N_29702);
nor UO_258 (O_258,N_29713,N_29896);
nor UO_259 (O_259,N_29572,N_29972);
or UO_260 (O_260,N_29270,N_29221);
or UO_261 (O_261,N_29630,N_29627);
or UO_262 (O_262,N_29472,N_29688);
and UO_263 (O_263,N_29665,N_29133);
nand UO_264 (O_264,N_29192,N_29672);
and UO_265 (O_265,N_29730,N_29885);
or UO_266 (O_266,N_29493,N_29926);
and UO_267 (O_267,N_29372,N_29919);
or UO_268 (O_268,N_29104,N_29129);
nand UO_269 (O_269,N_29060,N_29587);
and UO_270 (O_270,N_29717,N_29189);
xnor UO_271 (O_271,N_29924,N_29489);
xnor UO_272 (O_272,N_29592,N_29092);
or UO_273 (O_273,N_29486,N_29318);
xor UO_274 (O_274,N_29278,N_29352);
and UO_275 (O_275,N_29548,N_29814);
nor UO_276 (O_276,N_29449,N_29706);
nor UO_277 (O_277,N_29549,N_29081);
nor UO_278 (O_278,N_29528,N_29326);
or UO_279 (O_279,N_29429,N_29351);
and UO_280 (O_280,N_29439,N_29323);
xor UO_281 (O_281,N_29358,N_29302);
nand UO_282 (O_282,N_29761,N_29526);
and UO_283 (O_283,N_29300,N_29205);
nor UO_284 (O_284,N_29308,N_29644);
or UO_285 (O_285,N_29968,N_29294);
or UO_286 (O_286,N_29483,N_29950);
nor UO_287 (O_287,N_29349,N_29421);
nor UO_288 (O_288,N_29357,N_29927);
or UO_289 (O_289,N_29284,N_29140);
nor UO_290 (O_290,N_29947,N_29000);
xnor UO_291 (O_291,N_29378,N_29858);
or UO_292 (O_292,N_29875,N_29361);
nor UO_293 (O_293,N_29312,N_29292);
xor UO_294 (O_294,N_29500,N_29186);
nor UO_295 (O_295,N_29854,N_29102);
nand UO_296 (O_296,N_29460,N_29072);
nor UO_297 (O_297,N_29111,N_29190);
nand UO_298 (O_298,N_29652,N_29880);
and UO_299 (O_299,N_29338,N_29825);
or UO_300 (O_300,N_29037,N_29602);
nor UO_301 (O_301,N_29719,N_29231);
and UO_302 (O_302,N_29689,N_29262);
xor UO_303 (O_303,N_29734,N_29982);
and UO_304 (O_304,N_29769,N_29809);
nor UO_305 (O_305,N_29286,N_29784);
nand UO_306 (O_306,N_29922,N_29478);
nand UO_307 (O_307,N_29369,N_29808);
and UO_308 (O_308,N_29831,N_29269);
xnor UO_309 (O_309,N_29625,N_29501);
xor UO_310 (O_310,N_29272,N_29876);
nor UO_311 (O_311,N_29534,N_29183);
nand UO_312 (O_312,N_29157,N_29804);
nand UO_313 (O_313,N_29957,N_29799);
and UO_314 (O_314,N_29227,N_29387);
or UO_315 (O_315,N_29695,N_29962);
or UO_316 (O_316,N_29313,N_29913);
nor UO_317 (O_317,N_29797,N_29182);
nand UO_318 (O_318,N_29969,N_29889);
xor UO_319 (O_319,N_29266,N_29480);
nor UO_320 (O_320,N_29198,N_29944);
and UO_321 (O_321,N_29933,N_29010);
nor UO_322 (O_322,N_29575,N_29417);
nand UO_323 (O_323,N_29914,N_29829);
nor UO_324 (O_324,N_29447,N_29527);
or UO_325 (O_325,N_29546,N_29676);
or UO_326 (O_326,N_29930,N_29137);
nor UO_327 (O_327,N_29291,N_29428);
and UO_328 (O_328,N_29204,N_29423);
or UO_329 (O_329,N_29374,N_29206);
nand UO_330 (O_330,N_29011,N_29531);
nor UO_331 (O_331,N_29742,N_29867);
nor UO_332 (O_332,N_29100,N_29343);
nand UO_333 (O_333,N_29289,N_29263);
or UO_334 (O_334,N_29288,N_29568);
and UO_335 (O_335,N_29131,N_29147);
and UO_336 (O_336,N_29760,N_29790);
or UO_337 (O_337,N_29897,N_29260);
or UO_338 (O_338,N_29339,N_29295);
nor UO_339 (O_339,N_29552,N_29517);
nor UO_340 (O_340,N_29303,N_29795);
nor UO_341 (O_341,N_29293,N_29708);
or UO_342 (O_342,N_29918,N_29632);
and UO_343 (O_343,N_29175,N_29408);
or UO_344 (O_344,N_29557,N_29647);
or UO_345 (O_345,N_29796,N_29497);
nand UO_346 (O_346,N_29635,N_29337);
or UO_347 (O_347,N_29738,N_29234);
or UO_348 (O_348,N_29321,N_29994);
xor UO_349 (O_349,N_29145,N_29187);
and UO_350 (O_350,N_29409,N_29739);
and UO_351 (O_351,N_29492,N_29705);
xor UO_352 (O_352,N_29159,N_29846);
or UO_353 (O_353,N_29955,N_29362);
xnor UO_354 (O_354,N_29750,N_29332);
or UO_355 (O_355,N_29153,N_29934);
xor UO_356 (O_356,N_29330,N_29425);
and UO_357 (O_357,N_29901,N_29941);
nor UO_358 (O_358,N_29119,N_29946);
or UO_359 (O_359,N_29843,N_29588);
or UO_360 (O_360,N_29882,N_29494);
nor UO_361 (O_361,N_29544,N_29765);
nand UO_362 (O_362,N_29792,N_29740);
and UO_363 (O_363,N_29311,N_29322);
xnor UO_364 (O_364,N_29095,N_29048);
xnor UO_365 (O_365,N_29193,N_29992);
nor UO_366 (O_366,N_29167,N_29974);
and UO_367 (O_367,N_29028,N_29411);
xor UO_368 (O_368,N_29964,N_29271);
nand UO_369 (O_369,N_29624,N_29376);
and UO_370 (O_370,N_29315,N_29002);
or UO_371 (O_371,N_29410,N_29451);
nand UO_372 (O_372,N_29868,N_29700);
xnor UO_373 (O_373,N_29396,N_29027);
nand UO_374 (O_374,N_29356,N_29077);
or UO_375 (O_375,N_29052,N_29521);
xor UO_376 (O_376,N_29181,N_29432);
xor UO_377 (O_377,N_29683,N_29458);
xnor UO_378 (O_378,N_29731,N_29973);
nor UO_379 (O_379,N_29658,N_29902);
nand UO_380 (O_380,N_29383,N_29801);
nor UO_381 (O_381,N_29656,N_29487);
nor UO_382 (O_382,N_29241,N_29505);
or UO_383 (O_383,N_29188,N_29860);
nor UO_384 (O_384,N_29412,N_29975);
and UO_385 (O_385,N_29711,N_29988);
xor UO_386 (O_386,N_29006,N_29649);
xnor UO_387 (O_387,N_29298,N_29353);
or UO_388 (O_388,N_29980,N_29386);
and UO_389 (O_389,N_29218,N_29144);
nand UO_390 (O_390,N_29348,N_29570);
xor UO_391 (O_391,N_29007,N_29574);
xor UO_392 (O_392,N_29068,N_29462);
nand UO_393 (O_393,N_29275,N_29921);
nand UO_394 (O_394,N_29199,N_29222);
nor UO_395 (O_395,N_29191,N_29442);
nor UO_396 (O_396,N_29121,N_29124);
and UO_397 (O_397,N_29976,N_29399);
and UO_398 (O_398,N_29310,N_29954);
nor UO_399 (O_399,N_29959,N_29999);
or UO_400 (O_400,N_29607,N_29737);
or UO_401 (O_401,N_29014,N_29283);
nand UO_402 (O_402,N_29143,N_29743);
and UO_403 (O_403,N_29807,N_29791);
and UO_404 (O_404,N_29212,N_29851);
and UO_405 (O_405,N_29155,N_29047);
or UO_406 (O_406,N_29845,N_29727);
nand UO_407 (O_407,N_29253,N_29822);
and UO_408 (O_408,N_29113,N_29707);
nand UO_409 (O_409,N_29958,N_29775);
xnor UO_410 (O_410,N_29171,N_29589);
nor UO_411 (O_411,N_29788,N_29643);
and UO_412 (O_412,N_29306,N_29062);
and UO_413 (O_413,N_29674,N_29114);
nor UO_414 (O_414,N_29961,N_29022);
xor UO_415 (O_415,N_29903,N_29600);
nor UO_416 (O_416,N_29641,N_29400);
nor UO_417 (O_417,N_29800,N_29177);
and UO_418 (O_418,N_29948,N_29373);
nand UO_419 (O_419,N_29035,N_29375);
nor UO_420 (O_420,N_29051,N_29820);
xnor UO_421 (O_421,N_29655,N_29567);
nand UO_422 (O_422,N_29200,N_29041);
xor UO_423 (O_423,N_29653,N_29637);
xnor UO_424 (O_424,N_29767,N_29735);
nand UO_425 (O_425,N_29091,N_29457);
nor UO_426 (O_426,N_29196,N_29749);
xnor UO_427 (O_427,N_29810,N_29660);
nor UO_428 (O_428,N_29085,N_29728);
xnor UO_429 (O_429,N_29220,N_29667);
or UO_430 (O_430,N_29597,N_29754);
nor UO_431 (O_431,N_29782,N_29146);
nor UO_432 (O_432,N_29482,N_29236);
nand UO_433 (O_433,N_29139,N_29097);
nor UO_434 (O_434,N_29377,N_29907);
or UO_435 (O_435,N_29049,N_29299);
nand UO_436 (O_436,N_29584,N_29499);
or UO_437 (O_437,N_29433,N_29056);
or UO_438 (O_438,N_29481,N_29513);
and UO_439 (O_439,N_29603,N_29074);
and UO_440 (O_440,N_29437,N_29148);
xnor UO_441 (O_441,N_29381,N_29033);
and UO_442 (O_442,N_29088,N_29940);
nor UO_443 (O_443,N_29164,N_29606);
nand UO_444 (O_444,N_29058,N_29009);
nor UO_445 (O_445,N_29533,N_29614);
and UO_446 (O_446,N_29438,N_29774);
nor UO_447 (O_447,N_29141,N_29247);
or UO_448 (O_448,N_29368,N_29082);
xnor UO_449 (O_449,N_29938,N_29872);
or UO_450 (O_450,N_29826,N_29888);
nand UO_451 (O_451,N_29753,N_29013);
nand UO_452 (O_452,N_29830,N_29279);
and UO_453 (O_453,N_29450,N_29586);
nor UO_454 (O_454,N_29105,N_29251);
nand UO_455 (O_455,N_29640,N_29194);
nand UO_456 (O_456,N_29895,N_29636);
or UO_457 (O_457,N_29237,N_29297);
and UO_458 (O_458,N_29301,N_29834);
nand UO_459 (O_459,N_29287,N_29887);
xor UO_460 (O_460,N_29477,N_29488);
nand UO_461 (O_461,N_29122,N_29931);
nand UO_462 (O_462,N_29180,N_29821);
nor UO_463 (O_463,N_29169,N_29904);
nand UO_464 (O_464,N_29729,N_29254);
or UO_465 (O_465,N_29459,N_29285);
nor UO_466 (O_466,N_29722,N_29923);
nor UO_467 (O_467,N_29172,N_29773);
and UO_468 (O_468,N_29008,N_29550);
xnor UO_469 (O_469,N_29259,N_29985);
and UO_470 (O_470,N_29952,N_29639);
and UO_471 (O_471,N_29928,N_29094);
or UO_472 (O_472,N_29214,N_29609);
nand UO_473 (O_473,N_29666,N_29083);
xnor UO_474 (O_474,N_29327,N_29075);
nor UO_475 (O_475,N_29314,N_29987);
nor UO_476 (O_476,N_29989,N_29912);
or UO_477 (O_477,N_29406,N_29174);
or UO_478 (O_478,N_29057,N_29608);
xnor UO_479 (O_479,N_29066,N_29479);
xor UO_480 (O_480,N_29426,N_29359);
nand UO_481 (O_481,N_29853,N_29654);
nor UO_482 (O_482,N_29678,N_29648);
nand UO_483 (O_483,N_29553,N_29469);
and UO_484 (O_484,N_29967,N_29166);
xor UO_485 (O_485,N_29506,N_29165);
and UO_486 (O_486,N_29651,N_29758);
nand UO_487 (O_487,N_29884,N_29604);
nor UO_488 (O_488,N_29642,N_29511);
nor UO_489 (O_489,N_29069,N_29690);
nand UO_490 (O_490,N_29217,N_29663);
nand UO_491 (O_491,N_29610,N_29680);
nor UO_492 (O_492,N_29224,N_29290);
and UO_493 (O_493,N_29201,N_29844);
nor UO_494 (O_494,N_29692,N_29762);
nor UO_495 (O_495,N_29661,N_29569);
and UO_496 (O_496,N_29709,N_29045);
xor UO_497 (O_497,N_29850,N_29031);
nand UO_498 (O_498,N_29824,N_29965);
or UO_499 (O_499,N_29890,N_29346);
xor UO_500 (O_500,N_29136,N_29638);
nand UO_501 (O_501,N_29201,N_29860);
or UO_502 (O_502,N_29873,N_29300);
or UO_503 (O_503,N_29211,N_29451);
and UO_504 (O_504,N_29262,N_29664);
and UO_505 (O_505,N_29864,N_29135);
xor UO_506 (O_506,N_29381,N_29124);
and UO_507 (O_507,N_29398,N_29686);
and UO_508 (O_508,N_29426,N_29443);
nand UO_509 (O_509,N_29063,N_29825);
nor UO_510 (O_510,N_29913,N_29821);
or UO_511 (O_511,N_29120,N_29305);
or UO_512 (O_512,N_29819,N_29909);
and UO_513 (O_513,N_29737,N_29473);
nor UO_514 (O_514,N_29074,N_29987);
xnor UO_515 (O_515,N_29524,N_29979);
xor UO_516 (O_516,N_29700,N_29971);
xnor UO_517 (O_517,N_29280,N_29605);
and UO_518 (O_518,N_29438,N_29144);
xor UO_519 (O_519,N_29746,N_29073);
xnor UO_520 (O_520,N_29964,N_29494);
or UO_521 (O_521,N_29329,N_29249);
nor UO_522 (O_522,N_29509,N_29036);
nor UO_523 (O_523,N_29290,N_29617);
nand UO_524 (O_524,N_29882,N_29017);
nor UO_525 (O_525,N_29190,N_29966);
and UO_526 (O_526,N_29732,N_29138);
xor UO_527 (O_527,N_29944,N_29773);
nand UO_528 (O_528,N_29001,N_29264);
nor UO_529 (O_529,N_29958,N_29075);
or UO_530 (O_530,N_29975,N_29376);
nand UO_531 (O_531,N_29305,N_29571);
xnor UO_532 (O_532,N_29268,N_29067);
and UO_533 (O_533,N_29394,N_29154);
nand UO_534 (O_534,N_29118,N_29155);
nand UO_535 (O_535,N_29840,N_29424);
nor UO_536 (O_536,N_29062,N_29898);
and UO_537 (O_537,N_29386,N_29640);
nand UO_538 (O_538,N_29315,N_29483);
or UO_539 (O_539,N_29263,N_29902);
or UO_540 (O_540,N_29255,N_29774);
nand UO_541 (O_541,N_29251,N_29317);
nand UO_542 (O_542,N_29431,N_29690);
or UO_543 (O_543,N_29998,N_29023);
or UO_544 (O_544,N_29255,N_29029);
xnor UO_545 (O_545,N_29916,N_29365);
and UO_546 (O_546,N_29609,N_29971);
nor UO_547 (O_547,N_29601,N_29324);
nand UO_548 (O_548,N_29499,N_29777);
xnor UO_549 (O_549,N_29602,N_29133);
or UO_550 (O_550,N_29542,N_29710);
or UO_551 (O_551,N_29860,N_29341);
or UO_552 (O_552,N_29936,N_29314);
or UO_553 (O_553,N_29100,N_29556);
and UO_554 (O_554,N_29075,N_29023);
or UO_555 (O_555,N_29434,N_29220);
and UO_556 (O_556,N_29596,N_29451);
and UO_557 (O_557,N_29980,N_29202);
nand UO_558 (O_558,N_29340,N_29566);
or UO_559 (O_559,N_29037,N_29303);
nand UO_560 (O_560,N_29511,N_29551);
nand UO_561 (O_561,N_29938,N_29453);
xnor UO_562 (O_562,N_29254,N_29368);
and UO_563 (O_563,N_29211,N_29773);
nand UO_564 (O_564,N_29968,N_29018);
nand UO_565 (O_565,N_29255,N_29227);
and UO_566 (O_566,N_29880,N_29155);
nor UO_567 (O_567,N_29425,N_29587);
nand UO_568 (O_568,N_29937,N_29036);
xor UO_569 (O_569,N_29837,N_29500);
or UO_570 (O_570,N_29055,N_29443);
nand UO_571 (O_571,N_29034,N_29716);
or UO_572 (O_572,N_29496,N_29214);
nor UO_573 (O_573,N_29491,N_29137);
nor UO_574 (O_574,N_29922,N_29225);
and UO_575 (O_575,N_29189,N_29177);
nor UO_576 (O_576,N_29172,N_29523);
nand UO_577 (O_577,N_29889,N_29044);
and UO_578 (O_578,N_29939,N_29262);
nor UO_579 (O_579,N_29706,N_29377);
or UO_580 (O_580,N_29526,N_29610);
nand UO_581 (O_581,N_29571,N_29820);
xnor UO_582 (O_582,N_29678,N_29246);
xnor UO_583 (O_583,N_29904,N_29756);
and UO_584 (O_584,N_29466,N_29828);
or UO_585 (O_585,N_29287,N_29324);
or UO_586 (O_586,N_29797,N_29408);
nor UO_587 (O_587,N_29528,N_29199);
nand UO_588 (O_588,N_29479,N_29744);
or UO_589 (O_589,N_29213,N_29055);
and UO_590 (O_590,N_29403,N_29730);
nor UO_591 (O_591,N_29169,N_29763);
and UO_592 (O_592,N_29275,N_29964);
xor UO_593 (O_593,N_29315,N_29577);
or UO_594 (O_594,N_29580,N_29078);
or UO_595 (O_595,N_29148,N_29643);
or UO_596 (O_596,N_29010,N_29393);
and UO_597 (O_597,N_29066,N_29710);
nor UO_598 (O_598,N_29588,N_29344);
xnor UO_599 (O_599,N_29337,N_29045);
xor UO_600 (O_600,N_29075,N_29652);
and UO_601 (O_601,N_29672,N_29999);
xor UO_602 (O_602,N_29987,N_29208);
or UO_603 (O_603,N_29393,N_29821);
nand UO_604 (O_604,N_29848,N_29829);
nor UO_605 (O_605,N_29117,N_29895);
or UO_606 (O_606,N_29905,N_29902);
xor UO_607 (O_607,N_29514,N_29448);
nor UO_608 (O_608,N_29003,N_29727);
nor UO_609 (O_609,N_29977,N_29365);
nor UO_610 (O_610,N_29637,N_29279);
nor UO_611 (O_611,N_29935,N_29792);
xnor UO_612 (O_612,N_29828,N_29513);
nand UO_613 (O_613,N_29451,N_29419);
xnor UO_614 (O_614,N_29357,N_29693);
nand UO_615 (O_615,N_29909,N_29889);
or UO_616 (O_616,N_29371,N_29245);
nor UO_617 (O_617,N_29292,N_29422);
and UO_618 (O_618,N_29180,N_29603);
and UO_619 (O_619,N_29001,N_29385);
nor UO_620 (O_620,N_29898,N_29451);
nand UO_621 (O_621,N_29772,N_29232);
or UO_622 (O_622,N_29104,N_29878);
nor UO_623 (O_623,N_29886,N_29071);
nand UO_624 (O_624,N_29341,N_29840);
and UO_625 (O_625,N_29796,N_29916);
and UO_626 (O_626,N_29540,N_29202);
nand UO_627 (O_627,N_29948,N_29654);
nand UO_628 (O_628,N_29693,N_29606);
xor UO_629 (O_629,N_29697,N_29626);
or UO_630 (O_630,N_29495,N_29140);
nand UO_631 (O_631,N_29111,N_29442);
or UO_632 (O_632,N_29789,N_29321);
nand UO_633 (O_633,N_29869,N_29199);
nand UO_634 (O_634,N_29984,N_29666);
xnor UO_635 (O_635,N_29258,N_29928);
xor UO_636 (O_636,N_29080,N_29079);
xor UO_637 (O_637,N_29333,N_29666);
and UO_638 (O_638,N_29646,N_29976);
nor UO_639 (O_639,N_29191,N_29351);
or UO_640 (O_640,N_29076,N_29178);
nand UO_641 (O_641,N_29097,N_29886);
or UO_642 (O_642,N_29405,N_29831);
nor UO_643 (O_643,N_29275,N_29739);
or UO_644 (O_644,N_29964,N_29270);
xor UO_645 (O_645,N_29712,N_29855);
xnor UO_646 (O_646,N_29192,N_29962);
or UO_647 (O_647,N_29177,N_29446);
xnor UO_648 (O_648,N_29110,N_29624);
nand UO_649 (O_649,N_29764,N_29516);
nor UO_650 (O_650,N_29059,N_29936);
or UO_651 (O_651,N_29490,N_29552);
and UO_652 (O_652,N_29363,N_29798);
and UO_653 (O_653,N_29322,N_29154);
xnor UO_654 (O_654,N_29325,N_29781);
nand UO_655 (O_655,N_29854,N_29694);
or UO_656 (O_656,N_29593,N_29804);
and UO_657 (O_657,N_29297,N_29408);
nand UO_658 (O_658,N_29806,N_29296);
xnor UO_659 (O_659,N_29881,N_29956);
and UO_660 (O_660,N_29949,N_29264);
and UO_661 (O_661,N_29418,N_29339);
and UO_662 (O_662,N_29744,N_29031);
nand UO_663 (O_663,N_29778,N_29628);
xor UO_664 (O_664,N_29253,N_29422);
xnor UO_665 (O_665,N_29386,N_29579);
nand UO_666 (O_666,N_29952,N_29949);
xor UO_667 (O_667,N_29418,N_29224);
and UO_668 (O_668,N_29230,N_29607);
or UO_669 (O_669,N_29769,N_29669);
and UO_670 (O_670,N_29600,N_29669);
or UO_671 (O_671,N_29046,N_29230);
xnor UO_672 (O_672,N_29287,N_29271);
nand UO_673 (O_673,N_29742,N_29450);
nand UO_674 (O_674,N_29319,N_29147);
or UO_675 (O_675,N_29566,N_29941);
nand UO_676 (O_676,N_29101,N_29481);
nand UO_677 (O_677,N_29374,N_29929);
nor UO_678 (O_678,N_29245,N_29219);
or UO_679 (O_679,N_29328,N_29460);
and UO_680 (O_680,N_29959,N_29533);
or UO_681 (O_681,N_29210,N_29251);
nand UO_682 (O_682,N_29318,N_29707);
or UO_683 (O_683,N_29866,N_29020);
or UO_684 (O_684,N_29951,N_29397);
xnor UO_685 (O_685,N_29749,N_29963);
or UO_686 (O_686,N_29606,N_29375);
nand UO_687 (O_687,N_29993,N_29432);
and UO_688 (O_688,N_29058,N_29209);
nand UO_689 (O_689,N_29096,N_29709);
nand UO_690 (O_690,N_29506,N_29933);
xor UO_691 (O_691,N_29642,N_29174);
and UO_692 (O_692,N_29421,N_29265);
or UO_693 (O_693,N_29350,N_29988);
xor UO_694 (O_694,N_29039,N_29649);
or UO_695 (O_695,N_29281,N_29648);
xnor UO_696 (O_696,N_29750,N_29544);
nor UO_697 (O_697,N_29714,N_29827);
nor UO_698 (O_698,N_29600,N_29089);
nand UO_699 (O_699,N_29440,N_29596);
or UO_700 (O_700,N_29560,N_29999);
xnor UO_701 (O_701,N_29962,N_29073);
and UO_702 (O_702,N_29346,N_29908);
nand UO_703 (O_703,N_29577,N_29670);
or UO_704 (O_704,N_29142,N_29480);
and UO_705 (O_705,N_29298,N_29695);
and UO_706 (O_706,N_29894,N_29104);
xnor UO_707 (O_707,N_29831,N_29126);
and UO_708 (O_708,N_29891,N_29596);
xnor UO_709 (O_709,N_29952,N_29726);
xnor UO_710 (O_710,N_29305,N_29612);
or UO_711 (O_711,N_29519,N_29288);
xor UO_712 (O_712,N_29102,N_29158);
nor UO_713 (O_713,N_29020,N_29268);
or UO_714 (O_714,N_29049,N_29186);
nand UO_715 (O_715,N_29663,N_29012);
and UO_716 (O_716,N_29617,N_29933);
xor UO_717 (O_717,N_29443,N_29456);
xor UO_718 (O_718,N_29198,N_29063);
or UO_719 (O_719,N_29862,N_29082);
nand UO_720 (O_720,N_29114,N_29218);
nor UO_721 (O_721,N_29022,N_29226);
nand UO_722 (O_722,N_29232,N_29150);
nor UO_723 (O_723,N_29067,N_29179);
nor UO_724 (O_724,N_29840,N_29976);
xnor UO_725 (O_725,N_29111,N_29575);
nor UO_726 (O_726,N_29889,N_29761);
nand UO_727 (O_727,N_29371,N_29384);
and UO_728 (O_728,N_29303,N_29409);
or UO_729 (O_729,N_29228,N_29930);
nand UO_730 (O_730,N_29082,N_29871);
or UO_731 (O_731,N_29345,N_29943);
or UO_732 (O_732,N_29761,N_29291);
xnor UO_733 (O_733,N_29383,N_29384);
or UO_734 (O_734,N_29416,N_29104);
nand UO_735 (O_735,N_29934,N_29833);
and UO_736 (O_736,N_29556,N_29011);
nor UO_737 (O_737,N_29527,N_29229);
and UO_738 (O_738,N_29960,N_29215);
or UO_739 (O_739,N_29337,N_29564);
and UO_740 (O_740,N_29851,N_29913);
or UO_741 (O_741,N_29873,N_29961);
nor UO_742 (O_742,N_29841,N_29644);
nand UO_743 (O_743,N_29288,N_29795);
or UO_744 (O_744,N_29190,N_29677);
or UO_745 (O_745,N_29381,N_29604);
xnor UO_746 (O_746,N_29421,N_29895);
xor UO_747 (O_747,N_29216,N_29678);
or UO_748 (O_748,N_29183,N_29667);
nor UO_749 (O_749,N_29530,N_29377);
or UO_750 (O_750,N_29967,N_29428);
nor UO_751 (O_751,N_29509,N_29847);
xnor UO_752 (O_752,N_29573,N_29072);
nand UO_753 (O_753,N_29729,N_29773);
xnor UO_754 (O_754,N_29124,N_29499);
nor UO_755 (O_755,N_29290,N_29983);
nand UO_756 (O_756,N_29053,N_29311);
xnor UO_757 (O_757,N_29437,N_29477);
and UO_758 (O_758,N_29628,N_29202);
and UO_759 (O_759,N_29550,N_29888);
xnor UO_760 (O_760,N_29189,N_29666);
xnor UO_761 (O_761,N_29718,N_29522);
nor UO_762 (O_762,N_29431,N_29845);
xnor UO_763 (O_763,N_29609,N_29752);
or UO_764 (O_764,N_29781,N_29969);
or UO_765 (O_765,N_29649,N_29949);
and UO_766 (O_766,N_29918,N_29148);
nor UO_767 (O_767,N_29638,N_29039);
or UO_768 (O_768,N_29408,N_29228);
xor UO_769 (O_769,N_29720,N_29230);
and UO_770 (O_770,N_29164,N_29811);
xor UO_771 (O_771,N_29082,N_29059);
nand UO_772 (O_772,N_29365,N_29826);
nor UO_773 (O_773,N_29346,N_29940);
and UO_774 (O_774,N_29193,N_29351);
and UO_775 (O_775,N_29494,N_29654);
and UO_776 (O_776,N_29012,N_29708);
or UO_777 (O_777,N_29141,N_29098);
and UO_778 (O_778,N_29004,N_29003);
and UO_779 (O_779,N_29796,N_29180);
or UO_780 (O_780,N_29462,N_29655);
nand UO_781 (O_781,N_29962,N_29466);
xnor UO_782 (O_782,N_29424,N_29385);
nand UO_783 (O_783,N_29241,N_29285);
and UO_784 (O_784,N_29131,N_29670);
nor UO_785 (O_785,N_29699,N_29474);
nor UO_786 (O_786,N_29224,N_29499);
or UO_787 (O_787,N_29730,N_29489);
and UO_788 (O_788,N_29475,N_29941);
and UO_789 (O_789,N_29287,N_29614);
or UO_790 (O_790,N_29087,N_29591);
xor UO_791 (O_791,N_29033,N_29058);
and UO_792 (O_792,N_29653,N_29359);
or UO_793 (O_793,N_29644,N_29527);
and UO_794 (O_794,N_29654,N_29521);
nor UO_795 (O_795,N_29394,N_29178);
nand UO_796 (O_796,N_29469,N_29830);
nor UO_797 (O_797,N_29327,N_29022);
nor UO_798 (O_798,N_29932,N_29992);
xnor UO_799 (O_799,N_29223,N_29799);
nand UO_800 (O_800,N_29038,N_29480);
nand UO_801 (O_801,N_29050,N_29909);
xor UO_802 (O_802,N_29721,N_29792);
nor UO_803 (O_803,N_29891,N_29399);
or UO_804 (O_804,N_29374,N_29426);
nand UO_805 (O_805,N_29180,N_29607);
xor UO_806 (O_806,N_29492,N_29365);
and UO_807 (O_807,N_29664,N_29649);
or UO_808 (O_808,N_29454,N_29349);
nor UO_809 (O_809,N_29898,N_29433);
or UO_810 (O_810,N_29746,N_29082);
xor UO_811 (O_811,N_29828,N_29719);
or UO_812 (O_812,N_29988,N_29060);
xor UO_813 (O_813,N_29570,N_29415);
nor UO_814 (O_814,N_29474,N_29317);
xnor UO_815 (O_815,N_29335,N_29373);
xor UO_816 (O_816,N_29523,N_29056);
or UO_817 (O_817,N_29640,N_29783);
nand UO_818 (O_818,N_29052,N_29874);
xor UO_819 (O_819,N_29356,N_29716);
nand UO_820 (O_820,N_29169,N_29813);
xor UO_821 (O_821,N_29095,N_29624);
and UO_822 (O_822,N_29028,N_29583);
or UO_823 (O_823,N_29355,N_29622);
nor UO_824 (O_824,N_29342,N_29857);
xnor UO_825 (O_825,N_29236,N_29649);
nand UO_826 (O_826,N_29272,N_29422);
xnor UO_827 (O_827,N_29181,N_29875);
xor UO_828 (O_828,N_29337,N_29086);
xor UO_829 (O_829,N_29591,N_29657);
xnor UO_830 (O_830,N_29234,N_29879);
and UO_831 (O_831,N_29061,N_29028);
or UO_832 (O_832,N_29133,N_29595);
xnor UO_833 (O_833,N_29693,N_29017);
or UO_834 (O_834,N_29032,N_29119);
nand UO_835 (O_835,N_29487,N_29426);
and UO_836 (O_836,N_29220,N_29567);
and UO_837 (O_837,N_29968,N_29677);
xor UO_838 (O_838,N_29018,N_29183);
nand UO_839 (O_839,N_29956,N_29220);
and UO_840 (O_840,N_29795,N_29614);
xnor UO_841 (O_841,N_29652,N_29400);
xor UO_842 (O_842,N_29381,N_29290);
nor UO_843 (O_843,N_29962,N_29743);
nand UO_844 (O_844,N_29619,N_29490);
xnor UO_845 (O_845,N_29081,N_29909);
and UO_846 (O_846,N_29491,N_29684);
xnor UO_847 (O_847,N_29904,N_29306);
xnor UO_848 (O_848,N_29943,N_29972);
and UO_849 (O_849,N_29977,N_29924);
and UO_850 (O_850,N_29792,N_29917);
nor UO_851 (O_851,N_29893,N_29573);
and UO_852 (O_852,N_29657,N_29061);
nand UO_853 (O_853,N_29558,N_29330);
or UO_854 (O_854,N_29219,N_29259);
nor UO_855 (O_855,N_29328,N_29392);
xnor UO_856 (O_856,N_29618,N_29411);
nand UO_857 (O_857,N_29540,N_29704);
nand UO_858 (O_858,N_29704,N_29334);
and UO_859 (O_859,N_29369,N_29840);
xnor UO_860 (O_860,N_29829,N_29844);
nor UO_861 (O_861,N_29049,N_29300);
or UO_862 (O_862,N_29399,N_29017);
xor UO_863 (O_863,N_29291,N_29277);
and UO_864 (O_864,N_29822,N_29859);
or UO_865 (O_865,N_29266,N_29422);
nor UO_866 (O_866,N_29751,N_29098);
or UO_867 (O_867,N_29476,N_29499);
nand UO_868 (O_868,N_29545,N_29104);
nor UO_869 (O_869,N_29056,N_29442);
xor UO_870 (O_870,N_29382,N_29698);
nand UO_871 (O_871,N_29134,N_29392);
and UO_872 (O_872,N_29377,N_29232);
nor UO_873 (O_873,N_29203,N_29942);
xnor UO_874 (O_874,N_29585,N_29022);
xnor UO_875 (O_875,N_29112,N_29305);
and UO_876 (O_876,N_29851,N_29003);
nand UO_877 (O_877,N_29745,N_29303);
xor UO_878 (O_878,N_29288,N_29019);
and UO_879 (O_879,N_29938,N_29144);
nand UO_880 (O_880,N_29352,N_29808);
xnor UO_881 (O_881,N_29311,N_29226);
xor UO_882 (O_882,N_29327,N_29542);
xnor UO_883 (O_883,N_29948,N_29466);
xnor UO_884 (O_884,N_29716,N_29571);
or UO_885 (O_885,N_29854,N_29399);
xor UO_886 (O_886,N_29006,N_29941);
xnor UO_887 (O_887,N_29731,N_29063);
nand UO_888 (O_888,N_29748,N_29518);
nand UO_889 (O_889,N_29405,N_29903);
xor UO_890 (O_890,N_29848,N_29560);
xnor UO_891 (O_891,N_29338,N_29090);
nand UO_892 (O_892,N_29568,N_29949);
or UO_893 (O_893,N_29531,N_29108);
or UO_894 (O_894,N_29839,N_29692);
nand UO_895 (O_895,N_29831,N_29445);
nor UO_896 (O_896,N_29931,N_29664);
nor UO_897 (O_897,N_29358,N_29051);
or UO_898 (O_898,N_29534,N_29351);
nand UO_899 (O_899,N_29787,N_29954);
or UO_900 (O_900,N_29362,N_29480);
nand UO_901 (O_901,N_29736,N_29177);
and UO_902 (O_902,N_29395,N_29487);
nor UO_903 (O_903,N_29712,N_29523);
nand UO_904 (O_904,N_29828,N_29211);
xnor UO_905 (O_905,N_29778,N_29177);
or UO_906 (O_906,N_29372,N_29043);
xnor UO_907 (O_907,N_29937,N_29162);
and UO_908 (O_908,N_29816,N_29290);
xnor UO_909 (O_909,N_29989,N_29901);
and UO_910 (O_910,N_29591,N_29808);
nand UO_911 (O_911,N_29472,N_29992);
nor UO_912 (O_912,N_29130,N_29699);
nand UO_913 (O_913,N_29854,N_29068);
nor UO_914 (O_914,N_29706,N_29511);
nor UO_915 (O_915,N_29204,N_29767);
nor UO_916 (O_916,N_29467,N_29947);
and UO_917 (O_917,N_29595,N_29499);
and UO_918 (O_918,N_29436,N_29543);
or UO_919 (O_919,N_29735,N_29900);
nand UO_920 (O_920,N_29164,N_29856);
xor UO_921 (O_921,N_29272,N_29523);
xor UO_922 (O_922,N_29495,N_29197);
xnor UO_923 (O_923,N_29373,N_29880);
nor UO_924 (O_924,N_29110,N_29807);
nand UO_925 (O_925,N_29505,N_29194);
nand UO_926 (O_926,N_29765,N_29898);
nor UO_927 (O_927,N_29354,N_29373);
and UO_928 (O_928,N_29853,N_29270);
xnor UO_929 (O_929,N_29311,N_29385);
or UO_930 (O_930,N_29145,N_29611);
nor UO_931 (O_931,N_29545,N_29758);
or UO_932 (O_932,N_29164,N_29117);
nand UO_933 (O_933,N_29051,N_29107);
xnor UO_934 (O_934,N_29138,N_29832);
nand UO_935 (O_935,N_29800,N_29932);
nor UO_936 (O_936,N_29023,N_29429);
or UO_937 (O_937,N_29641,N_29294);
or UO_938 (O_938,N_29944,N_29723);
and UO_939 (O_939,N_29706,N_29988);
and UO_940 (O_940,N_29256,N_29878);
nor UO_941 (O_941,N_29070,N_29548);
nor UO_942 (O_942,N_29680,N_29803);
or UO_943 (O_943,N_29610,N_29681);
nand UO_944 (O_944,N_29634,N_29061);
and UO_945 (O_945,N_29464,N_29635);
or UO_946 (O_946,N_29363,N_29498);
and UO_947 (O_947,N_29081,N_29945);
xnor UO_948 (O_948,N_29611,N_29430);
nand UO_949 (O_949,N_29640,N_29229);
nor UO_950 (O_950,N_29526,N_29300);
and UO_951 (O_951,N_29135,N_29189);
nand UO_952 (O_952,N_29974,N_29285);
or UO_953 (O_953,N_29032,N_29105);
and UO_954 (O_954,N_29619,N_29110);
xnor UO_955 (O_955,N_29921,N_29313);
xor UO_956 (O_956,N_29957,N_29137);
xnor UO_957 (O_957,N_29881,N_29555);
nor UO_958 (O_958,N_29292,N_29040);
or UO_959 (O_959,N_29289,N_29658);
nand UO_960 (O_960,N_29192,N_29105);
and UO_961 (O_961,N_29125,N_29676);
and UO_962 (O_962,N_29365,N_29911);
or UO_963 (O_963,N_29208,N_29661);
nor UO_964 (O_964,N_29933,N_29784);
nor UO_965 (O_965,N_29751,N_29302);
nor UO_966 (O_966,N_29153,N_29104);
xor UO_967 (O_967,N_29764,N_29910);
nor UO_968 (O_968,N_29196,N_29014);
nand UO_969 (O_969,N_29266,N_29091);
nand UO_970 (O_970,N_29050,N_29149);
nand UO_971 (O_971,N_29805,N_29877);
xnor UO_972 (O_972,N_29581,N_29172);
or UO_973 (O_973,N_29726,N_29596);
and UO_974 (O_974,N_29580,N_29850);
xor UO_975 (O_975,N_29096,N_29164);
xor UO_976 (O_976,N_29413,N_29937);
xnor UO_977 (O_977,N_29451,N_29650);
or UO_978 (O_978,N_29483,N_29041);
and UO_979 (O_979,N_29076,N_29068);
and UO_980 (O_980,N_29008,N_29656);
nor UO_981 (O_981,N_29394,N_29331);
xor UO_982 (O_982,N_29077,N_29930);
or UO_983 (O_983,N_29009,N_29073);
nor UO_984 (O_984,N_29116,N_29352);
or UO_985 (O_985,N_29245,N_29134);
xnor UO_986 (O_986,N_29163,N_29459);
and UO_987 (O_987,N_29989,N_29577);
and UO_988 (O_988,N_29763,N_29788);
or UO_989 (O_989,N_29859,N_29900);
nor UO_990 (O_990,N_29674,N_29235);
or UO_991 (O_991,N_29435,N_29366);
and UO_992 (O_992,N_29442,N_29160);
nor UO_993 (O_993,N_29550,N_29189);
or UO_994 (O_994,N_29424,N_29719);
xor UO_995 (O_995,N_29060,N_29649);
or UO_996 (O_996,N_29131,N_29886);
xnor UO_997 (O_997,N_29298,N_29986);
nand UO_998 (O_998,N_29198,N_29481);
nor UO_999 (O_999,N_29471,N_29867);
nor UO_1000 (O_1000,N_29437,N_29874);
nand UO_1001 (O_1001,N_29732,N_29963);
nor UO_1002 (O_1002,N_29644,N_29008);
and UO_1003 (O_1003,N_29159,N_29062);
nor UO_1004 (O_1004,N_29137,N_29560);
nor UO_1005 (O_1005,N_29773,N_29859);
and UO_1006 (O_1006,N_29318,N_29265);
xnor UO_1007 (O_1007,N_29989,N_29267);
nand UO_1008 (O_1008,N_29018,N_29862);
xor UO_1009 (O_1009,N_29915,N_29598);
nand UO_1010 (O_1010,N_29545,N_29645);
nor UO_1011 (O_1011,N_29395,N_29097);
xor UO_1012 (O_1012,N_29471,N_29660);
xnor UO_1013 (O_1013,N_29282,N_29709);
or UO_1014 (O_1014,N_29416,N_29887);
xor UO_1015 (O_1015,N_29162,N_29031);
xnor UO_1016 (O_1016,N_29225,N_29947);
xor UO_1017 (O_1017,N_29512,N_29300);
nor UO_1018 (O_1018,N_29167,N_29404);
nand UO_1019 (O_1019,N_29217,N_29211);
or UO_1020 (O_1020,N_29571,N_29540);
or UO_1021 (O_1021,N_29246,N_29116);
or UO_1022 (O_1022,N_29216,N_29426);
nor UO_1023 (O_1023,N_29769,N_29710);
or UO_1024 (O_1024,N_29267,N_29213);
and UO_1025 (O_1025,N_29706,N_29339);
xnor UO_1026 (O_1026,N_29386,N_29060);
and UO_1027 (O_1027,N_29161,N_29939);
or UO_1028 (O_1028,N_29572,N_29425);
nor UO_1029 (O_1029,N_29002,N_29504);
or UO_1030 (O_1030,N_29475,N_29464);
or UO_1031 (O_1031,N_29165,N_29594);
and UO_1032 (O_1032,N_29834,N_29063);
xor UO_1033 (O_1033,N_29098,N_29311);
nor UO_1034 (O_1034,N_29777,N_29045);
nand UO_1035 (O_1035,N_29218,N_29240);
nand UO_1036 (O_1036,N_29076,N_29001);
and UO_1037 (O_1037,N_29829,N_29647);
nor UO_1038 (O_1038,N_29812,N_29641);
nand UO_1039 (O_1039,N_29300,N_29958);
nor UO_1040 (O_1040,N_29352,N_29957);
or UO_1041 (O_1041,N_29020,N_29269);
xor UO_1042 (O_1042,N_29309,N_29621);
xor UO_1043 (O_1043,N_29404,N_29265);
nand UO_1044 (O_1044,N_29417,N_29990);
or UO_1045 (O_1045,N_29612,N_29247);
nor UO_1046 (O_1046,N_29600,N_29202);
xnor UO_1047 (O_1047,N_29202,N_29584);
xor UO_1048 (O_1048,N_29625,N_29687);
xnor UO_1049 (O_1049,N_29341,N_29154);
or UO_1050 (O_1050,N_29778,N_29004);
and UO_1051 (O_1051,N_29191,N_29521);
and UO_1052 (O_1052,N_29407,N_29141);
nor UO_1053 (O_1053,N_29133,N_29473);
and UO_1054 (O_1054,N_29747,N_29286);
nand UO_1055 (O_1055,N_29976,N_29336);
nand UO_1056 (O_1056,N_29718,N_29425);
and UO_1057 (O_1057,N_29622,N_29190);
nor UO_1058 (O_1058,N_29101,N_29041);
and UO_1059 (O_1059,N_29492,N_29067);
nand UO_1060 (O_1060,N_29595,N_29476);
xnor UO_1061 (O_1061,N_29927,N_29868);
and UO_1062 (O_1062,N_29950,N_29621);
nand UO_1063 (O_1063,N_29707,N_29360);
or UO_1064 (O_1064,N_29769,N_29840);
or UO_1065 (O_1065,N_29086,N_29383);
nand UO_1066 (O_1066,N_29824,N_29237);
or UO_1067 (O_1067,N_29357,N_29621);
xor UO_1068 (O_1068,N_29433,N_29131);
xnor UO_1069 (O_1069,N_29787,N_29556);
xor UO_1070 (O_1070,N_29753,N_29999);
xnor UO_1071 (O_1071,N_29589,N_29832);
nand UO_1072 (O_1072,N_29655,N_29085);
or UO_1073 (O_1073,N_29487,N_29873);
and UO_1074 (O_1074,N_29662,N_29312);
xor UO_1075 (O_1075,N_29543,N_29098);
and UO_1076 (O_1076,N_29863,N_29662);
or UO_1077 (O_1077,N_29559,N_29079);
nand UO_1078 (O_1078,N_29568,N_29560);
nor UO_1079 (O_1079,N_29864,N_29368);
or UO_1080 (O_1080,N_29186,N_29428);
nor UO_1081 (O_1081,N_29424,N_29653);
nor UO_1082 (O_1082,N_29254,N_29975);
or UO_1083 (O_1083,N_29178,N_29995);
nand UO_1084 (O_1084,N_29543,N_29106);
nand UO_1085 (O_1085,N_29079,N_29677);
xnor UO_1086 (O_1086,N_29958,N_29061);
or UO_1087 (O_1087,N_29250,N_29487);
nand UO_1088 (O_1088,N_29788,N_29681);
and UO_1089 (O_1089,N_29808,N_29238);
nand UO_1090 (O_1090,N_29242,N_29324);
nand UO_1091 (O_1091,N_29002,N_29013);
and UO_1092 (O_1092,N_29371,N_29242);
nand UO_1093 (O_1093,N_29907,N_29318);
nand UO_1094 (O_1094,N_29720,N_29772);
and UO_1095 (O_1095,N_29942,N_29558);
nor UO_1096 (O_1096,N_29545,N_29885);
or UO_1097 (O_1097,N_29115,N_29931);
xor UO_1098 (O_1098,N_29637,N_29589);
and UO_1099 (O_1099,N_29345,N_29666);
nor UO_1100 (O_1100,N_29591,N_29171);
and UO_1101 (O_1101,N_29238,N_29886);
nor UO_1102 (O_1102,N_29174,N_29868);
nor UO_1103 (O_1103,N_29008,N_29555);
xor UO_1104 (O_1104,N_29474,N_29021);
nand UO_1105 (O_1105,N_29056,N_29258);
or UO_1106 (O_1106,N_29474,N_29142);
or UO_1107 (O_1107,N_29687,N_29375);
nor UO_1108 (O_1108,N_29942,N_29807);
nand UO_1109 (O_1109,N_29909,N_29840);
nand UO_1110 (O_1110,N_29364,N_29688);
or UO_1111 (O_1111,N_29984,N_29182);
nand UO_1112 (O_1112,N_29209,N_29793);
nand UO_1113 (O_1113,N_29940,N_29644);
xor UO_1114 (O_1114,N_29589,N_29599);
and UO_1115 (O_1115,N_29023,N_29807);
nor UO_1116 (O_1116,N_29278,N_29291);
or UO_1117 (O_1117,N_29317,N_29534);
xnor UO_1118 (O_1118,N_29627,N_29123);
nand UO_1119 (O_1119,N_29323,N_29404);
or UO_1120 (O_1120,N_29564,N_29660);
nor UO_1121 (O_1121,N_29327,N_29132);
and UO_1122 (O_1122,N_29765,N_29378);
nor UO_1123 (O_1123,N_29991,N_29076);
or UO_1124 (O_1124,N_29632,N_29992);
and UO_1125 (O_1125,N_29847,N_29935);
or UO_1126 (O_1126,N_29813,N_29504);
nor UO_1127 (O_1127,N_29893,N_29417);
and UO_1128 (O_1128,N_29877,N_29564);
and UO_1129 (O_1129,N_29413,N_29503);
xor UO_1130 (O_1130,N_29268,N_29075);
nor UO_1131 (O_1131,N_29948,N_29771);
or UO_1132 (O_1132,N_29248,N_29572);
xor UO_1133 (O_1133,N_29868,N_29743);
nor UO_1134 (O_1134,N_29118,N_29200);
and UO_1135 (O_1135,N_29119,N_29563);
xnor UO_1136 (O_1136,N_29147,N_29449);
or UO_1137 (O_1137,N_29747,N_29555);
or UO_1138 (O_1138,N_29853,N_29362);
nor UO_1139 (O_1139,N_29117,N_29141);
or UO_1140 (O_1140,N_29018,N_29554);
or UO_1141 (O_1141,N_29042,N_29854);
and UO_1142 (O_1142,N_29812,N_29937);
nand UO_1143 (O_1143,N_29993,N_29489);
or UO_1144 (O_1144,N_29405,N_29215);
or UO_1145 (O_1145,N_29380,N_29825);
and UO_1146 (O_1146,N_29766,N_29356);
nor UO_1147 (O_1147,N_29885,N_29229);
and UO_1148 (O_1148,N_29015,N_29834);
and UO_1149 (O_1149,N_29796,N_29111);
and UO_1150 (O_1150,N_29859,N_29059);
or UO_1151 (O_1151,N_29902,N_29058);
and UO_1152 (O_1152,N_29995,N_29689);
and UO_1153 (O_1153,N_29917,N_29651);
xor UO_1154 (O_1154,N_29512,N_29266);
nand UO_1155 (O_1155,N_29401,N_29364);
nor UO_1156 (O_1156,N_29812,N_29315);
nor UO_1157 (O_1157,N_29323,N_29186);
nor UO_1158 (O_1158,N_29425,N_29692);
nor UO_1159 (O_1159,N_29821,N_29548);
nor UO_1160 (O_1160,N_29179,N_29086);
and UO_1161 (O_1161,N_29601,N_29993);
xnor UO_1162 (O_1162,N_29425,N_29766);
nor UO_1163 (O_1163,N_29017,N_29612);
nand UO_1164 (O_1164,N_29751,N_29280);
xor UO_1165 (O_1165,N_29154,N_29085);
or UO_1166 (O_1166,N_29873,N_29462);
and UO_1167 (O_1167,N_29589,N_29104);
and UO_1168 (O_1168,N_29503,N_29810);
or UO_1169 (O_1169,N_29564,N_29918);
nor UO_1170 (O_1170,N_29129,N_29972);
and UO_1171 (O_1171,N_29362,N_29497);
or UO_1172 (O_1172,N_29497,N_29807);
or UO_1173 (O_1173,N_29271,N_29799);
xor UO_1174 (O_1174,N_29722,N_29456);
or UO_1175 (O_1175,N_29040,N_29084);
and UO_1176 (O_1176,N_29542,N_29550);
or UO_1177 (O_1177,N_29312,N_29580);
and UO_1178 (O_1178,N_29311,N_29603);
and UO_1179 (O_1179,N_29067,N_29933);
nand UO_1180 (O_1180,N_29183,N_29254);
nor UO_1181 (O_1181,N_29425,N_29828);
xnor UO_1182 (O_1182,N_29617,N_29391);
or UO_1183 (O_1183,N_29767,N_29322);
and UO_1184 (O_1184,N_29513,N_29362);
nor UO_1185 (O_1185,N_29024,N_29317);
nand UO_1186 (O_1186,N_29057,N_29828);
or UO_1187 (O_1187,N_29280,N_29258);
nor UO_1188 (O_1188,N_29924,N_29684);
nand UO_1189 (O_1189,N_29879,N_29878);
nand UO_1190 (O_1190,N_29001,N_29137);
xnor UO_1191 (O_1191,N_29161,N_29844);
xor UO_1192 (O_1192,N_29316,N_29013);
and UO_1193 (O_1193,N_29496,N_29506);
nand UO_1194 (O_1194,N_29289,N_29330);
and UO_1195 (O_1195,N_29505,N_29711);
or UO_1196 (O_1196,N_29691,N_29272);
nand UO_1197 (O_1197,N_29380,N_29804);
nor UO_1198 (O_1198,N_29971,N_29483);
nor UO_1199 (O_1199,N_29645,N_29553);
nand UO_1200 (O_1200,N_29319,N_29202);
nor UO_1201 (O_1201,N_29265,N_29362);
or UO_1202 (O_1202,N_29265,N_29934);
xor UO_1203 (O_1203,N_29971,N_29953);
and UO_1204 (O_1204,N_29731,N_29950);
nor UO_1205 (O_1205,N_29332,N_29787);
nand UO_1206 (O_1206,N_29664,N_29542);
nand UO_1207 (O_1207,N_29185,N_29111);
and UO_1208 (O_1208,N_29234,N_29732);
and UO_1209 (O_1209,N_29754,N_29728);
nand UO_1210 (O_1210,N_29650,N_29739);
and UO_1211 (O_1211,N_29441,N_29198);
xnor UO_1212 (O_1212,N_29801,N_29523);
xor UO_1213 (O_1213,N_29245,N_29076);
nand UO_1214 (O_1214,N_29130,N_29414);
nor UO_1215 (O_1215,N_29385,N_29439);
and UO_1216 (O_1216,N_29476,N_29349);
nor UO_1217 (O_1217,N_29988,N_29694);
nand UO_1218 (O_1218,N_29055,N_29079);
nor UO_1219 (O_1219,N_29773,N_29863);
and UO_1220 (O_1220,N_29090,N_29660);
nand UO_1221 (O_1221,N_29503,N_29551);
and UO_1222 (O_1222,N_29350,N_29958);
or UO_1223 (O_1223,N_29938,N_29967);
and UO_1224 (O_1224,N_29562,N_29558);
or UO_1225 (O_1225,N_29710,N_29109);
and UO_1226 (O_1226,N_29315,N_29619);
xnor UO_1227 (O_1227,N_29218,N_29495);
xnor UO_1228 (O_1228,N_29288,N_29563);
nor UO_1229 (O_1229,N_29410,N_29687);
and UO_1230 (O_1230,N_29750,N_29173);
nor UO_1231 (O_1231,N_29063,N_29090);
nor UO_1232 (O_1232,N_29079,N_29652);
and UO_1233 (O_1233,N_29499,N_29590);
and UO_1234 (O_1234,N_29499,N_29330);
nor UO_1235 (O_1235,N_29430,N_29015);
nand UO_1236 (O_1236,N_29627,N_29438);
or UO_1237 (O_1237,N_29743,N_29525);
nor UO_1238 (O_1238,N_29879,N_29172);
or UO_1239 (O_1239,N_29544,N_29590);
nor UO_1240 (O_1240,N_29118,N_29870);
nor UO_1241 (O_1241,N_29243,N_29348);
nand UO_1242 (O_1242,N_29390,N_29190);
nor UO_1243 (O_1243,N_29215,N_29600);
and UO_1244 (O_1244,N_29174,N_29045);
and UO_1245 (O_1245,N_29324,N_29866);
xnor UO_1246 (O_1246,N_29740,N_29969);
xor UO_1247 (O_1247,N_29175,N_29203);
or UO_1248 (O_1248,N_29136,N_29118);
nand UO_1249 (O_1249,N_29319,N_29841);
or UO_1250 (O_1250,N_29282,N_29596);
nor UO_1251 (O_1251,N_29641,N_29388);
nor UO_1252 (O_1252,N_29267,N_29649);
and UO_1253 (O_1253,N_29948,N_29608);
nor UO_1254 (O_1254,N_29655,N_29501);
nor UO_1255 (O_1255,N_29409,N_29529);
nor UO_1256 (O_1256,N_29707,N_29655);
nor UO_1257 (O_1257,N_29074,N_29896);
xor UO_1258 (O_1258,N_29760,N_29224);
and UO_1259 (O_1259,N_29329,N_29315);
nand UO_1260 (O_1260,N_29934,N_29580);
nand UO_1261 (O_1261,N_29189,N_29469);
or UO_1262 (O_1262,N_29572,N_29947);
nor UO_1263 (O_1263,N_29214,N_29128);
xor UO_1264 (O_1264,N_29254,N_29072);
nand UO_1265 (O_1265,N_29152,N_29550);
or UO_1266 (O_1266,N_29337,N_29123);
xor UO_1267 (O_1267,N_29472,N_29589);
nand UO_1268 (O_1268,N_29931,N_29719);
nor UO_1269 (O_1269,N_29345,N_29450);
nand UO_1270 (O_1270,N_29817,N_29279);
xnor UO_1271 (O_1271,N_29725,N_29357);
xnor UO_1272 (O_1272,N_29011,N_29768);
or UO_1273 (O_1273,N_29550,N_29799);
and UO_1274 (O_1274,N_29349,N_29831);
or UO_1275 (O_1275,N_29993,N_29359);
nor UO_1276 (O_1276,N_29263,N_29543);
and UO_1277 (O_1277,N_29996,N_29266);
and UO_1278 (O_1278,N_29035,N_29944);
nand UO_1279 (O_1279,N_29224,N_29165);
xnor UO_1280 (O_1280,N_29968,N_29769);
nor UO_1281 (O_1281,N_29584,N_29233);
xor UO_1282 (O_1282,N_29177,N_29330);
nand UO_1283 (O_1283,N_29314,N_29257);
and UO_1284 (O_1284,N_29383,N_29990);
nor UO_1285 (O_1285,N_29028,N_29598);
and UO_1286 (O_1286,N_29085,N_29318);
nor UO_1287 (O_1287,N_29368,N_29747);
or UO_1288 (O_1288,N_29430,N_29929);
or UO_1289 (O_1289,N_29308,N_29359);
xor UO_1290 (O_1290,N_29932,N_29660);
or UO_1291 (O_1291,N_29014,N_29704);
or UO_1292 (O_1292,N_29353,N_29194);
xor UO_1293 (O_1293,N_29074,N_29266);
or UO_1294 (O_1294,N_29208,N_29068);
or UO_1295 (O_1295,N_29920,N_29752);
or UO_1296 (O_1296,N_29930,N_29784);
nor UO_1297 (O_1297,N_29599,N_29070);
nor UO_1298 (O_1298,N_29797,N_29107);
nand UO_1299 (O_1299,N_29810,N_29894);
or UO_1300 (O_1300,N_29342,N_29478);
or UO_1301 (O_1301,N_29098,N_29257);
and UO_1302 (O_1302,N_29112,N_29758);
or UO_1303 (O_1303,N_29605,N_29016);
or UO_1304 (O_1304,N_29363,N_29062);
nand UO_1305 (O_1305,N_29502,N_29931);
nor UO_1306 (O_1306,N_29325,N_29172);
nor UO_1307 (O_1307,N_29841,N_29263);
nor UO_1308 (O_1308,N_29763,N_29475);
nand UO_1309 (O_1309,N_29055,N_29982);
nand UO_1310 (O_1310,N_29205,N_29419);
nand UO_1311 (O_1311,N_29270,N_29464);
and UO_1312 (O_1312,N_29365,N_29545);
nand UO_1313 (O_1313,N_29922,N_29692);
nor UO_1314 (O_1314,N_29143,N_29069);
nor UO_1315 (O_1315,N_29245,N_29608);
xnor UO_1316 (O_1316,N_29151,N_29336);
or UO_1317 (O_1317,N_29968,N_29304);
or UO_1318 (O_1318,N_29656,N_29499);
xor UO_1319 (O_1319,N_29990,N_29427);
nand UO_1320 (O_1320,N_29780,N_29451);
nand UO_1321 (O_1321,N_29342,N_29699);
or UO_1322 (O_1322,N_29144,N_29826);
xor UO_1323 (O_1323,N_29475,N_29161);
xor UO_1324 (O_1324,N_29690,N_29443);
and UO_1325 (O_1325,N_29646,N_29448);
nor UO_1326 (O_1326,N_29978,N_29901);
and UO_1327 (O_1327,N_29299,N_29849);
and UO_1328 (O_1328,N_29929,N_29583);
nand UO_1329 (O_1329,N_29355,N_29245);
and UO_1330 (O_1330,N_29328,N_29593);
nand UO_1331 (O_1331,N_29111,N_29029);
nor UO_1332 (O_1332,N_29681,N_29684);
nor UO_1333 (O_1333,N_29384,N_29162);
xor UO_1334 (O_1334,N_29009,N_29435);
xnor UO_1335 (O_1335,N_29928,N_29469);
nand UO_1336 (O_1336,N_29931,N_29016);
or UO_1337 (O_1337,N_29478,N_29329);
or UO_1338 (O_1338,N_29461,N_29031);
nor UO_1339 (O_1339,N_29392,N_29035);
nor UO_1340 (O_1340,N_29627,N_29195);
and UO_1341 (O_1341,N_29002,N_29693);
xnor UO_1342 (O_1342,N_29834,N_29113);
nor UO_1343 (O_1343,N_29786,N_29959);
and UO_1344 (O_1344,N_29816,N_29271);
or UO_1345 (O_1345,N_29064,N_29859);
xnor UO_1346 (O_1346,N_29329,N_29990);
xor UO_1347 (O_1347,N_29555,N_29137);
or UO_1348 (O_1348,N_29326,N_29651);
or UO_1349 (O_1349,N_29811,N_29424);
or UO_1350 (O_1350,N_29715,N_29637);
or UO_1351 (O_1351,N_29042,N_29976);
or UO_1352 (O_1352,N_29423,N_29274);
and UO_1353 (O_1353,N_29314,N_29578);
and UO_1354 (O_1354,N_29892,N_29879);
xnor UO_1355 (O_1355,N_29459,N_29334);
nand UO_1356 (O_1356,N_29639,N_29911);
nand UO_1357 (O_1357,N_29039,N_29396);
or UO_1358 (O_1358,N_29957,N_29058);
nor UO_1359 (O_1359,N_29890,N_29442);
xor UO_1360 (O_1360,N_29761,N_29805);
nand UO_1361 (O_1361,N_29928,N_29193);
or UO_1362 (O_1362,N_29879,N_29836);
nand UO_1363 (O_1363,N_29757,N_29679);
and UO_1364 (O_1364,N_29075,N_29762);
nor UO_1365 (O_1365,N_29451,N_29538);
nor UO_1366 (O_1366,N_29608,N_29044);
nand UO_1367 (O_1367,N_29927,N_29305);
or UO_1368 (O_1368,N_29003,N_29869);
xnor UO_1369 (O_1369,N_29845,N_29926);
nor UO_1370 (O_1370,N_29963,N_29600);
or UO_1371 (O_1371,N_29728,N_29168);
and UO_1372 (O_1372,N_29111,N_29632);
nand UO_1373 (O_1373,N_29123,N_29137);
or UO_1374 (O_1374,N_29794,N_29930);
or UO_1375 (O_1375,N_29180,N_29354);
nand UO_1376 (O_1376,N_29580,N_29519);
nor UO_1377 (O_1377,N_29174,N_29568);
or UO_1378 (O_1378,N_29476,N_29759);
nand UO_1379 (O_1379,N_29442,N_29812);
or UO_1380 (O_1380,N_29305,N_29918);
and UO_1381 (O_1381,N_29144,N_29632);
xnor UO_1382 (O_1382,N_29758,N_29761);
nor UO_1383 (O_1383,N_29295,N_29757);
nand UO_1384 (O_1384,N_29935,N_29037);
nor UO_1385 (O_1385,N_29745,N_29804);
and UO_1386 (O_1386,N_29713,N_29602);
and UO_1387 (O_1387,N_29900,N_29932);
nand UO_1388 (O_1388,N_29206,N_29692);
nand UO_1389 (O_1389,N_29521,N_29704);
or UO_1390 (O_1390,N_29865,N_29330);
xnor UO_1391 (O_1391,N_29744,N_29885);
and UO_1392 (O_1392,N_29733,N_29151);
and UO_1393 (O_1393,N_29068,N_29883);
and UO_1394 (O_1394,N_29874,N_29793);
and UO_1395 (O_1395,N_29544,N_29736);
xor UO_1396 (O_1396,N_29319,N_29156);
nor UO_1397 (O_1397,N_29025,N_29865);
nand UO_1398 (O_1398,N_29349,N_29815);
and UO_1399 (O_1399,N_29160,N_29505);
and UO_1400 (O_1400,N_29020,N_29525);
nand UO_1401 (O_1401,N_29956,N_29057);
and UO_1402 (O_1402,N_29149,N_29378);
and UO_1403 (O_1403,N_29703,N_29505);
nor UO_1404 (O_1404,N_29842,N_29928);
and UO_1405 (O_1405,N_29591,N_29436);
nand UO_1406 (O_1406,N_29994,N_29292);
and UO_1407 (O_1407,N_29350,N_29307);
and UO_1408 (O_1408,N_29887,N_29064);
xnor UO_1409 (O_1409,N_29284,N_29086);
or UO_1410 (O_1410,N_29760,N_29802);
nor UO_1411 (O_1411,N_29667,N_29414);
or UO_1412 (O_1412,N_29192,N_29563);
nor UO_1413 (O_1413,N_29912,N_29499);
xnor UO_1414 (O_1414,N_29274,N_29292);
nor UO_1415 (O_1415,N_29860,N_29034);
nand UO_1416 (O_1416,N_29062,N_29098);
xnor UO_1417 (O_1417,N_29235,N_29668);
nand UO_1418 (O_1418,N_29168,N_29147);
nor UO_1419 (O_1419,N_29294,N_29203);
and UO_1420 (O_1420,N_29684,N_29598);
xnor UO_1421 (O_1421,N_29849,N_29857);
or UO_1422 (O_1422,N_29641,N_29859);
nand UO_1423 (O_1423,N_29648,N_29651);
and UO_1424 (O_1424,N_29188,N_29096);
or UO_1425 (O_1425,N_29681,N_29452);
and UO_1426 (O_1426,N_29229,N_29215);
and UO_1427 (O_1427,N_29339,N_29671);
nor UO_1428 (O_1428,N_29298,N_29028);
xor UO_1429 (O_1429,N_29670,N_29098);
nor UO_1430 (O_1430,N_29774,N_29419);
xnor UO_1431 (O_1431,N_29362,N_29211);
nor UO_1432 (O_1432,N_29315,N_29460);
and UO_1433 (O_1433,N_29825,N_29233);
nor UO_1434 (O_1434,N_29823,N_29149);
nor UO_1435 (O_1435,N_29516,N_29573);
or UO_1436 (O_1436,N_29727,N_29210);
and UO_1437 (O_1437,N_29473,N_29603);
and UO_1438 (O_1438,N_29009,N_29099);
nand UO_1439 (O_1439,N_29652,N_29536);
nand UO_1440 (O_1440,N_29433,N_29219);
and UO_1441 (O_1441,N_29539,N_29417);
nor UO_1442 (O_1442,N_29619,N_29407);
nand UO_1443 (O_1443,N_29506,N_29371);
nand UO_1444 (O_1444,N_29773,N_29650);
nor UO_1445 (O_1445,N_29570,N_29267);
or UO_1446 (O_1446,N_29485,N_29014);
xnor UO_1447 (O_1447,N_29326,N_29248);
or UO_1448 (O_1448,N_29052,N_29090);
and UO_1449 (O_1449,N_29540,N_29839);
and UO_1450 (O_1450,N_29001,N_29214);
nand UO_1451 (O_1451,N_29130,N_29899);
nand UO_1452 (O_1452,N_29421,N_29866);
and UO_1453 (O_1453,N_29850,N_29488);
xnor UO_1454 (O_1454,N_29977,N_29193);
xor UO_1455 (O_1455,N_29171,N_29871);
xor UO_1456 (O_1456,N_29186,N_29287);
and UO_1457 (O_1457,N_29868,N_29526);
nor UO_1458 (O_1458,N_29136,N_29455);
and UO_1459 (O_1459,N_29487,N_29968);
nand UO_1460 (O_1460,N_29077,N_29483);
xnor UO_1461 (O_1461,N_29364,N_29781);
nor UO_1462 (O_1462,N_29819,N_29269);
nor UO_1463 (O_1463,N_29952,N_29360);
nor UO_1464 (O_1464,N_29882,N_29569);
and UO_1465 (O_1465,N_29710,N_29411);
nor UO_1466 (O_1466,N_29922,N_29845);
nand UO_1467 (O_1467,N_29494,N_29474);
or UO_1468 (O_1468,N_29321,N_29440);
nor UO_1469 (O_1469,N_29742,N_29756);
nand UO_1470 (O_1470,N_29711,N_29488);
or UO_1471 (O_1471,N_29995,N_29547);
nand UO_1472 (O_1472,N_29040,N_29427);
nand UO_1473 (O_1473,N_29366,N_29090);
nor UO_1474 (O_1474,N_29389,N_29033);
nor UO_1475 (O_1475,N_29375,N_29384);
xor UO_1476 (O_1476,N_29357,N_29666);
xnor UO_1477 (O_1477,N_29356,N_29253);
xor UO_1478 (O_1478,N_29936,N_29870);
or UO_1479 (O_1479,N_29175,N_29573);
and UO_1480 (O_1480,N_29280,N_29351);
nor UO_1481 (O_1481,N_29614,N_29633);
nor UO_1482 (O_1482,N_29028,N_29986);
or UO_1483 (O_1483,N_29703,N_29414);
and UO_1484 (O_1484,N_29196,N_29300);
and UO_1485 (O_1485,N_29943,N_29371);
or UO_1486 (O_1486,N_29063,N_29491);
and UO_1487 (O_1487,N_29049,N_29852);
or UO_1488 (O_1488,N_29412,N_29639);
xor UO_1489 (O_1489,N_29115,N_29023);
nand UO_1490 (O_1490,N_29566,N_29890);
nor UO_1491 (O_1491,N_29376,N_29999);
or UO_1492 (O_1492,N_29599,N_29308);
nand UO_1493 (O_1493,N_29906,N_29897);
nor UO_1494 (O_1494,N_29876,N_29610);
nand UO_1495 (O_1495,N_29019,N_29960);
xnor UO_1496 (O_1496,N_29300,N_29949);
or UO_1497 (O_1497,N_29759,N_29593);
or UO_1498 (O_1498,N_29939,N_29968);
and UO_1499 (O_1499,N_29356,N_29149);
nand UO_1500 (O_1500,N_29964,N_29916);
or UO_1501 (O_1501,N_29082,N_29225);
and UO_1502 (O_1502,N_29668,N_29406);
xor UO_1503 (O_1503,N_29590,N_29936);
nor UO_1504 (O_1504,N_29346,N_29018);
and UO_1505 (O_1505,N_29577,N_29460);
and UO_1506 (O_1506,N_29426,N_29752);
xor UO_1507 (O_1507,N_29784,N_29576);
nand UO_1508 (O_1508,N_29668,N_29404);
nand UO_1509 (O_1509,N_29392,N_29916);
xnor UO_1510 (O_1510,N_29992,N_29612);
nor UO_1511 (O_1511,N_29859,N_29495);
nand UO_1512 (O_1512,N_29885,N_29724);
or UO_1513 (O_1513,N_29111,N_29481);
and UO_1514 (O_1514,N_29095,N_29714);
or UO_1515 (O_1515,N_29306,N_29978);
or UO_1516 (O_1516,N_29576,N_29544);
nor UO_1517 (O_1517,N_29496,N_29409);
or UO_1518 (O_1518,N_29268,N_29879);
nor UO_1519 (O_1519,N_29558,N_29104);
or UO_1520 (O_1520,N_29671,N_29749);
nand UO_1521 (O_1521,N_29785,N_29036);
xor UO_1522 (O_1522,N_29292,N_29423);
nand UO_1523 (O_1523,N_29080,N_29904);
or UO_1524 (O_1524,N_29216,N_29932);
nor UO_1525 (O_1525,N_29703,N_29720);
xnor UO_1526 (O_1526,N_29615,N_29488);
or UO_1527 (O_1527,N_29511,N_29220);
xnor UO_1528 (O_1528,N_29976,N_29229);
nor UO_1529 (O_1529,N_29563,N_29043);
nor UO_1530 (O_1530,N_29153,N_29135);
nand UO_1531 (O_1531,N_29185,N_29166);
xor UO_1532 (O_1532,N_29050,N_29929);
or UO_1533 (O_1533,N_29916,N_29821);
and UO_1534 (O_1534,N_29128,N_29668);
nand UO_1535 (O_1535,N_29630,N_29802);
xor UO_1536 (O_1536,N_29602,N_29334);
nor UO_1537 (O_1537,N_29660,N_29773);
or UO_1538 (O_1538,N_29306,N_29471);
nor UO_1539 (O_1539,N_29271,N_29183);
nor UO_1540 (O_1540,N_29501,N_29020);
or UO_1541 (O_1541,N_29355,N_29685);
nand UO_1542 (O_1542,N_29796,N_29228);
or UO_1543 (O_1543,N_29675,N_29379);
xnor UO_1544 (O_1544,N_29828,N_29733);
xor UO_1545 (O_1545,N_29244,N_29502);
nor UO_1546 (O_1546,N_29943,N_29807);
nand UO_1547 (O_1547,N_29039,N_29498);
nand UO_1548 (O_1548,N_29748,N_29811);
xor UO_1549 (O_1549,N_29658,N_29730);
nand UO_1550 (O_1550,N_29027,N_29196);
or UO_1551 (O_1551,N_29270,N_29904);
and UO_1552 (O_1552,N_29035,N_29434);
or UO_1553 (O_1553,N_29699,N_29336);
and UO_1554 (O_1554,N_29147,N_29658);
or UO_1555 (O_1555,N_29555,N_29948);
xor UO_1556 (O_1556,N_29175,N_29337);
xor UO_1557 (O_1557,N_29868,N_29596);
or UO_1558 (O_1558,N_29603,N_29038);
or UO_1559 (O_1559,N_29860,N_29032);
and UO_1560 (O_1560,N_29080,N_29529);
xnor UO_1561 (O_1561,N_29836,N_29903);
xnor UO_1562 (O_1562,N_29522,N_29569);
xor UO_1563 (O_1563,N_29024,N_29270);
xnor UO_1564 (O_1564,N_29317,N_29307);
nand UO_1565 (O_1565,N_29374,N_29762);
nor UO_1566 (O_1566,N_29379,N_29346);
nand UO_1567 (O_1567,N_29808,N_29700);
nand UO_1568 (O_1568,N_29360,N_29772);
and UO_1569 (O_1569,N_29646,N_29723);
nand UO_1570 (O_1570,N_29337,N_29863);
and UO_1571 (O_1571,N_29004,N_29626);
nor UO_1572 (O_1572,N_29012,N_29884);
nand UO_1573 (O_1573,N_29531,N_29809);
xnor UO_1574 (O_1574,N_29053,N_29781);
nand UO_1575 (O_1575,N_29439,N_29488);
xor UO_1576 (O_1576,N_29928,N_29517);
xnor UO_1577 (O_1577,N_29302,N_29161);
nor UO_1578 (O_1578,N_29042,N_29106);
nand UO_1579 (O_1579,N_29808,N_29145);
nand UO_1580 (O_1580,N_29812,N_29974);
or UO_1581 (O_1581,N_29062,N_29691);
and UO_1582 (O_1582,N_29121,N_29962);
nor UO_1583 (O_1583,N_29808,N_29524);
and UO_1584 (O_1584,N_29975,N_29315);
nand UO_1585 (O_1585,N_29729,N_29798);
xor UO_1586 (O_1586,N_29452,N_29350);
nor UO_1587 (O_1587,N_29013,N_29480);
nor UO_1588 (O_1588,N_29325,N_29840);
and UO_1589 (O_1589,N_29874,N_29051);
and UO_1590 (O_1590,N_29120,N_29384);
and UO_1591 (O_1591,N_29118,N_29812);
nor UO_1592 (O_1592,N_29476,N_29204);
and UO_1593 (O_1593,N_29665,N_29111);
nand UO_1594 (O_1594,N_29552,N_29258);
xnor UO_1595 (O_1595,N_29865,N_29489);
xnor UO_1596 (O_1596,N_29294,N_29025);
nor UO_1597 (O_1597,N_29612,N_29450);
xnor UO_1598 (O_1598,N_29502,N_29320);
xor UO_1599 (O_1599,N_29192,N_29118);
nand UO_1600 (O_1600,N_29481,N_29393);
nor UO_1601 (O_1601,N_29058,N_29564);
nand UO_1602 (O_1602,N_29769,N_29770);
and UO_1603 (O_1603,N_29302,N_29964);
or UO_1604 (O_1604,N_29193,N_29602);
nand UO_1605 (O_1605,N_29945,N_29035);
or UO_1606 (O_1606,N_29410,N_29071);
or UO_1607 (O_1607,N_29858,N_29273);
nand UO_1608 (O_1608,N_29245,N_29399);
xnor UO_1609 (O_1609,N_29141,N_29985);
and UO_1610 (O_1610,N_29698,N_29536);
and UO_1611 (O_1611,N_29675,N_29141);
nand UO_1612 (O_1612,N_29682,N_29921);
or UO_1613 (O_1613,N_29148,N_29018);
and UO_1614 (O_1614,N_29647,N_29406);
nand UO_1615 (O_1615,N_29859,N_29719);
and UO_1616 (O_1616,N_29982,N_29434);
xor UO_1617 (O_1617,N_29479,N_29915);
and UO_1618 (O_1618,N_29895,N_29329);
and UO_1619 (O_1619,N_29484,N_29281);
nand UO_1620 (O_1620,N_29167,N_29889);
or UO_1621 (O_1621,N_29488,N_29535);
nor UO_1622 (O_1622,N_29256,N_29599);
nor UO_1623 (O_1623,N_29628,N_29822);
nand UO_1624 (O_1624,N_29832,N_29592);
and UO_1625 (O_1625,N_29526,N_29499);
nor UO_1626 (O_1626,N_29944,N_29554);
and UO_1627 (O_1627,N_29545,N_29707);
xnor UO_1628 (O_1628,N_29620,N_29328);
nor UO_1629 (O_1629,N_29943,N_29623);
or UO_1630 (O_1630,N_29262,N_29420);
nor UO_1631 (O_1631,N_29555,N_29744);
and UO_1632 (O_1632,N_29901,N_29618);
xnor UO_1633 (O_1633,N_29250,N_29639);
nand UO_1634 (O_1634,N_29381,N_29455);
nand UO_1635 (O_1635,N_29522,N_29714);
xor UO_1636 (O_1636,N_29915,N_29422);
nor UO_1637 (O_1637,N_29442,N_29583);
or UO_1638 (O_1638,N_29462,N_29620);
or UO_1639 (O_1639,N_29297,N_29284);
xor UO_1640 (O_1640,N_29795,N_29494);
and UO_1641 (O_1641,N_29140,N_29055);
nand UO_1642 (O_1642,N_29183,N_29215);
xor UO_1643 (O_1643,N_29658,N_29739);
nand UO_1644 (O_1644,N_29523,N_29574);
nor UO_1645 (O_1645,N_29585,N_29695);
xor UO_1646 (O_1646,N_29872,N_29949);
and UO_1647 (O_1647,N_29947,N_29549);
nand UO_1648 (O_1648,N_29574,N_29444);
xnor UO_1649 (O_1649,N_29781,N_29243);
nand UO_1650 (O_1650,N_29507,N_29634);
xor UO_1651 (O_1651,N_29982,N_29468);
xor UO_1652 (O_1652,N_29130,N_29486);
xnor UO_1653 (O_1653,N_29162,N_29892);
nor UO_1654 (O_1654,N_29531,N_29619);
xnor UO_1655 (O_1655,N_29184,N_29509);
nor UO_1656 (O_1656,N_29290,N_29739);
nor UO_1657 (O_1657,N_29175,N_29600);
and UO_1658 (O_1658,N_29769,N_29315);
or UO_1659 (O_1659,N_29163,N_29094);
or UO_1660 (O_1660,N_29252,N_29408);
nor UO_1661 (O_1661,N_29111,N_29752);
or UO_1662 (O_1662,N_29160,N_29043);
and UO_1663 (O_1663,N_29159,N_29270);
and UO_1664 (O_1664,N_29997,N_29995);
and UO_1665 (O_1665,N_29159,N_29860);
and UO_1666 (O_1666,N_29809,N_29582);
or UO_1667 (O_1667,N_29801,N_29219);
nand UO_1668 (O_1668,N_29049,N_29283);
nand UO_1669 (O_1669,N_29912,N_29664);
and UO_1670 (O_1670,N_29524,N_29526);
or UO_1671 (O_1671,N_29972,N_29122);
or UO_1672 (O_1672,N_29168,N_29944);
or UO_1673 (O_1673,N_29749,N_29701);
nand UO_1674 (O_1674,N_29904,N_29096);
nor UO_1675 (O_1675,N_29322,N_29319);
nor UO_1676 (O_1676,N_29358,N_29475);
or UO_1677 (O_1677,N_29638,N_29231);
nand UO_1678 (O_1678,N_29558,N_29729);
or UO_1679 (O_1679,N_29545,N_29701);
or UO_1680 (O_1680,N_29582,N_29606);
nor UO_1681 (O_1681,N_29304,N_29542);
xnor UO_1682 (O_1682,N_29436,N_29681);
nand UO_1683 (O_1683,N_29294,N_29166);
xor UO_1684 (O_1684,N_29521,N_29984);
or UO_1685 (O_1685,N_29727,N_29371);
nand UO_1686 (O_1686,N_29354,N_29527);
or UO_1687 (O_1687,N_29709,N_29365);
nand UO_1688 (O_1688,N_29109,N_29676);
xnor UO_1689 (O_1689,N_29210,N_29562);
and UO_1690 (O_1690,N_29484,N_29891);
and UO_1691 (O_1691,N_29186,N_29373);
nor UO_1692 (O_1692,N_29805,N_29019);
nor UO_1693 (O_1693,N_29872,N_29843);
or UO_1694 (O_1694,N_29387,N_29659);
or UO_1695 (O_1695,N_29713,N_29748);
nor UO_1696 (O_1696,N_29301,N_29388);
xor UO_1697 (O_1697,N_29727,N_29645);
nand UO_1698 (O_1698,N_29295,N_29178);
xnor UO_1699 (O_1699,N_29954,N_29353);
or UO_1700 (O_1700,N_29116,N_29159);
nor UO_1701 (O_1701,N_29848,N_29612);
xor UO_1702 (O_1702,N_29215,N_29755);
nand UO_1703 (O_1703,N_29399,N_29429);
nand UO_1704 (O_1704,N_29227,N_29996);
xnor UO_1705 (O_1705,N_29364,N_29717);
nand UO_1706 (O_1706,N_29214,N_29403);
or UO_1707 (O_1707,N_29034,N_29395);
xor UO_1708 (O_1708,N_29978,N_29802);
and UO_1709 (O_1709,N_29165,N_29709);
xor UO_1710 (O_1710,N_29969,N_29348);
xor UO_1711 (O_1711,N_29274,N_29702);
and UO_1712 (O_1712,N_29606,N_29104);
nor UO_1713 (O_1713,N_29200,N_29138);
and UO_1714 (O_1714,N_29929,N_29227);
nand UO_1715 (O_1715,N_29514,N_29122);
and UO_1716 (O_1716,N_29224,N_29331);
nand UO_1717 (O_1717,N_29056,N_29250);
xor UO_1718 (O_1718,N_29784,N_29593);
or UO_1719 (O_1719,N_29536,N_29341);
and UO_1720 (O_1720,N_29487,N_29880);
nor UO_1721 (O_1721,N_29512,N_29856);
nor UO_1722 (O_1722,N_29423,N_29630);
nand UO_1723 (O_1723,N_29655,N_29482);
or UO_1724 (O_1724,N_29928,N_29484);
nor UO_1725 (O_1725,N_29458,N_29083);
nand UO_1726 (O_1726,N_29744,N_29862);
xor UO_1727 (O_1727,N_29917,N_29726);
nand UO_1728 (O_1728,N_29762,N_29016);
nor UO_1729 (O_1729,N_29895,N_29139);
xor UO_1730 (O_1730,N_29301,N_29205);
xnor UO_1731 (O_1731,N_29842,N_29578);
or UO_1732 (O_1732,N_29519,N_29222);
xnor UO_1733 (O_1733,N_29537,N_29436);
xor UO_1734 (O_1734,N_29498,N_29106);
xnor UO_1735 (O_1735,N_29005,N_29513);
nand UO_1736 (O_1736,N_29743,N_29657);
nor UO_1737 (O_1737,N_29106,N_29888);
nand UO_1738 (O_1738,N_29598,N_29685);
nand UO_1739 (O_1739,N_29858,N_29177);
nor UO_1740 (O_1740,N_29292,N_29428);
xor UO_1741 (O_1741,N_29255,N_29980);
nand UO_1742 (O_1742,N_29326,N_29580);
or UO_1743 (O_1743,N_29824,N_29938);
and UO_1744 (O_1744,N_29970,N_29121);
and UO_1745 (O_1745,N_29084,N_29374);
or UO_1746 (O_1746,N_29503,N_29316);
nand UO_1747 (O_1747,N_29950,N_29673);
or UO_1748 (O_1748,N_29071,N_29778);
xnor UO_1749 (O_1749,N_29069,N_29248);
nand UO_1750 (O_1750,N_29198,N_29404);
nor UO_1751 (O_1751,N_29934,N_29898);
nor UO_1752 (O_1752,N_29117,N_29196);
xnor UO_1753 (O_1753,N_29435,N_29525);
xnor UO_1754 (O_1754,N_29694,N_29773);
or UO_1755 (O_1755,N_29673,N_29002);
or UO_1756 (O_1756,N_29190,N_29375);
xor UO_1757 (O_1757,N_29334,N_29448);
and UO_1758 (O_1758,N_29473,N_29003);
or UO_1759 (O_1759,N_29264,N_29191);
xnor UO_1760 (O_1760,N_29628,N_29857);
or UO_1761 (O_1761,N_29214,N_29863);
nand UO_1762 (O_1762,N_29974,N_29105);
and UO_1763 (O_1763,N_29955,N_29352);
nor UO_1764 (O_1764,N_29516,N_29993);
nand UO_1765 (O_1765,N_29607,N_29397);
and UO_1766 (O_1766,N_29281,N_29369);
nor UO_1767 (O_1767,N_29976,N_29032);
xor UO_1768 (O_1768,N_29462,N_29867);
and UO_1769 (O_1769,N_29315,N_29361);
nand UO_1770 (O_1770,N_29219,N_29085);
xnor UO_1771 (O_1771,N_29039,N_29852);
nor UO_1772 (O_1772,N_29641,N_29403);
xnor UO_1773 (O_1773,N_29087,N_29520);
or UO_1774 (O_1774,N_29882,N_29811);
nand UO_1775 (O_1775,N_29642,N_29406);
and UO_1776 (O_1776,N_29416,N_29262);
nand UO_1777 (O_1777,N_29016,N_29736);
or UO_1778 (O_1778,N_29715,N_29313);
xor UO_1779 (O_1779,N_29179,N_29858);
xnor UO_1780 (O_1780,N_29633,N_29904);
xnor UO_1781 (O_1781,N_29293,N_29291);
nor UO_1782 (O_1782,N_29412,N_29218);
and UO_1783 (O_1783,N_29918,N_29504);
nor UO_1784 (O_1784,N_29520,N_29655);
xor UO_1785 (O_1785,N_29197,N_29242);
nand UO_1786 (O_1786,N_29086,N_29849);
and UO_1787 (O_1787,N_29424,N_29980);
xnor UO_1788 (O_1788,N_29800,N_29353);
or UO_1789 (O_1789,N_29521,N_29597);
nand UO_1790 (O_1790,N_29112,N_29768);
or UO_1791 (O_1791,N_29932,N_29149);
nand UO_1792 (O_1792,N_29101,N_29025);
nand UO_1793 (O_1793,N_29241,N_29363);
nand UO_1794 (O_1794,N_29422,N_29187);
and UO_1795 (O_1795,N_29161,N_29148);
or UO_1796 (O_1796,N_29716,N_29609);
and UO_1797 (O_1797,N_29597,N_29685);
nor UO_1798 (O_1798,N_29926,N_29854);
nor UO_1799 (O_1799,N_29560,N_29789);
xnor UO_1800 (O_1800,N_29706,N_29848);
nor UO_1801 (O_1801,N_29983,N_29479);
nand UO_1802 (O_1802,N_29204,N_29164);
or UO_1803 (O_1803,N_29054,N_29658);
and UO_1804 (O_1804,N_29765,N_29049);
xnor UO_1805 (O_1805,N_29105,N_29219);
or UO_1806 (O_1806,N_29465,N_29906);
nor UO_1807 (O_1807,N_29874,N_29524);
nand UO_1808 (O_1808,N_29495,N_29855);
or UO_1809 (O_1809,N_29872,N_29991);
xor UO_1810 (O_1810,N_29093,N_29993);
xnor UO_1811 (O_1811,N_29479,N_29370);
nor UO_1812 (O_1812,N_29157,N_29371);
xnor UO_1813 (O_1813,N_29189,N_29261);
xor UO_1814 (O_1814,N_29548,N_29615);
and UO_1815 (O_1815,N_29023,N_29031);
nand UO_1816 (O_1816,N_29539,N_29086);
xnor UO_1817 (O_1817,N_29318,N_29302);
nand UO_1818 (O_1818,N_29289,N_29587);
nor UO_1819 (O_1819,N_29295,N_29095);
xnor UO_1820 (O_1820,N_29736,N_29142);
xor UO_1821 (O_1821,N_29666,N_29655);
and UO_1822 (O_1822,N_29509,N_29988);
and UO_1823 (O_1823,N_29643,N_29219);
xnor UO_1824 (O_1824,N_29958,N_29514);
or UO_1825 (O_1825,N_29416,N_29237);
xnor UO_1826 (O_1826,N_29012,N_29795);
or UO_1827 (O_1827,N_29239,N_29717);
nand UO_1828 (O_1828,N_29217,N_29650);
nand UO_1829 (O_1829,N_29216,N_29219);
xnor UO_1830 (O_1830,N_29972,N_29350);
or UO_1831 (O_1831,N_29266,N_29437);
nor UO_1832 (O_1832,N_29447,N_29462);
or UO_1833 (O_1833,N_29140,N_29801);
or UO_1834 (O_1834,N_29155,N_29827);
or UO_1835 (O_1835,N_29578,N_29834);
nor UO_1836 (O_1836,N_29528,N_29081);
or UO_1837 (O_1837,N_29296,N_29583);
and UO_1838 (O_1838,N_29181,N_29690);
or UO_1839 (O_1839,N_29971,N_29808);
and UO_1840 (O_1840,N_29566,N_29406);
nor UO_1841 (O_1841,N_29092,N_29978);
and UO_1842 (O_1842,N_29053,N_29099);
and UO_1843 (O_1843,N_29801,N_29832);
nor UO_1844 (O_1844,N_29780,N_29472);
nand UO_1845 (O_1845,N_29950,N_29489);
nor UO_1846 (O_1846,N_29510,N_29622);
or UO_1847 (O_1847,N_29963,N_29155);
or UO_1848 (O_1848,N_29340,N_29170);
xnor UO_1849 (O_1849,N_29739,N_29284);
nor UO_1850 (O_1850,N_29931,N_29447);
and UO_1851 (O_1851,N_29001,N_29132);
and UO_1852 (O_1852,N_29158,N_29764);
and UO_1853 (O_1853,N_29961,N_29158);
xor UO_1854 (O_1854,N_29879,N_29861);
and UO_1855 (O_1855,N_29465,N_29974);
and UO_1856 (O_1856,N_29543,N_29209);
nand UO_1857 (O_1857,N_29261,N_29169);
nand UO_1858 (O_1858,N_29582,N_29859);
or UO_1859 (O_1859,N_29695,N_29507);
nand UO_1860 (O_1860,N_29155,N_29218);
and UO_1861 (O_1861,N_29483,N_29588);
nand UO_1862 (O_1862,N_29034,N_29811);
or UO_1863 (O_1863,N_29177,N_29710);
xor UO_1864 (O_1864,N_29732,N_29250);
and UO_1865 (O_1865,N_29305,N_29050);
xor UO_1866 (O_1866,N_29244,N_29957);
or UO_1867 (O_1867,N_29098,N_29420);
nor UO_1868 (O_1868,N_29713,N_29183);
nor UO_1869 (O_1869,N_29471,N_29835);
xor UO_1870 (O_1870,N_29671,N_29093);
nand UO_1871 (O_1871,N_29497,N_29945);
and UO_1872 (O_1872,N_29742,N_29116);
and UO_1873 (O_1873,N_29959,N_29068);
xor UO_1874 (O_1874,N_29431,N_29255);
nor UO_1875 (O_1875,N_29320,N_29899);
nand UO_1876 (O_1876,N_29503,N_29445);
or UO_1877 (O_1877,N_29354,N_29702);
nor UO_1878 (O_1878,N_29363,N_29996);
and UO_1879 (O_1879,N_29423,N_29892);
and UO_1880 (O_1880,N_29185,N_29112);
xnor UO_1881 (O_1881,N_29329,N_29689);
or UO_1882 (O_1882,N_29497,N_29649);
or UO_1883 (O_1883,N_29417,N_29188);
and UO_1884 (O_1884,N_29414,N_29217);
nor UO_1885 (O_1885,N_29038,N_29389);
nor UO_1886 (O_1886,N_29432,N_29997);
and UO_1887 (O_1887,N_29233,N_29912);
or UO_1888 (O_1888,N_29855,N_29906);
or UO_1889 (O_1889,N_29433,N_29510);
nor UO_1890 (O_1890,N_29755,N_29243);
xnor UO_1891 (O_1891,N_29556,N_29109);
xnor UO_1892 (O_1892,N_29300,N_29328);
nand UO_1893 (O_1893,N_29584,N_29763);
nand UO_1894 (O_1894,N_29126,N_29298);
nor UO_1895 (O_1895,N_29072,N_29183);
nor UO_1896 (O_1896,N_29967,N_29165);
nand UO_1897 (O_1897,N_29488,N_29133);
and UO_1898 (O_1898,N_29242,N_29381);
xor UO_1899 (O_1899,N_29027,N_29510);
or UO_1900 (O_1900,N_29767,N_29789);
nor UO_1901 (O_1901,N_29984,N_29819);
nor UO_1902 (O_1902,N_29195,N_29967);
or UO_1903 (O_1903,N_29192,N_29202);
xor UO_1904 (O_1904,N_29962,N_29174);
and UO_1905 (O_1905,N_29295,N_29816);
xor UO_1906 (O_1906,N_29449,N_29331);
and UO_1907 (O_1907,N_29099,N_29502);
nand UO_1908 (O_1908,N_29777,N_29691);
nand UO_1909 (O_1909,N_29152,N_29710);
and UO_1910 (O_1910,N_29848,N_29572);
xnor UO_1911 (O_1911,N_29350,N_29806);
and UO_1912 (O_1912,N_29158,N_29005);
nor UO_1913 (O_1913,N_29636,N_29095);
or UO_1914 (O_1914,N_29015,N_29677);
or UO_1915 (O_1915,N_29145,N_29337);
and UO_1916 (O_1916,N_29160,N_29989);
xor UO_1917 (O_1917,N_29113,N_29179);
or UO_1918 (O_1918,N_29468,N_29565);
nor UO_1919 (O_1919,N_29821,N_29519);
or UO_1920 (O_1920,N_29359,N_29224);
nand UO_1921 (O_1921,N_29620,N_29501);
nand UO_1922 (O_1922,N_29399,N_29517);
and UO_1923 (O_1923,N_29400,N_29020);
xor UO_1924 (O_1924,N_29198,N_29990);
or UO_1925 (O_1925,N_29885,N_29752);
nor UO_1926 (O_1926,N_29273,N_29284);
xnor UO_1927 (O_1927,N_29778,N_29398);
nor UO_1928 (O_1928,N_29430,N_29346);
xor UO_1929 (O_1929,N_29370,N_29586);
nor UO_1930 (O_1930,N_29675,N_29815);
nor UO_1931 (O_1931,N_29763,N_29937);
xnor UO_1932 (O_1932,N_29214,N_29900);
or UO_1933 (O_1933,N_29955,N_29608);
and UO_1934 (O_1934,N_29244,N_29543);
or UO_1935 (O_1935,N_29037,N_29525);
xnor UO_1936 (O_1936,N_29939,N_29321);
nor UO_1937 (O_1937,N_29411,N_29504);
xnor UO_1938 (O_1938,N_29338,N_29854);
nor UO_1939 (O_1939,N_29151,N_29275);
and UO_1940 (O_1940,N_29927,N_29760);
or UO_1941 (O_1941,N_29240,N_29223);
nand UO_1942 (O_1942,N_29992,N_29698);
nand UO_1943 (O_1943,N_29683,N_29518);
nor UO_1944 (O_1944,N_29853,N_29118);
nor UO_1945 (O_1945,N_29272,N_29799);
nor UO_1946 (O_1946,N_29416,N_29393);
xnor UO_1947 (O_1947,N_29970,N_29608);
nor UO_1948 (O_1948,N_29055,N_29118);
or UO_1949 (O_1949,N_29234,N_29690);
nor UO_1950 (O_1950,N_29754,N_29255);
xnor UO_1951 (O_1951,N_29861,N_29719);
nor UO_1952 (O_1952,N_29740,N_29492);
xnor UO_1953 (O_1953,N_29680,N_29242);
xor UO_1954 (O_1954,N_29458,N_29311);
xor UO_1955 (O_1955,N_29812,N_29994);
or UO_1956 (O_1956,N_29462,N_29677);
and UO_1957 (O_1957,N_29852,N_29664);
xnor UO_1958 (O_1958,N_29012,N_29378);
nand UO_1959 (O_1959,N_29494,N_29319);
nand UO_1960 (O_1960,N_29455,N_29215);
xnor UO_1961 (O_1961,N_29613,N_29792);
nor UO_1962 (O_1962,N_29358,N_29452);
or UO_1963 (O_1963,N_29005,N_29325);
and UO_1964 (O_1964,N_29078,N_29446);
nand UO_1965 (O_1965,N_29163,N_29768);
nor UO_1966 (O_1966,N_29544,N_29561);
nand UO_1967 (O_1967,N_29885,N_29325);
or UO_1968 (O_1968,N_29499,N_29934);
nand UO_1969 (O_1969,N_29211,N_29469);
nand UO_1970 (O_1970,N_29745,N_29709);
or UO_1971 (O_1971,N_29204,N_29391);
nor UO_1972 (O_1972,N_29834,N_29632);
or UO_1973 (O_1973,N_29340,N_29938);
and UO_1974 (O_1974,N_29887,N_29412);
xor UO_1975 (O_1975,N_29454,N_29099);
and UO_1976 (O_1976,N_29385,N_29080);
nor UO_1977 (O_1977,N_29078,N_29084);
or UO_1978 (O_1978,N_29397,N_29633);
xor UO_1979 (O_1979,N_29897,N_29811);
and UO_1980 (O_1980,N_29738,N_29826);
nand UO_1981 (O_1981,N_29769,N_29434);
xnor UO_1982 (O_1982,N_29852,N_29211);
nand UO_1983 (O_1983,N_29903,N_29841);
nand UO_1984 (O_1984,N_29861,N_29756);
and UO_1985 (O_1985,N_29243,N_29870);
xnor UO_1986 (O_1986,N_29866,N_29139);
and UO_1987 (O_1987,N_29399,N_29554);
xor UO_1988 (O_1988,N_29974,N_29976);
nor UO_1989 (O_1989,N_29241,N_29283);
and UO_1990 (O_1990,N_29413,N_29322);
nor UO_1991 (O_1991,N_29253,N_29987);
nand UO_1992 (O_1992,N_29099,N_29210);
or UO_1993 (O_1993,N_29401,N_29248);
and UO_1994 (O_1994,N_29778,N_29329);
xor UO_1995 (O_1995,N_29919,N_29941);
and UO_1996 (O_1996,N_29857,N_29160);
or UO_1997 (O_1997,N_29280,N_29165);
or UO_1998 (O_1998,N_29997,N_29619);
xnor UO_1999 (O_1999,N_29958,N_29726);
or UO_2000 (O_2000,N_29454,N_29620);
nand UO_2001 (O_2001,N_29316,N_29810);
nor UO_2002 (O_2002,N_29212,N_29864);
nor UO_2003 (O_2003,N_29293,N_29310);
or UO_2004 (O_2004,N_29621,N_29789);
nor UO_2005 (O_2005,N_29379,N_29285);
and UO_2006 (O_2006,N_29622,N_29977);
nor UO_2007 (O_2007,N_29920,N_29668);
and UO_2008 (O_2008,N_29227,N_29830);
nand UO_2009 (O_2009,N_29525,N_29813);
or UO_2010 (O_2010,N_29672,N_29140);
nand UO_2011 (O_2011,N_29315,N_29104);
and UO_2012 (O_2012,N_29730,N_29270);
and UO_2013 (O_2013,N_29671,N_29829);
or UO_2014 (O_2014,N_29608,N_29143);
nor UO_2015 (O_2015,N_29426,N_29932);
nor UO_2016 (O_2016,N_29198,N_29290);
nand UO_2017 (O_2017,N_29480,N_29524);
nand UO_2018 (O_2018,N_29348,N_29160);
xnor UO_2019 (O_2019,N_29096,N_29007);
or UO_2020 (O_2020,N_29252,N_29172);
or UO_2021 (O_2021,N_29039,N_29231);
nand UO_2022 (O_2022,N_29531,N_29225);
and UO_2023 (O_2023,N_29036,N_29362);
or UO_2024 (O_2024,N_29209,N_29323);
nor UO_2025 (O_2025,N_29327,N_29380);
and UO_2026 (O_2026,N_29287,N_29339);
nor UO_2027 (O_2027,N_29958,N_29895);
xnor UO_2028 (O_2028,N_29990,N_29181);
nand UO_2029 (O_2029,N_29708,N_29862);
xnor UO_2030 (O_2030,N_29123,N_29469);
and UO_2031 (O_2031,N_29025,N_29085);
nand UO_2032 (O_2032,N_29327,N_29433);
or UO_2033 (O_2033,N_29212,N_29751);
xnor UO_2034 (O_2034,N_29335,N_29348);
xor UO_2035 (O_2035,N_29032,N_29405);
xnor UO_2036 (O_2036,N_29998,N_29341);
xnor UO_2037 (O_2037,N_29539,N_29828);
or UO_2038 (O_2038,N_29991,N_29698);
nand UO_2039 (O_2039,N_29702,N_29229);
xnor UO_2040 (O_2040,N_29092,N_29735);
xor UO_2041 (O_2041,N_29630,N_29791);
xnor UO_2042 (O_2042,N_29994,N_29063);
nand UO_2043 (O_2043,N_29644,N_29963);
or UO_2044 (O_2044,N_29786,N_29433);
xnor UO_2045 (O_2045,N_29488,N_29738);
and UO_2046 (O_2046,N_29212,N_29239);
xor UO_2047 (O_2047,N_29135,N_29062);
nor UO_2048 (O_2048,N_29334,N_29709);
and UO_2049 (O_2049,N_29261,N_29959);
nand UO_2050 (O_2050,N_29980,N_29673);
or UO_2051 (O_2051,N_29656,N_29889);
and UO_2052 (O_2052,N_29510,N_29208);
nor UO_2053 (O_2053,N_29216,N_29103);
and UO_2054 (O_2054,N_29823,N_29536);
or UO_2055 (O_2055,N_29776,N_29183);
xnor UO_2056 (O_2056,N_29427,N_29332);
nor UO_2057 (O_2057,N_29613,N_29999);
and UO_2058 (O_2058,N_29749,N_29959);
nor UO_2059 (O_2059,N_29252,N_29768);
xor UO_2060 (O_2060,N_29512,N_29188);
or UO_2061 (O_2061,N_29850,N_29340);
or UO_2062 (O_2062,N_29003,N_29106);
and UO_2063 (O_2063,N_29043,N_29403);
nand UO_2064 (O_2064,N_29417,N_29678);
nand UO_2065 (O_2065,N_29988,N_29973);
xor UO_2066 (O_2066,N_29644,N_29048);
and UO_2067 (O_2067,N_29705,N_29340);
and UO_2068 (O_2068,N_29602,N_29024);
and UO_2069 (O_2069,N_29153,N_29902);
nor UO_2070 (O_2070,N_29247,N_29298);
and UO_2071 (O_2071,N_29901,N_29474);
nand UO_2072 (O_2072,N_29724,N_29193);
nand UO_2073 (O_2073,N_29906,N_29229);
nand UO_2074 (O_2074,N_29832,N_29135);
nand UO_2075 (O_2075,N_29834,N_29506);
or UO_2076 (O_2076,N_29992,N_29951);
nor UO_2077 (O_2077,N_29582,N_29877);
xor UO_2078 (O_2078,N_29047,N_29269);
nor UO_2079 (O_2079,N_29238,N_29381);
nor UO_2080 (O_2080,N_29275,N_29853);
nor UO_2081 (O_2081,N_29985,N_29022);
nand UO_2082 (O_2082,N_29545,N_29288);
nand UO_2083 (O_2083,N_29982,N_29701);
nor UO_2084 (O_2084,N_29844,N_29254);
nor UO_2085 (O_2085,N_29143,N_29370);
or UO_2086 (O_2086,N_29266,N_29722);
nor UO_2087 (O_2087,N_29296,N_29631);
nor UO_2088 (O_2088,N_29322,N_29044);
xor UO_2089 (O_2089,N_29838,N_29482);
and UO_2090 (O_2090,N_29214,N_29424);
xnor UO_2091 (O_2091,N_29889,N_29169);
or UO_2092 (O_2092,N_29046,N_29827);
xnor UO_2093 (O_2093,N_29254,N_29663);
xnor UO_2094 (O_2094,N_29136,N_29087);
xor UO_2095 (O_2095,N_29921,N_29777);
xor UO_2096 (O_2096,N_29134,N_29707);
nand UO_2097 (O_2097,N_29435,N_29888);
nor UO_2098 (O_2098,N_29273,N_29139);
or UO_2099 (O_2099,N_29789,N_29892);
or UO_2100 (O_2100,N_29031,N_29360);
or UO_2101 (O_2101,N_29172,N_29370);
or UO_2102 (O_2102,N_29621,N_29633);
and UO_2103 (O_2103,N_29867,N_29247);
or UO_2104 (O_2104,N_29911,N_29849);
nor UO_2105 (O_2105,N_29967,N_29182);
xnor UO_2106 (O_2106,N_29369,N_29049);
nor UO_2107 (O_2107,N_29036,N_29117);
and UO_2108 (O_2108,N_29677,N_29570);
nor UO_2109 (O_2109,N_29517,N_29024);
nand UO_2110 (O_2110,N_29509,N_29658);
nor UO_2111 (O_2111,N_29874,N_29428);
xor UO_2112 (O_2112,N_29339,N_29189);
and UO_2113 (O_2113,N_29474,N_29108);
nand UO_2114 (O_2114,N_29941,N_29429);
and UO_2115 (O_2115,N_29066,N_29012);
nand UO_2116 (O_2116,N_29869,N_29291);
and UO_2117 (O_2117,N_29688,N_29388);
nor UO_2118 (O_2118,N_29090,N_29825);
or UO_2119 (O_2119,N_29194,N_29834);
nor UO_2120 (O_2120,N_29805,N_29292);
nor UO_2121 (O_2121,N_29221,N_29418);
or UO_2122 (O_2122,N_29906,N_29259);
or UO_2123 (O_2123,N_29271,N_29968);
xor UO_2124 (O_2124,N_29826,N_29753);
or UO_2125 (O_2125,N_29641,N_29495);
nor UO_2126 (O_2126,N_29637,N_29493);
or UO_2127 (O_2127,N_29123,N_29935);
nor UO_2128 (O_2128,N_29990,N_29227);
nand UO_2129 (O_2129,N_29729,N_29044);
xor UO_2130 (O_2130,N_29593,N_29351);
xor UO_2131 (O_2131,N_29442,N_29267);
nor UO_2132 (O_2132,N_29435,N_29654);
and UO_2133 (O_2133,N_29134,N_29261);
nor UO_2134 (O_2134,N_29525,N_29044);
or UO_2135 (O_2135,N_29042,N_29465);
or UO_2136 (O_2136,N_29079,N_29212);
or UO_2137 (O_2137,N_29122,N_29154);
nand UO_2138 (O_2138,N_29122,N_29069);
nor UO_2139 (O_2139,N_29347,N_29662);
and UO_2140 (O_2140,N_29751,N_29672);
or UO_2141 (O_2141,N_29408,N_29872);
or UO_2142 (O_2142,N_29607,N_29390);
nor UO_2143 (O_2143,N_29571,N_29336);
nand UO_2144 (O_2144,N_29060,N_29535);
and UO_2145 (O_2145,N_29350,N_29762);
xnor UO_2146 (O_2146,N_29613,N_29905);
nand UO_2147 (O_2147,N_29525,N_29179);
and UO_2148 (O_2148,N_29898,N_29450);
nor UO_2149 (O_2149,N_29553,N_29195);
and UO_2150 (O_2150,N_29009,N_29308);
nor UO_2151 (O_2151,N_29730,N_29633);
nor UO_2152 (O_2152,N_29439,N_29170);
and UO_2153 (O_2153,N_29660,N_29394);
or UO_2154 (O_2154,N_29728,N_29267);
nand UO_2155 (O_2155,N_29412,N_29610);
nor UO_2156 (O_2156,N_29739,N_29484);
and UO_2157 (O_2157,N_29602,N_29441);
or UO_2158 (O_2158,N_29014,N_29346);
xor UO_2159 (O_2159,N_29789,N_29870);
nor UO_2160 (O_2160,N_29666,N_29401);
nand UO_2161 (O_2161,N_29439,N_29414);
nand UO_2162 (O_2162,N_29730,N_29714);
nor UO_2163 (O_2163,N_29584,N_29630);
xor UO_2164 (O_2164,N_29287,N_29808);
or UO_2165 (O_2165,N_29841,N_29746);
nand UO_2166 (O_2166,N_29591,N_29124);
xor UO_2167 (O_2167,N_29629,N_29319);
nand UO_2168 (O_2168,N_29377,N_29565);
and UO_2169 (O_2169,N_29573,N_29560);
nor UO_2170 (O_2170,N_29528,N_29534);
xor UO_2171 (O_2171,N_29468,N_29529);
and UO_2172 (O_2172,N_29690,N_29797);
or UO_2173 (O_2173,N_29114,N_29172);
or UO_2174 (O_2174,N_29314,N_29026);
nor UO_2175 (O_2175,N_29105,N_29964);
nor UO_2176 (O_2176,N_29853,N_29943);
or UO_2177 (O_2177,N_29420,N_29450);
nand UO_2178 (O_2178,N_29119,N_29750);
or UO_2179 (O_2179,N_29894,N_29013);
nor UO_2180 (O_2180,N_29098,N_29482);
and UO_2181 (O_2181,N_29543,N_29757);
nand UO_2182 (O_2182,N_29152,N_29702);
xor UO_2183 (O_2183,N_29368,N_29542);
xnor UO_2184 (O_2184,N_29346,N_29748);
and UO_2185 (O_2185,N_29347,N_29992);
xnor UO_2186 (O_2186,N_29752,N_29313);
nor UO_2187 (O_2187,N_29902,N_29631);
nand UO_2188 (O_2188,N_29987,N_29043);
and UO_2189 (O_2189,N_29909,N_29802);
or UO_2190 (O_2190,N_29679,N_29011);
nor UO_2191 (O_2191,N_29718,N_29673);
nand UO_2192 (O_2192,N_29871,N_29267);
xor UO_2193 (O_2193,N_29905,N_29943);
and UO_2194 (O_2194,N_29497,N_29401);
xnor UO_2195 (O_2195,N_29636,N_29355);
xnor UO_2196 (O_2196,N_29513,N_29291);
or UO_2197 (O_2197,N_29835,N_29804);
nand UO_2198 (O_2198,N_29451,N_29858);
nor UO_2199 (O_2199,N_29303,N_29526);
nand UO_2200 (O_2200,N_29917,N_29951);
xor UO_2201 (O_2201,N_29754,N_29471);
and UO_2202 (O_2202,N_29222,N_29975);
and UO_2203 (O_2203,N_29523,N_29289);
and UO_2204 (O_2204,N_29082,N_29147);
xnor UO_2205 (O_2205,N_29560,N_29115);
xor UO_2206 (O_2206,N_29403,N_29912);
or UO_2207 (O_2207,N_29853,N_29365);
or UO_2208 (O_2208,N_29109,N_29856);
xor UO_2209 (O_2209,N_29737,N_29661);
xor UO_2210 (O_2210,N_29757,N_29486);
xnor UO_2211 (O_2211,N_29811,N_29788);
nor UO_2212 (O_2212,N_29761,N_29206);
or UO_2213 (O_2213,N_29316,N_29700);
xor UO_2214 (O_2214,N_29677,N_29568);
or UO_2215 (O_2215,N_29525,N_29368);
and UO_2216 (O_2216,N_29814,N_29249);
or UO_2217 (O_2217,N_29732,N_29507);
and UO_2218 (O_2218,N_29870,N_29103);
nand UO_2219 (O_2219,N_29608,N_29572);
nor UO_2220 (O_2220,N_29717,N_29134);
xnor UO_2221 (O_2221,N_29159,N_29351);
xor UO_2222 (O_2222,N_29022,N_29095);
and UO_2223 (O_2223,N_29859,N_29948);
nor UO_2224 (O_2224,N_29888,N_29746);
nand UO_2225 (O_2225,N_29401,N_29091);
nand UO_2226 (O_2226,N_29183,N_29695);
or UO_2227 (O_2227,N_29800,N_29845);
or UO_2228 (O_2228,N_29870,N_29053);
and UO_2229 (O_2229,N_29504,N_29799);
xnor UO_2230 (O_2230,N_29600,N_29360);
or UO_2231 (O_2231,N_29652,N_29107);
nor UO_2232 (O_2232,N_29977,N_29572);
xor UO_2233 (O_2233,N_29010,N_29979);
nor UO_2234 (O_2234,N_29452,N_29840);
and UO_2235 (O_2235,N_29502,N_29122);
or UO_2236 (O_2236,N_29151,N_29350);
and UO_2237 (O_2237,N_29554,N_29761);
and UO_2238 (O_2238,N_29827,N_29750);
or UO_2239 (O_2239,N_29141,N_29469);
and UO_2240 (O_2240,N_29939,N_29801);
or UO_2241 (O_2241,N_29344,N_29793);
nor UO_2242 (O_2242,N_29935,N_29972);
nand UO_2243 (O_2243,N_29341,N_29100);
and UO_2244 (O_2244,N_29788,N_29705);
and UO_2245 (O_2245,N_29064,N_29524);
nand UO_2246 (O_2246,N_29470,N_29582);
nand UO_2247 (O_2247,N_29359,N_29905);
and UO_2248 (O_2248,N_29241,N_29046);
or UO_2249 (O_2249,N_29444,N_29249);
and UO_2250 (O_2250,N_29159,N_29026);
nand UO_2251 (O_2251,N_29589,N_29300);
xor UO_2252 (O_2252,N_29784,N_29472);
nand UO_2253 (O_2253,N_29531,N_29170);
nor UO_2254 (O_2254,N_29297,N_29986);
xnor UO_2255 (O_2255,N_29412,N_29160);
and UO_2256 (O_2256,N_29277,N_29118);
xnor UO_2257 (O_2257,N_29023,N_29914);
and UO_2258 (O_2258,N_29646,N_29743);
nand UO_2259 (O_2259,N_29951,N_29919);
or UO_2260 (O_2260,N_29631,N_29138);
xnor UO_2261 (O_2261,N_29238,N_29932);
and UO_2262 (O_2262,N_29152,N_29128);
and UO_2263 (O_2263,N_29633,N_29847);
xnor UO_2264 (O_2264,N_29453,N_29254);
nor UO_2265 (O_2265,N_29266,N_29306);
or UO_2266 (O_2266,N_29809,N_29149);
nand UO_2267 (O_2267,N_29976,N_29668);
and UO_2268 (O_2268,N_29189,N_29015);
or UO_2269 (O_2269,N_29081,N_29926);
and UO_2270 (O_2270,N_29422,N_29130);
nand UO_2271 (O_2271,N_29732,N_29904);
xor UO_2272 (O_2272,N_29687,N_29973);
or UO_2273 (O_2273,N_29965,N_29450);
xor UO_2274 (O_2274,N_29431,N_29793);
nand UO_2275 (O_2275,N_29686,N_29349);
nand UO_2276 (O_2276,N_29497,N_29176);
nor UO_2277 (O_2277,N_29208,N_29127);
xnor UO_2278 (O_2278,N_29968,N_29666);
and UO_2279 (O_2279,N_29882,N_29366);
nand UO_2280 (O_2280,N_29100,N_29770);
or UO_2281 (O_2281,N_29989,N_29072);
nor UO_2282 (O_2282,N_29476,N_29289);
and UO_2283 (O_2283,N_29479,N_29899);
nand UO_2284 (O_2284,N_29796,N_29729);
xor UO_2285 (O_2285,N_29343,N_29198);
nor UO_2286 (O_2286,N_29889,N_29405);
or UO_2287 (O_2287,N_29550,N_29333);
or UO_2288 (O_2288,N_29816,N_29304);
or UO_2289 (O_2289,N_29967,N_29537);
and UO_2290 (O_2290,N_29975,N_29562);
and UO_2291 (O_2291,N_29083,N_29480);
xor UO_2292 (O_2292,N_29086,N_29027);
nand UO_2293 (O_2293,N_29522,N_29380);
or UO_2294 (O_2294,N_29269,N_29497);
nand UO_2295 (O_2295,N_29559,N_29507);
and UO_2296 (O_2296,N_29478,N_29097);
nand UO_2297 (O_2297,N_29961,N_29766);
and UO_2298 (O_2298,N_29333,N_29474);
xnor UO_2299 (O_2299,N_29535,N_29530);
and UO_2300 (O_2300,N_29365,N_29828);
nor UO_2301 (O_2301,N_29791,N_29297);
nand UO_2302 (O_2302,N_29810,N_29395);
nand UO_2303 (O_2303,N_29692,N_29787);
and UO_2304 (O_2304,N_29620,N_29964);
xnor UO_2305 (O_2305,N_29647,N_29351);
and UO_2306 (O_2306,N_29082,N_29781);
nand UO_2307 (O_2307,N_29366,N_29496);
nor UO_2308 (O_2308,N_29894,N_29698);
xnor UO_2309 (O_2309,N_29789,N_29412);
nand UO_2310 (O_2310,N_29031,N_29050);
nor UO_2311 (O_2311,N_29415,N_29138);
or UO_2312 (O_2312,N_29780,N_29059);
and UO_2313 (O_2313,N_29833,N_29616);
or UO_2314 (O_2314,N_29724,N_29617);
xnor UO_2315 (O_2315,N_29561,N_29630);
nor UO_2316 (O_2316,N_29109,N_29153);
or UO_2317 (O_2317,N_29891,N_29239);
xnor UO_2318 (O_2318,N_29598,N_29595);
nand UO_2319 (O_2319,N_29888,N_29847);
xnor UO_2320 (O_2320,N_29172,N_29901);
xor UO_2321 (O_2321,N_29618,N_29344);
xnor UO_2322 (O_2322,N_29753,N_29858);
nor UO_2323 (O_2323,N_29883,N_29204);
nand UO_2324 (O_2324,N_29759,N_29657);
xnor UO_2325 (O_2325,N_29627,N_29442);
and UO_2326 (O_2326,N_29626,N_29819);
nand UO_2327 (O_2327,N_29770,N_29473);
nor UO_2328 (O_2328,N_29337,N_29841);
nor UO_2329 (O_2329,N_29157,N_29400);
nor UO_2330 (O_2330,N_29762,N_29952);
nand UO_2331 (O_2331,N_29223,N_29681);
nor UO_2332 (O_2332,N_29017,N_29054);
nor UO_2333 (O_2333,N_29123,N_29714);
xor UO_2334 (O_2334,N_29698,N_29361);
nand UO_2335 (O_2335,N_29261,N_29245);
nor UO_2336 (O_2336,N_29699,N_29333);
or UO_2337 (O_2337,N_29543,N_29102);
and UO_2338 (O_2338,N_29009,N_29595);
or UO_2339 (O_2339,N_29975,N_29188);
nor UO_2340 (O_2340,N_29858,N_29516);
nor UO_2341 (O_2341,N_29836,N_29060);
and UO_2342 (O_2342,N_29678,N_29545);
xnor UO_2343 (O_2343,N_29976,N_29296);
nor UO_2344 (O_2344,N_29091,N_29271);
nand UO_2345 (O_2345,N_29261,N_29256);
nor UO_2346 (O_2346,N_29711,N_29063);
and UO_2347 (O_2347,N_29362,N_29623);
nand UO_2348 (O_2348,N_29466,N_29751);
and UO_2349 (O_2349,N_29303,N_29826);
and UO_2350 (O_2350,N_29218,N_29276);
or UO_2351 (O_2351,N_29027,N_29162);
and UO_2352 (O_2352,N_29793,N_29325);
or UO_2353 (O_2353,N_29568,N_29065);
xor UO_2354 (O_2354,N_29776,N_29576);
or UO_2355 (O_2355,N_29613,N_29102);
xnor UO_2356 (O_2356,N_29398,N_29936);
nor UO_2357 (O_2357,N_29902,N_29154);
xnor UO_2358 (O_2358,N_29761,N_29759);
xnor UO_2359 (O_2359,N_29161,N_29837);
nor UO_2360 (O_2360,N_29761,N_29711);
or UO_2361 (O_2361,N_29920,N_29098);
or UO_2362 (O_2362,N_29826,N_29618);
nor UO_2363 (O_2363,N_29684,N_29467);
nand UO_2364 (O_2364,N_29871,N_29187);
and UO_2365 (O_2365,N_29238,N_29184);
nand UO_2366 (O_2366,N_29074,N_29468);
nor UO_2367 (O_2367,N_29848,N_29748);
nor UO_2368 (O_2368,N_29155,N_29736);
xor UO_2369 (O_2369,N_29429,N_29811);
nand UO_2370 (O_2370,N_29730,N_29990);
and UO_2371 (O_2371,N_29890,N_29165);
nor UO_2372 (O_2372,N_29768,N_29406);
and UO_2373 (O_2373,N_29301,N_29680);
and UO_2374 (O_2374,N_29073,N_29818);
xnor UO_2375 (O_2375,N_29712,N_29389);
and UO_2376 (O_2376,N_29742,N_29210);
nor UO_2377 (O_2377,N_29127,N_29885);
nand UO_2378 (O_2378,N_29909,N_29680);
nor UO_2379 (O_2379,N_29273,N_29210);
xor UO_2380 (O_2380,N_29077,N_29608);
nand UO_2381 (O_2381,N_29943,N_29385);
and UO_2382 (O_2382,N_29433,N_29843);
xor UO_2383 (O_2383,N_29963,N_29258);
nor UO_2384 (O_2384,N_29866,N_29242);
or UO_2385 (O_2385,N_29927,N_29791);
nor UO_2386 (O_2386,N_29106,N_29855);
xor UO_2387 (O_2387,N_29422,N_29792);
xor UO_2388 (O_2388,N_29543,N_29229);
nor UO_2389 (O_2389,N_29798,N_29287);
xnor UO_2390 (O_2390,N_29763,N_29610);
nor UO_2391 (O_2391,N_29800,N_29251);
nand UO_2392 (O_2392,N_29110,N_29809);
nand UO_2393 (O_2393,N_29498,N_29818);
xor UO_2394 (O_2394,N_29808,N_29280);
and UO_2395 (O_2395,N_29872,N_29789);
and UO_2396 (O_2396,N_29914,N_29759);
nor UO_2397 (O_2397,N_29624,N_29075);
or UO_2398 (O_2398,N_29622,N_29642);
xnor UO_2399 (O_2399,N_29333,N_29669);
nor UO_2400 (O_2400,N_29292,N_29823);
nand UO_2401 (O_2401,N_29686,N_29751);
xnor UO_2402 (O_2402,N_29619,N_29409);
xor UO_2403 (O_2403,N_29529,N_29883);
xor UO_2404 (O_2404,N_29833,N_29790);
and UO_2405 (O_2405,N_29849,N_29382);
or UO_2406 (O_2406,N_29373,N_29884);
nand UO_2407 (O_2407,N_29632,N_29208);
nand UO_2408 (O_2408,N_29703,N_29614);
xnor UO_2409 (O_2409,N_29040,N_29519);
nor UO_2410 (O_2410,N_29116,N_29880);
xor UO_2411 (O_2411,N_29209,N_29829);
and UO_2412 (O_2412,N_29668,N_29337);
nor UO_2413 (O_2413,N_29648,N_29385);
nand UO_2414 (O_2414,N_29318,N_29484);
nor UO_2415 (O_2415,N_29861,N_29442);
nand UO_2416 (O_2416,N_29967,N_29902);
nor UO_2417 (O_2417,N_29961,N_29358);
nand UO_2418 (O_2418,N_29584,N_29622);
nor UO_2419 (O_2419,N_29706,N_29951);
nand UO_2420 (O_2420,N_29448,N_29189);
nor UO_2421 (O_2421,N_29600,N_29140);
nor UO_2422 (O_2422,N_29816,N_29197);
xnor UO_2423 (O_2423,N_29563,N_29131);
xor UO_2424 (O_2424,N_29242,N_29098);
xor UO_2425 (O_2425,N_29510,N_29438);
nand UO_2426 (O_2426,N_29922,N_29987);
xnor UO_2427 (O_2427,N_29554,N_29684);
or UO_2428 (O_2428,N_29133,N_29388);
nor UO_2429 (O_2429,N_29144,N_29775);
nor UO_2430 (O_2430,N_29102,N_29853);
xnor UO_2431 (O_2431,N_29288,N_29535);
and UO_2432 (O_2432,N_29285,N_29108);
or UO_2433 (O_2433,N_29472,N_29192);
xor UO_2434 (O_2434,N_29130,N_29473);
or UO_2435 (O_2435,N_29741,N_29025);
and UO_2436 (O_2436,N_29223,N_29878);
and UO_2437 (O_2437,N_29868,N_29897);
nand UO_2438 (O_2438,N_29265,N_29574);
xor UO_2439 (O_2439,N_29325,N_29554);
and UO_2440 (O_2440,N_29797,N_29721);
or UO_2441 (O_2441,N_29928,N_29907);
and UO_2442 (O_2442,N_29892,N_29335);
nor UO_2443 (O_2443,N_29687,N_29001);
and UO_2444 (O_2444,N_29174,N_29948);
xor UO_2445 (O_2445,N_29695,N_29598);
xor UO_2446 (O_2446,N_29742,N_29762);
nand UO_2447 (O_2447,N_29623,N_29981);
or UO_2448 (O_2448,N_29958,N_29080);
nor UO_2449 (O_2449,N_29898,N_29761);
xor UO_2450 (O_2450,N_29078,N_29321);
xor UO_2451 (O_2451,N_29437,N_29589);
and UO_2452 (O_2452,N_29841,N_29811);
nand UO_2453 (O_2453,N_29904,N_29638);
nand UO_2454 (O_2454,N_29900,N_29364);
xnor UO_2455 (O_2455,N_29830,N_29552);
nand UO_2456 (O_2456,N_29500,N_29453);
nand UO_2457 (O_2457,N_29472,N_29146);
and UO_2458 (O_2458,N_29788,N_29028);
nand UO_2459 (O_2459,N_29950,N_29297);
xor UO_2460 (O_2460,N_29836,N_29576);
nand UO_2461 (O_2461,N_29267,N_29907);
nand UO_2462 (O_2462,N_29493,N_29553);
xnor UO_2463 (O_2463,N_29079,N_29777);
nand UO_2464 (O_2464,N_29913,N_29328);
and UO_2465 (O_2465,N_29658,N_29919);
xor UO_2466 (O_2466,N_29308,N_29866);
xnor UO_2467 (O_2467,N_29543,N_29371);
nand UO_2468 (O_2468,N_29836,N_29501);
nor UO_2469 (O_2469,N_29141,N_29223);
nand UO_2470 (O_2470,N_29107,N_29966);
or UO_2471 (O_2471,N_29421,N_29523);
nor UO_2472 (O_2472,N_29129,N_29671);
nor UO_2473 (O_2473,N_29447,N_29619);
nor UO_2474 (O_2474,N_29309,N_29166);
xnor UO_2475 (O_2475,N_29213,N_29149);
and UO_2476 (O_2476,N_29536,N_29795);
nor UO_2477 (O_2477,N_29107,N_29398);
nand UO_2478 (O_2478,N_29260,N_29930);
nand UO_2479 (O_2479,N_29132,N_29851);
nand UO_2480 (O_2480,N_29356,N_29566);
or UO_2481 (O_2481,N_29926,N_29326);
nor UO_2482 (O_2482,N_29596,N_29903);
nand UO_2483 (O_2483,N_29857,N_29340);
or UO_2484 (O_2484,N_29804,N_29313);
nor UO_2485 (O_2485,N_29676,N_29982);
nand UO_2486 (O_2486,N_29717,N_29613);
xor UO_2487 (O_2487,N_29386,N_29877);
nand UO_2488 (O_2488,N_29675,N_29138);
xnor UO_2489 (O_2489,N_29811,N_29133);
xnor UO_2490 (O_2490,N_29017,N_29120);
or UO_2491 (O_2491,N_29687,N_29203);
or UO_2492 (O_2492,N_29052,N_29663);
or UO_2493 (O_2493,N_29821,N_29897);
nor UO_2494 (O_2494,N_29996,N_29159);
or UO_2495 (O_2495,N_29867,N_29966);
or UO_2496 (O_2496,N_29469,N_29038);
xor UO_2497 (O_2497,N_29647,N_29543);
nor UO_2498 (O_2498,N_29458,N_29241);
nor UO_2499 (O_2499,N_29207,N_29201);
and UO_2500 (O_2500,N_29335,N_29595);
xnor UO_2501 (O_2501,N_29080,N_29894);
and UO_2502 (O_2502,N_29643,N_29087);
or UO_2503 (O_2503,N_29414,N_29338);
nor UO_2504 (O_2504,N_29161,N_29626);
xnor UO_2505 (O_2505,N_29305,N_29079);
or UO_2506 (O_2506,N_29505,N_29211);
nand UO_2507 (O_2507,N_29075,N_29761);
nand UO_2508 (O_2508,N_29936,N_29744);
xnor UO_2509 (O_2509,N_29405,N_29300);
nand UO_2510 (O_2510,N_29230,N_29996);
and UO_2511 (O_2511,N_29919,N_29424);
or UO_2512 (O_2512,N_29525,N_29626);
and UO_2513 (O_2513,N_29607,N_29523);
xor UO_2514 (O_2514,N_29185,N_29435);
xor UO_2515 (O_2515,N_29017,N_29400);
nand UO_2516 (O_2516,N_29064,N_29770);
nor UO_2517 (O_2517,N_29373,N_29221);
or UO_2518 (O_2518,N_29310,N_29276);
or UO_2519 (O_2519,N_29498,N_29543);
nand UO_2520 (O_2520,N_29151,N_29864);
and UO_2521 (O_2521,N_29847,N_29113);
nand UO_2522 (O_2522,N_29501,N_29323);
nor UO_2523 (O_2523,N_29631,N_29198);
or UO_2524 (O_2524,N_29881,N_29101);
nor UO_2525 (O_2525,N_29903,N_29486);
and UO_2526 (O_2526,N_29938,N_29953);
and UO_2527 (O_2527,N_29700,N_29324);
and UO_2528 (O_2528,N_29190,N_29131);
or UO_2529 (O_2529,N_29468,N_29534);
and UO_2530 (O_2530,N_29029,N_29984);
or UO_2531 (O_2531,N_29708,N_29836);
nor UO_2532 (O_2532,N_29541,N_29253);
or UO_2533 (O_2533,N_29408,N_29817);
nor UO_2534 (O_2534,N_29295,N_29630);
nor UO_2535 (O_2535,N_29263,N_29882);
xnor UO_2536 (O_2536,N_29793,N_29258);
nor UO_2537 (O_2537,N_29541,N_29554);
xnor UO_2538 (O_2538,N_29421,N_29856);
xnor UO_2539 (O_2539,N_29209,N_29329);
xor UO_2540 (O_2540,N_29272,N_29601);
nand UO_2541 (O_2541,N_29881,N_29315);
nor UO_2542 (O_2542,N_29080,N_29549);
or UO_2543 (O_2543,N_29763,N_29541);
xor UO_2544 (O_2544,N_29406,N_29652);
and UO_2545 (O_2545,N_29427,N_29215);
nand UO_2546 (O_2546,N_29972,N_29172);
or UO_2547 (O_2547,N_29364,N_29286);
or UO_2548 (O_2548,N_29225,N_29056);
nor UO_2549 (O_2549,N_29154,N_29508);
and UO_2550 (O_2550,N_29830,N_29674);
and UO_2551 (O_2551,N_29882,N_29559);
xnor UO_2552 (O_2552,N_29800,N_29232);
or UO_2553 (O_2553,N_29966,N_29146);
and UO_2554 (O_2554,N_29226,N_29839);
nor UO_2555 (O_2555,N_29196,N_29311);
nor UO_2556 (O_2556,N_29079,N_29160);
nand UO_2557 (O_2557,N_29323,N_29957);
xnor UO_2558 (O_2558,N_29836,N_29703);
nor UO_2559 (O_2559,N_29112,N_29240);
xnor UO_2560 (O_2560,N_29063,N_29457);
xor UO_2561 (O_2561,N_29991,N_29519);
nand UO_2562 (O_2562,N_29202,N_29088);
nor UO_2563 (O_2563,N_29798,N_29059);
nand UO_2564 (O_2564,N_29257,N_29573);
xor UO_2565 (O_2565,N_29584,N_29871);
and UO_2566 (O_2566,N_29558,N_29814);
xor UO_2567 (O_2567,N_29143,N_29985);
nor UO_2568 (O_2568,N_29716,N_29655);
xnor UO_2569 (O_2569,N_29043,N_29264);
nor UO_2570 (O_2570,N_29588,N_29790);
and UO_2571 (O_2571,N_29452,N_29192);
nor UO_2572 (O_2572,N_29286,N_29776);
nor UO_2573 (O_2573,N_29141,N_29312);
or UO_2574 (O_2574,N_29636,N_29429);
or UO_2575 (O_2575,N_29586,N_29877);
xnor UO_2576 (O_2576,N_29941,N_29046);
xor UO_2577 (O_2577,N_29659,N_29018);
nand UO_2578 (O_2578,N_29633,N_29509);
nand UO_2579 (O_2579,N_29974,N_29644);
nand UO_2580 (O_2580,N_29983,N_29334);
nor UO_2581 (O_2581,N_29148,N_29888);
or UO_2582 (O_2582,N_29049,N_29149);
xnor UO_2583 (O_2583,N_29783,N_29328);
nor UO_2584 (O_2584,N_29446,N_29224);
xor UO_2585 (O_2585,N_29557,N_29507);
and UO_2586 (O_2586,N_29931,N_29370);
or UO_2587 (O_2587,N_29841,N_29156);
and UO_2588 (O_2588,N_29381,N_29342);
or UO_2589 (O_2589,N_29145,N_29852);
and UO_2590 (O_2590,N_29170,N_29910);
nor UO_2591 (O_2591,N_29957,N_29499);
or UO_2592 (O_2592,N_29080,N_29928);
xnor UO_2593 (O_2593,N_29920,N_29702);
or UO_2594 (O_2594,N_29808,N_29057);
or UO_2595 (O_2595,N_29938,N_29118);
or UO_2596 (O_2596,N_29162,N_29152);
and UO_2597 (O_2597,N_29978,N_29508);
and UO_2598 (O_2598,N_29021,N_29764);
nor UO_2599 (O_2599,N_29006,N_29581);
or UO_2600 (O_2600,N_29368,N_29591);
xnor UO_2601 (O_2601,N_29441,N_29019);
xor UO_2602 (O_2602,N_29250,N_29513);
xnor UO_2603 (O_2603,N_29156,N_29333);
nor UO_2604 (O_2604,N_29531,N_29408);
nor UO_2605 (O_2605,N_29843,N_29283);
or UO_2606 (O_2606,N_29731,N_29778);
nor UO_2607 (O_2607,N_29648,N_29155);
nand UO_2608 (O_2608,N_29507,N_29196);
or UO_2609 (O_2609,N_29604,N_29734);
nor UO_2610 (O_2610,N_29031,N_29603);
nand UO_2611 (O_2611,N_29601,N_29968);
nor UO_2612 (O_2612,N_29695,N_29075);
nand UO_2613 (O_2613,N_29283,N_29885);
xor UO_2614 (O_2614,N_29616,N_29150);
or UO_2615 (O_2615,N_29819,N_29156);
and UO_2616 (O_2616,N_29141,N_29457);
xnor UO_2617 (O_2617,N_29125,N_29894);
or UO_2618 (O_2618,N_29882,N_29089);
or UO_2619 (O_2619,N_29890,N_29124);
nor UO_2620 (O_2620,N_29525,N_29113);
and UO_2621 (O_2621,N_29104,N_29239);
nor UO_2622 (O_2622,N_29774,N_29083);
xnor UO_2623 (O_2623,N_29654,N_29518);
nand UO_2624 (O_2624,N_29119,N_29549);
nor UO_2625 (O_2625,N_29775,N_29925);
xnor UO_2626 (O_2626,N_29354,N_29606);
and UO_2627 (O_2627,N_29525,N_29443);
and UO_2628 (O_2628,N_29601,N_29439);
xor UO_2629 (O_2629,N_29944,N_29368);
and UO_2630 (O_2630,N_29157,N_29637);
nor UO_2631 (O_2631,N_29484,N_29036);
and UO_2632 (O_2632,N_29638,N_29554);
xnor UO_2633 (O_2633,N_29835,N_29356);
xnor UO_2634 (O_2634,N_29824,N_29616);
or UO_2635 (O_2635,N_29447,N_29397);
nand UO_2636 (O_2636,N_29214,N_29300);
nand UO_2637 (O_2637,N_29395,N_29695);
xor UO_2638 (O_2638,N_29340,N_29117);
nand UO_2639 (O_2639,N_29104,N_29350);
nand UO_2640 (O_2640,N_29498,N_29537);
and UO_2641 (O_2641,N_29238,N_29495);
nand UO_2642 (O_2642,N_29689,N_29953);
nor UO_2643 (O_2643,N_29099,N_29161);
xor UO_2644 (O_2644,N_29534,N_29879);
or UO_2645 (O_2645,N_29187,N_29782);
and UO_2646 (O_2646,N_29660,N_29111);
and UO_2647 (O_2647,N_29098,N_29178);
and UO_2648 (O_2648,N_29467,N_29710);
xor UO_2649 (O_2649,N_29768,N_29874);
nand UO_2650 (O_2650,N_29055,N_29501);
xor UO_2651 (O_2651,N_29060,N_29479);
nand UO_2652 (O_2652,N_29186,N_29742);
nand UO_2653 (O_2653,N_29391,N_29792);
xor UO_2654 (O_2654,N_29334,N_29216);
or UO_2655 (O_2655,N_29012,N_29000);
nor UO_2656 (O_2656,N_29296,N_29277);
and UO_2657 (O_2657,N_29576,N_29788);
nor UO_2658 (O_2658,N_29310,N_29095);
and UO_2659 (O_2659,N_29061,N_29644);
or UO_2660 (O_2660,N_29650,N_29367);
xor UO_2661 (O_2661,N_29980,N_29546);
and UO_2662 (O_2662,N_29626,N_29456);
xnor UO_2663 (O_2663,N_29102,N_29081);
nand UO_2664 (O_2664,N_29499,N_29853);
nor UO_2665 (O_2665,N_29552,N_29188);
nand UO_2666 (O_2666,N_29656,N_29364);
xnor UO_2667 (O_2667,N_29206,N_29892);
nor UO_2668 (O_2668,N_29927,N_29230);
nor UO_2669 (O_2669,N_29674,N_29859);
nand UO_2670 (O_2670,N_29463,N_29102);
xor UO_2671 (O_2671,N_29136,N_29125);
and UO_2672 (O_2672,N_29607,N_29278);
xnor UO_2673 (O_2673,N_29859,N_29777);
and UO_2674 (O_2674,N_29992,N_29654);
xor UO_2675 (O_2675,N_29674,N_29769);
xnor UO_2676 (O_2676,N_29750,N_29423);
xor UO_2677 (O_2677,N_29553,N_29591);
nand UO_2678 (O_2678,N_29557,N_29124);
nor UO_2679 (O_2679,N_29748,N_29214);
nor UO_2680 (O_2680,N_29926,N_29156);
and UO_2681 (O_2681,N_29120,N_29153);
and UO_2682 (O_2682,N_29422,N_29113);
nand UO_2683 (O_2683,N_29628,N_29350);
xor UO_2684 (O_2684,N_29403,N_29645);
nor UO_2685 (O_2685,N_29371,N_29763);
xnor UO_2686 (O_2686,N_29190,N_29262);
xor UO_2687 (O_2687,N_29024,N_29244);
xor UO_2688 (O_2688,N_29621,N_29051);
xnor UO_2689 (O_2689,N_29490,N_29294);
nand UO_2690 (O_2690,N_29346,N_29213);
xor UO_2691 (O_2691,N_29563,N_29584);
and UO_2692 (O_2692,N_29386,N_29808);
and UO_2693 (O_2693,N_29507,N_29881);
and UO_2694 (O_2694,N_29511,N_29273);
and UO_2695 (O_2695,N_29579,N_29750);
xnor UO_2696 (O_2696,N_29307,N_29346);
or UO_2697 (O_2697,N_29929,N_29739);
and UO_2698 (O_2698,N_29851,N_29002);
xor UO_2699 (O_2699,N_29805,N_29100);
and UO_2700 (O_2700,N_29692,N_29884);
or UO_2701 (O_2701,N_29003,N_29618);
xnor UO_2702 (O_2702,N_29052,N_29297);
nand UO_2703 (O_2703,N_29141,N_29365);
and UO_2704 (O_2704,N_29107,N_29094);
and UO_2705 (O_2705,N_29086,N_29322);
nor UO_2706 (O_2706,N_29143,N_29718);
and UO_2707 (O_2707,N_29988,N_29056);
nor UO_2708 (O_2708,N_29843,N_29071);
xor UO_2709 (O_2709,N_29816,N_29120);
nand UO_2710 (O_2710,N_29516,N_29235);
nand UO_2711 (O_2711,N_29017,N_29634);
and UO_2712 (O_2712,N_29307,N_29227);
or UO_2713 (O_2713,N_29189,N_29236);
and UO_2714 (O_2714,N_29834,N_29191);
xor UO_2715 (O_2715,N_29299,N_29391);
and UO_2716 (O_2716,N_29335,N_29317);
xor UO_2717 (O_2717,N_29009,N_29558);
or UO_2718 (O_2718,N_29841,N_29668);
and UO_2719 (O_2719,N_29812,N_29591);
nand UO_2720 (O_2720,N_29976,N_29225);
nor UO_2721 (O_2721,N_29148,N_29151);
xor UO_2722 (O_2722,N_29465,N_29259);
and UO_2723 (O_2723,N_29595,N_29377);
xor UO_2724 (O_2724,N_29750,N_29204);
nand UO_2725 (O_2725,N_29788,N_29876);
or UO_2726 (O_2726,N_29454,N_29539);
nor UO_2727 (O_2727,N_29495,N_29543);
xnor UO_2728 (O_2728,N_29106,N_29972);
nand UO_2729 (O_2729,N_29399,N_29930);
nand UO_2730 (O_2730,N_29740,N_29194);
or UO_2731 (O_2731,N_29266,N_29129);
xnor UO_2732 (O_2732,N_29236,N_29691);
nor UO_2733 (O_2733,N_29197,N_29385);
or UO_2734 (O_2734,N_29749,N_29578);
xnor UO_2735 (O_2735,N_29673,N_29537);
nand UO_2736 (O_2736,N_29040,N_29461);
xor UO_2737 (O_2737,N_29165,N_29238);
nand UO_2738 (O_2738,N_29143,N_29019);
and UO_2739 (O_2739,N_29122,N_29290);
nor UO_2740 (O_2740,N_29488,N_29470);
and UO_2741 (O_2741,N_29666,N_29161);
and UO_2742 (O_2742,N_29056,N_29271);
xnor UO_2743 (O_2743,N_29661,N_29898);
or UO_2744 (O_2744,N_29895,N_29780);
nand UO_2745 (O_2745,N_29147,N_29976);
or UO_2746 (O_2746,N_29260,N_29003);
nor UO_2747 (O_2747,N_29297,N_29538);
or UO_2748 (O_2748,N_29483,N_29437);
nor UO_2749 (O_2749,N_29907,N_29127);
and UO_2750 (O_2750,N_29424,N_29060);
or UO_2751 (O_2751,N_29815,N_29630);
and UO_2752 (O_2752,N_29480,N_29164);
nand UO_2753 (O_2753,N_29677,N_29838);
nand UO_2754 (O_2754,N_29506,N_29542);
nand UO_2755 (O_2755,N_29467,N_29984);
and UO_2756 (O_2756,N_29687,N_29397);
and UO_2757 (O_2757,N_29835,N_29720);
or UO_2758 (O_2758,N_29396,N_29073);
xor UO_2759 (O_2759,N_29775,N_29689);
nor UO_2760 (O_2760,N_29769,N_29138);
xor UO_2761 (O_2761,N_29015,N_29155);
or UO_2762 (O_2762,N_29499,N_29886);
and UO_2763 (O_2763,N_29315,N_29209);
nand UO_2764 (O_2764,N_29166,N_29409);
or UO_2765 (O_2765,N_29656,N_29358);
xnor UO_2766 (O_2766,N_29877,N_29860);
xnor UO_2767 (O_2767,N_29111,N_29724);
and UO_2768 (O_2768,N_29946,N_29521);
xor UO_2769 (O_2769,N_29767,N_29026);
nand UO_2770 (O_2770,N_29403,N_29822);
and UO_2771 (O_2771,N_29272,N_29585);
and UO_2772 (O_2772,N_29564,N_29295);
or UO_2773 (O_2773,N_29333,N_29505);
xnor UO_2774 (O_2774,N_29070,N_29502);
or UO_2775 (O_2775,N_29840,N_29462);
nor UO_2776 (O_2776,N_29344,N_29551);
nor UO_2777 (O_2777,N_29326,N_29263);
and UO_2778 (O_2778,N_29982,N_29674);
nor UO_2779 (O_2779,N_29668,N_29255);
and UO_2780 (O_2780,N_29723,N_29129);
and UO_2781 (O_2781,N_29933,N_29676);
and UO_2782 (O_2782,N_29104,N_29080);
nand UO_2783 (O_2783,N_29280,N_29691);
nand UO_2784 (O_2784,N_29934,N_29819);
nor UO_2785 (O_2785,N_29705,N_29412);
and UO_2786 (O_2786,N_29706,N_29775);
and UO_2787 (O_2787,N_29889,N_29756);
nand UO_2788 (O_2788,N_29242,N_29505);
nor UO_2789 (O_2789,N_29818,N_29920);
xor UO_2790 (O_2790,N_29307,N_29853);
nand UO_2791 (O_2791,N_29614,N_29789);
and UO_2792 (O_2792,N_29371,N_29397);
and UO_2793 (O_2793,N_29130,N_29235);
or UO_2794 (O_2794,N_29009,N_29725);
xnor UO_2795 (O_2795,N_29171,N_29650);
and UO_2796 (O_2796,N_29682,N_29558);
nor UO_2797 (O_2797,N_29974,N_29269);
nor UO_2798 (O_2798,N_29847,N_29907);
xnor UO_2799 (O_2799,N_29218,N_29281);
nor UO_2800 (O_2800,N_29304,N_29439);
nor UO_2801 (O_2801,N_29100,N_29298);
xnor UO_2802 (O_2802,N_29381,N_29643);
nand UO_2803 (O_2803,N_29630,N_29223);
nor UO_2804 (O_2804,N_29638,N_29074);
nand UO_2805 (O_2805,N_29381,N_29584);
nor UO_2806 (O_2806,N_29012,N_29664);
or UO_2807 (O_2807,N_29999,N_29167);
or UO_2808 (O_2808,N_29498,N_29215);
or UO_2809 (O_2809,N_29372,N_29074);
or UO_2810 (O_2810,N_29425,N_29893);
and UO_2811 (O_2811,N_29953,N_29278);
and UO_2812 (O_2812,N_29426,N_29031);
and UO_2813 (O_2813,N_29440,N_29622);
or UO_2814 (O_2814,N_29632,N_29191);
and UO_2815 (O_2815,N_29153,N_29613);
nor UO_2816 (O_2816,N_29475,N_29190);
nand UO_2817 (O_2817,N_29034,N_29130);
or UO_2818 (O_2818,N_29238,N_29569);
xnor UO_2819 (O_2819,N_29853,N_29258);
or UO_2820 (O_2820,N_29083,N_29239);
or UO_2821 (O_2821,N_29054,N_29812);
or UO_2822 (O_2822,N_29774,N_29501);
nor UO_2823 (O_2823,N_29505,N_29500);
or UO_2824 (O_2824,N_29187,N_29505);
xnor UO_2825 (O_2825,N_29902,N_29504);
xor UO_2826 (O_2826,N_29224,N_29876);
nand UO_2827 (O_2827,N_29578,N_29136);
or UO_2828 (O_2828,N_29958,N_29669);
nand UO_2829 (O_2829,N_29664,N_29450);
or UO_2830 (O_2830,N_29802,N_29620);
nand UO_2831 (O_2831,N_29401,N_29983);
nand UO_2832 (O_2832,N_29617,N_29793);
nand UO_2833 (O_2833,N_29197,N_29974);
nand UO_2834 (O_2834,N_29870,N_29396);
nor UO_2835 (O_2835,N_29855,N_29499);
nand UO_2836 (O_2836,N_29935,N_29258);
xor UO_2837 (O_2837,N_29293,N_29840);
or UO_2838 (O_2838,N_29973,N_29253);
nor UO_2839 (O_2839,N_29663,N_29582);
and UO_2840 (O_2840,N_29603,N_29590);
or UO_2841 (O_2841,N_29433,N_29871);
or UO_2842 (O_2842,N_29208,N_29275);
nor UO_2843 (O_2843,N_29480,N_29409);
nor UO_2844 (O_2844,N_29572,N_29263);
or UO_2845 (O_2845,N_29955,N_29013);
nand UO_2846 (O_2846,N_29806,N_29667);
nand UO_2847 (O_2847,N_29542,N_29155);
or UO_2848 (O_2848,N_29411,N_29088);
nand UO_2849 (O_2849,N_29914,N_29539);
or UO_2850 (O_2850,N_29122,N_29545);
xnor UO_2851 (O_2851,N_29067,N_29306);
and UO_2852 (O_2852,N_29689,N_29971);
xnor UO_2853 (O_2853,N_29532,N_29656);
xor UO_2854 (O_2854,N_29536,N_29030);
or UO_2855 (O_2855,N_29296,N_29981);
xnor UO_2856 (O_2856,N_29178,N_29706);
xor UO_2857 (O_2857,N_29863,N_29210);
nor UO_2858 (O_2858,N_29238,N_29189);
and UO_2859 (O_2859,N_29552,N_29384);
or UO_2860 (O_2860,N_29899,N_29645);
nand UO_2861 (O_2861,N_29738,N_29035);
xnor UO_2862 (O_2862,N_29582,N_29067);
and UO_2863 (O_2863,N_29490,N_29866);
or UO_2864 (O_2864,N_29471,N_29603);
nand UO_2865 (O_2865,N_29470,N_29224);
and UO_2866 (O_2866,N_29962,N_29732);
nand UO_2867 (O_2867,N_29536,N_29994);
nor UO_2868 (O_2868,N_29013,N_29711);
or UO_2869 (O_2869,N_29101,N_29228);
and UO_2870 (O_2870,N_29222,N_29516);
and UO_2871 (O_2871,N_29809,N_29015);
or UO_2872 (O_2872,N_29024,N_29567);
xnor UO_2873 (O_2873,N_29233,N_29359);
nor UO_2874 (O_2874,N_29086,N_29242);
nand UO_2875 (O_2875,N_29052,N_29872);
and UO_2876 (O_2876,N_29766,N_29956);
nand UO_2877 (O_2877,N_29118,N_29650);
xor UO_2878 (O_2878,N_29991,N_29561);
nand UO_2879 (O_2879,N_29278,N_29062);
and UO_2880 (O_2880,N_29913,N_29996);
and UO_2881 (O_2881,N_29562,N_29856);
and UO_2882 (O_2882,N_29561,N_29017);
nand UO_2883 (O_2883,N_29611,N_29846);
and UO_2884 (O_2884,N_29363,N_29530);
or UO_2885 (O_2885,N_29173,N_29164);
xor UO_2886 (O_2886,N_29261,N_29318);
nor UO_2887 (O_2887,N_29117,N_29919);
xnor UO_2888 (O_2888,N_29701,N_29108);
nor UO_2889 (O_2889,N_29152,N_29712);
or UO_2890 (O_2890,N_29397,N_29205);
nand UO_2891 (O_2891,N_29351,N_29751);
nor UO_2892 (O_2892,N_29706,N_29001);
nand UO_2893 (O_2893,N_29725,N_29140);
nor UO_2894 (O_2894,N_29602,N_29864);
and UO_2895 (O_2895,N_29632,N_29461);
nor UO_2896 (O_2896,N_29319,N_29963);
and UO_2897 (O_2897,N_29529,N_29673);
and UO_2898 (O_2898,N_29116,N_29335);
nand UO_2899 (O_2899,N_29750,N_29898);
nand UO_2900 (O_2900,N_29017,N_29425);
and UO_2901 (O_2901,N_29953,N_29903);
nand UO_2902 (O_2902,N_29849,N_29775);
and UO_2903 (O_2903,N_29457,N_29765);
nor UO_2904 (O_2904,N_29854,N_29790);
or UO_2905 (O_2905,N_29766,N_29159);
and UO_2906 (O_2906,N_29118,N_29027);
or UO_2907 (O_2907,N_29022,N_29371);
or UO_2908 (O_2908,N_29192,N_29838);
nand UO_2909 (O_2909,N_29018,N_29940);
nor UO_2910 (O_2910,N_29333,N_29392);
nand UO_2911 (O_2911,N_29546,N_29983);
and UO_2912 (O_2912,N_29844,N_29029);
xnor UO_2913 (O_2913,N_29568,N_29503);
nand UO_2914 (O_2914,N_29308,N_29137);
and UO_2915 (O_2915,N_29807,N_29632);
xor UO_2916 (O_2916,N_29236,N_29966);
nor UO_2917 (O_2917,N_29219,N_29838);
or UO_2918 (O_2918,N_29850,N_29151);
xor UO_2919 (O_2919,N_29030,N_29018);
nand UO_2920 (O_2920,N_29413,N_29743);
xor UO_2921 (O_2921,N_29352,N_29614);
xor UO_2922 (O_2922,N_29018,N_29107);
nand UO_2923 (O_2923,N_29470,N_29336);
xnor UO_2924 (O_2924,N_29121,N_29335);
xor UO_2925 (O_2925,N_29693,N_29187);
nand UO_2926 (O_2926,N_29412,N_29286);
and UO_2927 (O_2927,N_29006,N_29208);
xnor UO_2928 (O_2928,N_29601,N_29640);
xnor UO_2929 (O_2929,N_29082,N_29532);
xor UO_2930 (O_2930,N_29827,N_29291);
xor UO_2931 (O_2931,N_29051,N_29362);
or UO_2932 (O_2932,N_29331,N_29888);
and UO_2933 (O_2933,N_29302,N_29906);
or UO_2934 (O_2934,N_29884,N_29914);
xor UO_2935 (O_2935,N_29707,N_29308);
xnor UO_2936 (O_2936,N_29585,N_29653);
and UO_2937 (O_2937,N_29122,N_29689);
nor UO_2938 (O_2938,N_29795,N_29886);
or UO_2939 (O_2939,N_29153,N_29238);
nor UO_2940 (O_2940,N_29005,N_29954);
or UO_2941 (O_2941,N_29155,N_29526);
and UO_2942 (O_2942,N_29083,N_29027);
nor UO_2943 (O_2943,N_29350,N_29131);
nand UO_2944 (O_2944,N_29279,N_29117);
or UO_2945 (O_2945,N_29909,N_29095);
nand UO_2946 (O_2946,N_29358,N_29311);
and UO_2947 (O_2947,N_29143,N_29484);
and UO_2948 (O_2948,N_29828,N_29914);
nor UO_2949 (O_2949,N_29150,N_29459);
xor UO_2950 (O_2950,N_29402,N_29369);
nand UO_2951 (O_2951,N_29638,N_29896);
xnor UO_2952 (O_2952,N_29912,N_29945);
and UO_2953 (O_2953,N_29189,N_29983);
and UO_2954 (O_2954,N_29680,N_29014);
or UO_2955 (O_2955,N_29345,N_29520);
and UO_2956 (O_2956,N_29933,N_29762);
or UO_2957 (O_2957,N_29959,N_29889);
xor UO_2958 (O_2958,N_29870,N_29112);
nand UO_2959 (O_2959,N_29025,N_29082);
and UO_2960 (O_2960,N_29210,N_29178);
or UO_2961 (O_2961,N_29868,N_29461);
or UO_2962 (O_2962,N_29126,N_29226);
xor UO_2963 (O_2963,N_29319,N_29846);
or UO_2964 (O_2964,N_29200,N_29040);
nand UO_2965 (O_2965,N_29506,N_29387);
nand UO_2966 (O_2966,N_29646,N_29377);
nand UO_2967 (O_2967,N_29136,N_29590);
xor UO_2968 (O_2968,N_29215,N_29004);
nand UO_2969 (O_2969,N_29208,N_29217);
nand UO_2970 (O_2970,N_29693,N_29936);
nor UO_2971 (O_2971,N_29293,N_29996);
xor UO_2972 (O_2972,N_29505,N_29185);
nor UO_2973 (O_2973,N_29665,N_29975);
and UO_2974 (O_2974,N_29249,N_29529);
nand UO_2975 (O_2975,N_29151,N_29237);
or UO_2976 (O_2976,N_29958,N_29637);
or UO_2977 (O_2977,N_29729,N_29160);
nor UO_2978 (O_2978,N_29515,N_29077);
or UO_2979 (O_2979,N_29885,N_29452);
xor UO_2980 (O_2980,N_29625,N_29512);
xor UO_2981 (O_2981,N_29051,N_29058);
and UO_2982 (O_2982,N_29597,N_29660);
and UO_2983 (O_2983,N_29888,N_29831);
and UO_2984 (O_2984,N_29563,N_29072);
xnor UO_2985 (O_2985,N_29664,N_29289);
nand UO_2986 (O_2986,N_29346,N_29910);
or UO_2987 (O_2987,N_29144,N_29445);
and UO_2988 (O_2988,N_29128,N_29942);
or UO_2989 (O_2989,N_29022,N_29248);
nor UO_2990 (O_2990,N_29790,N_29512);
and UO_2991 (O_2991,N_29757,N_29912);
and UO_2992 (O_2992,N_29572,N_29036);
or UO_2993 (O_2993,N_29885,N_29732);
nand UO_2994 (O_2994,N_29160,N_29772);
nand UO_2995 (O_2995,N_29233,N_29129);
xnor UO_2996 (O_2996,N_29201,N_29947);
and UO_2997 (O_2997,N_29616,N_29045);
nand UO_2998 (O_2998,N_29255,N_29266);
or UO_2999 (O_2999,N_29503,N_29119);
or UO_3000 (O_3000,N_29729,N_29870);
and UO_3001 (O_3001,N_29955,N_29920);
nor UO_3002 (O_3002,N_29143,N_29230);
or UO_3003 (O_3003,N_29623,N_29805);
or UO_3004 (O_3004,N_29361,N_29194);
and UO_3005 (O_3005,N_29406,N_29600);
nand UO_3006 (O_3006,N_29164,N_29612);
nand UO_3007 (O_3007,N_29222,N_29470);
xor UO_3008 (O_3008,N_29473,N_29091);
or UO_3009 (O_3009,N_29717,N_29226);
nand UO_3010 (O_3010,N_29997,N_29755);
or UO_3011 (O_3011,N_29930,N_29280);
or UO_3012 (O_3012,N_29159,N_29022);
xnor UO_3013 (O_3013,N_29011,N_29435);
nand UO_3014 (O_3014,N_29311,N_29049);
nand UO_3015 (O_3015,N_29297,N_29080);
nand UO_3016 (O_3016,N_29840,N_29589);
or UO_3017 (O_3017,N_29407,N_29450);
or UO_3018 (O_3018,N_29647,N_29548);
or UO_3019 (O_3019,N_29609,N_29853);
nor UO_3020 (O_3020,N_29655,N_29493);
nand UO_3021 (O_3021,N_29271,N_29465);
xnor UO_3022 (O_3022,N_29334,N_29795);
and UO_3023 (O_3023,N_29085,N_29873);
nor UO_3024 (O_3024,N_29108,N_29642);
or UO_3025 (O_3025,N_29927,N_29302);
xnor UO_3026 (O_3026,N_29862,N_29910);
nor UO_3027 (O_3027,N_29818,N_29212);
nor UO_3028 (O_3028,N_29074,N_29261);
xor UO_3029 (O_3029,N_29401,N_29977);
or UO_3030 (O_3030,N_29988,N_29505);
xor UO_3031 (O_3031,N_29748,N_29571);
and UO_3032 (O_3032,N_29984,N_29457);
nor UO_3033 (O_3033,N_29693,N_29922);
or UO_3034 (O_3034,N_29142,N_29359);
and UO_3035 (O_3035,N_29698,N_29386);
nand UO_3036 (O_3036,N_29993,N_29355);
xnor UO_3037 (O_3037,N_29324,N_29289);
or UO_3038 (O_3038,N_29099,N_29367);
nand UO_3039 (O_3039,N_29618,N_29084);
xor UO_3040 (O_3040,N_29727,N_29705);
nand UO_3041 (O_3041,N_29674,N_29532);
and UO_3042 (O_3042,N_29533,N_29458);
nor UO_3043 (O_3043,N_29886,N_29398);
or UO_3044 (O_3044,N_29848,N_29058);
nor UO_3045 (O_3045,N_29706,N_29500);
or UO_3046 (O_3046,N_29933,N_29414);
xor UO_3047 (O_3047,N_29737,N_29374);
xor UO_3048 (O_3048,N_29408,N_29227);
or UO_3049 (O_3049,N_29869,N_29032);
or UO_3050 (O_3050,N_29690,N_29981);
nand UO_3051 (O_3051,N_29334,N_29012);
or UO_3052 (O_3052,N_29742,N_29775);
nor UO_3053 (O_3053,N_29526,N_29401);
nand UO_3054 (O_3054,N_29674,N_29319);
xnor UO_3055 (O_3055,N_29293,N_29417);
xor UO_3056 (O_3056,N_29982,N_29791);
and UO_3057 (O_3057,N_29107,N_29298);
nand UO_3058 (O_3058,N_29471,N_29497);
and UO_3059 (O_3059,N_29333,N_29179);
nand UO_3060 (O_3060,N_29376,N_29008);
nor UO_3061 (O_3061,N_29460,N_29762);
nand UO_3062 (O_3062,N_29844,N_29445);
nor UO_3063 (O_3063,N_29672,N_29325);
xor UO_3064 (O_3064,N_29615,N_29953);
xor UO_3065 (O_3065,N_29339,N_29709);
nand UO_3066 (O_3066,N_29259,N_29912);
nand UO_3067 (O_3067,N_29693,N_29962);
xnor UO_3068 (O_3068,N_29470,N_29630);
and UO_3069 (O_3069,N_29222,N_29725);
nor UO_3070 (O_3070,N_29199,N_29742);
nand UO_3071 (O_3071,N_29003,N_29325);
nor UO_3072 (O_3072,N_29298,N_29752);
nor UO_3073 (O_3073,N_29365,N_29170);
xor UO_3074 (O_3074,N_29171,N_29348);
nor UO_3075 (O_3075,N_29606,N_29135);
nor UO_3076 (O_3076,N_29153,N_29513);
and UO_3077 (O_3077,N_29805,N_29524);
and UO_3078 (O_3078,N_29753,N_29725);
nor UO_3079 (O_3079,N_29630,N_29393);
or UO_3080 (O_3080,N_29882,N_29963);
nor UO_3081 (O_3081,N_29168,N_29676);
nand UO_3082 (O_3082,N_29750,N_29145);
or UO_3083 (O_3083,N_29465,N_29708);
nor UO_3084 (O_3084,N_29059,N_29629);
nor UO_3085 (O_3085,N_29046,N_29590);
nor UO_3086 (O_3086,N_29631,N_29997);
or UO_3087 (O_3087,N_29971,N_29911);
xnor UO_3088 (O_3088,N_29924,N_29488);
nor UO_3089 (O_3089,N_29280,N_29067);
nand UO_3090 (O_3090,N_29393,N_29938);
nor UO_3091 (O_3091,N_29227,N_29493);
xnor UO_3092 (O_3092,N_29755,N_29989);
xor UO_3093 (O_3093,N_29821,N_29653);
nand UO_3094 (O_3094,N_29726,N_29970);
or UO_3095 (O_3095,N_29416,N_29079);
xnor UO_3096 (O_3096,N_29720,N_29246);
and UO_3097 (O_3097,N_29883,N_29483);
nand UO_3098 (O_3098,N_29426,N_29628);
or UO_3099 (O_3099,N_29748,N_29045);
nor UO_3100 (O_3100,N_29014,N_29718);
and UO_3101 (O_3101,N_29707,N_29387);
or UO_3102 (O_3102,N_29819,N_29809);
xor UO_3103 (O_3103,N_29612,N_29129);
or UO_3104 (O_3104,N_29315,N_29342);
or UO_3105 (O_3105,N_29308,N_29841);
xnor UO_3106 (O_3106,N_29379,N_29818);
xnor UO_3107 (O_3107,N_29246,N_29281);
and UO_3108 (O_3108,N_29778,N_29561);
xnor UO_3109 (O_3109,N_29595,N_29492);
and UO_3110 (O_3110,N_29250,N_29693);
nand UO_3111 (O_3111,N_29284,N_29125);
xnor UO_3112 (O_3112,N_29859,N_29099);
or UO_3113 (O_3113,N_29879,N_29245);
and UO_3114 (O_3114,N_29303,N_29865);
nand UO_3115 (O_3115,N_29023,N_29758);
or UO_3116 (O_3116,N_29647,N_29505);
and UO_3117 (O_3117,N_29878,N_29252);
and UO_3118 (O_3118,N_29511,N_29344);
and UO_3119 (O_3119,N_29083,N_29261);
nand UO_3120 (O_3120,N_29433,N_29385);
xor UO_3121 (O_3121,N_29995,N_29971);
and UO_3122 (O_3122,N_29266,N_29748);
and UO_3123 (O_3123,N_29904,N_29224);
nor UO_3124 (O_3124,N_29473,N_29382);
nand UO_3125 (O_3125,N_29398,N_29056);
or UO_3126 (O_3126,N_29913,N_29195);
nand UO_3127 (O_3127,N_29737,N_29901);
nor UO_3128 (O_3128,N_29340,N_29954);
and UO_3129 (O_3129,N_29785,N_29689);
xor UO_3130 (O_3130,N_29130,N_29635);
nand UO_3131 (O_3131,N_29970,N_29883);
and UO_3132 (O_3132,N_29938,N_29001);
nand UO_3133 (O_3133,N_29407,N_29260);
or UO_3134 (O_3134,N_29688,N_29034);
nor UO_3135 (O_3135,N_29023,N_29039);
and UO_3136 (O_3136,N_29297,N_29812);
xnor UO_3137 (O_3137,N_29773,N_29152);
nand UO_3138 (O_3138,N_29722,N_29571);
or UO_3139 (O_3139,N_29492,N_29344);
and UO_3140 (O_3140,N_29904,N_29110);
and UO_3141 (O_3141,N_29896,N_29318);
and UO_3142 (O_3142,N_29592,N_29814);
xor UO_3143 (O_3143,N_29951,N_29037);
xnor UO_3144 (O_3144,N_29282,N_29018);
or UO_3145 (O_3145,N_29655,N_29136);
nand UO_3146 (O_3146,N_29579,N_29609);
xor UO_3147 (O_3147,N_29270,N_29174);
nor UO_3148 (O_3148,N_29752,N_29682);
xor UO_3149 (O_3149,N_29352,N_29818);
or UO_3150 (O_3150,N_29287,N_29562);
and UO_3151 (O_3151,N_29906,N_29019);
and UO_3152 (O_3152,N_29871,N_29164);
nor UO_3153 (O_3153,N_29978,N_29595);
nor UO_3154 (O_3154,N_29850,N_29327);
and UO_3155 (O_3155,N_29416,N_29339);
nor UO_3156 (O_3156,N_29864,N_29274);
nor UO_3157 (O_3157,N_29248,N_29057);
and UO_3158 (O_3158,N_29632,N_29280);
and UO_3159 (O_3159,N_29687,N_29388);
and UO_3160 (O_3160,N_29106,N_29147);
and UO_3161 (O_3161,N_29993,N_29525);
and UO_3162 (O_3162,N_29442,N_29917);
or UO_3163 (O_3163,N_29730,N_29265);
nor UO_3164 (O_3164,N_29466,N_29484);
and UO_3165 (O_3165,N_29414,N_29021);
and UO_3166 (O_3166,N_29511,N_29144);
xor UO_3167 (O_3167,N_29801,N_29372);
xnor UO_3168 (O_3168,N_29374,N_29138);
xor UO_3169 (O_3169,N_29122,N_29527);
xor UO_3170 (O_3170,N_29345,N_29719);
or UO_3171 (O_3171,N_29817,N_29235);
and UO_3172 (O_3172,N_29541,N_29891);
xnor UO_3173 (O_3173,N_29832,N_29701);
and UO_3174 (O_3174,N_29338,N_29465);
nor UO_3175 (O_3175,N_29107,N_29579);
nor UO_3176 (O_3176,N_29733,N_29442);
nand UO_3177 (O_3177,N_29869,N_29054);
xor UO_3178 (O_3178,N_29426,N_29154);
or UO_3179 (O_3179,N_29230,N_29964);
or UO_3180 (O_3180,N_29268,N_29821);
or UO_3181 (O_3181,N_29500,N_29234);
nor UO_3182 (O_3182,N_29425,N_29862);
xnor UO_3183 (O_3183,N_29960,N_29976);
xnor UO_3184 (O_3184,N_29208,N_29683);
or UO_3185 (O_3185,N_29560,N_29672);
or UO_3186 (O_3186,N_29228,N_29931);
xnor UO_3187 (O_3187,N_29571,N_29919);
and UO_3188 (O_3188,N_29991,N_29318);
nor UO_3189 (O_3189,N_29577,N_29425);
nor UO_3190 (O_3190,N_29574,N_29348);
or UO_3191 (O_3191,N_29186,N_29832);
xor UO_3192 (O_3192,N_29903,N_29281);
nand UO_3193 (O_3193,N_29012,N_29197);
nor UO_3194 (O_3194,N_29873,N_29933);
xnor UO_3195 (O_3195,N_29887,N_29967);
nor UO_3196 (O_3196,N_29190,N_29973);
xnor UO_3197 (O_3197,N_29609,N_29289);
nand UO_3198 (O_3198,N_29625,N_29806);
xnor UO_3199 (O_3199,N_29220,N_29158);
or UO_3200 (O_3200,N_29471,N_29454);
nand UO_3201 (O_3201,N_29389,N_29575);
xor UO_3202 (O_3202,N_29488,N_29584);
or UO_3203 (O_3203,N_29440,N_29262);
and UO_3204 (O_3204,N_29269,N_29590);
and UO_3205 (O_3205,N_29459,N_29602);
xor UO_3206 (O_3206,N_29776,N_29866);
nor UO_3207 (O_3207,N_29854,N_29690);
and UO_3208 (O_3208,N_29895,N_29525);
nor UO_3209 (O_3209,N_29973,N_29760);
nor UO_3210 (O_3210,N_29251,N_29523);
nor UO_3211 (O_3211,N_29554,N_29026);
nand UO_3212 (O_3212,N_29665,N_29758);
xnor UO_3213 (O_3213,N_29576,N_29312);
xnor UO_3214 (O_3214,N_29067,N_29093);
xor UO_3215 (O_3215,N_29201,N_29840);
or UO_3216 (O_3216,N_29972,N_29251);
nand UO_3217 (O_3217,N_29123,N_29472);
and UO_3218 (O_3218,N_29821,N_29538);
nor UO_3219 (O_3219,N_29152,N_29035);
xor UO_3220 (O_3220,N_29485,N_29062);
or UO_3221 (O_3221,N_29640,N_29939);
nor UO_3222 (O_3222,N_29476,N_29419);
or UO_3223 (O_3223,N_29892,N_29147);
nor UO_3224 (O_3224,N_29472,N_29344);
xnor UO_3225 (O_3225,N_29576,N_29413);
nor UO_3226 (O_3226,N_29074,N_29954);
nand UO_3227 (O_3227,N_29174,N_29056);
or UO_3228 (O_3228,N_29211,N_29446);
or UO_3229 (O_3229,N_29573,N_29235);
nand UO_3230 (O_3230,N_29882,N_29647);
or UO_3231 (O_3231,N_29690,N_29883);
and UO_3232 (O_3232,N_29633,N_29583);
xnor UO_3233 (O_3233,N_29757,N_29669);
nor UO_3234 (O_3234,N_29986,N_29842);
xnor UO_3235 (O_3235,N_29017,N_29939);
and UO_3236 (O_3236,N_29358,N_29365);
and UO_3237 (O_3237,N_29149,N_29562);
xor UO_3238 (O_3238,N_29151,N_29210);
nand UO_3239 (O_3239,N_29354,N_29668);
and UO_3240 (O_3240,N_29652,N_29904);
and UO_3241 (O_3241,N_29919,N_29943);
nor UO_3242 (O_3242,N_29610,N_29674);
or UO_3243 (O_3243,N_29656,N_29109);
xor UO_3244 (O_3244,N_29116,N_29317);
nand UO_3245 (O_3245,N_29962,N_29724);
or UO_3246 (O_3246,N_29689,N_29600);
or UO_3247 (O_3247,N_29392,N_29901);
nand UO_3248 (O_3248,N_29946,N_29848);
or UO_3249 (O_3249,N_29185,N_29610);
nor UO_3250 (O_3250,N_29936,N_29295);
and UO_3251 (O_3251,N_29034,N_29945);
xor UO_3252 (O_3252,N_29439,N_29347);
xnor UO_3253 (O_3253,N_29234,N_29594);
and UO_3254 (O_3254,N_29625,N_29244);
and UO_3255 (O_3255,N_29015,N_29643);
xnor UO_3256 (O_3256,N_29042,N_29810);
xor UO_3257 (O_3257,N_29478,N_29055);
or UO_3258 (O_3258,N_29019,N_29966);
and UO_3259 (O_3259,N_29841,N_29189);
nor UO_3260 (O_3260,N_29676,N_29847);
nor UO_3261 (O_3261,N_29100,N_29504);
nor UO_3262 (O_3262,N_29999,N_29072);
xor UO_3263 (O_3263,N_29464,N_29013);
nand UO_3264 (O_3264,N_29489,N_29531);
nand UO_3265 (O_3265,N_29877,N_29140);
xor UO_3266 (O_3266,N_29328,N_29584);
and UO_3267 (O_3267,N_29901,N_29066);
and UO_3268 (O_3268,N_29530,N_29677);
or UO_3269 (O_3269,N_29321,N_29739);
xor UO_3270 (O_3270,N_29799,N_29256);
nor UO_3271 (O_3271,N_29578,N_29837);
xor UO_3272 (O_3272,N_29415,N_29863);
or UO_3273 (O_3273,N_29999,N_29926);
or UO_3274 (O_3274,N_29197,N_29670);
nand UO_3275 (O_3275,N_29602,N_29372);
and UO_3276 (O_3276,N_29130,N_29733);
and UO_3277 (O_3277,N_29671,N_29970);
nand UO_3278 (O_3278,N_29338,N_29726);
and UO_3279 (O_3279,N_29704,N_29308);
and UO_3280 (O_3280,N_29100,N_29983);
nand UO_3281 (O_3281,N_29970,N_29470);
xnor UO_3282 (O_3282,N_29898,N_29438);
nand UO_3283 (O_3283,N_29129,N_29001);
nor UO_3284 (O_3284,N_29858,N_29156);
nor UO_3285 (O_3285,N_29344,N_29497);
nor UO_3286 (O_3286,N_29726,N_29447);
and UO_3287 (O_3287,N_29210,N_29844);
and UO_3288 (O_3288,N_29716,N_29201);
or UO_3289 (O_3289,N_29384,N_29263);
xor UO_3290 (O_3290,N_29307,N_29535);
nand UO_3291 (O_3291,N_29806,N_29819);
nor UO_3292 (O_3292,N_29156,N_29706);
nand UO_3293 (O_3293,N_29598,N_29130);
or UO_3294 (O_3294,N_29646,N_29514);
nand UO_3295 (O_3295,N_29403,N_29067);
or UO_3296 (O_3296,N_29729,N_29660);
xor UO_3297 (O_3297,N_29132,N_29886);
and UO_3298 (O_3298,N_29186,N_29360);
nor UO_3299 (O_3299,N_29431,N_29578);
nor UO_3300 (O_3300,N_29358,N_29184);
xnor UO_3301 (O_3301,N_29526,N_29841);
and UO_3302 (O_3302,N_29803,N_29485);
nand UO_3303 (O_3303,N_29348,N_29157);
or UO_3304 (O_3304,N_29682,N_29400);
and UO_3305 (O_3305,N_29362,N_29616);
nor UO_3306 (O_3306,N_29689,N_29841);
and UO_3307 (O_3307,N_29074,N_29618);
and UO_3308 (O_3308,N_29122,N_29053);
and UO_3309 (O_3309,N_29711,N_29857);
xor UO_3310 (O_3310,N_29617,N_29339);
or UO_3311 (O_3311,N_29611,N_29472);
nor UO_3312 (O_3312,N_29318,N_29590);
xnor UO_3313 (O_3313,N_29718,N_29217);
nand UO_3314 (O_3314,N_29511,N_29198);
and UO_3315 (O_3315,N_29486,N_29398);
nor UO_3316 (O_3316,N_29713,N_29681);
nor UO_3317 (O_3317,N_29319,N_29186);
or UO_3318 (O_3318,N_29120,N_29737);
xor UO_3319 (O_3319,N_29274,N_29132);
and UO_3320 (O_3320,N_29529,N_29811);
or UO_3321 (O_3321,N_29321,N_29331);
or UO_3322 (O_3322,N_29321,N_29959);
and UO_3323 (O_3323,N_29136,N_29031);
and UO_3324 (O_3324,N_29741,N_29207);
or UO_3325 (O_3325,N_29113,N_29670);
nand UO_3326 (O_3326,N_29198,N_29762);
nor UO_3327 (O_3327,N_29346,N_29478);
xor UO_3328 (O_3328,N_29133,N_29004);
xnor UO_3329 (O_3329,N_29523,N_29507);
nand UO_3330 (O_3330,N_29413,N_29766);
or UO_3331 (O_3331,N_29411,N_29626);
nor UO_3332 (O_3332,N_29023,N_29211);
nor UO_3333 (O_3333,N_29043,N_29070);
nand UO_3334 (O_3334,N_29927,N_29414);
and UO_3335 (O_3335,N_29634,N_29980);
nand UO_3336 (O_3336,N_29242,N_29749);
or UO_3337 (O_3337,N_29448,N_29641);
nor UO_3338 (O_3338,N_29653,N_29682);
nor UO_3339 (O_3339,N_29985,N_29221);
nand UO_3340 (O_3340,N_29385,N_29983);
nand UO_3341 (O_3341,N_29946,N_29755);
nor UO_3342 (O_3342,N_29311,N_29101);
and UO_3343 (O_3343,N_29919,N_29346);
or UO_3344 (O_3344,N_29262,N_29349);
and UO_3345 (O_3345,N_29469,N_29648);
nor UO_3346 (O_3346,N_29562,N_29777);
xor UO_3347 (O_3347,N_29934,N_29414);
and UO_3348 (O_3348,N_29044,N_29621);
xor UO_3349 (O_3349,N_29893,N_29653);
or UO_3350 (O_3350,N_29801,N_29243);
and UO_3351 (O_3351,N_29553,N_29085);
and UO_3352 (O_3352,N_29678,N_29021);
nor UO_3353 (O_3353,N_29451,N_29181);
nor UO_3354 (O_3354,N_29740,N_29222);
nand UO_3355 (O_3355,N_29177,N_29684);
nor UO_3356 (O_3356,N_29591,N_29413);
nor UO_3357 (O_3357,N_29695,N_29810);
or UO_3358 (O_3358,N_29046,N_29111);
nor UO_3359 (O_3359,N_29434,N_29563);
nand UO_3360 (O_3360,N_29558,N_29296);
xor UO_3361 (O_3361,N_29287,N_29659);
and UO_3362 (O_3362,N_29439,N_29595);
and UO_3363 (O_3363,N_29173,N_29311);
and UO_3364 (O_3364,N_29588,N_29764);
and UO_3365 (O_3365,N_29313,N_29524);
xnor UO_3366 (O_3366,N_29414,N_29025);
or UO_3367 (O_3367,N_29869,N_29640);
nand UO_3368 (O_3368,N_29201,N_29170);
or UO_3369 (O_3369,N_29542,N_29135);
xnor UO_3370 (O_3370,N_29164,N_29039);
and UO_3371 (O_3371,N_29586,N_29270);
nor UO_3372 (O_3372,N_29298,N_29502);
nor UO_3373 (O_3373,N_29126,N_29091);
nor UO_3374 (O_3374,N_29823,N_29083);
or UO_3375 (O_3375,N_29828,N_29072);
xor UO_3376 (O_3376,N_29319,N_29666);
and UO_3377 (O_3377,N_29123,N_29637);
or UO_3378 (O_3378,N_29616,N_29387);
nor UO_3379 (O_3379,N_29413,N_29688);
and UO_3380 (O_3380,N_29549,N_29729);
nor UO_3381 (O_3381,N_29748,N_29034);
nor UO_3382 (O_3382,N_29293,N_29141);
xnor UO_3383 (O_3383,N_29275,N_29286);
xnor UO_3384 (O_3384,N_29492,N_29043);
and UO_3385 (O_3385,N_29321,N_29327);
and UO_3386 (O_3386,N_29500,N_29947);
nand UO_3387 (O_3387,N_29732,N_29468);
xnor UO_3388 (O_3388,N_29166,N_29485);
nor UO_3389 (O_3389,N_29473,N_29846);
nor UO_3390 (O_3390,N_29228,N_29564);
or UO_3391 (O_3391,N_29593,N_29642);
and UO_3392 (O_3392,N_29068,N_29741);
xnor UO_3393 (O_3393,N_29486,N_29634);
or UO_3394 (O_3394,N_29610,N_29096);
nand UO_3395 (O_3395,N_29377,N_29953);
nand UO_3396 (O_3396,N_29630,N_29997);
nor UO_3397 (O_3397,N_29906,N_29778);
and UO_3398 (O_3398,N_29689,N_29614);
and UO_3399 (O_3399,N_29034,N_29469);
xor UO_3400 (O_3400,N_29071,N_29051);
nor UO_3401 (O_3401,N_29439,N_29363);
and UO_3402 (O_3402,N_29679,N_29853);
and UO_3403 (O_3403,N_29906,N_29369);
or UO_3404 (O_3404,N_29438,N_29957);
xor UO_3405 (O_3405,N_29949,N_29864);
xnor UO_3406 (O_3406,N_29438,N_29890);
nor UO_3407 (O_3407,N_29312,N_29468);
nand UO_3408 (O_3408,N_29081,N_29078);
nand UO_3409 (O_3409,N_29899,N_29090);
or UO_3410 (O_3410,N_29933,N_29705);
nand UO_3411 (O_3411,N_29706,N_29647);
xor UO_3412 (O_3412,N_29871,N_29190);
xnor UO_3413 (O_3413,N_29965,N_29159);
or UO_3414 (O_3414,N_29117,N_29921);
nor UO_3415 (O_3415,N_29445,N_29619);
xnor UO_3416 (O_3416,N_29382,N_29617);
xnor UO_3417 (O_3417,N_29184,N_29235);
xnor UO_3418 (O_3418,N_29032,N_29369);
nand UO_3419 (O_3419,N_29185,N_29826);
nand UO_3420 (O_3420,N_29785,N_29951);
and UO_3421 (O_3421,N_29167,N_29100);
nand UO_3422 (O_3422,N_29869,N_29146);
xnor UO_3423 (O_3423,N_29839,N_29291);
nor UO_3424 (O_3424,N_29997,N_29350);
nor UO_3425 (O_3425,N_29759,N_29074);
and UO_3426 (O_3426,N_29073,N_29545);
nand UO_3427 (O_3427,N_29301,N_29318);
or UO_3428 (O_3428,N_29901,N_29610);
xnor UO_3429 (O_3429,N_29374,N_29207);
or UO_3430 (O_3430,N_29014,N_29880);
xnor UO_3431 (O_3431,N_29015,N_29424);
xnor UO_3432 (O_3432,N_29722,N_29366);
or UO_3433 (O_3433,N_29095,N_29792);
and UO_3434 (O_3434,N_29823,N_29066);
xor UO_3435 (O_3435,N_29531,N_29267);
nor UO_3436 (O_3436,N_29339,N_29982);
nor UO_3437 (O_3437,N_29441,N_29260);
nor UO_3438 (O_3438,N_29215,N_29866);
and UO_3439 (O_3439,N_29037,N_29242);
nor UO_3440 (O_3440,N_29627,N_29199);
xor UO_3441 (O_3441,N_29771,N_29469);
or UO_3442 (O_3442,N_29573,N_29049);
nand UO_3443 (O_3443,N_29061,N_29895);
nor UO_3444 (O_3444,N_29078,N_29611);
nand UO_3445 (O_3445,N_29891,N_29720);
xnor UO_3446 (O_3446,N_29850,N_29989);
nand UO_3447 (O_3447,N_29564,N_29333);
nor UO_3448 (O_3448,N_29130,N_29157);
xnor UO_3449 (O_3449,N_29738,N_29142);
xnor UO_3450 (O_3450,N_29179,N_29508);
xnor UO_3451 (O_3451,N_29704,N_29898);
nand UO_3452 (O_3452,N_29756,N_29761);
or UO_3453 (O_3453,N_29459,N_29634);
or UO_3454 (O_3454,N_29560,N_29028);
nor UO_3455 (O_3455,N_29271,N_29687);
nor UO_3456 (O_3456,N_29960,N_29640);
nand UO_3457 (O_3457,N_29692,N_29013);
nand UO_3458 (O_3458,N_29028,N_29074);
nand UO_3459 (O_3459,N_29651,N_29280);
and UO_3460 (O_3460,N_29238,N_29605);
and UO_3461 (O_3461,N_29943,N_29410);
and UO_3462 (O_3462,N_29688,N_29344);
or UO_3463 (O_3463,N_29660,N_29663);
xnor UO_3464 (O_3464,N_29894,N_29030);
and UO_3465 (O_3465,N_29682,N_29892);
and UO_3466 (O_3466,N_29874,N_29555);
and UO_3467 (O_3467,N_29497,N_29976);
and UO_3468 (O_3468,N_29196,N_29175);
and UO_3469 (O_3469,N_29492,N_29302);
and UO_3470 (O_3470,N_29327,N_29351);
nand UO_3471 (O_3471,N_29550,N_29374);
and UO_3472 (O_3472,N_29639,N_29892);
xor UO_3473 (O_3473,N_29463,N_29158);
or UO_3474 (O_3474,N_29703,N_29156);
xnor UO_3475 (O_3475,N_29204,N_29533);
nor UO_3476 (O_3476,N_29226,N_29035);
nand UO_3477 (O_3477,N_29556,N_29888);
or UO_3478 (O_3478,N_29649,N_29111);
and UO_3479 (O_3479,N_29660,N_29375);
or UO_3480 (O_3480,N_29217,N_29416);
or UO_3481 (O_3481,N_29265,N_29120);
and UO_3482 (O_3482,N_29180,N_29025);
nor UO_3483 (O_3483,N_29846,N_29895);
nor UO_3484 (O_3484,N_29716,N_29312);
nand UO_3485 (O_3485,N_29273,N_29852);
nor UO_3486 (O_3486,N_29386,N_29551);
and UO_3487 (O_3487,N_29786,N_29322);
and UO_3488 (O_3488,N_29670,N_29511);
nand UO_3489 (O_3489,N_29777,N_29475);
xor UO_3490 (O_3490,N_29760,N_29175);
or UO_3491 (O_3491,N_29351,N_29230);
or UO_3492 (O_3492,N_29789,N_29618);
nor UO_3493 (O_3493,N_29881,N_29691);
xor UO_3494 (O_3494,N_29858,N_29562);
nand UO_3495 (O_3495,N_29170,N_29635);
xnor UO_3496 (O_3496,N_29225,N_29257);
nor UO_3497 (O_3497,N_29734,N_29295);
nand UO_3498 (O_3498,N_29729,N_29987);
xor UO_3499 (O_3499,N_29246,N_29694);
endmodule