module basic_2500_25000_3000_40_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1352,In_2193);
xor U1 (N_1,In_1053,In_1748);
nand U2 (N_2,In_272,In_2315);
nor U3 (N_3,In_742,In_679);
xnor U4 (N_4,In_2441,In_897);
xnor U5 (N_5,In_2322,In_2395);
and U6 (N_6,In_806,In_759);
or U7 (N_7,In_1735,In_732);
nand U8 (N_8,In_1091,In_106);
xor U9 (N_9,In_1027,In_517);
nor U10 (N_10,In_825,In_2396);
nand U11 (N_11,In_324,In_1775);
xor U12 (N_12,In_386,In_1719);
nand U13 (N_13,In_1797,In_75);
and U14 (N_14,In_2151,In_1988);
and U15 (N_15,In_677,In_2344);
xor U16 (N_16,In_1169,In_495);
nor U17 (N_17,In_133,In_1236);
and U18 (N_18,In_1534,In_1782);
and U19 (N_19,In_1394,In_208);
and U20 (N_20,In_181,In_746);
and U21 (N_21,In_1376,In_691);
nor U22 (N_22,In_2120,In_1133);
nor U23 (N_23,In_422,In_125);
xor U24 (N_24,In_493,In_20);
and U25 (N_25,In_156,In_2316);
and U26 (N_26,In_520,In_790);
nand U27 (N_27,In_1472,In_65);
and U28 (N_28,In_1300,In_2062);
or U29 (N_29,In_874,In_1229);
and U30 (N_30,In_49,In_882);
and U31 (N_31,In_1431,In_2083);
and U32 (N_32,In_1101,In_311);
xnor U33 (N_33,In_37,In_1622);
nand U34 (N_34,In_2004,In_1208);
nand U35 (N_35,In_484,In_1720);
and U36 (N_36,In_2483,In_1466);
nand U37 (N_37,In_1817,In_1018);
nand U38 (N_38,In_2058,In_417);
nand U39 (N_39,In_1390,In_2241);
nand U40 (N_40,In_1890,In_1827);
and U41 (N_41,In_953,In_1627);
or U42 (N_42,In_2370,In_301);
nor U43 (N_43,In_260,In_1752);
and U44 (N_44,In_1128,In_1665);
or U45 (N_45,In_604,In_54);
and U46 (N_46,In_1322,In_1517);
nand U47 (N_47,In_1326,In_1649);
nor U48 (N_48,In_722,In_1807);
or U49 (N_49,In_1971,In_2367);
nand U50 (N_50,In_590,In_1366);
nor U51 (N_51,In_2172,In_1951);
nor U52 (N_52,In_1370,In_881);
and U53 (N_53,In_2457,In_640);
nand U54 (N_54,In_680,In_1878);
or U55 (N_55,In_780,In_1621);
and U56 (N_56,In_2436,In_1082);
and U57 (N_57,In_264,In_1280);
or U58 (N_58,In_756,In_1793);
and U59 (N_59,In_999,In_1289);
or U60 (N_60,In_1253,In_250);
and U61 (N_61,In_623,In_2131);
nand U62 (N_62,In_2328,In_330);
xor U63 (N_63,In_1417,In_1154);
and U64 (N_64,In_2117,In_580);
nor U65 (N_65,In_326,In_700);
or U66 (N_66,In_1100,In_2497);
and U67 (N_67,In_589,In_1533);
nor U68 (N_68,In_2213,In_507);
or U69 (N_69,In_2017,In_1578);
nand U70 (N_70,In_455,In_1781);
or U71 (N_71,In_1997,In_1028);
nand U72 (N_72,In_136,In_636);
xnor U73 (N_73,In_1172,In_427);
or U74 (N_74,In_148,In_114);
xor U75 (N_75,In_2076,In_409);
nor U76 (N_76,In_1731,In_436);
and U77 (N_77,In_1338,In_1846);
and U78 (N_78,In_968,In_384);
nor U79 (N_79,In_2499,In_627);
or U80 (N_80,In_498,In_309);
or U81 (N_81,In_1362,In_73);
and U82 (N_82,In_1174,In_2188);
nand U83 (N_83,In_1774,In_1502);
nor U84 (N_84,In_1697,In_2036);
nand U85 (N_85,In_2332,In_434);
nor U86 (N_86,In_2493,In_1221);
nand U87 (N_87,In_929,In_739);
or U88 (N_88,In_1840,In_2192);
or U89 (N_89,In_41,In_2018);
xnor U90 (N_90,In_1007,In_421);
xnor U91 (N_91,In_1337,In_594);
and U92 (N_92,In_1479,In_1702);
or U93 (N_93,In_792,In_843);
xor U94 (N_94,In_2264,In_1302);
and U95 (N_95,In_773,In_1411);
nand U96 (N_96,In_1469,In_1666);
nand U97 (N_97,In_2429,In_2066);
nand U98 (N_98,In_1835,In_723);
nor U99 (N_99,In_62,In_147);
xnor U100 (N_100,In_1911,In_1150);
and U101 (N_101,In_703,In_2187);
xor U102 (N_102,In_903,In_1132);
and U103 (N_103,In_1332,In_1497);
nor U104 (N_104,In_522,In_204);
nor U105 (N_105,In_104,In_475);
and U106 (N_106,In_2158,In_474);
nand U107 (N_107,In_1647,In_1836);
nand U108 (N_108,In_849,In_2362);
xnor U109 (N_109,In_942,In_2383);
or U110 (N_110,In_1601,In_1989);
nor U111 (N_111,In_2425,In_2454);
and U112 (N_112,In_396,In_2046);
nand U113 (N_113,In_103,In_1565);
nand U114 (N_114,In_2140,In_2416);
or U115 (N_115,In_820,In_29);
and U116 (N_116,In_1684,In_1899);
xor U117 (N_117,In_2221,In_2051);
and U118 (N_118,In_331,In_738);
nor U119 (N_119,In_767,In_976);
and U120 (N_120,In_365,In_1645);
nor U121 (N_121,In_1372,In_998);
and U122 (N_122,In_1135,In_115);
or U123 (N_123,In_46,In_298);
and U124 (N_124,In_270,In_1328);
xnor U125 (N_125,In_1025,In_2252);
or U126 (N_126,In_1607,In_1616);
xnor U127 (N_127,In_1405,In_2024);
xnor U128 (N_128,In_277,In_1355);
xor U129 (N_129,In_225,In_1023);
and U130 (N_130,In_374,In_1889);
nor U131 (N_131,In_1718,In_2400);
xnor U132 (N_132,In_232,In_315);
and U133 (N_133,In_2167,In_1083);
and U134 (N_134,In_950,In_1375);
or U135 (N_135,In_2081,In_1151);
or U136 (N_136,In_320,In_2164);
nor U137 (N_137,In_1768,In_2444);
xnor U138 (N_138,In_128,In_1408);
xnor U139 (N_139,In_2271,In_1651);
and U140 (N_140,In_1130,In_1239);
and U141 (N_141,In_1194,In_634);
or U142 (N_142,In_647,In_951);
nor U143 (N_143,In_912,In_1558);
nand U144 (N_144,In_715,In_711);
or U145 (N_145,In_72,In_1822);
nor U146 (N_146,In_120,In_1808);
nor U147 (N_147,In_2157,In_76);
xor U148 (N_148,In_2054,In_1410);
nand U149 (N_149,In_2148,In_2078);
xnor U150 (N_150,In_1769,In_496);
nor U151 (N_151,In_823,In_1068);
or U152 (N_152,In_2126,In_2009);
and U153 (N_153,In_1036,In_302);
or U154 (N_154,In_1085,In_1316);
or U155 (N_155,In_1409,In_213);
and U156 (N_156,In_240,In_752);
and U157 (N_157,In_1104,In_2353);
or U158 (N_158,In_481,In_763);
xnor U159 (N_159,In_1490,In_2410);
nor U160 (N_160,In_2155,In_1734);
and U161 (N_161,In_2084,In_1032);
nand U162 (N_162,In_1143,In_380);
xor U163 (N_163,In_2190,In_1920);
nand U164 (N_164,In_1215,In_788);
nand U165 (N_165,In_1333,In_588);
nor U166 (N_166,In_398,In_2006);
or U167 (N_167,In_2308,In_1004);
or U168 (N_168,In_488,In_1311);
and U169 (N_169,In_1541,In_555);
or U170 (N_170,In_472,In_984);
xor U171 (N_171,In_2432,In_2053);
nand U172 (N_172,In_1804,In_90);
or U173 (N_173,In_459,In_757);
nor U174 (N_174,In_1166,In_373);
nor U175 (N_175,In_1430,In_1560);
and U176 (N_176,In_100,In_940);
xnor U177 (N_177,In_891,In_827);
nand U178 (N_178,In_1675,In_1015);
and U179 (N_179,In_195,In_871);
nor U180 (N_180,In_2237,In_359);
xnor U181 (N_181,In_1139,In_888);
nor U182 (N_182,In_2105,In_2266);
and U183 (N_183,In_219,In_1464);
nand U184 (N_184,In_2405,In_1599);
xor U185 (N_185,In_57,In_2008);
and U186 (N_186,In_1526,In_2250);
nand U187 (N_187,In_1219,In_1939);
nand U188 (N_188,In_2179,In_2375);
nand U189 (N_189,In_1245,In_1287);
nand U190 (N_190,In_568,In_2130);
and U191 (N_191,In_2235,In_1155);
nand U192 (N_192,In_1250,In_1973);
xnor U193 (N_193,In_1763,In_1033);
nand U194 (N_194,In_2364,In_675);
nor U195 (N_195,In_1325,In_2458);
nand U196 (N_196,In_1984,In_227);
nor U197 (N_197,In_836,In_753);
nand U198 (N_198,In_1255,In_971);
or U199 (N_199,In_1981,In_1914);
nand U200 (N_200,In_808,In_123);
xnor U201 (N_201,In_457,In_562);
xor U202 (N_202,In_1696,In_23);
nor U203 (N_203,In_1330,In_770);
nor U204 (N_204,In_2477,In_1639);
nand U205 (N_205,In_1866,In_813);
or U206 (N_206,In_447,In_1515);
or U207 (N_207,In_1286,In_1730);
xor U208 (N_208,In_1324,In_571);
xnor U209 (N_209,In_406,In_176);
and U210 (N_210,In_560,In_2207);
or U211 (N_211,In_1514,In_401);
nor U212 (N_212,In_1746,In_197);
and U213 (N_213,In_1237,In_138);
or U214 (N_214,In_1893,In_2225);
and U215 (N_215,In_173,In_719);
nand U216 (N_216,In_124,In_1365);
nand U217 (N_217,In_748,In_2323);
nand U218 (N_218,In_1611,In_467);
nand U219 (N_219,In_111,In_1373);
or U220 (N_220,In_2049,In_2013);
and U221 (N_221,In_2333,In_924);
or U222 (N_222,In_1264,In_913);
and U223 (N_223,In_1868,In_599);
xor U224 (N_224,In_280,In_1281);
or U225 (N_225,In_2015,In_686);
nand U226 (N_226,In_892,In_2034);
nor U227 (N_227,In_2166,In_2104);
nor U228 (N_228,In_1545,In_787);
nand U229 (N_229,In_2388,In_273);
nand U230 (N_230,In_433,In_1121);
xor U231 (N_231,In_2277,In_153);
nor U232 (N_232,In_852,In_109);
nor U233 (N_233,In_2480,In_2135);
and U234 (N_234,In_1788,In_2397);
and U235 (N_235,In_1432,In_291);
xor U236 (N_236,In_1970,In_596);
xnor U237 (N_237,In_1875,In_1379);
xor U238 (N_238,In_1240,In_2020);
nor U239 (N_239,In_1400,In_1642);
or U240 (N_240,In_1880,In_1771);
xor U241 (N_241,In_1640,In_316);
or U242 (N_242,In_2303,In_2371);
nand U243 (N_243,In_1934,In_658);
nor U244 (N_244,In_205,In_622);
and U245 (N_245,In_1953,In_980);
or U246 (N_246,In_1717,In_463);
or U247 (N_247,In_1576,In_1780);
nand U248 (N_248,In_1884,In_1223);
xnor U249 (N_249,In_2401,In_1757);
and U250 (N_250,In_947,In_2378);
nand U251 (N_251,In_1729,In_1709);
nand U252 (N_252,In_650,In_978);
and U253 (N_253,In_694,In_1905);
nand U254 (N_254,In_554,In_1940);
xor U255 (N_255,In_1672,In_941);
and U256 (N_256,In_2299,In_2334);
nor U257 (N_257,In_171,In_1636);
nor U258 (N_258,In_721,In_1873);
xor U259 (N_259,In_6,In_2111);
and U260 (N_260,In_1276,In_31);
and U261 (N_261,In_1026,In_271);
nor U262 (N_262,In_426,In_629);
nand U263 (N_263,In_314,In_1447);
nor U264 (N_264,In_439,In_412);
or U265 (N_265,In_657,In_2168);
or U266 (N_266,In_766,In_1423);
xnor U267 (N_267,In_206,In_403);
nor U268 (N_268,In_1246,In_2263);
and U269 (N_269,In_1820,In_2283);
nor U270 (N_270,In_350,In_2014);
nor U271 (N_271,In_126,In_1902);
nor U272 (N_272,In_2350,In_1163);
nor U273 (N_273,In_1575,In_118);
and U274 (N_274,In_829,In_909);
xnor U275 (N_275,In_253,In_2447);
or U276 (N_276,In_1648,In_1310);
nor U277 (N_277,In_900,In_784);
xor U278 (N_278,In_2339,In_1059);
or U279 (N_279,In_1402,In_1109);
xnor U280 (N_280,In_1529,In_51);
nor U281 (N_281,In_189,In_1535);
xor U282 (N_282,In_531,In_1420);
xor U283 (N_283,In_1364,In_333);
xor U284 (N_284,In_2185,In_1888);
nand U285 (N_285,In_2301,In_855);
and U286 (N_286,In_1441,In_1047);
xnor U287 (N_287,In_712,In_2481);
xnor U288 (N_288,In_1187,In_2318);
and U289 (N_289,In_696,In_2340);
or U290 (N_290,In_239,In_1499);
xnor U291 (N_291,In_12,In_1921);
nand U292 (N_292,In_1094,In_1368);
nor U293 (N_293,In_2124,In_2482);
or U294 (N_294,In_229,In_966);
and U295 (N_295,In_2214,In_2421);
nor U296 (N_296,In_774,In_95);
or U297 (N_297,In_2202,In_2109);
nand U298 (N_298,In_2199,In_1153);
nor U299 (N_299,In_2035,In_2132);
or U300 (N_300,In_2331,In_297);
or U301 (N_301,In_1975,In_1103);
nor U302 (N_302,In_1102,In_987);
nor U303 (N_303,In_973,In_856);
nand U304 (N_304,In_193,In_1791);
nor U305 (N_305,In_1284,In_144);
or U306 (N_306,In_1290,In_2305);
nand U307 (N_307,In_294,In_1738);
nand U308 (N_308,In_1643,In_1900);
nor U309 (N_309,In_1474,In_1256);
xnor U310 (N_310,In_2108,In_247);
or U311 (N_311,In_117,In_1061);
or U312 (N_312,In_1307,In_538);
nor U313 (N_313,In_1380,In_342);
and U314 (N_314,In_948,In_1713);
nor U315 (N_315,In_2141,In_473);
and U316 (N_316,In_2442,In_2260);
or U317 (N_317,In_527,In_269);
and U318 (N_318,In_1670,In_710);
xor U319 (N_319,In_1896,In_1353);
or U320 (N_320,In_1839,In_1937);
xor U321 (N_321,In_2094,In_1413);
or U322 (N_322,In_2244,In_1983);
nor U323 (N_323,In_1871,In_915);
and U324 (N_324,In_744,In_1354);
and U325 (N_325,In_2359,In_1870);
nand U326 (N_326,In_2259,In_857);
nor U327 (N_327,In_949,In_186);
nor U328 (N_328,In_376,In_1434);
and U329 (N_329,In_754,In_1632);
or U330 (N_330,In_1120,In_551);
xnor U331 (N_331,In_553,In_2440);
or U332 (N_332,In_2142,In_83);
xor U333 (N_333,In_1573,In_2476);
nand U334 (N_334,In_656,In_1152);
nor U335 (N_335,In_1475,In_284);
and U336 (N_336,In_513,In_1570);
xor U337 (N_337,In_2437,In_1220);
xnor U338 (N_338,In_378,In_477);
nor U339 (N_339,In_2492,In_509);
xnor U340 (N_340,In_1553,In_167);
nor U341 (N_341,In_2282,In_28);
nand U342 (N_342,In_1021,In_1996);
or U343 (N_343,In_1987,In_1844);
nor U344 (N_344,In_2327,In_918);
or U345 (N_345,In_1427,In_441);
xnor U346 (N_346,In_772,In_163);
or U347 (N_347,In_1743,In_2460);
and U348 (N_348,In_1539,In_875);
or U349 (N_349,In_1903,In_340);
xnor U350 (N_350,In_556,In_1218);
or U351 (N_351,In_1357,In_1660);
nand U352 (N_352,In_2281,In_2267);
nor U353 (N_353,In_1389,In_2195);
and U354 (N_354,In_85,In_1667);
and U355 (N_355,In_783,In_2240);
nand U356 (N_356,In_745,In_851);
nand U357 (N_357,In_521,In_955);
and U358 (N_358,In_2358,In_500);
or U359 (N_359,In_1603,In_653);
nor U360 (N_360,In_1242,In_1954);
nor U361 (N_361,In_1606,In_448);
nor U362 (N_362,In_1504,In_1279);
or U363 (N_363,In_648,In_1048);
xor U364 (N_364,In_1227,In_2293);
nor U365 (N_365,In_2402,In_826);
nor U366 (N_366,In_2077,In_428);
and U367 (N_367,In_1478,In_1727);
nand U368 (N_368,In_1961,In_1428);
or U369 (N_369,In_285,In_2038);
or U370 (N_370,In_946,In_1456);
xnor U371 (N_371,In_1489,In_322);
xnor U372 (N_372,In_1600,In_1313);
nand U373 (N_373,In_1964,In_867);
xnor U374 (N_374,In_885,In_39);
and U375 (N_375,In_737,In_1561);
or U376 (N_376,In_61,In_685);
nand U377 (N_377,In_1841,In_524);
nand U378 (N_378,In_352,In_997);
xor U379 (N_379,In_2204,In_209);
nand U380 (N_380,In_1777,In_1929);
xnor U381 (N_381,In_353,In_740);
nor U382 (N_382,In_275,In_765);
or U383 (N_383,In_47,In_2251);
nor U384 (N_384,In_642,In_56);
xor U385 (N_385,In_2335,In_2230);
or U386 (N_386,In_2438,In_923);
nand U387 (N_387,In_246,In_2205);
xor U388 (N_388,In_50,In_9);
nand U389 (N_389,In_681,In_2183);
nor U390 (N_390,In_1708,In_778);
nand U391 (N_391,In_1142,In_1060);
nand U392 (N_392,In_1892,In_1234);
nor U393 (N_393,In_2298,In_1525);
or U394 (N_394,In_1031,In_2426);
nand U395 (N_395,In_442,In_425);
nor U396 (N_396,In_55,In_1909);
nand U397 (N_397,In_1105,In_1522);
or U398 (N_398,In_505,In_1378);
and U399 (N_399,In_1831,In_2466);
nand U400 (N_400,In_1090,In_728);
nor U401 (N_401,In_1704,In_1095);
and U402 (N_402,In_1002,In_1010);
nor U403 (N_403,In_1876,In_2433);
nor U404 (N_404,In_1823,In_497);
and U405 (N_405,In_768,In_1308);
xor U406 (N_406,In_1055,In_1495);
nor U407 (N_407,In_1853,In_802);
nor U408 (N_408,In_2103,In_336);
or U409 (N_409,In_979,In_981);
nand U410 (N_410,In_637,In_2178);
nor U411 (N_411,In_318,In_2469);
and U412 (N_412,In_1331,In_2355);
or U413 (N_413,In_190,In_431);
nand U414 (N_414,In_231,In_1124);
xnor U415 (N_415,In_2491,In_2464);
or U416 (N_416,In_1941,In_2227);
or U417 (N_417,In_1736,In_1359);
nor U418 (N_418,In_819,In_1885);
xor U419 (N_419,In_1180,In_1744);
or U420 (N_420,In_919,In_2079);
xnor U421 (N_421,In_149,In_503);
nor U422 (N_422,In_1480,In_1345);
or U423 (N_423,In_1559,In_1019);
nand U424 (N_424,In_389,In_1081);
nor U425 (N_425,In_2150,In_796);
nor U426 (N_426,In_476,In_1789);
or U427 (N_427,In_1107,In_161);
xor U428 (N_428,In_2422,In_1257);
nand U429 (N_429,In_1238,In_288);
or U430 (N_430,In_945,In_501);
and U431 (N_431,In_16,In_1228);
and U432 (N_432,In_1269,In_2095);
or U433 (N_433,In_1923,In_1557);
and U434 (N_434,In_541,In_105);
nand U435 (N_435,In_1682,In_1449);
nand U436 (N_436,In_1993,In_145);
or U437 (N_437,In_600,In_276);
nand U438 (N_438,In_595,In_958);
xnor U439 (N_439,In_1894,In_224);
xor U440 (N_440,In_140,In_1580);
xnor U441 (N_441,In_1344,In_69);
xor U442 (N_442,In_2110,In_43);
xnor U443 (N_443,In_988,In_174);
or U444 (N_444,In_1029,In_1127);
nor U445 (N_445,In_906,In_1196);
nor U446 (N_446,In_504,In_122);
or U447 (N_447,In_169,In_614);
and U448 (N_448,In_1425,In_2033);
nand U449 (N_449,In_734,In_2098);
nor U450 (N_450,In_11,In_1419);
or U451 (N_451,In_1520,In_1977);
nand U452 (N_452,In_1259,In_139);
nand U453 (N_453,In_1825,In_1761);
nand U454 (N_454,In_1008,In_2099);
or U455 (N_455,In_1756,In_2387);
nand U456 (N_456,In_1271,In_2390);
and U457 (N_457,In_1056,In_162);
and U458 (N_458,In_499,In_970);
xor U459 (N_459,In_619,In_1784);
or U460 (N_460,In_429,In_2212);
xnor U461 (N_461,In_2085,In_969);
and U462 (N_462,In_1904,In_1552);
and U463 (N_463,In_858,In_432);
or U464 (N_464,In_2428,In_1204);
nand U465 (N_465,In_628,In_542);
nor U466 (N_466,In_2041,In_854);
nor U467 (N_467,In_1547,In_2351);
xnor U468 (N_468,In_2253,In_1676);
or U469 (N_469,In_884,In_2101);
nand U470 (N_470,In_586,In_860);
nor U471 (N_471,In_926,In_2113);
xor U472 (N_472,In_2336,In_731);
or U473 (N_473,In_2498,In_2129);
nor U474 (N_474,In_667,In_801);
nor U475 (N_475,In_1303,In_1585);
xor U476 (N_476,In_1395,In_616);
xnor U477 (N_477,In_2249,In_1254);
or U478 (N_478,In_939,In_1452);
xnor U479 (N_479,In_2,In_638);
and U480 (N_480,In_873,In_361);
nor U481 (N_481,In_1733,In_714);
or U482 (N_482,In_492,In_1778);
nand U483 (N_483,In_2463,In_654);
or U484 (N_484,In_2025,In_1815);
and U485 (N_485,In_347,In_1213);
or U486 (N_486,In_107,In_2485);
or U487 (N_487,In_2102,In_370);
nand U488 (N_488,In_137,In_2310);
xor U489 (N_489,In_1272,In_1908);
or U490 (N_490,In_178,In_534);
xor U491 (N_491,In_2423,In_612);
and U492 (N_492,In_674,In_1834);
nor U493 (N_493,In_621,In_1700);
and U494 (N_494,In_2186,In_2145);
and U495 (N_495,In_1548,In_1296);
xor U496 (N_496,In_200,In_573);
or U497 (N_497,In_606,In_2484);
xor U498 (N_498,In_1092,In_363);
and U499 (N_499,In_419,In_1267);
xnor U500 (N_500,In_1845,In_1519);
nor U501 (N_501,In_2399,In_727);
xor U502 (N_502,In_1314,In_151);
or U503 (N_503,In_1506,In_1623);
and U504 (N_504,In_1931,In_610);
xor U505 (N_505,In_1810,In_1701);
or U506 (N_506,In_2326,In_392);
nand U507 (N_507,In_332,In_2097);
nand U508 (N_508,In_1114,In_1438);
and U509 (N_509,In_1699,In_40);
nand U510 (N_510,In_526,In_1192);
xor U511 (N_511,In_1283,In_1562);
nor U512 (N_512,In_1546,In_539);
or U513 (N_513,In_1942,In_279);
nor U514 (N_514,In_1753,In_177);
nor U515 (N_515,In_1646,In_1518);
and U516 (N_516,In_1596,In_932);
and U517 (N_517,In_1110,In_821);
nor U518 (N_518,In_2010,In_228);
and U519 (N_519,In_413,In_418);
nand U520 (N_520,In_1188,In_461);
xor U521 (N_521,In_701,In_366);
nand U522 (N_522,In_2261,In_689);
xnor U523 (N_523,In_397,In_93);
nand U524 (N_524,In_669,In_2292);
xnor U525 (N_525,In_977,In_188);
nor U526 (N_526,In_853,In_1473);
nand U527 (N_527,In_1363,In_1426);
and U528 (N_528,In_1098,In_2342);
nor U529 (N_529,In_1972,In_2265);
xnor U530 (N_530,In_2291,In_511);
xnor U531 (N_531,In_214,In_1149);
or U532 (N_532,In_961,In_2487);
nor U533 (N_533,In_367,In_670);
or U534 (N_534,In_908,In_1637);
and U535 (N_535,In_2044,In_1544);
or U536 (N_536,In_1891,In_2496);
xnor U537 (N_537,In_317,In_1088);
xor U538 (N_538,In_182,In_1195);
nand U539 (N_539,In_2413,In_1164);
nand U540 (N_540,In_848,In_2452);
nor U541 (N_541,In_750,In_1662);
and U542 (N_542,In_452,In_1343);
nand U543 (N_543,In_34,In_1001);
or U544 (N_544,In_921,In_1723);
or U545 (N_545,In_1586,In_2273);
or U546 (N_546,In_785,In_2037);
xnor U547 (N_547,In_2019,In_1455);
xor U548 (N_548,In_1715,In_2000);
or U549 (N_549,In_1398,In_259);
or U550 (N_550,In_1315,In_393);
nand U551 (N_551,In_2012,In_2138);
and U552 (N_552,In_688,In_2324);
xnor U553 (N_553,In_1,In_1175);
nand U554 (N_554,In_1598,In_1030);
nor U555 (N_555,In_1850,In_2021);
nand U556 (N_556,In_207,In_1323);
xor U557 (N_557,In_2448,In_603);
nor U558 (N_558,In_1512,In_2107);
nor U559 (N_559,In_566,In_1882);
nand U560 (N_560,In_705,In_1336);
and U561 (N_561,In_310,In_2163);
nand U562 (N_562,In_127,In_19);
nor U563 (N_563,In_2022,In_536);
nor U564 (N_564,In_1986,In_1862);
xnor U565 (N_565,In_355,In_2269);
nand U566 (N_566,In_2473,In_1079);
xor U567 (N_567,In_2206,In_440);
nor U568 (N_568,In_491,In_17);
nand U569 (N_569,In_613,In_1244);
nand U570 (N_570,In_1136,In_60);
or U571 (N_571,In_1138,In_1626);
nor U572 (N_572,In_203,In_13);
nor U573 (N_573,In_424,In_832);
or U574 (N_574,In_838,In_687);
nor U575 (N_575,In_337,In_956);
or U576 (N_576,In_2380,In_1161);
xnor U577 (N_577,In_4,In_2320);
xor U578 (N_578,In_2043,In_1930);
nor U579 (N_579,In_1072,In_287);
or U580 (N_580,In_764,In_1016);
and U581 (N_581,In_278,In_1484);
nor U582 (N_582,In_2486,In_2317);
or U583 (N_583,In_134,In_914);
nand U584 (N_584,In_2361,In_965);
and U585 (N_585,In_2382,In_2439);
or U586 (N_586,In_535,In_1439);
nand U587 (N_587,In_2082,In_251);
nand U588 (N_588,In_1935,In_81);
nor U589 (N_589,In_995,In_1842);
or U590 (N_590,In_1064,In_191);
xnor U591 (N_591,In_1216,In_771);
and U592 (N_592,In_2368,In_1895);
xor U593 (N_593,In_1171,In_1832);
and U594 (N_594,In_1830,In_462);
xnor U595 (N_595,In_1446,In_1650);
nand U596 (N_596,In_2404,In_143);
and U597 (N_597,In_1041,In_1273);
nor U598 (N_598,In_842,In_348);
or U599 (N_599,In_716,In_1349);
nor U600 (N_600,In_1812,In_165);
xor U601 (N_601,In_2075,In_1086);
nand U602 (N_602,In_1358,In_1168);
and U603 (N_603,In_2071,In_1073);
nand U604 (N_604,In_664,In_1231);
and U605 (N_605,In_1470,In_1681);
xor U606 (N_606,In_672,In_1304);
and U607 (N_607,In_2023,In_27);
nand U608 (N_608,In_292,In_1351);
nand U609 (N_609,In_2233,In_1248);
or U610 (N_610,In_290,In_1966);
and U611 (N_611,In_199,In_2220);
and U612 (N_612,In_155,In_1183);
xor U613 (N_613,In_1783,In_706);
xnor U614 (N_614,In_690,In_281);
and U615 (N_615,In_729,In_242);
or U616 (N_616,In_2288,In_2450);
or U617 (N_617,In_1843,In_2030);
nand U618 (N_618,In_533,In_1505);
nand U619 (N_619,In_71,In_1605);
nor U620 (N_620,In_508,In_2352);
and U621 (N_621,In_87,In_121);
xor U622 (N_622,In_449,In_430);
and U623 (N_623,In_2343,In_1457);
xnor U624 (N_624,In_2005,In_67);
nor U625 (N_625,In_702,In_889);
and U626 (N_626,In_1014,In_1070);
nor U627 (N_627,In_1851,In_1712);
xor U628 (N_628,N_275,In_1078);
nand U629 (N_629,In_2285,N_496);
nor U630 (N_630,N_148,N_497);
xor U631 (N_631,In_1587,N_481);
or U632 (N_632,In_799,In_1872);
xnor U633 (N_633,N_45,In_1301);
xor U634 (N_634,N_249,In_1907);
or U635 (N_635,In_1412,In_2247);
nor U636 (N_636,In_1758,In_1531);
nand U637 (N_637,N_419,N_454);
xor U638 (N_638,In_1022,In_934);
xor U639 (N_639,In_1721,In_709);
xor U640 (N_640,In_2245,N_549);
or U641 (N_641,In_1117,In_2379);
xor U642 (N_642,In_2106,In_2194);
or U643 (N_643,In_2307,N_75);
or U644 (N_644,N_290,N_615);
xor U645 (N_645,N_282,In_1619);
nand U646 (N_646,In_1879,In_1404);
and U647 (N_647,In_354,N_308);
xor U648 (N_648,N_73,In_1134);
or U649 (N_649,In_659,In_465);
or U650 (N_650,N_293,In_1126);
nor U651 (N_651,In_2197,In_546);
or U652 (N_652,N_581,N_318);
nor U653 (N_653,N_90,N_239);
or U654 (N_654,In_683,In_282);
nand U655 (N_655,N_68,N_622);
xnor U656 (N_656,In_1184,In_2424);
xnor U657 (N_657,In_2258,N_234);
or U658 (N_658,N_528,In_1927);
nor U659 (N_659,In_886,N_217);
or U660 (N_660,In_2341,N_379);
or U661 (N_661,In_1549,In_1309);
nor U662 (N_662,In_1691,In_175);
nor U663 (N_663,N_142,In_74);
nand U664 (N_664,In_168,In_1992);
and U665 (N_665,In_2086,N_563);
nand U666 (N_666,N_594,In_1631);
and U667 (N_667,In_1181,In_1792);
nand U668 (N_668,In_1462,N_238);
nand U669 (N_669,In_1926,In_2134);
xnor U670 (N_670,In_357,In_485);
xor U671 (N_671,In_645,In_1230);
nand U672 (N_672,In_1679,In_1145);
nor U673 (N_673,In_30,N_325);
and U674 (N_674,N_228,In_180);
xnor U675 (N_675,In_236,In_1429);
xnor U676 (N_676,In_2016,In_237);
nor U677 (N_677,In_1924,In_545);
xnor U678 (N_678,N_447,In_2357);
and U679 (N_679,In_751,In_1638);
xor U680 (N_680,In_718,In_1084);
xnor U681 (N_681,In_896,N_368);
and U682 (N_682,In_368,In_249);
or U683 (N_683,N_456,In_1985);
nand U684 (N_684,In_1725,In_1440);
nor U685 (N_685,In_811,In_1779);
nand U686 (N_686,In_1837,In_299);
nor U687 (N_687,In_1826,N_138);
nand U688 (N_688,In_1507,In_102);
nor U689 (N_689,N_477,In_2222);
xnor U690 (N_690,In_1624,In_2032);
or U691 (N_691,N_403,In_1341);
or U692 (N_692,N_258,In_898);
xnor U693 (N_693,In_1212,In_824);
nand U694 (N_694,N_585,In_1040);
xnor U695 (N_695,In_720,In_1692);
nand U696 (N_696,N_272,N_543);
and U697 (N_697,N_190,In_2027);
or U698 (N_698,In_1960,N_40);
and U699 (N_699,In_364,In_887);
nor U700 (N_700,N_401,N_386);
or U701 (N_701,In_1450,In_1397);
xnor U702 (N_702,N_313,In_868);
nor U703 (N_703,In_1922,In_1755);
nor U704 (N_704,N_226,N_539);
and U705 (N_705,N_112,In_1339);
nand U706 (N_706,In_1157,N_84);
xnor U707 (N_707,In_2052,In_1160);
nand U708 (N_708,In_1582,In_2255);
xnor U709 (N_709,N_338,N_606);
nor U710 (N_710,N_515,N_546);
nor U711 (N_711,N_46,In_295);
xor U712 (N_712,In_1569,In_458);
and U713 (N_713,N_151,N_101);
and U714 (N_714,In_238,In_1952);
xnor U715 (N_715,N_437,N_186);
xnor U716 (N_716,In_1262,In_1054);
xor U717 (N_717,In_2153,In_2278);
nor U718 (N_718,N_455,In_289);
or U719 (N_719,In_2348,In_304);
nor U720 (N_720,In_2211,In_2398);
nand U721 (N_721,In_1006,N_276);
or U722 (N_722,In_1407,N_559);
and U723 (N_723,N_233,In_1910);
xnor U724 (N_724,In_2112,In_233);
xor U725 (N_725,In_1946,In_385);
and U726 (N_726,In_1595,In_518);
or U727 (N_727,In_665,In_959);
nand U728 (N_728,N_411,In_878);
nor U729 (N_729,N_257,In_1350);
and U730 (N_730,In_2162,In_2289);
and U731 (N_731,In_698,In_2297);
and U732 (N_732,In_609,N_81);
and U733 (N_733,N_146,In_828);
nor U734 (N_734,In_494,N_416);
nor U735 (N_735,N_48,In_101);
xor U736 (N_736,In_1459,In_202);
or U737 (N_737,In_2309,In_1297);
xnor U738 (N_738,N_518,In_572);
xor U739 (N_739,In_876,In_1865);
or U740 (N_740,In_1994,In_201);
nor U741 (N_741,N_610,N_444);
nor U742 (N_742,In_185,In_591);
nor U743 (N_743,In_1625,In_537);
xor U744 (N_744,In_1444,N_369);
or U745 (N_745,In_1564,In_967);
or U746 (N_746,N_345,In_935);
and U747 (N_747,In_408,In_2088);
or U748 (N_748,N_591,In_708);
nand U749 (N_749,In_443,In_550);
or U750 (N_750,N_443,In_451);
and U751 (N_751,N_457,In_2060);
nor U752 (N_752,In_991,In_804);
nand U753 (N_753,In_98,In_1906);
nor U754 (N_754,N_578,N_87);
nand U755 (N_755,In_32,In_346);
nor U756 (N_756,In_607,In_1146);
nand U757 (N_757,In_631,In_2039);
or U758 (N_758,In_2209,In_1813);
nor U759 (N_759,N_195,In_1751);
nand U760 (N_760,N_270,In_2154);
and U761 (N_761,In_1683,In_1819);
nor U762 (N_762,In_755,In_1978);
xor U763 (N_763,N_202,In_660);
nor U764 (N_764,N_114,In_692);
and U765 (N_765,N_450,In_2338);
xor U766 (N_766,In_1067,In_1540);
and U767 (N_767,N_501,N_245);
nor U768 (N_768,In_2268,In_1202);
nor U769 (N_769,In_1391,In_2279);
nand U770 (N_770,In_1392,In_1674);
and U771 (N_771,In_1141,N_38);
or U772 (N_772,N_584,In_2451);
and U773 (N_773,N_179,In_1863);
nand U774 (N_774,In_319,N_378);
nor U775 (N_775,In_2069,In_1588);
xnor U776 (N_776,In_1193,In_1802);
nor U777 (N_777,In_761,In_625);
or U778 (N_778,In_839,In_1465);
or U779 (N_779,N_434,N_418);
and U780 (N_780,N_157,N_343);
nand U781 (N_781,In_1206,In_1685);
or U782 (N_782,In_1956,In_1243);
nor U783 (N_783,In_212,N_392);
nand U784 (N_784,N_50,In_1860);
nand U785 (N_785,In_1173,In_1065);
xor U786 (N_786,N_96,In_782);
and U787 (N_787,In_818,In_2048);
or U788 (N_788,In_684,N_25);
and U789 (N_789,N_32,N_211);
or U790 (N_790,In_2470,N_82);
and U791 (N_791,N_519,N_145);
and U792 (N_792,In_576,In_2047);
and U793 (N_793,In_879,In_960);
nor U794 (N_794,N_13,N_18);
and U795 (N_795,In_671,N_570);
nor U796 (N_796,In_1591,In_1342);
or U797 (N_797,In_1772,N_163);
or U798 (N_798,In_1293,In_2210);
or U799 (N_799,In_286,In_916);
nand U800 (N_800,N_110,In_402);
nand U801 (N_801,In_2122,In_1454);
or U802 (N_802,N_511,In_187);
nor U803 (N_803,N_352,In_1521);
or U804 (N_804,In_1165,In_358);
nand U805 (N_805,In_552,N_587);
nor U806 (N_806,In_78,In_1912);
and U807 (N_807,In_1224,In_1680);
nand U808 (N_808,N_216,In_809);
nand U809 (N_809,N_564,In_506);
nor U810 (N_810,In_1037,N_199);
nand U811 (N_811,N_230,In_1577);
nand U812 (N_812,In_2136,In_8);
nor U813 (N_813,N_430,In_1000);
nor U814 (N_814,N_473,In_306);
or U815 (N_815,In_1020,In_1277);
xnor U816 (N_816,N_404,In_1694);
nor U817 (N_817,N_126,In_1249);
nor U818 (N_818,In_830,N_147);
nor U819 (N_819,In_2096,N_162);
nand U820 (N_820,N_330,In_2374);
nor U821 (N_821,In_964,In_1809);
nand U822 (N_822,In_704,In_2354);
or U823 (N_823,N_49,In_1498);
or U824 (N_824,In_1799,In_1968);
nor U825 (N_825,N_588,In_1275);
xor U826 (N_826,N_312,In_1422);
nor U827 (N_827,In_1785,In_2057);
or U828 (N_828,In_391,N_280);
nor U829 (N_829,In_94,In_480);
or U830 (N_830,N_458,In_2391);
nand U831 (N_831,In_1786,N_452);
and U832 (N_832,N_253,N_507);
nor U833 (N_833,In_339,In_1485);
xor U834 (N_834,N_494,In_1693);
nand U835 (N_835,N_149,N_175);
nand U836 (N_836,In_1200,In_2040);
xor U837 (N_837,In_1108,In_415);
nor U838 (N_838,N_144,In_1115);
nand U839 (N_839,In_1913,In_1741);
xnor U840 (N_840,N_505,In_66);
xnor U841 (N_841,N_123,In_1747);
and U842 (N_842,N_83,N_76);
nand U843 (N_843,In_1099,In_1416);
or U844 (N_844,N_53,N_486);
xor U845 (N_845,N_43,N_139);
or U846 (N_846,N_592,In_1306);
or U847 (N_847,In_407,In_1974);
nor U848 (N_848,In_2165,In_1144);
or U849 (N_849,In_1491,In_2415);
nor U850 (N_850,In_2286,In_815);
nand U851 (N_851,N_347,In_1374);
or U852 (N_852,N_530,N_471);
nor U853 (N_853,N_106,N_105);
or U854 (N_854,In_2238,In_2056);
or U855 (N_855,In_1435,In_1468);
xor U856 (N_856,N_244,N_509);
xor U857 (N_857,N_17,In_775);
or U858 (N_858,N_281,N_618);
or U859 (N_859,N_374,N_609);
nand U860 (N_860,In_1897,N_246);
or U861 (N_861,In_420,N_260);
and U862 (N_862,In_1371,N_356);
nor U863 (N_863,In_1097,In_807);
nand U864 (N_864,In_1773,In_1189);
or U865 (N_865,In_1948,N_184);
or U866 (N_866,N_520,In_1012);
and U867 (N_867,In_110,In_1610);
xnor U868 (N_868,In_112,In_1916);
or U869 (N_869,In_1917,N_522);
nor U870 (N_870,N_78,N_33);
nor U871 (N_871,In_2411,N_319);
or U872 (N_872,In_992,In_1051);
xor U873 (N_873,N_580,In_2248);
xnor U874 (N_874,In_1159,In_2189);
and U875 (N_875,In_255,In_266);
nand U876 (N_876,In_2182,N_598);
nor U877 (N_877,In_1754,N_362);
and U878 (N_878,In_963,N_116);
or U879 (N_879,In_1035,N_367);
or U880 (N_880,In_1800,N_174);
xnor U881 (N_881,In_256,In_438);
and U882 (N_882,In_170,N_200);
and U883 (N_883,In_2184,In_840);
or U884 (N_884,In_2201,N_115);
and U885 (N_885,In_1555,In_44);
nor U886 (N_886,N_31,In_2296);
or U887 (N_887,N_420,N_534);
xor U888 (N_888,N_269,In_726);
nor U889 (N_889,N_196,In_2161);
xnor U890 (N_890,N_267,In_1261);
or U891 (N_891,In_1158,In_699);
nand U892 (N_892,In_994,N_423);
nor U893 (N_893,N_213,In_910);
xnor U894 (N_894,In_1445,In_2133);
xnor U895 (N_895,In_1285,In_2217);
xor U896 (N_896,N_476,In_2459);
nand U897 (N_897,In_2366,In_928);
nor U898 (N_898,In_2311,In_1936);
nor U899 (N_899,In_2313,N_243);
nor U900 (N_900,N_479,In_1678);
and U901 (N_901,N_574,In_1705);
and U902 (N_902,In_1958,N_209);
nand U903 (N_903,N_548,In_1433);
or U904 (N_904,In_1080,In_1633);
or U905 (N_905,In_585,In_1076);
xor U906 (N_906,N_324,N_540);
nand U907 (N_907,In_2216,In_1965);
nand U908 (N_908,In_1291,N_601);
nor U909 (N_909,In_130,In_1299);
xor U910 (N_910,In_2226,In_1335);
and U911 (N_911,In_328,In_1787);
xnor U912 (N_912,In_1453,In_404);
and U913 (N_913,In_482,In_693);
or U914 (N_914,In_1969,In_2223);
and U915 (N_915,In_1848,In_1063);
nor U916 (N_916,In_1233,N_26);
or U917 (N_917,In_2028,In_1045);
nor U918 (N_918,In_1998,In_800);
or U919 (N_919,In_483,In_760);
nand U920 (N_920,N_394,In_235);
xor U921 (N_921,N_611,In_741);
nor U922 (N_922,In_2372,N_487);
xor U923 (N_923,N_93,N_366);
nor U924 (N_924,N_317,In_2489);
xor U925 (N_925,N_133,N_541);
and U926 (N_926,In_135,N_339);
or U927 (N_927,N_391,N_532);
and U928 (N_928,N_254,In_1537);
and U929 (N_929,N_129,In_450);
and U930 (N_930,In_2408,In_581);
nor U931 (N_931,N_252,In_1131);
nand U932 (N_932,N_484,N_306);
nand U933 (N_933,N_172,In_1990);
or U934 (N_934,In_1111,N_582);
or U935 (N_935,In_179,In_1628);
nor U936 (N_936,In_1003,N_499);
nor U937 (N_937,In_108,N_376);
and U938 (N_938,In_865,In_561);
nor U939 (N_939,In_1944,N_117);
nor U940 (N_940,N_135,N_316);
nand U941 (N_941,In_1933,N_399);
xnor U942 (N_942,N_346,In_308);
xnor U943 (N_943,N_396,In_1496);
xnor U944 (N_944,N_71,N_506);
nor U945 (N_945,In_1919,N_62);
nor U946 (N_946,In_1232,In_578);
or U947 (N_947,In_769,N_223);
nor U948 (N_948,In_1901,N_562);
or U949 (N_949,In_445,N_371);
nor U950 (N_950,N_554,In_1673);
nand U951 (N_951,In_2137,In_850);
and U952 (N_952,In_2064,In_323);
nand U953 (N_953,In_602,In_1609);
and U954 (N_954,In_146,In_1932);
nor U955 (N_955,In_1069,In_1319);
nor U956 (N_956,In_2300,N_7);
xor U957 (N_957,In_615,In_641);
and U958 (N_958,N_607,In_893);
nor U959 (N_959,In_22,N_264);
nand U960 (N_960,In_1125,N_287);
or U961 (N_961,In_1266,N_201);
or U962 (N_962,In_131,In_1554);
and U963 (N_963,In_1044,N_576);
nor U964 (N_964,In_611,In_2218);
xnor U965 (N_965,In_1657,N_55);
xor U966 (N_966,N_121,In_1590);
nor U967 (N_967,N_19,N_314);
and U968 (N_968,In_781,N_44);
nand U969 (N_969,In_1298,In_184);
nor U970 (N_970,In_1798,N_173);
nand U971 (N_971,In_1703,N_185);
nand U972 (N_972,In_1096,N_355);
and U973 (N_973,In_86,In_558);
nand U974 (N_974,N_74,In_1689);
xor U975 (N_975,In_2384,N_85);
nand U976 (N_976,In_1811,N_536);
or U977 (N_977,In_437,N_417);
or U978 (N_978,N_279,N_165);
or U979 (N_979,N_586,In_911);
xnor U980 (N_980,In_1530,In_1928);
nand U981 (N_981,N_459,In_1235);
and U982 (N_982,N_544,In_962);
nor U983 (N_983,N_359,In_943);
nand U984 (N_984,In_157,In_116);
nand U985 (N_985,N_525,In_1436);
and U986 (N_986,In_1005,In_1690);
nand U987 (N_987,N_331,N_448);
nand U988 (N_988,In_2434,N_159);
nand U989 (N_989,In_877,N_322);
xnor U990 (N_990,N_514,In_1615);
nand U991 (N_991,In_454,N_560);
nor U992 (N_992,N_590,In_944);
or U993 (N_993,In_1367,N_94);
nor U994 (N_994,In_1074,N_132);
nand U995 (N_995,N_4,In_1050);
nand U996 (N_996,In_565,In_1604);
nand U997 (N_997,In_682,N_357);
xnor U998 (N_998,In_1017,N_27);
or U999 (N_999,N_99,In_525);
and U1000 (N_1000,In_835,In_1824);
and U1001 (N_1001,In_2128,In_986);
and U1002 (N_1002,N_98,In_1818);
nand U1003 (N_1003,In_1945,N_69);
and U1004 (N_1004,N_206,In_99);
or U1005 (N_1005,In_789,N_298);
or U1006 (N_1006,In_1062,N_189);
nand U1007 (N_1007,In_1207,In_2031);
or U1008 (N_1008,N_266,N_155);
nand U1009 (N_1009,In_1963,In_5);
nor U1010 (N_1010,N_111,In_479);
or U1011 (N_1011,N_182,In_63);
and U1012 (N_1012,In_584,In_2373);
nor U1013 (N_1013,In_24,N_571);
xor U1014 (N_1014,N_288,N_198);
and U1015 (N_1015,In_52,In_736);
nand U1016 (N_1016,In_2445,In_394);
or U1017 (N_1017,In_91,In_2243);
or U1018 (N_1018,In_274,In_730);
and U1019 (N_1019,In_1858,In_975);
or U1020 (N_1020,In_1726,In_2050);
and U1021 (N_1021,N_136,In_1038);
and U1022 (N_1022,N_205,In_416);
or U1023 (N_1023,N_375,In_982);
and U1024 (N_1024,In_577,N_320);
or U1025 (N_1025,In_1644,In_1198);
nand U1026 (N_1026,N_194,In_937);
nor U1027 (N_1027,In_1869,N_614);
nand U1028 (N_1028,N_523,N_168);
or U1029 (N_1029,N_208,N_241);
and U1030 (N_1030,N_542,In_1137);
nand U1031 (N_1031,N_24,In_2092);
nor U1032 (N_1032,N_310,N_161);
nor U1033 (N_1033,In_575,In_1503);
nor U1034 (N_1034,N_551,In_2284);
nor U1035 (N_1035,In_1185,In_2175);
and U1036 (N_1036,In_460,N_524);
nand U1037 (N_1037,In_345,N_255);
xor U1038 (N_1038,In_1278,In_2419);
and U1039 (N_1039,In_1052,N_436);
or U1040 (N_1040,N_231,N_500);
and U1041 (N_1041,In_2478,N_251);
nand U1042 (N_1042,In_267,In_183);
nand U1043 (N_1043,In_890,N_166);
and U1044 (N_1044,In_1251,In_2246);
or U1045 (N_1045,In_2449,N_227);
or U1046 (N_1046,In_2091,In_490);
or U1047 (N_1047,In_1481,In_866);
nor U1048 (N_1048,In_1641,In_446);
nor U1049 (N_1049,In_82,N_91);
or U1050 (N_1050,N_229,N_140);
and U1051 (N_1051,In_2276,N_412);
or U1052 (N_1052,In_564,In_257);
nor U1053 (N_1053,In_21,N_464);
nand U1054 (N_1054,N_302,In_263);
or U1055 (N_1055,N_169,In_2093);
and U1056 (N_1056,In_617,In_2080);
nand U1057 (N_1057,In_2143,N_303);
nor U1058 (N_1058,In_758,In_1377);
xnor U1059 (N_1059,In_2389,N_285);
and U1060 (N_1060,In_574,In_2346);
and U1061 (N_1061,N_365,In_2287);
xor U1062 (N_1062,In_2254,In_847);
or U1063 (N_1063,In_2116,In_216);
nor U1064 (N_1064,In_159,N_273);
nand U1065 (N_1065,In_2319,N_183);
and U1066 (N_1066,In_1838,In_803);
or U1067 (N_1067,In_662,In_70);
or U1068 (N_1068,In_1737,In_1177);
nor U1069 (N_1069,In_1629,In_1634);
nand U1070 (N_1070,In_2330,In_1209);
nand U1071 (N_1071,In_1042,In_487);
nand U1072 (N_1072,N_335,In_1493);
xnor U1073 (N_1073,N_382,In_1513);
and U1074 (N_1074,In_221,In_1421);
nor U1075 (N_1075,In_2347,In_663);
nand U1076 (N_1076,N_408,N_619);
nand U1077 (N_1077,In_470,In_2045);
and U1078 (N_1078,In_464,In_160);
nor U1079 (N_1079,In_1814,In_2173);
or U1080 (N_1080,In_1327,In_1077);
nand U1081 (N_1081,In_661,In_1116);
and U1082 (N_1082,N_535,In_529);
nand U1083 (N_1083,N_435,In_1443);
xnor U1084 (N_1084,In_2224,N_309);
or U1085 (N_1085,In_907,In_1528);
nand U1086 (N_1086,In_540,In_646);
or U1087 (N_1087,In_2294,N_440);
xor U1088 (N_1088,N_573,In_1140);
nor U1089 (N_1089,In_36,In_296);
nor U1090 (N_1090,In_2365,In_1854);
xnor U1091 (N_1091,In_2229,In_605);
xor U1092 (N_1092,N_415,In_141);
xor U1093 (N_1093,N_214,In_92);
xnor U1094 (N_1094,In_210,In_2418);
nor U1095 (N_1095,In_2073,In_307);
or U1096 (N_1096,N_120,N_192);
or U1097 (N_1097,In_515,In_2001);
and U1098 (N_1098,In_863,In_1790);
nand U1099 (N_1099,In_1361,In_1509);
and U1100 (N_1100,N_153,N_593);
nor U1101 (N_1101,N_222,N_623);
and U1102 (N_1102,N_589,N_383);
and U1103 (N_1103,N_472,N_224);
xnor U1104 (N_1104,In_2474,N_572);
nor U1105 (N_1105,In_936,N_261);
and U1106 (N_1106,N_315,In_377);
nor U1107 (N_1107,N_15,In_268);
or U1108 (N_1108,In_2377,In_1089);
xnor U1109 (N_1109,N_600,In_1671);
nand U1110 (N_1110,In_1523,N_107);
nand U1111 (N_1111,In_1387,In_920);
nor U1112 (N_1112,In_1760,In_1855);
and U1113 (N_1113,N_152,In_2063);
and U1114 (N_1114,N_529,N_475);
nor U1115 (N_1115,In_132,In_1762);
and U1116 (N_1116,In_1388,N_22);
or U1117 (N_1117,In_360,N_334);
nand U1118 (N_1118,In_516,In_2461);
nand U1119 (N_1119,N_512,In_749);
or U1120 (N_1120,In_2360,In_1112);
xnor U1121 (N_1121,N_97,In_1602);
xnor U1122 (N_1122,In_713,In_1551);
or U1123 (N_1123,N_328,In_390);
or U1124 (N_1124,In_1659,In_666);
nand U1125 (N_1125,In_557,In_1263);
and U1126 (N_1126,In_2072,In_215);
xor U1127 (N_1127,In_676,N_427);
or U1128 (N_1128,N_34,N_483);
nor U1129 (N_1129,In_444,In_1655);
nand U1130 (N_1130,In_902,N_402);
or U1131 (N_1131,N_568,In_1508);
xnor U1132 (N_1132,In_194,In_1759);
nor U1133 (N_1133,N_495,N_545);
nor U1134 (N_1134,In_1766,In_1980);
or U1135 (N_1135,In_1210,In_1034);
nor U1136 (N_1136,In_223,In_1222);
and U1137 (N_1137,In_2329,N_240);
nand U1138 (N_1138,In_582,N_277);
nand U1139 (N_1139,In_1252,In_252);
nand U1140 (N_1140,In_335,In_1442);
xnor U1141 (N_1141,N_156,In_1516);
nand U1142 (N_1142,In_626,In_2176);
or U1143 (N_1143,In_1947,In_119);
and U1144 (N_1144,In_2406,N_550);
or U1145 (N_1145,N_109,N_52);
and U1146 (N_1146,In_1563,In_1698);
xor U1147 (N_1147,In_624,In_543);
xnor U1148 (N_1148,In_1396,In_2409);
xnor U1149 (N_1149,In_38,N_250);
nand U1150 (N_1150,In_1574,N_292);
and U1151 (N_1151,In_2125,In_89);
xor U1152 (N_1152,N_12,In_1049);
xnor U1153 (N_1153,N_204,N_389);
xnor U1154 (N_1154,In_837,N_360);
nor U1155 (N_1155,In_1943,N_351);
nand U1156 (N_1156,N_624,N_265);
nand U1157 (N_1157,N_89,In_375);
nor U1158 (N_1158,In_262,In_371);
nor U1159 (N_1159,In_2272,N_177);
nor U1160 (N_1160,In_794,In_2385);
xnor U1161 (N_1161,N_425,In_2159);
xor U1162 (N_1162,In_1268,In_1589);
nor U1163 (N_1163,In_305,In_633);
or U1164 (N_1164,In_880,In_1384);
and U1165 (N_1165,N_321,N_336);
xor U1166 (N_1166,In_795,N_187);
nand U1167 (N_1167,In_220,In_1658);
nor U1168 (N_1168,In_2417,N_616);
xnor U1169 (N_1169,In_1543,In_2002);
xnor U1170 (N_1170,N_236,N_441);
xor U1171 (N_1171,In_651,N_513);
nor U1172 (N_1172,N_478,In_2420);
and U1173 (N_1173,In_1448,N_323);
or U1174 (N_1174,In_954,In_1617);
nor U1175 (N_1175,N_384,In_1401);
or U1176 (N_1176,In_1492,In_1156);
nor U1177 (N_1177,In_1039,N_381);
nand U1178 (N_1178,In_1794,In_1476);
and U1179 (N_1179,N_428,N_54);
nand U1180 (N_1180,In_211,In_1214);
nand U1181 (N_1181,In_2231,N_510);
nor U1182 (N_1182,N_221,N_406);
xor U1183 (N_1183,In_1162,In_1382);
xnor U1184 (N_1184,N_63,N_36);
and U1185 (N_1185,In_1959,N_304);
and U1186 (N_1186,In_1057,In_2443);
xnor U1187 (N_1187,In_2115,In_2180);
nor U1188 (N_1188,In_983,In_895);
xnor U1189 (N_1189,N_3,N_370);
xor U1190 (N_1190,In_2306,In_2393);
nand U1191 (N_1191,In_1656,In_405);
and U1192 (N_1192,In_904,N_262);
nor U1193 (N_1193,N_125,In_356);
or U1194 (N_1194,In_1663,In_2215);
nand U1195 (N_1195,N_466,N_188);
nand U1196 (N_1196,In_1501,N_617);
xor U1197 (N_1197,In_1579,In_817);
xnor U1198 (N_1198,In_1418,In_154);
nor U1199 (N_1199,In_53,In_1714);
or U1200 (N_1200,In_1739,In_2139);
or U1201 (N_1201,N_556,In_164);
xor U1202 (N_1202,In_2011,In_864);
and U1203 (N_1203,In_1043,N_395);
xor U1204 (N_1204,In_2321,N_88);
or U1205 (N_1205,N_327,In_512);
xnor U1206 (N_1206,In_2274,In_362);
or U1207 (N_1207,In_1488,N_268);
xor U1208 (N_1208,In_283,In_1511);
xnor U1209 (N_1209,In_1524,N_259);
xnor U1210 (N_1210,In_1295,In_831);
nand U1211 (N_1211,In_343,In_313);
xnor U1212 (N_1212,In_1317,In_2191);
xnor U1213 (N_1213,In_593,In_2236);
nand U1214 (N_1214,In_1796,In_411);
nor U1215 (N_1215,N_143,In_1724);
nor U1216 (N_1216,In_226,In_2147);
nor U1217 (N_1217,In_1321,In_2312);
xor U1218 (N_1218,In_1630,In_1856);
or U1219 (N_1219,In_1527,N_393);
and U1220 (N_1220,In_1566,In_1716);
or U1221 (N_1221,N_526,N_491);
nor U1222 (N_1222,In_2059,N_141);
xnor U1223 (N_1223,N_289,N_6);
and U1224 (N_1224,In_18,In_3);
or U1225 (N_1225,In_58,In_1765);
xnor U1226 (N_1226,In_996,N_47);
nor U1227 (N_1227,In_1686,In_1874);
and U1228 (N_1228,In_1967,N_2);
nor U1229 (N_1229,In_1849,In_1688);
nand U1230 (N_1230,In_1687,N_439);
or U1231 (N_1231,In_1816,In_859);
or U1232 (N_1232,In_1274,In_2386);
nand U1233 (N_1233,In_1167,N_604);
or U1234 (N_1234,N_59,In_1999);
or U1235 (N_1235,N_0,N_503);
xor U1236 (N_1236,In_1461,N_620);
and U1237 (N_1237,N_414,In_1205);
nand U1238 (N_1238,In_2427,In_1241);
or U1239 (N_1239,N_10,N_176);
xnor U1240 (N_1240,N_599,In_2203);
nor U1241 (N_1241,N_533,N_295);
xnor U1242 (N_1242,In_1770,In_1661);
and U1243 (N_1243,N_461,N_555);
nand U1244 (N_1244,In_2087,In_2171);
nand U1245 (N_1245,In_192,In_1197);
nand U1246 (N_1246,In_2392,In_2146);
nor U1247 (N_1247,N_353,In_1201);
nand U1248 (N_1248,In_1191,N_11);
and U1249 (N_1249,In_1356,In_933);
nand U1250 (N_1250,N_39,N_833);
nand U1251 (N_1251,N_299,N_769);
nor U1252 (N_1252,N_1070,N_170);
or U1253 (N_1253,In_48,N_820);
and U1254 (N_1254,In_1360,N_803);
xor U1255 (N_1255,N_809,In_844);
xor U1256 (N_1256,N_861,N_908);
xor U1257 (N_1257,In_985,N_407);
and U1258 (N_1258,N_891,N_297);
xnor U1259 (N_1259,N_900,N_1014);
nor U1260 (N_1260,N_158,N_332);
nor U1261 (N_1261,In_2270,N_815);
or U1262 (N_1262,N_1003,N_978);
nor U1263 (N_1263,In_1424,N_1060);
and U1264 (N_1264,N_717,In_423);
nor U1265 (N_1265,N_921,N_735);
nor U1266 (N_1266,N_877,N_687);
nand U1267 (N_1267,N_1165,N_795);
and U1268 (N_1268,N_1219,In_142);
or U1269 (N_1269,In_1463,In_2196);
nand U1270 (N_1270,N_489,N_807);
or U1271 (N_1271,In_400,N_558);
and U1272 (N_1272,In_1211,N_1052);
or U1273 (N_1273,In_329,N_349);
and U1274 (N_1274,In_172,In_2381);
nor U1275 (N_1275,N_1126,In_735);
and U1276 (N_1276,In_639,N_1193);
xor U1277 (N_1277,N_1128,N_1145);
and U1278 (N_1278,N_1185,N_1215);
and U1279 (N_1279,N_1137,In_786);
xnor U1280 (N_1280,N_761,N_79);
nor U1281 (N_1281,N_892,N_685);
nand U1282 (N_1282,N_993,In_1066);
or U1283 (N_1283,N_970,In_1270);
or U1284 (N_1284,In_1122,N_719);
nor U1285 (N_1285,N_1053,In_2074);
nor U1286 (N_1286,In_351,N_372);
nor U1287 (N_1287,N_344,In_469);
and U1288 (N_1288,N_1043,In_1265);
xnor U1289 (N_1289,N_1113,In_1536);
and U1290 (N_1290,In_1859,N_668);
nor U1291 (N_1291,In_388,In_579);
and U1292 (N_1292,N_866,N_806);
nand U1293 (N_1293,N_639,N_836);
nand U1294 (N_1294,In_630,N_808);
nand U1295 (N_1295,N_1107,In_2262);
xor U1296 (N_1296,N_790,N_923);
or U1297 (N_1297,In_618,In_96);
nand U1298 (N_1298,N_492,N_983);
or U1299 (N_1299,In_456,N_703);
or U1300 (N_1300,In_2152,N_648);
xnor U1301 (N_1301,In_1597,In_1305);
or U1302 (N_1302,In_861,N_1155);
and U1303 (N_1303,In_486,N_661);
nand U1304 (N_1304,In_678,N_889);
and U1305 (N_1305,In_1113,N_911);
nand U1306 (N_1306,N_294,N_942);
xor U1307 (N_1307,N_1085,N_814);
nand U1308 (N_1308,N_164,N_1064);
nor U1309 (N_1309,N_669,In_1024);
nand U1310 (N_1310,In_548,N_118);
nand U1311 (N_1311,N_941,In_196);
and U1312 (N_1312,N_882,N_732);
nor U1313 (N_1313,N_113,N_834);
nand U1314 (N_1314,In_1414,In_530);
or U1315 (N_1315,In_1571,N_839);
and U1316 (N_1316,N_671,In_870);
and U1317 (N_1317,N_657,N_734);
nor U1318 (N_1318,In_1593,N_493);
xor U1319 (N_1319,In_841,N_1181);
nor U1320 (N_1320,N_1041,In_26);
nand U1321 (N_1321,In_25,N_350);
nor U1322 (N_1322,N_127,N_28);
or U1323 (N_1323,N_237,N_130);
or U1324 (N_1324,In_974,N_898);
nand U1325 (N_1325,N_1109,N_797);
nand U1326 (N_1326,In_1292,N_781);
and U1327 (N_1327,N_841,N_1115);
or U1328 (N_1328,N_1100,In_1852);
nor U1329 (N_1329,In_834,N_16);
or U1330 (N_1330,N_874,In_1740);
or U1331 (N_1331,In_1538,N_256);
nor U1332 (N_1332,In_1123,N_1171);
or U1333 (N_1333,In_1883,N_1013);
nor U1334 (N_1334,In_791,N_1132);
xnor U1335 (N_1335,N_934,N_1143);
or U1336 (N_1336,N_801,In_2118);
or U1337 (N_1337,In_917,N_937);
nand U1338 (N_1338,N_1178,N_659);
xor U1339 (N_1339,In_1918,In_608);
and U1340 (N_1340,N_1182,In_1801);
xor U1341 (N_1341,N_625,N_602);
nor U1342 (N_1342,N_1068,N_862);
or U1343 (N_1343,N_631,N_644);
or U1344 (N_1344,N_1120,N_982);
or U1345 (N_1345,In_2200,N_1147);
nor U1346 (N_1346,In_1071,In_777);
nor U1347 (N_1347,N_1158,N_1062);
or U1348 (N_1348,In_502,N_1057);
and U1349 (N_1349,N_1227,N_566);
nor U1350 (N_1350,N_924,N_1);
nand U1351 (N_1351,In_1613,In_2181);
nor U1352 (N_1352,N_361,In_369);
or U1353 (N_1353,N_1196,In_338);
nand U1354 (N_1354,In_2003,N_897);
nand U1355 (N_1355,N_1172,N_1209);
or U1356 (N_1356,N_1129,N_134);
nand U1357 (N_1357,N_778,N_662);
nor U1358 (N_1358,N_945,N_1116);
nand U1359 (N_1359,In_673,In_1460);
and U1360 (N_1360,In_2208,In_2257);
and U1361 (N_1361,In_1877,N_858);
nor U1362 (N_1362,In_649,In_303);
nor U1363 (N_1363,In_1318,N_424);
nand U1364 (N_1364,N_1212,In_234);
and U1365 (N_1365,In_570,N_235);
and U1366 (N_1366,In_1829,N_1038);
nand U1367 (N_1367,N_998,N_787);
nand U1368 (N_1368,N_857,In_64);
xor U1369 (N_1369,N_718,N_1229);
nor U1370 (N_1370,N_561,N_652);
or U1371 (N_1371,N_341,N_1130);
nor U1372 (N_1372,N_912,In_643);
nand U1373 (N_1373,In_2123,N_637);
nor U1374 (N_1374,N_1162,In_1329);
nand U1375 (N_1375,N_677,N_670);
or U1376 (N_1376,In_1288,In_1767);
nor U1377 (N_1377,N_633,N_171);
nand U1378 (N_1378,N_673,N_1066);
nand U1379 (N_1379,N_1069,N_1067);
nand U1380 (N_1380,N_827,N_651);
or U1381 (N_1381,In_547,N_838);
xnor U1382 (N_1382,N_1046,N_1106);
or U1383 (N_1383,In_1294,In_1009);
nand U1384 (N_1384,N_1032,In_1949);
xor U1385 (N_1385,N_1202,In_1669);
or U1386 (N_1386,N_421,N_780);
xnor U1387 (N_1387,N_1170,N_57);
xor U1388 (N_1388,N_756,N_950);
nand U1389 (N_1389,N_880,In_2455);
and U1390 (N_1390,In_779,N_8);
nor U1391 (N_1391,N_992,N_1002);
or U1392 (N_1392,N_968,In_2475);
and U1393 (N_1393,N_1198,N_1012);
xnor U1394 (N_1394,N_1025,N_1160);
or U1395 (N_1395,N_1189,In_1764);
nand U1396 (N_1396,N_77,N_627);
nor U1397 (N_1397,In_1635,In_1957);
xor U1398 (N_1398,N_832,N_569);
xor U1399 (N_1399,In_1950,N_812);
nor U1400 (N_1400,N_794,In_747);
or U1401 (N_1401,N_41,In_1406);
nor U1402 (N_1402,In_42,N_796);
nand U1403 (N_1403,N_212,In_872);
nand U1404 (N_1404,In_972,N_467);
nand U1405 (N_1405,N_1033,N_1077);
nor U1406 (N_1406,N_713,N_885);
xnor U1407 (N_1407,In_2055,N_763);
nand U1408 (N_1408,In_2431,N_1114);
or U1409 (N_1409,In_812,N_1099);
and U1410 (N_1410,In_563,N_773);
and U1411 (N_1411,N_655,N_180);
and U1412 (N_1412,In_258,In_383);
and U1413 (N_1413,N_686,In_1013);
nand U1414 (N_1414,N_1029,In_1745);
and U1415 (N_1415,N_1179,N_961);
nand U1416 (N_1416,N_80,N_917);
or U1417 (N_1417,N_1183,N_1020);
nand U1418 (N_1418,N_1059,N_438);
or U1419 (N_1419,N_744,In_2275);
nor U1420 (N_1420,In_2356,N_1234);
or U1421 (N_1421,In_334,N_1011);
nor U1422 (N_1422,In_1385,In_1148);
or U1423 (N_1423,In_952,N_242);
xnor U1424 (N_1424,In_2302,N_1236);
and U1425 (N_1425,In_218,In_632);
nor U1426 (N_1426,In_1199,N_225);
xor U1427 (N_1427,In_1170,N_1119);
and U1428 (N_1428,N_755,N_634);
nand U1429 (N_1429,In_2029,In_293);
xor U1430 (N_1430,N_772,N_658);
nor U1431 (N_1431,N_167,In_1584);
and U1432 (N_1432,N_893,N_1190);
or U1433 (N_1433,N_516,N_1037);
nor U1434 (N_1434,N_736,N_690);
nand U1435 (N_1435,In_1568,N_986);
or U1436 (N_1436,In_1915,In_2495);
nand U1437 (N_1437,N_1026,N_1221);
nor U1438 (N_1438,N_1203,N_1122);
xnor U1439 (N_1439,N_1127,In_414);
xor U1440 (N_1440,N_37,N_884);
nand U1441 (N_1441,N_666,N_1015);
xnor U1442 (N_1442,N_776,N_1136);
nor U1443 (N_1443,N_363,In_327);
xnor U1444 (N_1444,N_463,In_549);
nor U1445 (N_1445,N_291,N_65);
nand U1446 (N_1446,N_855,In_2363);
nand U1447 (N_1447,In_2174,In_635);
nand U1448 (N_1448,In_1186,In_1795);
nand U1449 (N_1449,N_608,N_218);
nor U1450 (N_1450,N_840,N_193);
nor U1451 (N_1451,N_626,In_901);
and U1452 (N_1452,In_2065,In_1664);
xnor U1453 (N_1453,N_498,In_1106);
nand U1454 (N_1454,N_1249,N_1177);
or U1455 (N_1455,N_354,N_741);
or U1456 (N_1456,N_488,N_770);
xnor U1457 (N_1457,N_1246,In_1592);
or U1458 (N_1458,In_1677,N_67);
nor U1459 (N_1459,In_1118,N_767);
xor U1460 (N_1460,N_725,In_1500);
and U1461 (N_1461,In_2467,In_810);
or U1462 (N_1462,In_2468,In_1312);
and U1463 (N_1463,N_753,N_1175);
xnor U1464 (N_1464,N_845,N_972);
and U1465 (N_1465,N_1180,In_1653);
and U1466 (N_1466,N_469,In_559);
and U1467 (N_1467,N_1081,N_869);
or U1468 (N_1468,N_846,N_1006);
and U1469 (N_1469,N_1123,N_829);
nor U1470 (N_1470,N_1240,N_870);
nand U1471 (N_1471,N_837,N_1096);
or U1472 (N_1472,In_569,In_395);
or U1473 (N_1473,N_1086,In_989);
or U1474 (N_1474,In_2061,N_903);
nor U1475 (N_1475,In_805,N_985);
and U1476 (N_1476,N_1091,In_243);
and U1477 (N_1477,In_1058,N_696);
or U1478 (N_1478,N_612,N_980);
or U1479 (N_1479,In_2407,In_1203);
nand U1480 (N_1480,In_2070,N_642);
nor U1481 (N_1481,N_957,N_485);
or U1482 (N_1482,N_14,N_854);
xor U1483 (N_1483,In_528,N_377);
nand U1484 (N_1484,In_1567,N_1187);
or U1485 (N_1485,N_567,In_1867);
and U1486 (N_1486,N_1241,In_697);
and U1487 (N_1487,In_489,N_813);
xor U1488 (N_1488,In_717,In_597);
or U1489 (N_1489,N_920,In_2349);
and U1490 (N_1490,N_758,N_987);
nor U1491 (N_1491,N_1042,In_1486);
nor U1492 (N_1492,N_1161,In_2026);
nand U1493 (N_1493,In_1176,N_699);
xor U1494 (N_1494,In_2446,N_29);
or U1495 (N_1495,In_15,N_1010);
or U1496 (N_1496,N_848,N_1083);
and U1497 (N_1497,In_14,In_59);
nor U1498 (N_1498,In_1995,N_1076);
xor U1499 (N_1499,In_957,N_597);
xor U1500 (N_1500,In_265,N_989);
xnor U1501 (N_1501,N_274,N_737);
xnor U1502 (N_1502,N_844,N_958);
xnor U1503 (N_1503,N_688,N_1007);
xnor U1504 (N_1504,N_936,In_2114);
nor U1505 (N_1505,N_553,N_1142);
xnor U1506 (N_1506,N_654,In_1864);
nor U1507 (N_1507,In_931,N_628);
and U1508 (N_1508,In_1346,N_1167);
nand U1509 (N_1509,In_1340,N_804);
nor U1510 (N_1510,N_679,In_2456);
nand U1511 (N_1511,In_2412,In_2177);
nand U1512 (N_1512,N_940,In_198);
nand U1513 (N_1513,In_567,N_1016);
nand U1514 (N_1514,N_842,N_66);
nand U1515 (N_1515,In_341,N_1201);
nand U1516 (N_1516,N_721,N_1075);
and U1517 (N_1517,N_210,N_1048);
and U1518 (N_1518,N_95,N_791);
xnor U1519 (N_1519,In_862,In_2149);
or U1520 (N_1520,In_1881,N_1163);
nand U1521 (N_1521,N_751,N_960);
nand U1522 (N_1522,In_1821,N_1028);
nand U1523 (N_1523,In_33,In_1258);
nor U1524 (N_1524,N_706,In_1046);
nand U1525 (N_1525,N_782,N_710);
xnor U1526 (N_1526,N_397,N_527);
and U1527 (N_1527,N_1153,In_2430);
nor U1528 (N_1528,N_300,In_1075);
or U1529 (N_1529,In_2435,N_1230);
and U1530 (N_1530,N_823,N_1073);
nand U1531 (N_1531,In_1581,N_785);
xnor U1532 (N_1532,N_405,N_521);
nor U1533 (N_1533,N_629,N_977);
or U1534 (N_1534,N_1072,N_1144);
nand U1535 (N_1535,In_1225,In_793);
nor U1536 (N_1536,N_711,N_1087);
xor U1537 (N_1537,In_2169,In_938);
nand U1538 (N_1538,N_1118,N_1049);
nand U1539 (N_1539,N_340,N_364);
nand U1540 (N_1540,N_248,N_1031);
nor U1541 (N_1541,N_1018,In_822);
xor U1542 (N_1542,N_1245,N_963);
nor U1543 (N_1543,N_799,N_410);
and U1544 (N_1544,N_100,N_531);
nand U1545 (N_1545,N_358,In_2234);
nor U1546 (N_1546,In_1119,N_973);
and U1547 (N_1547,In_2090,N_453);
xor U1548 (N_1548,In_2403,N_680);
nand U1549 (N_1549,In_1381,N_724);
xnor U1550 (N_1550,In_1467,N_465);
nand U1551 (N_1551,In_1742,N_1117);
nor U1552 (N_1552,In_1618,N_872);
or U1553 (N_1553,N_232,N_678);
nand U1554 (N_1554,In_814,N_714);
or U1555 (N_1555,N_278,N_1009);
nor U1556 (N_1556,N_689,N_831);
or U1557 (N_1557,N_727,N_826);
and U1558 (N_1558,In_471,In_379);
or U1559 (N_1559,N_904,In_905);
and U1560 (N_1560,N_1195,N_1017);
or U1561 (N_1561,In_88,N_72);
nor U1562 (N_1562,N_938,In_84);
or U1563 (N_1563,N_850,N_800);
and U1564 (N_1564,In_1979,In_1803);
xor U1565 (N_1565,In_1728,N_1019);
nor U1566 (N_1566,N_777,In_1451);
or U1567 (N_1567,N_811,N_789);
xnor U1568 (N_1568,N_1174,N_783);
xnor U1569 (N_1569,In_344,In_300);
nand U1570 (N_1570,N_307,N_1121);
and U1571 (N_1571,In_321,N_997);
and U1572 (N_1572,In_514,N_388);
nor U1573 (N_1573,N_547,N_1200);
and U1574 (N_1574,N_1125,N_1135);
xnor U1575 (N_1575,N_746,N_909);
and U1576 (N_1576,In_1487,In_2290);
and U1577 (N_1577,N_694,N_798);
or U1578 (N_1578,In_1369,N_932);
xor U1579 (N_1579,N_1080,In_1898);
xnor U1580 (N_1580,N_342,In_2453);
or U1581 (N_1581,In_922,N_971);
and U1582 (N_1582,In_1654,N_745);
nand U1583 (N_1583,N_552,In_668);
or U1584 (N_1584,In_97,N_104);
nand U1585 (N_1585,N_726,N_398);
nand U1586 (N_1586,In_1458,N_788);
xnor U1587 (N_1587,N_843,In_1991);
and U1588 (N_1588,In_7,N_1133);
nand U1589 (N_1589,In_1129,N_1131);
nor U1590 (N_1590,N_692,In_1614);
or U1591 (N_1591,In_925,N_380);
xnor U1592 (N_1592,In_2156,N_895);
xnor U1593 (N_1593,In_2369,In_2394);
xnor U1594 (N_1594,N_422,In_1612);
xnor U1595 (N_1595,N_131,N_1111);
or U1596 (N_1596,N_649,N_859);
xor U1597 (N_1597,N_160,In_2042);
or U1598 (N_1598,In_113,N_1084);
nand U1599 (N_1599,N_60,N_1207);
and U1600 (N_1600,N_1093,N_660);
nor U1601 (N_1601,N_1055,In_1805);
and U1602 (N_1602,N_640,N_1244);
or U1603 (N_1603,N_868,N_1138);
and U1604 (N_1604,In_1260,N_1151);
nand U1605 (N_1605,N_1110,N_856);
nor U1606 (N_1606,In_1532,N_748);
and U1607 (N_1607,In_1594,N_284);
xor U1608 (N_1608,N_931,In_79);
and U1609 (N_1609,N_1173,N_959);
nor U1610 (N_1610,N_1097,N_890);
and U1611 (N_1611,In_1711,N_771);
nor U1612 (N_1612,N_1226,N_1184);
or U1613 (N_1613,N_881,N_583);
and U1614 (N_1614,In_724,N_873);
or U1615 (N_1615,N_1168,N_1235);
nand U1616 (N_1616,N_446,In_381);
xnor U1617 (N_1617,N_1063,N_792);
and U1618 (N_1618,N_1050,N_1079);
and U1619 (N_1619,In_382,In_2068);
nand U1620 (N_1620,N_1108,N_922);
or U1621 (N_1621,N_1157,N_990);
and U1622 (N_1622,In_695,N_538);
and U1623 (N_1623,In_743,N_878);
or U1624 (N_1624,In_1722,In_1178);
nor U1625 (N_1625,N_517,N_426);
nor U1626 (N_1626,In_2119,In_2304);
and U1627 (N_1627,N_886,N_1134);
nor U1628 (N_1628,N_181,N_828);
xnor U1629 (N_1629,N_596,N_759);
and U1630 (N_1630,N_1214,N_348);
or U1631 (N_1631,N_191,In_2488);
nor U1632 (N_1632,In_312,In_1147);
and U1633 (N_1633,In_1477,N_1021);
or U1634 (N_1634,N_701,N_853);
or U1635 (N_1635,In_845,In_532);
or U1636 (N_1636,In_1550,In_129);
or U1637 (N_1637,In_1749,N_715);
and U1638 (N_1638,N_9,N_333);
and U1639 (N_1639,N_1223,N_1169);
nand U1640 (N_1640,N_409,N_764);
and U1641 (N_1641,N_1140,N_691);
nor U1642 (N_1642,In_1399,N_1217);
xnor U1643 (N_1643,N_784,N_664);
or U1644 (N_1644,N_667,N_603);
xor U1645 (N_1645,N_871,N_879);
and U1646 (N_1646,N_385,In_1857);
and U1647 (N_1647,In_435,In_644);
nand U1648 (N_1648,N_442,In_725);
or U1649 (N_1649,In_733,In_544);
nor U1650 (N_1650,N_951,N_676);
and U1651 (N_1651,In_2242,N_1092);
nand U1652 (N_1652,N_847,N_647);
xor U1653 (N_1653,In_2376,N_1224);
and U1654 (N_1654,N_896,N_621);
nor U1655 (N_1655,N_1065,N_645);
nand U1656 (N_1656,In_1510,N_311);
xnor U1657 (N_1657,In_883,N_490);
and U1658 (N_1658,N_1124,N_1154);
nor U1659 (N_1659,N_913,N_712);
and U1660 (N_1660,N_991,N_1248);
or U1661 (N_1661,In_372,In_261);
or U1662 (N_1662,N_1088,In_601);
xnor U1663 (N_1663,N_1210,N_124);
or U1664 (N_1664,N_863,N_818);
and U1665 (N_1665,N_1034,N_1148);
xor U1666 (N_1666,In_798,N_1102);
xnor U1667 (N_1667,In_2337,In_1093);
and U1668 (N_1668,In_2280,N_1208);
xnor U1669 (N_1669,N_779,N_1247);
nand U1670 (N_1670,N_967,N_577);
nor U1671 (N_1671,In_1348,N_956);
and U1672 (N_1672,In_1828,N_247);
or U1673 (N_1673,In_241,In_166);
nand U1674 (N_1674,N_976,N_1228);
nand U1675 (N_1675,N_643,N_952);
xor U1676 (N_1676,In_399,N_1089);
xor U1677 (N_1677,N_1233,N_786);
and U1678 (N_1678,N_1090,N_665);
nand U1679 (N_1679,N_1192,In_1938);
or U1680 (N_1680,N_1082,N_852);
and U1681 (N_1681,N_955,In_1583);
nor U1682 (N_1682,In_1403,In_762);
and U1683 (N_1683,N_946,N_1152);
or U1684 (N_1684,N_329,N_108);
or U1685 (N_1685,N_1213,N_301);
xor U1686 (N_1686,N_21,N_1243);
nor U1687 (N_1687,In_816,N_137);
nand U1688 (N_1688,N_508,N_636);
and U1689 (N_1689,In_1542,N_1232);
or U1690 (N_1690,In_930,N_925);
nor U1691 (N_1691,N_775,N_953);
and U1692 (N_1692,N_1001,N_30);
nand U1693 (N_1693,In_222,N_1039);
xnor U1694 (N_1694,N_768,N_641);
nand U1695 (N_1695,In_1861,In_244);
and U1696 (N_1696,N_757,N_557);
or U1697 (N_1697,N_1051,N_64);
and U1698 (N_1698,N_835,N_906);
nor U1699 (N_1699,N_749,N_565);
or U1700 (N_1700,In_2170,N_901);
nand U1701 (N_1701,In_869,In_1190);
or U1702 (N_1702,N_305,In_2462);
and U1703 (N_1703,N_830,N_752);
xnor U1704 (N_1704,N_819,N_996);
nand U1705 (N_1705,N_1211,N_400);
nor U1706 (N_1706,N_1197,In_1347);
and U1707 (N_1707,In_652,In_899);
nand U1708 (N_1708,In_1217,N_203);
nand U1709 (N_1709,In_1887,In_1334);
and U1710 (N_1710,In_1011,N_1218);
or U1711 (N_1711,N_1071,N_705);
and U1712 (N_1712,In_245,N_930);
nor U1713 (N_1713,In_1732,In_776);
or U1714 (N_1714,N_1191,N_675);
nor U1715 (N_1715,N_708,N_697);
xor U1716 (N_1716,N_207,In_2414);
and U1717 (N_1717,N_728,In_2239);
or U1718 (N_1718,N_954,In_158);
nand U1719 (N_1719,In_10,N_326);
nand U1720 (N_1720,N_579,N_263);
xnor U1721 (N_1721,N_178,N_974);
or U1722 (N_1722,N_944,N_432);
and U1723 (N_1723,In_1620,N_150);
nand U1724 (N_1724,N_271,N_86);
and U1725 (N_1725,N_738,In_1572);
xor U1726 (N_1726,N_750,N_1000);
nand U1727 (N_1727,N_197,In_2160);
xor U1728 (N_1728,N_887,N_899);
nand U1729 (N_1729,N_964,N_860);
and U1730 (N_1730,N_1176,In_349);
nand U1731 (N_1731,N_1056,N_638);
xor U1732 (N_1732,N_1194,N_650);
nand U1733 (N_1733,N_888,In_248);
or U1734 (N_1734,N_1149,In_1776);
nand U1735 (N_1735,In_1483,In_2256);
nor U1736 (N_1736,N_337,In_1710);
xnor U1737 (N_1737,N_373,In_387);
and U1738 (N_1738,In_894,N_947);
xor U1739 (N_1739,N_1074,In_1393);
nor U1740 (N_1740,N_51,N_817);
xor U1741 (N_1741,N_1030,N_935);
or U1742 (N_1742,In_707,N_995);
nor U1743 (N_1743,In_510,N_1040);
and U1744 (N_1744,In_1982,N_910);
or U1745 (N_1745,N_154,N_929);
nor U1746 (N_1746,N_1204,N_1164);
nand U1747 (N_1747,N_722,N_1216);
xnor U1748 (N_1748,N_1141,In_1806);
or U1749 (N_1749,In_1179,N_468);
nor U1750 (N_1750,In_2100,N_215);
or U1751 (N_1751,N_1150,In_1383);
and U1752 (N_1752,In_2121,N_656);
nand U1753 (N_1753,N_1101,In_453);
nor U1754 (N_1754,N_1242,N_632);
nor U1755 (N_1755,N_1045,N_1239);
nor U1756 (N_1756,N_390,In_1386);
and U1757 (N_1757,N_793,In_592);
nand U1758 (N_1758,N_474,In_1494);
xor U1759 (N_1759,In_2472,N_672);
or U1760 (N_1760,N_698,N_613);
or U1761 (N_1761,N_1054,In_152);
or U1762 (N_1762,In_2127,N_92);
nor U1763 (N_1763,In_2067,N_449);
nand U1764 (N_1764,In_1471,N_1098);
or U1765 (N_1765,N_709,N_296);
or U1766 (N_1766,In_1962,N_883);
xor U1767 (N_1767,N_816,In_927);
and U1768 (N_1768,N_1061,N_1237);
and U1769 (N_1769,In_620,N_1103);
and U1770 (N_1770,In_2465,N_875);
nand U1771 (N_1771,N_5,N_1146);
and U1772 (N_1772,In_1437,In_1955);
nand U1773 (N_1773,N_480,In_1707);
xnor U1774 (N_1774,N_682,N_56);
or U1775 (N_1775,N_431,In_2345);
and U1776 (N_1776,N_825,N_1035);
and U1777 (N_1777,In_1282,N_876);
nor U1778 (N_1778,N_821,In_1886);
or U1779 (N_1779,N_739,In_1847);
nor U1780 (N_1780,N_1156,N_743);
xor U1781 (N_1781,N_700,N_219);
and U1782 (N_1782,N_760,N_704);
nand U1783 (N_1783,N_683,N_1023);
xor U1784 (N_1784,In_230,N_61);
xnor U1785 (N_1785,N_1004,N_988);
and U1786 (N_1786,N_851,N_927);
nand U1787 (N_1787,N_653,In_1976);
or U1788 (N_1788,N_681,N_754);
xnor U1789 (N_1789,N_1159,N_1058);
and U1790 (N_1790,N_220,N_762);
and U1791 (N_1791,N_387,N_716);
nand U1792 (N_1792,N_702,In_254);
or U1793 (N_1793,N_984,N_537);
nand U1794 (N_1794,N_1199,N_283);
xor U1795 (N_1795,In_150,In_598);
nor U1796 (N_1796,N_918,In_1750);
nand U1797 (N_1797,N_723,N_1225);
xor U1798 (N_1798,N_646,In_2490);
nor U1799 (N_1799,N_128,N_730);
xor U1800 (N_1800,N_695,N_1186);
nor U1801 (N_1801,N_1166,N_919);
and U1802 (N_1802,N_1095,In_583);
xor U1803 (N_1803,N_20,In_1415);
nor U1804 (N_1804,N_1104,N_867);
xnor U1805 (N_1805,N_674,N_1238);
nand U1806 (N_1806,In_410,N_1044);
and U1807 (N_1807,N_575,N_928);
nor U1808 (N_1808,N_1008,N_731);
or U1809 (N_1809,N_663,N_966);
and U1810 (N_1810,In_2198,N_1094);
and U1811 (N_1811,In_1695,N_765);
xor U1812 (N_1812,N_766,N_747);
nor U1813 (N_1813,N_1206,N_445);
nor U1814 (N_1814,N_965,N_595);
xnor U1815 (N_1815,In_797,N_905);
xnor U1816 (N_1816,In_1652,N_822);
and U1817 (N_1817,N_429,N_1188);
xnor U1818 (N_1818,N_35,N_482);
and U1819 (N_1819,N_849,N_975);
and U1820 (N_1820,N_58,N_907);
and U1821 (N_1821,In_2295,In_833);
nand U1822 (N_1822,In_1226,In_478);
nor U1823 (N_1823,N_1027,In_519);
or U1824 (N_1824,N_824,N_122);
nand U1825 (N_1825,N_915,N_916);
xor U1826 (N_1826,N_433,In_0);
nor U1827 (N_1827,In_1182,N_969);
nor U1828 (N_1828,N_1220,N_23);
or U1829 (N_1829,In_68,N_733);
nand U1830 (N_1830,N_902,In_1925);
nor U1831 (N_1831,N_1036,N_1112);
nor U1832 (N_1832,In_587,In_523);
nand U1833 (N_1833,N_1222,In_468);
or U1834 (N_1834,In_45,N_462);
nand U1835 (N_1835,In_80,N_42);
nand U1836 (N_1836,N_502,N_119);
or U1837 (N_1837,In_466,N_805);
nand U1838 (N_1838,N_1105,N_1231);
xnor U1839 (N_1839,N_810,In_2228);
nor U1840 (N_1840,N_413,In_1706);
nor U1841 (N_1841,In_846,In_35);
and U1842 (N_1842,N_635,N_103);
nor U1843 (N_1843,N_864,In_1320);
nor U1844 (N_1844,N_70,N_693);
or U1845 (N_1845,N_979,In_1087);
nand U1846 (N_1846,N_999,In_217);
and U1847 (N_1847,In_2232,N_451);
nor U1848 (N_1848,N_102,N_949);
xnor U1849 (N_1849,N_460,N_1005);
or U1850 (N_1850,In_2007,In_2325);
nor U1851 (N_1851,In_2494,N_1078);
or U1852 (N_1852,In_655,N_470);
xnor U1853 (N_1853,N_981,In_1668);
xnor U1854 (N_1854,N_1047,N_684);
xnor U1855 (N_1855,N_774,N_926);
or U1856 (N_1856,N_504,N_1022);
xnor U1857 (N_1857,N_962,In_1247);
or U1858 (N_1858,N_605,N_630);
or U1859 (N_1859,In_993,N_994);
and U1860 (N_1860,N_286,N_1024);
nand U1861 (N_1861,N_948,N_707);
nor U1862 (N_1862,N_894,N_939);
nand U1863 (N_1863,N_802,In_77);
nor U1864 (N_1864,In_1608,N_943);
or U1865 (N_1865,In_2219,N_740);
and U1866 (N_1866,N_914,In_2089);
and U1867 (N_1867,In_1833,In_2471);
or U1868 (N_1868,In_2479,N_1139);
or U1869 (N_1869,N_720,In_1482);
nor U1870 (N_1870,In_2144,N_865);
and U1871 (N_1871,In_325,In_1556);
nand U1872 (N_1872,N_742,N_1205);
xor U1873 (N_1873,In_990,In_2314);
or U1874 (N_1874,N_933,N_729);
or U1875 (N_1875,N_1316,N_1537);
or U1876 (N_1876,N_1357,N_1533);
xnor U1877 (N_1877,N_1631,N_1842);
xnor U1878 (N_1878,N_1565,N_1776);
nand U1879 (N_1879,N_1477,N_1779);
and U1880 (N_1880,N_1584,N_1841);
xor U1881 (N_1881,N_1784,N_1598);
or U1882 (N_1882,N_1692,N_1723);
or U1883 (N_1883,N_1614,N_1321);
or U1884 (N_1884,N_1564,N_1496);
nand U1885 (N_1885,N_1253,N_1580);
or U1886 (N_1886,N_1857,N_1782);
or U1887 (N_1887,N_1840,N_1536);
nand U1888 (N_1888,N_1299,N_1291);
nor U1889 (N_1889,N_1540,N_1517);
or U1890 (N_1890,N_1510,N_1481);
or U1891 (N_1891,N_1396,N_1870);
nor U1892 (N_1892,N_1759,N_1793);
or U1893 (N_1893,N_1535,N_1399);
xnor U1894 (N_1894,N_1549,N_1874);
xnor U1895 (N_1895,N_1780,N_1669);
nand U1896 (N_1896,N_1625,N_1442);
or U1897 (N_1897,N_1781,N_1376);
or U1898 (N_1898,N_1482,N_1425);
nand U1899 (N_1899,N_1346,N_1377);
and U1900 (N_1900,N_1741,N_1837);
nand U1901 (N_1901,N_1401,N_1498);
nand U1902 (N_1902,N_1457,N_1324);
xor U1903 (N_1903,N_1761,N_1254);
nand U1904 (N_1904,N_1368,N_1635);
and U1905 (N_1905,N_1666,N_1591);
xnor U1906 (N_1906,N_1538,N_1507);
nor U1907 (N_1907,N_1483,N_1774);
xor U1908 (N_1908,N_1455,N_1786);
nor U1909 (N_1909,N_1516,N_1500);
or U1910 (N_1910,N_1819,N_1677);
xnor U1911 (N_1911,N_1742,N_1672);
xnor U1912 (N_1912,N_1756,N_1460);
or U1913 (N_1913,N_1662,N_1532);
or U1914 (N_1914,N_1395,N_1826);
nand U1915 (N_1915,N_1257,N_1812);
and U1916 (N_1916,N_1822,N_1392);
or U1917 (N_1917,N_1380,N_1262);
xnor U1918 (N_1918,N_1655,N_1449);
nand U1919 (N_1919,N_1468,N_1578);
nand U1920 (N_1920,N_1573,N_1852);
nor U1921 (N_1921,N_1526,N_1319);
xor U1922 (N_1922,N_1544,N_1790);
or U1923 (N_1923,N_1271,N_1372);
or U1924 (N_1924,N_1349,N_1588);
nor U1925 (N_1925,N_1367,N_1652);
or U1926 (N_1926,N_1589,N_1845);
and U1927 (N_1927,N_1701,N_1665);
xor U1928 (N_1928,N_1513,N_1465);
nand U1929 (N_1929,N_1716,N_1547);
xor U1930 (N_1930,N_1753,N_1659);
or U1931 (N_1931,N_1452,N_1648);
xor U1932 (N_1932,N_1274,N_1358);
and U1933 (N_1933,N_1270,N_1521);
or U1934 (N_1934,N_1637,N_1329);
nor U1935 (N_1935,N_1379,N_1288);
and U1936 (N_1936,N_1647,N_1417);
and U1937 (N_1937,N_1423,N_1607);
nand U1938 (N_1938,N_1581,N_1502);
nand U1939 (N_1939,N_1304,N_1788);
or U1940 (N_1940,N_1794,N_1369);
nor U1941 (N_1941,N_1767,N_1545);
nand U1942 (N_1942,N_1272,N_1301);
nor U1943 (N_1943,N_1736,N_1599);
or U1944 (N_1944,N_1830,N_1436);
nand U1945 (N_1945,N_1339,N_1527);
and U1946 (N_1946,N_1644,N_1809);
xor U1947 (N_1947,N_1287,N_1518);
nor U1948 (N_1948,N_1471,N_1493);
and U1949 (N_1949,N_1778,N_1338);
or U1950 (N_1950,N_1709,N_1429);
or U1951 (N_1951,N_1832,N_1715);
or U1952 (N_1952,N_1724,N_1863);
nand U1953 (N_1953,N_1649,N_1785);
nand U1954 (N_1954,N_1706,N_1726);
nor U1955 (N_1955,N_1360,N_1622);
and U1956 (N_1956,N_1294,N_1760);
xnor U1957 (N_1957,N_1438,N_1453);
xnor U1958 (N_1958,N_1322,N_1663);
or U1959 (N_1959,N_1735,N_1290);
nand U1960 (N_1960,N_1577,N_1285);
nor U1961 (N_1961,N_1411,N_1310);
nor U1962 (N_1962,N_1266,N_1654);
nor U1963 (N_1963,N_1859,N_1466);
xor U1964 (N_1964,N_1628,N_1464);
xor U1965 (N_1965,N_1683,N_1630);
nor U1966 (N_1966,N_1491,N_1697);
nand U1967 (N_1967,N_1639,N_1678);
and U1968 (N_1968,N_1766,N_1601);
or U1969 (N_1969,N_1501,N_1725);
nand U1970 (N_1970,N_1559,N_1375);
xor U1971 (N_1971,N_1624,N_1612);
or U1972 (N_1972,N_1543,N_1371);
xnor U1973 (N_1973,N_1755,N_1381);
xor U1974 (N_1974,N_1712,N_1770);
or U1975 (N_1975,N_1394,N_1440);
nand U1976 (N_1976,N_1443,N_1326);
or U1977 (N_1977,N_1611,N_1831);
and U1978 (N_1978,N_1676,N_1872);
xnor U1979 (N_1979,N_1408,N_1503);
or U1980 (N_1980,N_1576,N_1562);
or U1981 (N_1981,N_1733,N_1638);
or U1982 (N_1982,N_1490,N_1340);
xor U1983 (N_1983,N_1582,N_1415);
nand U1984 (N_1984,N_1839,N_1480);
or U1985 (N_1985,N_1560,N_1497);
and U1986 (N_1986,N_1439,N_1768);
or U1987 (N_1987,N_1749,N_1388);
xor U1988 (N_1988,N_1795,N_1504);
xnor U1989 (N_1989,N_1426,N_1805);
nand U1990 (N_1990,N_1593,N_1714);
nor U1991 (N_1991,N_1311,N_1556);
and U1992 (N_1992,N_1539,N_1444);
xnor U1993 (N_1993,N_1393,N_1352);
xor U1994 (N_1994,N_1834,N_1296);
nand U1995 (N_1995,N_1844,N_1681);
or U1996 (N_1996,N_1680,N_1259);
nand U1997 (N_1997,N_1846,N_1308);
nand U1998 (N_1998,N_1470,N_1657);
nor U1999 (N_1999,N_1359,N_1670);
or U2000 (N_2000,N_1341,N_1705);
or U2001 (N_2001,N_1345,N_1300);
xor U2002 (N_2002,N_1469,N_1587);
nand U2003 (N_2003,N_1519,N_1667);
nand U2004 (N_2004,N_1553,N_1318);
nand U2005 (N_2005,N_1397,N_1816);
nand U2006 (N_2006,N_1387,N_1428);
nand U2007 (N_2007,N_1806,N_1525);
nor U2008 (N_2008,N_1462,N_1330);
nand U2009 (N_2009,N_1484,N_1263);
nor U2010 (N_2010,N_1277,N_1686);
nand U2011 (N_2011,N_1864,N_1719);
nor U2012 (N_2012,N_1434,N_1658);
nand U2013 (N_2013,N_1685,N_1463);
or U2014 (N_2014,N_1848,N_1608);
nand U2015 (N_2015,N_1374,N_1555);
or U2016 (N_2016,N_1251,N_1302);
xnor U2017 (N_2017,N_1252,N_1298);
xnor U2018 (N_2018,N_1627,N_1492);
nor U2019 (N_2019,N_1574,N_1721);
and U2020 (N_2020,N_1682,N_1378);
nand U2021 (N_2021,N_1604,N_1632);
nor U2022 (N_2022,N_1617,N_1337);
or U2023 (N_2023,N_1868,N_1334);
xnor U2024 (N_2024,N_1810,N_1499);
and U2025 (N_2025,N_1698,N_1646);
or U2026 (N_2026,N_1447,N_1656);
and U2027 (N_2027,N_1430,N_1514);
nor U2028 (N_2028,N_1276,N_1597);
nor U2029 (N_2029,N_1451,N_1403);
and U2030 (N_2030,N_1303,N_1297);
or U2031 (N_2031,N_1282,N_1320);
and U2032 (N_2032,N_1641,N_1554);
xor U2033 (N_2033,N_1413,N_1815);
nand U2034 (N_2034,N_1331,N_1569);
and U2035 (N_2035,N_1813,N_1688);
or U2036 (N_2036,N_1548,N_1590);
xnor U2037 (N_2037,N_1508,N_1406);
nand U2038 (N_2038,N_1441,N_1867);
and U2039 (N_2039,N_1566,N_1747);
xor U2040 (N_2040,N_1472,N_1629);
xnor U2041 (N_2041,N_1487,N_1746);
xnor U2042 (N_2042,N_1636,N_1528);
nand U2043 (N_2043,N_1802,N_1700);
nor U2044 (N_2044,N_1275,N_1823);
nand U2045 (N_2045,N_1347,N_1264);
xor U2046 (N_2046,N_1255,N_1355);
nand U2047 (N_2047,N_1476,N_1718);
or U2048 (N_2048,N_1744,N_1798);
nor U2049 (N_2049,N_1722,N_1595);
and U2050 (N_2050,N_1594,N_1454);
nand U2051 (N_2051,N_1762,N_1505);
nand U2052 (N_2052,N_1281,N_1353);
xor U2053 (N_2053,N_1695,N_1280);
nand U2054 (N_2054,N_1687,N_1422);
xnor U2055 (N_2055,N_1713,N_1350);
nand U2056 (N_2056,N_1534,N_1801);
and U2057 (N_2057,N_1268,N_1745);
nor U2058 (N_2058,N_1383,N_1634);
nor U2059 (N_2059,N_1432,N_1583);
or U2060 (N_2060,N_1783,N_1509);
and U2061 (N_2061,N_1550,N_1871);
nor U2062 (N_2062,N_1354,N_1704);
xnor U2063 (N_2063,N_1585,N_1684);
and U2064 (N_2064,N_1407,N_1856);
or U2065 (N_2065,N_1858,N_1362);
and U2066 (N_2066,N_1603,N_1445);
xnor U2067 (N_2067,N_1551,N_1366);
or U2068 (N_2068,N_1609,N_1279);
nand U2069 (N_2069,N_1833,N_1365);
or U2070 (N_2070,N_1750,N_1356);
or U2071 (N_2071,N_1506,N_1328);
nand U2072 (N_2072,N_1699,N_1344);
or U2073 (N_2073,N_1703,N_1727);
or U2074 (N_2074,N_1313,N_1410);
nand U2075 (N_2075,N_1616,N_1552);
and U2076 (N_2076,N_1619,N_1317);
xor U2077 (N_2077,N_1650,N_1335);
or U2078 (N_2078,N_1694,N_1579);
nor U2079 (N_2079,N_1811,N_1446);
nor U2080 (N_2080,N_1572,N_1799);
nor U2081 (N_2081,N_1416,N_1531);
or U2082 (N_2082,N_1772,N_1702);
nor U2083 (N_2083,N_1382,N_1278);
and U2084 (N_2084,N_1398,N_1620);
and U2085 (N_2085,N_1748,N_1295);
nor U2086 (N_2086,N_1847,N_1691);
nor U2087 (N_2087,N_1307,N_1265);
and U2088 (N_2088,N_1389,N_1789);
and U2089 (N_2089,N_1739,N_1459);
xor U2090 (N_2090,N_1561,N_1474);
and U2091 (N_2091,N_1796,N_1673);
nor U2092 (N_2092,N_1437,N_1558);
nor U2093 (N_2093,N_1289,N_1850);
and U2094 (N_2094,N_1523,N_1390);
nand U2095 (N_2095,N_1803,N_1256);
xor U2096 (N_2096,N_1828,N_1314);
nand U2097 (N_2097,N_1640,N_1763);
xor U2098 (N_2098,N_1419,N_1618);
and U2099 (N_2099,N_1853,N_1386);
and U2100 (N_2100,N_1729,N_1485);
and U2101 (N_2101,N_1524,N_1512);
nand U2102 (N_2102,N_1792,N_1568);
and U2103 (N_2103,N_1570,N_1606);
or U2104 (N_2104,N_1351,N_1851);
xnor U2105 (N_2105,N_1348,N_1814);
nand U2106 (N_2106,N_1414,N_1610);
or U2107 (N_2107,N_1567,N_1520);
and U2108 (N_2108,N_1373,N_1400);
nor U2109 (N_2109,N_1424,N_1653);
and U2110 (N_2110,N_1711,N_1495);
and U2111 (N_2111,N_1511,N_1804);
xor U2112 (N_2112,N_1791,N_1671);
and U2113 (N_2113,N_1849,N_1325);
xor U2114 (N_2114,N_1752,N_1405);
or U2115 (N_2115,N_1777,N_1708);
nand U2116 (N_2116,N_1467,N_1771);
xor U2117 (N_2117,N_1664,N_1651);
and U2118 (N_2118,N_1293,N_1309);
or U2119 (N_2119,N_1494,N_1728);
nor U2120 (N_2120,N_1689,N_1557);
or U2121 (N_2121,N_1738,N_1690);
nor U2122 (N_2122,N_1575,N_1258);
and U2123 (N_2123,N_1861,N_1563);
and U2124 (N_2124,N_1642,N_1626);
xnor U2125 (N_2125,N_1435,N_1458);
xor U2126 (N_2126,N_1261,N_1855);
or U2127 (N_2127,N_1332,N_1333);
and U2128 (N_2128,N_1734,N_1586);
nor U2129 (N_2129,N_1315,N_1284);
nor U2130 (N_2130,N_1343,N_1306);
xor U2131 (N_2131,N_1613,N_1869);
xor U2132 (N_2132,N_1717,N_1621);
nand U2133 (N_2133,N_1836,N_1515);
nand U2134 (N_2134,N_1808,N_1800);
or U2135 (N_2135,N_1409,N_1260);
and U2136 (N_2136,N_1743,N_1286);
nand U2137 (N_2137,N_1843,N_1361);
and U2138 (N_2138,N_1807,N_1862);
and U2139 (N_2139,N_1488,N_1546);
and U2140 (N_2140,N_1530,N_1433);
or U2141 (N_2141,N_1758,N_1764);
nand U2142 (N_2142,N_1775,N_1473);
xnor U2143 (N_2143,N_1448,N_1675);
nor U2144 (N_2144,N_1765,N_1827);
and U2145 (N_2145,N_1456,N_1754);
and U2146 (N_2146,N_1838,N_1820);
and U2147 (N_2147,N_1571,N_1873);
or U2148 (N_2148,N_1707,N_1450);
xor U2149 (N_2149,N_1363,N_1720);
xor U2150 (N_2150,N_1421,N_1825);
nand U2151 (N_2151,N_1327,N_1769);
or U2152 (N_2152,N_1489,N_1693);
and U2153 (N_2153,N_1596,N_1336);
nor U2154 (N_2154,N_1600,N_1829);
nand U2155 (N_2155,N_1865,N_1757);
xor U2156 (N_2156,N_1602,N_1592);
and U2157 (N_2157,N_1732,N_1605);
nand U2158 (N_2158,N_1312,N_1461);
nand U2159 (N_2159,N_1364,N_1821);
and U2160 (N_2160,N_1478,N_1323);
or U2161 (N_2161,N_1679,N_1696);
nand U2162 (N_2162,N_1370,N_1342);
or U2163 (N_2163,N_1740,N_1615);
or U2164 (N_2164,N_1384,N_1305);
xnor U2165 (N_2165,N_1475,N_1660);
nor U2166 (N_2166,N_1385,N_1529);
nand U2167 (N_2167,N_1730,N_1737);
nor U2168 (N_2168,N_1710,N_1751);
or U2169 (N_2169,N_1250,N_1731);
or U2170 (N_2170,N_1402,N_1643);
nand U2171 (N_2171,N_1542,N_1427);
nand U2172 (N_2172,N_1292,N_1404);
xnor U2173 (N_2173,N_1835,N_1645);
or U2174 (N_2174,N_1824,N_1431);
nor U2175 (N_2175,N_1674,N_1773);
and U2176 (N_2176,N_1541,N_1269);
nand U2177 (N_2177,N_1486,N_1668);
or U2178 (N_2178,N_1479,N_1817);
or U2179 (N_2179,N_1418,N_1854);
nor U2180 (N_2180,N_1797,N_1633);
or U2181 (N_2181,N_1818,N_1522);
nand U2182 (N_2182,N_1420,N_1866);
nor U2183 (N_2183,N_1273,N_1623);
and U2184 (N_2184,N_1267,N_1283);
nand U2185 (N_2185,N_1412,N_1860);
xor U2186 (N_2186,N_1661,N_1391);
or U2187 (N_2187,N_1787,N_1361);
nand U2188 (N_2188,N_1270,N_1808);
xor U2189 (N_2189,N_1646,N_1262);
or U2190 (N_2190,N_1363,N_1535);
xnor U2191 (N_2191,N_1820,N_1294);
xor U2192 (N_2192,N_1487,N_1414);
and U2193 (N_2193,N_1398,N_1499);
nor U2194 (N_2194,N_1795,N_1733);
xnor U2195 (N_2195,N_1548,N_1463);
xnor U2196 (N_2196,N_1420,N_1693);
or U2197 (N_2197,N_1544,N_1332);
or U2198 (N_2198,N_1688,N_1441);
nor U2199 (N_2199,N_1647,N_1292);
nor U2200 (N_2200,N_1341,N_1570);
and U2201 (N_2201,N_1593,N_1537);
nand U2202 (N_2202,N_1472,N_1277);
xnor U2203 (N_2203,N_1695,N_1528);
and U2204 (N_2204,N_1415,N_1753);
nor U2205 (N_2205,N_1468,N_1843);
and U2206 (N_2206,N_1841,N_1524);
nor U2207 (N_2207,N_1606,N_1276);
xor U2208 (N_2208,N_1305,N_1593);
and U2209 (N_2209,N_1443,N_1704);
xnor U2210 (N_2210,N_1734,N_1712);
nand U2211 (N_2211,N_1541,N_1400);
nor U2212 (N_2212,N_1324,N_1649);
xnor U2213 (N_2213,N_1576,N_1354);
or U2214 (N_2214,N_1528,N_1250);
nor U2215 (N_2215,N_1446,N_1314);
xor U2216 (N_2216,N_1388,N_1289);
and U2217 (N_2217,N_1311,N_1453);
or U2218 (N_2218,N_1349,N_1727);
xnor U2219 (N_2219,N_1503,N_1849);
xnor U2220 (N_2220,N_1308,N_1686);
or U2221 (N_2221,N_1317,N_1401);
nand U2222 (N_2222,N_1626,N_1394);
and U2223 (N_2223,N_1370,N_1726);
or U2224 (N_2224,N_1493,N_1802);
or U2225 (N_2225,N_1506,N_1371);
nor U2226 (N_2226,N_1864,N_1760);
xnor U2227 (N_2227,N_1535,N_1379);
xnor U2228 (N_2228,N_1698,N_1392);
xnor U2229 (N_2229,N_1790,N_1705);
nand U2230 (N_2230,N_1354,N_1387);
or U2231 (N_2231,N_1838,N_1397);
nand U2232 (N_2232,N_1453,N_1428);
or U2233 (N_2233,N_1725,N_1629);
nand U2234 (N_2234,N_1669,N_1864);
or U2235 (N_2235,N_1365,N_1292);
or U2236 (N_2236,N_1531,N_1824);
and U2237 (N_2237,N_1611,N_1783);
xnor U2238 (N_2238,N_1670,N_1468);
xnor U2239 (N_2239,N_1524,N_1597);
or U2240 (N_2240,N_1525,N_1771);
xnor U2241 (N_2241,N_1673,N_1716);
nor U2242 (N_2242,N_1274,N_1769);
nand U2243 (N_2243,N_1570,N_1346);
xor U2244 (N_2244,N_1543,N_1407);
nand U2245 (N_2245,N_1373,N_1437);
and U2246 (N_2246,N_1635,N_1812);
nand U2247 (N_2247,N_1329,N_1742);
nand U2248 (N_2248,N_1348,N_1806);
and U2249 (N_2249,N_1778,N_1387);
xor U2250 (N_2250,N_1526,N_1766);
or U2251 (N_2251,N_1717,N_1601);
xnor U2252 (N_2252,N_1269,N_1456);
and U2253 (N_2253,N_1619,N_1338);
nand U2254 (N_2254,N_1825,N_1488);
and U2255 (N_2255,N_1849,N_1717);
and U2256 (N_2256,N_1622,N_1325);
nor U2257 (N_2257,N_1854,N_1266);
nor U2258 (N_2258,N_1776,N_1775);
and U2259 (N_2259,N_1641,N_1597);
xor U2260 (N_2260,N_1839,N_1824);
nand U2261 (N_2261,N_1530,N_1538);
and U2262 (N_2262,N_1375,N_1301);
xor U2263 (N_2263,N_1378,N_1828);
nand U2264 (N_2264,N_1485,N_1543);
and U2265 (N_2265,N_1658,N_1459);
or U2266 (N_2266,N_1607,N_1872);
nand U2267 (N_2267,N_1840,N_1473);
and U2268 (N_2268,N_1375,N_1728);
and U2269 (N_2269,N_1482,N_1388);
nor U2270 (N_2270,N_1608,N_1315);
and U2271 (N_2271,N_1459,N_1723);
or U2272 (N_2272,N_1276,N_1474);
xor U2273 (N_2273,N_1317,N_1762);
nor U2274 (N_2274,N_1684,N_1611);
and U2275 (N_2275,N_1750,N_1532);
and U2276 (N_2276,N_1774,N_1591);
nand U2277 (N_2277,N_1839,N_1343);
and U2278 (N_2278,N_1648,N_1339);
nor U2279 (N_2279,N_1625,N_1257);
nor U2280 (N_2280,N_1705,N_1359);
nor U2281 (N_2281,N_1666,N_1647);
xor U2282 (N_2282,N_1589,N_1631);
xnor U2283 (N_2283,N_1462,N_1611);
and U2284 (N_2284,N_1751,N_1836);
xnor U2285 (N_2285,N_1797,N_1749);
nand U2286 (N_2286,N_1647,N_1275);
nor U2287 (N_2287,N_1644,N_1864);
nand U2288 (N_2288,N_1542,N_1789);
nand U2289 (N_2289,N_1378,N_1257);
nand U2290 (N_2290,N_1764,N_1371);
and U2291 (N_2291,N_1581,N_1374);
nand U2292 (N_2292,N_1350,N_1439);
nor U2293 (N_2293,N_1422,N_1353);
xor U2294 (N_2294,N_1844,N_1732);
and U2295 (N_2295,N_1825,N_1717);
nor U2296 (N_2296,N_1506,N_1484);
and U2297 (N_2297,N_1795,N_1670);
or U2298 (N_2298,N_1409,N_1354);
nor U2299 (N_2299,N_1355,N_1493);
xor U2300 (N_2300,N_1378,N_1630);
or U2301 (N_2301,N_1773,N_1593);
or U2302 (N_2302,N_1506,N_1250);
nand U2303 (N_2303,N_1405,N_1845);
and U2304 (N_2304,N_1704,N_1321);
or U2305 (N_2305,N_1819,N_1792);
nand U2306 (N_2306,N_1823,N_1495);
or U2307 (N_2307,N_1272,N_1841);
nor U2308 (N_2308,N_1707,N_1430);
nand U2309 (N_2309,N_1457,N_1412);
or U2310 (N_2310,N_1267,N_1327);
nor U2311 (N_2311,N_1408,N_1784);
nor U2312 (N_2312,N_1417,N_1444);
or U2313 (N_2313,N_1726,N_1711);
and U2314 (N_2314,N_1800,N_1487);
xor U2315 (N_2315,N_1434,N_1348);
and U2316 (N_2316,N_1391,N_1589);
or U2317 (N_2317,N_1338,N_1330);
or U2318 (N_2318,N_1455,N_1797);
nor U2319 (N_2319,N_1792,N_1417);
and U2320 (N_2320,N_1488,N_1849);
xor U2321 (N_2321,N_1639,N_1293);
nand U2322 (N_2322,N_1665,N_1538);
nor U2323 (N_2323,N_1702,N_1411);
nand U2324 (N_2324,N_1863,N_1462);
and U2325 (N_2325,N_1605,N_1698);
and U2326 (N_2326,N_1338,N_1702);
nand U2327 (N_2327,N_1503,N_1487);
and U2328 (N_2328,N_1834,N_1749);
and U2329 (N_2329,N_1546,N_1332);
or U2330 (N_2330,N_1527,N_1718);
xnor U2331 (N_2331,N_1771,N_1628);
nand U2332 (N_2332,N_1765,N_1384);
nand U2333 (N_2333,N_1769,N_1404);
or U2334 (N_2334,N_1256,N_1738);
xnor U2335 (N_2335,N_1357,N_1687);
xnor U2336 (N_2336,N_1277,N_1786);
nor U2337 (N_2337,N_1398,N_1779);
nand U2338 (N_2338,N_1585,N_1809);
nor U2339 (N_2339,N_1840,N_1410);
or U2340 (N_2340,N_1425,N_1722);
xnor U2341 (N_2341,N_1640,N_1472);
nor U2342 (N_2342,N_1350,N_1472);
or U2343 (N_2343,N_1767,N_1724);
nand U2344 (N_2344,N_1761,N_1324);
nand U2345 (N_2345,N_1657,N_1261);
nand U2346 (N_2346,N_1367,N_1299);
nor U2347 (N_2347,N_1808,N_1363);
or U2348 (N_2348,N_1603,N_1705);
nor U2349 (N_2349,N_1472,N_1479);
xor U2350 (N_2350,N_1603,N_1686);
nor U2351 (N_2351,N_1624,N_1759);
nor U2352 (N_2352,N_1507,N_1722);
and U2353 (N_2353,N_1500,N_1792);
nor U2354 (N_2354,N_1511,N_1707);
and U2355 (N_2355,N_1305,N_1492);
xor U2356 (N_2356,N_1596,N_1869);
or U2357 (N_2357,N_1453,N_1363);
nor U2358 (N_2358,N_1413,N_1785);
xnor U2359 (N_2359,N_1593,N_1316);
and U2360 (N_2360,N_1365,N_1418);
xnor U2361 (N_2361,N_1767,N_1841);
and U2362 (N_2362,N_1854,N_1450);
nor U2363 (N_2363,N_1304,N_1489);
nand U2364 (N_2364,N_1637,N_1633);
xnor U2365 (N_2365,N_1440,N_1790);
nand U2366 (N_2366,N_1289,N_1326);
nand U2367 (N_2367,N_1439,N_1635);
and U2368 (N_2368,N_1707,N_1611);
xor U2369 (N_2369,N_1254,N_1644);
xor U2370 (N_2370,N_1595,N_1858);
nand U2371 (N_2371,N_1643,N_1568);
or U2372 (N_2372,N_1258,N_1287);
nor U2373 (N_2373,N_1254,N_1251);
or U2374 (N_2374,N_1619,N_1674);
or U2375 (N_2375,N_1737,N_1630);
or U2376 (N_2376,N_1277,N_1626);
or U2377 (N_2377,N_1782,N_1376);
or U2378 (N_2378,N_1367,N_1718);
nand U2379 (N_2379,N_1587,N_1807);
xor U2380 (N_2380,N_1660,N_1469);
nand U2381 (N_2381,N_1665,N_1568);
and U2382 (N_2382,N_1866,N_1385);
xor U2383 (N_2383,N_1287,N_1268);
or U2384 (N_2384,N_1315,N_1506);
nor U2385 (N_2385,N_1478,N_1622);
xnor U2386 (N_2386,N_1509,N_1396);
or U2387 (N_2387,N_1701,N_1858);
xnor U2388 (N_2388,N_1857,N_1557);
or U2389 (N_2389,N_1815,N_1802);
or U2390 (N_2390,N_1562,N_1702);
nand U2391 (N_2391,N_1296,N_1267);
xnor U2392 (N_2392,N_1600,N_1722);
nor U2393 (N_2393,N_1615,N_1312);
xnor U2394 (N_2394,N_1541,N_1624);
and U2395 (N_2395,N_1791,N_1412);
or U2396 (N_2396,N_1844,N_1851);
nor U2397 (N_2397,N_1566,N_1608);
or U2398 (N_2398,N_1442,N_1708);
xor U2399 (N_2399,N_1531,N_1528);
and U2400 (N_2400,N_1791,N_1727);
xnor U2401 (N_2401,N_1333,N_1732);
xor U2402 (N_2402,N_1453,N_1821);
and U2403 (N_2403,N_1378,N_1259);
nand U2404 (N_2404,N_1611,N_1348);
or U2405 (N_2405,N_1802,N_1386);
and U2406 (N_2406,N_1361,N_1370);
or U2407 (N_2407,N_1752,N_1831);
or U2408 (N_2408,N_1559,N_1851);
nor U2409 (N_2409,N_1853,N_1327);
and U2410 (N_2410,N_1868,N_1320);
or U2411 (N_2411,N_1524,N_1536);
and U2412 (N_2412,N_1474,N_1702);
nand U2413 (N_2413,N_1454,N_1702);
nand U2414 (N_2414,N_1267,N_1704);
xnor U2415 (N_2415,N_1779,N_1306);
nand U2416 (N_2416,N_1632,N_1633);
nand U2417 (N_2417,N_1560,N_1693);
nor U2418 (N_2418,N_1331,N_1855);
nand U2419 (N_2419,N_1616,N_1539);
nand U2420 (N_2420,N_1751,N_1861);
xor U2421 (N_2421,N_1351,N_1731);
nand U2422 (N_2422,N_1620,N_1384);
nand U2423 (N_2423,N_1639,N_1561);
and U2424 (N_2424,N_1558,N_1718);
or U2425 (N_2425,N_1359,N_1332);
or U2426 (N_2426,N_1379,N_1666);
or U2427 (N_2427,N_1557,N_1607);
xor U2428 (N_2428,N_1376,N_1732);
xor U2429 (N_2429,N_1391,N_1852);
nand U2430 (N_2430,N_1450,N_1389);
nand U2431 (N_2431,N_1308,N_1834);
and U2432 (N_2432,N_1474,N_1587);
nor U2433 (N_2433,N_1591,N_1460);
or U2434 (N_2434,N_1353,N_1659);
nor U2435 (N_2435,N_1270,N_1811);
xor U2436 (N_2436,N_1276,N_1838);
nor U2437 (N_2437,N_1769,N_1679);
or U2438 (N_2438,N_1564,N_1696);
xor U2439 (N_2439,N_1673,N_1328);
nor U2440 (N_2440,N_1497,N_1415);
and U2441 (N_2441,N_1397,N_1342);
nand U2442 (N_2442,N_1479,N_1740);
and U2443 (N_2443,N_1626,N_1610);
xor U2444 (N_2444,N_1613,N_1331);
xnor U2445 (N_2445,N_1546,N_1775);
xnor U2446 (N_2446,N_1598,N_1351);
and U2447 (N_2447,N_1664,N_1621);
xnor U2448 (N_2448,N_1499,N_1496);
nor U2449 (N_2449,N_1588,N_1609);
or U2450 (N_2450,N_1845,N_1577);
nor U2451 (N_2451,N_1542,N_1734);
nor U2452 (N_2452,N_1720,N_1656);
xor U2453 (N_2453,N_1589,N_1645);
and U2454 (N_2454,N_1353,N_1872);
xnor U2455 (N_2455,N_1685,N_1735);
xnor U2456 (N_2456,N_1279,N_1472);
nor U2457 (N_2457,N_1623,N_1374);
and U2458 (N_2458,N_1356,N_1847);
and U2459 (N_2459,N_1349,N_1441);
and U2460 (N_2460,N_1600,N_1423);
xor U2461 (N_2461,N_1871,N_1823);
or U2462 (N_2462,N_1367,N_1568);
or U2463 (N_2463,N_1558,N_1523);
or U2464 (N_2464,N_1794,N_1672);
and U2465 (N_2465,N_1288,N_1761);
and U2466 (N_2466,N_1765,N_1497);
xnor U2467 (N_2467,N_1267,N_1414);
nand U2468 (N_2468,N_1362,N_1656);
nor U2469 (N_2469,N_1572,N_1623);
or U2470 (N_2470,N_1397,N_1376);
xor U2471 (N_2471,N_1370,N_1649);
xnor U2472 (N_2472,N_1580,N_1583);
nor U2473 (N_2473,N_1853,N_1709);
or U2474 (N_2474,N_1326,N_1710);
nor U2475 (N_2475,N_1811,N_1570);
or U2476 (N_2476,N_1609,N_1667);
xnor U2477 (N_2477,N_1507,N_1551);
nor U2478 (N_2478,N_1279,N_1825);
and U2479 (N_2479,N_1566,N_1355);
or U2480 (N_2480,N_1543,N_1400);
and U2481 (N_2481,N_1691,N_1489);
or U2482 (N_2482,N_1594,N_1844);
nor U2483 (N_2483,N_1412,N_1765);
xor U2484 (N_2484,N_1782,N_1384);
or U2485 (N_2485,N_1271,N_1296);
nor U2486 (N_2486,N_1382,N_1559);
xnor U2487 (N_2487,N_1293,N_1706);
nand U2488 (N_2488,N_1562,N_1469);
nand U2489 (N_2489,N_1638,N_1322);
nor U2490 (N_2490,N_1688,N_1669);
and U2491 (N_2491,N_1307,N_1728);
nor U2492 (N_2492,N_1551,N_1800);
nand U2493 (N_2493,N_1415,N_1298);
nor U2494 (N_2494,N_1287,N_1871);
nand U2495 (N_2495,N_1497,N_1871);
nand U2496 (N_2496,N_1263,N_1454);
and U2497 (N_2497,N_1712,N_1719);
nor U2498 (N_2498,N_1440,N_1266);
nor U2499 (N_2499,N_1618,N_1872);
nor U2500 (N_2500,N_1938,N_2187);
xnor U2501 (N_2501,N_1956,N_2106);
nor U2502 (N_2502,N_2358,N_1946);
and U2503 (N_2503,N_1981,N_2251);
nor U2504 (N_2504,N_2269,N_2385);
xnor U2505 (N_2505,N_2092,N_2252);
or U2506 (N_2506,N_2102,N_1900);
nor U2507 (N_2507,N_2451,N_2105);
or U2508 (N_2508,N_2420,N_2235);
nor U2509 (N_2509,N_2029,N_2154);
nand U2510 (N_2510,N_2320,N_2403);
or U2511 (N_2511,N_2076,N_2069);
and U2512 (N_2512,N_1961,N_2273);
and U2513 (N_2513,N_2415,N_2381);
nor U2514 (N_2514,N_2421,N_1947);
and U2515 (N_2515,N_2321,N_2088);
xnor U2516 (N_2516,N_2126,N_2429);
nand U2517 (N_2517,N_1970,N_2045);
nand U2518 (N_2518,N_2144,N_2363);
or U2519 (N_2519,N_1892,N_2293);
nor U2520 (N_2520,N_2387,N_2116);
and U2521 (N_2521,N_2449,N_2450);
or U2522 (N_2522,N_1943,N_2139);
nor U2523 (N_2523,N_2177,N_2280);
and U2524 (N_2524,N_1915,N_2444);
or U2525 (N_2525,N_2243,N_1886);
xor U2526 (N_2526,N_1983,N_2165);
or U2527 (N_2527,N_1924,N_2496);
nand U2528 (N_2528,N_2226,N_2111);
xnor U2529 (N_2529,N_2162,N_2422);
or U2530 (N_2530,N_1936,N_2315);
or U2531 (N_2531,N_2404,N_2191);
and U2532 (N_2532,N_2410,N_2434);
or U2533 (N_2533,N_2136,N_2484);
xnor U2534 (N_2534,N_1879,N_2264);
or U2535 (N_2535,N_1906,N_2114);
and U2536 (N_2536,N_2194,N_2219);
nand U2537 (N_2537,N_2331,N_1966);
or U2538 (N_2538,N_2205,N_2272);
and U2539 (N_2539,N_2072,N_2042);
nand U2540 (N_2540,N_2085,N_1905);
or U2541 (N_2541,N_2065,N_2183);
nor U2542 (N_2542,N_2155,N_1888);
xor U2543 (N_2543,N_2201,N_2281);
nand U2544 (N_2544,N_2498,N_2290);
nand U2545 (N_2545,N_2458,N_2365);
or U2546 (N_2546,N_2161,N_2433);
nor U2547 (N_2547,N_2117,N_2148);
nor U2548 (N_2548,N_2466,N_2078);
nand U2549 (N_2549,N_1891,N_2279);
or U2550 (N_2550,N_2068,N_2224);
xor U2551 (N_2551,N_2071,N_2104);
nor U2552 (N_2552,N_2334,N_2423);
xnor U2553 (N_2553,N_2033,N_2371);
nand U2554 (N_2554,N_2412,N_2206);
nor U2555 (N_2555,N_2198,N_2055);
or U2556 (N_2556,N_2200,N_2347);
or U2557 (N_2557,N_2047,N_2238);
and U2558 (N_2558,N_2103,N_1883);
nor U2559 (N_2559,N_2160,N_2081);
and U2560 (N_2560,N_2095,N_1885);
nand U2561 (N_2561,N_2241,N_2390);
xnor U2562 (N_2562,N_2010,N_2374);
nand U2563 (N_2563,N_2419,N_1917);
nand U2564 (N_2564,N_2460,N_2479);
nor U2565 (N_2565,N_2164,N_2312);
xnor U2566 (N_2566,N_2445,N_2378);
or U2567 (N_2567,N_1903,N_1921);
xnor U2568 (N_2568,N_2471,N_1968);
or U2569 (N_2569,N_2020,N_1976);
and U2570 (N_2570,N_2147,N_2207);
or U2571 (N_2571,N_2352,N_2353);
or U2572 (N_2572,N_2212,N_2247);
nand U2573 (N_2573,N_2377,N_2325);
nand U2574 (N_2574,N_2003,N_2488);
or U2575 (N_2575,N_1959,N_2294);
nor U2576 (N_2576,N_1985,N_2487);
and U2577 (N_2577,N_2493,N_1940);
nor U2578 (N_2578,N_2125,N_2196);
and U2579 (N_2579,N_2399,N_1992);
or U2580 (N_2580,N_2351,N_1953);
xnor U2581 (N_2581,N_2425,N_2060);
nand U2582 (N_2582,N_2019,N_2311);
nor U2583 (N_2583,N_1971,N_1988);
nand U2584 (N_2584,N_2338,N_2395);
or U2585 (N_2585,N_1875,N_2394);
or U2586 (N_2586,N_2248,N_2005);
nor U2587 (N_2587,N_2128,N_2140);
xor U2588 (N_2588,N_2250,N_1965);
nor U2589 (N_2589,N_2163,N_2180);
xor U2590 (N_2590,N_2063,N_2316);
and U2591 (N_2591,N_2296,N_2455);
nor U2592 (N_2592,N_1896,N_2375);
or U2593 (N_2593,N_2239,N_1960);
nor U2594 (N_2594,N_1934,N_2392);
nor U2595 (N_2595,N_2052,N_1916);
xor U2596 (N_2596,N_2166,N_2268);
nand U2597 (N_2597,N_2297,N_1951);
xor U2598 (N_2598,N_2237,N_2361);
or U2599 (N_2599,N_2443,N_1930);
and U2600 (N_2600,N_2083,N_2380);
nand U2601 (N_2601,N_2469,N_2211);
nor U2602 (N_2602,N_2027,N_2285);
nand U2603 (N_2603,N_2324,N_2082);
xnor U2604 (N_2604,N_1980,N_2499);
nand U2605 (N_2605,N_2266,N_2044);
and U2606 (N_2606,N_2291,N_2428);
or U2607 (N_2607,N_2061,N_1982);
nor U2608 (N_2608,N_2234,N_2432);
and U2609 (N_2609,N_2232,N_1967);
and U2610 (N_2610,N_2329,N_1909);
xnor U2611 (N_2611,N_2463,N_2064);
nand U2612 (N_2612,N_2303,N_2382);
or U2613 (N_2613,N_2299,N_2464);
xnor U2614 (N_2614,N_2298,N_2202);
nand U2615 (N_2615,N_2473,N_2090);
nor U2616 (N_2616,N_2284,N_2057);
xnor U2617 (N_2617,N_2339,N_2300);
and U2618 (N_2618,N_1958,N_2149);
nor U2619 (N_2619,N_2034,N_2467);
or U2620 (N_2620,N_2195,N_2157);
nor U2621 (N_2621,N_2490,N_2040);
or U2622 (N_2622,N_2492,N_2059);
nor U2623 (N_2623,N_2448,N_2384);
or U2624 (N_2624,N_2388,N_2110);
nor U2625 (N_2625,N_1899,N_2260);
and U2626 (N_2626,N_2062,N_2159);
nor U2627 (N_2627,N_2204,N_2058);
nand U2628 (N_2628,N_2230,N_2413);
or U2629 (N_2629,N_2213,N_2319);
nand U2630 (N_2630,N_2407,N_2454);
xnor U2631 (N_2631,N_2430,N_2357);
and U2632 (N_2632,N_1994,N_2209);
and U2633 (N_2633,N_2309,N_2091);
xnor U2634 (N_2634,N_2015,N_2097);
nand U2635 (N_2635,N_2344,N_1939);
nand U2636 (N_2636,N_2409,N_2222);
or U2637 (N_2637,N_2115,N_1944);
nand U2638 (N_2638,N_2369,N_2295);
and U2639 (N_2639,N_2024,N_2447);
xor U2640 (N_2640,N_2397,N_2168);
xnor U2641 (N_2641,N_2393,N_2427);
nand U2642 (N_2642,N_1895,N_1991);
nand U2643 (N_2643,N_2008,N_2332);
or U2644 (N_2644,N_2002,N_2244);
nand U2645 (N_2645,N_2112,N_2342);
xnor U2646 (N_2646,N_2245,N_1902);
nand U2647 (N_2647,N_2276,N_1890);
or U2648 (N_2648,N_1975,N_2080);
xnor U2649 (N_2649,N_2453,N_1919);
nand U2650 (N_2650,N_1990,N_2262);
or U2651 (N_2651,N_1882,N_2240);
nor U2652 (N_2652,N_2215,N_1926);
and U2653 (N_2653,N_2431,N_2481);
nor U2654 (N_2654,N_2127,N_2121);
or U2655 (N_2655,N_2411,N_2283);
nand U2656 (N_2656,N_2337,N_2383);
nand U2657 (N_2657,N_2118,N_2292);
nand U2658 (N_2658,N_2133,N_1979);
and U2659 (N_2659,N_1893,N_2176);
and U2660 (N_2660,N_2462,N_2152);
nand U2661 (N_2661,N_2025,N_2099);
or U2662 (N_2662,N_2491,N_1998);
xnor U2663 (N_2663,N_2477,N_2486);
xor U2664 (N_2664,N_2253,N_2396);
nand U2665 (N_2665,N_2199,N_2259);
or U2666 (N_2666,N_2098,N_2185);
xor U2667 (N_2667,N_1925,N_2203);
xor U2668 (N_2668,N_2373,N_2016);
or U2669 (N_2669,N_2070,N_2414);
nor U2670 (N_2670,N_2468,N_1952);
nand U2671 (N_2671,N_2093,N_2129);
nand U2672 (N_2672,N_2470,N_2313);
nor U2673 (N_2673,N_2391,N_2485);
xor U2674 (N_2674,N_2326,N_2246);
nand U2675 (N_2675,N_2101,N_2265);
and U2676 (N_2676,N_2330,N_2054);
xnor U2677 (N_2677,N_1901,N_2402);
or U2678 (N_2678,N_2075,N_2441);
nor U2679 (N_2679,N_1932,N_1962);
or U2680 (N_2680,N_2341,N_2188);
nand U2681 (N_2681,N_2023,N_2236);
and U2682 (N_2682,N_2172,N_1914);
xor U2683 (N_2683,N_2231,N_1922);
nand U2684 (N_2684,N_1931,N_2386);
nor U2685 (N_2685,N_2079,N_2474);
nand U2686 (N_2686,N_2398,N_2340);
xnor U2687 (N_2687,N_2077,N_2416);
and U2688 (N_2688,N_1928,N_2014);
nand U2689 (N_2689,N_2327,N_2261);
or U2690 (N_2690,N_2000,N_1929);
or U2691 (N_2691,N_2087,N_1887);
nor U2692 (N_2692,N_2356,N_2305);
and U2693 (N_2693,N_2270,N_2189);
xor U2694 (N_2694,N_2288,N_2084);
and U2695 (N_2695,N_2035,N_2026);
nand U2696 (N_2696,N_2435,N_1977);
and U2697 (N_2697,N_2368,N_2107);
nor U2698 (N_2698,N_2011,N_2495);
and U2699 (N_2699,N_2046,N_2307);
nor U2700 (N_2700,N_2028,N_2457);
nand U2701 (N_2701,N_2184,N_2178);
nor U2702 (N_2702,N_2113,N_2089);
or U2703 (N_2703,N_2401,N_2436);
nor U2704 (N_2704,N_1997,N_2370);
nor U2705 (N_2705,N_2446,N_1923);
nand U2706 (N_2706,N_2036,N_2406);
xor U2707 (N_2707,N_2287,N_2362);
nand U2708 (N_2708,N_2346,N_2349);
nand U2709 (N_2709,N_2173,N_1907);
nor U2710 (N_2710,N_2304,N_2282);
or U2711 (N_2711,N_2169,N_2379);
nor U2712 (N_2712,N_2130,N_2475);
or U2713 (N_2713,N_2355,N_2263);
nor U2714 (N_2714,N_1996,N_1948);
nand U2715 (N_2715,N_2151,N_1969);
nor U2716 (N_2716,N_2459,N_2138);
nor U2717 (N_2717,N_2009,N_2174);
xnor U2718 (N_2718,N_2360,N_2257);
nor U2719 (N_2719,N_2258,N_2233);
nand U2720 (N_2720,N_1918,N_2038);
or U2721 (N_2721,N_1912,N_2367);
nor U2722 (N_2722,N_2094,N_2145);
or U2723 (N_2723,N_2141,N_1884);
nor U2724 (N_2724,N_2175,N_1993);
nor U2725 (N_2725,N_1954,N_1908);
or U2726 (N_2726,N_2120,N_2037);
nor U2727 (N_2727,N_2153,N_2218);
nand U2728 (N_2728,N_2197,N_2190);
nand U2729 (N_2729,N_2056,N_2323);
and U2730 (N_2730,N_1974,N_2408);
xnor U2731 (N_2731,N_2017,N_2494);
nor U2732 (N_2732,N_2074,N_2439);
xnor U2733 (N_2733,N_2437,N_2225);
and U2734 (N_2734,N_2442,N_2376);
nor U2735 (N_2735,N_2333,N_2221);
or U2736 (N_2736,N_1978,N_1904);
xor U2737 (N_2737,N_2220,N_2124);
nor U2738 (N_2738,N_1987,N_2227);
and U2739 (N_2739,N_2004,N_2372);
xnor U2740 (N_2740,N_2228,N_1898);
nand U2741 (N_2741,N_2007,N_2426);
xnor U2742 (N_2742,N_2066,N_2271);
or U2743 (N_2743,N_2167,N_1973);
nand U2744 (N_2744,N_1878,N_2249);
xor U2745 (N_2745,N_2256,N_2278);
nor U2746 (N_2746,N_2400,N_2302);
nor U2747 (N_2747,N_2286,N_1935);
and U2748 (N_2748,N_2006,N_2208);
nor U2749 (N_2749,N_1949,N_2021);
nor U2750 (N_2750,N_2223,N_2354);
and U2751 (N_2751,N_1989,N_2275);
or U2752 (N_2752,N_1933,N_2452);
xnor U2753 (N_2753,N_2182,N_2041);
and U2754 (N_2754,N_2465,N_2336);
or U2755 (N_2755,N_2108,N_1894);
nand U2756 (N_2756,N_1945,N_2193);
or U2757 (N_2757,N_2048,N_1911);
nor U2758 (N_2758,N_2308,N_2100);
or U2759 (N_2759,N_1927,N_2186);
xor U2760 (N_2760,N_2440,N_2229);
or U2761 (N_2761,N_2343,N_2242);
or U2762 (N_2762,N_2031,N_2073);
nand U2763 (N_2763,N_1897,N_2086);
nand U2764 (N_2764,N_2456,N_2348);
or U2765 (N_2765,N_1986,N_1910);
nand U2766 (N_2766,N_2123,N_2314);
nor U2767 (N_2767,N_2067,N_2438);
nor U2768 (N_2768,N_1995,N_2267);
nand U2769 (N_2769,N_2478,N_2350);
nor U2770 (N_2770,N_1920,N_1881);
or U2771 (N_2771,N_2322,N_1937);
nand U2772 (N_2772,N_2461,N_2497);
xnor U2773 (N_2773,N_2032,N_2043);
nand U2774 (N_2774,N_2318,N_2158);
nor U2775 (N_2775,N_1877,N_2310);
nor U2776 (N_2776,N_2472,N_2483);
nor U2777 (N_2777,N_1913,N_1963);
nor U2778 (N_2778,N_2171,N_2192);
xor U2779 (N_2779,N_1950,N_2137);
nor U2780 (N_2780,N_2482,N_2214);
xnor U2781 (N_2781,N_2001,N_2216);
xnor U2782 (N_2782,N_1972,N_2335);
nand U2783 (N_2783,N_2417,N_2150);
or U2784 (N_2784,N_2050,N_2142);
xor U2785 (N_2785,N_2405,N_2018);
nor U2786 (N_2786,N_1889,N_2131);
and U2787 (N_2787,N_1876,N_1984);
nand U2788 (N_2788,N_2418,N_2274);
nand U2789 (N_2789,N_2012,N_2096);
xnor U2790 (N_2790,N_2119,N_2328);
nand U2791 (N_2791,N_2051,N_2217);
xor U2792 (N_2792,N_2039,N_2156);
nand U2793 (N_2793,N_1957,N_2049);
and U2794 (N_2794,N_2022,N_2135);
nor U2795 (N_2795,N_2345,N_2179);
xnor U2796 (N_2796,N_1999,N_2254);
and U2797 (N_2797,N_2122,N_2053);
or U2798 (N_2798,N_2389,N_2476);
or U2799 (N_2799,N_1942,N_2255);
xnor U2800 (N_2800,N_2306,N_2480);
xor U2801 (N_2801,N_2359,N_1880);
xnor U2802 (N_2802,N_2210,N_2181);
nor U2803 (N_2803,N_2317,N_2424);
nor U2804 (N_2804,N_2489,N_2170);
and U2805 (N_2805,N_2277,N_2109);
nor U2806 (N_2806,N_1941,N_2134);
and U2807 (N_2807,N_2013,N_1955);
xor U2808 (N_2808,N_2364,N_2030);
or U2809 (N_2809,N_2143,N_1964);
nand U2810 (N_2810,N_2146,N_2301);
nor U2811 (N_2811,N_2132,N_2366);
nor U2812 (N_2812,N_2289,N_2021);
xor U2813 (N_2813,N_2316,N_2262);
xnor U2814 (N_2814,N_1965,N_2251);
xnor U2815 (N_2815,N_1931,N_2210);
or U2816 (N_2816,N_1924,N_1990);
xor U2817 (N_2817,N_2206,N_1963);
nand U2818 (N_2818,N_2426,N_2420);
and U2819 (N_2819,N_2206,N_2398);
nor U2820 (N_2820,N_2418,N_2455);
nor U2821 (N_2821,N_2298,N_2125);
and U2822 (N_2822,N_1996,N_2094);
xor U2823 (N_2823,N_1965,N_2143);
xnor U2824 (N_2824,N_2459,N_2239);
or U2825 (N_2825,N_2417,N_2447);
xnor U2826 (N_2826,N_2162,N_1919);
nor U2827 (N_2827,N_2187,N_1971);
or U2828 (N_2828,N_2447,N_2341);
nor U2829 (N_2829,N_2383,N_1879);
nand U2830 (N_2830,N_2135,N_2305);
or U2831 (N_2831,N_2425,N_2373);
nand U2832 (N_2832,N_2311,N_1997);
or U2833 (N_2833,N_2472,N_2193);
and U2834 (N_2834,N_2282,N_2052);
xor U2835 (N_2835,N_2150,N_2251);
and U2836 (N_2836,N_2374,N_2183);
and U2837 (N_2837,N_2214,N_2086);
or U2838 (N_2838,N_2430,N_2491);
or U2839 (N_2839,N_2237,N_2442);
nand U2840 (N_2840,N_2324,N_1992);
nor U2841 (N_2841,N_2203,N_2472);
or U2842 (N_2842,N_1931,N_2423);
xnor U2843 (N_2843,N_2421,N_2080);
xor U2844 (N_2844,N_1910,N_2277);
nor U2845 (N_2845,N_1945,N_2494);
nor U2846 (N_2846,N_2320,N_2233);
nor U2847 (N_2847,N_2263,N_2296);
and U2848 (N_2848,N_2002,N_2359);
nor U2849 (N_2849,N_2019,N_1912);
or U2850 (N_2850,N_1967,N_2173);
or U2851 (N_2851,N_2487,N_2361);
or U2852 (N_2852,N_1971,N_2093);
xnor U2853 (N_2853,N_2327,N_2007);
or U2854 (N_2854,N_2013,N_2209);
and U2855 (N_2855,N_2238,N_1989);
nor U2856 (N_2856,N_2406,N_2056);
or U2857 (N_2857,N_2486,N_2439);
or U2858 (N_2858,N_1929,N_2368);
nor U2859 (N_2859,N_2354,N_1882);
xnor U2860 (N_2860,N_2268,N_1917);
or U2861 (N_2861,N_2428,N_1901);
nor U2862 (N_2862,N_2360,N_1970);
nor U2863 (N_2863,N_2131,N_2020);
or U2864 (N_2864,N_2040,N_2476);
xor U2865 (N_2865,N_1933,N_2406);
xor U2866 (N_2866,N_2230,N_2186);
nor U2867 (N_2867,N_2490,N_1937);
nor U2868 (N_2868,N_1956,N_2373);
and U2869 (N_2869,N_2057,N_2117);
and U2870 (N_2870,N_2204,N_2234);
nand U2871 (N_2871,N_2196,N_2361);
nand U2872 (N_2872,N_2380,N_2088);
nor U2873 (N_2873,N_2172,N_2109);
xor U2874 (N_2874,N_2042,N_2198);
nand U2875 (N_2875,N_2077,N_2027);
or U2876 (N_2876,N_2136,N_1904);
or U2877 (N_2877,N_2348,N_2277);
xor U2878 (N_2878,N_2377,N_2493);
nor U2879 (N_2879,N_1971,N_2467);
nand U2880 (N_2880,N_2473,N_2198);
nand U2881 (N_2881,N_2346,N_2398);
or U2882 (N_2882,N_2118,N_2413);
nand U2883 (N_2883,N_2310,N_1964);
xnor U2884 (N_2884,N_2475,N_2440);
or U2885 (N_2885,N_1957,N_2170);
nor U2886 (N_2886,N_2033,N_1896);
nand U2887 (N_2887,N_2466,N_1977);
and U2888 (N_2888,N_2115,N_2108);
and U2889 (N_2889,N_2374,N_2201);
nor U2890 (N_2890,N_2004,N_1955);
and U2891 (N_2891,N_2069,N_2331);
nor U2892 (N_2892,N_2421,N_2035);
xnor U2893 (N_2893,N_2108,N_1901);
nor U2894 (N_2894,N_2438,N_2468);
nor U2895 (N_2895,N_1919,N_2197);
nor U2896 (N_2896,N_2484,N_2400);
and U2897 (N_2897,N_1974,N_2260);
or U2898 (N_2898,N_2007,N_2435);
nor U2899 (N_2899,N_2104,N_2179);
nor U2900 (N_2900,N_1982,N_2461);
and U2901 (N_2901,N_2148,N_2016);
or U2902 (N_2902,N_2074,N_2482);
nand U2903 (N_2903,N_2354,N_1970);
xnor U2904 (N_2904,N_2139,N_2062);
xor U2905 (N_2905,N_2007,N_2233);
nand U2906 (N_2906,N_2314,N_2284);
nor U2907 (N_2907,N_2433,N_2011);
nand U2908 (N_2908,N_2361,N_2376);
or U2909 (N_2909,N_2074,N_2365);
or U2910 (N_2910,N_1991,N_2432);
or U2911 (N_2911,N_2109,N_2405);
and U2912 (N_2912,N_2284,N_2293);
or U2913 (N_2913,N_1988,N_2300);
nor U2914 (N_2914,N_2209,N_2240);
and U2915 (N_2915,N_2211,N_2314);
nor U2916 (N_2916,N_2071,N_2007);
nand U2917 (N_2917,N_1879,N_2074);
or U2918 (N_2918,N_1929,N_2460);
or U2919 (N_2919,N_2185,N_2068);
nand U2920 (N_2920,N_2258,N_2008);
and U2921 (N_2921,N_2486,N_1974);
xor U2922 (N_2922,N_2034,N_1980);
nor U2923 (N_2923,N_2210,N_2366);
and U2924 (N_2924,N_2202,N_2163);
and U2925 (N_2925,N_2031,N_2223);
and U2926 (N_2926,N_2340,N_1885);
nor U2927 (N_2927,N_1959,N_2350);
nor U2928 (N_2928,N_1996,N_1899);
nor U2929 (N_2929,N_2361,N_2362);
nor U2930 (N_2930,N_2058,N_2492);
nor U2931 (N_2931,N_2414,N_2427);
and U2932 (N_2932,N_1919,N_2053);
or U2933 (N_2933,N_2264,N_2105);
nor U2934 (N_2934,N_1878,N_1993);
and U2935 (N_2935,N_2424,N_2104);
nand U2936 (N_2936,N_2499,N_2237);
nand U2937 (N_2937,N_2279,N_2370);
nand U2938 (N_2938,N_2113,N_2461);
or U2939 (N_2939,N_2375,N_2406);
and U2940 (N_2940,N_2048,N_1974);
nand U2941 (N_2941,N_2291,N_2146);
xnor U2942 (N_2942,N_2453,N_2302);
or U2943 (N_2943,N_2145,N_2004);
xnor U2944 (N_2944,N_2408,N_1926);
nor U2945 (N_2945,N_1893,N_2152);
nand U2946 (N_2946,N_2070,N_2497);
and U2947 (N_2947,N_2419,N_2242);
xor U2948 (N_2948,N_2435,N_2309);
and U2949 (N_2949,N_2412,N_1878);
and U2950 (N_2950,N_2097,N_2284);
nand U2951 (N_2951,N_2086,N_2343);
and U2952 (N_2952,N_2116,N_2385);
or U2953 (N_2953,N_2178,N_2035);
nand U2954 (N_2954,N_2430,N_2282);
xor U2955 (N_2955,N_2187,N_2050);
xnor U2956 (N_2956,N_2406,N_2229);
nand U2957 (N_2957,N_2417,N_1995);
and U2958 (N_2958,N_2014,N_2269);
xor U2959 (N_2959,N_2146,N_2440);
and U2960 (N_2960,N_2464,N_2144);
or U2961 (N_2961,N_1900,N_2095);
or U2962 (N_2962,N_2112,N_2141);
xnor U2963 (N_2963,N_2088,N_2423);
xnor U2964 (N_2964,N_2175,N_2299);
and U2965 (N_2965,N_2299,N_2286);
or U2966 (N_2966,N_2130,N_2470);
nor U2967 (N_2967,N_2293,N_2466);
nand U2968 (N_2968,N_2187,N_1890);
xnor U2969 (N_2969,N_2328,N_2463);
nor U2970 (N_2970,N_2406,N_2476);
or U2971 (N_2971,N_1887,N_2016);
xnor U2972 (N_2972,N_2088,N_2446);
nand U2973 (N_2973,N_1915,N_2083);
xnor U2974 (N_2974,N_1934,N_2447);
and U2975 (N_2975,N_2477,N_2025);
or U2976 (N_2976,N_2196,N_2329);
or U2977 (N_2977,N_2360,N_2174);
nor U2978 (N_2978,N_2331,N_1928);
xor U2979 (N_2979,N_1943,N_2070);
or U2980 (N_2980,N_2472,N_2399);
xor U2981 (N_2981,N_2182,N_2071);
or U2982 (N_2982,N_2359,N_2474);
nor U2983 (N_2983,N_1980,N_2043);
and U2984 (N_2984,N_2318,N_2372);
and U2985 (N_2985,N_1955,N_2368);
nor U2986 (N_2986,N_2491,N_1988);
or U2987 (N_2987,N_2395,N_2216);
nand U2988 (N_2988,N_2204,N_1922);
xor U2989 (N_2989,N_2198,N_2216);
or U2990 (N_2990,N_2296,N_1875);
nand U2991 (N_2991,N_1989,N_2067);
xnor U2992 (N_2992,N_2152,N_2154);
nand U2993 (N_2993,N_2134,N_2136);
or U2994 (N_2994,N_2143,N_2176);
nor U2995 (N_2995,N_2245,N_2176);
xnor U2996 (N_2996,N_2212,N_2037);
xnor U2997 (N_2997,N_2410,N_2301);
nand U2998 (N_2998,N_2118,N_2058);
nor U2999 (N_2999,N_2288,N_1998);
nor U3000 (N_3000,N_1924,N_2433);
xnor U3001 (N_3001,N_2449,N_2281);
nor U3002 (N_3002,N_2046,N_2277);
and U3003 (N_3003,N_2303,N_2389);
and U3004 (N_3004,N_2240,N_2290);
or U3005 (N_3005,N_2416,N_2193);
xnor U3006 (N_3006,N_2223,N_2287);
or U3007 (N_3007,N_2495,N_2443);
xor U3008 (N_3008,N_2232,N_2077);
nor U3009 (N_3009,N_2122,N_2036);
nand U3010 (N_3010,N_1930,N_2222);
and U3011 (N_3011,N_2329,N_2296);
nand U3012 (N_3012,N_2092,N_2483);
nor U3013 (N_3013,N_1957,N_2084);
nor U3014 (N_3014,N_1933,N_2108);
nor U3015 (N_3015,N_2194,N_2313);
xor U3016 (N_3016,N_1936,N_2187);
nor U3017 (N_3017,N_2366,N_2032);
and U3018 (N_3018,N_2105,N_1985);
or U3019 (N_3019,N_2437,N_1910);
nand U3020 (N_3020,N_1978,N_2064);
xor U3021 (N_3021,N_2463,N_1878);
xnor U3022 (N_3022,N_2069,N_2362);
nor U3023 (N_3023,N_2252,N_2458);
nand U3024 (N_3024,N_2431,N_2110);
xor U3025 (N_3025,N_2410,N_2244);
nand U3026 (N_3026,N_2052,N_2113);
xnor U3027 (N_3027,N_2352,N_2325);
nand U3028 (N_3028,N_2073,N_2049);
xor U3029 (N_3029,N_2073,N_2202);
and U3030 (N_3030,N_2465,N_2379);
and U3031 (N_3031,N_2159,N_2089);
nand U3032 (N_3032,N_2201,N_2088);
or U3033 (N_3033,N_2204,N_1941);
nand U3034 (N_3034,N_2322,N_2097);
or U3035 (N_3035,N_2109,N_2040);
nor U3036 (N_3036,N_1953,N_2485);
nand U3037 (N_3037,N_1910,N_2300);
nand U3038 (N_3038,N_1891,N_2391);
or U3039 (N_3039,N_2320,N_2261);
xor U3040 (N_3040,N_1878,N_2233);
nor U3041 (N_3041,N_2220,N_2404);
nor U3042 (N_3042,N_2251,N_2304);
nand U3043 (N_3043,N_2118,N_2441);
and U3044 (N_3044,N_2080,N_2427);
nand U3045 (N_3045,N_2294,N_2095);
and U3046 (N_3046,N_1997,N_2476);
and U3047 (N_3047,N_2266,N_2003);
xor U3048 (N_3048,N_2361,N_1967);
nand U3049 (N_3049,N_2236,N_2442);
nand U3050 (N_3050,N_2029,N_1905);
nand U3051 (N_3051,N_2182,N_2391);
and U3052 (N_3052,N_2324,N_2366);
nand U3053 (N_3053,N_2450,N_2290);
nor U3054 (N_3054,N_2236,N_2158);
or U3055 (N_3055,N_2175,N_2071);
nand U3056 (N_3056,N_2397,N_2344);
or U3057 (N_3057,N_2183,N_2151);
nand U3058 (N_3058,N_2009,N_2013);
or U3059 (N_3059,N_1990,N_2220);
nor U3060 (N_3060,N_2474,N_2048);
nor U3061 (N_3061,N_2357,N_1989);
nor U3062 (N_3062,N_1949,N_2254);
nand U3063 (N_3063,N_2443,N_2304);
nand U3064 (N_3064,N_2139,N_2250);
and U3065 (N_3065,N_2352,N_1900);
nor U3066 (N_3066,N_2301,N_2386);
xor U3067 (N_3067,N_2160,N_2336);
xor U3068 (N_3068,N_1948,N_2392);
xor U3069 (N_3069,N_2379,N_2041);
nand U3070 (N_3070,N_2189,N_2396);
or U3071 (N_3071,N_2380,N_2203);
and U3072 (N_3072,N_2189,N_2400);
or U3073 (N_3073,N_1922,N_2100);
nand U3074 (N_3074,N_2481,N_1955);
nand U3075 (N_3075,N_2024,N_2348);
and U3076 (N_3076,N_2284,N_2326);
nor U3077 (N_3077,N_2436,N_2063);
nand U3078 (N_3078,N_1879,N_1904);
nor U3079 (N_3079,N_1947,N_2053);
or U3080 (N_3080,N_2096,N_2480);
or U3081 (N_3081,N_2229,N_2372);
and U3082 (N_3082,N_2260,N_1888);
or U3083 (N_3083,N_2368,N_2192);
or U3084 (N_3084,N_1952,N_2304);
xor U3085 (N_3085,N_1921,N_2033);
and U3086 (N_3086,N_2465,N_1931);
and U3087 (N_3087,N_2259,N_2396);
and U3088 (N_3088,N_2043,N_1902);
xor U3089 (N_3089,N_2033,N_2099);
nor U3090 (N_3090,N_2226,N_2472);
or U3091 (N_3091,N_1974,N_2261);
and U3092 (N_3092,N_2353,N_2120);
xnor U3093 (N_3093,N_2085,N_2189);
and U3094 (N_3094,N_2167,N_2209);
or U3095 (N_3095,N_1884,N_2429);
nor U3096 (N_3096,N_2257,N_2131);
and U3097 (N_3097,N_2430,N_1885);
nand U3098 (N_3098,N_2115,N_2270);
nor U3099 (N_3099,N_2292,N_2137);
and U3100 (N_3100,N_1939,N_1945);
and U3101 (N_3101,N_1987,N_2128);
or U3102 (N_3102,N_2255,N_2339);
xnor U3103 (N_3103,N_2151,N_2242);
nand U3104 (N_3104,N_2109,N_2233);
and U3105 (N_3105,N_2484,N_2200);
nand U3106 (N_3106,N_2410,N_1878);
and U3107 (N_3107,N_2288,N_1934);
or U3108 (N_3108,N_2118,N_1889);
xnor U3109 (N_3109,N_2189,N_2384);
xor U3110 (N_3110,N_2338,N_1961);
and U3111 (N_3111,N_2482,N_2287);
nand U3112 (N_3112,N_2016,N_2045);
nor U3113 (N_3113,N_1927,N_1913);
and U3114 (N_3114,N_2437,N_1928);
nand U3115 (N_3115,N_1992,N_1974);
or U3116 (N_3116,N_1967,N_2179);
and U3117 (N_3117,N_2109,N_2054);
or U3118 (N_3118,N_2036,N_1983);
or U3119 (N_3119,N_2458,N_2339);
xor U3120 (N_3120,N_2006,N_2333);
nor U3121 (N_3121,N_1946,N_2057);
nand U3122 (N_3122,N_2172,N_2414);
or U3123 (N_3123,N_1952,N_2150);
nand U3124 (N_3124,N_2181,N_1889);
nand U3125 (N_3125,N_2526,N_2622);
and U3126 (N_3126,N_2635,N_2788);
and U3127 (N_3127,N_2720,N_2854);
xor U3128 (N_3128,N_2739,N_2549);
nor U3129 (N_3129,N_2920,N_2940);
nor U3130 (N_3130,N_3124,N_2670);
xor U3131 (N_3131,N_3112,N_2891);
or U3132 (N_3132,N_2745,N_2909);
nor U3133 (N_3133,N_2935,N_2693);
or U3134 (N_3134,N_2765,N_2582);
nor U3135 (N_3135,N_2540,N_2984);
and U3136 (N_3136,N_2933,N_2959);
and U3137 (N_3137,N_3013,N_2981);
nor U3138 (N_3138,N_2966,N_2912);
nand U3139 (N_3139,N_2753,N_3017);
or U3140 (N_3140,N_2595,N_2560);
nand U3141 (N_3141,N_3034,N_2599);
nand U3142 (N_3142,N_2881,N_2820);
and U3143 (N_3143,N_2954,N_3093);
and U3144 (N_3144,N_2544,N_2642);
nand U3145 (N_3145,N_2616,N_2849);
or U3146 (N_3146,N_2521,N_2563);
or U3147 (N_3147,N_2871,N_2829);
nand U3148 (N_3148,N_2677,N_2624);
nand U3149 (N_3149,N_3044,N_2839);
and U3150 (N_3150,N_2750,N_2573);
or U3151 (N_3151,N_2887,N_2698);
nor U3152 (N_3152,N_3088,N_2752);
nand U3153 (N_3153,N_2532,N_3082);
nand U3154 (N_3154,N_2749,N_2787);
or U3155 (N_3155,N_2650,N_2922);
xnor U3156 (N_3156,N_2980,N_2971);
nand U3157 (N_3157,N_3030,N_2592);
nor U3158 (N_3158,N_2657,N_2558);
xor U3159 (N_3159,N_2786,N_2627);
or U3160 (N_3160,N_2536,N_2692);
xor U3161 (N_3161,N_2872,N_2575);
xnor U3162 (N_3162,N_3102,N_2856);
or U3163 (N_3163,N_3097,N_3007);
nand U3164 (N_3164,N_2983,N_3103);
and U3165 (N_3165,N_2561,N_2934);
nand U3166 (N_3166,N_2842,N_3109);
and U3167 (N_3167,N_2632,N_2524);
and U3168 (N_3168,N_2664,N_2836);
or U3169 (N_3169,N_2795,N_2837);
xor U3170 (N_3170,N_2918,N_2991);
nor U3171 (N_3171,N_2902,N_2665);
and U3172 (N_3172,N_2628,N_3018);
nor U3173 (N_3173,N_2744,N_2614);
nor U3174 (N_3174,N_2557,N_2611);
and U3175 (N_3175,N_3100,N_2673);
nor U3176 (N_3176,N_2944,N_2525);
nand U3177 (N_3177,N_2522,N_3121);
or U3178 (N_3178,N_2993,N_2732);
and U3179 (N_3179,N_2681,N_2726);
nor U3180 (N_3180,N_2579,N_3117);
xor U3181 (N_3181,N_3006,N_2784);
or U3182 (N_3182,N_2814,N_2571);
and U3183 (N_3183,N_2580,N_2961);
and U3184 (N_3184,N_2974,N_2884);
and U3185 (N_3185,N_3036,N_2979);
or U3186 (N_3186,N_2699,N_3067);
and U3187 (N_3187,N_2858,N_2798);
nand U3188 (N_3188,N_2761,N_2668);
or U3189 (N_3189,N_2669,N_2606);
or U3190 (N_3190,N_3004,N_2867);
nand U3191 (N_3191,N_2683,N_2734);
xor U3192 (N_3192,N_2827,N_3028);
and U3193 (N_3193,N_3065,N_3051);
nand U3194 (N_3194,N_2631,N_2535);
nor U3195 (N_3195,N_3031,N_2904);
nor U3196 (N_3196,N_2537,N_2957);
and U3197 (N_3197,N_3073,N_3054);
or U3198 (N_3198,N_3012,N_2718);
or U3199 (N_3199,N_2586,N_2717);
and U3200 (N_3200,N_2930,N_2691);
nand U3201 (N_3201,N_2850,N_2649);
nor U3202 (N_3202,N_2972,N_2715);
nand U3203 (N_3203,N_2658,N_3086);
or U3204 (N_3204,N_2915,N_2723);
xnor U3205 (N_3205,N_3015,N_2523);
nand U3206 (N_3206,N_2848,N_2770);
and U3207 (N_3207,N_2874,N_2607);
nor U3208 (N_3208,N_3038,N_2682);
nand U3209 (N_3209,N_3009,N_2502);
and U3210 (N_3210,N_3055,N_2948);
xnor U3211 (N_3211,N_2950,N_2680);
nand U3212 (N_3212,N_3053,N_2710);
nand U3213 (N_3213,N_2828,N_2530);
and U3214 (N_3214,N_2851,N_2916);
nor U3215 (N_3215,N_2879,N_2751);
or U3216 (N_3216,N_3063,N_2554);
xor U3217 (N_3217,N_2728,N_2587);
nor U3218 (N_3218,N_3049,N_2647);
or U3219 (N_3219,N_2973,N_2804);
and U3220 (N_3220,N_2946,N_3089);
nand U3221 (N_3221,N_3005,N_2538);
and U3222 (N_3222,N_2953,N_3079);
nor U3223 (N_3223,N_2712,N_2529);
xor U3224 (N_3224,N_2646,N_3090);
or U3225 (N_3225,N_3105,N_2987);
and U3226 (N_3226,N_3002,N_2629);
or U3227 (N_3227,N_2706,N_2731);
nand U3228 (N_3228,N_3113,N_3092);
xor U3229 (N_3229,N_2771,N_2762);
nand U3230 (N_3230,N_3096,N_2548);
xor U3231 (N_3231,N_2782,N_2763);
xnor U3232 (N_3232,N_2951,N_3010);
nand U3233 (N_3233,N_2805,N_3008);
nor U3234 (N_3234,N_2725,N_2927);
or U3235 (N_3235,N_2754,N_2690);
and U3236 (N_3236,N_3021,N_2662);
nor U3237 (N_3237,N_2504,N_2577);
and U3238 (N_3238,N_2671,N_2541);
nor U3239 (N_3239,N_2713,N_2534);
and U3240 (N_3240,N_3057,N_2988);
xnor U3241 (N_3241,N_2510,N_2822);
and U3242 (N_3242,N_2604,N_2511);
xnor U3243 (N_3243,N_3108,N_2823);
or U3244 (N_3244,N_2546,N_3037);
nor U3245 (N_3245,N_2864,N_2703);
nand U3246 (N_3246,N_2896,N_2997);
or U3247 (N_3247,N_2892,N_2711);
nand U3248 (N_3248,N_2766,N_2970);
or U3249 (N_3249,N_2964,N_3024);
nor U3250 (N_3250,N_2833,N_2519);
or U3251 (N_3251,N_3043,N_2889);
or U3252 (N_3252,N_2603,N_2897);
xor U3253 (N_3253,N_2768,N_3061);
nand U3254 (N_3254,N_2746,N_3098);
and U3255 (N_3255,N_2901,N_2808);
and U3256 (N_3256,N_2992,N_3000);
nand U3257 (N_3257,N_2738,N_2947);
and U3258 (N_3258,N_2776,N_2531);
nand U3259 (N_3259,N_2873,N_2694);
and U3260 (N_3260,N_2568,N_2630);
nor U3261 (N_3261,N_3064,N_2716);
and U3262 (N_3262,N_2797,N_2862);
xnor U3263 (N_3263,N_2928,N_2921);
and U3264 (N_3264,N_2855,N_2772);
xor U3265 (N_3265,N_2636,N_2612);
nor U3266 (N_3266,N_3016,N_2885);
nor U3267 (N_3267,N_2996,N_3122);
xor U3268 (N_3268,N_2796,N_2733);
or U3269 (N_3269,N_2569,N_2809);
or U3270 (N_3270,N_2807,N_2617);
or U3271 (N_3271,N_2719,N_3052);
xor U3272 (N_3272,N_3014,N_2623);
xor U3273 (N_3273,N_2644,N_2547);
and U3274 (N_3274,N_2643,N_2594);
or U3275 (N_3275,N_2825,N_2937);
or U3276 (N_3276,N_2767,N_2602);
nor U3277 (N_3277,N_2818,N_2986);
nand U3278 (N_3278,N_2799,N_3025);
or U3279 (N_3279,N_2919,N_2741);
and U3280 (N_3280,N_2955,N_3123);
nand U3281 (N_3281,N_2967,N_2899);
nor U3282 (N_3282,N_2697,N_2663);
xor U3283 (N_3283,N_2824,N_2517);
or U3284 (N_3284,N_2830,N_3120);
and U3285 (N_3285,N_2886,N_2832);
nand U3286 (N_3286,N_2543,N_2625);
nor U3287 (N_3287,N_2562,N_2923);
nand U3288 (N_3288,N_2574,N_3032);
xnor U3289 (N_3289,N_2806,N_2975);
or U3290 (N_3290,N_2672,N_2990);
and U3291 (N_3291,N_2876,N_2666);
xor U3292 (N_3292,N_2679,N_2659);
nor U3293 (N_3293,N_2903,N_2695);
nand U3294 (N_3294,N_3078,N_2515);
or U3295 (N_3295,N_2926,N_3085);
xor U3296 (N_3296,N_2597,N_2736);
nor U3297 (N_3297,N_2709,N_2501);
or U3298 (N_3298,N_3033,N_2593);
nor U3299 (N_3299,N_3041,N_2610);
xnor U3300 (N_3300,N_3106,N_3116);
nor U3301 (N_3301,N_2507,N_2963);
xnor U3302 (N_3302,N_3077,N_2633);
and U3303 (N_3303,N_2952,N_2994);
nor U3304 (N_3304,N_2559,N_2769);
xnor U3305 (N_3305,N_2705,N_2877);
or U3306 (N_3306,N_2760,N_2977);
xnor U3307 (N_3307,N_2840,N_2939);
and U3308 (N_3308,N_2656,N_2591);
xor U3309 (N_3309,N_2865,N_2508);
and U3310 (N_3310,N_2500,N_2801);
xor U3311 (N_3311,N_3001,N_2539);
nand U3312 (N_3312,N_2958,N_2908);
xnor U3313 (N_3313,N_3060,N_2601);
and U3314 (N_3314,N_2512,N_2900);
xnor U3315 (N_3315,N_2949,N_2700);
and U3316 (N_3316,N_2619,N_2914);
and U3317 (N_3317,N_2998,N_2505);
nand U3318 (N_3318,N_2578,N_2590);
and U3319 (N_3319,N_2618,N_2742);
xor U3320 (N_3320,N_2956,N_3094);
nor U3321 (N_3321,N_2868,N_2701);
nor U3322 (N_3322,N_3062,N_2789);
nor U3323 (N_3323,N_2724,N_2686);
xor U3324 (N_3324,N_2565,N_2812);
xnor U3325 (N_3325,N_2834,N_3019);
xnor U3326 (N_3326,N_2678,N_2882);
xnor U3327 (N_3327,N_2727,N_2514);
nor U3328 (N_3328,N_2550,N_3020);
or U3329 (N_3329,N_2552,N_2572);
and U3330 (N_3330,N_2778,N_2518);
and U3331 (N_3331,N_2516,N_2942);
nor U3332 (N_3332,N_2702,N_2925);
xor U3333 (N_3333,N_2924,N_2821);
nor U3334 (N_3334,N_2775,N_3083);
nor U3335 (N_3335,N_2687,N_2689);
and U3336 (N_3336,N_2800,N_2929);
xor U3337 (N_3337,N_3074,N_2995);
and U3338 (N_3338,N_2816,N_2846);
or U3339 (N_3339,N_2652,N_2566);
nand U3340 (N_3340,N_3042,N_2857);
xor U3341 (N_3341,N_3075,N_3023);
xnor U3342 (N_3342,N_2684,N_3068);
nand U3343 (N_3343,N_2564,N_2645);
or U3344 (N_3344,N_2755,N_2513);
nand U3345 (N_3345,N_2581,N_2802);
nand U3346 (N_3346,N_3072,N_3027);
or U3347 (N_3347,N_2729,N_2931);
xnor U3348 (N_3348,N_2576,N_2785);
xnor U3349 (N_3349,N_2609,N_2913);
and U3350 (N_3350,N_2815,N_2835);
xnor U3351 (N_3351,N_3099,N_3087);
and U3352 (N_3352,N_2875,N_2898);
or U3353 (N_3353,N_2570,N_2978);
nor U3354 (N_3354,N_2748,N_2598);
and U3355 (N_3355,N_2863,N_2969);
nand U3356 (N_3356,N_2893,N_2758);
nand U3357 (N_3357,N_3080,N_2811);
nor U3358 (N_3358,N_2621,N_2869);
or U3359 (N_3359,N_2790,N_2932);
nand U3360 (N_3360,N_2708,N_2945);
nor U3361 (N_3361,N_2793,N_3003);
nand U3362 (N_3362,N_2596,N_2743);
or U3363 (N_3363,N_3022,N_2783);
nor U3364 (N_3364,N_2757,N_2792);
xor U3365 (N_3365,N_2620,N_2735);
and U3366 (N_3366,N_2528,N_2870);
nand U3367 (N_3367,N_3026,N_3114);
or U3368 (N_3368,N_3071,N_3119);
and U3369 (N_3369,N_2759,N_2841);
nand U3370 (N_3370,N_2962,N_2791);
nand U3371 (N_3371,N_2740,N_2527);
xnor U3372 (N_3372,N_2813,N_2826);
or U3373 (N_3373,N_3110,N_3029);
nor U3374 (N_3374,N_2883,N_2838);
and U3375 (N_3375,N_2641,N_2817);
and U3376 (N_3376,N_3059,N_3058);
nand U3377 (N_3377,N_2905,N_2675);
nor U3378 (N_3378,N_2696,N_3050);
and U3379 (N_3379,N_2756,N_2730);
xnor U3380 (N_3380,N_2779,N_2588);
nor U3381 (N_3381,N_2637,N_2660);
nand U3382 (N_3382,N_2747,N_2721);
nor U3383 (N_3383,N_2888,N_3095);
or U3384 (N_3384,N_3091,N_2941);
nor U3385 (N_3385,N_2843,N_2844);
or U3386 (N_3386,N_2985,N_2638);
or U3387 (N_3387,N_2640,N_2608);
nand U3388 (N_3388,N_2845,N_2589);
or U3389 (N_3389,N_2674,N_2938);
xnor U3390 (N_3390,N_2910,N_2764);
and U3391 (N_3391,N_3084,N_2583);
xor U3392 (N_3392,N_2960,N_2545);
and U3393 (N_3393,N_2533,N_2906);
and U3394 (N_3394,N_2794,N_2506);
nor U3395 (N_3395,N_2651,N_2989);
or U3396 (N_3396,N_2853,N_2866);
nor U3397 (N_3397,N_2509,N_2847);
nor U3398 (N_3398,N_2707,N_2819);
nor U3399 (N_3399,N_3104,N_3048);
nand U3400 (N_3400,N_2654,N_2626);
nand U3401 (N_3401,N_3070,N_3039);
or U3402 (N_3402,N_2878,N_2917);
xor U3403 (N_3403,N_2803,N_2860);
xor U3404 (N_3404,N_2685,N_2968);
or U3405 (N_3405,N_2936,N_2653);
nand U3406 (N_3406,N_3081,N_2859);
xnor U3407 (N_3407,N_2880,N_3101);
or U3408 (N_3408,N_2890,N_2551);
nand U3409 (N_3409,N_2600,N_3056);
nor U3410 (N_3410,N_2999,N_2503);
or U3411 (N_3411,N_2556,N_2831);
nor U3412 (N_3412,N_2605,N_3047);
nand U3413 (N_3413,N_2667,N_2982);
xor U3414 (N_3414,N_3111,N_2911);
and U3415 (N_3415,N_3069,N_2585);
nand U3416 (N_3416,N_2553,N_2676);
nor U3417 (N_3417,N_2737,N_2555);
nand U3418 (N_3418,N_3118,N_3040);
xnor U3419 (N_3419,N_2894,N_2810);
nor U3420 (N_3420,N_2520,N_3046);
nand U3421 (N_3421,N_3076,N_2722);
nor U3422 (N_3422,N_2774,N_2661);
nand U3423 (N_3423,N_2688,N_2861);
nand U3424 (N_3424,N_2965,N_3045);
or U3425 (N_3425,N_2648,N_2907);
nand U3426 (N_3426,N_2634,N_2895);
nand U3427 (N_3427,N_2852,N_2781);
nor U3428 (N_3428,N_2542,N_2714);
xnor U3429 (N_3429,N_3115,N_2584);
xor U3430 (N_3430,N_2777,N_2655);
xor U3431 (N_3431,N_2615,N_2773);
nand U3432 (N_3432,N_3035,N_2639);
nor U3433 (N_3433,N_3011,N_2567);
and U3434 (N_3434,N_3066,N_2780);
nor U3435 (N_3435,N_3107,N_2976);
nand U3436 (N_3436,N_2943,N_2613);
and U3437 (N_3437,N_2704,N_2567);
xor U3438 (N_3438,N_2523,N_2719);
nor U3439 (N_3439,N_3061,N_3046);
xnor U3440 (N_3440,N_2874,N_2814);
nand U3441 (N_3441,N_3066,N_2646);
nand U3442 (N_3442,N_2956,N_3090);
nand U3443 (N_3443,N_3019,N_2817);
nor U3444 (N_3444,N_2602,N_2851);
nand U3445 (N_3445,N_2532,N_3010);
and U3446 (N_3446,N_2953,N_2682);
or U3447 (N_3447,N_2885,N_2713);
nor U3448 (N_3448,N_3075,N_2907);
or U3449 (N_3449,N_2969,N_3116);
nor U3450 (N_3450,N_2964,N_3100);
nand U3451 (N_3451,N_3108,N_2588);
or U3452 (N_3452,N_2875,N_2573);
nor U3453 (N_3453,N_2662,N_2604);
or U3454 (N_3454,N_2901,N_2812);
nand U3455 (N_3455,N_2712,N_2847);
xor U3456 (N_3456,N_2717,N_2912);
or U3457 (N_3457,N_2862,N_2842);
nand U3458 (N_3458,N_2973,N_2538);
xor U3459 (N_3459,N_2692,N_2981);
nand U3460 (N_3460,N_2658,N_2673);
nand U3461 (N_3461,N_3021,N_2637);
or U3462 (N_3462,N_2624,N_2850);
nor U3463 (N_3463,N_2536,N_2903);
or U3464 (N_3464,N_2549,N_2592);
nand U3465 (N_3465,N_2772,N_2791);
or U3466 (N_3466,N_2683,N_2729);
nand U3467 (N_3467,N_2504,N_2801);
or U3468 (N_3468,N_2840,N_3049);
nor U3469 (N_3469,N_3004,N_3029);
and U3470 (N_3470,N_3012,N_2533);
nand U3471 (N_3471,N_3090,N_2764);
or U3472 (N_3472,N_2764,N_2738);
or U3473 (N_3473,N_2726,N_2751);
nand U3474 (N_3474,N_2937,N_2826);
and U3475 (N_3475,N_2722,N_2542);
and U3476 (N_3476,N_2792,N_3035);
or U3477 (N_3477,N_2939,N_3086);
nor U3478 (N_3478,N_3067,N_2547);
nand U3479 (N_3479,N_2972,N_2773);
and U3480 (N_3480,N_2609,N_2608);
and U3481 (N_3481,N_2501,N_2930);
or U3482 (N_3482,N_2757,N_2818);
or U3483 (N_3483,N_2760,N_2828);
nand U3484 (N_3484,N_2660,N_2648);
and U3485 (N_3485,N_2793,N_2895);
or U3486 (N_3486,N_2885,N_2939);
or U3487 (N_3487,N_2613,N_2757);
and U3488 (N_3488,N_2906,N_2544);
and U3489 (N_3489,N_2694,N_2961);
nor U3490 (N_3490,N_2826,N_2828);
xnor U3491 (N_3491,N_3030,N_2938);
nand U3492 (N_3492,N_2917,N_2946);
or U3493 (N_3493,N_2565,N_2772);
nand U3494 (N_3494,N_2797,N_2854);
xnor U3495 (N_3495,N_2617,N_2658);
xor U3496 (N_3496,N_2874,N_2995);
or U3497 (N_3497,N_2990,N_2547);
nand U3498 (N_3498,N_2863,N_2848);
xor U3499 (N_3499,N_2950,N_2822);
xnor U3500 (N_3500,N_2562,N_2797);
or U3501 (N_3501,N_2872,N_2979);
xnor U3502 (N_3502,N_2528,N_2962);
or U3503 (N_3503,N_2512,N_2649);
or U3504 (N_3504,N_2789,N_2941);
or U3505 (N_3505,N_3086,N_2926);
or U3506 (N_3506,N_3091,N_3008);
nand U3507 (N_3507,N_2534,N_2839);
nand U3508 (N_3508,N_2618,N_3059);
and U3509 (N_3509,N_2619,N_2734);
nor U3510 (N_3510,N_2616,N_2720);
nor U3511 (N_3511,N_3061,N_2739);
and U3512 (N_3512,N_2695,N_2834);
xor U3513 (N_3513,N_2951,N_2779);
and U3514 (N_3514,N_2838,N_2863);
nor U3515 (N_3515,N_3121,N_2796);
and U3516 (N_3516,N_3028,N_2924);
nand U3517 (N_3517,N_3001,N_2588);
or U3518 (N_3518,N_3014,N_2509);
nand U3519 (N_3519,N_2769,N_2517);
nor U3520 (N_3520,N_2918,N_2742);
nor U3521 (N_3521,N_2957,N_3050);
nor U3522 (N_3522,N_2820,N_2955);
or U3523 (N_3523,N_3124,N_2610);
or U3524 (N_3524,N_2687,N_3112);
and U3525 (N_3525,N_2974,N_2635);
or U3526 (N_3526,N_2890,N_2866);
or U3527 (N_3527,N_3034,N_2563);
and U3528 (N_3528,N_2958,N_2676);
nand U3529 (N_3529,N_2585,N_2829);
and U3530 (N_3530,N_2526,N_2775);
nor U3531 (N_3531,N_2642,N_2637);
nand U3532 (N_3532,N_2879,N_2882);
nand U3533 (N_3533,N_2654,N_2505);
and U3534 (N_3534,N_2886,N_2566);
xnor U3535 (N_3535,N_2633,N_2816);
and U3536 (N_3536,N_2611,N_2987);
or U3537 (N_3537,N_3023,N_2893);
and U3538 (N_3538,N_2840,N_2618);
or U3539 (N_3539,N_2528,N_2606);
xor U3540 (N_3540,N_2504,N_2786);
nor U3541 (N_3541,N_2553,N_2755);
xnor U3542 (N_3542,N_2970,N_2524);
nand U3543 (N_3543,N_3109,N_2667);
xor U3544 (N_3544,N_2739,N_2798);
nor U3545 (N_3545,N_2582,N_3006);
nor U3546 (N_3546,N_2800,N_2732);
nor U3547 (N_3547,N_2808,N_3104);
xor U3548 (N_3548,N_3095,N_2852);
xnor U3549 (N_3549,N_2660,N_2911);
nor U3550 (N_3550,N_2830,N_2982);
nand U3551 (N_3551,N_2945,N_2562);
xnor U3552 (N_3552,N_3053,N_2552);
nand U3553 (N_3553,N_2785,N_2805);
nor U3554 (N_3554,N_2534,N_2703);
nor U3555 (N_3555,N_3033,N_2925);
xor U3556 (N_3556,N_2508,N_2579);
or U3557 (N_3557,N_2583,N_2889);
nand U3558 (N_3558,N_2787,N_2843);
nor U3559 (N_3559,N_2635,N_2602);
nor U3560 (N_3560,N_3045,N_2872);
nand U3561 (N_3561,N_2787,N_2748);
nand U3562 (N_3562,N_2528,N_3036);
xnor U3563 (N_3563,N_2731,N_2595);
and U3564 (N_3564,N_3113,N_2799);
nor U3565 (N_3565,N_2763,N_2948);
or U3566 (N_3566,N_2765,N_2603);
and U3567 (N_3567,N_2588,N_3016);
or U3568 (N_3568,N_2686,N_2773);
nand U3569 (N_3569,N_2884,N_2847);
or U3570 (N_3570,N_2967,N_3097);
or U3571 (N_3571,N_3082,N_2662);
xnor U3572 (N_3572,N_3081,N_2829);
or U3573 (N_3573,N_2604,N_3105);
xnor U3574 (N_3574,N_3019,N_2630);
nor U3575 (N_3575,N_2697,N_2513);
nand U3576 (N_3576,N_2558,N_2509);
nand U3577 (N_3577,N_2796,N_2839);
and U3578 (N_3578,N_3086,N_2928);
nor U3579 (N_3579,N_2653,N_2814);
or U3580 (N_3580,N_2669,N_2706);
or U3581 (N_3581,N_2838,N_2974);
nand U3582 (N_3582,N_2545,N_2728);
nor U3583 (N_3583,N_2579,N_2718);
nor U3584 (N_3584,N_2667,N_2697);
and U3585 (N_3585,N_2655,N_2841);
and U3586 (N_3586,N_3036,N_2611);
nand U3587 (N_3587,N_2832,N_3107);
xor U3588 (N_3588,N_2751,N_3085);
nand U3589 (N_3589,N_2634,N_2852);
or U3590 (N_3590,N_2575,N_2559);
xor U3591 (N_3591,N_2843,N_2818);
xor U3592 (N_3592,N_3090,N_2612);
xnor U3593 (N_3593,N_3008,N_2943);
and U3594 (N_3594,N_3032,N_2703);
nand U3595 (N_3595,N_3051,N_2672);
or U3596 (N_3596,N_2720,N_3085);
nand U3597 (N_3597,N_2791,N_3051);
or U3598 (N_3598,N_2849,N_2622);
and U3599 (N_3599,N_2559,N_2747);
and U3600 (N_3600,N_2596,N_2899);
and U3601 (N_3601,N_2689,N_2828);
and U3602 (N_3602,N_2615,N_2941);
nand U3603 (N_3603,N_2833,N_2630);
nand U3604 (N_3604,N_2674,N_2904);
nor U3605 (N_3605,N_2701,N_2592);
nor U3606 (N_3606,N_2625,N_3122);
nand U3607 (N_3607,N_2914,N_2551);
xnor U3608 (N_3608,N_2678,N_2549);
nand U3609 (N_3609,N_2622,N_3055);
nand U3610 (N_3610,N_3105,N_2523);
and U3611 (N_3611,N_2514,N_2925);
or U3612 (N_3612,N_2738,N_2878);
and U3613 (N_3613,N_3011,N_3020);
nor U3614 (N_3614,N_2771,N_3104);
nand U3615 (N_3615,N_2987,N_2732);
or U3616 (N_3616,N_2585,N_2521);
xor U3617 (N_3617,N_2957,N_2825);
and U3618 (N_3618,N_2519,N_3048);
nor U3619 (N_3619,N_2812,N_2669);
nor U3620 (N_3620,N_3087,N_3012);
xnor U3621 (N_3621,N_2512,N_2895);
xor U3622 (N_3622,N_2634,N_2969);
xor U3623 (N_3623,N_2979,N_2949);
nor U3624 (N_3624,N_2934,N_2950);
xor U3625 (N_3625,N_2503,N_2877);
and U3626 (N_3626,N_2685,N_2651);
or U3627 (N_3627,N_2830,N_2584);
nand U3628 (N_3628,N_2807,N_2942);
xnor U3629 (N_3629,N_2527,N_3034);
nor U3630 (N_3630,N_2582,N_2716);
nand U3631 (N_3631,N_2673,N_3033);
nor U3632 (N_3632,N_2989,N_2523);
and U3633 (N_3633,N_2574,N_2691);
or U3634 (N_3634,N_2670,N_2880);
and U3635 (N_3635,N_2583,N_2784);
and U3636 (N_3636,N_2529,N_2651);
and U3637 (N_3637,N_3020,N_3071);
and U3638 (N_3638,N_2954,N_2963);
nor U3639 (N_3639,N_2540,N_2844);
or U3640 (N_3640,N_2681,N_2808);
or U3641 (N_3641,N_3111,N_2956);
and U3642 (N_3642,N_2730,N_2792);
nor U3643 (N_3643,N_2753,N_2990);
nand U3644 (N_3644,N_2510,N_2900);
and U3645 (N_3645,N_2904,N_2637);
xor U3646 (N_3646,N_2798,N_2941);
xnor U3647 (N_3647,N_2714,N_2985);
xor U3648 (N_3648,N_3114,N_2848);
and U3649 (N_3649,N_2696,N_2539);
nor U3650 (N_3650,N_2526,N_2596);
nor U3651 (N_3651,N_2611,N_2508);
xor U3652 (N_3652,N_2625,N_2977);
nand U3653 (N_3653,N_2775,N_2777);
and U3654 (N_3654,N_3104,N_2695);
and U3655 (N_3655,N_3114,N_2704);
and U3656 (N_3656,N_2600,N_3050);
nand U3657 (N_3657,N_3055,N_2580);
nand U3658 (N_3658,N_2680,N_3021);
or U3659 (N_3659,N_2911,N_2800);
and U3660 (N_3660,N_2883,N_3084);
xnor U3661 (N_3661,N_2621,N_2807);
and U3662 (N_3662,N_2770,N_2563);
and U3663 (N_3663,N_3075,N_3026);
nand U3664 (N_3664,N_2666,N_2681);
or U3665 (N_3665,N_3076,N_2858);
and U3666 (N_3666,N_2733,N_2702);
nand U3667 (N_3667,N_2783,N_2526);
xnor U3668 (N_3668,N_3041,N_2856);
nor U3669 (N_3669,N_3043,N_2894);
or U3670 (N_3670,N_2798,N_2989);
nor U3671 (N_3671,N_3041,N_2718);
or U3672 (N_3672,N_2849,N_2673);
xnor U3673 (N_3673,N_3098,N_2788);
xnor U3674 (N_3674,N_2559,N_2861);
or U3675 (N_3675,N_3043,N_2857);
or U3676 (N_3676,N_2760,N_2895);
xor U3677 (N_3677,N_3009,N_2622);
xnor U3678 (N_3678,N_3083,N_3111);
nand U3679 (N_3679,N_2920,N_2513);
or U3680 (N_3680,N_2914,N_2720);
and U3681 (N_3681,N_2938,N_2670);
xnor U3682 (N_3682,N_2651,N_2871);
xnor U3683 (N_3683,N_2884,N_2900);
xnor U3684 (N_3684,N_2933,N_2964);
xnor U3685 (N_3685,N_2791,N_2947);
nor U3686 (N_3686,N_2560,N_3057);
or U3687 (N_3687,N_2832,N_2567);
xnor U3688 (N_3688,N_2882,N_2739);
and U3689 (N_3689,N_2838,N_2796);
or U3690 (N_3690,N_2951,N_2690);
nand U3691 (N_3691,N_2988,N_2766);
nand U3692 (N_3692,N_2680,N_3059);
nand U3693 (N_3693,N_2645,N_2655);
xor U3694 (N_3694,N_2604,N_2571);
or U3695 (N_3695,N_2815,N_2573);
or U3696 (N_3696,N_2774,N_2663);
xor U3697 (N_3697,N_2933,N_3102);
and U3698 (N_3698,N_2570,N_2711);
and U3699 (N_3699,N_2629,N_2759);
and U3700 (N_3700,N_2856,N_2732);
xnor U3701 (N_3701,N_2852,N_2793);
nor U3702 (N_3702,N_2745,N_3089);
xnor U3703 (N_3703,N_2518,N_2797);
nor U3704 (N_3704,N_2982,N_2729);
nor U3705 (N_3705,N_2835,N_2563);
and U3706 (N_3706,N_2793,N_3037);
xnor U3707 (N_3707,N_2835,N_2929);
nand U3708 (N_3708,N_2928,N_2562);
xor U3709 (N_3709,N_2663,N_2810);
nand U3710 (N_3710,N_3010,N_2691);
nand U3711 (N_3711,N_2794,N_2606);
nor U3712 (N_3712,N_2555,N_3068);
nor U3713 (N_3713,N_3040,N_2562);
and U3714 (N_3714,N_3034,N_3063);
xnor U3715 (N_3715,N_2789,N_3103);
nand U3716 (N_3716,N_3064,N_3025);
or U3717 (N_3717,N_2811,N_2767);
or U3718 (N_3718,N_2612,N_2875);
xnor U3719 (N_3719,N_2700,N_2974);
nor U3720 (N_3720,N_2597,N_3083);
or U3721 (N_3721,N_2687,N_2623);
and U3722 (N_3722,N_2754,N_2912);
xnor U3723 (N_3723,N_2771,N_3094);
nand U3724 (N_3724,N_2951,N_2898);
or U3725 (N_3725,N_3078,N_2799);
and U3726 (N_3726,N_3014,N_3090);
nand U3727 (N_3727,N_2540,N_2686);
xnor U3728 (N_3728,N_3026,N_2535);
xnor U3729 (N_3729,N_2733,N_2547);
nand U3730 (N_3730,N_3062,N_2704);
nor U3731 (N_3731,N_2651,N_2545);
xor U3732 (N_3732,N_2941,N_2757);
nor U3733 (N_3733,N_2975,N_2712);
xnor U3734 (N_3734,N_2889,N_3004);
nand U3735 (N_3735,N_2736,N_2546);
xnor U3736 (N_3736,N_2515,N_2546);
or U3737 (N_3737,N_2760,N_2675);
nor U3738 (N_3738,N_2804,N_2941);
or U3739 (N_3739,N_2747,N_2572);
or U3740 (N_3740,N_3066,N_2587);
nand U3741 (N_3741,N_2846,N_2594);
and U3742 (N_3742,N_2713,N_2812);
or U3743 (N_3743,N_2582,N_2844);
or U3744 (N_3744,N_2951,N_2810);
or U3745 (N_3745,N_2535,N_2919);
xnor U3746 (N_3746,N_2769,N_2877);
nor U3747 (N_3747,N_3102,N_2838);
nor U3748 (N_3748,N_2581,N_2840);
xor U3749 (N_3749,N_3096,N_3114);
nor U3750 (N_3750,N_3222,N_3496);
xnor U3751 (N_3751,N_3326,N_3285);
or U3752 (N_3752,N_3692,N_3453);
or U3753 (N_3753,N_3275,N_3637);
nor U3754 (N_3754,N_3740,N_3641);
and U3755 (N_3755,N_3373,N_3162);
xor U3756 (N_3756,N_3554,N_3584);
nor U3757 (N_3757,N_3708,N_3601);
or U3758 (N_3758,N_3623,N_3344);
and U3759 (N_3759,N_3359,N_3325);
or U3760 (N_3760,N_3257,N_3190);
nand U3761 (N_3761,N_3363,N_3445);
or U3762 (N_3762,N_3318,N_3742);
and U3763 (N_3763,N_3152,N_3675);
and U3764 (N_3764,N_3610,N_3519);
nor U3765 (N_3765,N_3308,N_3727);
nand U3766 (N_3766,N_3415,N_3165);
nor U3767 (N_3767,N_3220,N_3487);
and U3768 (N_3768,N_3357,N_3309);
nor U3769 (N_3769,N_3566,N_3316);
and U3770 (N_3770,N_3545,N_3322);
and U3771 (N_3771,N_3413,N_3243);
and U3772 (N_3772,N_3151,N_3592);
nand U3773 (N_3773,N_3369,N_3175);
nor U3774 (N_3774,N_3194,N_3185);
nand U3775 (N_3775,N_3382,N_3256);
or U3776 (N_3776,N_3150,N_3724);
or U3777 (N_3777,N_3435,N_3330);
and U3778 (N_3778,N_3507,N_3235);
and U3779 (N_3779,N_3139,N_3229);
xor U3780 (N_3780,N_3291,N_3443);
or U3781 (N_3781,N_3549,N_3405);
and U3782 (N_3782,N_3594,N_3276);
xor U3783 (N_3783,N_3631,N_3618);
or U3784 (N_3784,N_3379,N_3704);
and U3785 (N_3785,N_3624,N_3437);
nand U3786 (N_3786,N_3553,N_3749);
or U3787 (N_3787,N_3206,N_3505);
or U3788 (N_3788,N_3645,N_3176);
nand U3789 (N_3789,N_3391,N_3729);
xnor U3790 (N_3790,N_3733,N_3191);
nor U3791 (N_3791,N_3232,N_3538);
nor U3792 (N_3792,N_3690,N_3494);
and U3793 (N_3793,N_3705,N_3398);
or U3794 (N_3794,N_3512,N_3284);
nor U3795 (N_3795,N_3657,N_3573);
nand U3796 (N_3796,N_3468,N_3723);
nand U3797 (N_3797,N_3451,N_3649);
and U3798 (N_3798,N_3493,N_3524);
nor U3799 (N_3799,N_3575,N_3201);
and U3800 (N_3800,N_3476,N_3608);
and U3801 (N_3801,N_3492,N_3539);
and U3802 (N_3802,N_3676,N_3252);
and U3803 (N_3803,N_3368,N_3170);
or U3804 (N_3804,N_3163,N_3598);
nand U3805 (N_3805,N_3313,N_3720);
or U3806 (N_3806,N_3699,N_3726);
or U3807 (N_3807,N_3745,N_3134);
and U3808 (N_3808,N_3366,N_3181);
nand U3809 (N_3809,N_3423,N_3665);
or U3810 (N_3810,N_3239,N_3427);
or U3811 (N_3811,N_3396,N_3130);
xor U3812 (N_3812,N_3634,N_3362);
nand U3813 (N_3813,N_3590,N_3630);
or U3814 (N_3814,N_3739,N_3455);
nand U3815 (N_3815,N_3157,N_3364);
nor U3816 (N_3816,N_3551,N_3462);
xor U3817 (N_3817,N_3638,N_3254);
nor U3818 (N_3818,N_3214,N_3365);
and U3819 (N_3819,N_3467,N_3557);
and U3820 (N_3820,N_3342,N_3619);
nor U3821 (N_3821,N_3523,N_3390);
nand U3822 (N_3822,N_3650,N_3211);
or U3823 (N_3823,N_3138,N_3567);
and U3824 (N_3824,N_3355,N_3574);
nand U3825 (N_3825,N_3329,N_3412);
nand U3826 (N_3826,N_3367,N_3346);
and U3827 (N_3827,N_3188,N_3597);
nand U3828 (N_3828,N_3678,N_3295);
xor U3829 (N_3829,N_3454,N_3743);
nor U3830 (N_3830,N_3228,N_3502);
nor U3831 (N_3831,N_3240,N_3444);
nor U3832 (N_3832,N_3570,N_3639);
nor U3833 (N_3833,N_3663,N_3155);
nand U3834 (N_3834,N_3140,N_3732);
nor U3835 (N_3835,N_3700,N_3563);
nor U3836 (N_3836,N_3506,N_3522);
nand U3837 (N_3837,N_3450,N_3253);
and U3838 (N_3838,N_3560,N_3304);
nor U3839 (N_3839,N_3255,N_3516);
or U3840 (N_3840,N_3298,N_3319);
or U3841 (N_3841,N_3360,N_3161);
nor U3842 (N_3842,N_3466,N_3338);
nor U3843 (N_3843,N_3555,N_3281);
or U3844 (N_3844,N_3274,N_3137);
or U3845 (N_3845,N_3670,N_3528);
or U3846 (N_3846,N_3408,N_3658);
or U3847 (N_3847,N_3534,N_3677);
or U3848 (N_3848,N_3414,N_3456);
nand U3849 (N_3849,N_3470,N_3612);
xor U3850 (N_3850,N_3210,N_3581);
nor U3851 (N_3851,N_3707,N_3301);
xor U3852 (N_3852,N_3474,N_3218);
nor U3853 (N_3853,N_3636,N_3579);
or U3854 (N_3854,N_3350,N_3683);
or U3855 (N_3855,N_3404,N_3387);
nand U3856 (N_3856,N_3230,N_3282);
xor U3857 (N_3857,N_3583,N_3389);
or U3858 (N_3858,N_3400,N_3629);
nand U3859 (N_3859,N_3717,N_3548);
xor U3860 (N_3860,N_3447,N_3544);
or U3861 (N_3861,N_3627,N_3302);
and U3862 (N_3862,N_3374,N_3688);
or U3863 (N_3863,N_3153,N_3486);
nand U3864 (N_3864,N_3244,N_3307);
nand U3865 (N_3865,N_3543,N_3179);
and U3866 (N_3866,N_3681,N_3686);
and U3867 (N_3867,N_3578,N_3283);
xor U3868 (N_3868,N_3353,N_3697);
nor U3869 (N_3869,N_3489,N_3438);
nand U3870 (N_3870,N_3217,N_3261);
nand U3871 (N_3871,N_3320,N_3406);
nand U3872 (N_3872,N_3526,N_3585);
xnor U3873 (N_3873,N_3241,N_3540);
nor U3874 (N_3874,N_3334,N_3303);
or U3875 (N_3875,N_3602,N_3485);
nor U3876 (N_3876,N_3737,N_3336);
nand U3877 (N_3877,N_3399,N_3682);
or U3878 (N_3878,N_3383,N_3345);
nor U3879 (N_3879,N_3317,N_3187);
and U3880 (N_3880,N_3127,N_3694);
nand U3881 (N_3881,N_3245,N_3576);
nor U3882 (N_3882,N_3591,N_3497);
nand U3883 (N_3883,N_3656,N_3258);
nand U3884 (N_3884,N_3464,N_3648);
nor U3885 (N_3885,N_3515,N_3718);
nor U3886 (N_3886,N_3393,N_3469);
or U3887 (N_3887,N_3333,N_3710);
nand U3888 (N_3888,N_3171,N_3478);
nand U3889 (N_3889,N_3148,N_3132);
xnor U3890 (N_3890,N_3738,N_3609);
nand U3891 (N_3891,N_3735,N_3324);
xnor U3892 (N_3892,N_3586,N_3503);
and U3893 (N_3893,N_3457,N_3674);
nand U3894 (N_3894,N_3625,N_3558);
nand U3895 (N_3895,N_3352,N_3472);
nor U3896 (N_3896,N_3606,N_3263);
or U3897 (N_3897,N_3626,N_3268);
nor U3898 (N_3898,N_3440,N_3696);
xor U3899 (N_3899,N_3529,N_3667);
nand U3900 (N_3900,N_3380,N_3193);
nor U3901 (N_3901,N_3501,N_3397);
xor U3902 (N_3902,N_3533,N_3418);
or U3903 (N_3903,N_3593,N_3315);
nand U3904 (N_3904,N_3465,N_3141);
and U3905 (N_3905,N_3296,N_3142);
nand U3906 (N_3906,N_3673,N_3247);
nor U3907 (N_3907,N_3265,N_3358);
or U3908 (N_3908,N_3215,N_3266);
or U3909 (N_3909,N_3668,N_3728);
xor U3910 (N_3910,N_3323,N_3143);
nor U3911 (N_3911,N_3203,N_3286);
or U3912 (N_3912,N_3335,N_3174);
nor U3913 (N_3913,N_3480,N_3577);
nand U3914 (N_3914,N_3731,N_3747);
or U3915 (N_3915,N_3173,N_3482);
and U3916 (N_3916,N_3411,N_3518);
nor U3917 (N_3917,N_3279,N_3483);
or U3918 (N_3918,N_3491,N_3426);
nand U3919 (N_3919,N_3633,N_3653);
xor U3920 (N_3920,N_3300,N_3388);
nor U3921 (N_3921,N_3199,N_3164);
xnor U3922 (N_3922,N_3647,N_3730);
or U3923 (N_3923,N_3223,N_3290);
nand U3924 (N_3924,N_3622,N_3292);
nor U3925 (N_3925,N_3655,N_3213);
nand U3926 (N_3926,N_3452,N_3734);
nor U3927 (N_3927,N_3209,N_3154);
nor U3928 (N_3928,N_3706,N_3589);
nor U3929 (N_3929,N_3477,N_3632);
nor U3930 (N_3930,N_3640,N_3672);
nand U3931 (N_3931,N_3685,N_3499);
nor U3932 (N_3932,N_3273,N_3378);
nand U3933 (N_3933,N_3687,N_3237);
nand U3934 (N_3934,N_3416,N_3702);
and U3935 (N_3935,N_3736,N_3371);
and U3936 (N_3936,N_3607,N_3536);
and U3937 (N_3937,N_3337,N_3488);
or U3938 (N_3938,N_3661,N_3125);
nand U3939 (N_3939,N_3375,N_3495);
or U3940 (N_3940,N_3725,N_3156);
nor U3941 (N_3941,N_3160,N_3180);
nor U3942 (N_3942,N_3703,N_3272);
xnor U3943 (N_3943,N_3225,N_3294);
nand U3944 (N_3944,N_3565,N_3562);
xnor U3945 (N_3945,N_3711,N_3613);
nor U3946 (N_3946,N_3611,N_3689);
xnor U3947 (N_3947,N_3394,N_3410);
or U3948 (N_3948,N_3131,N_3401);
xnor U3949 (N_3949,N_3671,N_3662);
nand U3950 (N_3950,N_3428,N_3429);
or U3951 (N_3951,N_3666,N_3644);
xor U3952 (N_3952,N_3182,N_3587);
and U3953 (N_3953,N_3509,N_3569);
xnor U3954 (N_3954,N_3270,N_3475);
nand U3955 (N_3955,N_3521,N_3490);
nand U3956 (N_3956,N_3133,N_3189);
nor U3957 (N_3957,N_3441,N_3424);
xor U3958 (N_3958,N_3425,N_3145);
nand U3959 (N_3959,N_3341,N_3205);
nand U3960 (N_3960,N_3340,N_3541);
xor U3961 (N_3961,N_3432,N_3236);
or U3962 (N_3962,N_3433,N_3719);
nand U3963 (N_3963,N_3159,N_3234);
nand U3964 (N_3964,N_3348,N_3635);
nor U3965 (N_3965,N_3321,N_3517);
xor U3966 (N_3966,N_3278,N_3714);
nand U3967 (N_3967,N_3224,N_3530);
or U3968 (N_3968,N_3402,N_3208);
or U3969 (N_3969,N_3376,N_3126);
nor U3970 (N_3970,N_3616,N_3604);
nor U3971 (N_3971,N_3546,N_3242);
or U3972 (N_3972,N_3233,N_3596);
xnor U3973 (N_3973,N_3332,N_3259);
or U3974 (N_3974,N_3392,N_3463);
xnor U3975 (N_3975,N_3356,N_3471);
nand U3976 (N_3976,N_3547,N_3385);
or U3977 (N_3977,N_3314,N_3354);
nor U3978 (N_3978,N_3514,N_3484);
nor U3979 (N_3979,N_3395,N_3741);
xnor U3980 (N_3980,N_3449,N_3621);
or U3981 (N_3981,N_3407,N_3204);
and U3982 (N_3982,N_3197,N_3461);
nor U3983 (N_3983,N_3654,N_3498);
or U3984 (N_3984,N_3542,N_3599);
nor U3985 (N_3985,N_3246,N_3167);
nor U3986 (N_3986,N_3479,N_3251);
nand U3987 (N_3987,N_3693,N_3250);
nand U3988 (N_3988,N_3198,N_3660);
nand U3989 (N_3989,N_3299,N_3481);
or U3990 (N_3990,N_3691,N_3178);
nand U3991 (N_3991,N_3327,N_3709);
nand U3992 (N_3992,N_3559,N_3361);
xnor U3993 (N_3993,N_3520,N_3531);
nor U3994 (N_3994,N_3177,N_3664);
and U3995 (N_3995,N_3422,N_3381);
or U3996 (N_3996,N_3288,N_3147);
or U3997 (N_3997,N_3409,N_3716);
nor U3998 (N_3998,N_3202,N_3473);
or U3999 (N_3999,N_3311,N_3262);
xnor U4000 (N_4000,N_3564,N_3200);
or U4001 (N_4001,N_3168,N_3669);
xnor U4002 (N_4002,N_3504,N_3746);
xnor U4003 (N_4003,N_3216,N_3128);
nand U4004 (N_4004,N_3620,N_3588);
or U4005 (N_4005,N_3701,N_3417);
nor U4006 (N_4006,N_3527,N_3431);
or U4007 (N_4007,N_3525,N_3196);
or U4008 (N_4008,N_3508,N_3386);
and U4009 (N_4009,N_3331,N_3561);
or U4010 (N_4010,N_3603,N_3744);
and U4011 (N_4011,N_3459,N_3277);
nand U4012 (N_4012,N_3537,N_3582);
nand U4013 (N_4013,N_3721,N_3219);
nand U4014 (N_4014,N_3183,N_3651);
nor U4015 (N_4015,N_3146,N_3227);
and U4016 (N_4016,N_3184,N_3614);
nand U4017 (N_4017,N_3446,N_3195);
xnor U4018 (N_4018,N_3448,N_3231);
and U4019 (N_4019,N_3172,N_3430);
and U4020 (N_4020,N_3436,N_3421);
nor U4021 (N_4021,N_3420,N_3748);
and U4022 (N_4022,N_3552,N_3166);
nor U4023 (N_4023,N_3510,N_3238);
or U4024 (N_4024,N_3679,N_3600);
xnor U4025 (N_4025,N_3249,N_3269);
or U4026 (N_4026,N_3550,N_3271);
and U4027 (N_4027,N_3434,N_3642);
nor U4028 (N_4028,N_3698,N_3248);
and U4029 (N_4029,N_3377,N_3267);
nand U4030 (N_4030,N_3192,N_3144);
and U4031 (N_4031,N_3722,N_3615);
or U4032 (N_4032,N_3580,N_3511);
or U4033 (N_4033,N_3403,N_3646);
or U4034 (N_4034,N_3628,N_3169);
xor U4035 (N_4035,N_3617,N_3339);
or U4036 (N_4036,N_3343,N_3535);
xnor U4037 (N_4037,N_3328,N_3556);
or U4038 (N_4038,N_3370,N_3136);
xor U4039 (N_4039,N_3572,N_3135);
or U4040 (N_4040,N_3221,N_3680);
or U4041 (N_4041,N_3643,N_3306);
and U4042 (N_4042,N_3439,N_3568);
nand U4043 (N_4043,N_3460,N_3207);
and U4044 (N_4044,N_3349,N_3513);
xnor U4045 (N_4045,N_3260,N_3532);
or U4046 (N_4046,N_3226,N_3571);
xnor U4047 (N_4047,N_3129,N_3419);
and U4048 (N_4048,N_3458,N_3280);
nand U4049 (N_4049,N_3442,N_3713);
nand U4050 (N_4050,N_3659,N_3287);
nor U4051 (N_4051,N_3652,N_3351);
nand U4052 (N_4052,N_3312,N_3712);
or U4053 (N_4053,N_3605,N_3293);
nand U4054 (N_4054,N_3384,N_3310);
xor U4055 (N_4055,N_3595,N_3297);
and U4056 (N_4056,N_3289,N_3695);
nand U4057 (N_4057,N_3715,N_3264);
nor U4058 (N_4058,N_3372,N_3684);
nor U4059 (N_4059,N_3186,N_3212);
nor U4060 (N_4060,N_3149,N_3158);
and U4061 (N_4061,N_3500,N_3347);
and U4062 (N_4062,N_3305,N_3374);
xor U4063 (N_4063,N_3402,N_3159);
or U4064 (N_4064,N_3160,N_3522);
or U4065 (N_4065,N_3185,N_3220);
and U4066 (N_4066,N_3150,N_3334);
or U4067 (N_4067,N_3500,N_3265);
xnor U4068 (N_4068,N_3471,N_3299);
nand U4069 (N_4069,N_3394,N_3206);
nor U4070 (N_4070,N_3176,N_3607);
and U4071 (N_4071,N_3715,N_3669);
nor U4072 (N_4072,N_3137,N_3457);
xor U4073 (N_4073,N_3315,N_3228);
and U4074 (N_4074,N_3299,N_3633);
xor U4075 (N_4075,N_3622,N_3703);
and U4076 (N_4076,N_3563,N_3159);
or U4077 (N_4077,N_3643,N_3384);
and U4078 (N_4078,N_3568,N_3496);
or U4079 (N_4079,N_3597,N_3621);
or U4080 (N_4080,N_3676,N_3521);
nand U4081 (N_4081,N_3344,N_3331);
xor U4082 (N_4082,N_3325,N_3660);
and U4083 (N_4083,N_3517,N_3411);
and U4084 (N_4084,N_3180,N_3640);
nor U4085 (N_4085,N_3483,N_3593);
xnor U4086 (N_4086,N_3557,N_3278);
nor U4087 (N_4087,N_3421,N_3153);
and U4088 (N_4088,N_3213,N_3708);
nand U4089 (N_4089,N_3227,N_3585);
and U4090 (N_4090,N_3277,N_3348);
nand U4091 (N_4091,N_3452,N_3483);
and U4092 (N_4092,N_3351,N_3235);
and U4093 (N_4093,N_3477,N_3259);
or U4094 (N_4094,N_3479,N_3131);
nand U4095 (N_4095,N_3165,N_3564);
or U4096 (N_4096,N_3154,N_3615);
and U4097 (N_4097,N_3210,N_3253);
xnor U4098 (N_4098,N_3433,N_3499);
xor U4099 (N_4099,N_3515,N_3656);
and U4100 (N_4100,N_3328,N_3543);
nor U4101 (N_4101,N_3608,N_3680);
nor U4102 (N_4102,N_3634,N_3503);
or U4103 (N_4103,N_3278,N_3692);
nor U4104 (N_4104,N_3421,N_3325);
nand U4105 (N_4105,N_3604,N_3637);
or U4106 (N_4106,N_3605,N_3697);
or U4107 (N_4107,N_3573,N_3564);
or U4108 (N_4108,N_3483,N_3242);
or U4109 (N_4109,N_3497,N_3396);
nand U4110 (N_4110,N_3542,N_3240);
and U4111 (N_4111,N_3227,N_3596);
nor U4112 (N_4112,N_3448,N_3559);
or U4113 (N_4113,N_3649,N_3729);
nand U4114 (N_4114,N_3450,N_3591);
and U4115 (N_4115,N_3627,N_3170);
or U4116 (N_4116,N_3354,N_3228);
nor U4117 (N_4117,N_3169,N_3500);
and U4118 (N_4118,N_3379,N_3639);
xor U4119 (N_4119,N_3690,N_3216);
nand U4120 (N_4120,N_3671,N_3308);
nand U4121 (N_4121,N_3691,N_3600);
xor U4122 (N_4122,N_3414,N_3200);
xor U4123 (N_4123,N_3525,N_3639);
xnor U4124 (N_4124,N_3517,N_3418);
xnor U4125 (N_4125,N_3251,N_3331);
xnor U4126 (N_4126,N_3487,N_3252);
xnor U4127 (N_4127,N_3143,N_3636);
nand U4128 (N_4128,N_3446,N_3234);
or U4129 (N_4129,N_3486,N_3705);
and U4130 (N_4130,N_3336,N_3723);
xnor U4131 (N_4131,N_3585,N_3461);
nand U4132 (N_4132,N_3317,N_3420);
nor U4133 (N_4133,N_3132,N_3561);
nor U4134 (N_4134,N_3271,N_3718);
nor U4135 (N_4135,N_3656,N_3267);
or U4136 (N_4136,N_3590,N_3693);
nor U4137 (N_4137,N_3324,N_3385);
nor U4138 (N_4138,N_3540,N_3711);
nand U4139 (N_4139,N_3448,N_3476);
or U4140 (N_4140,N_3341,N_3474);
and U4141 (N_4141,N_3528,N_3461);
nor U4142 (N_4142,N_3398,N_3163);
or U4143 (N_4143,N_3575,N_3458);
nor U4144 (N_4144,N_3707,N_3641);
and U4145 (N_4145,N_3663,N_3333);
or U4146 (N_4146,N_3469,N_3466);
and U4147 (N_4147,N_3641,N_3655);
or U4148 (N_4148,N_3522,N_3691);
and U4149 (N_4149,N_3282,N_3136);
or U4150 (N_4150,N_3434,N_3396);
nor U4151 (N_4151,N_3714,N_3573);
or U4152 (N_4152,N_3387,N_3371);
and U4153 (N_4153,N_3358,N_3293);
or U4154 (N_4154,N_3601,N_3384);
or U4155 (N_4155,N_3197,N_3621);
nand U4156 (N_4156,N_3555,N_3426);
and U4157 (N_4157,N_3586,N_3444);
xnor U4158 (N_4158,N_3295,N_3376);
nand U4159 (N_4159,N_3522,N_3703);
nor U4160 (N_4160,N_3511,N_3437);
or U4161 (N_4161,N_3395,N_3517);
nand U4162 (N_4162,N_3413,N_3693);
or U4163 (N_4163,N_3687,N_3149);
or U4164 (N_4164,N_3428,N_3474);
xnor U4165 (N_4165,N_3359,N_3126);
or U4166 (N_4166,N_3460,N_3738);
nor U4167 (N_4167,N_3602,N_3563);
nor U4168 (N_4168,N_3595,N_3507);
or U4169 (N_4169,N_3461,N_3704);
or U4170 (N_4170,N_3458,N_3176);
xor U4171 (N_4171,N_3182,N_3222);
nor U4172 (N_4172,N_3445,N_3142);
or U4173 (N_4173,N_3361,N_3713);
xor U4174 (N_4174,N_3125,N_3432);
nor U4175 (N_4175,N_3191,N_3255);
nor U4176 (N_4176,N_3310,N_3346);
or U4177 (N_4177,N_3721,N_3170);
xor U4178 (N_4178,N_3199,N_3390);
or U4179 (N_4179,N_3539,N_3628);
or U4180 (N_4180,N_3226,N_3720);
xnor U4181 (N_4181,N_3413,N_3586);
or U4182 (N_4182,N_3219,N_3475);
xnor U4183 (N_4183,N_3733,N_3421);
nor U4184 (N_4184,N_3368,N_3326);
nor U4185 (N_4185,N_3400,N_3229);
nand U4186 (N_4186,N_3474,N_3686);
nor U4187 (N_4187,N_3484,N_3679);
and U4188 (N_4188,N_3406,N_3378);
nor U4189 (N_4189,N_3144,N_3674);
and U4190 (N_4190,N_3430,N_3452);
nor U4191 (N_4191,N_3475,N_3472);
or U4192 (N_4192,N_3499,N_3396);
xnor U4193 (N_4193,N_3481,N_3358);
and U4194 (N_4194,N_3466,N_3587);
nand U4195 (N_4195,N_3684,N_3570);
nor U4196 (N_4196,N_3320,N_3619);
nor U4197 (N_4197,N_3652,N_3392);
and U4198 (N_4198,N_3708,N_3203);
xnor U4199 (N_4199,N_3437,N_3567);
nand U4200 (N_4200,N_3514,N_3367);
xnor U4201 (N_4201,N_3679,N_3635);
and U4202 (N_4202,N_3461,N_3550);
and U4203 (N_4203,N_3727,N_3244);
and U4204 (N_4204,N_3280,N_3555);
and U4205 (N_4205,N_3471,N_3712);
xor U4206 (N_4206,N_3524,N_3396);
and U4207 (N_4207,N_3287,N_3295);
or U4208 (N_4208,N_3653,N_3252);
nand U4209 (N_4209,N_3667,N_3393);
xnor U4210 (N_4210,N_3580,N_3265);
nand U4211 (N_4211,N_3161,N_3561);
or U4212 (N_4212,N_3218,N_3568);
nand U4213 (N_4213,N_3266,N_3553);
nor U4214 (N_4214,N_3185,N_3238);
nor U4215 (N_4215,N_3326,N_3579);
or U4216 (N_4216,N_3499,N_3170);
nand U4217 (N_4217,N_3278,N_3306);
or U4218 (N_4218,N_3584,N_3289);
and U4219 (N_4219,N_3485,N_3685);
nand U4220 (N_4220,N_3466,N_3152);
or U4221 (N_4221,N_3265,N_3164);
or U4222 (N_4222,N_3290,N_3150);
nor U4223 (N_4223,N_3585,N_3630);
xnor U4224 (N_4224,N_3470,N_3747);
nor U4225 (N_4225,N_3391,N_3529);
or U4226 (N_4226,N_3487,N_3225);
or U4227 (N_4227,N_3597,N_3539);
nor U4228 (N_4228,N_3671,N_3333);
nand U4229 (N_4229,N_3206,N_3550);
nor U4230 (N_4230,N_3411,N_3415);
and U4231 (N_4231,N_3524,N_3721);
xnor U4232 (N_4232,N_3676,N_3212);
xnor U4233 (N_4233,N_3301,N_3203);
xnor U4234 (N_4234,N_3661,N_3611);
nor U4235 (N_4235,N_3651,N_3740);
nor U4236 (N_4236,N_3247,N_3530);
nor U4237 (N_4237,N_3366,N_3325);
nor U4238 (N_4238,N_3666,N_3719);
and U4239 (N_4239,N_3299,N_3476);
nor U4240 (N_4240,N_3330,N_3157);
nand U4241 (N_4241,N_3457,N_3571);
and U4242 (N_4242,N_3342,N_3273);
nand U4243 (N_4243,N_3724,N_3382);
nor U4244 (N_4244,N_3383,N_3281);
nor U4245 (N_4245,N_3385,N_3437);
or U4246 (N_4246,N_3342,N_3639);
or U4247 (N_4247,N_3439,N_3671);
nand U4248 (N_4248,N_3416,N_3288);
nand U4249 (N_4249,N_3708,N_3306);
nor U4250 (N_4250,N_3562,N_3607);
xor U4251 (N_4251,N_3531,N_3579);
nand U4252 (N_4252,N_3630,N_3315);
and U4253 (N_4253,N_3623,N_3478);
and U4254 (N_4254,N_3740,N_3647);
or U4255 (N_4255,N_3385,N_3130);
and U4256 (N_4256,N_3596,N_3471);
nand U4257 (N_4257,N_3280,N_3271);
nor U4258 (N_4258,N_3646,N_3323);
xor U4259 (N_4259,N_3589,N_3407);
nand U4260 (N_4260,N_3261,N_3546);
or U4261 (N_4261,N_3417,N_3741);
and U4262 (N_4262,N_3632,N_3251);
nand U4263 (N_4263,N_3433,N_3470);
xnor U4264 (N_4264,N_3531,N_3146);
or U4265 (N_4265,N_3539,N_3687);
nor U4266 (N_4266,N_3491,N_3524);
or U4267 (N_4267,N_3217,N_3513);
xnor U4268 (N_4268,N_3314,N_3540);
or U4269 (N_4269,N_3701,N_3489);
and U4270 (N_4270,N_3511,N_3396);
nor U4271 (N_4271,N_3634,N_3688);
and U4272 (N_4272,N_3400,N_3699);
or U4273 (N_4273,N_3136,N_3335);
and U4274 (N_4274,N_3298,N_3493);
and U4275 (N_4275,N_3417,N_3307);
xor U4276 (N_4276,N_3411,N_3685);
or U4277 (N_4277,N_3385,N_3231);
nor U4278 (N_4278,N_3390,N_3737);
and U4279 (N_4279,N_3726,N_3551);
nor U4280 (N_4280,N_3667,N_3504);
and U4281 (N_4281,N_3557,N_3619);
xnor U4282 (N_4282,N_3528,N_3518);
xor U4283 (N_4283,N_3446,N_3398);
xnor U4284 (N_4284,N_3240,N_3494);
xnor U4285 (N_4285,N_3647,N_3632);
xor U4286 (N_4286,N_3602,N_3596);
or U4287 (N_4287,N_3149,N_3519);
nor U4288 (N_4288,N_3382,N_3659);
or U4289 (N_4289,N_3586,N_3271);
xnor U4290 (N_4290,N_3274,N_3449);
xnor U4291 (N_4291,N_3533,N_3186);
and U4292 (N_4292,N_3663,N_3558);
xor U4293 (N_4293,N_3235,N_3338);
xnor U4294 (N_4294,N_3465,N_3182);
xnor U4295 (N_4295,N_3195,N_3353);
and U4296 (N_4296,N_3545,N_3258);
xnor U4297 (N_4297,N_3207,N_3733);
or U4298 (N_4298,N_3274,N_3348);
nor U4299 (N_4299,N_3227,N_3427);
xnor U4300 (N_4300,N_3201,N_3527);
or U4301 (N_4301,N_3273,N_3676);
or U4302 (N_4302,N_3489,N_3512);
or U4303 (N_4303,N_3218,N_3336);
and U4304 (N_4304,N_3242,N_3606);
and U4305 (N_4305,N_3514,N_3741);
nand U4306 (N_4306,N_3440,N_3450);
nand U4307 (N_4307,N_3260,N_3601);
xor U4308 (N_4308,N_3670,N_3689);
and U4309 (N_4309,N_3514,N_3708);
nand U4310 (N_4310,N_3592,N_3566);
nand U4311 (N_4311,N_3711,N_3640);
or U4312 (N_4312,N_3132,N_3581);
nand U4313 (N_4313,N_3452,N_3346);
nor U4314 (N_4314,N_3336,N_3178);
or U4315 (N_4315,N_3149,N_3235);
xor U4316 (N_4316,N_3194,N_3348);
nand U4317 (N_4317,N_3172,N_3730);
nor U4318 (N_4318,N_3261,N_3207);
xnor U4319 (N_4319,N_3425,N_3646);
xnor U4320 (N_4320,N_3208,N_3181);
xnor U4321 (N_4321,N_3615,N_3669);
or U4322 (N_4322,N_3256,N_3748);
nand U4323 (N_4323,N_3315,N_3195);
or U4324 (N_4324,N_3335,N_3191);
nand U4325 (N_4325,N_3377,N_3416);
and U4326 (N_4326,N_3721,N_3273);
nor U4327 (N_4327,N_3478,N_3543);
or U4328 (N_4328,N_3548,N_3261);
nand U4329 (N_4329,N_3636,N_3323);
nor U4330 (N_4330,N_3297,N_3186);
nand U4331 (N_4331,N_3642,N_3322);
nand U4332 (N_4332,N_3431,N_3450);
nor U4333 (N_4333,N_3623,N_3287);
xnor U4334 (N_4334,N_3536,N_3639);
nand U4335 (N_4335,N_3197,N_3129);
and U4336 (N_4336,N_3639,N_3212);
and U4337 (N_4337,N_3365,N_3300);
or U4338 (N_4338,N_3212,N_3159);
nor U4339 (N_4339,N_3602,N_3325);
nand U4340 (N_4340,N_3530,N_3715);
and U4341 (N_4341,N_3397,N_3384);
nor U4342 (N_4342,N_3190,N_3516);
or U4343 (N_4343,N_3348,N_3480);
and U4344 (N_4344,N_3424,N_3198);
and U4345 (N_4345,N_3333,N_3226);
or U4346 (N_4346,N_3601,N_3741);
nor U4347 (N_4347,N_3241,N_3411);
xor U4348 (N_4348,N_3376,N_3358);
nor U4349 (N_4349,N_3464,N_3192);
or U4350 (N_4350,N_3152,N_3361);
nor U4351 (N_4351,N_3247,N_3620);
nand U4352 (N_4352,N_3392,N_3387);
or U4353 (N_4353,N_3229,N_3132);
and U4354 (N_4354,N_3289,N_3641);
xor U4355 (N_4355,N_3164,N_3497);
and U4356 (N_4356,N_3404,N_3646);
nand U4357 (N_4357,N_3410,N_3184);
and U4358 (N_4358,N_3311,N_3524);
and U4359 (N_4359,N_3284,N_3632);
nor U4360 (N_4360,N_3459,N_3591);
nor U4361 (N_4361,N_3254,N_3601);
and U4362 (N_4362,N_3420,N_3136);
nand U4363 (N_4363,N_3663,N_3344);
and U4364 (N_4364,N_3173,N_3150);
nand U4365 (N_4365,N_3216,N_3414);
nor U4366 (N_4366,N_3127,N_3158);
or U4367 (N_4367,N_3186,N_3192);
or U4368 (N_4368,N_3615,N_3219);
nand U4369 (N_4369,N_3405,N_3167);
nor U4370 (N_4370,N_3247,N_3684);
or U4371 (N_4371,N_3503,N_3140);
and U4372 (N_4372,N_3504,N_3266);
or U4373 (N_4373,N_3658,N_3461);
xor U4374 (N_4374,N_3663,N_3548);
or U4375 (N_4375,N_3951,N_4355);
and U4376 (N_4376,N_4335,N_3913);
nor U4377 (N_4377,N_4341,N_3933);
xnor U4378 (N_4378,N_4037,N_4329);
xor U4379 (N_4379,N_3904,N_4297);
and U4380 (N_4380,N_3874,N_3751);
and U4381 (N_4381,N_4151,N_4209);
nand U4382 (N_4382,N_4241,N_3909);
or U4383 (N_4383,N_4169,N_4350);
or U4384 (N_4384,N_4084,N_4236);
nand U4385 (N_4385,N_3830,N_4283);
and U4386 (N_4386,N_4332,N_3801);
and U4387 (N_4387,N_4003,N_4277);
nor U4388 (N_4388,N_4027,N_3984);
nor U4389 (N_4389,N_4343,N_3838);
or U4390 (N_4390,N_4345,N_3910);
xor U4391 (N_4391,N_3976,N_4161);
xnor U4392 (N_4392,N_3990,N_4136);
nor U4393 (N_4393,N_4020,N_4077);
nand U4394 (N_4394,N_3760,N_3899);
nor U4395 (N_4395,N_3887,N_4285);
nand U4396 (N_4396,N_4170,N_4134);
nand U4397 (N_4397,N_4087,N_4102);
nand U4398 (N_4398,N_4204,N_3870);
nand U4399 (N_4399,N_4127,N_4305);
and U4400 (N_4400,N_3817,N_3989);
nand U4401 (N_4401,N_3805,N_4255);
and U4402 (N_4402,N_4230,N_3831);
xor U4403 (N_4403,N_3950,N_4122);
nand U4404 (N_4404,N_3856,N_3977);
and U4405 (N_4405,N_4271,N_4357);
nor U4406 (N_4406,N_4330,N_4146);
or U4407 (N_4407,N_4059,N_3929);
xor U4408 (N_4408,N_3793,N_4064);
nand U4409 (N_4409,N_4165,N_4094);
and U4410 (N_4410,N_3762,N_4337);
and U4411 (N_4411,N_3768,N_3982);
xor U4412 (N_4412,N_4289,N_4017);
nand U4413 (N_4413,N_3936,N_3814);
nor U4414 (N_4414,N_4254,N_4183);
nand U4415 (N_4415,N_3935,N_3795);
and U4416 (N_4416,N_3975,N_4257);
xor U4417 (N_4417,N_4286,N_4206);
xor U4418 (N_4418,N_3809,N_4348);
and U4419 (N_4419,N_4125,N_4298);
xnor U4420 (N_4420,N_3850,N_4320);
nor U4421 (N_4421,N_3774,N_3857);
nor U4422 (N_4422,N_4242,N_3894);
and U4423 (N_4423,N_3993,N_4062);
nand U4424 (N_4424,N_4089,N_4083);
or U4425 (N_4425,N_3833,N_4006);
or U4426 (N_4426,N_3859,N_4051);
xor U4427 (N_4427,N_4314,N_4155);
nor U4428 (N_4428,N_4253,N_3781);
nor U4429 (N_4429,N_4181,N_3869);
xnor U4430 (N_4430,N_4123,N_4187);
nand U4431 (N_4431,N_3867,N_4328);
or U4432 (N_4432,N_4312,N_4024);
nor U4433 (N_4433,N_3962,N_3901);
nand U4434 (N_4434,N_4069,N_4226);
nand U4435 (N_4435,N_3794,N_3862);
or U4436 (N_4436,N_3879,N_4260);
nor U4437 (N_4437,N_4115,N_4245);
and U4438 (N_4438,N_3773,N_4081);
xnor U4439 (N_4439,N_4036,N_3979);
xnor U4440 (N_4440,N_3953,N_4019);
and U4441 (N_4441,N_4216,N_4126);
or U4442 (N_4442,N_3758,N_4067);
xnor U4443 (N_4443,N_4053,N_3841);
nor U4444 (N_4444,N_4198,N_3797);
nor U4445 (N_4445,N_3789,N_4291);
nor U4446 (N_4446,N_4353,N_4093);
or U4447 (N_4447,N_3853,N_4150);
or U4448 (N_4448,N_4045,N_3945);
and U4449 (N_4449,N_4360,N_4124);
and U4450 (N_4450,N_4352,N_3983);
nand U4451 (N_4451,N_4221,N_4303);
nor U4452 (N_4452,N_3848,N_4208);
or U4453 (N_4453,N_4218,N_4046);
and U4454 (N_4454,N_3966,N_4296);
or U4455 (N_4455,N_4055,N_4004);
or U4456 (N_4456,N_4143,N_4160);
or U4457 (N_4457,N_4080,N_3931);
and U4458 (N_4458,N_4304,N_3985);
and U4459 (N_4459,N_4131,N_4050);
nand U4460 (N_4460,N_4092,N_4032);
and U4461 (N_4461,N_4354,N_4294);
and U4462 (N_4462,N_3974,N_3996);
or U4463 (N_4463,N_3852,N_4322);
or U4464 (N_4464,N_3865,N_3769);
and U4465 (N_4465,N_4044,N_4340);
and U4466 (N_4466,N_4323,N_4261);
or U4467 (N_4467,N_4212,N_3961);
or U4468 (N_4468,N_3821,N_4367);
and U4469 (N_4469,N_4248,N_3861);
and U4470 (N_4470,N_4295,N_4108);
nor U4471 (N_4471,N_3855,N_4147);
and U4472 (N_4472,N_3854,N_4041);
xnor U4473 (N_4473,N_4109,N_3788);
and U4474 (N_4474,N_4047,N_4188);
xnor U4475 (N_4475,N_4210,N_4023);
and U4476 (N_4476,N_3766,N_3750);
or U4477 (N_4477,N_3836,N_4072);
nand U4478 (N_4478,N_3928,N_3900);
and U4479 (N_4479,N_4268,N_3778);
nor U4480 (N_4480,N_4192,N_4293);
xnor U4481 (N_4481,N_3994,N_4244);
nor U4482 (N_4482,N_3969,N_4334);
or U4483 (N_4483,N_3888,N_4316);
and U4484 (N_4484,N_4030,N_4139);
nand U4485 (N_4485,N_4272,N_4356);
or U4486 (N_4486,N_4365,N_3905);
or U4487 (N_4487,N_3756,N_4052);
and U4488 (N_4488,N_3823,N_3753);
or U4489 (N_4489,N_4137,N_3840);
nor U4490 (N_4490,N_3921,N_4145);
or U4491 (N_4491,N_4144,N_4232);
nand U4492 (N_4492,N_4065,N_4318);
nand U4493 (N_4493,N_3816,N_3834);
xor U4494 (N_4494,N_4156,N_3924);
and U4495 (N_4495,N_3889,N_3949);
or U4496 (N_4496,N_4358,N_4313);
nand U4497 (N_4497,N_3860,N_3818);
or U4498 (N_4498,N_4056,N_3824);
and U4499 (N_4499,N_4120,N_3959);
nand U4500 (N_4500,N_3897,N_4190);
nor U4501 (N_4501,N_4153,N_4194);
xnor U4502 (N_4502,N_4372,N_4104);
xor U4503 (N_4503,N_4308,N_4008);
xnor U4504 (N_4504,N_3926,N_3971);
xnor U4505 (N_4505,N_4038,N_4091);
nor U4506 (N_4506,N_4284,N_3934);
or U4507 (N_4507,N_3792,N_4005);
nand U4508 (N_4508,N_4217,N_3881);
xor U4509 (N_4509,N_3783,N_4012);
and U4510 (N_4510,N_3822,N_4185);
or U4511 (N_4511,N_4173,N_4040);
nand U4512 (N_4512,N_4176,N_3954);
or U4513 (N_4513,N_4063,N_3845);
xor U4514 (N_4514,N_4148,N_4225);
and U4515 (N_4515,N_3967,N_3946);
and U4516 (N_4516,N_3991,N_3930);
xor U4517 (N_4517,N_4162,N_3780);
nand U4518 (N_4518,N_4324,N_4347);
nand U4519 (N_4519,N_3875,N_4220);
nor U4520 (N_4520,N_4110,N_3957);
and U4521 (N_4521,N_4259,N_4351);
and U4522 (N_4522,N_3842,N_4199);
and U4523 (N_4523,N_3851,N_4211);
xnor U4524 (N_4524,N_4118,N_4274);
nor U4525 (N_4525,N_4112,N_4158);
or U4526 (N_4526,N_4202,N_4214);
xor U4527 (N_4527,N_4264,N_4085);
nand U4528 (N_4528,N_3863,N_3790);
nand U4529 (N_4529,N_4142,N_4031);
nor U4530 (N_4530,N_4090,N_3799);
and U4531 (N_4531,N_3885,N_4266);
or U4532 (N_4532,N_4010,N_4238);
xnor U4533 (N_4533,N_4193,N_4100);
nand U4534 (N_4534,N_4265,N_4105);
nor U4535 (N_4535,N_3791,N_3973);
nor U4536 (N_4536,N_4177,N_4326);
nor U4537 (N_4537,N_4159,N_4088);
xor U4538 (N_4538,N_3903,N_4026);
nor U4539 (N_4539,N_3896,N_3886);
xor U4540 (N_4540,N_4021,N_4175);
or U4541 (N_4541,N_3864,N_4061);
xor U4542 (N_4542,N_4302,N_4179);
and U4543 (N_4543,N_4371,N_3876);
or U4544 (N_4544,N_4288,N_4205);
nor U4545 (N_4545,N_4121,N_4075);
nor U4546 (N_4546,N_4203,N_3826);
nand U4547 (N_4547,N_4262,N_3872);
nor U4548 (N_4548,N_4078,N_3980);
and U4549 (N_4549,N_3981,N_4267);
xnor U4550 (N_4550,N_4207,N_3844);
nand U4551 (N_4551,N_4073,N_4034);
and U4552 (N_4552,N_4007,N_4130);
nor U4553 (N_4553,N_3858,N_4189);
and U4554 (N_4554,N_4222,N_4166);
nor U4555 (N_4555,N_3972,N_3890);
nor U4556 (N_4556,N_4279,N_4363);
and U4557 (N_4557,N_3835,N_4086);
nand U4558 (N_4558,N_4074,N_4346);
xnor U4559 (N_4559,N_3952,N_3802);
nand U4560 (N_4560,N_4229,N_4042);
nor U4561 (N_4561,N_4128,N_4361);
or U4562 (N_4562,N_3938,N_4022);
and U4563 (N_4563,N_4278,N_4068);
or U4564 (N_4564,N_3968,N_3914);
or U4565 (N_4565,N_4154,N_4164);
and U4566 (N_4566,N_4106,N_3782);
xor U4567 (N_4567,N_3806,N_4325);
or U4568 (N_4568,N_4336,N_4001);
or U4569 (N_4569,N_3918,N_4138);
or U4570 (N_4570,N_3947,N_3892);
or U4571 (N_4571,N_4373,N_4300);
xor U4572 (N_4572,N_4258,N_3804);
nor U4573 (N_4573,N_4263,N_3755);
nand U4574 (N_4574,N_4163,N_4369);
nor U4575 (N_4575,N_3884,N_3798);
xor U4576 (N_4576,N_4256,N_3877);
and U4577 (N_4577,N_4215,N_3883);
and U4578 (N_4578,N_4171,N_3777);
or U4579 (N_4579,N_4269,N_3839);
nand U4580 (N_4580,N_3882,N_4013);
and U4581 (N_4581,N_3937,N_4079);
or U4582 (N_4582,N_4224,N_4114);
xnor U4583 (N_4583,N_3812,N_4066);
xnor U4584 (N_4584,N_4157,N_4252);
or U4585 (N_4585,N_3776,N_4096);
xor U4586 (N_4586,N_4076,N_4374);
xnor U4587 (N_4587,N_4191,N_3803);
and U4588 (N_4588,N_4321,N_4098);
and U4589 (N_4589,N_3764,N_3757);
or U4590 (N_4590,N_4290,N_4338);
or U4591 (N_4591,N_3763,N_3787);
or U4592 (N_4592,N_4095,N_4025);
and U4593 (N_4593,N_4233,N_3891);
xnor U4594 (N_4594,N_3942,N_3911);
nand U4595 (N_4595,N_3956,N_4301);
nand U4596 (N_4596,N_4117,N_4311);
or U4597 (N_4597,N_4273,N_4029);
xor U4598 (N_4598,N_4035,N_3965);
or U4599 (N_4599,N_4141,N_3825);
nand U4600 (N_4600,N_3796,N_4281);
and U4601 (N_4601,N_3939,N_4116);
nand U4602 (N_4602,N_3868,N_3944);
nor U4603 (N_4603,N_3878,N_3927);
nor U4604 (N_4604,N_3775,N_3871);
nand U4605 (N_4605,N_3808,N_4319);
and U4606 (N_4606,N_4082,N_4307);
xor U4607 (N_4607,N_4016,N_3998);
and U4608 (N_4608,N_4057,N_3987);
or U4609 (N_4609,N_4227,N_4097);
nor U4610 (N_4610,N_4002,N_4223);
and U4611 (N_4611,N_3964,N_4282);
or U4612 (N_4612,N_4070,N_4270);
nand U4613 (N_4613,N_4103,N_3813);
xnor U4614 (N_4614,N_4219,N_3919);
xnor U4615 (N_4615,N_3846,N_3906);
or U4616 (N_4616,N_4339,N_4197);
xor U4617 (N_4617,N_3932,N_3866);
nand U4618 (N_4618,N_3785,N_3772);
nor U4619 (N_4619,N_4246,N_4182);
and U4620 (N_4620,N_3765,N_4028);
xnor U4621 (N_4621,N_3828,N_4180);
xnor U4622 (N_4622,N_4276,N_4309);
nand U4623 (N_4623,N_3970,N_4196);
nand U4624 (N_4624,N_3827,N_3759);
nand U4625 (N_4625,N_4344,N_4249);
or U4626 (N_4626,N_4119,N_3925);
or U4627 (N_4627,N_3908,N_4133);
nand U4628 (N_4628,N_4048,N_4331);
and U4629 (N_4629,N_3920,N_4200);
or U4630 (N_4630,N_4368,N_4018);
nor U4631 (N_4631,N_4287,N_4054);
and U4632 (N_4632,N_3915,N_4247);
nor U4633 (N_4633,N_3770,N_4228);
nor U4634 (N_4634,N_4149,N_3829);
and U4635 (N_4635,N_4213,N_3807);
nand U4636 (N_4636,N_4275,N_3800);
nand U4637 (N_4637,N_3988,N_3843);
nand U4638 (N_4638,N_3997,N_4299);
or U4639 (N_4639,N_4172,N_4014);
nand U4640 (N_4640,N_3820,N_4135);
xor U4641 (N_4641,N_4129,N_4201);
nand U4642 (N_4642,N_3902,N_3958);
nand U4643 (N_4643,N_3895,N_4000);
and U4644 (N_4644,N_3761,N_4060);
nor U4645 (N_4645,N_4107,N_4237);
or U4646 (N_4646,N_3948,N_4315);
nand U4647 (N_4647,N_3916,N_4362);
xor U4648 (N_4648,N_3810,N_3922);
or U4649 (N_4649,N_3819,N_4366);
nor U4650 (N_4650,N_3811,N_4280);
and U4651 (N_4651,N_4292,N_3995);
or U4652 (N_4652,N_3923,N_3880);
nor U4653 (N_4653,N_4058,N_3784);
xor U4654 (N_4654,N_3752,N_3771);
and U4655 (N_4655,N_4327,N_3912);
nand U4656 (N_4656,N_3754,N_3907);
or U4657 (N_4657,N_3943,N_3941);
nor U4658 (N_4658,N_4364,N_3786);
xnor U4659 (N_4659,N_4240,N_4140);
and U4660 (N_4660,N_4101,N_4342);
and U4661 (N_4661,N_4015,N_3779);
nand U4662 (N_4662,N_4243,N_3960);
and U4663 (N_4663,N_4370,N_4011);
xnor U4664 (N_4664,N_3955,N_4009);
nand U4665 (N_4665,N_4349,N_4306);
xor U4666 (N_4666,N_4250,N_3917);
and U4667 (N_4667,N_3849,N_4239);
and U4668 (N_4668,N_4113,N_4310);
nor U4669 (N_4669,N_4174,N_3893);
xor U4670 (N_4670,N_4033,N_4043);
or U4671 (N_4671,N_3898,N_3873);
nor U4672 (N_4672,N_4251,N_4049);
nor U4673 (N_4673,N_4235,N_4039);
or U4674 (N_4674,N_3767,N_4333);
nor U4675 (N_4675,N_3815,N_4178);
nand U4676 (N_4676,N_3837,N_4359);
and U4677 (N_4677,N_3847,N_4195);
and U4678 (N_4678,N_4111,N_3978);
nand U4679 (N_4679,N_3832,N_4234);
or U4680 (N_4680,N_3992,N_4071);
and U4681 (N_4681,N_4152,N_3999);
xor U4682 (N_4682,N_3940,N_3986);
and U4683 (N_4683,N_4231,N_4167);
nor U4684 (N_4684,N_3963,N_4184);
and U4685 (N_4685,N_4186,N_4317);
nand U4686 (N_4686,N_4132,N_4168);
nor U4687 (N_4687,N_4099,N_3867);
and U4688 (N_4688,N_3944,N_3908);
xor U4689 (N_4689,N_3816,N_4206);
nor U4690 (N_4690,N_3831,N_3835);
nand U4691 (N_4691,N_4134,N_4119);
xor U4692 (N_4692,N_3944,N_4026);
and U4693 (N_4693,N_4261,N_4198);
xor U4694 (N_4694,N_3929,N_4040);
xnor U4695 (N_4695,N_3800,N_4053);
and U4696 (N_4696,N_3803,N_4225);
and U4697 (N_4697,N_4071,N_4077);
nor U4698 (N_4698,N_3925,N_3913);
nor U4699 (N_4699,N_4015,N_4227);
nand U4700 (N_4700,N_4097,N_3803);
nand U4701 (N_4701,N_4277,N_4139);
xor U4702 (N_4702,N_3767,N_4257);
nand U4703 (N_4703,N_4007,N_4297);
and U4704 (N_4704,N_3774,N_4123);
nand U4705 (N_4705,N_4031,N_3787);
nand U4706 (N_4706,N_3892,N_3972);
or U4707 (N_4707,N_4209,N_4235);
and U4708 (N_4708,N_3877,N_3908);
or U4709 (N_4709,N_4013,N_4104);
xor U4710 (N_4710,N_4006,N_3986);
and U4711 (N_4711,N_4293,N_4351);
and U4712 (N_4712,N_3896,N_4234);
xnor U4713 (N_4713,N_3899,N_4201);
xnor U4714 (N_4714,N_4116,N_4075);
xnor U4715 (N_4715,N_3955,N_4032);
nor U4716 (N_4716,N_4352,N_4056);
and U4717 (N_4717,N_4215,N_3914);
or U4718 (N_4718,N_4082,N_4207);
and U4719 (N_4719,N_4315,N_3870);
nor U4720 (N_4720,N_3799,N_3959);
nor U4721 (N_4721,N_4033,N_4235);
nand U4722 (N_4722,N_3942,N_4003);
and U4723 (N_4723,N_3869,N_4086);
nand U4724 (N_4724,N_3913,N_3843);
nor U4725 (N_4725,N_4031,N_3839);
and U4726 (N_4726,N_3863,N_3782);
nand U4727 (N_4727,N_4090,N_4239);
xor U4728 (N_4728,N_3850,N_3806);
xnor U4729 (N_4729,N_4310,N_4361);
xor U4730 (N_4730,N_4219,N_3920);
nand U4731 (N_4731,N_3922,N_4114);
or U4732 (N_4732,N_3925,N_4138);
nand U4733 (N_4733,N_3971,N_3959);
xor U4734 (N_4734,N_4179,N_3858);
nand U4735 (N_4735,N_4045,N_4154);
xnor U4736 (N_4736,N_4099,N_3841);
xor U4737 (N_4737,N_3943,N_4164);
and U4738 (N_4738,N_3951,N_4312);
xnor U4739 (N_4739,N_3921,N_3942);
nand U4740 (N_4740,N_4172,N_4155);
nor U4741 (N_4741,N_4087,N_4217);
nand U4742 (N_4742,N_4330,N_4277);
xnor U4743 (N_4743,N_3778,N_4330);
or U4744 (N_4744,N_4105,N_3793);
xnor U4745 (N_4745,N_3864,N_4029);
and U4746 (N_4746,N_3953,N_4191);
nand U4747 (N_4747,N_3846,N_3868);
nand U4748 (N_4748,N_4013,N_4030);
or U4749 (N_4749,N_4331,N_3930);
xor U4750 (N_4750,N_4367,N_4095);
xnor U4751 (N_4751,N_3780,N_4111);
and U4752 (N_4752,N_4284,N_3801);
nor U4753 (N_4753,N_4367,N_3911);
nand U4754 (N_4754,N_4110,N_3792);
nor U4755 (N_4755,N_3896,N_4032);
nor U4756 (N_4756,N_4129,N_3838);
xnor U4757 (N_4757,N_4099,N_3992);
nor U4758 (N_4758,N_4010,N_4206);
or U4759 (N_4759,N_3892,N_4237);
nor U4760 (N_4760,N_4054,N_3856);
and U4761 (N_4761,N_3782,N_3961);
nand U4762 (N_4762,N_4241,N_3868);
nand U4763 (N_4763,N_3889,N_4124);
nand U4764 (N_4764,N_3933,N_4032);
or U4765 (N_4765,N_3767,N_3830);
or U4766 (N_4766,N_3940,N_4338);
or U4767 (N_4767,N_4218,N_4270);
or U4768 (N_4768,N_4293,N_4031);
and U4769 (N_4769,N_4340,N_4165);
or U4770 (N_4770,N_4173,N_3913);
xor U4771 (N_4771,N_3949,N_3792);
and U4772 (N_4772,N_4317,N_4090);
and U4773 (N_4773,N_4257,N_3911);
or U4774 (N_4774,N_4310,N_4120);
xor U4775 (N_4775,N_3922,N_4039);
xnor U4776 (N_4776,N_3928,N_4054);
xnor U4777 (N_4777,N_4258,N_3987);
nand U4778 (N_4778,N_4153,N_3906);
nand U4779 (N_4779,N_4157,N_3806);
nand U4780 (N_4780,N_4335,N_4148);
and U4781 (N_4781,N_4056,N_4100);
and U4782 (N_4782,N_4280,N_4372);
nor U4783 (N_4783,N_3765,N_4291);
nand U4784 (N_4784,N_4017,N_4037);
or U4785 (N_4785,N_4053,N_3765);
nor U4786 (N_4786,N_3894,N_3897);
and U4787 (N_4787,N_4175,N_4265);
and U4788 (N_4788,N_3952,N_4180);
and U4789 (N_4789,N_4341,N_4293);
nor U4790 (N_4790,N_4117,N_4280);
xnor U4791 (N_4791,N_4039,N_4360);
and U4792 (N_4792,N_3947,N_3899);
or U4793 (N_4793,N_4097,N_3999);
nor U4794 (N_4794,N_3808,N_4083);
or U4795 (N_4795,N_3774,N_4105);
nor U4796 (N_4796,N_4078,N_4076);
nor U4797 (N_4797,N_3868,N_3777);
xnor U4798 (N_4798,N_3760,N_3999);
or U4799 (N_4799,N_3933,N_4298);
or U4800 (N_4800,N_3926,N_3835);
nor U4801 (N_4801,N_3875,N_3829);
nor U4802 (N_4802,N_3989,N_3887);
nand U4803 (N_4803,N_4228,N_4357);
xnor U4804 (N_4804,N_3917,N_4153);
and U4805 (N_4805,N_3980,N_4089);
xnor U4806 (N_4806,N_3787,N_4210);
nor U4807 (N_4807,N_4040,N_4331);
nor U4808 (N_4808,N_4163,N_4320);
and U4809 (N_4809,N_4051,N_3866);
nor U4810 (N_4810,N_3963,N_3877);
and U4811 (N_4811,N_3862,N_4060);
nor U4812 (N_4812,N_4157,N_3981);
nor U4813 (N_4813,N_3947,N_3837);
nand U4814 (N_4814,N_3820,N_3857);
nand U4815 (N_4815,N_4224,N_3780);
and U4816 (N_4816,N_4071,N_4057);
nor U4817 (N_4817,N_4009,N_4035);
or U4818 (N_4818,N_4140,N_4266);
and U4819 (N_4819,N_3777,N_3756);
and U4820 (N_4820,N_3961,N_3977);
nand U4821 (N_4821,N_3837,N_4155);
xnor U4822 (N_4822,N_3857,N_3987);
or U4823 (N_4823,N_4152,N_4177);
and U4824 (N_4824,N_4195,N_4365);
or U4825 (N_4825,N_4091,N_3942);
xor U4826 (N_4826,N_3945,N_4096);
nand U4827 (N_4827,N_4089,N_4165);
nand U4828 (N_4828,N_4020,N_4314);
and U4829 (N_4829,N_3996,N_4304);
nor U4830 (N_4830,N_4292,N_3889);
xnor U4831 (N_4831,N_3840,N_4135);
and U4832 (N_4832,N_4321,N_3953);
or U4833 (N_4833,N_3881,N_3763);
nor U4834 (N_4834,N_3902,N_4158);
and U4835 (N_4835,N_3778,N_4313);
nor U4836 (N_4836,N_4137,N_4155);
or U4837 (N_4837,N_4056,N_4340);
or U4838 (N_4838,N_4255,N_4038);
and U4839 (N_4839,N_4284,N_4088);
xnor U4840 (N_4840,N_4073,N_3804);
nor U4841 (N_4841,N_4162,N_4077);
nor U4842 (N_4842,N_3775,N_4016);
nand U4843 (N_4843,N_4174,N_3808);
or U4844 (N_4844,N_4106,N_3880);
or U4845 (N_4845,N_4196,N_4181);
or U4846 (N_4846,N_4365,N_3754);
and U4847 (N_4847,N_4349,N_3953);
or U4848 (N_4848,N_3767,N_3775);
or U4849 (N_4849,N_3799,N_4323);
or U4850 (N_4850,N_4100,N_4006);
and U4851 (N_4851,N_3946,N_4342);
nor U4852 (N_4852,N_4083,N_3838);
nor U4853 (N_4853,N_4149,N_3921);
or U4854 (N_4854,N_4108,N_4049);
nor U4855 (N_4855,N_4336,N_4084);
xor U4856 (N_4856,N_3888,N_4024);
or U4857 (N_4857,N_4312,N_4145);
nand U4858 (N_4858,N_4101,N_4240);
nor U4859 (N_4859,N_3946,N_4198);
xnor U4860 (N_4860,N_4115,N_4138);
nor U4861 (N_4861,N_3891,N_3982);
or U4862 (N_4862,N_4183,N_3978);
nand U4863 (N_4863,N_4132,N_4257);
or U4864 (N_4864,N_4016,N_4208);
nor U4865 (N_4865,N_3832,N_4289);
xor U4866 (N_4866,N_3756,N_4362);
xor U4867 (N_4867,N_4250,N_3827);
nand U4868 (N_4868,N_3947,N_4085);
nand U4869 (N_4869,N_3865,N_4227);
and U4870 (N_4870,N_3770,N_3906);
or U4871 (N_4871,N_3858,N_3978);
or U4872 (N_4872,N_4096,N_3973);
nor U4873 (N_4873,N_3866,N_4266);
nor U4874 (N_4874,N_4278,N_4093);
nand U4875 (N_4875,N_3758,N_3919);
xnor U4876 (N_4876,N_3887,N_3850);
or U4877 (N_4877,N_4111,N_3879);
or U4878 (N_4878,N_4250,N_4358);
xnor U4879 (N_4879,N_4059,N_4153);
or U4880 (N_4880,N_3888,N_4124);
and U4881 (N_4881,N_4259,N_4165);
nand U4882 (N_4882,N_4342,N_4001);
and U4883 (N_4883,N_4123,N_4140);
and U4884 (N_4884,N_4037,N_3790);
nor U4885 (N_4885,N_4306,N_3871);
and U4886 (N_4886,N_3998,N_3758);
and U4887 (N_4887,N_4032,N_3776);
xnor U4888 (N_4888,N_3920,N_4280);
nand U4889 (N_4889,N_3756,N_3953);
xnor U4890 (N_4890,N_4009,N_4166);
nor U4891 (N_4891,N_3985,N_4292);
xnor U4892 (N_4892,N_4147,N_3833);
and U4893 (N_4893,N_4148,N_4057);
or U4894 (N_4894,N_3915,N_4110);
and U4895 (N_4895,N_4319,N_3765);
xor U4896 (N_4896,N_4112,N_4146);
and U4897 (N_4897,N_4067,N_4098);
nor U4898 (N_4898,N_4245,N_4352);
nor U4899 (N_4899,N_3880,N_3755);
or U4900 (N_4900,N_4362,N_3794);
nor U4901 (N_4901,N_4013,N_3807);
or U4902 (N_4902,N_4224,N_4159);
and U4903 (N_4903,N_3954,N_3866);
xnor U4904 (N_4904,N_4270,N_4054);
xnor U4905 (N_4905,N_4326,N_4259);
xnor U4906 (N_4906,N_3813,N_4096);
nand U4907 (N_4907,N_4084,N_4321);
and U4908 (N_4908,N_4044,N_4080);
nand U4909 (N_4909,N_4039,N_4052);
nor U4910 (N_4910,N_4161,N_4083);
and U4911 (N_4911,N_4241,N_4068);
and U4912 (N_4912,N_3911,N_4074);
and U4913 (N_4913,N_3900,N_3905);
xor U4914 (N_4914,N_3864,N_4251);
nand U4915 (N_4915,N_4217,N_4089);
and U4916 (N_4916,N_4189,N_4053);
nand U4917 (N_4917,N_4286,N_3773);
nand U4918 (N_4918,N_3868,N_3919);
nand U4919 (N_4919,N_3797,N_3876);
or U4920 (N_4920,N_4347,N_3850);
and U4921 (N_4921,N_3996,N_3872);
nand U4922 (N_4922,N_4260,N_3925);
or U4923 (N_4923,N_4204,N_4297);
xor U4924 (N_4924,N_4244,N_4025);
xor U4925 (N_4925,N_3934,N_4370);
and U4926 (N_4926,N_3806,N_3807);
nor U4927 (N_4927,N_4225,N_4302);
nor U4928 (N_4928,N_4065,N_3893);
xnor U4929 (N_4929,N_3849,N_3858);
nand U4930 (N_4930,N_4215,N_3869);
and U4931 (N_4931,N_3794,N_4130);
and U4932 (N_4932,N_4368,N_4309);
and U4933 (N_4933,N_4197,N_4080);
xnor U4934 (N_4934,N_4085,N_4356);
nor U4935 (N_4935,N_4167,N_3888);
nor U4936 (N_4936,N_4146,N_3944);
and U4937 (N_4937,N_4035,N_4194);
and U4938 (N_4938,N_4182,N_4211);
nor U4939 (N_4939,N_3884,N_3791);
xor U4940 (N_4940,N_3819,N_3884);
nor U4941 (N_4941,N_4155,N_4060);
and U4942 (N_4942,N_3942,N_4353);
nand U4943 (N_4943,N_4329,N_4001);
nor U4944 (N_4944,N_3854,N_4231);
nand U4945 (N_4945,N_3870,N_4236);
xor U4946 (N_4946,N_4292,N_3950);
or U4947 (N_4947,N_4329,N_4222);
xor U4948 (N_4948,N_4139,N_3908);
xnor U4949 (N_4949,N_4312,N_3845);
or U4950 (N_4950,N_4156,N_4366);
nor U4951 (N_4951,N_4103,N_3802);
xor U4952 (N_4952,N_4044,N_3952);
nor U4953 (N_4953,N_4139,N_3766);
and U4954 (N_4954,N_4021,N_3850);
and U4955 (N_4955,N_4303,N_4202);
nand U4956 (N_4956,N_4351,N_4198);
xor U4957 (N_4957,N_4298,N_4040);
nand U4958 (N_4958,N_4302,N_3815);
nor U4959 (N_4959,N_4076,N_3896);
nand U4960 (N_4960,N_4130,N_3945);
or U4961 (N_4961,N_4307,N_4242);
or U4962 (N_4962,N_3784,N_4204);
nor U4963 (N_4963,N_3969,N_4043);
nor U4964 (N_4964,N_4249,N_4154);
nor U4965 (N_4965,N_4333,N_4276);
nand U4966 (N_4966,N_4131,N_3936);
or U4967 (N_4967,N_4017,N_4368);
and U4968 (N_4968,N_4367,N_3926);
and U4969 (N_4969,N_4026,N_4221);
nand U4970 (N_4970,N_3997,N_4266);
nand U4971 (N_4971,N_3849,N_3977);
xor U4972 (N_4972,N_4309,N_3820);
xnor U4973 (N_4973,N_4072,N_3891);
and U4974 (N_4974,N_3959,N_4199);
or U4975 (N_4975,N_3948,N_4121);
or U4976 (N_4976,N_4286,N_3898);
or U4977 (N_4977,N_4273,N_3991);
and U4978 (N_4978,N_3817,N_4091);
nor U4979 (N_4979,N_4252,N_3916);
xor U4980 (N_4980,N_3997,N_4098);
nand U4981 (N_4981,N_4213,N_4254);
and U4982 (N_4982,N_3813,N_4240);
nand U4983 (N_4983,N_4224,N_4088);
and U4984 (N_4984,N_4004,N_4001);
nand U4985 (N_4985,N_3965,N_4336);
xor U4986 (N_4986,N_4137,N_4371);
nand U4987 (N_4987,N_4294,N_4250);
nor U4988 (N_4988,N_4187,N_3994);
xnor U4989 (N_4989,N_4324,N_4197);
or U4990 (N_4990,N_4366,N_3801);
nor U4991 (N_4991,N_4064,N_4059);
xnor U4992 (N_4992,N_3758,N_4103);
and U4993 (N_4993,N_3964,N_4269);
xnor U4994 (N_4994,N_3896,N_3969);
nor U4995 (N_4995,N_3756,N_3791);
nor U4996 (N_4996,N_4209,N_4113);
xnor U4997 (N_4997,N_3955,N_3840);
or U4998 (N_4998,N_4346,N_4352);
nor U4999 (N_4999,N_4237,N_3894);
and U5000 (N_5000,N_4397,N_4958);
or U5001 (N_5001,N_4499,N_4393);
nor U5002 (N_5002,N_4480,N_4975);
xnor U5003 (N_5003,N_4651,N_4999);
and U5004 (N_5004,N_4802,N_4494);
nor U5005 (N_5005,N_4929,N_4609);
nand U5006 (N_5006,N_4948,N_4508);
nor U5007 (N_5007,N_4517,N_4427);
nor U5008 (N_5008,N_4390,N_4557);
and U5009 (N_5009,N_4669,N_4799);
xor U5010 (N_5010,N_4811,N_4420);
or U5011 (N_5011,N_4518,N_4689);
nand U5012 (N_5012,N_4566,N_4759);
nor U5013 (N_5013,N_4906,N_4626);
nand U5014 (N_5014,N_4588,N_4946);
xnor U5015 (N_5015,N_4475,N_4467);
or U5016 (N_5016,N_4389,N_4398);
or U5017 (N_5017,N_4732,N_4970);
or U5018 (N_5018,N_4431,N_4784);
nand U5019 (N_5019,N_4548,N_4536);
nor U5020 (N_5020,N_4856,N_4954);
or U5021 (N_5021,N_4823,N_4641);
or U5022 (N_5022,N_4919,N_4449);
nand U5023 (N_5023,N_4715,N_4845);
xnor U5024 (N_5024,N_4493,N_4640);
xor U5025 (N_5025,N_4525,N_4439);
xor U5026 (N_5026,N_4926,N_4468);
or U5027 (N_5027,N_4540,N_4704);
or U5028 (N_5028,N_4567,N_4619);
nand U5029 (N_5029,N_4874,N_4624);
or U5030 (N_5030,N_4996,N_4966);
nor U5031 (N_5031,N_4591,N_4697);
nand U5032 (N_5032,N_4809,N_4713);
and U5033 (N_5033,N_4978,N_4711);
nor U5034 (N_5034,N_4558,N_4739);
or U5035 (N_5035,N_4406,N_4812);
and U5036 (N_5036,N_4514,N_4719);
nor U5037 (N_5037,N_4531,N_4457);
nor U5038 (N_5038,N_4944,N_4528);
nand U5039 (N_5039,N_4997,N_4498);
or U5040 (N_5040,N_4887,N_4601);
nand U5041 (N_5041,N_4962,N_4898);
or U5042 (N_5042,N_4648,N_4775);
nor U5043 (N_5043,N_4578,N_4888);
nand U5044 (N_5044,N_4864,N_4741);
nor U5045 (N_5045,N_4532,N_4871);
xnor U5046 (N_5046,N_4671,N_4804);
or U5047 (N_5047,N_4838,N_4496);
xnor U5048 (N_5048,N_4527,N_4501);
nand U5049 (N_5049,N_4524,N_4989);
and U5050 (N_5050,N_4375,N_4407);
and U5051 (N_5051,N_4597,N_4947);
and U5052 (N_5052,N_4585,N_4754);
nand U5053 (N_5053,N_4894,N_4632);
nand U5054 (N_5054,N_4502,N_4990);
nand U5055 (N_5055,N_4429,N_4852);
xnor U5056 (N_5056,N_4665,N_4376);
and U5057 (N_5057,N_4684,N_4638);
nor U5058 (N_5058,N_4676,N_4963);
nand U5059 (N_5059,N_4967,N_4628);
xnor U5060 (N_5060,N_4829,N_4593);
or U5061 (N_5061,N_4603,N_4629);
or U5062 (N_5062,N_4916,N_4780);
nand U5063 (N_5063,N_4483,N_4938);
nand U5064 (N_5064,N_4452,N_4981);
and U5065 (N_5065,N_4659,N_4773);
and U5066 (N_5066,N_4965,N_4700);
nand U5067 (N_5067,N_4830,N_4824);
and U5068 (N_5068,N_4918,N_4458);
nand U5069 (N_5069,N_4788,N_4821);
nor U5070 (N_5070,N_4466,N_4396);
and U5071 (N_5071,N_4696,N_4504);
xor U5072 (N_5072,N_4599,N_4520);
and U5073 (N_5073,N_4644,N_4589);
nand U5074 (N_5074,N_4403,N_4728);
nor U5075 (N_5075,N_4855,N_4955);
and U5076 (N_5076,N_4418,N_4833);
and U5077 (N_5077,N_4616,N_4455);
nand U5078 (N_5078,N_4622,N_4596);
nand U5079 (N_5079,N_4826,N_4819);
or U5080 (N_5080,N_4915,N_4565);
nand U5081 (N_5081,N_4464,N_4760);
nand U5082 (N_5082,N_4986,N_4988);
or U5083 (N_5083,N_4571,N_4649);
xor U5084 (N_5084,N_4974,N_4613);
or U5085 (N_5085,N_4408,N_4801);
nand U5086 (N_5086,N_4952,N_4860);
xor U5087 (N_5087,N_4712,N_4994);
xnor U5088 (N_5088,N_4905,N_4647);
or U5089 (N_5089,N_4383,N_4580);
xor U5090 (N_5090,N_4459,N_4507);
and U5091 (N_5091,N_4949,N_4983);
or U5092 (N_5092,N_4576,N_4738);
or U5093 (N_5093,N_4512,N_4409);
or U5094 (N_5094,N_4973,N_4932);
nand U5095 (N_5095,N_4476,N_4951);
nor U5096 (N_5096,N_4847,N_4904);
nor U5097 (N_5097,N_4834,N_4831);
xnor U5098 (N_5098,N_4980,N_4652);
xor U5099 (N_5099,N_4562,N_4998);
and U5100 (N_5100,N_4426,N_4846);
nand U5101 (N_5101,N_4914,N_4755);
or U5102 (N_5102,N_4683,N_4432);
or U5103 (N_5103,N_4423,N_4937);
and U5104 (N_5104,N_4816,N_4634);
or U5105 (N_5105,N_4556,N_4579);
or U5106 (N_5106,N_4515,N_4768);
or U5107 (N_5107,N_4893,N_4382);
nand U5108 (N_5108,N_4810,N_4699);
and U5109 (N_5109,N_4896,N_4487);
or U5110 (N_5110,N_4884,N_4569);
nand U5111 (N_5111,N_4796,N_4471);
nor U5112 (N_5112,N_4542,N_4680);
xor U5113 (N_5113,N_4503,N_4931);
nor U5114 (N_5114,N_4960,N_4749);
and U5115 (N_5115,N_4943,N_4460);
or U5116 (N_5116,N_4767,N_4379);
and U5117 (N_5117,N_4706,N_4900);
and U5118 (N_5118,N_4993,N_4545);
xnor U5119 (N_5119,N_4882,N_4798);
nor U5120 (N_5120,N_4443,N_4587);
and U5121 (N_5121,N_4869,N_4463);
xor U5122 (N_5122,N_4940,N_4674);
or U5123 (N_5123,N_4698,N_4901);
or U5124 (N_5124,N_4912,N_4839);
nand U5125 (N_5125,N_4481,N_4703);
or U5126 (N_5126,N_4633,N_4752);
nand U5127 (N_5127,N_4777,N_4691);
and U5128 (N_5128,N_4727,N_4465);
and U5129 (N_5129,N_4662,N_4484);
nor U5130 (N_5130,N_4522,N_4645);
nand U5131 (N_5131,N_4794,N_4664);
nor U5132 (N_5132,N_4737,N_4836);
nor U5133 (N_5133,N_4422,N_4708);
or U5134 (N_5134,N_4440,N_4730);
nor U5135 (N_5135,N_4497,N_4682);
nand U5136 (N_5136,N_4611,N_4681);
and U5137 (N_5137,N_4763,N_4987);
and U5138 (N_5138,N_4729,N_4656);
xor U5139 (N_5139,N_4957,N_4984);
or U5140 (N_5140,N_4550,N_4677);
nor U5141 (N_5141,N_4414,N_4654);
and U5142 (N_5142,N_4472,N_4885);
nor U5143 (N_5143,N_4400,N_4658);
nor U5144 (N_5144,N_4380,N_4535);
nand U5145 (N_5145,N_4892,N_4552);
and U5146 (N_5146,N_4621,N_4602);
nor U5147 (N_5147,N_4553,N_4735);
nand U5148 (N_5148,N_4485,N_4606);
xor U5149 (N_5149,N_4462,N_4724);
or U5150 (N_5150,N_4818,N_4491);
nor U5151 (N_5151,N_4897,N_4742);
and U5152 (N_5152,N_4620,N_4608);
or U5153 (N_5153,N_4586,N_4857);
nand U5154 (N_5154,N_4774,N_4843);
or U5155 (N_5155,N_4705,N_4961);
and U5156 (N_5156,N_4549,N_4631);
and U5157 (N_5157,N_4817,N_4436);
nand U5158 (N_5158,N_4559,N_4679);
or U5159 (N_5159,N_4433,N_4653);
or U5160 (N_5160,N_4663,N_4451);
nor U5161 (N_5161,N_4492,N_4863);
nor U5162 (N_5162,N_4934,N_4721);
and U5163 (N_5163,N_4404,N_4410);
nand U5164 (N_5164,N_4509,N_4820);
and U5165 (N_5165,N_4911,N_4908);
xnor U5166 (N_5166,N_4907,N_4537);
xnor U5167 (N_5167,N_4785,N_4544);
xor U5168 (N_5168,N_4861,N_4770);
and U5169 (N_5169,N_4746,N_4825);
nor U5170 (N_5170,N_4546,N_4758);
xor U5171 (N_5171,N_4902,N_4555);
and U5172 (N_5172,N_4995,N_4849);
nand U5173 (N_5173,N_4594,N_4604);
nand U5174 (N_5174,N_4625,N_4617);
nand U5175 (N_5175,N_4950,N_4793);
nand U5176 (N_5176,N_4572,N_4880);
nor U5177 (N_5177,N_4827,N_4969);
nand U5178 (N_5178,N_4800,N_4757);
or U5179 (N_5179,N_4766,N_4964);
nor U5180 (N_5180,N_4511,N_4387);
and U5181 (N_5181,N_4750,N_4392);
nand U5182 (N_5182,N_4636,N_4854);
or U5183 (N_5183,N_4521,N_4474);
nand U5184 (N_5184,N_4513,N_4769);
xor U5185 (N_5185,N_4385,N_4976);
or U5186 (N_5186,N_4787,N_4953);
nand U5187 (N_5187,N_4605,N_4442);
or U5188 (N_5188,N_4441,N_4672);
nand U5189 (N_5189,N_4828,N_4598);
nand U5190 (N_5190,N_4917,N_4670);
nor U5191 (N_5191,N_4384,N_4879);
nand U5192 (N_5192,N_4692,N_4437);
and U5193 (N_5193,N_4778,N_4607);
and U5194 (N_5194,N_4723,N_4920);
and U5195 (N_5195,N_4506,N_4667);
nor U5196 (N_5196,N_4790,N_4717);
nor U5197 (N_5197,N_4479,N_4386);
nor U5198 (N_5198,N_4642,N_4772);
and U5199 (N_5199,N_4878,N_4707);
xnor U5200 (N_5200,N_4614,N_4421);
nor U5201 (N_5201,N_4630,N_4941);
or U5202 (N_5202,N_4394,N_4564);
and U5203 (N_5203,N_4405,N_4968);
and U5204 (N_5204,N_4734,N_4618);
nand U5205 (N_5205,N_4922,N_4771);
nand U5206 (N_5206,N_4877,N_4971);
or U5207 (N_5207,N_4473,N_4858);
xnor U5208 (N_5208,N_4500,N_4600);
nor U5209 (N_5209,N_4875,N_4714);
xnor U5210 (N_5210,N_4701,N_4388);
xnor U5211 (N_5211,N_4891,N_4868);
nand U5212 (N_5212,N_4716,N_4985);
nand U5213 (N_5213,N_4853,N_4982);
or U5214 (N_5214,N_4581,N_4751);
and U5215 (N_5215,N_4563,N_4745);
and U5216 (N_5216,N_4806,N_4543);
nor U5217 (N_5217,N_4837,N_4428);
or U5218 (N_5218,N_4523,N_4844);
nor U5219 (N_5219,N_4972,N_4541);
nand U5220 (N_5220,N_4554,N_4813);
or U5221 (N_5221,N_4639,N_4687);
and U5222 (N_5222,N_4395,N_4903);
or U5223 (N_5223,N_4477,N_4446);
or U5224 (N_5224,N_4688,N_4765);
or U5225 (N_5225,N_4533,N_4534);
or U5226 (N_5226,N_4568,N_4740);
nor U5227 (N_5227,N_4538,N_4842);
or U5228 (N_5228,N_4661,N_4782);
xor U5229 (N_5229,N_4928,N_4482);
and U5230 (N_5230,N_4761,N_4822);
nand U5231 (N_5231,N_4425,N_4456);
xor U5232 (N_5232,N_4650,N_4519);
xnor U5233 (N_5233,N_4381,N_4490);
nand U5234 (N_5234,N_4870,N_4805);
nor U5235 (N_5235,N_4447,N_4709);
nand U5236 (N_5236,N_4574,N_4921);
or U5237 (N_5237,N_4377,N_4646);
nor U5238 (N_5238,N_4851,N_4694);
and U5239 (N_5239,N_4776,N_4469);
nor U5240 (N_5240,N_4505,N_4445);
or U5241 (N_5241,N_4733,N_4417);
xnor U5242 (N_5242,N_4979,N_4413);
nor U5243 (N_5243,N_4655,N_4551);
nand U5244 (N_5244,N_4668,N_4530);
and U5245 (N_5245,N_4575,N_4448);
and U5246 (N_5246,N_4726,N_4945);
xor U5247 (N_5247,N_4424,N_4850);
nor U5248 (N_5248,N_4781,N_4924);
nand U5249 (N_5249,N_4722,N_4675);
or U5250 (N_5250,N_4401,N_4872);
nor U5251 (N_5251,N_4873,N_4762);
and U5252 (N_5252,N_4444,N_4807);
nor U5253 (N_5253,N_4927,N_4415);
nor U5254 (N_5254,N_4378,N_4808);
and U5255 (N_5255,N_4595,N_4547);
nand U5256 (N_5256,N_4913,N_4859);
xor U5257 (N_5257,N_4584,N_4612);
xor U5258 (N_5258,N_4673,N_4747);
xor U5259 (N_5259,N_4789,N_4942);
nor U5260 (N_5260,N_4815,N_4610);
or U5261 (N_5261,N_4435,N_4695);
nor U5262 (N_5262,N_4450,N_4592);
nor U5263 (N_5263,N_4615,N_4489);
and U5264 (N_5264,N_4909,N_4453);
or U5265 (N_5265,N_4956,N_4560);
or U5266 (N_5266,N_4718,N_4582);
nand U5267 (N_5267,N_4570,N_4748);
nor U5268 (N_5268,N_4495,N_4529);
nor U5269 (N_5269,N_4992,N_4865);
xor U5270 (N_5270,N_4510,N_4725);
or U5271 (N_5271,N_4786,N_4889);
nand U5272 (N_5272,N_4840,N_4832);
and U5273 (N_5273,N_4895,N_4416);
nor U5274 (N_5274,N_4573,N_4890);
nand U5275 (N_5275,N_4881,N_4743);
xor U5276 (N_5276,N_4867,N_4666);
nand U5277 (N_5277,N_4470,N_4702);
nand U5278 (N_5278,N_4779,N_4577);
nor U5279 (N_5279,N_4991,N_4430);
or U5280 (N_5280,N_4933,N_4803);
nand U5281 (N_5281,N_4486,N_4936);
and U5282 (N_5282,N_4583,N_4693);
nor U5283 (N_5283,N_4848,N_4539);
nor U5284 (N_5284,N_4438,N_4883);
nand U5285 (N_5285,N_4930,N_4925);
or U5286 (N_5286,N_4678,N_4623);
nor U5287 (N_5287,N_4876,N_4686);
or U5288 (N_5288,N_4434,N_4411);
and U5289 (N_5289,N_4685,N_4764);
xor U5290 (N_5290,N_4454,N_4720);
nand U5291 (N_5291,N_4783,N_4590);
or U5292 (N_5292,N_4710,N_4660);
and U5293 (N_5293,N_4959,N_4795);
xor U5294 (N_5294,N_4835,N_4637);
xnor U5295 (N_5295,N_4814,N_4657);
or U5296 (N_5296,N_4797,N_4923);
nand U5297 (N_5297,N_4391,N_4412);
xor U5298 (N_5298,N_4402,N_4792);
nor U5299 (N_5299,N_4643,N_4753);
xnor U5300 (N_5300,N_4744,N_4526);
nor U5301 (N_5301,N_4935,N_4635);
nand U5302 (N_5302,N_4488,N_4866);
nor U5303 (N_5303,N_4939,N_4399);
xnor U5304 (N_5304,N_4862,N_4977);
nor U5305 (N_5305,N_4561,N_4731);
nor U5306 (N_5306,N_4690,N_4756);
nand U5307 (N_5307,N_4627,N_4516);
nand U5308 (N_5308,N_4886,N_4461);
nor U5309 (N_5309,N_4478,N_4899);
or U5310 (N_5310,N_4419,N_4841);
or U5311 (N_5311,N_4736,N_4910);
and U5312 (N_5312,N_4791,N_4616);
and U5313 (N_5313,N_4678,N_4931);
nand U5314 (N_5314,N_4744,N_4678);
or U5315 (N_5315,N_4620,N_4532);
nor U5316 (N_5316,N_4997,N_4400);
nand U5317 (N_5317,N_4949,N_4810);
or U5318 (N_5318,N_4536,N_4537);
or U5319 (N_5319,N_4913,N_4375);
nand U5320 (N_5320,N_4829,N_4934);
xnor U5321 (N_5321,N_4734,N_4820);
or U5322 (N_5322,N_4489,N_4569);
nand U5323 (N_5323,N_4854,N_4886);
or U5324 (N_5324,N_4858,N_4692);
xor U5325 (N_5325,N_4482,N_4927);
nor U5326 (N_5326,N_4421,N_4580);
nand U5327 (N_5327,N_4898,N_4668);
nand U5328 (N_5328,N_4455,N_4625);
and U5329 (N_5329,N_4519,N_4768);
or U5330 (N_5330,N_4479,N_4830);
nor U5331 (N_5331,N_4927,N_4470);
nand U5332 (N_5332,N_4460,N_4475);
xnor U5333 (N_5333,N_4821,N_4628);
nor U5334 (N_5334,N_4791,N_4628);
and U5335 (N_5335,N_4948,N_4673);
or U5336 (N_5336,N_4900,N_4564);
and U5337 (N_5337,N_4762,N_4715);
xnor U5338 (N_5338,N_4657,N_4768);
xnor U5339 (N_5339,N_4686,N_4765);
nor U5340 (N_5340,N_4715,N_4524);
xor U5341 (N_5341,N_4557,N_4655);
and U5342 (N_5342,N_4892,N_4711);
nand U5343 (N_5343,N_4835,N_4445);
or U5344 (N_5344,N_4821,N_4873);
or U5345 (N_5345,N_4668,N_4719);
nand U5346 (N_5346,N_4700,N_4667);
nor U5347 (N_5347,N_4761,N_4783);
or U5348 (N_5348,N_4655,N_4989);
and U5349 (N_5349,N_4900,N_4920);
xnor U5350 (N_5350,N_4745,N_4857);
and U5351 (N_5351,N_4720,N_4474);
xnor U5352 (N_5352,N_4720,N_4922);
and U5353 (N_5353,N_4558,N_4995);
or U5354 (N_5354,N_4658,N_4418);
or U5355 (N_5355,N_4731,N_4483);
or U5356 (N_5356,N_4632,N_4969);
nand U5357 (N_5357,N_4714,N_4609);
nor U5358 (N_5358,N_4375,N_4911);
nor U5359 (N_5359,N_4922,N_4696);
nand U5360 (N_5360,N_4535,N_4402);
and U5361 (N_5361,N_4467,N_4715);
nand U5362 (N_5362,N_4549,N_4838);
nor U5363 (N_5363,N_4473,N_4383);
nor U5364 (N_5364,N_4586,N_4498);
and U5365 (N_5365,N_4784,N_4406);
nand U5366 (N_5366,N_4463,N_4381);
and U5367 (N_5367,N_4446,N_4816);
nand U5368 (N_5368,N_4911,N_4941);
nand U5369 (N_5369,N_4518,N_4673);
or U5370 (N_5370,N_4887,N_4412);
xnor U5371 (N_5371,N_4412,N_4545);
or U5372 (N_5372,N_4780,N_4441);
xnor U5373 (N_5373,N_4833,N_4627);
nand U5374 (N_5374,N_4495,N_4856);
nor U5375 (N_5375,N_4435,N_4541);
xor U5376 (N_5376,N_4871,N_4569);
or U5377 (N_5377,N_4570,N_4404);
nand U5378 (N_5378,N_4752,N_4592);
or U5379 (N_5379,N_4469,N_4612);
nand U5380 (N_5380,N_4999,N_4521);
nand U5381 (N_5381,N_4580,N_4489);
xor U5382 (N_5382,N_4506,N_4484);
xnor U5383 (N_5383,N_4808,N_4819);
nor U5384 (N_5384,N_4560,N_4849);
and U5385 (N_5385,N_4532,N_4680);
xor U5386 (N_5386,N_4714,N_4673);
or U5387 (N_5387,N_4594,N_4743);
nor U5388 (N_5388,N_4464,N_4948);
xnor U5389 (N_5389,N_4817,N_4834);
and U5390 (N_5390,N_4625,N_4378);
xnor U5391 (N_5391,N_4430,N_4673);
nand U5392 (N_5392,N_4689,N_4663);
nand U5393 (N_5393,N_4605,N_4739);
or U5394 (N_5394,N_4470,N_4898);
nand U5395 (N_5395,N_4733,N_4579);
xnor U5396 (N_5396,N_4837,N_4875);
or U5397 (N_5397,N_4491,N_4435);
or U5398 (N_5398,N_4662,N_4672);
xor U5399 (N_5399,N_4632,N_4964);
nor U5400 (N_5400,N_4545,N_4804);
nor U5401 (N_5401,N_4861,N_4451);
nor U5402 (N_5402,N_4958,N_4979);
nand U5403 (N_5403,N_4865,N_4902);
nor U5404 (N_5404,N_4792,N_4701);
xnor U5405 (N_5405,N_4837,N_4911);
nand U5406 (N_5406,N_4512,N_4953);
nor U5407 (N_5407,N_4986,N_4905);
or U5408 (N_5408,N_4646,N_4964);
and U5409 (N_5409,N_4602,N_4791);
xor U5410 (N_5410,N_4849,N_4843);
xor U5411 (N_5411,N_4438,N_4700);
and U5412 (N_5412,N_4642,N_4552);
xnor U5413 (N_5413,N_4915,N_4519);
or U5414 (N_5414,N_4969,N_4823);
nor U5415 (N_5415,N_4410,N_4607);
or U5416 (N_5416,N_4991,N_4858);
nor U5417 (N_5417,N_4969,N_4950);
nand U5418 (N_5418,N_4463,N_4452);
or U5419 (N_5419,N_4885,N_4743);
nand U5420 (N_5420,N_4835,N_4650);
xnor U5421 (N_5421,N_4573,N_4701);
or U5422 (N_5422,N_4589,N_4416);
and U5423 (N_5423,N_4544,N_4430);
nand U5424 (N_5424,N_4501,N_4546);
nor U5425 (N_5425,N_4465,N_4940);
and U5426 (N_5426,N_4699,N_4541);
or U5427 (N_5427,N_4654,N_4930);
nand U5428 (N_5428,N_4815,N_4444);
xnor U5429 (N_5429,N_4688,N_4618);
or U5430 (N_5430,N_4879,N_4740);
xnor U5431 (N_5431,N_4857,N_4867);
nand U5432 (N_5432,N_4515,N_4981);
or U5433 (N_5433,N_4963,N_4738);
nand U5434 (N_5434,N_4634,N_4473);
xnor U5435 (N_5435,N_4453,N_4420);
nor U5436 (N_5436,N_4974,N_4778);
nand U5437 (N_5437,N_4686,N_4612);
nor U5438 (N_5438,N_4410,N_4840);
and U5439 (N_5439,N_4949,N_4724);
or U5440 (N_5440,N_4737,N_4850);
xnor U5441 (N_5441,N_4473,N_4454);
or U5442 (N_5442,N_4623,N_4408);
nand U5443 (N_5443,N_4726,N_4380);
nor U5444 (N_5444,N_4590,N_4812);
nor U5445 (N_5445,N_4410,N_4771);
nor U5446 (N_5446,N_4703,N_4470);
nor U5447 (N_5447,N_4889,N_4794);
nand U5448 (N_5448,N_4591,N_4467);
nand U5449 (N_5449,N_4592,N_4566);
and U5450 (N_5450,N_4789,N_4959);
or U5451 (N_5451,N_4697,N_4998);
nand U5452 (N_5452,N_4869,N_4782);
nand U5453 (N_5453,N_4969,N_4692);
xnor U5454 (N_5454,N_4905,N_4978);
nand U5455 (N_5455,N_4636,N_4733);
and U5456 (N_5456,N_4521,N_4741);
or U5457 (N_5457,N_4727,N_4597);
xnor U5458 (N_5458,N_4666,N_4902);
nor U5459 (N_5459,N_4787,N_4659);
xor U5460 (N_5460,N_4410,N_4637);
xor U5461 (N_5461,N_4687,N_4719);
nand U5462 (N_5462,N_4955,N_4563);
or U5463 (N_5463,N_4779,N_4474);
xnor U5464 (N_5464,N_4674,N_4409);
or U5465 (N_5465,N_4732,N_4983);
nand U5466 (N_5466,N_4784,N_4895);
xnor U5467 (N_5467,N_4949,N_4908);
nand U5468 (N_5468,N_4561,N_4689);
nor U5469 (N_5469,N_4983,N_4821);
and U5470 (N_5470,N_4608,N_4409);
nor U5471 (N_5471,N_4969,N_4451);
nand U5472 (N_5472,N_4794,N_4670);
xor U5473 (N_5473,N_4614,N_4484);
nor U5474 (N_5474,N_4467,N_4983);
and U5475 (N_5475,N_4699,N_4691);
nor U5476 (N_5476,N_4737,N_4816);
nand U5477 (N_5477,N_4679,N_4478);
and U5478 (N_5478,N_4936,N_4785);
and U5479 (N_5479,N_4973,N_4692);
and U5480 (N_5480,N_4644,N_4617);
nor U5481 (N_5481,N_4613,N_4912);
xnor U5482 (N_5482,N_4895,N_4405);
or U5483 (N_5483,N_4378,N_4988);
and U5484 (N_5484,N_4752,N_4601);
and U5485 (N_5485,N_4643,N_4388);
and U5486 (N_5486,N_4833,N_4605);
xor U5487 (N_5487,N_4880,N_4396);
nor U5488 (N_5488,N_4594,N_4533);
nor U5489 (N_5489,N_4390,N_4732);
nand U5490 (N_5490,N_4822,N_4923);
xor U5491 (N_5491,N_4566,N_4947);
and U5492 (N_5492,N_4416,N_4937);
xnor U5493 (N_5493,N_4636,N_4417);
xnor U5494 (N_5494,N_4792,N_4744);
nor U5495 (N_5495,N_4784,N_4674);
nand U5496 (N_5496,N_4830,N_4875);
nand U5497 (N_5497,N_4523,N_4961);
and U5498 (N_5498,N_4642,N_4479);
nor U5499 (N_5499,N_4650,N_4841);
nand U5500 (N_5500,N_4519,N_4693);
and U5501 (N_5501,N_4982,N_4551);
or U5502 (N_5502,N_4970,N_4822);
or U5503 (N_5503,N_4511,N_4874);
xnor U5504 (N_5504,N_4875,N_4894);
and U5505 (N_5505,N_4995,N_4696);
nor U5506 (N_5506,N_4653,N_4934);
and U5507 (N_5507,N_4739,N_4777);
or U5508 (N_5508,N_4727,N_4953);
or U5509 (N_5509,N_4420,N_4432);
and U5510 (N_5510,N_4474,N_4587);
nand U5511 (N_5511,N_4983,N_4404);
nand U5512 (N_5512,N_4697,N_4392);
or U5513 (N_5513,N_4735,N_4951);
nand U5514 (N_5514,N_4667,N_4906);
and U5515 (N_5515,N_4583,N_4988);
and U5516 (N_5516,N_4967,N_4541);
and U5517 (N_5517,N_4459,N_4994);
xnor U5518 (N_5518,N_4536,N_4614);
nand U5519 (N_5519,N_4886,N_4498);
nor U5520 (N_5520,N_4971,N_4822);
nor U5521 (N_5521,N_4456,N_4510);
or U5522 (N_5522,N_4649,N_4948);
nor U5523 (N_5523,N_4495,N_4396);
xor U5524 (N_5524,N_4479,N_4908);
and U5525 (N_5525,N_4651,N_4921);
or U5526 (N_5526,N_4559,N_4959);
and U5527 (N_5527,N_4846,N_4539);
and U5528 (N_5528,N_4390,N_4898);
or U5529 (N_5529,N_4776,N_4542);
and U5530 (N_5530,N_4639,N_4856);
nand U5531 (N_5531,N_4559,N_4836);
xnor U5532 (N_5532,N_4863,N_4906);
or U5533 (N_5533,N_4951,N_4937);
or U5534 (N_5534,N_4375,N_4638);
or U5535 (N_5535,N_4639,N_4813);
nor U5536 (N_5536,N_4525,N_4806);
nand U5537 (N_5537,N_4900,N_4773);
nor U5538 (N_5538,N_4604,N_4893);
or U5539 (N_5539,N_4492,N_4452);
nand U5540 (N_5540,N_4761,N_4998);
and U5541 (N_5541,N_4520,N_4441);
nand U5542 (N_5542,N_4671,N_4488);
or U5543 (N_5543,N_4436,N_4533);
nor U5544 (N_5544,N_4471,N_4595);
and U5545 (N_5545,N_4563,N_4473);
nand U5546 (N_5546,N_4464,N_4722);
xnor U5547 (N_5547,N_4845,N_4798);
and U5548 (N_5548,N_4606,N_4500);
nand U5549 (N_5549,N_4951,N_4985);
nor U5550 (N_5550,N_4777,N_4447);
nor U5551 (N_5551,N_4401,N_4790);
or U5552 (N_5552,N_4867,N_4686);
nor U5553 (N_5553,N_4545,N_4635);
xor U5554 (N_5554,N_4741,N_4558);
or U5555 (N_5555,N_4904,N_4434);
nand U5556 (N_5556,N_4588,N_4387);
or U5557 (N_5557,N_4567,N_4708);
xor U5558 (N_5558,N_4417,N_4747);
xnor U5559 (N_5559,N_4866,N_4439);
nor U5560 (N_5560,N_4618,N_4756);
nand U5561 (N_5561,N_4990,N_4641);
nand U5562 (N_5562,N_4895,N_4436);
xor U5563 (N_5563,N_4504,N_4833);
or U5564 (N_5564,N_4906,N_4703);
xnor U5565 (N_5565,N_4683,N_4597);
or U5566 (N_5566,N_4847,N_4609);
nor U5567 (N_5567,N_4389,N_4936);
and U5568 (N_5568,N_4614,N_4969);
or U5569 (N_5569,N_4529,N_4451);
nor U5570 (N_5570,N_4449,N_4475);
nand U5571 (N_5571,N_4514,N_4549);
and U5572 (N_5572,N_4490,N_4530);
nor U5573 (N_5573,N_4684,N_4764);
nand U5574 (N_5574,N_4830,N_4681);
nor U5575 (N_5575,N_4826,N_4659);
nor U5576 (N_5576,N_4717,N_4599);
nor U5577 (N_5577,N_4660,N_4648);
or U5578 (N_5578,N_4567,N_4691);
xor U5579 (N_5579,N_4908,N_4486);
or U5580 (N_5580,N_4581,N_4864);
nand U5581 (N_5581,N_4724,N_4929);
nand U5582 (N_5582,N_4531,N_4387);
nor U5583 (N_5583,N_4865,N_4426);
nand U5584 (N_5584,N_4931,N_4890);
xnor U5585 (N_5585,N_4960,N_4715);
nand U5586 (N_5586,N_4463,N_4612);
xor U5587 (N_5587,N_4518,N_4893);
or U5588 (N_5588,N_4456,N_4450);
nor U5589 (N_5589,N_4746,N_4682);
nor U5590 (N_5590,N_4927,N_4437);
nand U5591 (N_5591,N_4596,N_4765);
xnor U5592 (N_5592,N_4653,N_4454);
or U5593 (N_5593,N_4576,N_4604);
and U5594 (N_5594,N_4843,N_4551);
or U5595 (N_5595,N_4985,N_4892);
xnor U5596 (N_5596,N_4643,N_4919);
xor U5597 (N_5597,N_4463,N_4889);
xor U5598 (N_5598,N_4935,N_4525);
nor U5599 (N_5599,N_4645,N_4437);
or U5600 (N_5600,N_4383,N_4624);
nand U5601 (N_5601,N_4746,N_4799);
and U5602 (N_5602,N_4384,N_4687);
and U5603 (N_5603,N_4756,N_4686);
and U5604 (N_5604,N_4891,N_4534);
nand U5605 (N_5605,N_4680,N_4993);
or U5606 (N_5606,N_4696,N_4781);
and U5607 (N_5607,N_4749,N_4692);
xnor U5608 (N_5608,N_4385,N_4975);
xnor U5609 (N_5609,N_4889,N_4831);
nor U5610 (N_5610,N_4707,N_4485);
and U5611 (N_5611,N_4442,N_4896);
xor U5612 (N_5612,N_4477,N_4674);
nand U5613 (N_5613,N_4603,N_4573);
nor U5614 (N_5614,N_4868,N_4827);
or U5615 (N_5615,N_4930,N_4786);
and U5616 (N_5616,N_4820,N_4688);
nor U5617 (N_5617,N_4684,N_4993);
or U5618 (N_5618,N_4468,N_4966);
and U5619 (N_5619,N_4619,N_4956);
nand U5620 (N_5620,N_4637,N_4671);
xnor U5621 (N_5621,N_4880,N_4917);
nor U5622 (N_5622,N_4873,N_4539);
or U5623 (N_5623,N_4850,N_4610);
nand U5624 (N_5624,N_4729,N_4748);
nor U5625 (N_5625,N_5326,N_5470);
xnor U5626 (N_5626,N_5460,N_5510);
nor U5627 (N_5627,N_5304,N_5048);
nor U5628 (N_5628,N_5603,N_5187);
and U5629 (N_5629,N_5531,N_5329);
nand U5630 (N_5630,N_5581,N_5497);
xor U5631 (N_5631,N_5574,N_5298);
nand U5632 (N_5632,N_5611,N_5166);
or U5633 (N_5633,N_5554,N_5387);
or U5634 (N_5634,N_5135,N_5553);
and U5635 (N_5635,N_5025,N_5544);
nand U5636 (N_5636,N_5509,N_5494);
nand U5637 (N_5637,N_5065,N_5405);
xor U5638 (N_5638,N_5511,N_5588);
or U5639 (N_5639,N_5317,N_5277);
nor U5640 (N_5640,N_5348,N_5491);
nor U5641 (N_5641,N_5243,N_5161);
or U5642 (N_5642,N_5552,N_5534);
nand U5643 (N_5643,N_5120,N_5044);
or U5644 (N_5644,N_5462,N_5256);
nand U5645 (N_5645,N_5620,N_5394);
nand U5646 (N_5646,N_5075,N_5282);
nor U5647 (N_5647,N_5076,N_5582);
nor U5648 (N_5648,N_5035,N_5302);
nand U5649 (N_5649,N_5176,N_5296);
nand U5650 (N_5650,N_5252,N_5440);
and U5651 (N_5651,N_5518,N_5205);
nand U5652 (N_5652,N_5441,N_5308);
xor U5653 (N_5653,N_5098,N_5040);
or U5654 (N_5654,N_5358,N_5384);
nor U5655 (N_5655,N_5274,N_5433);
nand U5656 (N_5656,N_5332,N_5002);
xor U5657 (N_5657,N_5072,N_5013);
nand U5658 (N_5658,N_5220,N_5335);
nor U5659 (N_5659,N_5269,N_5170);
nor U5660 (N_5660,N_5221,N_5356);
nand U5661 (N_5661,N_5601,N_5112);
xor U5662 (N_5662,N_5505,N_5287);
and U5663 (N_5663,N_5105,N_5436);
and U5664 (N_5664,N_5539,N_5536);
xnor U5665 (N_5665,N_5041,N_5343);
and U5666 (N_5666,N_5472,N_5344);
nor U5667 (N_5667,N_5144,N_5503);
or U5668 (N_5668,N_5283,N_5226);
and U5669 (N_5669,N_5514,N_5237);
nor U5670 (N_5670,N_5430,N_5006);
and U5671 (N_5671,N_5489,N_5571);
and U5672 (N_5672,N_5416,N_5443);
or U5673 (N_5673,N_5610,N_5125);
and U5674 (N_5674,N_5190,N_5371);
and U5675 (N_5675,N_5078,N_5306);
and U5676 (N_5676,N_5540,N_5527);
nor U5677 (N_5677,N_5342,N_5026);
nor U5678 (N_5678,N_5107,N_5385);
nor U5679 (N_5679,N_5070,N_5369);
nand U5680 (N_5680,N_5357,N_5521);
or U5681 (N_5681,N_5268,N_5207);
xnor U5682 (N_5682,N_5160,N_5073);
nor U5683 (N_5683,N_5355,N_5362);
nor U5684 (N_5684,N_5379,N_5297);
xnor U5685 (N_5685,N_5364,N_5437);
and U5686 (N_5686,N_5255,N_5001);
or U5687 (N_5687,N_5007,N_5613);
or U5688 (N_5688,N_5047,N_5557);
xnor U5689 (N_5689,N_5471,N_5608);
nand U5690 (N_5690,N_5110,N_5151);
and U5691 (N_5691,N_5173,N_5483);
nand U5692 (N_5692,N_5109,N_5008);
xnor U5693 (N_5693,N_5270,N_5087);
nand U5694 (N_5694,N_5427,N_5417);
nor U5695 (N_5695,N_5147,N_5012);
and U5696 (N_5696,N_5447,N_5508);
and U5697 (N_5697,N_5215,N_5542);
or U5698 (N_5698,N_5003,N_5623);
or U5699 (N_5699,N_5402,N_5555);
and U5700 (N_5700,N_5301,N_5398);
nor U5701 (N_5701,N_5543,N_5590);
and U5702 (N_5702,N_5568,N_5476);
or U5703 (N_5703,N_5077,N_5278);
nor U5704 (N_5704,N_5396,N_5030);
nor U5705 (N_5705,N_5023,N_5501);
xor U5706 (N_5706,N_5341,N_5480);
nor U5707 (N_5707,N_5088,N_5114);
xnor U5708 (N_5708,N_5216,N_5324);
nand U5709 (N_5709,N_5349,N_5272);
nand U5710 (N_5710,N_5591,N_5352);
xnor U5711 (N_5711,N_5456,N_5119);
nand U5712 (N_5712,N_5366,N_5411);
nor U5713 (N_5713,N_5530,N_5225);
and U5714 (N_5714,N_5218,N_5285);
nand U5715 (N_5715,N_5127,N_5015);
or U5716 (N_5716,N_5260,N_5280);
xnor U5717 (N_5717,N_5235,N_5361);
and U5718 (N_5718,N_5528,N_5318);
nand U5719 (N_5719,N_5422,N_5165);
xor U5720 (N_5720,N_5336,N_5079);
and U5721 (N_5721,N_5570,N_5419);
nand U5722 (N_5722,N_5210,N_5597);
and U5723 (N_5723,N_5195,N_5082);
xnor U5724 (N_5724,N_5271,N_5551);
or U5725 (N_5725,N_5016,N_5463);
nor U5726 (N_5726,N_5180,N_5381);
nor U5727 (N_5727,N_5535,N_5525);
xor U5728 (N_5728,N_5621,N_5523);
nor U5729 (N_5729,N_5467,N_5484);
xor U5730 (N_5730,N_5259,N_5089);
xnor U5731 (N_5731,N_5322,N_5186);
and U5732 (N_5732,N_5141,N_5258);
and U5733 (N_5733,N_5395,N_5547);
and U5734 (N_5734,N_5262,N_5616);
nor U5735 (N_5735,N_5377,N_5245);
and U5736 (N_5736,N_5313,N_5010);
and U5737 (N_5737,N_5131,N_5512);
nand U5738 (N_5738,N_5101,N_5222);
nor U5739 (N_5739,N_5071,N_5241);
nor U5740 (N_5740,N_5049,N_5307);
nor U5741 (N_5741,N_5019,N_5290);
xnor U5742 (N_5742,N_5011,N_5199);
nand U5743 (N_5743,N_5202,N_5624);
and U5744 (N_5744,N_5042,N_5085);
and U5745 (N_5745,N_5375,N_5099);
xnor U5746 (N_5746,N_5248,N_5171);
nand U5747 (N_5747,N_5567,N_5622);
and U5748 (N_5748,N_5407,N_5168);
and U5749 (N_5749,N_5498,N_5090);
nand U5750 (N_5750,N_5583,N_5565);
xnor U5751 (N_5751,N_5064,N_5577);
nor U5752 (N_5752,N_5121,N_5572);
and U5753 (N_5753,N_5055,N_5486);
or U5754 (N_5754,N_5424,N_5293);
nand U5755 (N_5755,N_5589,N_5445);
nand U5756 (N_5756,N_5315,N_5517);
nor U5757 (N_5757,N_5281,N_5431);
nand U5758 (N_5758,N_5206,N_5247);
nand U5759 (N_5759,N_5400,N_5350);
nand U5760 (N_5760,N_5333,N_5057);
nand U5761 (N_5761,N_5029,N_5148);
or U5762 (N_5762,N_5466,N_5435);
nand U5763 (N_5763,N_5576,N_5236);
and U5764 (N_5764,N_5607,N_5178);
nand U5765 (N_5765,N_5397,N_5428);
and U5766 (N_5766,N_5383,N_5038);
xor U5767 (N_5767,N_5198,N_5478);
or U5768 (N_5768,N_5227,N_5106);
xor U5769 (N_5769,N_5123,N_5414);
and U5770 (N_5770,N_5338,N_5091);
nand U5771 (N_5771,N_5179,N_5558);
nand U5772 (N_5772,N_5132,N_5140);
or U5773 (N_5773,N_5124,N_5139);
nand U5774 (N_5774,N_5153,N_5056);
and U5775 (N_5775,N_5021,N_5291);
nand U5776 (N_5776,N_5507,N_5059);
nand U5777 (N_5777,N_5134,N_5500);
nor U5778 (N_5778,N_5410,N_5152);
nor U5779 (N_5779,N_5446,N_5081);
and U5780 (N_5780,N_5031,N_5244);
and U5781 (N_5781,N_5193,N_5217);
xnor U5782 (N_5782,N_5309,N_5230);
nor U5783 (N_5783,N_5201,N_5284);
nor U5784 (N_5784,N_5191,N_5005);
nor U5785 (N_5785,N_5239,N_5150);
or U5786 (N_5786,N_5550,N_5420);
xnor U5787 (N_5787,N_5212,N_5519);
nor U5788 (N_5788,N_5374,N_5325);
nor U5789 (N_5789,N_5457,N_5122);
nor U5790 (N_5790,N_5063,N_5563);
or U5791 (N_5791,N_5382,N_5323);
nand U5792 (N_5792,N_5182,N_5156);
nand U5793 (N_5793,N_5312,N_5067);
xor U5794 (N_5794,N_5213,N_5051);
nor U5795 (N_5795,N_5251,N_5328);
or U5796 (N_5796,N_5368,N_5022);
and U5797 (N_5797,N_5254,N_5017);
or U5798 (N_5798,N_5200,N_5275);
xnor U5799 (N_5799,N_5592,N_5181);
or U5800 (N_5800,N_5286,N_5545);
xor U5801 (N_5801,N_5203,N_5584);
and U5802 (N_5802,N_5533,N_5189);
and U5803 (N_5803,N_5432,N_5231);
and U5804 (N_5804,N_5609,N_5619);
nand U5805 (N_5805,N_5249,N_5188);
and U5806 (N_5806,N_5115,N_5177);
nand U5807 (N_5807,N_5175,N_5103);
xor U5808 (N_5808,N_5403,N_5050);
nand U5809 (N_5809,N_5204,N_5224);
and U5810 (N_5810,N_5459,N_5000);
nand U5811 (N_5811,N_5464,N_5184);
nor U5812 (N_5812,N_5606,N_5526);
or U5813 (N_5813,N_5311,N_5365);
nand U5814 (N_5814,N_5455,N_5367);
and U5815 (N_5815,N_5288,N_5549);
xor U5816 (N_5816,N_5043,N_5209);
xnor U5817 (N_5817,N_5569,N_5066);
and U5818 (N_5818,N_5585,N_5492);
xor U5819 (N_5819,N_5600,N_5265);
xor U5820 (N_5820,N_5575,N_5439);
or U5821 (N_5821,N_5094,N_5593);
or U5822 (N_5822,N_5453,N_5093);
xnor U5823 (N_5823,N_5538,N_5363);
and U5824 (N_5824,N_5174,N_5353);
and U5825 (N_5825,N_5034,N_5359);
and U5826 (N_5826,N_5253,N_5334);
and U5827 (N_5827,N_5228,N_5421);
nand U5828 (N_5828,N_5018,N_5409);
xnor U5829 (N_5829,N_5149,N_5305);
nand U5830 (N_5830,N_5164,N_5194);
nor U5831 (N_5831,N_5319,N_5442);
nor U5832 (N_5832,N_5111,N_5426);
xor U5833 (N_5833,N_5234,N_5586);
and U5834 (N_5834,N_5157,N_5504);
nor U5835 (N_5835,N_5027,N_5303);
nand U5836 (N_5836,N_5145,N_5337);
and U5837 (N_5837,N_5321,N_5423);
nand U5838 (N_5838,N_5473,N_5246);
and U5839 (N_5839,N_5448,N_5595);
nor U5840 (N_5840,N_5104,N_5133);
nand U5841 (N_5841,N_5391,N_5300);
xnor U5842 (N_5842,N_5159,N_5295);
xor U5843 (N_5843,N_5564,N_5580);
nor U5844 (N_5844,N_5273,N_5605);
or U5845 (N_5845,N_5039,N_5331);
xnor U5846 (N_5846,N_5211,N_5418);
or U5847 (N_5847,N_5354,N_5380);
nor U5848 (N_5848,N_5158,N_5434);
and U5849 (N_5849,N_5292,N_5232);
nor U5850 (N_5850,N_5294,N_5024);
and U5851 (N_5851,N_5095,N_5172);
nor U5852 (N_5852,N_5559,N_5392);
and U5853 (N_5853,N_5192,N_5429);
nor U5854 (N_5854,N_5233,N_5425);
nand U5855 (N_5855,N_5458,N_5412);
nor U5856 (N_5856,N_5345,N_5046);
and U5857 (N_5857,N_5495,N_5546);
nor U5858 (N_5858,N_5155,N_5515);
and U5859 (N_5859,N_5481,N_5136);
nand U5860 (N_5860,N_5548,N_5068);
nand U5861 (N_5861,N_5524,N_5080);
and U5862 (N_5862,N_5346,N_5477);
or U5863 (N_5863,N_5163,N_5537);
nor U5864 (N_5864,N_5242,N_5566);
nand U5865 (N_5865,N_5360,N_5037);
xor U5866 (N_5866,N_5154,N_5485);
nand U5867 (N_5867,N_5378,N_5062);
nor U5868 (N_5868,N_5386,N_5413);
xnor U5869 (N_5869,N_5061,N_5113);
nand U5870 (N_5870,N_5074,N_5320);
or U5871 (N_5871,N_5452,N_5474);
nor U5872 (N_5872,N_5351,N_5108);
or U5873 (N_5873,N_5408,N_5240);
xnor U5874 (N_5874,N_5506,N_5614);
nor U5875 (N_5875,N_5069,N_5579);
nand U5876 (N_5876,N_5594,N_5615);
and U5877 (N_5877,N_5482,N_5496);
or U5878 (N_5878,N_5314,N_5562);
or U5879 (N_5879,N_5347,N_5261);
xor U5880 (N_5880,N_5465,N_5117);
or U5881 (N_5881,N_5529,N_5185);
xor U5882 (N_5882,N_5014,N_5196);
and U5883 (N_5883,N_5561,N_5223);
or U5884 (N_5884,N_5266,N_5138);
and U5885 (N_5885,N_5146,N_5004);
nand U5886 (N_5886,N_5461,N_5310);
nand U5887 (N_5887,N_5479,N_5263);
nand U5888 (N_5888,N_5143,N_5167);
xnor U5889 (N_5889,N_5052,N_5129);
xor U5890 (N_5890,N_5475,N_5388);
or U5891 (N_5891,N_5116,N_5370);
xor U5892 (N_5892,N_5264,N_5401);
and U5893 (N_5893,N_5451,N_5490);
nand U5894 (N_5894,N_5276,N_5267);
nor U5895 (N_5895,N_5084,N_5086);
and U5896 (N_5896,N_5522,N_5100);
or U5897 (N_5897,N_5541,N_5045);
xor U5898 (N_5898,N_5208,N_5009);
or U5899 (N_5899,N_5599,N_5340);
xnor U5900 (N_5900,N_5053,N_5036);
nand U5901 (N_5901,N_5032,N_5330);
nor U5902 (N_5902,N_5556,N_5617);
or U5903 (N_5903,N_5299,N_5372);
nand U5904 (N_5904,N_5137,N_5142);
nor U5905 (N_5905,N_5560,N_5169);
nand U5906 (N_5906,N_5454,N_5126);
nand U5907 (N_5907,N_5183,N_5596);
xor U5908 (N_5908,N_5573,N_5118);
nand U5909 (N_5909,N_5092,N_5612);
or U5910 (N_5910,N_5487,N_5130);
nand U5911 (N_5911,N_5097,N_5469);
or U5912 (N_5912,N_5393,N_5618);
nand U5913 (N_5913,N_5229,N_5602);
nand U5914 (N_5914,N_5096,N_5083);
nor U5915 (N_5915,N_5028,N_5578);
nor U5916 (N_5916,N_5493,N_5058);
xor U5917 (N_5917,N_5102,N_5238);
and U5918 (N_5918,N_5339,N_5449);
or U5919 (N_5919,N_5390,N_5373);
nand U5920 (N_5920,N_5404,N_5250);
xnor U5921 (N_5921,N_5499,N_5327);
and U5922 (N_5922,N_5438,N_5316);
xnor U5923 (N_5923,N_5197,N_5598);
and U5924 (N_5924,N_5468,N_5279);
or U5925 (N_5925,N_5502,N_5532);
nand U5926 (N_5926,N_5060,N_5162);
xnor U5927 (N_5927,N_5033,N_5399);
and U5928 (N_5928,N_5020,N_5128);
nand U5929 (N_5929,N_5376,N_5289);
nor U5930 (N_5930,N_5219,N_5406);
or U5931 (N_5931,N_5587,N_5450);
nor U5932 (N_5932,N_5415,N_5257);
nor U5933 (N_5933,N_5516,N_5389);
nand U5934 (N_5934,N_5444,N_5054);
nand U5935 (N_5935,N_5520,N_5488);
or U5936 (N_5936,N_5214,N_5513);
nand U5937 (N_5937,N_5604,N_5485);
or U5938 (N_5938,N_5117,N_5134);
or U5939 (N_5939,N_5014,N_5001);
xnor U5940 (N_5940,N_5579,N_5472);
nand U5941 (N_5941,N_5360,N_5116);
nor U5942 (N_5942,N_5156,N_5266);
xor U5943 (N_5943,N_5174,N_5308);
or U5944 (N_5944,N_5577,N_5523);
nor U5945 (N_5945,N_5574,N_5078);
or U5946 (N_5946,N_5068,N_5410);
and U5947 (N_5947,N_5366,N_5478);
or U5948 (N_5948,N_5158,N_5121);
or U5949 (N_5949,N_5537,N_5043);
and U5950 (N_5950,N_5504,N_5618);
xnor U5951 (N_5951,N_5034,N_5154);
and U5952 (N_5952,N_5353,N_5618);
and U5953 (N_5953,N_5229,N_5086);
nand U5954 (N_5954,N_5544,N_5170);
nand U5955 (N_5955,N_5286,N_5293);
nor U5956 (N_5956,N_5095,N_5177);
xor U5957 (N_5957,N_5213,N_5463);
nand U5958 (N_5958,N_5192,N_5579);
or U5959 (N_5959,N_5287,N_5610);
and U5960 (N_5960,N_5187,N_5117);
nand U5961 (N_5961,N_5322,N_5107);
nand U5962 (N_5962,N_5490,N_5138);
nor U5963 (N_5963,N_5018,N_5170);
nor U5964 (N_5964,N_5018,N_5175);
or U5965 (N_5965,N_5431,N_5591);
xor U5966 (N_5966,N_5286,N_5225);
and U5967 (N_5967,N_5616,N_5003);
xor U5968 (N_5968,N_5106,N_5182);
xor U5969 (N_5969,N_5243,N_5262);
nand U5970 (N_5970,N_5042,N_5264);
nor U5971 (N_5971,N_5443,N_5004);
nor U5972 (N_5972,N_5032,N_5423);
xnor U5973 (N_5973,N_5603,N_5216);
and U5974 (N_5974,N_5380,N_5321);
xor U5975 (N_5975,N_5364,N_5018);
nand U5976 (N_5976,N_5296,N_5232);
xnor U5977 (N_5977,N_5116,N_5035);
and U5978 (N_5978,N_5305,N_5402);
nand U5979 (N_5979,N_5445,N_5070);
and U5980 (N_5980,N_5523,N_5210);
xnor U5981 (N_5981,N_5461,N_5297);
nand U5982 (N_5982,N_5023,N_5514);
nor U5983 (N_5983,N_5039,N_5485);
nor U5984 (N_5984,N_5059,N_5170);
nor U5985 (N_5985,N_5594,N_5493);
nor U5986 (N_5986,N_5423,N_5570);
and U5987 (N_5987,N_5350,N_5100);
and U5988 (N_5988,N_5215,N_5079);
nand U5989 (N_5989,N_5258,N_5106);
or U5990 (N_5990,N_5478,N_5341);
xnor U5991 (N_5991,N_5507,N_5266);
or U5992 (N_5992,N_5393,N_5372);
nor U5993 (N_5993,N_5505,N_5121);
and U5994 (N_5994,N_5388,N_5158);
or U5995 (N_5995,N_5031,N_5618);
nor U5996 (N_5996,N_5600,N_5575);
and U5997 (N_5997,N_5400,N_5320);
nand U5998 (N_5998,N_5293,N_5053);
or U5999 (N_5999,N_5148,N_5547);
xor U6000 (N_6000,N_5514,N_5500);
and U6001 (N_6001,N_5047,N_5599);
xor U6002 (N_6002,N_5176,N_5318);
or U6003 (N_6003,N_5513,N_5088);
or U6004 (N_6004,N_5049,N_5570);
or U6005 (N_6005,N_5552,N_5344);
nor U6006 (N_6006,N_5604,N_5020);
xnor U6007 (N_6007,N_5153,N_5448);
nor U6008 (N_6008,N_5474,N_5224);
nand U6009 (N_6009,N_5586,N_5228);
and U6010 (N_6010,N_5045,N_5568);
nor U6011 (N_6011,N_5372,N_5545);
nand U6012 (N_6012,N_5373,N_5472);
nand U6013 (N_6013,N_5181,N_5506);
and U6014 (N_6014,N_5470,N_5457);
nor U6015 (N_6015,N_5413,N_5016);
nand U6016 (N_6016,N_5421,N_5386);
nor U6017 (N_6017,N_5159,N_5031);
nor U6018 (N_6018,N_5587,N_5463);
xor U6019 (N_6019,N_5142,N_5219);
and U6020 (N_6020,N_5472,N_5228);
xnor U6021 (N_6021,N_5498,N_5308);
or U6022 (N_6022,N_5039,N_5352);
xor U6023 (N_6023,N_5222,N_5171);
nand U6024 (N_6024,N_5525,N_5434);
or U6025 (N_6025,N_5080,N_5114);
xor U6026 (N_6026,N_5583,N_5060);
nand U6027 (N_6027,N_5495,N_5108);
xnor U6028 (N_6028,N_5348,N_5221);
nand U6029 (N_6029,N_5388,N_5319);
nand U6030 (N_6030,N_5379,N_5385);
nand U6031 (N_6031,N_5103,N_5213);
and U6032 (N_6032,N_5277,N_5342);
and U6033 (N_6033,N_5061,N_5489);
or U6034 (N_6034,N_5571,N_5414);
or U6035 (N_6035,N_5365,N_5510);
and U6036 (N_6036,N_5579,N_5412);
xor U6037 (N_6037,N_5149,N_5518);
and U6038 (N_6038,N_5352,N_5205);
and U6039 (N_6039,N_5427,N_5246);
nand U6040 (N_6040,N_5029,N_5425);
or U6041 (N_6041,N_5502,N_5422);
and U6042 (N_6042,N_5087,N_5546);
nand U6043 (N_6043,N_5566,N_5082);
xor U6044 (N_6044,N_5578,N_5060);
and U6045 (N_6045,N_5322,N_5004);
or U6046 (N_6046,N_5333,N_5603);
or U6047 (N_6047,N_5413,N_5222);
xor U6048 (N_6048,N_5314,N_5307);
and U6049 (N_6049,N_5550,N_5597);
nor U6050 (N_6050,N_5610,N_5187);
nor U6051 (N_6051,N_5290,N_5413);
nor U6052 (N_6052,N_5287,N_5310);
xnor U6053 (N_6053,N_5310,N_5368);
xnor U6054 (N_6054,N_5411,N_5432);
and U6055 (N_6055,N_5428,N_5454);
or U6056 (N_6056,N_5512,N_5132);
nand U6057 (N_6057,N_5439,N_5535);
nand U6058 (N_6058,N_5382,N_5227);
and U6059 (N_6059,N_5560,N_5544);
nand U6060 (N_6060,N_5577,N_5067);
xor U6061 (N_6061,N_5588,N_5358);
nor U6062 (N_6062,N_5516,N_5029);
or U6063 (N_6063,N_5394,N_5281);
and U6064 (N_6064,N_5140,N_5287);
xnor U6065 (N_6065,N_5266,N_5002);
nand U6066 (N_6066,N_5611,N_5030);
and U6067 (N_6067,N_5153,N_5172);
nor U6068 (N_6068,N_5076,N_5574);
nand U6069 (N_6069,N_5045,N_5184);
nor U6070 (N_6070,N_5373,N_5226);
xnor U6071 (N_6071,N_5298,N_5337);
nand U6072 (N_6072,N_5435,N_5600);
and U6073 (N_6073,N_5207,N_5116);
and U6074 (N_6074,N_5140,N_5602);
xnor U6075 (N_6075,N_5488,N_5003);
nand U6076 (N_6076,N_5434,N_5261);
and U6077 (N_6077,N_5035,N_5325);
nor U6078 (N_6078,N_5321,N_5127);
and U6079 (N_6079,N_5130,N_5420);
nor U6080 (N_6080,N_5578,N_5285);
nand U6081 (N_6081,N_5622,N_5021);
nand U6082 (N_6082,N_5402,N_5128);
nand U6083 (N_6083,N_5197,N_5300);
nand U6084 (N_6084,N_5614,N_5598);
nor U6085 (N_6085,N_5247,N_5053);
nor U6086 (N_6086,N_5619,N_5512);
and U6087 (N_6087,N_5520,N_5382);
xnor U6088 (N_6088,N_5362,N_5108);
xor U6089 (N_6089,N_5069,N_5239);
nand U6090 (N_6090,N_5196,N_5114);
xnor U6091 (N_6091,N_5133,N_5362);
nor U6092 (N_6092,N_5111,N_5406);
nor U6093 (N_6093,N_5556,N_5229);
xnor U6094 (N_6094,N_5175,N_5128);
and U6095 (N_6095,N_5403,N_5324);
or U6096 (N_6096,N_5161,N_5142);
nor U6097 (N_6097,N_5152,N_5168);
xnor U6098 (N_6098,N_5439,N_5240);
or U6099 (N_6099,N_5239,N_5548);
nor U6100 (N_6100,N_5553,N_5184);
nor U6101 (N_6101,N_5154,N_5542);
or U6102 (N_6102,N_5301,N_5028);
nor U6103 (N_6103,N_5275,N_5589);
nand U6104 (N_6104,N_5560,N_5475);
and U6105 (N_6105,N_5451,N_5240);
or U6106 (N_6106,N_5613,N_5122);
nand U6107 (N_6107,N_5125,N_5349);
nor U6108 (N_6108,N_5484,N_5593);
nand U6109 (N_6109,N_5374,N_5256);
nor U6110 (N_6110,N_5154,N_5168);
and U6111 (N_6111,N_5561,N_5447);
nand U6112 (N_6112,N_5331,N_5091);
nor U6113 (N_6113,N_5594,N_5312);
nand U6114 (N_6114,N_5153,N_5014);
and U6115 (N_6115,N_5367,N_5257);
nand U6116 (N_6116,N_5223,N_5484);
nand U6117 (N_6117,N_5104,N_5538);
nor U6118 (N_6118,N_5454,N_5579);
and U6119 (N_6119,N_5527,N_5090);
nor U6120 (N_6120,N_5478,N_5559);
and U6121 (N_6121,N_5469,N_5031);
nand U6122 (N_6122,N_5349,N_5574);
xnor U6123 (N_6123,N_5341,N_5531);
and U6124 (N_6124,N_5314,N_5421);
nor U6125 (N_6125,N_5216,N_5597);
xnor U6126 (N_6126,N_5186,N_5528);
nor U6127 (N_6127,N_5327,N_5421);
nor U6128 (N_6128,N_5423,N_5075);
and U6129 (N_6129,N_5610,N_5431);
nor U6130 (N_6130,N_5195,N_5207);
or U6131 (N_6131,N_5079,N_5177);
xor U6132 (N_6132,N_5557,N_5497);
nor U6133 (N_6133,N_5603,N_5191);
or U6134 (N_6134,N_5015,N_5357);
nand U6135 (N_6135,N_5161,N_5269);
xnor U6136 (N_6136,N_5535,N_5577);
nand U6137 (N_6137,N_5212,N_5339);
xnor U6138 (N_6138,N_5194,N_5336);
xor U6139 (N_6139,N_5505,N_5066);
xnor U6140 (N_6140,N_5309,N_5368);
nand U6141 (N_6141,N_5032,N_5193);
nand U6142 (N_6142,N_5575,N_5373);
xor U6143 (N_6143,N_5221,N_5193);
nor U6144 (N_6144,N_5300,N_5348);
and U6145 (N_6145,N_5548,N_5533);
nand U6146 (N_6146,N_5283,N_5372);
nor U6147 (N_6147,N_5360,N_5427);
xnor U6148 (N_6148,N_5281,N_5102);
xnor U6149 (N_6149,N_5125,N_5209);
nand U6150 (N_6150,N_5420,N_5326);
or U6151 (N_6151,N_5607,N_5319);
nor U6152 (N_6152,N_5412,N_5047);
nand U6153 (N_6153,N_5610,N_5302);
and U6154 (N_6154,N_5583,N_5192);
and U6155 (N_6155,N_5538,N_5124);
nor U6156 (N_6156,N_5212,N_5124);
nor U6157 (N_6157,N_5114,N_5382);
nand U6158 (N_6158,N_5152,N_5187);
or U6159 (N_6159,N_5364,N_5405);
nand U6160 (N_6160,N_5526,N_5608);
and U6161 (N_6161,N_5508,N_5130);
nand U6162 (N_6162,N_5018,N_5546);
nand U6163 (N_6163,N_5375,N_5400);
nor U6164 (N_6164,N_5179,N_5473);
xnor U6165 (N_6165,N_5539,N_5439);
or U6166 (N_6166,N_5270,N_5617);
nor U6167 (N_6167,N_5392,N_5428);
and U6168 (N_6168,N_5492,N_5353);
and U6169 (N_6169,N_5173,N_5472);
and U6170 (N_6170,N_5498,N_5343);
xor U6171 (N_6171,N_5308,N_5145);
nor U6172 (N_6172,N_5161,N_5412);
nor U6173 (N_6173,N_5105,N_5569);
xor U6174 (N_6174,N_5620,N_5354);
xnor U6175 (N_6175,N_5218,N_5319);
nand U6176 (N_6176,N_5380,N_5386);
and U6177 (N_6177,N_5060,N_5561);
nor U6178 (N_6178,N_5216,N_5551);
nand U6179 (N_6179,N_5188,N_5245);
and U6180 (N_6180,N_5405,N_5439);
nand U6181 (N_6181,N_5066,N_5116);
or U6182 (N_6182,N_5449,N_5518);
or U6183 (N_6183,N_5460,N_5155);
xnor U6184 (N_6184,N_5263,N_5378);
nor U6185 (N_6185,N_5281,N_5335);
xor U6186 (N_6186,N_5544,N_5279);
nor U6187 (N_6187,N_5554,N_5364);
nor U6188 (N_6188,N_5035,N_5042);
nand U6189 (N_6189,N_5613,N_5034);
and U6190 (N_6190,N_5566,N_5382);
or U6191 (N_6191,N_5531,N_5391);
nand U6192 (N_6192,N_5306,N_5265);
nand U6193 (N_6193,N_5148,N_5185);
or U6194 (N_6194,N_5040,N_5400);
nor U6195 (N_6195,N_5494,N_5053);
nor U6196 (N_6196,N_5075,N_5582);
nand U6197 (N_6197,N_5493,N_5575);
xor U6198 (N_6198,N_5537,N_5563);
nor U6199 (N_6199,N_5385,N_5436);
xor U6200 (N_6200,N_5536,N_5004);
nor U6201 (N_6201,N_5246,N_5265);
nor U6202 (N_6202,N_5168,N_5198);
nor U6203 (N_6203,N_5552,N_5073);
nor U6204 (N_6204,N_5288,N_5026);
nand U6205 (N_6205,N_5209,N_5247);
nand U6206 (N_6206,N_5373,N_5604);
nand U6207 (N_6207,N_5570,N_5244);
or U6208 (N_6208,N_5177,N_5431);
nor U6209 (N_6209,N_5040,N_5269);
or U6210 (N_6210,N_5214,N_5518);
nand U6211 (N_6211,N_5365,N_5554);
nor U6212 (N_6212,N_5385,N_5123);
or U6213 (N_6213,N_5579,N_5148);
xor U6214 (N_6214,N_5291,N_5484);
xnor U6215 (N_6215,N_5600,N_5492);
xnor U6216 (N_6216,N_5215,N_5337);
xnor U6217 (N_6217,N_5595,N_5161);
xor U6218 (N_6218,N_5066,N_5606);
or U6219 (N_6219,N_5324,N_5221);
nand U6220 (N_6220,N_5155,N_5000);
xnor U6221 (N_6221,N_5116,N_5589);
nor U6222 (N_6222,N_5605,N_5560);
nand U6223 (N_6223,N_5585,N_5229);
or U6224 (N_6224,N_5201,N_5447);
and U6225 (N_6225,N_5381,N_5408);
xnor U6226 (N_6226,N_5500,N_5198);
nand U6227 (N_6227,N_5457,N_5336);
nor U6228 (N_6228,N_5270,N_5414);
nand U6229 (N_6229,N_5192,N_5116);
or U6230 (N_6230,N_5020,N_5041);
nor U6231 (N_6231,N_5409,N_5275);
nor U6232 (N_6232,N_5174,N_5453);
and U6233 (N_6233,N_5442,N_5510);
xor U6234 (N_6234,N_5202,N_5173);
nor U6235 (N_6235,N_5142,N_5251);
or U6236 (N_6236,N_5213,N_5202);
and U6237 (N_6237,N_5392,N_5188);
nor U6238 (N_6238,N_5597,N_5040);
xnor U6239 (N_6239,N_5443,N_5403);
nand U6240 (N_6240,N_5368,N_5294);
nor U6241 (N_6241,N_5443,N_5110);
or U6242 (N_6242,N_5124,N_5342);
nand U6243 (N_6243,N_5570,N_5556);
and U6244 (N_6244,N_5614,N_5318);
or U6245 (N_6245,N_5243,N_5139);
or U6246 (N_6246,N_5023,N_5065);
or U6247 (N_6247,N_5339,N_5086);
nand U6248 (N_6248,N_5326,N_5409);
or U6249 (N_6249,N_5411,N_5038);
and U6250 (N_6250,N_6073,N_5780);
nand U6251 (N_6251,N_6067,N_5712);
or U6252 (N_6252,N_6207,N_5814);
and U6253 (N_6253,N_5739,N_5965);
xor U6254 (N_6254,N_5848,N_5974);
xor U6255 (N_6255,N_6171,N_6153);
nor U6256 (N_6256,N_5864,N_5805);
xor U6257 (N_6257,N_6064,N_5783);
xnor U6258 (N_6258,N_5660,N_6039);
xnor U6259 (N_6259,N_6142,N_5710);
xor U6260 (N_6260,N_5694,N_5999);
or U6261 (N_6261,N_6045,N_5868);
xnor U6262 (N_6262,N_5996,N_5829);
xnor U6263 (N_6263,N_5917,N_6175);
or U6264 (N_6264,N_6030,N_5765);
or U6265 (N_6265,N_5909,N_5919);
xnor U6266 (N_6266,N_5859,N_5920);
nor U6267 (N_6267,N_5964,N_6110);
nor U6268 (N_6268,N_5994,N_5857);
or U6269 (N_6269,N_6076,N_5702);
nor U6270 (N_6270,N_6140,N_5792);
xnor U6271 (N_6271,N_5926,N_6230);
xnor U6272 (N_6272,N_5952,N_5757);
nand U6273 (N_6273,N_5652,N_5899);
xnor U6274 (N_6274,N_5930,N_5880);
nand U6275 (N_6275,N_6037,N_6132);
xnor U6276 (N_6276,N_5759,N_6246);
and U6277 (N_6277,N_5627,N_6018);
nand U6278 (N_6278,N_5657,N_6227);
nand U6279 (N_6279,N_5643,N_6221);
nand U6280 (N_6280,N_6034,N_5878);
and U6281 (N_6281,N_5680,N_6103);
nand U6282 (N_6282,N_6029,N_5916);
xor U6283 (N_6283,N_6178,N_6081);
and U6284 (N_6284,N_5847,N_5774);
xnor U6285 (N_6285,N_6150,N_5750);
nand U6286 (N_6286,N_6233,N_5747);
or U6287 (N_6287,N_5762,N_6088);
xnor U6288 (N_6288,N_5677,N_6024);
xnor U6289 (N_6289,N_5670,N_6104);
and U6290 (N_6290,N_6111,N_5778);
xor U6291 (N_6291,N_6137,N_6136);
and U6292 (N_6292,N_6209,N_5998);
and U6293 (N_6293,N_5675,N_5978);
or U6294 (N_6294,N_5701,N_6231);
nand U6295 (N_6295,N_5914,N_6046);
nand U6296 (N_6296,N_6077,N_6145);
and U6297 (N_6297,N_5696,N_6109);
nor U6298 (N_6298,N_6214,N_6082);
nor U6299 (N_6299,N_6011,N_6022);
and U6300 (N_6300,N_5826,N_6149);
and U6301 (N_6301,N_6044,N_6107);
xor U6302 (N_6302,N_5938,N_5997);
xor U6303 (N_6303,N_5649,N_6168);
xor U6304 (N_6304,N_5953,N_5713);
xnor U6305 (N_6305,N_5790,N_5659);
nand U6306 (N_6306,N_6213,N_6200);
nand U6307 (N_6307,N_5863,N_5960);
and U6308 (N_6308,N_6133,N_6186);
nand U6309 (N_6309,N_5800,N_5718);
and U6310 (N_6310,N_6249,N_5844);
nor U6311 (N_6311,N_5889,N_5976);
xor U6312 (N_6312,N_5937,N_5959);
and U6313 (N_6313,N_5834,N_5954);
or U6314 (N_6314,N_5895,N_5648);
or U6315 (N_6315,N_6206,N_5798);
nor U6316 (N_6316,N_6123,N_6162);
xor U6317 (N_6317,N_6156,N_6098);
xnor U6318 (N_6318,N_5647,N_5898);
and U6319 (N_6319,N_5927,N_5979);
nor U6320 (N_6320,N_6157,N_6166);
nand U6321 (N_6321,N_6247,N_5951);
and U6322 (N_6322,N_6095,N_5716);
nand U6323 (N_6323,N_6129,N_6054);
xor U6324 (N_6324,N_5676,N_5804);
xor U6325 (N_6325,N_6210,N_5632);
nand U6326 (N_6326,N_6012,N_5946);
nor U6327 (N_6327,N_5856,N_5745);
nor U6328 (N_6328,N_5654,N_6138);
or U6329 (N_6329,N_6079,N_6074);
and U6330 (N_6330,N_6196,N_6031);
xor U6331 (N_6331,N_6224,N_5653);
nor U6332 (N_6332,N_6236,N_6078);
or U6333 (N_6333,N_5687,N_6190);
or U6334 (N_6334,N_5874,N_5813);
nand U6335 (N_6335,N_6248,N_6052);
or U6336 (N_6336,N_5714,N_5931);
nor U6337 (N_6337,N_5781,N_5948);
xor U6338 (N_6338,N_5634,N_6155);
and U6339 (N_6339,N_5865,N_5761);
nand U6340 (N_6340,N_5981,N_5907);
and U6341 (N_6341,N_5892,N_5725);
and U6342 (N_6342,N_5934,N_5752);
xnor U6343 (N_6343,N_6219,N_5727);
nor U6344 (N_6344,N_6223,N_5855);
xnor U6345 (N_6345,N_6014,N_5949);
or U6346 (N_6346,N_5830,N_5630);
nand U6347 (N_6347,N_5886,N_5968);
and U6348 (N_6348,N_6043,N_5756);
and U6349 (N_6349,N_6013,N_5722);
nor U6350 (N_6350,N_6183,N_5656);
and U6351 (N_6351,N_6173,N_5950);
and U6352 (N_6352,N_6065,N_5900);
or U6353 (N_6353,N_6106,N_5625);
and U6354 (N_6354,N_6160,N_6120);
and U6355 (N_6355,N_5728,N_5658);
xnor U6356 (N_6356,N_5875,N_5985);
nor U6357 (N_6357,N_6174,N_6069);
nor U6358 (N_6358,N_5983,N_6100);
or U6359 (N_6359,N_5955,N_5901);
nor U6360 (N_6360,N_5906,N_5709);
nor U6361 (N_6361,N_6005,N_5651);
xnor U6362 (N_6362,N_6072,N_6003);
xor U6363 (N_6363,N_5662,N_5945);
and U6364 (N_6364,N_6068,N_5911);
or U6365 (N_6365,N_5681,N_6188);
xnor U6366 (N_6366,N_5980,N_5973);
xnor U6367 (N_6367,N_5704,N_5815);
and U6368 (N_6368,N_5683,N_5736);
xnor U6369 (N_6369,N_5962,N_5991);
and U6370 (N_6370,N_5754,N_5650);
or U6371 (N_6371,N_5833,N_5876);
nor U6372 (N_6372,N_6225,N_6125);
nor U6373 (N_6373,N_6047,N_5822);
xor U6374 (N_6374,N_5904,N_5843);
nand U6375 (N_6375,N_5738,N_6164);
or U6376 (N_6376,N_5885,N_6117);
xor U6377 (N_6377,N_5860,N_6180);
xnor U6378 (N_6378,N_5646,N_6205);
nor U6379 (N_6379,N_5672,N_6194);
or U6380 (N_6380,N_6135,N_5633);
or U6381 (N_6381,N_5720,N_5923);
xor U6382 (N_6382,N_5846,N_6185);
xor U6383 (N_6383,N_6114,N_5665);
nand U6384 (N_6384,N_5990,N_6017);
nand U6385 (N_6385,N_5912,N_6193);
or U6386 (N_6386,N_5777,N_5724);
xor U6387 (N_6387,N_5785,N_6050);
nand U6388 (N_6388,N_6038,N_5812);
or U6389 (N_6389,N_5682,N_5684);
nor U6390 (N_6390,N_6102,N_6176);
xor U6391 (N_6391,N_5883,N_5820);
and U6392 (N_6392,N_5775,N_5816);
nand U6393 (N_6393,N_5825,N_6062);
nand U6394 (N_6394,N_5989,N_6116);
nor U6395 (N_6395,N_5845,N_6232);
xor U6396 (N_6396,N_6222,N_6001);
and U6397 (N_6397,N_5849,N_6070);
nand U6398 (N_6398,N_6056,N_6090);
and U6399 (N_6399,N_5769,N_6241);
nor U6400 (N_6400,N_5903,N_6147);
nand U6401 (N_6401,N_5733,N_6226);
or U6402 (N_6402,N_6179,N_5636);
nor U6403 (N_6403,N_6189,N_5799);
xor U6404 (N_6404,N_5743,N_5664);
and U6405 (N_6405,N_5944,N_5741);
and U6406 (N_6406,N_5828,N_6032);
and U6407 (N_6407,N_6139,N_5890);
nand U6408 (N_6408,N_5933,N_5854);
or U6409 (N_6409,N_6218,N_5891);
nand U6410 (N_6410,N_5742,N_6115);
and U6411 (N_6411,N_6096,N_6009);
nor U6412 (N_6412,N_5821,N_5674);
or U6413 (N_6413,N_5786,N_6025);
nand U6414 (N_6414,N_6151,N_5689);
nand U6415 (N_6415,N_5666,N_6208);
and U6416 (N_6416,N_5852,N_5668);
xor U6417 (N_6417,N_5987,N_6126);
nor U6418 (N_6418,N_6143,N_6216);
xor U6419 (N_6419,N_6131,N_5717);
or U6420 (N_6420,N_5913,N_6134);
nand U6421 (N_6421,N_6075,N_5908);
nor U6422 (N_6422,N_5842,N_6177);
nand U6423 (N_6423,N_5663,N_6007);
and U6424 (N_6424,N_5966,N_6217);
and U6425 (N_6425,N_5640,N_5862);
or U6426 (N_6426,N_6000,N_6182);
nor U6427 (N_6427,N_6019,N_6093);
nor U6428 (N_6428,N_6041,N_6202);
or U6429 (N_6429,N_6124,N_5993);
nor U6430 (N_6430,N_5732,N_6199);
xnor U6431 (N_6431,N_6026,N_6119);
xor U6432 (N_6432,N_6023,N_5629);
xor U6433 (N_6433,N_5787,N_5635);
nand U6434 (N_6434,N_5928,N_5755);
xnor U6435 (N_6435,N_5877,N_5698);
nand U6436 (N_6436,N_6033,N_5735);
xor U6437 (N_6437,N_5961,N_6027);
nor U6438 (N_6438,N_6215,N_6235);
xnor U6439 (N_6439,N_5749,N_5888);
nand U6440 (N_6440,N_5823,N_5943);
nor U6441 (N_6441,N_5986,N_6159);
and U6442 (N_6442,N_5797,N_6191);
xnor U6443 (N_6443,N_5708,N_6020);
and U6444 (N_6444,N_6089,N_6148);
nor U6445 (N_6445,N_6201,N_6002);
and U6446 (N_6446,N_5782,N_6112);
xor U6447 (N_6447,N_5801,N_5695);
or U6448 (N_6448,N_5690,N_5924);
and U6449 (N_6449,N_5918,N_5984);
nand U6450 (N_6450,N_5706,N_5884);
xnor U6451 (N_6451,N_5887,N_6016);
nor U6452 (N_6452,N_6105,N_5809);
nor U6453 (N_6453,N_5638,N_6170);
or U6454 (N_6454,N_5837,N_5673);
or U6455 (N_6455,N_5867,N_5784);
and U6456 (N_6456,N_5831,N_6015);
or U6457 (N_6457,N_5958,N_6083);
nor U6458 (N_6458,N_5861,N_5982);
nand U6459 (N_6459,N_5679,N_6060);
nor U6460 (N_6460,N_5970,N_6245);
nor U6461 (N_6461,N_6080,N_6161);
or U6462 (N_6462,N_5626,N_6121);
and U6463 (N_6463,N_6169,N_6097);
xnor U6464 (N_6464,N_5751,N_6211);
xnor U6465 (N_6465,N_6028,N_5791);
and U6466 (N_6466,N_5776,N_5832);
nand U6467 (N_6467,N_5992,N_5671);
nor U6468 (N_6468,N_5929,N_5808);
nor U6469 (N_6469,N_5763,N_6099);
nand U6470 (N_6470,N_6053,N_6040);
or U6471 (N_6471,N_5731,N_5915);
nand U6472 (N_6472,N_5942,N_5678);
nand U6473 (N_6473,N_5703,N_6238);
or U6474 (N_6474,N_6010,N_6146);
nor U6475 (N_6475,N_5975,N_5905);
or U6476 (N_6476,N_6167,N_5721);
and U6477 (N_6477,N_6085,N_5873);
nor U6478 (N_6478,N_5939,N_5853);
nand U6479 (N_6479,N_5744,N_6152);
and U6480 (N_6480,N_5644,N_6240);
and U6481 (N_6481,N_5838,N_5803);
nand U6482 (N_6482,N_6244,N_5866);
or U6483 (N_6483,N_5957,N_5705);
and U6484 (N_6484,N_6006,N_5788);
or U6485 (N_6485,N_5645,N_5697);
xnor U6486 (N_6486,N_6058,N_5637);
xor U6487 (N_6487,N_5807,N_5719);
or U6488 (N_6488,N_5988,N_5779);
xnor U6489 (N_6489,N_6113,N_5921);
nand U6490 (N_6490,N_5858,N_6172);
or U6491 (N_6491,N_5771,N_6061);
nor U6492 (N_6492,N_6048,N_5700);
and U6493 (N_6493,N_5806,N_6066);
or U6494 (N_6494,N_5841,N_5839);
xor U6495 (N_6495,N_6212,N_5693);
xnor U6496 (N_6496,N_6021,N_5734);
and U6497 (N_6497,N_6128,N_5850);
and U6498 (N_6498,N_5758,N_5935);
nor U6499 (N_6499,N_6057,N_5764);
nand U6500 (N_6500,N_5870,N_5767);
and U6501 (N_6501,N_6163,N_5824);
and U6502 (N_6502,N_5688,N_5882);
nor U6503 (N_6503,N_6051,N_5766);
and U6504 (N_6504,N_5851,N_5642);
nor U6505 (N_6505,N_5685,N_5773);
and U6506 (N_6506,N_6187,N_5768);
or U6507 (N_6507,N_5967,N_6181);
or U6508 (N_6508,N_5936,N_6008);
and U6509 (N_6509,N_6063,N_6239);
nor U6510 (N_6510,N_5723,N_5802);
or U6511 (N_6511,N_5972,N_6042);
nor U6512 (N_6512,N_6118,N_5947);
and U6513 (N_6513,N_5686,N_5753);
or U6514 (N_6514,N_6192,N_6198);
nor U6515 (N_6515,N_5810,N_5794);
nand U6516 (N_6516,N_5730,N_5969);
nand U6517 (N_6517,N_5869,N_5896);
nand U6518 (N_6518,N_6154,N_5817);
and U6519 (N_6519,N_6184,N_5715);
xor U6520 (N_6520,N_5737,N_5631);
or U6521 (N_6521,N_5977,N_5691);
or U6522 (N_6522,N_6035,N_6141);
nand U6523 (N_6523,N_5925,N_6036);
nor U6524 (N_6524,N_5746,N_5796);
or U6525 (N_6525,N_6144,N_5894);
and U6526 (N_6526,N_6234,N_5692);
nor U6527 (N_6527,N_6071,N_6092);
nand U6528 (N_6528,N_5628,N_6108);
and U6529 (N_6529,N_5941,N_5835);
nand U6530 (N_6530,N_5740,N_5836);
or U6531 (N_6531,N_5956,N_5871);
nand U6532 (N_6532,N_5661,N_6197);
and U6533 (N_6533,N_6242,N_5811);
nand U6534 (N_6534,N_6203,N_5655);
and U6535 (N_6535,N_5819,N_6049);
nand U6536 (N_6536,N_5639,N_5922);
nand U6537 (N_6537,N_6055,N_5726);
nor U6538 (N_6538,N_6204,N_6229);
xnor U6539 (N_6539,N_5881,N_6086);
nor U6540 (N_6540,N_6237,N_6087);
and U6541 (N_6541,N_5711,N_6004);
nor U6542 (N_6542,N_6243,N_5707);
nor U6543 (N_6543,N_5902,N_5971);
nand U6544 (N_6544,N_6130,N_6220);
or U6545 (N_6545,N_5963,N_5827);
xor U6546 (N_6546,N_5932,N_5641);
xnor U6547 (N_6547,N_5793,N_6158);
nand U6548 (N_6548,N_5893,N_5772);
or U6549 (N_6549,N_5940,N_5770);
or U6550 (N_6550,N_6165,N_5729);
and U6551 (N_6551,N_6127,N_5699);
nand U6552 (N_6552,N_5667,N_6195);
xnor U6553 (N_6553,N_5879,N_5910);
nor U6554 (N_6554,N_6091,N_6228);
or U6555 (N_6555,N_5897,N_5669);
and U6556 (N_6556,N_5840,N_6122);
xor U6557 (N_6557,N_6094,N_5818);
or U6558 (N_6558,N_6101,N_5795);
nand U6559 (N_6559,N_6059,N_5995);
nand U6560 (N_6560,N_5789,N_5872);
nor U6561 (N_6561,N_5748,N_6084);
xor U6562 (N_6562,N_5760,N_6166);
and U6563 (N_6563,N_6064,N_6065);
nand U6564 (N_6564,N_6188,N_5939);
or U6565 (N_6565,N_5874,N_5778);
xor U6566 (N_6566,N_5756,N_5945);
or U6567 (N_6567,N_5987,N_6079);
or U6568 (N_6568,N_5876,N_5896);
xnor U6569 (N_6569,N_5754,N_5749);
nand U6570 (N_6570,N_5752,N_6112);
xor U6571 (N_6571,N_5675,N_6055);
or U6572 (N_6572,N_5722,N_5892);
and U6573 (N_6573,N_6179,N_5885);
nand U6574 (N_6574,N_6049,N_5786);
xnor U6575 (N_6575,N_6116,N_6100);
nand U6576 (N_6576,N_6034,N_5978);
and U6577 (N_6577,N_6169,N_5874);
or U6578 (N_6578,N_5916,N_5823);
and U6579 (N_6579,N_5626,N_6231);
xnor U6580 (N_6580,N_5705,N_5899);
xnor U6581 (N_6581,N_5911,N_5749);
nand U6582 (N_6582,N_6129,N_6019);
nor U6583 (N_6583,N_6223,N_6174);
nor U6584 (N_6584,N_5692,N_5733);
nand U6585 (N_6585,N_6244,N_6148);
nand U6586 (N_6586,N_5744,N_5965);
nor U6587 (N_6587,N_6090,N_5745);
nand U6588 (N_6588,N_5769,N_6014);
or U6589 (N_6589,N_5906,N_6190);
nor U6590 (N_6590,N_5903,N_5775);
nand U6591 (N_6591,N_6169,N_6087);
nand U6592 (N_6592,N_5789,N_6195);
nor U6593 (N_6593,N_6245,N_5703);
nand U6594 (N_6594,N_5911,N_5899);
xor U6595 (N_6595,N_5923,N_5952);
and U6596 (N_6596,N_6066,N_5677);
and U6597 (N_6597,N_6098,N_5819);
or U6598 (N_6598,N_5676,N_5835);
or U6599 (N_6599,N_5664,N_5795);
xnor U6600 (N_6600,N_5735,N_5658);
and U6601 (N_6601,N_6192,N_5951);
nor U6602 (N_6602,N_5966,N_5841);
nor U6603 (N_6603,N_5779,N_6051);
nand U6604 (N_6604,N_5745,N_6116);
or U6605 (N_6605,N_6016,N_5989);
nor U6606 (N_6606,N_5692,N_6164);
or U6607 (N_6607,N_5704,N_6168);
or U6608 (N_6608,N_5999,N_5990);
xnor U6609 (N_6609,N_5729,N_5681);
nand U6610 (N_6610,N_5749,N_5975);
xnor U6611 (N_6611,N_6076,N_5763);
and U6612 (N_6612,N_6107,N_6169);
nand U6613 (N_6613,N_5637,N_5794);
nor U6614 (N_6614,N_5631,N_5752);
nand U6615 (N_6615,N_6010,N_5774);
nand U6616 (N_6616,N_6133,N_5723);
xnor U6617 (N_6617,N_6086,N_6028);
and U6618 (N_6618,N_5727,N_5937);
and U6619 (N_6619,N_5932,N_5783);
and U6620 (N_6620,N_5874,N_6009);
nand U6621 (N_6621,N_6200,N_6132);
nor U6622 (N_6622,N_5826,N_5862);
and U6623 (N_6623,N_5987,N_6164);
nand U6624 (N_6624,N_6021,N_5739);
xnor U6625 (N_6625,N_5802,N_5783);
and U6626 (N_6626,N_5774,N_6212);
or U6627 (N_6627,N_5769,N_5909);
nor U6628 (N_6628,N_6227,N_6024);
and U6629 (N_6629,N_6027,N_5931);
nand U6630 (N_6630,N_5708,N_6050);
and U6631 (N_6631,N_6243,N_5945);
xnor U6632 (N_6632,N_5935,N_5650);
nand U6633 (N_6633,N_5872,N_5962);
xor U6634 (N_6634,N_5948,N_5792);
nor U6635 (N_6635,N_5990,N_5807);
or U6636 (N_6636,N_5740,N_5719);
nor U6637 (N_6637,N_5634,N_5641);
xnor U6638 (N_6638,N_6226,N_5895);
and U6639 (N_6639,N_5630,N_6107);
xor U6640 (N_6640,N_6207,N_5702);
or U6641 (N_6641,N_6035,N_5890);
and U6642 (N_6642,N_5978,N_5765);
xor U6643 (N_6643,N_5853,N_5792);
or U6644 (N_6644,N_6090,N_5646);
or U6645 (N_6645,N_6086,N_5741);
or U6646 (N_6646,N_6034,N_6050);
nor U6647 (N_6647,N_6158,N_5842);
or U6648 (N_6648,N_5847,N_5764);
xnor U6649 (N_6649,N_6092,N_6227);
xnor U6650 (N_6650,N_5903,N_6208);
and U6651 (N_6651,N_5760,N_5913);
nand U6652 (N_6652,N_6119,N_5652);
nor U6653 (N_6653,N_6046,N_5791);
and U6654 (N_6654,N_5858,N_6090);
nor U6655 (N_6655,N_6077,N_5718);
nor U6656 (N_6656,N_5720,N_5656);
xor U6657 (N_6657,N_6231,N_5864);
or U6658 (N_6658,N_6104,N_6153);
or U6659 (N_6659,N_6032,N_6128);
or U6660 (N_6660,N_5836,N_5722);
xnor U6661 (N_6661,N_6043,N_5914);
or U6662 (N_6662,N_5799,N_6102);
and U6663 (N_6663,N_5866,N_5773);
or U6664 (N_6664,N_5899,N_5989);
nand U6665 (N_6665,N_6089,N_6068);
and U6666 (N_6666,N_5740,N_6126);
nand U6667 (N_6667,N_5876,N_5798);
nor U6668 (N_6668,N_5774,N_5736);
and U6669 (N_6669,N_6018,N_6147);
nor U6670 (N_6670,N_6088,N_6084);
and U6671 (N_6671,N_5652,N_6192);
xnor U6672 (N_6672,N_6107,N_5741);
xnor U6673 (N_6673,N_6223,N_5752);
nor U6674 (N_6674,N_5734,N_5673);
or U6675 (N_6675,N_6156,N_5692);
or U6676 (N_6676,N_5966,N_5769);
xnor U6677 (N_6677,N_5691,N_5805);
or U6678 (N_6678,N_6084,N_5813);
xnor U6679 (N_6679,N_6200,N_6038);
xor U6680 (N_6680,N_6144,N_6201);
or U6681 (N_6681,N_5883,N_6160);
nand U6682 (N_6682,N_6072,N_6024);
and U6683 (N_6683,N_6101,N_5696);
nor U6684 (N_6684,N_5899,N_6207);
xor U6685 (N_6685,N_6242,N_6148);
nor U6686 (N_6686,N_5842,N_6142);
nand U6687 (N_6687,N_5976,N_6155);
nor U6688 (N_6688,N_5899,N_5875);
xnor U6689 (N_6689,N_6204,N_5844);
nand U6690 (N_6690,N_6016,N_6062);
nand U6691 (N_6691,N_6062,N_6226);
or U6692 (N_6692,N_5685,N_5961);
nand U6693 (N_6693,N_5760,N_5939);
or U6694 (N_6694,N_6109,N_5902);
or U6695 (N_6695,N_5935,N_5925);
xnor U6696 (N_6696,N_6132,N_5960);
xnor U6697 (N_6697,N_5886,N_6205);
or U6698 (N_6698,N_6107,N_6235);
nor U6699 (N_6699,N_5977,N_6234);
xnor U6700 (N_6700,N_5920,N_6147);
nor U6701 (N_6701,N_6115,N_6110);
nor U6702 (N_6702,N_5971,N_6038);
nor U6703 (N_6703,N_6040,N_5929);
nand U6704 (N_6704,N_5744,N_5920);
or U6705 (N_6705,N_5993,N_6037);
and U6706 (N_6706,N_5718,N_6104);
nor U6707 (N_6707,N_6162,N_6016);
nand U6708 (N_6708,N_6152,N_6110);
nor U6709 (N_6709,N_6166,N_6130);
xor U6710 (N_6710,N_5717,N_6116);
nor U6711 (N_6711,N_5731,N_6080);
nor U6712 (N_6712,N_6040,N_6162);
or U6713 (N_6713,N_5682,N_5748);
or U6714 (N_6714,N_6238,N_5805);
nor U6715 (N_6715,N_6176,N_5856);
nand U6716 (N_6716,N_5790,N_5686);
nor U6717 (N_6717,N_5766,N_5733);
xnor U6718 (N_6718,N_6172,N_5724);
nand U6719 (N_6719,N_5637,N_5719);
nand U6720 (N_6720,N_6017,N_6212);
xnor U6721 (N_6721,N_6249,N_5663);
nor U6722 (N_6722,N_6192,N_5828);
or U6723 (N_6723,N_5921,N_5923);
nand U6724 (N_6724,N_6036,N_6114);
nor U6725 (N_6725,N_5746,N_6234);
and U6726 (N_6726,N_6178,N_6204);
and U6727 (N_6727,N_6048,N_5863);
xor U6728 (N_6728,N_5972,N_5832);
or U6729 (N_6729,N_5788,N_5957);
or U6730 (N_6730,N_5856,N_6186);
and U6731 (N_6731,N_5902,N_5788);
nor U6732 (N_6732,N_5974,N_5668);
and U6733 (N_6733,N_5816,N_5860);
and U6734 (N_6734,N_5685,N_6046);
nor U6735 (N_6735,N_5845,N_5954);
nand U6736 (N_6736,N_6175,N_6113);
nand U6737 (N_6737,N_5866,N_6101);
or U6738 (N_6738,N_5960,N_5703);
or U6739 (N_6739,N_5950,N_6174);
and U6740 (N_6740,N_6197,N_6094);
nor U6741 (N_6741,N_5653,N_5898);
and U6742 (N_6742,N_5889,N_5652);
and U6743 (N_6743,N_5872,N_6173);
and U6744 (N_6744,N_6084,N_5809);
and U6745 (N_6745,N_6124,N_5958);
nand U6746 (N_6746,N_5883,N_5722);
nor U6747 (N_6747,N_5722,N_6176);
xnor U6748 (N_6748,N_5916,N_5917);
nor U6749 (N_6749,N_5888,N_6048);
nor U6750 (N_6750,N_5655,N_5654);
xnor U6751 (N_6751,N_5940,N_6035);
nor U6752 (N_6752,N_6135,N_6147);
and U6753 (N_6753,N_5905,N_6198);
xnor U6754 (N_6754,N_5867,N_5803);
or U6755 (N_6755,N_5713,N_6122);
nor U6756 (N_6756,N_6164,N_6241);
or U6757 (N_6757,N_6121,N_6190);
or U6758 (N_6758,N_6151,N_6245);
and U6759 (N_6759,N_5930,N_5706);
xor U6760 (N_6760,N_6243,N_6005);
nand U6761 (N_6761,N_6141,N_5911);
and U6762 (N_6762,N_6118,N_5754);
xor U6763 (N_6763,N_5887,N_5923);
nor U6764 (N_6764,N_5837,N_6140);
nor U6765 (N_6765,N_6044,N_5939);
xor U6766 (N_6766,N_6091,N_5794);
nand U6767 (N_6767,N_6100,N_6207);
nand U6768 (N_6768,N_6190,N_5805);
or U6769 (N_6769,N_5682,N_6201);
or U6770 (N_6770,N_6176,N_5626);
and U6771 (N_6771,N_6207,N_6187);
nand U6772 (N_6772,N_5675,N_5690);
nand U6773 (N_6773,N_6172,N_5663);
nand U6774 (N_6774,N_5707,N_5741);
and U6775 (N_6775,N_6141,N_6019);
nand U6776 (N_6776,N_6136,N_6111);
and U6777 (N_6777,N_5683,N_6008);
or U6778 (N_6778,N_6059,N_5713);
or U6779 (N_6779,N_6134,N_5943);
nor U6780 (N_6780,N_5724,N_6024);
nor U6781 (N_6781,N_5717,N_6047);
nor U6782 (N_6782,N_5692,N_5792);
nand U6783 (N_6783,N_5769,N_5716);
nor U6784 (N_6784,N_5970,N_6145);
xnor U6785 (N_6785,N_5766,N_5943);
and U6786 (N_6786,N_5661,N_6088);
and U6787 (N_6787,N_5901,N_5836);
nor U6788 (N_6788,N_6105,N_5763);
nand U6789 (N_6789,N_6120,N_6148);
or U6790 (N_6790,N_6175,N_6214);
xnor U6791 (N_6791,N_6002,N_6111);
xnor U6792 (N_6792,N_5989,N_5681);
xnor U6793 (N_6793,N_5671,N_5873);
nor U6794 (N_6794,N_5921,N_5813);
and U6795 (N_6795,N_6209,N_5907);
nand U6796 (N_6796,N_5805,N_5926);
nor U6797 (N_6797,N_6180,N_5817);
or U6798 (N_6798,N_5629,N_6154);
and U6799 (N_6799,N_5711,N_5898);
and U6800 (N_6800,N_5694,N_6181);
nor U6801 (N_6801,N_5900,N_5970);
nor U6802 (N_6802,N_6027,N_6025);
nand U6803 (N_6803,N_6118,N_5800);
and U6804 (N_6804,N_6202,N_5792);
and U6805 (N_6805,N_6012,N_6046);
nand U6806 (N_6806,N_5648,N_5815);
xor U6807 (N_6807,N_5947,N_5808);
and U6808 (N_6808,N_6114,N_6085);
nor U6809 (N_6809,N_5695,N_5666);
nor U6810 (N_6810,N_5992,N_5896);
xnor U6811 (N_6811,N_5659,N_5713);
and U6812 (N_6812,N_5758,N_5789);
or U6813 (N_6813,N_5819,N_6181);
and U6814 (N_6814,N_6175,N_5906);
and U6815 (N_6815,N_6015,N_5669);
nor U6816 (N_6816,N_6133,N_6171);
nor U6817 (N_6817,N_5772,N_5627);
xnor U6818 (N_6818,N_6068,N_5660);
and U6819 (N_6819,N_5698,N_6071);
or U6820 (N_6820,N_6057,N_5754);
xor U6821 (N_6821,N_5806,N_5756);
nor U6822 (N_6822,N_5718,N_6079);
or U6823 (N_6823,N_6014,N_6163);
and U6824 (N_6824,N_6106,N_5627);
xor U6825 (N_6825,N_5752,N_6016);
and U6826 (N_6826,N_6130,N_5869);
and U6827 (N_6827,N_5896,N_5945);
nand U6828 (N_6828,N_5677,N_6187);
and U6829 (N_6829,N_5871,N_5845);
or U6830 (N_6830,N_5764,N_6117);
nand U6831 (N_6831,N_5935,N_5869);
xnor U6832 (N_6832,N_6169,N_6076);
nor U6833 (N_6833,N_6069,N_5646);
xor U6834 (N_6834,N_5746,N_5834);
and U6835 (N_6835,N_6196,N_6247);
xor U6836 (N_6836,N_5716,N_5897);
nor U6837 (N_6837,N_6164,N_5899);
and U6838 (N_6838,N_5660,N_5695);
nand U6839 (N_6839,N_6167,N_6104);
xor U6840 (N_6840,N_6002,N_5858);
or U6841 (N_6841,N_5973,N_5872);
nor U6842 (N_6842,N_6175,N_6073);
nand U6843 (N_6843,N_6038,N_5713);
xnor U6844 (N_6844,N_6044,N_5730);
or U6845 (N_6845,N_5957,N_5821);
xor U6846 (N_6846,N_5728,N_6066);
xor U6847 (N_6847,N_6056,N_6125);
nor U6848 (N_6848,N_6103,N_5971);
or U6849 (N_6849,N_6015,N_5956);
and U6850 (N_6850,N_5687,N_6204);
or U6851 (N_6851,N_6081,N_5933);
or U6852 (N_6852,N_5690,N_5834);
nor U6853 (N_6853,N_5808,N_5662);
nand U6854 (N_6854,N_6086,N_6236);
xor U6855 (N_6855,N_6037,N_6162);
and U6856 (N_6856,N_5926,N_6194);
nand U6857 (N_6857,N_5902,N_5913);
and U6858 (N_6858,N_5915,N_6033);
nand U6859 (N_6859,N_6113,N_6223);
nand U6860 (N_6860,N_5954,N_6135);
nand U6861 (N_6861,N_6108,N_5876);
xor U6862 (N_6862,N_6117,N_5718);
xnor U6863 (N_6863,N_5677,N_6046);
nand U6864 (N_6864,N_5979,N_5906);
xor U6865 (N_6865,N_5989,N_6137);
and U6866 (N_6866,N_6192,N_5985);
or U6867 (N_6867,N_6045,N_6018);
and U6868 (N_6868,N_6244,N_5808);
nand U6869 (N_6869,N_6203,N_5904);
or U6870 (N_6870,N_5955,N_5791);
or U6871 (N_6871,N_6080,N_6078);
nor U6872 (N_6872,N_5727,N_5667);
xor U6873 (N_6873,N_5816,N_6121);
nand U6874 (N_6874,N_5977,N_5805);
nand U6875 (N_6875,N_6699,N_6641);
or U6876 (N_6876,N_6677,N_6655);
nor U6877 (N_6877,N_6381,N_6346);
xor U6878 (N_6878,N_6251,N_6866);
or U6879 (N_6879,N_6874,N_6706);
nand U6880 (N_6880,N_6370,N_6290);
xor U6881 (N_6881,N_6653,N_6808);
nand U6882 (N_6882,N_6562,N_6661);
xor U6883 (N_6883,N_6293,N_6263);
nor U6884 (N_6884,N_6681,N_6329);
and U6885 (N_6885,N_6621,N_6578);
nor U6886 (N_6886,N_6851,N_6532);
nand U6887 (N_6887,N_6734,N_6516);
nand U6888 (N_6888,N_6524,N_6745);
and U6889 (N_6889,N_6482,N_6485);
or U6890 (N_6890,N_6719,N_6644);
nand U6891 (N_6891,N_6404,N_6519);
nor U6892 (N_6892,N_6702,N_6441);
and U6893 (N_6893,N_6316,N_6758);
or U6894 (N_6894,N_6791,N_6725);
xnor U6895 (N_6895,N_6318,N_6757);
or U6896 (N_6896,N_6774,N_6576);
xnor U6897 (N_6897,N_6543,N_6304);
nand U6898 (N_6898,N_6744,N_6609);
nor U6899 (N_6899,N_6669,N_6600);
or U6900 (N_6900,N_6623,N_6267);
nor U6901 (N_6901,N_6255,N_6831);
or U6902 (N_6902,N_6473,N_6793);
xnor U6903 (N_6903,N_6338,N_6559);
or U6904 (N_6904,N_6280,N_6646);
nor U6905 (N_6905,N_6515,N_6872);
nor U6906 (N_6906,N_6588,N_6358);
and U6907 (N_6907,N_6738,N_6612);
or U6908 (N_6908,N_6603,N_6323);
xnor U6909 (N_6909,N_6778,N_6460);
nand U6910 (N_6910,N_6801,N_6579);
xor U6911 (N_6911,N_6788,N_6514);
nand U6912 (N_6912,N_6683,N_6818);
xnor U6913 (N_6913,N_6393,N_6360);
xnor U6914 (N_6914,N_6703,N_6488);
or U6915 (N_6915,N_6447,N_6815);
xor U6916 (N_6916,N_6637,N_6635);
nand U6917 (N_6917,N_6610,N_6762);
nor U6918 (N_6918,N_6523,N_6763);
nor U6919 (N_6919,N_6281,N_6504);
nand U6920 (N_6920,N_6567,N_6313);
xor U6921 (N_6921,N_6387,N_6792);
nor U6922 (N_6922,N_6396,N_6326);
and U6923 (N_6923,N_6401,N_6727);
nor U6924 (N_6924,N_6604,N_6265);
nand U6925 (N_6925,N_6771,N_6794);
or U6926 (N_6926,N_6707,N_6333);
nand U6927 (N_6927,N_6695,N_6282);
or U6928 (N_6928,N_6581,N_6736);
nand U6929 (N_6929,N_6746,N_6419);
nand U6930 (N_6930,N_6841,N_6619);
nor U6931 (N_6931,N_6735,N_6849);
nor U6932 (N_6932,N_6608,N_6638);
nor U6933 (N_6933,N_6493,N_6781);
nand U6934 (N_6934,N_6420,N_6310);
xor U6935 (N_6935,N_6498,N_6747);
and U6936 (N_6936,N_6779,N_6691);
or U6937 (N_6937,N_6446,N_6479);
nand U6938 (N_6938,N_6806,N_6795);
nor U6939 (N_6939,N_6714,N_6631);
nor U6940 (N_6940,N_6303,N_6723);
xor U6941 (N_6941,N_6667,N_6713);
xnor U6942 (N_6942,N_6803,N_6258);
nand U6943 (N_6943,N_6555,N_6327);
nor U6944 (N_6944,N_6798,N_6508);
and U6945 (N_6945,N_6787,N_6395);
xnor U6946 (N_6946,N_6607,N_6440);
or U6947 (N_6947,N_6595,N_6693);
nor U6948 (N_6948,N_6520,N_6606);
and U6949 (N_6949,N_6306,N_6585);
or U6950 (N_6950,N_6495,N_6605);
nor U6951 (N_6951,N_6743,N_6668);
xnor U6952 (N_6952,N_6843,N_6477);
nand U6953 (N_6953,N_6648,N_6569);
and U6954 (N_6954,N_6785,N_6535);
and U6955 (N_6955,N_6406,N_6348);
and U6956 (N_6956,N_6853,N_6690);
nand U6957 (N_6957,N_6299,N_6616);
nand U6958 (N_6958,N_6867,N_6686);
and U6959 (N_6959,N_6461,N_6542);
nand U6960 (N_6960,N_6362,N_6522);
or U6961 (N_6961,N_6528,N_6278);
and U6962 (N_6962,N_6259,N_6587);
or U6963 (N_6963,N_6636,N_6368);
or U6964 (N_6964,N_6730,N_6764);
nand U6965 (N_6965,N_6413,N_6659);
and U6966 (N_6966,N_6343,N_6268);
nor U6967 (N_6967,N_6846,N_6684);
nor U6968 (N_6968,N_6257,N_6314);
nand U6969 (N_6969,N_6852,N_6620);
xor U6970 (N_6970,N_6742,N_6652);
nor U6971 (N_6971,N_6674,N_6296);
or U6972 (N_6972,N_6311,N_6836);
or U6973 (N_6973,N_6570,N_6463);
and U6974 (N_6974,N_6422,N_6740);
xnor U6975 (N_6975,N_6692,N_6317);
nand U6976 (N_6976,N_6383,N_6300);
and U6977 (N_6977,N_6283,N_6642);
nand U6978 (N_6978,N_6573,N_6708);
and U6979 (N_6979,N_6390,N_6301);
xor U6980 (N_6980,N_6544,N_6591);
and U6981 (N_6981,N_6733,N_6676);
and U6982 (N_6982,N_6782,N_6731);
xor U6983 (N_6983,N_6525,N_6826);
or U6984 (N_6984,N_6371,N_6494);
or U6985 (N_6985,N_6513,N_6860);
or U6986 (N_6986,N_6364,N_6429);
nand U6987 (N_6987,N_6536,N_6672);
nor U6988 (N_6988,N_6855,N_6339);
or U6989 (N_6989,N_6698,N_6469);
or U6990 (N_6990,N_6820,N_6700);
xnor U6991 (N_6991,N_6353,N_6583);
and U6992 (N_6992,N_6505,N_6799);
nand U6993 (N_6993,N_6537,N_6614);
xor U6994 (N_6994,N_6720,N_6776);
nand U6995 (N_6995,N_6431,N_6250);
or U6996 (N_6996,N_6775,N_6835);
and U6997 (N_6997,N_6709,N_6320);
nor U6998 (N_6998,N_6418,N_6470);
xnor U6999 (N_6999,N_6858,N_6483);
or U7000 (N_7000,N_6434,N_6292);
nand U7001 (N_7001,N_6445,N_6710);
nor U7002 (N_7002,N_6496,N_6398);
nand U7003 (N_7003,N_6366,N_6597);
nand U7004 (N_7004,N_6666,N_6718);
nor U7005 (N_7005,N_6444,N_6436);
and U7006 (N_7006,N_6540,N_6832);
xnor U7007 (N_7007,N_6466,N_6545);
and U7008 (N_7008,N_6269,N_6367);
and U7009 (N_7009,N_6767,N_6298);
nand U7010 (N_7010,N_6856,N_6673);
nand U7011 (N_7011,N_6722,N_6392);
nor U7012 (N_7012,N_6384,N_6601);
xor U7013 (N_7013,N_6768,N_6582);
nand U7014 (N_7014,N_6550,N_6405);
nor U7015 (N_7015,N_6816,N_6772);
nor U7016 (N_7016,N_6837,N_6862);
nand U7017 (N_7017,N_6751,N_6685);
nand U7018 (N_7018,N_6340,N_6696);
or U7019 (N_7019,N_6594,N_6334);
and U7020 (N_7020,N_6554,N_6748);
nor U7021 (N_7021,N_6511,N_6380);
and U7022 (N_7022,N_6671,N_6256);
nor U7023 (N_7023,N_6342,N_6427);
or U7024 (N_7024,N_6486,N_6819);
nor U7025 (N_7025,N_6432,N_6593);
nor U7026 (N_7026,N_6321,N_6344);
or U7027 (N_7027,N_6552,N_6632);
nand U7028 (N_7028,N_6752,N_6489);
or U7029 (N_7029,N_6639,N_6551);
nor U7030 (N_7030,N_6805,N_6332);
nor U7031 (N_7031,N_6662,N_6500);
nand U7032 (N_7032,N_6679,N_6421);
xnor U7033 (N_7033,N_6359,N_6560);
nor U7034 (N_7034,N_6732,N_6739);
xnor U7035 (N_7035,N_6870,N_6821);
nand U7036 (N_7036,N_6454,N_6665);
or U7037 (N_7037,N_6331,N_6789);
nand U7038 (N_7038,N_6471,N_6721);
nand U7039 (N_7039,N_6277,N_6497);
and U7040 (N_7040,N_6307,N_6760);
nand U7041 (N_7041,N_6645,N_6330);
or U7042 (N_7042,N_6625,N_6840);
nor U7043 (N_7043,N_6602,N_6487);
nor U7044 (N_7044,N_6628,N_6842);
nor U7045 (N_7045,N_6548,N_6319);
nor U7046 (N_7046,N_6354,N_6556);
or U7047 (N_7047,N_6351,N_6811);
nand U7048 (N_7048,N_6272,N_6825);
xnor U7049 (N_7049,N_6561,N_6571);
xnor U7050 (N_7050,N_6424,N_6412);
nor U7051 (N_7051,N_6823,N_6834);
xnor U7052 (N_7052,N_6449,N_6481);
nand U7053 (N_7053,N_6517,N_6577);
nand U7054 (N_7054,N_6357,N_6688);
nor U7055 (N_7055,N_6812,N_6388);
and U7056 (N_7056,N_6617,N_6575);
nand U7057 (N_7057,N_6833,N_6822);
and U7058 (N_7058,N_6759,N_6848);
nor U7059 (N_7059,N_6780,N_6270);
and U7060 (N_7060,N_6385,N_6572);
nor U7061 (N_7061,N_6375,N_6379);
xnor U7062 (N_7062,N_6309,N_6506);
and U7063 (N_7063,N_6724,N_6262);
nor U7064 (N_7064,N_6455,N_6557);
xnor U7065 (N_7065,N_6715,N_6804);
or U7066 (N_7066,N_6417,N_6654);
and U7067 (N_7067,N_6374,N_6527);
or U7068 (N_7068,N_6288,N_6618);
xnor U7069 (N_7069,N_6664,N_6765);
and U7070 (N_7070,N_6786,N_6783);
or U7071 (N_7071,N_6450,N_6302);
nand U7072 (N_7072,N_6287,N_6408);
nor U7073 (N_7073,N_6467,N_6650);
nand U7074 (N_7074,N_6297,N_6274);
and U7075 (N_7075,N_6503,N_6538);
xor U7076 (N_7076,N_6361,N_6402);
and U7077 (N_7077,N_6439,N_6491);
or U7078 (N_7078,N_6480,N_6324);
nor U7079 (N_7079,N_6871,N_6711);
xor U7080 (N_7080,N_6397,N_6291);
or U7081 (N_7081,N_6328,N_6830);
or U7082 (N_7082,N_6337,N_6626);
or U7083 (N_7083,N_6531,N_6430);
nor U7084 (N_7084,N_6425,N_6356);
or U7085 (N_7085,N_6378,N_6717);
or U7086 (N_7086,N_6629,N_6844);
xor U7087 (N_7087,N_6873,N_6868);
and U7088 (N_7088,N_6634,N_6802);
or U7089 (N_7089,N_6284,N_6589);
xor U7090 (N_7090,N_6474,N_6777);
and U7091 (N_7091,N_6526,N_6761);
and U7092 (N_7092,N_6660,N_6464);
and U7093 (N_7093,N_6701,N_6415);
nor U7094 (N_7094,N_6435,N_6428);
or U7095 (N_7095,N_6458,N_6729);
nor U7096 (N_7096,N_6512,N_6426);
nand U7097 (N_7097,N_6549,N_6847);
or U7098 (N_7098,N_6814,N_6295);
nor U7099 (N_7099,N_6433,N_6423);
nor U7100 (N_7100,N_6737,N_6754);
and U7101 (N_7101,N_6838,N_6845);
xor U7102 (N_7102,N_6712,N_6452);
or U7103 (N_7103,N_6462,N_6565);
nand U7104 (N_7104,N_6409,N_6275);
nand U7105 (N_7105,N_6689,N_6694);
xnor U7106 (N_7106,N_6365,N_6649);
and U7107 (N_7107,N_6350,N_6682);
and U7108 (N_7108,N_6566,N_6382);
xor U7109 (N_7109,N_6643,N_6797);
and U7110 (N_7110,N_6501,N_6502);
nand U7111 (N_7111,N_6657,N_6615);
nor U7112 (N_7112,N_6530,N_6564);
nor U7113 (N_7113,N_6854,N_6704);
xnor U7114 (N_7114,N_6766,N_6266);
and U7115 (N_7115,N_6271,N_6824);
nor U7116 (N_7116,N_6534,N_6443);
or U7117 (N_7117,N_6386,N_6558);
and U7118 (N_7118,N_6864,N_6322);
xor U7119 (N_7119,N_6574,N_6391);
or U7120 (N_7120,N_6741,N_6622);
nor U7121 (N_7121,N_6411,N_6325);
nor U7122 (N_7122,N_6305,N_6663);
nand U7123 (N_7123,N_6539,N_6336);
or U7124 (N_7124,N_6475,N_6349);
or U7125 (N_7125,N_6790,N_6403);
or U7126 (N_7126,N_6770,N_6457);
nor U7127 (N_7127,N_6753,N_6533);
nor U7128 (N_7128,N_6437,N_6264);
xor U7129 (N_7129,N_6658,N_6400);
and U7130 (N_7130,N_6553,N_6547);
xnor U7131 (N_7131,N_6613,N_6451);
or U7132 (N_7132,N_6252,N_6509);
xor U7133 (N_7133,N_6347,N_6254);
or U7134 (N_7134,N_6651,N_6563);
and U7135 (N_7135,N_6341,N_6352);
and U7136 (N_7136,N_6492,N_6670);
xnor U7137 (N_7137,N_6859,N_6315);
or U7138 (N_7138,N_6599,N_6373);
or U7139 (N_7139,N_6376,N_6499);
nand U7140 (N_7140,N_6453,N_6442);
and U7141 (N_7141,N_6468,N_6773);
and U7142 (N_7142,N_6507,N_6656);
and U7143 (N_7143,N_6286,N_6518);
nor U7144 (N_7144,N_6372,N_6410);
and U7145 (N_7145,N_6448,N_6705);
or U7146 (N_7146,N_6716,N_6726);
nand U7147 (N_7147,N_6827,N_6546);
xor U7148 (N_7148,N_6817,N_6529);
nand U7149 (N_7149,N_6586,N_6438);
and U7150 (N_7150,N_6389,N_6465);
or U7151 (N_7151,N_6394,N_6828);
xor U7152 (N_7152,N_6407,N_6647);
or U7153 (N_7153,N_6261,N_6809);
nor U7154 (N_7154,N_6580,N_6624);
or U7155 (N_7155,N_6633,N_6829);
or U7156 (N_7156,N_6335,N_6478);
or U7157 (N_7157,N_6355,N_6416);
nor U7158 (N_7158,N_6279,N_6627);
xor U7159 (N_7159,N_6800,N_6850);
and U7160 (N_7160,N_6796,N_6697);
and U7161 (N_7161,N_6861,N_6728);
xor U7162 (N_7162,N_6630,N_6510);
xor U7163 (N_7163,N_6592,N_6289);
nor U7164 (N_7164,N_6584,N_6839);
or U7165 (N_7165,N_6456,N_6459);
xnor U7166 (N_7166,N_6541,N_6260);
xor U7167 (N_7167,N_6414,N_6640);
nand U7168 (N_7168,N_6294,N_6399);
and U7169 (N_7169,N_6784,N_6869);
nor U7170 (N_7170,N_6285,N_6308);
or U7171 (N_7171,N_6678,N_6377);
xnor U7172 (N_7172,N_6611,N_6521);
xor U7173 (N_7173,N_6749,N_6276);
xnor U7174 (N_7174,N_6472,N_6476);
xnor U7175 (N_7175,N_6865,N_6598);
and U7176 (N_7176,N_6813,N_6675);
or U7177 (N_7177,N_6687,N_6312);
and U7178 (N_7178,N_6857,N_6810);
xnor U7179 (N_7179,N_6680,N_6750);
and U7180 (N_7180,N_6484,N_6596);
or U7181 (N_7181,N_6863,N_6253);
xnor U7182 (N_7182,N_6769,N_6755);
xor U7183 (N_7183,N_6568,N_6369);
and U7184 (N_7184,N_6590,N_6490);
nor U7185 (N_7185,N_6345,N_6273);
or U7186 (N_7186,N_6756,N_6807);
and U7187 (N_7187,N_6363,N_6395);
xor U7188 (N_7188,N_6498,N_6572);
nand U7189 (N_7189,N_6488,N_6371);
nand U7190 (N_7190,N_6264,N_6284);
and U7191 (N_7191,N_6639,N_6662);
or U7192 (N_7192,N_6383,N_6723);
xnor U7193 (N_7193,N_6770,N_6658);
or U7194 (N_7194,N_6808,N_6449);
nand U7195 (N_7195,N_6493,N_6341);
xor U7196 (N_7196,N_6667,N_6734);
nand U7197 (N_7197,N_6486,N_6411);
or U7198 (N_7198,N_6483,N_6353);
xor U7199 (N_7199,N_6669,N_6775);
and U7200 (N_7200,N_6473,N_6624);
or U7201 (N_7201,N_6641,N_6640);
or U7202 (N_7202,N_6494,N_6696);
and U7203 (N_7203,N_6612,N_6264);
or U7204 (N_7204,N_6333,N_6473);
xnor U7205 (N_7205,N_6449,N_6419);
xnor U7206 (N_7206,N_6518,N_6351);
xnor U7207 (N_7207,N_6727,N_6655);
nor U7208 (N_7208,N_6594,N_6351);
nand U7209 (N_7209,N_6369,N_6608);
or U7210 (N_7210,N_6823,N_6497);
or U7211 (N_7211,N_6710,N_6424);
and U7212 (N_7212,N_6347,N_6778);
or U7213 (N_7213,N_6554,N_6423);
or U7214 (N_7214,N_6574,N_6682);
nor U7215 (N_7215,N_6427,N_6636);
nor U7216 (N_7216,N_6648,N_6268);
or U7217 (N_7217,N_6389,N_6599);
nand U7218 (N_7218,N_6517,N_6690);
xnor U7219 (N_7219,N_6513,N_6268);
nand U7220 (N_7220,N_6774,N_6480);
or U7221 (N_7221,N_6397,N_6483);
xnor U7222 (N_7222,N_6853,N_6523);
or U7223 (N_7223,N_6528,N_6650);
and U7224 (N_7224,N_6454,N_6261);
nand U7225 (N_7225,N_6404,N_6324);
xor U7226 (N_7226,N_6610,N_6384);
xnor U7227 (N_7227,N_6859,N_6621);
and U7228 (N_7228,N_6521,N_6671);
nand U7229 (N_7229,N_6809,N_6773);
and U7230 (N_7230,N_6728,N_6659);
or U7231 (N_7231,N_6692,N_6343);
or U7232 (N_7232,N_6647,N_6781);
xor U7233 (N_7233,N_6454,N_6545);
and U7234 (N_7234,N_6491,N_6266);
nor U7235 (N_7235,N_6308,N_6275);
nand U7236 (N_7236,N_6575,N_6568);
xor U7237 (N_7237,N_6561,N_6624);
or U7238 (N_7238,N_6763,N_6566);
or U7239 (N_7239,N_6276,N_6750);
or U7240 (N_7240,N_6570,N_6613);
or U7241 (N_7241,N_6404,N_6747);
nor U7242 (N_7242,N_6350,N_6628);
and U7243 (N_7243,N_6417,N_6521);
nor U7244 (N_7244,N_6683,N_6437);
nand U7245 (N_7245,N_6560,N_6357);
nor U7246 (N_7246,N_6480,N_6487);
and U7247 (N_7247,N_6798,N_6320);
or U7248 (N_7248,N_6836,N_6764);
and U7249 (N_7249,N_6446,N_6573);
nand U7250 (N_7250,N_6274,N_6518);
and U7251 (N_7251,N_6331,N_6798);
and U7252 (N_7252,N_6420,N_6349);
or U7253 (N_7253,N_6321,N_6420);
nor U7254 (N_7254,N_6588,N_6338);
nand U7255 (N_7255,N_6657,N_6465);
and U7256 (N_7256,N_6472,N_6548);
nor U7257 (N_7257,N_6464,N_6573);
nand U7258 (N_7258,N_6365,N_6820);
nand U7259 (N_7259,N_6595,N_6539);
and U7260 (N_7260,N_6394,N_6399);
nand U7261 (N_7261,N_6609,N_6486);
or U7262 (N_7262,N_6613,N_6326);
or U7263 (N_7263,N_6854,N_6481);
and U7264 (N_7264,N_6301,N_6411);
nand U7265 (N_7265,N_6800,N_6724);
nand U7266 (N_7266,N_6804,N_6262);
nor U7267 (N_7267,N_6737,N_6461);
or U7268 (N_7268,N_6759,N_6660);
xor U7269 (N_7269,N_6736,N_6600);
xor U7270 (N_7270,N_6598,N_6784);
nor U7271 (N_7271,N_6508,N_6397);
nor U7272 (N_7272,N_6799,N_6840);
xor U7273 (N_7273,N_6822,N_6611);
xor U7274 (N_7274,N_6601,N_6289);
nand U7275 (N_7275,N_6636,N_6852);
nand U7276 (N_7276,N_6820,N_6610);
and U7277 (N_7277,N_6657,N_6400);
or U7278 (N_7278,N_6375,N_6480);
nor U7279 (N_7279,N_6791,N_6414);
xnor U7280 (N_7280,N_6283,N_6467);
and U7281 (N_7281,N_6674,N_6857);
xnor U7282 (N_7282,N_6609,N_6417);
nand U7283 (N_7283,N_6513,N_6740);
or U7284 (N_7284,N_6688,N_6820);
nand U7285 (N_7285,N_6381,N_6296);
and U7286 (N_7286,N_6785,N_6650);
nand U7287 (N_7287,N_6554,N_6766);
nor U7288 (N_7288,N_6817,N_6839);
or U7289 (N_7289,N_6746,N_6332);
or U7290 (N_7290,N_6405,N_6542);
and U7291 (N_7291,N_6498,N_6402);
and U7292 (N_7292,N_6368,N_6722);
xor U7293 (N_7293,N_6598,N_6652);
xnor U7294 (N_7294,N_6852,N_6382);
or U7295 (N_7295,N_6587,N_6840);
and U7296 (N_7296,N_6299,N_6815);
or U7297 (N_7297,N_6320,N_6797);
or U7298 (N_7298,N_6434,N_6795);
or U7299 (N_7299,N_6874,N_6376);
nor U7300 (N_7300,N_6488,N_6272);
or U7301 (N_7301,N_6679,N_6365);
and U7302 (N_7302,N_6373,N_6611);
or U7303 (N_7303,N_6277,N_6265);
nand U7304 (N_7304,N_6550,N_6258);
and U7305 (N_7305,N_6285,N_6587);
and U7306 (N_7306,N_6790,N_6769);
nand U7307 (N_7307,N_6836,N_6819);
nor U7308 (N_7308,N_6568,N_6755);
nand U7309 (N_7309,N_6486,N_6835);
nand U7310 (N_7310,N_6839,N_6868);
nor U7311 (N_7311,N_6374,N_6383);
xor U7312 (N_7312,N_6670,N_6701);
nor U7313 (N_7313,N_6683,N_6705);
nor U7314 (N_7314,N_6791,N_6702);
or U7315 (N_7315,N_6843,N_6525);
or U7316 (N_7316,N_6467,N_6674);
nor U7317 (N_7317,N_6787,N_6692);
and U7318 (N_7318,N_6663,N_6317);
or U7319 (N_7319,N_6467,N_6438);
nor U7320 (N_7320,N_6715,N_6774);
and U7321 (N_7321,N_6311,N_6308);
or U7322 (N_7322,N_6418,N_6812);
or U7323 (N_7323,N_6385,N_6740);
or U7324 (N_7324,N_6805,N_6756);
nand U7325 (N_7325,N_6333,N_6606);
nor U7326 (N_7326,N_6252,N_6561);
nand U7327 (N_7327,N_6780,N_6576);
nor U7328 (N_7328,N_6422,N_6836);
nor U7329 (N_7329,N_6670,N_6778);
nor U7330 (N_7330,N_6853,N_6857);
or U7331 (N_7331,N_6773,N_6254);
and U7332 (N_7332,N_6255,N_6325);
or U7333 (N_7333,N_6856,N_6779);
nand U7334 (N_7334,N_6688,N_6674);
nand U7335 (N_7335,N_6480,N_6745);
and U7336 (N_7336,N_6540,N_6718);
and U7337 (N_7337,N_6789,N_6753);
xor U7338 (N_7338,N_6461,N_6854);
nor U7339 (N_7339,N_6341,N_6555);
nand U7340 (N_7340,N_6697,N_6311);
nand U7341 (N_7341,N_6844,N_6673);
xnor U7342 (N_7342,N_6671,N_6365);
or U7343 (N_7343,N_6250,N_6628);
and U7344 (N_7344,N_6515,N_6661);
or U7345 (N_7345,N_6342,N_6670);
nand U7346 (N_7346,N_6595,N_6848);
xnor U7347 (N_7347,N_6349,N_6709);
and U7348 (N_7348,N_6266,N_6480);
nor U7349 (N_7349,N_6616,N_6710);
nor U7350 (N_7350,N_6450,N_6545);
xor U7351 (N_7351,N_6591,N_6674);
xnor U7352 (N_7352,N_6510,N_6636);
xor U7353 (N_7353,N_6256,N_6335);
and U7354 (N_7354,N_6360,N_6382);
nor U7355 (N_7355,N_6446,N_6315);
and U7356 (N_7356,N_6702,N_6692);
or U7357 (N_7357,N_6708,N_6475);
and U7358 (N_7358,N_6597,N_6620);
xnor U7359 (N_7359,N_6598,N_6341);
xor U7360 (N_7360,N_6536,N_6570);
nand U7361 (N_7361,N_6403,N_6311);
or U7362 (N_7362,N_6329,N_6862);
nor U7363 (N_7363,N_6496,N_6252);
nor U7364 (N_7364,N_6364,N_6873);
and U7365 (N_7365,N_6518,N_6335);
nand U7366 (N_7366,N_6685,N_6411);
nor U7367 (N_7367,N_6489,N_6599);
xnor U7368 (N_7368,N_6822,N_6345);
and U7369 (N_7369,N_6603,N_6838);
nand U7370 (N_7370,N_6590,N_6843);
and U7371 (N_7371,N_6705,N_6621);
xor U7372 (N_7372,N_6778,N_6417);
nand U7373 (N_7373,N_6497,N_6492);
nor U7374 (N_7374,N_6748,N_6855);
xnor U7375 (N_7375,N_6583,N_6600);
nand U7376 (N_7376,N_6529,N_6842);
and U7377 (N_7377,N_6643,N_6405);
and U7378 (N_7378,N_6723,N_6357);
xor U7379 (N_7379,N_6767,N_6717);
nor U7380 (N_7380,N_6273,N_6793);
or U7381 (N_7381,N_6542,N_6303);
nand U7382 (N_7382,N_6641,N_6409);
nand U7383 (N_7383,N_6568,N_6521);
or U7384 (N_7384,N_6793,N_6368);
nand U7385 (N_7385,N_6688,N_6739);
nand U7386 (N_7386,N_6685,N_6833);
and U7387 (N_7387,N_6748,N_6665);
and U7388 (N_7388,N_6742,N_6546);
nand U7389 (N_7389,N_6734,N_6356);
nor U7390 (N_7390,N_6308,N_6684);
or U7391 (N_7391,N_6594,N_6432);
nor U7392 (N_7392,N_6300,N_6420);
xnor U7393 (N_7393,N_6578,N_6749);
or U7394 (N_7394,N_6555,N_6265);
nor U7395 (N_7395,N_6348,N_6397);
xor U7396 (N_7396,N_6279,N_6866);
or U7397 (N_7397,N_6744,N_6771);
nand U7398 (N_7398,N_6779,N_6623);
or U7399 (N_7399,N_6718,N_6717);
nor U7400 (N_7400,N_6385,N_6603);
nand U7401 (N_7401,N_6854,N_6646);
and U7402 (N_7402,N_6429,N_6283);
and U7403 (N_7403,N_6607,N_6811);
nand U7404 (N_7404,N_6846,N_6817);
or U7405 (N_7405,N_6452,N_6320);
xor U7406 (N_7406,N_6269,N_6744);
nand U7407 (N_7407,N_6371,N_6384);
nor U7408 (N_7408,N_6581,N_6305);
nand U7409 (N_7409,N_6529,N_6740);
or U7410 (N_7410,N_6305,N_6313);
nand U7411 (N_7411,N_6569,N_6298);
nor U7412 (N_7412,N_6556,N_6441);
and U7413 (N_7413,N_6367,N_6652);
or U7414 (N_7414,N_6429,N_6607);
nand U7415 (N_7415,N_6502,N_6301);
nand U7416 (N_7416,N_6540,N_6863);
or U7417 (N_7417,N_6377,N_6315);
or U7418 (N_7418,N_6848,N_6413);
nor U7419 (N_7419,N_6364,N_6350);
nor U7420 (N_7420,N_6546,N_6550);
or U7421 (N_7421,N_6734,N_6638);
and U7422 (N_7422,N_6472,N_6363);
nor U7423 (N_7423,N_6651,N_6755);
nor U7424 (N_7424,N_6822,N_6477);
and U7425 (N_7425,N_6770,N_6804);
nand U7426 (N_7426,N_6653,N_6432);
nor U7427 (N_7427,N_6843,N_6871);
nor U7428 (N_7428,N_6633,N_6598);
or U7429 (N_7429,N_6793,N_6339);
xnor U7430 (N_7430,N_6356,N_6485);
nand U7431 (N_7431,N_6407,N_6607);
nor U7432 (N_7432,N_6623,N_6799);
nand U7433 (N_7433,N_6524,N_6389);
xnor U7434 (N_7434,N_6500,N_6765);
nor U7435 (N_7435,N_6634,N_6724);
nor U7436 (N_7436,N_6689,N_6525);
xor U7437 (N_7437,N_6488,N_6448);
and U7438 (N_7438,N_6381,N_6265);
nor U7439 (N_7439,N_6800,N_6329);
nor U7440 (N_7440,N_6673,N_6753);
nor U7441 (N_7441,N_6459,N_6741);
nand U7442 (N_7442,N_6760,N_6775);
xor U7443 (N_7443,N_6859,N_6538);
nor U7444 (N_7444,N_6766,N_6318);
nor U7445 (N_7445,N_6278,N_6828);
or U7446 (N_7446,N_6402,N_6610);
nor U7447 (N_7447,N_6759,N_6650);
nand U7448 (N_7448,N_6851,N_6309);
xnor U7449 (N_7449,N_6375,N_6394);
xor U7450 (N_7450,N_6865,N_6804);
nor U7451 (N_7451,N_6577,N_6560);
nor U7452 (N_7452,N_6643,N_6568);
xnor U7453 (N_7453,N_6683,N_6606);
and U7454 (N_7454,N_6413,N_6443);
xnor U7455 (N_7455,N_6335,N_6453);
nand U7456 (N_7456,N_6415,N_6676);
xnor U7457 (N_7457,N_6576,N_6482);
or U7458 (N_7458,N_6589,N_6604);
or U7459 (N_7459,N_6406,N_6482);
nor U7460 (N_7460,N_6559,N_6796);
or U7461 (N_7461,N_6507,N_6593);
xor U7462 (N_7462,N_6731,N_6605);
xor U7463 (N_7463,N_6504,N_6694);
or U7464 (N_7464,N_6809,N_6616);
or U7465 (N_7465,N_6870,N_6436);
xor U7466 (N_7466,N_6615,N_6500);
xnor U7467 (N_7467,N_6481,N_6370);
or U7468 (N_7468,N_6807,N_6452);
and U7469 (N_7469,N_6404,N_6439);
nor U7470 (N_7470,N_6616,N_6546);
and U7471 (N_7471,N_6474,N_6824);
nand U7472 (N_7472,N_6466,N_6325);
nor U7473 (N_7473,N_6725,N_6540);
nor U7474 (N_7474,N_6520,N_6666);
nor U7475 (N_7475,N_6744,N_6289);
xor U7476 (N_7476,N_6774,N_6555);
nor U7477 (N_7477,N_6465,N_6538);
nor U7478 (N_7478,N_6822,N_6259);
xor U7479 (N_7479,N_6767,N_6703);
and U7480 (N_7480,N_6516,N_6570);
xnor U7481 (N_7481,N_6618,N_6739);
and U7482 (N_7482,N_6828,N_6463);
or U7483 (N_7483,N_6294,N_6582);
or U7484 (N_7484,N_6434,N_6556);
nor U7485 (N_7485,N_6602,N_6811);
and U7486 (N_7486,N_6315,N_6364);
xor U7487 (N_7487,N_6418,N_6564);
or U7488 (N_7488,N_6495,N_6580);
xnor U7489 (N_7489,N_6512,N_6640);
or U7490 (N_7490,N_6762,N_6756);
nand U7491 (N_7491,N_6323,N_6630);
and U7492 (N_7492,N_6855,N_6417);
xnor U7493 (N_7493,N_6668,N_6599);
or U7494 (N_7494,N_6612,N_6697);
and U7495 (N_7495,N_6736,N_6407);
or U7496 (N_7496,N_6675,N_6272);
or U7497 (N_7497,N_6541,N_6363);
nor U7498 (N_7498,N_6308,N_6543);
or U7499 (N_7499,N_6362,N_6714);
or U7500 (N_7500,N_7397,N_6878);
nand U7501 (N_7501,N_7461,N_7050);
or U7502 (N_7502,N_7352,N_6927);
nor U7503 (N_7503,N_7118,N_7300);
and U7504 (N_7504,N_7140,N_7180);
xor U7505 (N_7505,N_7464,N_7177);
or U7506 (N_7506,N_6966,N_7164);
xnor U7507 (N_7507,N_7216,N_7381);
nand U7508 (N_7508,N_7110,N_7452);
and U7509 (N_7509,N_7175,N_6922);
and U7510 (N_7510,N_7139,N_7292);
and U7511 (N_7511,N_7046,N_7290);
nand U7512 (N_7512,N_7478,N_7296);
or U7513 (N_7513,N_7102,N_7451);
xor U7514 (N_7514,N_6923,N_7053);
nor U7515 (N_7515,N_6928,N_7198);
or U7516 (N_7516,N_6982,N_7161);
and U7517 (N_7517,N_7299,N_7295);
or U7518 (N_7518,N_7042,N_7472);
and U7519 (N_7519,N_7242,N_7430);
nand U7520 (N_7520,N_6935,N_7458);
nand U7521 (N_7521,N_7293,N_7469);
nor U7522 (N_7522,N_7051,N_7455);
nor U7523 (N_7523,N_7272,N_7243);
nand U7524 (N_7524,N_6889,N_7260);
nor U7525 (N_7525,N_6937,N_7089);
xnor U7526 (N_7526,N_6919,N_7067);
or U7527 (N_7527,N_7069,N_7280);
or U7528 (N_7528,N_7447,N_7221);
nor U7529 (N_7529,N_7390,N_7207);
nand U7530 (N_7530,N_6904,N_7291);
xor U7531 (N_7531,N_7385,N_7277);
or U7532 (N_7532,N_6977,N_7211);
and U7533 (N_7533,N_6985,N_7453);
and U7534 (N_7534,N_6913,N_7318);
or U7535 (N_7535,N_6894,N_6951);
or U7536 (N_7536,N_7147,N_7012);
xor U7537 (N_7537,N_7262,N_7034);
xnor U7538 (N_7538,N_7479,N_7080);
nand U7539 (N_7539,N_7462,N_7073);
or U7540 (N_7540,N_6897,N_7206);
nor U7541 (N_7541,N_7439,N_7255);
or U7542 (N_7542,N_7244,N_7486);
nand U7543 (N_7543,N_7226,N_7239);
xnor U7544 (N_7544,N_7388,N_6995);
or U7545 (N_7545,N_6912,N_7403);
xnor U7546 (N_7546,N_6952,N_6997);
nor U7547 (N_7547,N_7412,N_7470);
or U7548 (N_7548,N_7218,N_7285);
and U7549 (N_7549,N_6883,N_7096);
xnor U7550 (N_7550,N_7040,N_7298);
xor U7551 (N_7551,N_7329,N_7025);
nor U7552 (N_7552,N_6989,N_6971);
or U7553 (N_7553,N_7105,N_7029);
nor U7554 (N_7554,N_6947,N_7032);
xnor U7555 (N_7555,N_7353,N_7444);
and U7556 (N_7556,N_7016,N_7440);
nor U7557 (N_7557,N_6980,N_6993);
or U7558 (N_7558,N_6938,N_6892);
nand U7559 (N_7559,N_7436,N_7488);
xor U7560 (N_7560,N_7045,N_7245);
xor U7561 (N_7561,N_6973,N_6968);
or U7562 (N_7562,N_7492,N_7074);
xor U7563 (N_7563,N_7271,N_7038);
nor U7564 (N_7564,N_7126,N_7010);
xnor U7565 (N_7565,N_7375,N_7117);
nand U7566 (N_7566,N_7011,N_7205);
nand U7567 (N_7567,N_7106,N_6903);
and U7568 (N_7568,N_7151,N_7182);
xor U7569 (N_7569,N_7176,N_7030);
and U7570 (N_7570,N_7049,N_6978);
or U7571 (N_7571,N_7362,N_7442);
nand U7572 (N_7572,N_7201,N_7020);
or U7573 (N_7573,N_7121,N_7495);
xnor U7574 (N_7574,N_6957,N_7340);
xnor U7575 (N_7575,N_7428,N_7099);
or U7576 (N_7576,N_7332,N_6899);
or U7577 (N_7577,N_7072,N_7189);
nor U7578 (N_7578,N_7411,N_7409);
xnor U7579 (N_7579,N_6884,N_7471);
nand U7580 (N_7580,N_7389,N_7487);
nor U7581 (N_7581,N_7359,N_7449);
and U7582 (N_7582,N_7484,N_7265);
xnor U7583 (N_7583,N_7423,N_7047);
and U7584 (N_7584,N_7071,N_7348);
nand U7585 (N_7585,N_7311,N_7114);
nand U7586 (N_7586,N_6953,N_7079);
nand U7587 (N_7587,N_7497,N_6921);
or U7588 (N_7588,N_7361,N_7426);
nor U7589 (N_7589,N_7355,N_7191);
xor U7590 (N_7590,N_7056,N_7212);
or U7591 (N_7591,N_7491,N_7467);
xnor U7592 (N_7592,N_7227,N_7456);
xnor U7593 (N_7593,N_7209,N_7082);
xnor U7594 (N_7594,N_7024,N_7392);
and U7595 (N_7595,N_7398,N_7119);
nand U7596 (N_7596,N_7217,N_7008);
xor U7597 (N_7597,N_6880,N_7163);
nor U7598 (N_7598,N_7234,N_7386);
nand U7599 (N_7599,N_7123,N_7199);
nor U7600 (N_7600,N_6891,N_7345);
and U7601 (N_7601,N_6940,N_7181);
or U7602 (N_7602,N_7434,N_7107);
xnor U7603 (N_7603,N_7120,N_7100);
nand U7604 (N_7604,N_7153,N_7269);
or U7605 (N_7605,N_7257,N_7223);
nor U7606 (N_7606,N_6955,N_6876);
nand U7607 (N_7607,N_7168,N_7135);
and U7608 (N_7608,N_7408,N_7322);
nand U7609 (N_7609,N_6907,N_7376);
or U7610 (N_7610,N_7429,N_6916);
or U7611 (N_7611,N_6905,N_7092);
nand U7612 (N_7612,N_7331,N_7202);
nor U7613 (N_7613,N_7334,N_7261);
and U7614 (N_7614,N_7077,N_7279);
nand U7615 (N_7615,N_7335,N_7017);
and U7616 (N_7616,N_6917,N_7367);
and U7617 (N_7617,N_6964,N_7377);
or U7618 (N_7618,N_7372,N_7185);
xor U7619 (N_7619,N_7437,N_7490);
xnor U7620 (N_7620,N_6895,N_7027);
nand U7621 (N_7621,N_6909,N_7220);
nor U7622 (N_7622,N_6885,N_7132);
xnor U7623 (N_7623,N_7324,N_6900);
nand U7624 (N_7624,N_7267,N_7039);
nor U7625 (N_7625,N_7339,N_7315);
xnor U7626 (N_7626,N_7112,N_7263);
xnor U7627 (N_7627,N_7094,N_7405);
xnor U7628 (N_7628,N_7286,N_6879);
nor U7629 (N_7629,N_7004,N_6967);
nor U7630 (N_7630,N_7307,N_7278);
or U7631 (N_7631,N_7448,N_6945);
xnor U7632 (N_7632,N_7178,N_6887);
or U7633 (N_7633,N_7419,N_7197);
nor U7634 (N_7634,N_7005,N_7041);
xor U7635 (N_7635,N_7438,N_7143);
nand U7636 (N_7636,N_7460,N_7435);
and U7637 (N_7637,N_7404,N_7350);
and U7638 (N_7638,N_7413,N_7021);
nand U7639 (N_7639,N_7258,N_7000);
nand U7640 (N_7640,N_7309,N_7368);
xor U7641 (N_7641,N_7059,N_7036);
and U7642 (N_7642,N_7146,N_7317);
nand U7643 (N_7643,N_6877,N_7288);
xor U7644 (N_7644,N_7129,N_7433);
nand U7645 (N_7645,N_7224,N_7457);
nor U7646 (N_7646,N_7219,N_7327);
xor U7647 (N_7647,N_7459,N_7159);
nor U7648 (N_7648,N_6936,N_7276);
nor U7649 (N_7649,N_7160,N_7483);
and U7650 (N_7650,N_7001,N_7358);
and U7651 (N_7651,N_7144,N_7065);
xor U7652 (N_7652,N_7194,N_7225);
nor U7653 (N_7653,N_7009,N_7018);
nor U7654 (N_7654,N_7060,N_7137);
or U7655 (N_7655,N_6932,N_7169);
nor U7656 (N_7656,N_7289,N_7130);
nor U7657 (N_7657,N_7095,N_6988);
nor U7658 (N_7658,N_7445,N_7063);
nor U7659 (N_7659,N_7078,N_7314);
nand U7660 (N_7660,N_7252,N_7357);
or U7661 (N_7661,N_7195,N_7058);
and U7662 (N_7662,N_7190,N_7473);
and U7663 (N_7663,N_7128,N_7075);
or U7664 (N_7664,N_6898,N_7402);
or U7665 (N_7665,N_7333,N_7142);
xnor U7666 (N_7666,N_6976,N_6911);
nand U7667 (N_7667,N_7346,N_7363);
xnor U7668 (N_7668,N_7167,N_7305);
or U7669 (N_7669,N_7351,N_7310);
or U7670 (N_7670,N_7133,N_6970);
xnor U7671 (N_7671,N_7006,N_7066);
xor U7672 (N_7672,N_7418,N_6915);
or U7673 (N_7673,N_7157,N_7399);
and U7674 (N_7674,N_7134,N_7281);
or U7675 (N_7675,N_7476,N_7313);
or U7676 (N_7676,N_6974,N_7215);
or U7677 (N_7677,N_6983,N_6875);
and U7678 (N_7678,N_6996,N_7248);
nor U7679 (N_7679,N_7347,N_7237);
and U7680 (N_7680,N_7330,N_7382);
nor U7681 (N_7681,N_6943,N_7124);
xor U7682 (N_7682,N_7417,N_6882);
and U7683 (N_7683,N_6950,N_7481);
xnor U7684 (N_7684,N_7303,N_6925);
and U7685 (N_7685,N_7055,N_6975);
and U7686 (N_7686,N_7373,N_7301);
or U7687 (N_7687,N_7356,N_7253);
or U7688 (N_7688,N_7454,N_6908);
nand U7689 (N_7689,N_7098,N_7468);
xor U7690 (N_7690,N_7282,N_7186);
and U7691 (N_7691,N_7183,N_7304);
nor U7692 (N_7692,N_7249,N_7431);
and U7693 (N_7693,N_7489,N_7364);
nor U7694 (N_7694,N_6963,N_7165);
and U7695 (N_7695,N_6961,N_6902);
or U7696 (N_7696,N_7443,N_7229);
nor U7697 (N_7697,N_6890,N_7002);
xnor U7698 (N_7698,N_7023,N_7113);
nor U7699 (N_7699,N_7236,N_7238);
or U7700 (N_7700,N_7208,N_7294);
or U7701 (N_7701,N_7328,N_6965);
xor U7702 (N_7702,N_7235,N_7427);
nand U7703 (N_7703,N_6956,N_6999);
or U7704 (N_7704,N_7415,N_6949);
nor U7705 (N_7705,N_7284,N_6939);
or U7706 (N_7706,N_7316,N_7370);
nor U7707 (N_7707,N_7148,N_7342);
and U7708 (N_7708,N_7374,N_7193);
xnor U7709 (N_7709,N_7270,N_7410);
nor U7710 (N_7710,N_6954,N_6942);
xor U7711 (N_7711,N_6933,N_7028);
xor U7712 (N_7712,N_7097,N_7111);
nor U7713 (N_7713,N_7171,N_7275);
xor U7714 (N_7714,N_7407,N_6930);
or U7715 (N_7715,N_6929,N_7420);
nor U7716 (N_7716,N_6924,N_7086);
nand U7717 (N_7717,N_7064,N_7104);
nand U7718 (N_7718,N_7084,N_7406);
and U7719 (N_7719,N_7158,N_7391);
xor U7720 (N_7720,N_7325,N_6972);
and U7721 (N_7721,N_7421,N_7338);
nor U7722 (N_7722,N_7154,N_7187);
nor U7723 (N_7723,N_6914,N_7393);
or U7724 (N_7724,N_7319,N_7088);
or U7725 (N_7725,N_7365,N_6958);
and U7726 (N_7726,N_7425,N_7228);
nor U7727 (N_7727,N_7192,N_7349);
or U7728 (N_7728,N_6986,N_7015);
nand U7729 (N_7729,N_6948,N_7326);
and U7730 (N_7730,N_7337,N_7203);
nand U7731 (N_7731,N_6992,N_7463);
xor U7732 (N_7732,N_7394,N_7152);
nand U7733 (N_7733,N_7274,N_7173);
and U7734 (N_7734,N_7122,N_6941);
nor U7735 (N_7735,N_7019,N_7155);
xnor U7736 (N_7736,N_7268,N_7477);
nand U7737 (N_7737,N_7465,N_7170);
xnor U7738 (N_7738,N_7083,N_7441);
and U7739 (N_7739,N_6888,N_7283);
or U7740 (N_7740,N_7379,N_7166);
or U7741 (N_7741,N_7214,N_7387);
xor U7742 (N_7742,N_7496,N_7312);
nor U7743 (N_7743,N_7131,N_6918);
nand U7744 (N_7744,N_7068,N_7156);
nand U7745 (N_7745,N_7336,N_7432);
and U7746 (N_7746,N_7240,N_7091);
nand U7747 (N_7747,N_6991,N_7400);
and U7748 (N_7748,N_7213,N_7343);
nor U7749 (N_7749,N_7022,N_7087);
nand U7750 (N_7750,N_7250,N_6960);
nor U7751 (N_7751,N_7174,N_7341);
xnor U7752 (N_7752,N_6998,N_7360);
or U7753 (N_7753,N_7210,N_6962);
or U7754 (N_7754,N_7127,N_7035);
and U7755 (N_7755,N_7052,N_6994);
xor U7756 (N_7756,N_7101,N_7043);
nor U7757 (N_7757,N_7116,N_6944);
nand U7758 (N_7758,N_7085,N_7383);
and U7759 (N_7759,N_7204,N_6886);
xor U7760 (N_7760,N_7366,N_7371);
nand U7761 (N_7761,N_7344,N_7378);
nand U7762 (N_7762,N_7200,N_7273);
nor U7763 (N_7763,N_7048,N_7093);
nand U7764 (N_7764,N_7306,N_7061);
nand U7765 (N_7765,N_7401,N_7145);
nor U7766 (N_7766,N_7482,N_7499);
or U7767 (N_7767,N_7416,N_7081);
and U7768 (N_7768,N_7070,N_6893);
nand U7769 (N_7769,N_7172,N_6934);
or U7770 (N_7770,N_7115,N_6920);
or U7771 (N_7771,N_7422,N_7031);
xnor U7772 (N_7772,N_6969,N_7384);
xor U7773 (N_7773,N_7125,N_7090);
or U7774 (N_7774,N_7450,N_6981);
xnor U7775 (N_7775,N_6926,N_7062);
xnor U7776 (N_7776,N_7013,N_7466);
or U7777 (N_7777,N_7054,N_7474);
nor U7778 (N_7778,N_7138,N_7485);
xor U7779 (N_7779,N_7026,N_7354);
and U7780 (N_7780,N_6931,N_7424);
nand U7781 (N_7781,N_6990,N_7149);
or U7782 (N_7782,N_7323,N_6906);
xor U7783 (N_7783,N_6959,N_6946);
and U7784 (N_7784,N_7480,N_7179);
nor U7785 (N_7785,N_7446,N_6901);
or U7786 (N_7786,N_7308,N_7033);
and U7787 (N_7787,N_7014,N_7247);
nor U7788 (N_7788,N_7057,N_7232);
nand U7789 (N_7789,N_7184,N_7241);
xnor U7790 (N_7790,N_7254,N_6896);
and U7791 (N_7791,N_7494,N_7141);
or U7792 (N_7792,N_7037,N_7297);
and U7793 (N_7793,N_7108,N_7231);
or U7794 (N_7794,N_7256,N_7320);
or U7795 (N_7795,N_7076,N_6979);
nor U7796 (N_7796,N_7380,N_7414);
nand U7797 (N_7797,N_7287,N_7498);
or U7798 (N_7798,N_7264,N_6987);
nor U7799 (N_7799,N_7321,N_7369);
xnor U7800 (N_7800,N_6881,N_6984);
or U7801 (N_7801,N_7230,N_7044);
xnor U7802 (N_7802,N_7302,N_7103);
nand U7803 (N_7803,N_7222,N_7246);
xnor U7804 (N_7804,N_6910,N_7396);
or U7805 (N_7805,N_7493,N_7395);
xor U7806 (N_7806,N_7259,N_7475);
nand U7807 (N_7807,N_7266,N_7003);
nand U7808 (N_7808,N_7136,N_7162);
nor U7809 (N_7809,N_7251,N_7150);
nor U7810 (N_7810,N_7188,N_7007);
and U7811 (N_7811,N_7109,N_7233);
nor U7812 (N_7812,N_7196,N_7004);
and U7813 (N_7813,N_7242,N_6980);
and U7814 (N_7814,N_7420,N_6965);
and U7815 (N_7815,N_7198,N_7488);
or U7816 (N_7816,N_6923,N_7378);
or U7817 (N_7817,N_7246,N_7044);
nand U7818 (N_7818,N_6889,N_7487);
nand U7819 (N_7819,N_7088,N_7437);
xor U7820 (N_7820,N_6974,N_7163);
nand U7821 (N_7821,N_7243,N_7217);
xor U7822 (N_7822,N_7063,N_7296);
and U7823 (N_7823,N_7413,N_7314);
or U7824 (N_7824,N_7235,N_7234);
xnor U7825 (N_7825,N_7225,N_7110);
and U7826 (N_7826,N_7486,N_7462);
xnor U7827 (N_7827,N_7000,N_7405);
or U7828 (N_7828,N_7355,N_7086);
xnor U7829 (N_7829,N_7304,N_7360);
or U7830 (N_7830,N_7070,N_7285);
and U7831 (N_7831,N_7362,N_7203);
nor U7832 (N_7832,N_7246,N_6886);
or U7833 (N_7833,N_6989,N_6996);
xor U7834 (N_7834,N_7413,N_7466);
xnor U7835 (N_7835,N_6903,N_7181);
xor U7836 (N_7836,N_7161,N_7345);
nor U7837 (N_7837,N_7242,N_7125);
nor U7838 (N_7838,N_7469,N_7389);
and U7839 (N_7839,N_6960,N_7469);
nor U7840 (N_7840,N_6948,N_7136);
nand U7841 (N_7841,N_7007,N_7478);
nor U7842 (N_7842,N_6926,N_6948);
nand U7843 (N_7843,N_6925,N_7384);
xor U7844 (N_7844,N_6952,N_7497);
or U7845 (N_7845,N_7407,N_7309);
or U7846 (N_7846,N_7303,N_7410);
or U7847 (N_7847,N_7117,N_7396);
or U7848 (N_7848,N_7312,N_6991);
and U7849 (N_7849,N_6963,N_6876);
xnor U7850 (N_7850,N_7450,N_7172);
nor U7851 (N_7851,N_6910,N_7447);
nor U7852 (N_7852,N_7295,N_7228);
nand U7853 (N_7853,N_7406,N_7071);
and U7854 (N_7854,N_7236,N_7486);
nand U7855 (N_7855,N_7140,N_6986);
and U7856 (N_7856,N_7122,N_6972);
nor U7857 (N_7857,N_7328,N_7128);
nand U7858 (N_7858,N_7035,N_7378);
and U7859 (N_7859,N_7054,N_7299);
nand U7860 (N_7860,N_6935,N_7088);
or U7861 (N_7861,N_7092,N_7428);
nand U7862 (N_7862,N_7409,N_6924);
nand U7863 (N_7863,N_7162,N_7306);
nor U7864 (N_7864,N_7295,N_7023);
or U7865 (N_7865,N_7175,N_7464);
or U7866 (N_7866,N_7237,N_7342);
xor U7867 (N_7867,N_7071,N_7380);
xnor U7868 (N_7868,N_6943,N_7461);
xor U7869 (N_7869,N_7024,N_7226);
xnor U7870 (N_7870,N_6993,N_7272);
nor U7871 (N_7871,N_7484,N_7404);
xnor U7872 (N_7872,N_7077,N_6915);
nor U7873 (N_7873,N_7458,N_6889);
xnor U7874 (N_7874,N_7183,N_7037);
nor U7875 (N_7875,N_6937,N_7447);
nor U7876 (N_7876,N_7314,N_6995);
and U7877 (N_7877,N_7052,N_6928);
xor U7878 (N_7878,N_7146,N_7434);
xor U7879 (N_7879,N_7101,N_6974);
nand U7880 (N_7880,N_7372,N_7311);
nor U7881 (N_7881,N_7483,N_7249);
or U7882 (N_7882,N_6958,N_7356);
nand U7883 (N_7883,N_7218,N_7062);
xor U7884 (N_7884,N_7084,N_7030);
nand U7885 (N_7885,N_7112,N_7029);
nor U7886 (N_7886,N_7309,N_7363);
or U7887 (N_7887,N_7374,N_7150);
xor U7888 (N_7888,N_7231,N_7225);
and U7889 (N_7889,N_7142,N_7320);
or U7890 (N_7890,N_7129,N_7365);
nor U7891 (N_7891,N_6880,N_7391);
or U7892 (N_7892,N_7216,N_7008);
or U7893 (N_7893,N_6998,N_7248);
nor U7894 (N_7894,N_7024,N_7061);
and U7895 (N_7895,N_7484,N_7126);
or U7896 (N_7896,N_7259,N_7417);
nor U7897 (N_7897,N_6914,N_7234);
xnor U7898 (N_7898,N_7229,N_7368);
and U7899 (N_7899,N_7424,N_7167);
or U7900 (N_7900,N_7318,N_7232);
or U7901 (N_7901,N_7453,N_7344);
nor U7902 (N_7902,N_7050,N_7231);
and U7903 (N_7903,N_6881,N_6920);
xnor U7904 (N_7904,N_7145,N_7354);
nor U7905 (N_7905,N_7186,N_7012);
nand U7906 (N_7906,N_6974,N_7482);
nand U7907 (N_7907,N_7321,N_7151);
or U7908 (N_7908,N_7410,N_7220);
nor U7909 (N_7909,N_7101,N_7221);
nor U7910 (N_7910,N_7155,N_7016);
or U7911 (N_7911,N_7110,N_7140);
and U7912 (N_7912,N_7299,N_6980);
xnor U7913 (N_7913,N_7097,N_7297);
nor U7914 (N_7914,N_7415,N_7385);
and U7915 (N_7915,N_7135,N_6950);
nor U7916 (N_7916,N_7214,N_7498);
nand U7917 (N_7917,N_6904,N_6958);
and U7918 (N_7918,N_7000,N_7453);
xor U7919 (N_7919,N_6933,N_7343);
and U7920 (N_7920,N_7309,N_6914);
or U7921 (N_7921,N_6928,N_6985);
nor U7922 (N_7922,N_6882,N_7103);
nor U7923 (N_7923,N_7175,N_7120);
nand U7924 (N_7924,N_7396,N_7113);
nand U7925 (N_7925,N_7083,N_6910);
or U7926 (N_7926,N_7002,N_6945);
xnor U7927 (N_7927,N_6966,N_6992);
or U7928 (N_7928,N_7120,N_7256);
and U7929 (N_7929,N_7127,N_7188);
nand U7930 (N_7930,N_7082,N_7345);
nor U7931 (N_7931,N_6983,N_6896);
or U7932 (N_7932,N_7038,N_7276);
nand U7933 (N_7933,N_7070,N_7240);
and U7934 (N_7934,N_7213,N_7307);
nand U7935 (N_7935,N_7364,N_7260);
xnor U7936 (N_7936,N_6948,N_7199);
or U7937 (N_7937,N_7237,N_7010);
and U7938 (N_7938,N_6889,N_7035);
or U7939 (N_7939,N_7075,N_6974);
and U7940 (N_7940,N_7180,N_7014);
nand U7941 (N_7941,N_7166,N_7465);
xnor U7942 (N_7942,N_7488,N_7196);
nor U7943 (N_7943,N_7362,N_7249);
and U7944 (N_7944,N_7203,N_7360);
or U7945 (N_7945,N_7093,N_7394);
and U7946 (N_7946,N_7407,N_6896);
nor U7947 (N_7947,N_6960,N_7098);
and U7948 (N_7948,N_7188,N_7060);
xor U7949 (N_7949,N_7142,N_7294);
or U7950 (N_7950,N_7281,N_6920);
nand U7951 (N_7951,N_7450,N_7447);
nor U7952 (N_7952,N_7284,N_6917);
and U7953 (N_7953,N_7293,N_7403);
nand U7954 (N_7954,N_6916,N_7469);
nand U7955 (N_7955,N_7068,N_6880);
xor U7956 (N_7956,N_7082,N_7177);
nor U7957 (N_7957,N_7464,N_7081);
xnor U7958 (N_7958,N_6917,N_7152);
or U7959 (N_7959,N_7329,N_6892);
xor U7960 (N_7960,N_7222,N_7334);
and U7961 (N_7961,N_7275,N_7486);
xnor U7962 (N_7962,N_6961,N_7380);
and U7963 (N_7963,N_7356,N_7378);
and U7964 (N_7964,N_7335,N_6884);
and U7965 (N_7965,N_6956,N_7468);
nor U7966 (N_7966,N_7454,N_7409);
or U7967 (N_7967,N_6997,N_7482);
nand U7968 (N_7968,N_7187,N_7400);
nor U7969 (N_7969,N_7311,N_7083);
and U7970 (N_7970,N_7391,N_6882);
and U7971 (N_7971,N_7182,N_6995);
and U7972 (N_7972,N_7277,N_7214);
nand U7973 (N_7973,N_7420,N_7148);
or U7974 (N_7974,N_6946,N_6986);
nor U7975 (N_7975,N_7350,N_7095);
and U7976 (N_7976,N_7070,N_7182);
and U7977 (N_7977,N_7046,N_7348);
and U7978 (N_7978,N_7344,N_7086);
xor U7979 (N_7979,N_7051,N_7023);
nand U7980 (N_7980,N_7431,N_6968);
xor U7981 (N_7981,N_7183,N_7296);
nor U7982 (N_7982,N_7180,N_7023);
xnor U7983 (N_7983,N_7353,N_7155);
or U7984 (N_7984,N_7321,N_7317);
nand U7985 (N_7985,N_7274,N_7384);
and U7986 (N_7986,N_6910,N_7049);
and U7987 (N_7987,N_7397,N_7261);
and U7988 (N_7988,N_7377,N_6948);
or U7989 (N_7989,N_7399,N_6980);
nor U7990 (N_7990,N_6957,N_7426);
nand U7991 (N_7991,N_7344,N_7372);
xnor U7992 (N_7992,N_7010,N_6911);
nand U7993 (N_7993,N_7014,N_7346);
xnor U7994 (N_7994,N_7017,N_7291);
and U7995 (N_7995,N_7191,N_7086);
and U7996 (N_7996,N_7107,N_7242);
nor U7997 (N_7997,N_6998,N_7487);
nor U7998 (N_7998,N_7116,N_6969);
and U7999 (N_7999,N_7130,N_7495);
xnor U8000 (N_8000,N_7263,N_7169);
nor U8001 (N_8001,N_7226,N_6942);
or U8002 (N_8002,N_7260,N_7257);
xnor U8003 (N_8003,N_7244,N_7214);
xnor U8004 (N_8004,N_6875,N_7251);
and U8005 (N_8005,N_7187,N_7438);
xnor U8006 (N_8006,N_7035,N_7185);
or U8007 (N_8007,N_7210,N_7183);
nand U8008 (N_8008,N_7072,N_7109);
nor U8009 (N_8009,N_7324,N_6937);
nand U8010 (N_8010,N_7416,N_6903);
nand U8011 (N_8011,N_7279,N_7327);
xor U8012 (N_8012,N_7082,N_7465);
xor U8013 (N_8013,N_7187,N_7291);
nor U8014 (N_8014,N_7340,N_7105);
xnor U8015 (N_8015,N_7360,N_6902);
nor U8016 (N_8016,N_7023,N_6949);
nor U8017 (N_8017,N_6938,N_7283);
nand U8018 (N_8018,N_7008,N_7267);
nand U8019 (N_8019,N_7254,N_6882);
and U8020 (N_8020,N_7070,N_6939);
nor U8021 (N_8021,N_7487,N_7363);
or U8022 (N_8022,N_7294,N_7089);
xor U8023 (N_8023,N_7435,N_7024);
xnor U8024 (N_8024,N_7051,N_7287);
nand U8025 (N_8025,N_7048,N_7252);
and U8026 (N_8026,N_6906,N_7245);
and U8027 (N_8027,N_7216,N_7016);
nand U8028 (N_8028,N_7259,N_7235);
or U8029 (N_8029,N_7010,N_6975);
xnor U8030 (N_8030,N_6996,N_7286);
and U8031 (N_8031,N_7061,N_7223);
xnor U8032 (N_8032,N_7108,N_7003);
nor U8033 (N_8033,N_7441,N_6915);
and U8034 (N_8034,N_7490,N_7390);
and U8035 (N_8035,N_7376,N_6943);
and U8036 (N_8036,N_7068,N_7093);
nand U8037 (N_8037,N_7366,N_7200);
nand U8038 (N_8038,N_7166,N_6924);
and U8039 (N_8039,N_7449,N_6958);
xor U8040 (N_8040,N_7470,N_7279);
and U8041 (N_8041,N_7138,N_7142);
or U8042 (N_8042,N_7001,N_6882);
nor U8043 (N_8043,N_7273,N_7020);
nand U8044 (N_8044,N_7209,N_7294);
or U8045 (N_8045,N_7354,N_7140);
and U8046 (N_8046,N_7162,N_7147);
or U8047 (N_8047,N_7172,N_7298);
or U8048 (N_8048,N_7038,N_7127);
nand U8049 (N_8049,N_7475,N_7126);
nand U8050 (N_8050,N_7470,N_7242);
nand U8051 (N_8051,N_7249,N_7481);
and U8052 (N_8052,N_7367,N_6995);
nor U8053 (N_8053,N_7266,N_7151);
nand U8054 (N_8054,N_7103,N_7123);
nand U8055 (N_8055,N_6890,N_7084);
nor U8056 (N_8056,N_7380,N_7348);
and U8057 (N_8057,N_7186,N_7137);
and U8058 (N_8058,N_7380,N_6938);
and U8059 (N_8059,N_7301,N_7278);
and U8060 (N_8060,N_7475,N_7406);
or U8061 (N_8061,N_7467,N_7320);
or U8062 (N_8062,N_7061,N_7382);
nor U8063 (N_8063,N_6963,N_6919);
or U8064 (N_8064,N_7229,N_7404);
and U8065 (N_8065,N_7058,N_7054);
xor U8066 (N_8066,N_7248,N_7069);
and U8067 (N_8067,N_7258,N_7162);
and U8068 (N_8068,N_7122,N_7309);
nand U8069 (N_8069,N_7268,N_7143);
or U8070 (N_8070,N_7211,N_7331);
nand U8071 (N_8071,N_7423,N_7254);
or U8072 (N_8072,N_7443,N_7101);
or U8073 (N_8073,N_7424,N_7061);
and U8074 (N_8074,N_7258,N_7350);
xor U8075 (N_8075,N_7008,N_7035);
nand U8076 (N_8076,N_7060,N_7484);
nor U8077 (N_8077,N_6878,N_7370);
xor U8078 (N_8078,N_7120,N_6911);
or U8079 (N_8079,N_7439,N_7427);
and U8080 (N_8080,N_7057,N_7197);
nor U8081 (N_8081,N_6967,N_7310);
or U8082 (N_8082,N_7007,N_7368);
nand U8083 (N_8083,N_7137,N_7083);
nor U8084 (N_8084,N_7344,N_6955);
or U8085 (N_8085,N_7133,N_7111);
nand U8086 (N_8086,N_7140,N_7446);
xnor U8087 (N_8087,N_7256,N_7193);
xnor U8088 (N_8088,N_7116,N_7473);
xor U8089 (N_8089,N_7058,N_7061);
and U8090 (N_8090,N_6959,N_7134);
nand U8091 (N_8091,N_7095,N_7125);
or U8092 (N_8092,N_7477,N_7061);
or U8093 (N_8093,N_7067,N_7169);
and U8094 (N_8094,N_7208,N_7282);
nor U8095 (N_8095,N_7243,N_7429);
xor U8096 (N_8096,N_6947,N_6907);
nor U8097 (N_8097,N_7000,N_6975);
or U8098 (N_8098,N_7149,N_7172);
nor U8099 (N_8099,N_7236,N_7027);
and U8100 (N_8100,N_7371,N_7347);
and U8101 (N_8101,N_6959,N_6978);
or U8102 (N_8102,N_7064,N_7499);
xnor U8103 (N_8103,N_7409,N_7150);
xor U8104 (N_8104,N_7326,N_7013);
xnor U8105 (N_8105,N_7195,N_6985);
nand U8106 (N_8106,N_7036,N_7026);
and U8107 (N_8107,N_6935,N_6901);
or U8108 (N_8108,N_7068,N_6877);
nor U8109 (N_8109,N_7362,N_6948);
xnor U8110 (N_8110,N_7360,N_7083);
xnor U8111 (N_8111,N_7069,N_7218);
and U8112 (N_8112,N_7499,N_7188);
or U8113 (N_8113,N_7495,N_7481);
nand U8114 (N_8114,N_6876,N_7387);
and U8115 (N_8115,N_7014,N_7118);
and U8116 (N_8116,N_7444,N_7251);
or U8117 (N_8117,N_7058,N_7196);
nor U8118 (N_8118,N_7016,N_7029);
xor U8119 (N_8119,N_6943,N_7362);
xor U8120 (N_8120,N_7456,N_7105);
xor U8121 (N_8121,N_7355,N_7165);
nor U8122 (N_8122,N_7304,N_6982);
or U8123 (N_8123,N_7182,N_7421);
nor U8124 (N_8124,N_6947,N_7252);
nor U8125 (N_8125,N_7649,N_7930);
and U8126 (N_8126,N_7650,N_7934);
and U8127 (N_8127,N_7865,N_7733);
or U8128 (N_8128,N_8029,N_7715);
nor U8129 (N_8129,N_7957,N_8096);
xor U8130 (N_8130,N_8008,N_7942);
or U8131 (N_8131,N_7707,N_7785);
and U8132 (N_8132,N_8067,N_7555);
and U8133 (N_8133,N_7594,N_7545);
xnor U8134 (N_8134,N_7864,N_7968);
or U8135 (N_8135,N_7516,N_7807);
and U8136 (N_8136,N_7795,N_8048);
nand U8137 (N_8137,N_8061,N_7967);
nor U8138 (N_8138,N_7791,N_7953);
and U8139 (N_8139,N_7861,N_7568);
and U8140 (N_8140,N_7991,N_7582);
and U8141 (N_8141,N_8099,N_7681);
nand U8142 (N_8142,N_8076,N_7872);
nor U8143 (N_8143,N_8068,N_7808);
or U8144 (N_8144,N_7614,N_7718);
nand U8145 (N_8145,N_7546,N_7743);
nand U8146 (N_8146,N_7829,N_7810);
nand U8147 (N_8147,N_7887,N_8051);
xor U8148 (N_8148,N_7759,N_8025);
xor U8149 (N_8149,N_8090,N_7731);
nand U8150 (N_8150,N_7600,N_7607);
or U8151 (N_8151,N_8038,N_7653);
or U8152 (N_8152,N_7907,N_7534);
nor U8153 (N_8153,N_7971,N_7925);
xor U8154 (N_8154,N_7560,N_7672);
or U8155 (N_8155,N_7659,N_7690);
or U8156 (N_8156,N_7993,N_7914);
and U8157 (N_8157,N_7622,N_7851);
or U8158 (N_8158,N_7879,N_8036);
nand U8159 (N_8159,N_8024,N_7855);
xnor U8160 (N_8160,N_7884,N_8082);
or U8161 (N_8161,N_7714,N_7984);
xor U8162 (N_8162,N_7557,N_7951);
xor U8163 (N_8163,N_7547,N_7794);
nand U8164 (N_8164,N_7933,N_7770);
nand U8165 (N_8165,N_7592,N_7799);
and U8166 (N_8166,N_7945,N_8101);
and U8167 (N_8167,N_7746,N_8077);
or U8168 (N_8168,N_7542,N_7937);
xor U8169 (N_8169,N_7742,N_7676);
nor U8170 (N_8170,N_7705,N_7540);
and U8171 (N_8171,N_8100,N_8124);
or U8172 (N_8172,N_7593,N_7577);
and U8173 (N_8173,N_7686,N_7543);
nand U8174 (N_8174,N_7633,N_7862);
xor U8175 (N_8175,N_7973,N_7848);
nand U8176 (N_8176,N_7623,N_8045);
or U8177 (N_8177,N_7868,N_7652);
or U8178 (N_8178,N_7943,N_7918);
or U8179 (N_8179,N_8047,N_7575);
xnor U8180 (N_8180,N_7580,N_7752);
nand U8181 (N_8181,N_7936,N_8005);
nand U8182 (N_8182,N_7767,N_7517);
nor U8183 (N_8183,N_8083,N_8054);
and U8184 (N_8184,N_7701,N_7806);
or U8185 (N_8185,N_7610,N_7667);
nand U8186 (N_8186,N_7663,N_7741);
or U8187 (N_8187,N_7768,N_7771);
or U8188 (N_8188,N_7627,N_7927);
and U8189 (N_8189,N_7751,N_8030);
nor U8190 (N_8190,N_7763,N_7589);
nor U8191 (N_8191,N_7734,N_7565);
xnor U8192 (N_8192,N_7717,N_7809);
xnor U8193 (N_8193,N_7689,N_7790);
or U8194 (N_8194,N_7842,N_7657);
nand U8195 (N_8195,N_8010,N_7959);
and U8196 (N_8196,N_7812,N_7845);
xnor U8197 (N_8197,N_8088,N_7617);
or U8198 (N_8198,N_7780,N_7856);
nand U8199 (N_8199,N_7896,N_7635);
nor U8200 (N_8200,N_7749,N_7738);
xnor U8201 (N_8201,N_7670,N_8015);
xor U8202 (N_8202,N_7588,N_7559);
nand U8203 (N_8203,N_8056,N_7551);
and U8204 (N_8204,N_8074,N_7917);
nand U8205 (N_8205,N_7928,N_7569);
and U8206 (N_8206,N_7818,N_7815);
nor U8207 (N_8207,N_7988,N_7518);
or U8208 (N_8208,N_8106,N_7624);
xnor U8209 (N_8209,N_7834,N_7677);
and U8210 (N_8210,N_7946,N_7924);
and U8211 (N_8211,N_8012,N_8001);
nor U8212 (N_8212,N_7688,N_7660);
or U8213 (N_8213,N_8057,N_7537);
and U8214 (N_8214,N_7802,N_7612);
nor U8215 (N_8215,N_7880,N_7827);
nand U8216 (N_8216,N_7507,N_7964);
or U8217 (N_8217,N_8037,N_8011);
nand U8218 (N_8218,N_8107,N_8066);
xor U8219 (N_8219,N_7905,N_7995);
nor U8220 (N_8220,N_7506,N_7538);
and U8221 (N_8221,N_7509,N_7773);
nand U8222 (N_8222,N_7858,N_7618);
nand U8223 (N_8223,N_7631,N_7950);
or U8224 (N_8224,N_7893,N_7695);
nand U8225 (N_8225,N_7755,N_7748);
xnor U8226 (N_8226,N_7990,N_7515);
xnor U8227 (N_8227,N_7669,N_7643);
and U8228 (N_8228,N_7826,N_8122);
or U8229 (N_8229,N_7713,N_7904);
xor U8230 (N_8230,N_8123,N_8042);
xor U8231 (N_8231,N_7940,N_7673);
nand U8232 (N_8232,N_7720,N_7836);
nor U8233 (N_8233,N_7760,N_7691);
nor U8234 (N_8234,N_7835,N_7919);
xor U8235 (N_8235,N_7938,N_8018);
xor U8236 (N_8236,N_7709,N_7792);
nand U8237 (N_8237,N_8043,N_7952);
nand U8238 (N_8238,N_7874,N_7970);
nor U8239 (N_8239,N_7522,N_7974);
or U8240 (N_8240,N_7753,N_7573);
nor U8241 (N_8241,N_7888,N_7541);
and U8242 (N_8242,N_7894,N_7825);
or U8243 (N_8243,N_8022,N_8095);
nor U8244 (N_8244,N_7897,N_7583);
xor U8245 (N_8245,N_7616,N_7831);
or U8246 (N_8246,N_7869,N_8112);
xor U8247 (N_8247,N_7889,N_7931);
and U8248 (N_8248,N_7615,N_7939);
or U8249 (N_8249,N_7566,N_7822);
nor U8250 (N_8250,N_8085,N_7661);
and U8251 (N_8251,N_7563,N_7723);
nand U8252 (N_8252,N_7619,N_7696);
and U8253 (N_8253,N_8027,N_7601);
or U8254 (N_8254,N_7776,N_8009);
xor U8255 (N_8255,N_8064,N_7781);
xor U8256 (N_8256,N_7620,N_8075);
and U8257 (N_8257,N_7986,N_8111);
and U8258 (N_8258,N_7671,N_7687);
or U8259 (N_8259,N_7700,N_8115);
and U8260 (N_8260,N_8071,N_7960);
nor U8261 (N_8261,N_7639,N_7598);
nand U8262 (N_8262,N_8117,N_8097);
xnor U8263 (N_8263,N_7722,N_7531);
nand U8264 (N_8264,N_7975,N_7944);
nand U8265 (N_8265,N_7866,N_8035);
nand U8266 (N_8266,N_7912,N_7564);
or U8267 (N_8267,N_7976,N_7504);
or U8268 (N_8268,N_7909,N_7916);
nand U8269 (N_8269,N_7996,N_7824);
nand U8270 (N_8270,N_7634,N_7920);
or U8271 (N_8271,N_7740,N_7535);
xnor U8272 (N_8272,N_7640,N_8032);
and U8273 (N_8273,N_7630,N_7621);
xor U8274 (N_8274,N_7730,N_8105);
nand U8275 (N_8275,N_8053,N_8006);
or U8276 (N_8276,N_8040,N_7777);
or U8277 (N_8277,N_8120,N_7766);
and U8278 (N_8278,N_8060,N_7756);
nor U8279 (N_8279,N_7502,N_7524);
or U8280 (N_8280,N_7638,N_7536);
or U8281 (N_8281,N_8084,N_7977);
and U8282 (N_8282,N_8019,N_7579);
or U8283 (N_8283,N_8121,N_7562);
xor U8284 (N_8284,N_7699,N_7883);
xnor U8285 (N_8285,N_8108,N_7523);
nor U8286 (N_8286,N_7632,N_8081);
or U8287 (N_8287,N_7911,N_7500);
and U8288 (N_8288,N_8014,N_7881);
xnor U8289 (N_8289,N_7932,N_7587);
and U8290 (N_8290,N_8003,N_7702);
or U8291 (N_8291,N_7739,N_7817);
nand U8292 (N_8292,N_7902,N_8087);
or U8293 (N_8293,N_7778,N_8055);
and U8294 (N_8294,N_7838,N_7764);
or U8295 (N_8295,N_8073,N_7526);
and U8296 (N_8296,N_7844,N_7982);
nand U8297 (N_8297,N_7591,N_7706);
nor U8298 (N_8298,N_8103,N_7665);
xnor U8299 (N_8299,N_8091,N_7839);
nand U8300 (N_8300,N_7508,N_8098);
or U8301 (N_8301,N_8118,N_7765);
and U8302 (N_8302,N_7729,N_7958);
or U8303 (N_8303,N_7684,N_7782);
nand U8304 (N_8304,N_7989,N_7901);
xor U8305 (N_8305,N_7774,N_7850);
or U8306 (N_8306,N_7606,N_7609);
or U8307 (N_8307,N_7948,N_7814);
xor U8308 (N_8308,N_7685,N_7513);
nor U8309 (N_8309,N_8046,N_7821);
and U8310 (N_8310,N_7693,N_7668);
and U8311 (N_8311,N_7886,N_7793);
nor U8312 (N_8312,N_8079,N_8044);
nor U8313 (N_8313,N_8033,N_7599);
nand U8314 (N_8314,N_7854,N_7962);
or U8315 (N_8315,N_7510,N_7692);
or U8316 (N_8316,N_7611,N_7570);
xor U8317 (N_8317,N_7520,N_8104);
and U8318 (N_8318,N_7801,N_7697);
or U8319 (N_8319,N_7750,N_7529);
nor U8320 (N_8320,N_7721,N_7726);
or U8321 (N_8321,N_7549,N_7954);
or U8322 (N_8322,N_7891,N_7737);
nand U8323 (N_8323,N_8065,N_8007);
or U8324 (N_8324,N_8016,N_7949);
or U8325 (N_8325,N_7788,N_7978);
nor U8326 (N_8326,N_7816,N_7747);
and U8327 (N_8327,N_7527,N_7603);
xor U8328 (N_8328,N_7556,N_7625);
or U8329 (N_8329,N_8023,N_7596);
nor U8330 (N_8330,N_8094,N_7629);
and U8331 (N_8331,N_7963,N_7533);
and U8332 (N_8332,N_7830,N_7608);
xnor U8333 (N_8333,N_8041,N_7727);
nand U8334 (N_8334,N_7985,N_7796);
and U8335 (N_8335,N_7525,N_7735);
nor U8336 (N_8336,N_8080,N_7820);
nand U8337 (N_8337,N_7980,N_7784);
and U8338 (N_8338,N_7955,N_7656);
and U8339 (N_8339,N_7719,N_7941);
or U8340 (N_8340,N_7605,N_7552);
and U8341 (N_8341,N_7833,N_7539);
nor U8342 (N_8342,N_7597,N_7595);
and U8343 (N_8343,N_7698,N_7885);
nor U8344 (N_8344,N_7772,N_7921);
nand U8345 (N_8345,N_7999,N_7553);
or U8346 (N_8346,N_7501,N_7875);
and U8347 (N_8347,N_8034,N_8116);
xnor U8348 (N_8348,N_7704,N_7994);
xor U8349 (N_8349,N_7849,N_7898);
and U8350 (N_8350,N_7890,N_7956);
nor U8351 (N_8351,N_7578,N_8109);
nor U8352 (N_8352,N_7910,N_8092);
nor U8353 (N_8353,N_7992,N_7680);
nor U8354 (N_8354,N_8052,N_7574);
nand U8355 (N_8355,N_8113,N_7514);
nand U8356 (N_8356,N_7644,N_7895);
nor U8357 (N_8357,N_7604,N_7892);
xnor U8358 (N_8358,N_7966,N_8013);
and U8359 (N_8359,N_7554,N_8086);
or U8360 (N_8360,N_8039,N_7658);
or U8361 (N_8361,N_7732,N_7882);
xor U8362 (N_8362,N_7997,N_7602);
or U8363 (N_8363,N_7636,N_7811);
or U8364 (N_8364,N_7915,N_7998);
and U8365 (N_8365,N_8021,N_7646);
nand U8366 (N_8366,N_7655,N_7528);
xor U8367 (N_8367,N_7754,N_8004);
nor U8368 (N_8368,N_7761,N_7900);
xor U8369 (N_8369,N_7648,N_7969);
nand U8370 (N_8370,N_7762,N_7789);
nor U8371 (N_8371,N_8089,N_8031);
nand U8372 (N_8372,N_7877,N_7736);
nand U8373 (N_8373,N_7972,N_7846);
xnor U8374 (N_8374,N_7783,N_7852);
nand U8375 (N_8375,N_7832,N_7876);
or U8376 (N_8376,N_7981,N_7935);
and U8377 (N_8377,N_8059,N_7803);
and U8378 (N_8378,N_7679,N_7870);
nor U8379 (N_8379,N_7585,N_7871);
or U8380 (N_8380,N_7853,N_7694);
and U8381 (N_8381,N_8119,N_7572);
and U8382 (N_8382,N_8017,N_7682);
or U8383 (N_8383,N_7922,N_7923);
or U8384 (N_8384,N_7511,N_7857);
xnor U8385 (N_8385,N_7666,N_7961);
nor U8386 (N_8386,N_7847,N_7654);
nor U8387 (N_8387,N_7683,N_7787);
and U8388 (N_8388,N_7503,N_7548);
nand U8389 (N_8389,N_7550,N_8028);
xnor U8390 (N_8390,N_8072,N_7613);
nor U8391 (N_8391,N_7819,N_7716);
and U8392 (N_8392,N_7947,N_7571);
nand U8393 (N_8393,N_7906,N_7926);
xnor U8394 (N_8394,N_8110,N_7544);
or U8395 (N_8395,N_7724,N_7899);
or U8396 (N_8396,N_7837,N_7711);
nand U8397 (N_8397,N_7532,N_7521);
xnor U8398 (N_8398,N_7823,N_8058);
nand U8399 (N_8399,N_7584,N_7867);
and U8400 (N_8400,N_7903,N_7841);
nor U8401 (N_8401,N_7813,N_7863);
or U8402 (N_8402,N_7745,N_7908);
nand U8403 (N_8403,N_7641,N_7561);
xnor U8404 (N_8404,N_7637,N_7769);
nand U8405 (N_8405,N_7505,N_7965);
or U8406 (N_8406,N_7987,N_7878);
nand U8407 (N_8407,N_7708,N_7710);
xnor U8408 (N_8408,N_7804,N_8114);
xor U8409 (N_8409,N_7628,N_7728);
or U8410 (N_8410,N_7800,N_7797);
xor U8411 (N_8411,N_7586,N_7651);
nor U8412 (N_8412,N_7662,N_7703);
and U8413 (N_8413,N_8002,N_8020);
nor U8414 (N_8414,N_7642,N_7558);
nand U8415 (N_8415,N_7725,N_8049);
xor U8416 (N_8416,N_7758,N_7929);
and U8417 (N_8417,N_7840,N_7645);
xnor U8418 (N_8418,N_8050,N_8069);
nand U8419 (N_8419,N_7805,N_8026);
and U8420 (N_8420,N_7712,N_7675);
nor U8421 (N_8421,N_8062,N_7664);
or U8422 (N_8422,N_7786,N_8070);
or U8423 (N_8423,N_7913,N_7860);
xnor U8424 (N_8424,N_7512,N_8000);
xnor U8425 (N_8425,N_7744,N_7757);
or U8426 (N_8426,N_7530,N_7576);
nand U8427 (N_8427,N_7843,N_8093);
and U8428 (N_8428,N_7678,N_7979);
and U8429 (N_8429,N_8102,N_7519);
nand U8430 (N_8430,N_7873,N_7590);
xor U8431 (N_8431,N_7674,N_7983);
and U8432 (N_8432,N_8078,N_7626);
nor U8433 (N_8433,N_7798,N_7859);
and U8434 (N_8434,N_7581,N_7567);
and U8435 (N_8435,N_7828,N_7779);
and U8436 (N_8436,N_8063,N_7775);
xnor U8437 (N_8437,N_7647,N_7942);
nor U8438 (N_8438,N_7517,N_7833);
and U8439 (N_8439,N_7604,N_7561);
nand U8440 (N_8440,N_7959,N_7701);
and U8441 (N_8441,N_7884,N_7576);
nor U8442 (N_8442,N_7968,N_8066);
or U8443 (N_8443,N_7737,N_7682);
or U8444 (N_8444,N_7779,N_7585);
or U8445 (N_8445,N_7801,N_7506);
xor U8446 (N_8446,N_7537,N_7844);
and U8447 (N_8447,N_7943,N_7764);
nor U8448 (N_8448,N_8066,N_7806);
or U8449 (N_8449,N_7891,N_7824);
or U8450 (N_8450,N_8102,N_7815);
or U8451 (N_8451,N_7740,N_8049);
or U8452 (N_8452,N_7894,N_8113);
xor U8453 (N_8453,N_7692,N_7879);
xnor U8454 (N_8454,N_7980,N_7758);
nand U8455 (N_8455,N_8008,N_7996);
or U8456 (N_8456,N_7936,N_7927);
and U8457 (N_8457,N_8059,N_8119);
xor U8458 (N_8458,N_7520,N_8068);
nor U8459 (N_8459,N_8102,N_7651);
and U8460 (N_8460,N_7578,N_7662);
xnor U8461 (N_8461,N_7568,N_7637);
nor U8462 (N_8462,N_8038,N_7990);
or U8463 (N_8463,N_7828,N_7756);
nand U8464 (N_8464,N_7861,N_8079);
xor U8465 (N_8465,N_7783,N_7737);
and U8466 (N_8466,N_7612,N_8033);
nor U8467 (N_8467,N_7983,N_7703);
nor U8468 (N_8468,N_7664,N_7739);
nor U8469 (N_8469,N_7763,N_7775);
nor U8470 (N_8470,N_7873,N_8103);
nand U8471 (N_8471,N_7741,N_7800);
or U8472 (N_8472,N_8035,N_7729);
nand U8473 (N_8473,N_8080,N_7823);
or U8474 (N_8474,N_7918,N_7906);
nor U8475 (N_8475,N_8027,N_8114);
xnor U8476 (N_8476,N_7955,N_7661);
nor U8477 (N_8477,N_8098,N_7886);
nand U8478 (N_8478,N_7573,N_7613);
xor U8479 (N_8479,N_8071,N_7809);
nand U8480 (N_8480,N_8119,N_7625);
and U8481 (N_8481,N_7582,N_7689);
nor U8482 (N_8482,N_7732,N_8005);
or U8483 (N_8483,N_7858,N_7764);
nand U8484 (N_8484,N_8001,N_7578);
nor U8485 (N_8485,N_7819,N_7995);
nor U8486 (N_8486,N_7942,N_8073);
or U8487 (N_8487,N_7647,N_8118);
or U8488 (N_8488,N_8009,N_8050);
and U8489 (N_8489,N_7637,N_7765);
nand U8490 (N_8490,N_7792,N_7755);
and U8491 (N_8491,N_8108,N_7586);
xnor U8492 (N_8492,N_7607,N_8002);
nand U8493 (N_8493,N_7758,N_8035);
and U8494 (N_8494,N_7973,N_7937);
or U8495 (N_8495,N_7525,N_7504);
xnor U8496 (N_8496,N_7697,N_7818);
and U8497 (N_8497,N_7742,N_7865);
or U8498 (N_8498,N_7542,N_7585);
nand U8499 (N_8499,N_7809,N_7575);
and U8500 (N_8500,N_7717,N_8081);
xnor U8501 (N_8501,N_7570,N_7888);
nand U8502 (N_8502,N_7525,N_7906);
xnor U8503 (N_8503,N_7768,N_7703);
nor U8504 (N_8504,N_7841,N_7682);
and U8505 (N_8505,N_7724,N_8086);
nand U8506 (N_8506,N_7781,N_7599);
or U8507 (N_8507,N_7849,N_7992);
or U8508 (N_8508,N_8040,N_7534);
and U8509 (N_8509,N_7965,N_7789);
and U8510 (N_8510,N_7737,N_7814);
nand U8511 (N_8511,N_7980,N_7636);
xnor U8512 (N_8512,N_7914,N_7861);
nor U8513 (N_8513,N_7642,N_7978);
or U8514 (N_8514,N_7563,N_7967);
or U8515 (N_8515,N_7616,N_8083);
and U8516 (N_8516,N_7622,N_7741);
or U8517 (N_8517,N_7516,N_7995);
nand U8518 (N_8518,N_7894,N_7554);
and U8519 (N_8519,N_7713,N_7799);
and U8520 (N_8520,N_7812,N_7853);
or U8521 (N_8521,N_7803,N_7850);
or U8522 (N_8522,N_7705,N_7890);
and U8523 (N_8523,N_7709,N_7679);
nor U8524 (N_8524,N_7930,N_8041);
or U8525 (N_8525,N_7524,N_7856);
and U8526 (N_8526,N_7589,N_7607);
and U8527 (N_8527,N_7814,N_7589);
or U8528 (N_8528,N_7963,N_8060);
xnor U8529 (N_8529,N_7719,N_8013);
nand U8530 (N_8530,N_7775,N_7587);
or U8531 (N_8531,N_7534,N_7815);
and U8532 (N_8532,N_7947,N_8019);
or U8533 (N_8533,N_7552,N_7729);
xnor U8534 (N_8534,N_7710,N_7535);
xor U8535 (N_8535,N_7876,N_7695);
nor U8536 (N_8536,N_7932,N_8012);
or U8537 (N_8537,N_7566,N_7855);
nor U8538 (N_8538,N_8066,N_7878);
or U8539 (N_8539,N_7665,N_7924);
nor U8540 (N_8540,N_7812,N_7882);
and U8541 (N_8541,N_7760,N_7753);
nand U8542 (N_8542,N_7773,N_7759);
xnor U8543 (N_8543,N_7506,N_7949);
nand U8544 (N_8544,N_7649,N_7860);
and U8545 (N_8545,N_7936,N_7548);
or U8546 (N_8546,N_7727,N_7895);
nand U8547 (N_8547,N_7554,N_7753);
xor U8548 (N_8548,N_7990,N_7620);
nor U8549 (N_8549,N_7695,N_7541);
xnor U8550 (N_8550,N_7850,N_7966);
nand U8551 (N_8551,N_7868,N_7894);
nor U8552 (N_8552,N_7950,N_7863);
nor U8553 (N_8553,N_7684,N_7850);
nor U8554 (N_8554,N_8006,N_7505);
nor U8555 (N_8555,N_7817,N_7873);
nand U8556 (N_8556,N_7603,N_8081);
nand U8557 (N_8557,N_7527,N_8033);
nor U8558 (N_8558,N_7701,N_7656);
and U8559 (N_8559,N_8085,N_7737);
nor U8560 (N_8560,N_7601,N_7546);
nor U8561 (N_8561,N_7676,N_7720);
nand U8562 (N_8562,N_7962,N_7945);
nand U8563 (N_8563,N_7707,N_7780);
or U8564 (N_8564,N_7708,N_7972);
nor U8565 (N_8565,N_7592,N_8083);
nand U8566 (N_8566,N_8025,N_7852);
nand U8567 (N_8567,N_8120,N_8097);
and U8568 (N_8568,N_8005,N_7867);
or U8569 (N_8569,N_7932,N_8114);
xnor U8570 (N_8570,N_7981,N_8059);
or U8571 (N_8571,N_8035,N_8050);
nor U8572 (N_8572,N_8114,N_7780);
nand U8573 (N_8573,N_7866,N_7523);
nor U8574 (N_8574,N_7642,N_7565);
nor U8575 (N_8575,N_7899,N_8095);
or U8576 (N_8576,N_7876,N_7808);
xor U8577 (N_8577,N_7573,N_7681);
xor U8578 (N_8578,N_7844,N_7641);
nor U8579 (N_8579,N_7608,N_7566);
nand U8580 (N_8580,N_7978,N_7750);
and U8581 (N_8581,N_7780,N_8082);
nor U8582 (N_8582,N_7729,N_8096);
xnor U8583 (N_8583,N_7961,N_7706);
xor U8584 (N_8584,N_7900,N_7636);
and U8585 (N_8585,N_7676,N_7882);
or U8586 (N_8586,N_7841,N_7623);
and U8587 (N_8587,N_8115,N_7629);
xnor U8588 (N_8588,N_7917,N_7980);
nor U8589 (N_8589,N_7501,N_7740);
nor U8590 (N_8590,N_7941,N_7922);
nand U8591 (N_8591,N_7634,N_7853);
nand U8592 (N_8592,N_7977,N_7522);
and U8593 (N_8593,N_7831,N_7929);
nand U8594 (N_8594,N_7510,N_7991);
nand U8595 (N_8595,N_7894,N_7725);
nor U8596 (N_8596,N_7665,N_7769);
nand U8597 (N_8597,N_7887,N_7768);
xor U8598 (N_8598,N_8044,N_7917);
or U8599 (N_8599,N_7592,N_7843);
and U8600 (N_8600,N_8039,N_7724);
xnor U8601 (N_8601,N_8026,N_7799);
or U8602 (N_8602,N_8020,N_7914);
nor U8603 (N_8603,N_7708,N_7807);
or U8604 (N_8604,N_7836,N_7654);
and U8605 (N_8605,N_7713,N_7855);
nand U8606 (N_8606,N_7808,N_8086);
xor U8607 (N_8607,N_7937,N_7986);
nand U8608 (N_8608,N_8049,N_7842);
and U8609 (N_8609,N_7862,N_7594);
nor U8610 (N_8610,N_8117,N_7609);
nor U8611 (N_8611,N_7688,N_7572);
and U8612 (N_8612,N_7661,N_7662);
xnor U8613 (N_8613,N_7603,N_7969);
nor U8614 (N_8614,N_7997,N_8077);
or U8615 (N_8615,N_7813,N_7513);
and U8616 (N_8616,N_7929,N_8055);
nand U8617 (N_8617,N_8082,N_7837);
nand U8618 (N_8618,N_7994,N_7717);
xnor U8619 (N_8619,N_7547,N_7574);
nor U8620 (N_8620,N_7726,N_7561);
or U8621 (N_8621,N_7843,N_8081);
and U8622 (N_8622,N_7999,N_7744);
and U8623 (N_8623,N_7634,N_7802);
nor U8624 (N_8624,N_7858,N_7694);
and U8625 (N_8625,N_7979,N_7958);
nor U8626 (N_8626,N_7849,N_7725);
and U8627 (N_8627,N_7696,N_8012);
and U8628 (N_8628,N_7630,N_7552);
xnor U8629 (N_8629,N_8012,N_7954);
or U8630 (N_8630,N_7935,N_8057);
xor U8631 (N_8631,N_7847,N_7613);
xnor U8632 (N_8632,N_8010,N_7878);
or U8633 (N_8633,N_7827,N_7759);
and U8634 (N_8634,N_8027,N_7582);
or U8635 (N_8635,N_7780,N_7923);
or U8636 (N_8636,N_7745,N_7511);
nor U8637 (N_8637,N_7738,N_8096);
and U8638 (N_8638,N_7714,N_8023);
nor U8639 (N_8639,N_7730,N_7665);
nand U8640 (N_8640,N_8048,N_7551);
xor U8641 (N_8641,N_7779,N_7528);
or U8642 (N_8642,N_7699,N_7959);
nand U8643 (N_8643,N_7620,N_7503);
nand U8644 (N_8644,N_7996,N_7584);
nand U8645 (N_8645,N_7697,N_7957);
and U8646 (N_8646,N_7731,N_7821);
xnor U8647 (N_8647,N_8043,N_7993);
nor U8648 (N_8648,N_7599,N_7842);
nand U8649 (N_8649,N_7792,N_7741);
xor U8650 (N_8650,N_7866,N_7964);
nand U8651 (N_8651,N_7782,N_8024);
xnor U8652 (N_8652,N_8110,N_8035);
nand U8653 (N_8653,N_8059,N_7658);
or U8654 (N_8654,N_7902,N_7859);
or U8655 (N_8655,N_8013,N_8093);
and U8656 (N_8656,N_7702,N_7782);
xnor U8657 (N_8657,N_7861,N_7701);
nor U8658 (N_8658,N_7670,N_8058);
and U8659 (N_8659,N_7553,N_8122);
nand U8660 (N_8660,N_7925,N_7730);
nor U8661 (N_8661,N_7564,N_7938);
nand U8662 (N_8662,N_7579,N_7784);
nor U8663 (N_8663,N_7729,N_7903);
nor U8664 (N_8664,N_7938,N_7760);
xnor U8665 (N_8665,N_7975,N_7865);
and U8666 (N_8666,N_7887,N_7799);
or U8667 (N_8667,N_7541,N_7849);
and U8668 (N_8668,N_7519,N_7640);
xor U8669 (N_8669,N_7983,N_7950);
nor U8670 (N_8670,N_7836,N_7663);
xor U8671 (N_8671,N_7558,N_8095);
xnor U8672 (N_8672,N_8039,N_8093);
and U8673 (N_8673,N_7662,N_7723);
or U8674 (N_8674,N_7536,N_7696);
nand U8675 (N_8675,N_7925,N_7737);
nand U8676 (N_8676,N_8066,N_7577);
xor U8677 (N_8677,N_7653,N_7981);
nand U8678 (N_8678,N_7667,N_7816);
or U8679 (N_8679,N_7667,N_8013);
nor U8680 (N_8680,N_7905,N_7767);
nor U8681 (N_8681,N_7917,N_7617);
and U8682 (N_8682,N_7526,N_7817);
and U8683 (N_8683,N_7747,N_7518);
xnor U8684 (N_8684,N_7511,N_7650);
nor U8685 (N_8685,N_7556,N_7742);
nand U8686 (N_8686,N_7663,N_7991);
or U8687 (N_8687,N_7867,N_7672);
xnor U8688 (N_8688,N_7652,N_7620);
and U8689 (N_8689,N_8099,N_8002);
nand U8690 (N_8690,N_8002,N_7721);
and U8691 (N_8691,N_7730,N_7648);
and U8692 (N_8692,N_7975,N_8020);
xor U8693 (N_8693,N_7526,N_7952);
or U8694 (N_8694,N_7536,N_7912);
nor U8695 (N_8695,N_7974,N_7606);
xnor U8696 (N_8696,N_7666,N_7691);
and U8697 (N_8697,N_7804,N_7629);
and U8698 (N_8698,N_7728,N_7937);
nor U8699 (N_8699,N_7916,N_8079);
xor U8700 (N_8700,N_7783,N_8074);
and U8701 (N_8701,N_7528,N_8060);
nand U8702 (N_8702,N_7662,N_8082);
and U8703 (N_8703,N_7932,N_7651);
nand U8704 (N_8704,N_7590,N_7596);
and U8705 (N_8705,N_7952,N_7570);
nor U8706 (N_8706,N_7788,N_7551);
and U8707 (N_8707,N_7789,N_7858);
nand U8708 (N_8708,N_7767,N_7685);
or U8709 (N_8709,N_7855,N_7937);
nand U8710 (N_8710,N_7737,N_7898);
xor U8711 (N_8711,N_7765,N_7805);
and U8712 (N_8712,N_7734,N_7697);
and U8713 (N_8713,N_7839,N_7989);
and U8714 (N_8714,N_7780,N_8014);
xor U8715 (N_8715,N_7606,N_7650);
and U8716 (N_8716,N_7631,N_7869);
nor U8717 (N_8717,N_8124,N_8019);
xnor U8718 (N_8718,N_7800,N_8036);
and U8719 (N_8719,N_7782,N_7852);
xnor U8720 (N_8720,N_7820,N_7607);
nand U8721 (N_8721,N_7973,N_7801);
and U8722 (N_8722,N_7530,N_7824);
nor U8723 (N_8723,N_7688,N_7739);
and U8724 (N_8724,N_8121,N_7994);
xor U8725 (N_8725,N_7557,N_7728);
or U8726 (N_8726,N_7820,N_7700);
nor U8727 (N_8727,N_7576,N_7970);
nand U8728 (N_8728,N_7885,N_8113);
nand U8729 (N_8729,N_7961,N_7619);
nor U8730 (N_8730,N_7924,N_7717);
nor U8731 (N_8731,N_8114,N_7885);
nor U8732 (N_8732,N_7915,N_7818);
nand U8733 (N_8733,N_8122,N_7911);
xnor U8734 (N_8734,N_7583,N_7562);
nor U8735 (N_8735,N_7517,N_8116);
xnor U8736 (N_8736,N_7852,N_8113);
nand U8737 (N_8737,N_8041,N_7994);
nor U8738 (N_8738,N_7947,N_7677);
and U8739 (N_8739,N_7940,N_7768);
nand U8740 (N_8740,N_7692,N_8038);
nand U8741 (N_8741,N_7977,N_7874);
and U8742 (N_8742,N_8023,N_7579);
and U8743 (N_8743,N_7661,N_8105);
nand U8744 (N_8744,N_7894,N_7974);
nand U8745 (N_8745,N_7553,N_8000);
nor U8746 (N_8746,N_7944,N_7598);
and U8747 (N_8747,N_7657,N_7648);
nor U8748 (N_8748,N_7958,N_7703);
nor U8749 (N_8749,N_7897,N_8001);
or U8750 (N_8750,N_8440,N_8574);
xnor U8751 (N_8751,N_8609,N_8424);
and U8752 (N_8752,N_8353,N_8737);
xor U8753 (N_8753,N_8473,N_8731);
and U8754 (N_8754,N_8418,N_8295);
xor U8755 (N_8755,N_8326,N_8144);
or U8756 (N_8756,N_8539,N_8673);
or U8757 (N_8757,N_8314,N_8416);
nand U8758 (N_8758,N_8245,N_8451);
and U8759 (N_8759,N_8478,N_8554);
or U8760 (N_8760,N_8330,N_8743);
nor U8761 (N_8761,N_8584,N_8710);
or U8762 (N_8762,N_8448,N_8193);
or U8763 (N_8763,N_8586,N_8238);
nand U8764 (N_8764,N_8361,N_8380);
xnor U8765 (N_8765,N_8542,N_8627);
and U8766 (N_8766,N_8517,N_8501);
xnor U8767 (N_8767,N_8626,N_8475);
nor U8768 (N_8768,N_8212,N_8508);
or U8769 (N_8769,N_8615,N_8339);
and U8770 (N_8770,N_8611,N_8393);
or U8771 (N_8771,N_8131,N_8715);
xor U8772 (N_8772,N_8665,N_8499);
and U8773 (N_8773,N_8494,N_8605);
nand U8774 (N_8774,N_8397,N_8218);
or U8775 (N_8775,N_8739,N_8137);
xnor U8776 (N_8776,N_8370,N_8298);
nand U8777 (N_8777,N_8301,N_8532);
xor U8778 (N_8778,N_8273,N_8650);
nand U8779 (N_8779,N_8625,N_8631);
xor U8780 (N_8780,N_8429,N_8745);
nor U8781 (N_8781,N_8324,N_8319);
nor U8782 (N_8782,N_8580,N_8576);
xor U8783 (N_8783,N_8682,N_8700);
xor U8784 (N_8784,N_8523,N_8307);
nor U8785 (N_8785,N_8192,N_8232);
nand U8786 (N_8786,N_8321,N_8642);
nand U8787 (N_8787,N_8602,N_8356);
nand U8788 (N_8788,N_8256,N_8342);
nor U8789 (N_8789,N_8322,N_8667);
and U8790 (N_8790,N_8589,N_8389);
xnor U8791 (N_8791,N_8606,N_8350);
and U8792 (N_8792,N_8262,N_8194);
and U8793 (N_8793,N_8660,N_8210);
nand U8794 (N_8794,N_8684,N_8138);
or U8795 (N_8795,N_8741,N_8555);
xnor U8796 (N_8796,N_8161,N_8513);
nand U8797 (N_8797,N_8723,N_8159);
or U8798 (N_8798,N_8509,N_8247);
and U8799 (N_8799,N_8169,N_8510);
xor U8800 (N_8800,N_8279,N_8672);
nand U8801 (N_8801,N_8711,N_8402);
and U8802 (N_8802,N_8414,N_8622);
xnor U8803 (N_8803,N_8549,N_8221);
xor U8804 (N_8804,N_8717,N_8514);
xor U8805 (N_8805,N_8306,N_8209);
nor U8806 (N_8806,N_8676,N_8135);
or U8807 (N_8807,N_8472,N_8726);
or U8808 (N_8808,N_8152,N_8263);
nor U8809 (N_8809,N_8354,N_8456);
and U8810 (N_8810,N_8671,N_8433);
and U8811 (N_8811,N_8381,N_8713);
or U8812 (N_8812,N_8577,N_8204);
and U8813 (N_8813,N_8228,N_8636);
nor U8814 (N_8814,N_8492,N_8734);
nor U8815 (N_8815,N_8647,N_8153);
and U8816 (N_8816,N_8729,N_8200);
nor U8817 (N_8817,N_8688,N_8657);
xnor U8818 (N_8818,N_8404,N_8173);
and U8819 (N_8819,N_8694,N_8638);
or U8820 (N_8820,N_8308,N_8629);
xnor U8821 (N_8821,N_8335,N_8543);
nand U8822 (N_8822,N_8243,N_8336);
nand U8823 (N_8823,N_8454,N_8744);
or U8824 (N_8824,N_8248,N_8362);
xnor U8825 (N_8825,N_8359,N_8242);
nor U8826 (N_8826,N_8220,N_8612);
xnor U8827 (N_8827,N_8390,N_8406);
nor U8828 (N_8828,N_8325,N_8365);
nand U8829 (N_8829,N_8477,N_8530);
or U8830 (N_8830,N_8255,N_8378);
nand U8831 (N_8831,N_8223,N_8702);
xor U8832 (N_8832,N_8323,N_8490);
or U8833 (N_8833,N_8136,N_8360);
or U8834 (N_8834,N_8208,N_8441);
xnor U8835 (N_8835,N_8703,N_8143);
nand U8836 (N_8836,N_8317,N_8377);
nand U8837 (N_8837,N_8338,N_8181);
or U8838 (N_8838,N_8716,N_8344);
or U8839 (N_8839,N_8593,N_8563);
nand U8840 (N_8840,N_8155,N_8480);
nand U8841 (N_8841,N_8373,N_8386);
and U8842 (N_8842,N_8655,N_8432);
nor U8843 (N_8843,N_8413,N_8640);
or U8844 (N_8844,N_8670,N_8746);
and U8845 (N_8845,N_8613,N_8195);
xor U8846 (N_8846,N_8229,N_8649);
xor U8847 (N_8847,N_8226,N_8468);
or U8848 (N_8848,N_8412,N_8348);
xnor U8849 (N_8849,N_8578,N_8595);
and U8850 (N_8850,N_8415,N_8654);
nor U8851 (N_8851,N_8411,N_8151);
and U8852 (N_8852,N_8610,N_8701);
xnor U8853 (N_8853,N_8343,N_8740);
nor U8854 (N_8854,N_8458,N_8240);
or U8855 (N_8855,N_8747,N_8296);
nand U8856 (N_8856,N_8363,N_8453);
nand U8857 (N_8857,N_8383,N_8132);
nand U8858 (N_8858,N_8529,N_8544);
and U8859 (N_8859,N_8461,N_8434);
xor U8860 (N_8860,N_8730,N_8460);
or U8861 (N_8861,N_8559,N_8297);
and U8862 (N_8862,N_8316,N_8225);
or U8863 (N_8863,N_8185,N_8355);
nand U8864 (N_8864,N_8674,N_8669);
nand U8865 (N_8865,N_8624,N_8430);
or U8866 (N_8866,N_8251,N_8698);
nor U8867 (N_8867,N_8175,N_8621);
nor U8868 (N_8868,N_8732,N_8180);
nand U8869 (N_8869,N_8214,N_8166);
nor U8870 (N_8870,N_8467,N_8568);
or U8871 (N_8871,N_8244,N_8565);
xnor U8872 (N_8872,N_8571,N_8372);
xor U8873 (N_8873,N_8252,N_8720);
nand U8874 (N_8874,N_8447,N_8455);
and U8875 (N_8875,N_8189,N_8696);
and U8876 (N_8876,N_8259,N_8556);
nand U8877 (N_8877,N_8130,N_8471);
or U8878 (N_8878,N_8553,N_8628);
xor U8879 (N_8879,N_8483,N_8619);
nand U8880 (N_8880,N_8444,N_8582);
xnor U8881 (N_8881,N_8401,N_8659);
nor U8882 (N_8882,N_8535,N_8643);
and U8883 (N_8883,N_8207,N_8391);
nor U8884 (N_8884,N_8721,N_8289);
nor U8885 (N_8885,N_8462,N_8283);
nor U8886 (N_8886,N_8522,N_8235);
and U8887 (N_8887,N_8352,N_8241);
xnor U8888 (N_8888,N_8215,N_8533);
nand U8889 (N_8889,N_8531,N_8234);
and U8890 (N_8890,N_8179,N_8504);
or U8891 (N_8891,N_8197,N_8253);
and U8892 (N_8892,N_8579,N_8691);
nor U8893 (N_8893,N_8641,N_8465);
and U8894 (N_8894,N_8186,N_8205);
xor U8895 (N_8895,N_8442,N_8603);
nand U8896 (N_8896,N_8709,N_8272);
or U8897 (N_8897,N_8267,N_8417);
and U8898 (N_8898,N_8176,N_8329);
nor U8899 (N_8899,N_8735,N_8512);
or U8900 (N_8900,N_8213,N_8566);
and U8901 (N_8901,N_8187,N_8435);
nor U8902 (N_8902,N_8598,N_8320);
nand U8903 (N_8903,N_8575,N_8632);
nand U8904 (N_8904,N_8463,N_8191);
nor U8905 (N_8905,N_8400,N_8217);
or U8906 (N_8906,N_8488,N_8171);
nand U8907 (N_8907,N_8617,N_8367);
nor U8908 (N_8908,N_8675,N_8570);
nand U8909 (N_8909,N_8170,N_8493);
xnor U8910 (N_8910,N_8183,N_8270);
and U8911 (N_8911,N_8608,N_8371);
and U8912 (N_8912,N_8592,N_8560);
xnor U8913 (N_8913,N_8311,N_8420);
and U8914 (N_8914,N_8485,N_8421);
nand U8915 (N_8915,N_8190,N_8573);
or U8916 (N_8916,N_8548,N_8382);
nor U8917 (N_8917,N_8409,N_8596);
nor U8918 (N_8918,N_8639,N_8351);
xnor U8919 (N_8919,N_8250,N_8257);
xnor U8920 (N_8920,N_8474,N_8695);
nand U8921 (N_8921,N_8552,N_8302);
or U8922 (N_8922,N_8260,N_8633);
nor U8923 (N_8923,N_8140,N_8630);
xor U8924 (N_8924,N_8310,N_8534);
nand U8925 (N_8925,N_8690,N_8237);
or U8926 (N_8926,N_8149,N_8516);
xor U8927 (N_8927,N_8206,N_8349);
nand U8928 (N_8928,N_8146,N_8422);
nand U8929 (N_8929,N_8203,N_8450);
nor U8930 (N_8930,N_8699,N_8287);
nand U8931 (N_8931,N_8452,N_8284);
or U8932 (N_8932,N_8182,N_8724);
or U8933 (N_8933,N_8249,N_8384);
or U8934 (N_8934,N_8196,N_8599);
and U8935 (N_8935,N_8133,N_8318);
or U8936 (N_8936,N_8469,N_8294);
nand U8937 (N_8937,N_8374,N_8268);
nand U8938 (N_8938,N_8585,N_8738);
or U8939 (N_8939,N_8511,N_8211);
nor U8940 (N_8940,N_8558,N_8728);
and U8941 (N_8941,N_8293,N_8347);
and U8942 (N_8942,N_8261,N_8150);
nand U8943 (N_8943,N_8459,N_8129);
xor U8944 (N_8944,N_8506,N_8594);
or U8945 (N_8945,N_8160,N_8644);
xnor U8946 (N_8946,N_8718,N_8680);
nand U8947 (N_8947,N_8286,N_8697);
nand U8948 (N_8948,N_8683,N_8346);
or U8949 (N_8949,N_8503,N_8276);
nor U8950 (N_8950,N_8663,N_8125);
nor U8951 (N_8951,N_8388,N_8174);
and U8952 (N_8952,N_8345,N_8491);
nand U8953 (N_8953,N_8677,N_8277);
and U8954 (N_8954,N_8484,N_8300);
xor U8955 (N_8955,N_8395,N_8614);
xor U8956 (N_8956,N_8188,N_8645);
nor U8957 (N_8957,N_8705,N_8487);
nand U8958 (N_8958,N_8496,N_8134);
nand U8959 (N_8959,N_8507,N_8445);
or U8960 (N_8960,N_8661,N_8288);
and U8961 (N_8961,N_8403,N_8162);
and U8962 (N_8962,N_8154,N_8495);
nor U8963 (N_8963,N_8457,N_8588);
xor U8964 (N_8964,N_8254,N_8222);
nand U8965 (N_8965,N_8227,N_8664);
or U8966 (N_8966,N_8540,N_8727);
or U8967 (N_8967,N_8303,N_8431);
and U8968 (N_8968,N_8258,N_8604);
or U8969 (N_8969,N_8419,N_8708);
xnor U8970 (N_8970,N_8398,N_8315);
nor U8971 (N_8971,N_8281,N_8646);
nor U8972 (N_8972,N_8437,N_8178);
xnor U8973 (N_8973,N_8526,N_8500);
or U8974 (N_8974,N_8357,N_8299);
or U8975 (N_8975,N_8337,N_8662);
nand U8976 (N_8976,N_8264,N_8387);
nand U8977 (N_8977,N_8305,N_8165);
xnor U8978 (N_8978,N_8428,N_8479);
nand U8979 (N_8979,N_8498,N_8706);
xnor U8980 (N_8980,N_8358,N_8742);
and U8981 (N_8981,N_8748,N_8396);
nand U8982 (N_8982,N_8607,N_8634);
and U8983 (N_8983,N_8309,N_8278);
or U8984 (N_8984,N_8439,N_8236);
nor U8985 (N_8985,N_8231,N_8280);
nor U8986 (N_8986,N_8521,N_8581);
and U8987 (N_8987,N_8658,N_8145);
and U8988 (N_8988,N_8591,N_8719);
nor U8989 (N_8989,N_8572,N_8545);
nand U8990 (N_8990,N_8285,N_8168);
or U8991 (N_8991,N_8620,N_8550);
xnor U8992 (N_8992,N_8333,N_8148);
nand U8993 (N_8993,N_8184,N_8518);
xnor U8994 (N_8994,N_8327,N_8142);
nor U8995 (N_8995,N_8464,N_8537);
or U8996 (N_8996,N_8569,N_8519);
or U8997 (N_8997,N_8635,N_8141);
nand U8998 (N_8998,N_8172,N_8551);
xnor U8999 (N_8999,N_8427,N_8425);
xnor U9000 (N_9000,N_8541,N_8466);
and U9001 (N_9001,N_8265,N_8527);
or U9002 (N_9002,N_8449,N_8177);
nand U9003 (N_9003,N_8266,N_8366);
or U9004 (N_9004,N_8271,N_8364);
nand U9005 (N_9005,N_8749,N_8557);
xnor U9006 (N_9006,N_8341,N_8167);
xnor U9007 (N_9007,N_8436,N_8497);
and U9008 (N_9008,N_8369,N_8282);
xor U9009 (N_9009,N_8666,N_8394);
and U9010 (N_9010,N_8637,N_8686);
nand U9011 (N_9011,N_8139,N_8426);
and U9012 (N_9012,N_8201,N_8618);
nor U9013 (N_9013,N_8233,N_8505);
xor U9014 (N_9014,N_8656,N_8410);
nor U9015 (N_9015,N_8126,N_8601);
nor U9016 (N_9016,N_8334,N_8147);
nand U9017 (N_9017,N_8304,N_8725);
xnor U9018 (N_9018,N_8399,N_8368);
xnor U9019 (N_9019,N_8547,N_8128);
nor U9020 (N_9020,N_8470,N_8156);
xnor U9021 (N_9021,N_8224,N_8687);
nor U9022 (N_9022,N_8269,N_8405);
nand U9023 (N_9023,N_8597,N_8546);
nor U9024 (N_9024,N_8438,N_8652);
and U9025 (N_9025,N_8482,N_8515);
or U9026 (N_9026,N_8291,N_8379);
or U9027 (N_9027,N_8481,N_8712);
or U9028 (N_9028,N_8736,N_8164);
nand U9029 (N_9029,N_8489,N_8681);
and U9030 (N_9030,N_8392,N_8332);
and U9031 (N_9031,N_8158,N_8536);
nor U9032 (N_9032,N_8590,N_8127);
and U9033 (N_9033,N_8219,N_8733);
nor U9034 (N_9034,N_8443,N_8564);
xnor U9035 (N_9035,N_8163,N_8685);
or U9036 (N_9036,N_8562,N_8538);
or U9037 (N_9037,N_8407,N_8376);
or U9038 (N_9038,N_8331,N_8239);
nand U9039 (N_9039,N_8616,N_8486);
xnor U9040 (N_9040,N_8524,N_8230);
nor U9041 (N_9041,N_8678,N_8340);
and U9042 (N_9042,N_8567,N_8583);
nand U9043 (N_9043,N_8290,N_8274);
or U9044 (N_9044,N_8600,N_8292);
nand U9045 (N_9045,N_8707,N_8313);
and U9046 (N_9046,N_8528,N_8679);
or U9047 (N_9047,N_8693,N_8704);
or U9048 (N_9048,N_8689,N_8408);
and U9049 (N_9049,N_8587,N_8668);
and U9050 (N_9050,N_8525,N_8385);
nor U9051 (N_9051,N_8692,N_8722);
nor U9052 (N_9052,N_8502,N_8648);
xnor U9053 (N_9053,N_8216,N_8328);
or U9054 (N_9054,N_8312,N_8476);
nor U9055 (N_9055,N_8275,N_8423);
and U9056 (N_9056,N_8246,N_8199);
and U9057 (N_9057,N_8202,N_8561);
nand U9058 (N_9058,N_8198,N_8446);
nor U9059 (N_9059,N_8651,N_8623);
xor U9060 (N_9060,N_8653,N_8714);
xor U9061 (N_9061,N_8157,N_8520);
and U9062 (N_9062,N_8375,N_8640);
nor U9063 (N_9063,N_8544,N_8431);
and U9064 (N_9064,N_8710,N_8418);
nand U9065 (N_9065,N_8603,N_8292);
nor U9066 (N_9066,N_8178,N_8549);
and U9067 (N_9067,N_8715,N_8441);
nand U9068 (N_9068,N_8668,N_8728);
nand U9069 (N_9069,N_8496,N_8670);
xor U9070 (N_9070,N_8173,N_8424);
xnor U9071 (N_9071,N_8280,N_8590);
nand U9072 (N_9072,N_8707,N_8653);
xnor U9073 (N_9073,N_8202,N_8218);
and U9074 (N_9074,N_8733,N_8225);
and U9075 (N_9075,N_8727,N_8315);
and U9076 (N_9076,N_8643,N_8633);
xor U9077 (N_9077,N_8387,N_8392);
nand U9078 (N_9078,N_8504,N_8204);
nor U9079 (N_9079,N_8250,N_8572);
xnor U9080 (N_9080,N_8484,N_8312);
nand U9081 (N_9081,N_8561,N_8433);
nand U9082 (N_9082,N_8580,N_8410);
or U9083 (N_9083,N_8489,N_8694);
nand U9084 (N_9084,N_8193,N_8606);
xor U9085 (N_9085,N_8268,N_8334);
or U9086 (N_9086,N_8241,N_8531);
and U9087 (N_9087,N_8397,N_8521);
and U9088 (N_9088,N_8215,N_8656);
nand U9089 (N_9089,N_8662,N_8484);
xor U9090 (N_9090,N_8606,N_8408);
or U9091 (N_9091,N_8471,N_8714);
and U9092 (N_9092,N_8401,N_8499);
nand U9093 (N_9093,N_8646,N_8227);
or U9094 (N_9094,N_8676,N_8180);
nor U9095 (N_9095,N_8486,N_8459);
nand U9096 (N_9096,N_8621,N_8516);
nand U9097 (N_9097,N_8700,N_8485);
and U9098 (N_9098,N_8498,N_8220);
or U9099 (N_9099,N_8620,N_8270);
xnor U9100 (N_9100,N_8201,N_8285);
nand U9101 (N_9101,N_8456,N_8600);
and U9102 (N_9102,N_8711,N_8353);
nor U9103 (N_9103,N_8363,N_8570);
xor U9104 (N_9104,N_8532,N_8339);
or U9105 (N_9105,N_8220,N_8350);
nand U9106 (N_9106,N_8498,N_8280);
and U9107 (N_9107,N_8555,N_8514);
and U9108 (N_9108,N_8677,N_8295);
and U9109 (N_9109,N_8588,N_8238);
or U9110 (N_9110,N_8532,N_8267);
and U9111 (N_9111,N_8594,N_8429);
or U9112 (N_9112,N_8338,N_8551);
or U9113 (N_9113,N_8130,N_8386);
nand U9114 (N_9114,N_8649,N_8728);
and U9115 (N_9115,N_8615,N_8272);
or U9116 (N_9116,N_8640,N_8580);
nand U9117 (N_9117,N_8591,N_8706);
xor U9118 (N_9118,N_8660,N_8597);
xor U9119 (N_9119,N_8297,N_8713);
xor U9120 (N_9120,N_8582,N_8354);
xor U9121 (N_9121,N_8180,N_8402);
xnor U9122 (N_9122,N_8603,N_8632);
xor U9123 (N_9123,N_8374,N_8447);
and U9124 (N_9124,N_8187,N_8180);
or U9125 (N_9125,N_8322,N_8700);
and U9126 (N_9126,N_8319,N_8125);
nand U9127 (N_9127,N_8561,N_8607);
nand U9128 (N_9128,N_8690,N_8462);
and U9129 (N_9129,N_8632,N_8501);
and U9130 (N_9130,N_8624,N_8362);
or U9131 (N_9131,N_8394,N_8738);
or U9132 (N_9132,N_8311,N_8139);
xor U9133 (N_9133,N_8580,N_8727);
and U9134 (N_9134,N_8589,N_8170);
nor U9135 (N_9135,N_8662,N_8475);
xnor U9136 (N_9136,N_8343,N_8221);
or U9137 (N_9137,N_8290,N_8718);
nand U9138 (N_9138,N_8631,N_8361);
xnor U9139 (N_9139,N_8299,N_8209);
nor U9140 (N_9140,N_8137,N_8136);
and U9141 (N_9141,N_8485,N_8710);
xnor U9142 (N_9142,N_8236,N_8233);
xor U9143 (N_9143,N_8501,N_8265);
xor U9144 (N_9144,N_8607,N_8749);
or U9145 (N_9145,N_8391,N_8605);
nand U9146 (N_9146,N_8535,N_8386);
or U9147 (N_9147,N_8459,N_8649);
xnor U9148 (N_9148,N_8298,N_8290);
xnor U9149 (N_9149,N_8721,N_8180);
nor U9150 (N_9150,N_8257,N_8583);
or U9151 (N_9151,N_8145,N_8705);
nand U9152 (N_9152,N_8730,N_8443);
xnor U9153 (N_9153,N_8522,N_8313);
nand U9154 (N_9154,N_8439,N_8285);
nand U9155 (N_9155,N_8375,N_8407);
nor U9156 (N_9156,N_8386,N_8746);
or U9157 (N_9157,N_8195,N_8352);
and U9158 (N_9158,N_8129,N_8619);
nand U9159 (N_9159,N_8684,N_8604);
xor U9160 (N_9160,N_8525,N_8719);
nand U9161 (N_9161,N_8260,N_8347);
nor U9162 (N_9162,N_8468,N_8255);
xnor U9163 (N_9163,N_8592,N_8285);
xor U9164 (N_9164,N_8247,N_8179);
or U9165 (N_9165,N_8150,N_8419);
nor U9166 (N_9166,N_8502,N_8437);
nand U9167 (N_9167,N_8554,N_8392);
xor U9168 (N_9168,N_8504,N_8429);
and U9169 (N_9169,N_8491,N_8131);
nor U9170 (N_9170,N_8539,N_8393);
nand U9171 (N_9171,N_8345,N_8677);
nor U9172 (N_9172,N_8712,N_8551);
nand U9173 (N_9173,N_8582,N_8373);
nand U9174 (N_9174,N_8645,N_8311);
or U9175 (N_9175,N_8732,N_8552);
nor U9176 (N_9176,N_8586,N_8463);
nor U9177 (N_9177,N_8556,N_8515);
or U9178 (N_9178,N_8495,N_8127);
or U9179 (N_9179,N_8428,N_8586);
and U9180 (N_9180,N_8584,N_8236);
or U9181 (N_9181,N_8314,N_8584);
or U9182 (N_9182,N_8384,N_8734);
and U9183 (N_9183,N_8749,N_8332);
nand U9184 (N_9184,N_8638,N_8709);
or U9185 (N_9185,N_8511,N_8726);
nor U9186 (N_9186,N_8617,N_8127);
nor U9187 (N_9187,N_8479,N_8501);
nor U9188 (N_9188,N_8505,N_8608);
and U9189 (N_9189,N_8158,N_8148);
xnor U9190 (N_9190,N_8265,N_8722);
and U9191 (N_9191,N_8420,N_8403);
nor U9192 (N_9192,N_8656,N_8746);
or U9193 (N_9193,N_8742,N_8212);
nor U9194 (N_9194,N_8419,N_8136);
nand U9195 (N_9195,N_8574,N_8389);
and U9196 (N_9196,N_8650,N_8582);
nor U9197 (N_9197,N_8265,N_8706);
nand U9198 (N_9198,N_8667,N_8196);
nand U9199 (N_9199,N_8455,N_8409);
and U9200 (N_9200,N_8170,N_8505);
or U9201 (N_9201,N_8310,N_8495);
or U9202 (N_9202,N_8283,N_8288);
and U9203 (N_9203,N_8447,N_8170);
nand U9204 (N_9204,N_8673,N_8195);
nand U9205 (N_9205,N_8659,N_8601);
nand U9206 (N_9206,N_8572,N_8541);
and U9207 (N_9207,N_8604,N_8515);
and U9208 (N_9208,N_8555,N_8275);
or U9209 (N_9209,N_8567,N_8676);
nand U9210 (N_9210,N_8405,N_8191);
or U9211 (N_9211,N_8552,N_8416);
or U9212 (N_9212,N_8278,N_8373);
and U9213 (N_9213,N_8570,N_8731);
xor U9214 (N_9214,N_8146,N_8561);
nand U9215 (N_9215,N_8460,N_8565);
nor U9216 (N_9216,N_8452,N_8140);
and U9217 (N_9217,N_8558,N_8178);
xor U9218 (N_9218,N_8418,N_8233);
and U9219 (N_9219,N_8151,N_8507);
xnor U9220 (N_9220,N_8556,N_8644);
xnor U9221 (N_9221,N_8598,N_8555);
xnor U9222 (N_9222,N_8210,N_8636);
xor U9223 (N_9223,N_8528,N_8279);
nand U9224 (N_9224,N_8515,N_8559);
xor U9225 (N_9225,N_8157,N_8363);
and U9226 (N_9226,N_8453,N_8309);
or U9227 (N_9227,N_8354,N_8303);
and U9228 (N_9228,N_8717,N_8570);
xnor U9229 (N_9229,N_8513,N_8278);
nor U9230 (N_9230,N_8508,N_8340);
and U9231 (N_9231,N_8349,N_8343);
and U9232 (N_9232,N_8711,N_8312);
and U9233 (N_9233,N_8157,N_8523);
and U9234 (N_9234,N_8439,N_8329);
nor U9235 (N_9235,N_8301,N_8224);
or U9236 (N_9236,N_8386,N_8400);
or U9237 (N_9237,N_8259,N_8439);
and U9238 (N_9238,N_8618,N_8157);
or U9239 (N_9239,N_8393,N_8369);
nand U9240 (N_9240,N_8253,N_8366);
or U9241 (N_9241,N_8674,N_8157);
xor U9242 (N_9242,N_8291,N_8521);
xnor U9243 (N_9243,N_8669,N_8698);
nor U9244 (N_9244,N_8458,N_8178);
nand U9245 (N_9245,N_8615,N_8613);
and U9246 (N_9246,N_8595,N_8198);
nand U9247 (N_9247,N_8587,N_8489);
nand U9248 (N_9248,N_8285,N_8619);
and U9249 (N_9249,N_8206,N_8716);
nand U9250 (N_9250,N_8462,N_8219);
and U9251 (N_9251,N_8446,N_8533);
or U9252 (N_9252,N_8593,N_8568);
nor U9253 (N_9253,N_8165,N_8190);
nor U9254 (N_9254,N_8546,N_8231);
nor U9255 (N_9255,N_8565,N_8534);
and U9256 (N_9256,N_8580,N_8524);
nor U9257 (N_9257,N_8156,N_8212);
nor U9258 (N_9258,N_8651,N_8469);
nor U9259 (N_9259,N_8680,N_8449);
nand U9260 (N_9260,N_8206,N_8741);
nand U9261 (N_9261,N_8626,N_8301);
nor U9262 (N_9262,N_8420,N_8710);
or U9263 (N_9263,N_8651,N_8335);
or U9264 (N_9264,N_8680,N_8703);
nand U9265 (N_9265,N_8531,N_8413);
or U9266 (N_9266,N_8494,N_8205);
and U9267 (N_9267,N_8729,N_8502);
xnor U9268 (N_9268,N_8224,N_8491);
and U9269 (N_9269,N_8629,N_8144);
nand U9270 (N_9270,N_8464,N_8182);
nand U9271 (N_9271,N_8367,N_8203);
nand U9272 (N_9272,N_8163,N_8267);
nand U9273 (N_9273,N_8148,N_8302);
or U9274 (N_9274,N_8305,N_8389);
or U9275 (N_9275,N_8486,N_8637);
and U9276 (N_9276,N_8685,N_8735);
or U9277 (N_9277,N_8350,N_8715);
xor U9278 (N_9278,N_8679,N_8635);
or U9279 (N_9279,N_8405,N_8404);
and U9280 (N_9280,N_8342,N_8591);
or U9281 (N_9281,N_8574,N_8279);
or U9282 (N_9282,N_8261,N_8165);
nor U9283 (N_9283,N_8479,N_8284);
xor U9284 (N_9284,N_8294,N_8558);
or U9285 (N_9285,N_8510,N_8578);
nand U9286 (N_9286,N_8448,N_8398);
and U9287 (N_9287,N_8252,N_8680);
or U9288 (N_9288,N_8240,N_8388);
or U9289 (N_9289,N_8179,N_8168);
and U9290 (N_9290,N_8550,N_8421);
nor U9291 (N_9291,N_8378,N_8229);
nand U9292 (N_9292,N_8645,N_8563);
or U9293 (N_9293,N_8246,N_8584);
and U9294 (N_9294,N_8668,N_8710);
xnor U9295 (N_9295,N_8239,N_8538);
nand U9296 (N_9296,N_8285,N_8353);
or U9297 (N_9297,N_8306,N_8438);
xnor U9298 (N_9298,N_8701,N_8189);
and U9299 (N_9299,N_8457,N_8281);
nand U9300 (N_9300,N_8413,N_8465);
or U9301 (N_9301,N_8612,N_8286);
nor U9302 (N_9302,N_8420,N_8673);
or U9303 (N_9303,N_8745,N_8172);
and U9304 (N_9304,N_8239,N_8516);
nor U9305 (N_9305,N_8580,N_8515);
or U9306 (N_9306,N_8403,N_8539);
and U9307 (N_9307,N_8453,N_8227);
or U9308 (N_9308,N_8216,N_8496);
nand U9309 (N_9309,N_8438,N_8521);
nor U9310 (N_9310,N_8279,N_8743);
nand U9311 (N_9311,N_8285,N_8502);
nand U9312 (N_9312,N_8534,N_8550);
nand U9313 (N_9313,N_8385,N_8558);
or U9314 (N_9314,N_8375,N_8623);
and U9315 (N_9315,N_8161,N_8277);
xnor U9316 (N_9316,N_8439,N_8701);
nor U9317 (N_9317,N_8459,N_8685);
xnor U9318 (N_9318,N_8134,N_8422);
xnor U9319 (N_9319,N_8271,N_8689);
xor U9320 (N_9320,N_8509,N_8482);
or U9321 (N_9321,N_8146,N_8268);
nand U9322 (N_9322,N_8525,N_8491);
xor U9323 (N_9323,N_8293,N_8332);
nor U9324 (N_9324,N_8567,N_8619);
nand U9325 (N_9325,N_8731,N_8516);
and U9326 (N_9326,N_8625,N_8485);
nor U9327 (N_9327,N_8656,N_8609);
nor U9328 (N_9328,N_8422,N_8503);
nand U9329 (N_9329,N_8665,N_8219);
nand U9330 (N_9330,N_8126,N_8692);
xor U9331 (N_9331,N_8482,N_8697);
nor U9332 (N_9332,N_8536,N_8295);
nand U9333 (N_9333,N_8471,N_8655);
nand U9334 (N_9334,N_8485,N_8733);
nor U9335 (N_9335,N_8151,N_8624);
nand U9336 (N_9336,N_8481,N_8479);
nor U9337 (N_9337,N_8261,N_8413);
nand U9338 (N_9338,N_8447,N_8134);
xnor U9339 (N_9339,N_8382,N_8538);
and U9340 (N_9340,N_8406,N_8543);
and U9341 (N_9341,N_8167,N_8437);
or U9342 (N_9342,N_8635,N_8215);
nand U9343 (N_9343,N_8272,N_8166);
nor U9344 (N_9344,N_8652,N_8380);
xor U9345 (N_9345,N_8173,N_8360);
nand U9346 (N_9346,N_8535,N_8320);
nor U9347 (N_9347,N_8673,N_8612);
nand U9348 (N_9348,N_8250,N_8742);
nor U9349 (N_9349,N_8230,N_8128);
nand U9350 (N_9350,N_8671,N_8193);
or U9351 (N_9351,N_8582,N_8282);
and U9352 (N_9352,N_8317,N_8709);
nand U9353 (N_9353,N_8141,N_8409);
xor U9354 (N_9354,N_8610,N_8556);
xor U9355 (N_9355,N_8415,N_8299);
xor U9356 (N_9356,N_8209,N_8384);
or U9357 (N_9357,N_8419,N_8481);
nand U9358 (N_9358,N_8132,N_8745);
nor U9359 (N_9359,N_8683,N_8598);
nor U9360 (N_9360,N_8382,N_8504);
nand U9361 (N_9361,N_8417,N_8543);
xor U9362 (N_9362,N_8688,N_8389);
nand U9363 (N_9363,N_8376,N_8385);
and U9364 (N_9364,N_8737,N_8516);
xor U9365 (N_9365,N_8212,N_8710);
and U9366 (N_9366,N_8649,N_8481);
or U9367 (N_9367,N_8129,N_8574);
nor U9368 (N_9368,N_8599,N_8316);
nor U9369 (N_9369,N_8399,N_8690);
and U9370 (N_9370,N_8368,N_8563);
or U9371 (N_9371,N_8525,N_8656);
nand U9372 (N_9372,N_8454,N_8161);
nor U9373 (N_9373,N_8653,N_8568);
xor U9374 (N_9374,N_8314,N_8747);
nor U9375 (N_9375,N_9185,N_9034);
and U9376 (N_9376,N_8957,N_8830);
xnor U9377 (N_9377,N_9148,N_8887);
nor U9378 (N_9378,N_9289,N_8763);
nand U9379 (N_9379,N_8949,N_8845);
nand U9380 (N_9380,N_9004,N_9090);
nand U9381 (N_9381,N_8786,N_9254);
and U9382 (N_9382,N_9044,N_9039);
nand U9383 (N_9383,N_8753,N_9010);
and U9384 (N_9384,N_9271,N_8883);
nand U9385 (N_9385,N_9323,N_9241);
and U9386 (N_9386,N_9312,N_9325);
xor U9387 (N_9387,N_9250,N_8965);
or U9388 (N_9388,N_9013,N_8781);
nand U9389 (N_9389,N_8877,N_8927);
and U9390 (N_9390,N_8969,N_8913);
and U9391 (N_9391,N_9098,N_8878);
or U9392 (N_9392,N_9103,N_8922);
or U9393 (N_9393,N_9248,N_9278);
xor U9394 (N_9394,N_9131,N_9057);
or U9395 (N_9395,N_9333,N_8910);
or U9396 (N_9396,N_8842,N_9163);
or U9397 (N_9397,N_9229,N_9372);
and U9398 (N_9398,N_8987,N_8950);
nor U9399 (N_9399,N_8793,N_9210);
or U9400 (N_9400,N_8779,N_9201);
nor U9401 (N_9401,N_8975,N_9240);
nand U9402 (N_9402,N_9005,N_9180);
or U9403 (N_9403,N_9128,N_8798);
nand U9404 (N_9404,N_9002,N_8939);
nor U9405 (N_9405,N_8903,N_8967);
and U9406 (N_9406,N_9107,N_9202);
nand U9407 (N_9407,N_9172,N_9169);
and U9408 (N_9408,N_9161,N_8937);
and U9409 (N_9409,N_9233,N_9246);
nand U9410 (N_9410,N_8925,N_9188);
nor U9411 (N_9411,N_9213,N_9125);
xor U9412 (N_9412,N_9313,N_9072);
nand U9413 (N_9413,N_8963,N_9030);
nand U9414 (N_9414,N_9339,N_9369);
nand U9415 (N_9415,N_9095,N_8876);
and U9416 (N_9416,N_8964,N_9287);
xnor U9417 (N_9417,N_9165,N_9054);
xnor U9418 (N_9418,N_9171,N_9359);
xor U9419 (N_9419,N_8797,N_8759);
and U9420 (N_9420,N_9176,N_8974);
nor U9421 (N_9421,N_9156,N_9230);
xnor U9422 (N_9422,N_9087,N_8981);
nor U9423 (N_9423,N_8778,N_9177);
and U9424 (N_9424,N_8962,N_8853);
and U9425 (N_9425,N_8912,N_9194);
or U9426 (N_9426,N_9112,N_9298);
or U9427 (N_9427,N_8952,N_8995);
or U9428 (N_9428,N_8931,N_9282);
xor U9429 (N_9429,N_8914,N_9129);
and U9430 (N_9430,N_8960,N_8791);
nor U9431 (N_9431,N_9108,N_9138);
or U9432 (N_9432,N_9249,N_8892);
nor U9433 (N_9433,N_9170,N_8889);
or U9434 (N_9434,N_8896,N_8776);
and U9435 (N_9435,N_8806,N_9243);
or U9436 (N_9436,N_9142,N_8819);
nand U9437 (N_9437,N_9206,N_9269);
or U9438 (N_9438,N_8758,N_9152);
nand U9439 (N_9439,N_9050,N_8849);
xnor U9440 (N_9440,N_8770,N_8788);
xnor U9441 (N_9441,N_9062,N_9196);
xnor U9442 (N_9442,N_9366,N_8915);
xor U9443 (N_9443,N_9264,N_9024);
nor U9444 (N_9444,N_9012,N_8924);
nor U9445 (N_9445,N_9166,N_9017);
nor U9446 (N_9446,N_9292,N_8886);
xnor U9447 (N_9447,N_9370,N_8795);
or U9448 (N_9448,N_9094,N_9299);
nor U9449 (N_9449,N_9231,N_9154);
and U9450 (N_9450,N_9190,N_9173);
and U9451 (N_9451,N_9367,N_9046);
and U9452 (N_9452,N_9033,N_8901);
or U9453 (N_9453,N_8800,N_9355);
nand U9454 (N_9454,N_8751,N_9056);
or U9455 (N_9455,N_9191,N_8787);
or U9456 (N_9456,N_9330,N_9295);
nand U9457 (N_9457,N_8916,N_9351);
or U9458 (N_9458,N_8828,N_9350);
xor U9459 (N_9459,N_8909,N_9018);
or U9460 (N_9460,N_9209,N_9025);
and U9461 (N_9461,N_9301,N_9096);
xnor U9462 (N_9462,N_9263,N_8769);
or U9463 (N_9463,N_9327,N_8900);
and U9464 (N_9464,N_9253,N_9212);
nand U9465 (N_9465,N_8825,N_8832);
nor U9466 (N_9466,N_9311,N_8820);
or U9467 (N_9467,N_9214,N_8941);
nor U9468 (N_9468,N_8888,N_9146);
xor U9469 (N_9469,N_9257,N_9360);
or U9470 (N_9470,N_9089,N_8784);
nor U9471 (N_9471,N_9110,N_8998);
and U9472 (N_9472,N_8997,N_8902);
nand U9473 (N_9473,N_9310,N_8771);
xor U9474 (N_9474,N_8891,N_9097);
nand U9475 (N_9475,N_9309,N_9133);
xor U9476 (N_9476,N_8934,N_9260);
nor U9477 (N_9477,N_8968,N_9078);
or U9478 (N_9478,N_9184,N_9265);
nand U9479 (N_9479,N_9235,N_8955);
or U9480 (N_9480,N_8948,N_8966);
or U9481 (N_9481,N_9092,N_9134);
nand U9482 (N_9482,N_8993,N_8996);
nand U9483 (N_9483,N_8855,N_9199);
xnor U9484 (N_9484,N_8928,N_8917);
and U9485 (N_9485,N_8821,N_8765);
or U9486 (N_9486,N_9223,N_9071);
and U9487 (N_9487,N_9181,N_8761);
nand U9488 (N_9488,N_9014,N_8813);
and U9489 (N_9489,N_8864,N_9284);
xnor U9490 (N_9490,N_8989,N_9322);
nand U9491 (N_9491,N_9186,N_9140);
xnor U9492 (N_9492,N_9337,N_8834);
nor U9493 (N_9493,N_8847,N_9279);
nand U9494 (N_9494,N_8792,N_9127);
nor U9495 (N_9495,N_8810,N_8841);
nor U9496 (N_9496,N_8890,N_8873);
nor U9497 (N_9497,N_9053,N_9082);
and U9498 (N_9498,N_9200,N_8768);
and U9499 (N_9499,N_9346,N_9175);
or U9500 (N_9500,N_9160,N_9075);
or U9501 (N_9501,N_8844,N_9373);
xor U9502 (N_9502,N_9168,N_8794);
or U9503 (N_9503,N_8971,N_9300);
nor U9504 (N_9504,N_8951,N_9315);
nand U9505 (N_9505,N_9036,N_8970);
and U9506 (N_9506,N_8846,N_9136);
and U9507 (N_9507,N_8838,N_9028);
xnor U9508 (N_9508,N_8837,N_8980);
xor U9509 (N_9509,N_9324,N_8992);
nor U9510 (N_9510,N_9023,N_9042);
xnor U9511 (N_9511,N_9363,N_9218);
and U9512 (N_9512,N_9041,N_8945);
nand U9513 (N_9513,N_9354,N_8946);
nor U9514 (N_9514,N_8857,N_8852);
xnor U9515 (N_9515,N_8803,N_8918);
or U9516 (N_9516,N_8826,N_8868);
nand U9517 (N_9517,N_9123,N_9204);
or U9518 (N_9518,N_9081,N_9321);
and U9519 (N_9519,N_8920,N_9247);
nor U9520 (N_9520,N_8822,N_9357);
and U9521 (N_9521,N_8907,N_8984);
or U9522 (N_9522,N_8760,N_8986);
nand U9523 (N_9523,N_8782,N_9232);
and U9524 (N_9524,N_9043,N_9244);
nand U9525 (N_9525,N_9085,N_9007);
nor U9526 (N_9526,N_8942,N_9045);
xnor U9527 (N_9527,N_8783,N_9109);
and U9528 (N_9528,N_9114,N_8932);
and U9529 (N_9529,N_8839,N_9280);
nand U9530 (N_9530,N_9237,N_9022);
and U9531 (N_9531,N_9008,N_9368);
and U9532 (N_9532,N_8911,N_9353);
and U9533 (N_9533,N_9222,N_8898);
and U9534 (N_9534,N_8988,N_8956);
xnor U9535 (N_9535,N_9197,N_9015);
nor U9536 (N_9536,N_8843,N_9352);
nand U9537 (N_9537,N_8812,N_8863);
or U9538 (N_9538,N_9126,N_9162);
and U9539 (N_9539,N_9091,N_8789);
and U9540 (N_9540,N_9343,N_8762);
and U9541 (N_9541,N_9066,N_8978);
xor U9542 (N_9542,N_9093,N_9281);
nor U9543 (N_9543,N_9297,N_9167);
nor U9544 (N_9544,N_9317,N_8840);
and U9545 (N_9545,N_9319,N_8895);
xnor U9546 (N_9546,N_9258,N_8954);
xnor U9547 (N_9547,N_9285,N_9100);
nor U9548 (N_9548,N_8919,N_8767);
or U9549 (N_9549,N_9151,N_9203);
and U9550 (N_9550,N_8985,N_8860);
or U9551 (N_9551,N_9251,N_9195);
nand U9552 (N_9552,N_9228,N_8871);
nor U9553 (N_9553,N_9088,N_8755);
and U9554 (N_9554,N_9174,N_9051);
nand U9555 (N_9555,N_9032,N_8959);
and U9556 (N_9556,N_8850,N_8930);
and U9557 (N_9557,N_8811,N_9349);
and U9558 (N_9558,N_8777,N_9242);
and U9559 (N_9559,N_9335,N_9155);
or U9560 (N_9560,N_8817,N_8823);
xor U9561 (N_9561,N_9238,N_9067);
nand U9562 (N_9562,N_8833,N_9358);
xnor U9563 (N_9563,N_8929,N_8874);
or U9564 (N_9564,N_9193,N_8861);
or U9565 (N_9565,N_8867,N_8879);
nor U9566 (N_9566,N_9104,N_8936);
and U9567 (N_9567,N_8977,N_8953);
and U9568 (N_9568,N_8870,N_8897);
nor U9569 (N_9569,N_9048,N_9275);
or U9570 (N_9570,N_9326,N_9117);
nand U9571 (N_9571,N_9000,N_9187);
or U9572 (N_9572,N_9020,N_9016);
or U9573 (N_9573,N_9215,N_9049);
xor U9574 (N_9574,N_8872,N_8848);
or U9575 (N_9575,N_9189,N_9274);
or U9576 (N_9576,N_9118,N_9307);
or U9577 (N_9577,N_8772,N_9304);
xor U9578 (N_9578,N_8836,N_8869);
nor U9579 (N_9579,N_9113,N_8815);
and U9580 (N_9580,N_9021,N_9308);
nand U9581 (N_9581,N_9080,N_9035);
xnor U9582 (N_9582,N_9273,N_8906);
nand U9583 (N_9583,N_9306,N_9320);
nand U9584 (N_9584,N_8799,N_9341);
nand U9585 (N_9585,N_8804,N_8790);
and U9586 (N_9586,N_9141,N_9277);
and U9587 (N_9587,N_9347,N_8851);
or U9588 (N_9588,N_9120,N_9064);
nand U9589 (N_9589,N_8809,N_9219);
or U9590 (N_9590,N_9101,N_9009);
nand U9591 (N_9591,N_9291,N_9083);
nor U9592 (N_9592,N_9374,N_9122);
xnor U9593 (N_9593,N_8994,N_9371);
nor U9594 (N_9594,N_8827,N_9314);
nor U9595 (N_9595,N_9236,N_8785);
nand U9596 (N_9596,N_9331,N_9006);
and U9597 (N_9597,N_8983,N_9038);
or U9598 (N_9598,N_8979,N_8862);
nor U9599 (N_9599,N_9255,N_9065);
and U9600 (N_9600,N_9305,N_9245);
or U9601 (N_9601,N_9059,N_8858);
nor U9602 (N_9602,N_8866,N_8766);
or U9603 (N_9603,N_9058,N_9261);
nand U9604 (N_9604,N_9061,N_9227);
nand U9605 (N_9605,N_9149,N_8961);
and U9606 (N_9606,N_9001,N_8816);
and U9607 (N_9607,N_9115,N_9294);
and U9608 (N_9608,N_9124,N_8921);
nor U9609 (N_9609,N_9040,N_9029);
nor U9610 (N_9610,N_9334,N_8775);
and U9611 (N_9611,N_9060,N_9052);
and U9612 (N_9612,N_8835,N_8808);
or U9613 (N_9613,N_9147,N_9198);
or U9614 (N_9614,N_9266,N_9365);
and U9615 (N_9615,N_8893,N_8947);
or U9616 (N_9616,N_9074,N_8976);
xnor U9617 (N_9617,N_9328,N_9150);
nor U9618 (N_9618,N_9272,N_9207);
or U9619 (N_9619,N_9217,N_8814);
or U9620 (N_9620,N_8773,N_9132);
xor U9621 (N_9621,N_9216,N_8973);
and U9622 (N_9622,N_8894,N_8859);
and U9623 (N_9623,N_9340,N_9288);
nand U9624 (N_9624,N_8764,N_9286);
nor U9625 (N_9625,N_8885,N_9031);
nand U9626 (N_9626,N_8756,N_9290);
or U9627 (N_9627,N_9073,N_9135);
xor U9628 (N_9628,N_9178,N_9296);
and U9629 (N_9629,N_9262,N_8865);
xor U9630 (N_9630,N_9111,N_8935);
or U9631 (N_9631,N_9205,N_9344);
or U9632 (N_9632,N_8750,N_9130);
or U9633 (N_9633,N_9342,N_9119);
or U9634 (N_9634,N_9037,N_8940);
and U9635 (N_9635,N_8933,N_9106);
nor U9636 (N_9636,N_8801,N_9164);
or U9637 (N_9637,N_9077,N_9293);
xnor U9638 (N_9638,N_9143,N_9268);
xnor U9639 (N_9639,N_9179,N_9139);
or U9640 (N_9640,N_9105,N_9225);
xnor U9641 (N_9641,N_9283,N_8829);
xor U9642 (N_9642,N_9026,N_9157);
and U9643 (N_9643,N_9084,N_9027);
nor U9644 (N_9644,N_9302,N_9356);
or U9645 (N_9645,N_9332,N_8831);
or U9646 (N_9646,N_9137,N_8752);
nor U9647 (N_9647,N_8854,N_9252);
or U9648 (N_9648,N_9364,N_8944);
or U9649 (N_9649,N_8904,N_9259);
nand U9650 (N_9650,N_8880,N_9086);
nand U9651 (N_9651,N_8926,N_9336);
xnor U9652 (N_9652,N_9220,N_8991);
nand U9653 (N_9653,N_9158,N_9182);
xor U9654 (N_9654,N_9318,N_8884);
and U9655 (N_9655,N_9145,N_8818);
nor U9656 (N_9656,N_9361,N_8982);
and U9657 (N_9657,N_8958,N_8938);
nand U9658 (N_9658,N_9121,N_9076);
nand U9659 (N_9659,N_9270,N_9047);
nor U9660 (N_9660,N_9102,N_9063);
and U9661 (N_9661,N_8875,N_9226);
and U9662 (N_9662,N_9192,N_8999);
and U9663 (N_9663,N_9153,N_8780);
xor U9664 (N_9664,N_9348,N_9316);
nor U9665 (N_9665,N_9068,N_9211);
or U9666 (N_9666,N_8796,N_9003);
nor U9667 (N_9667,N_9338,N_9276);
nor U9668 (N_9668,N_8923,N_9099);
nand U9669 (N_9669,N_9224,N_9329);
xnor U9670 (N_9670,N_9303,N_8757);
and U9671 (N_9671,N_8754,N_9234);
and U9672 (N_9672,N_9362,N_9019);
or U9673 (N_9673,N_8943,N_9011);
or U9674 (N_9674,N_9183,N_9069);
xnor U9675 (N_9675,N_9159,N_8881);
or U9676 (N_9676,N_8824,N_8990);
and U9677 (N_9677,N_8972,N_9055);
or U9678 (N_9678,N_9256,N_8805);
xnor U9679 (N_9679,N_9208,N_8882);
nand U9680 (N_9680,N_9221,N_8908);
nand U9681 (N_9681,N_9239,N_9116);
and U9682 (N_9682,N_8899,N_8905);
or U9683 (N_9683,N_8802,N_9144);
nor U9684 (N_9684,N_8856,N_9070);
and U9685 (N_9685,N_9267,N_8807);
nor U9686 (N_9686,N_8774,N_9079);
xor U9687 (N_9687,N_9345,N_8799);
or U9688 (N_9688,N_8945,N_8808);
nand U9689 (N_9689,N_9033,N_8767);
xnor U9690 (N_9690,N_9100,N_9262);
nor U9691 (N_9691,N_8849,N_9106);
and U9692 (N_9692,N_9226,N_9367);
nand U9693 (N_9693,N_8792,N_8870);
and U9694 (N_9694,N_9162,N_9005);
nor U9695 (N_9695,N_9124,N_9031);
nand U9696 (N_9696,N_8861,N_8901);
or U9697 (N_9697,N_9052,N_8989);
nor U9698 (N_9698,N_9287,N_9109);
and U9699 (N_9699,N_8831,N_8914);
xor U9700 (N_9700,N_8988,N_8960);
or U9701 (N_9701,N_9201,N_8754);
xor U9702 (N_9702,N_9050,N_9082);
or U9703 (N_9703,N_9183,N_8807);
and U9704 (N_9704,N_8942,N_8868);
nor U9705 (N_9705,N_9245,N_9044);
nand U9706 (N_9706,N_9266,N_9082);
nor U9707 (N_9707,N_9083,N_8769);
xnor U9708 (N_9708,N_9104,N_8871);
and U9709 (N_9709,N_9181,N_9209);
or U9710 (N_9710,N_8779,N_9066);
and U9711 (N_9711,N_8843,N_9137);
or U9712 (N_9712,N_9049,N_9128);
or U9713 (N_9713,N_9321,N_9106);
and U9714 (N_9714,N_8819,N_9233);
nor U9715 (N_9715,N_8961,N_8998);
nor U9716 (N_9716,N_8799,N_8800);
nand U9717 (N_9717,N_8905,N_8804);
and U9718 (N_9718,N_9321,N_9047);
xor U9719 (N_9719,N_8956,N_9124);
and U9720 (N_9720,N_9012,N_9303);
nand U9721 (N_9721,N_9098,N_8984);
nand U9722 (N_9722,N_9056,N_9340);
and U9723 (N_9723,N_9079,N_9204);
or U9724 (N_9724,N_8994,N_9281);
and U9725 (N_9725,N_9291,N_8869);
xor U9726 (N_9726,N_9290,N_9115);
nor U9727 (N_9727,N_8796,N_8988);
and U9728 (N_9728,N_8972,N_9009);
and U9729 (N_9729,N_8980,N_9105);
or U9730 (N_9730,N_8893,N_9011);
xnor U9731 (N_9731,N_8799,N_9182);
nor U9732 (N_9732,N_9014,N_9133);
xnor U9733 (N_9733,N_8837,N_8853);
nand U9734 (N_9734,N_9080,N_9139);
and U9735 (N_9735,N_9370,N_9173);
or U9736 (N_9736,N_8886,N_8984);
xnor U9737 (N_9737,N_8971,N_9018);
xnor U9738 (N_9738,N_8949,N_8948);
nor U9739 (N_9739,N_9029,N_9236);
xor U9740 (N_9740,N_9090,N_8966);
or U9741 (N_9741,N_9282,N_9236);
and U9742 (N_9742,N_9225,N_8920);
nand U9743 (N_9743,N_9333,N_8973);
and U9744 (N_9744,N_8999,N_8989);
and U9745 (N_9745,N_9248,N_8830);
or U9746 (N_9746,N_9087,N_8816);
nor U9747 (N_9747,N_8933,N_9191);
nor U9748 (N_9748,N_9143,N_9248);
or U9749 (N_9749,N_9197,N_8999);
and U9750 (N_9750,N_8815,N_8838);
nor U9751 (N_9751,N_8893,N_9338);
nand U9752 (N_9752,N_9027,N_8931);
nor U9753 (N_9753,N_8782,N_8940);
or U9754 (N_9754,N_9203,N_9193);
nor U9755 (N_9755,N_8928,N_8984);
nand U9756 (N_9756,N_8782,N_8985);
nor U9757 (N_9757,N_9151,N_8958);
nor U9758 (N_9758,N_9344,N_9079);
or U9759 (N_9759,N_8920,N_8751);
and U9760 (N_9760,N_8966,N_9187);
xnor U9761 (N_9761,N_8891,N_8847);
nor U9762 (N_9762,N_9108,N_9230);
and U9763 (N_9763,N_9317,N_8761);
nand U9764 (N_9764,N_9271,N_8891);
and U9765 (N_9765,N_8875,N_8836);
xor U9766 (N_9766,N_9307,N_9272);
nand U9767 (N_9767,N_8846,N_8797);
or U9768 (N_9768,N_9004,N_8925);
nand U9769 (N_9769,N_9351,N_9061);
and U9770 (N_9770,N_8884,N_9137);
nor U9771 (N_9771,N_8807,N_9178);
nor U9772 (N_9772,N_8875,N_9224);
nor U9773 (N_9773,N_9201,N_9119);
or U9774 (N_9774,N_9055,N_9208);
or U9775 (N_9775,N_9241,N_9021);
nor U9776 (N_9776,N_9295,N_9006);
nor U9777 (N_9777,N_9290,N_9298);
nor U9778 (N_9778,N_8942,N_8874);
or U9779 (N_9779,N_9218,N_9265);
nand U9780 (N_9780,N_9345,N_9245);
and U9781 (N_9781,N_9258,N_8839);
nor U9782 (N_9782,N_9213,N_9315);
xnor U9783 (N_9783,N_9325,N_8764);
nand U9784 (N_9784,N_9081,N_9240);
nand U9785 (N_9785,N_9335,N_9305);
xnor U9786 (N_9786,N_9051,N_9256);
xnor U9787 (N_9787,N_8979,N_9290);
and U9788 (N_9788,N_8864,N_8791);
xor U9789 (N_9789,N_8760,N_9277);
nor U9790 (N_9790,N_9046,N_9081);
or U9791 (N_9791,N_9228,N_9076);
nor U9792 (N_9792,N_8969,N_8833);
nand U9793 (N_9793,N_9110,N_8751);
nor U9794 (N_9794,N_8776,N_9318);
xor U9795 (N_9795,N_9031,N_8867);
and U9796 (N_9796,N_9257,N_8781);
nor U9797 (N_9797,N_8805,N_9027);
and U9798 (N_9798,N_9064,N_8825);
nor U9799 (N_9799,N_9001,N_8805);
nor U9800 (N_9800,N_8775,N_9352);
xnor U9801 (N_9801,N_8860,N_9353);
or U9802 (N_9802,N_8932,N_9302);
and U9803 (N_9803,N_8904,N_9226);
and U9804 (N_9804,N_9016,N_8988);
or U9805 (N_9805,N_8871,N_9137);
xor U9806 (N_9806,N_9179,N_9300);
or U9807 (N_9807,N_9007,N_8988);
nor U9808 (N_9808,N_9001,N_8830);
xnor U9809 (N_9809,N_8766,N_8821);
nand U9810 (N_9810,N_9052,N_8830);
xor U9811 (N_9811,N_8910,N_9325);
nand U9812 (N_9812,N_9169,N_9363);
nand U9813 (N_9813,N_8968,N_8907);
or U9814 (N_9814,N_9354,N_9029);
nor U9815 (N_9815,N_9304,N_8983);
or U9816 (N_9816,N_8959,N_9113);
xnor U9817 (N_9817,N_8986,N_9333);
nand U9818 (N_9818,N_8845,N_9062);
nand U9819 (N_9819,N_9059,N_9037);
xor U9820 (N_9820,N_9097,N_9049);
nand U9821 (N_9821,N_9189,N_9210);
nand U9822 (N_9822,N_8988,N_9160);
xnor U9823 (N_9823,N_9295,N_8969);
nand U9824 (N_9824,N_9035,N_9152);
xor U9825 (N_9825,N_8858,N_8752);
xnor U9826 (N_9826,N_9130,N_8863);
nor U9827 (N_9827,N_9355,N_9182);
and U9828 (N_9828,N_8948,N_9176);
nor U9829 (N_9829,N_9062,N_9117);
xor U9830 (N_9830,N_8799,N_9152);
xor U9831 (N_9831,N_8782,N_9240);
and U9832 (N_9832,N_9276,N_9218);
xnor U9833 (N_9833,N_9105,N_9114);
nor U9834 (N_9834,N_9141,N_9317);
or U9835 (N_9835,N_9058,N_9352);
and U9836 (N_9836,N_9130,N_8868);
nor U9837 (N_9837,N_9324,N_8832);
nor U9838 (N_9838,N_9158,N_9336);
or U9839 (N_9839,N_9235,N_8943);
nand U9840 (N_9840,N_9359,N_8787);
or U9841 (N_9841,N_9139,N_8983);
nor U9842 (N_9842,N_9007,N_8758);
or U9843 (N_9843,N_8798,N_8983);
xnor U9844 (N_9844,N_9223,N_9068);
nand U9845 (N_9845,N_8958,N_9012);
and U9846 (N_9846,N_8843,N_9083);
nand U9847 (N_9847,N_8973,N_8761);
nor U9848 (N_9848,N_9364,N_9300);
and U9849 (N_9849,N_9280,N_8851);
xnor U9850 (N_9850,N_8776,N_9347);
xnor U9851 (N_9851,N_8934,N_9023);
nand U9852 (N_9852,N_9036,N_9030);
or U9853 (N_9853,N_9050,N_8756);
and U9854 (N_9854,N_9320,N_8904);
xnor U9855 (N_9855,N_8822,N_9085);
nor U9856 (N_9856,N_9080,N_9234);
and U9857 (N_9857,N_9064,N_8874);
nor U9858 (N_9858,N_9105,N_9368);
nor U9859 (N_9859,N_8792,N_8807);
and U9860 (N_9860,N_8810,N_8947);
or U9861 (N_9861,N_9268,N_9157);
and U9862 (N_9862,N_9188,N_8757);
nand U9863 (N_9863,N_9009,N_9075);
xor U9864 (N_9864,N_9123,N_9024);
and U9865 (N_9865,N_9279,N_9326);
nor U9866 (N_9866,N_8852,N_9237);
and U9867 (N_9867,N_8817,N_8973);
nand U9868 (N_9868,N_8790,N_9213);
or U9869 (N_9869,N_9241,N_9102);
and U9870 (N_9870,N_8838,N_9284);
nand U9871 (N_9871,N_8990,N_9295);
nor U9872 (N_9872,N_9344,N_9234);
and U9873 (N_9873,N_8879,N_9003);
xor U9874 (N_9874,N_9130,N_8860);
and U9875 (N_9875,N_8779,N_9117);
or U9876 (N_9876,N_9041,N_9023);
xnor U9877 (N_9877,N_9186,N_9204);
nor U9878 (N_9878,N_8765,N_9282);
xor U9879 (N_9879,N_9295,N_8834);
nor U9880 (N_9880,N_9199,N_8997);
and U9881 (N_9881,N_8918,N_8989);
nand U9882 (N_9882,N_8913,N_8892);
and U9883 (N_9883,N_9193,N_9212);
nor U9884 (N_9884,N_8803,N_9313);
nand U9885 (N_9885,N_9088,N_8765);
or U9886 (N_9886,N_8899,N_9186);
nand U9887 (N_9887,N_9194,N_9082);
and U9888 (N_9888,N_9271,N_8991);
nand U9889 (N_9889,N_9034,N_9096);
or U9890 (N_9890,N_9212,N_8842);
nand U9891 (N_9891,N_9045,N_9022);
nor U9892 (N_9892,N_9274,N_9266);
or U9893 (N_9893,N_9073,N_9303);
and U9894 (N_9894,N_8994,N_9042);
or U9895 (N_9895,N_8844,N_8956);
or U9896 (N_9896,N_9367,N_8770);
and U9897 (N_9897,N_9048,N_8892);
or U9898 (N_9898,N_8784,N_9126);
nor U9899 (N_9899,N_9161,N_8930);
and U9900 (N_9900,N_9010,N_9278);
or U9901 (N_9901,N_8835,N_9197);
xnor U9902 (N_9902,N_8855,N_9277);
nand U9903 (N_9903,N_9173,N_8830);
and U9904 (N_9904,N_9368,N_8792);
or U9905 (N_9905,N_8893,N_9185);
nor U9906 (N_9906,N_8841,N_9205);
or U9907 (N_9907,N_9214,N_9300);
nand U9908 (N_9908,N_8970,N_9104);
xor U9909 (N_9909,N_9371,N_9164);
and U9910 (N_9910,N_8815,N_9071);
and U9911 (N_9911,N_9208,N_8821);
nand U9912 (N_9912,N_9153,N_9041);
nor U9913 (N_9913,N_9247,N_9178);
nor U9914 (N_9914,N_9044,N_9101);
xor U9915 (N_9915,N_9259,N_8857);
nand U9916 (N_9916,N_9071,N_9231);
nor U9917 (N_9917,N_9035,N_9001);
xor U9918 (N_9918,N_8870,N_9192);
or U9919 (N_9919,N_9212,N_8958);
and U9920 (N_9920,N_9135,N_9245);
or U9921 (N_9921,N_9140,N_8975);
and U9922 (N_9922,N_8780,N_9339);
nand U9923 (N_9923,N_9196,N_8829);
nand U9924 (N_9924,N_9074,N_8925);
and U9925 (N_9925,N_8969,N_9177);
nor U9926 (N_9926,N_9075,N_9352);
xor U9927 (N_9927,N_8979,N_9150);
and U9928 (N_9928,N_9054,N_9309);
nor U9929 (N_9929,N_8829,N_8901);
xor U9930 (N_9930,N_9087,N_9264);
or U9931 (N_9931,N_9252,N_8952);
and U9932 (N_9932,N_9272,N_8869);
or U9933 (N_9933,N_8821,N_8987);
nand U9934 (N_9934,N_9237,N_9186);
nand U9935 (N_9935,N_9064,N_9141);
and U9936 (N_9936,N_9119,N_8808);
nor U9937 (N_9937,N_9082,N_9025);
nor U9938 (N_9938,N_9283,N_9314);
and U9939 (N_9939,N_9143,N_8917);
nor U9940 (N_9940,N_9259,N_9116);
xnor U9941 (N_9941,N_8759,N_8949);
nand U9942 (N_9942,N_8869,N_9012);
and U9943 (N_9943,N_9219,N_8825);
nor U9944 (N_9944,N_9034,N_9307);
xor U9945 (N_9945,N_9356,N_9371);
xnor U9946 (N_9946,N_8804,N_8987);
or U9947 (N_9947,N_9189,N_8892);
xnor U9948 (N_9948,N_9014,N_9015);
xor U9949 (N_9949,N_9304,N_8783);
nand U9950 (N_9950,N_9123,N_8996);
xor U9951 (N_9951,N_9202,N_9024);
nand U9952 (N_9952,N_8958,N_8822);
nand U9953 (N_9953,N_9354,N_9124);
and U9954 (N_9954,N_8998,N_9146);
or U9955 (N_9955,N_8805,N_9130);
nor U9956 (N_9956,N_9137,N_9243);
nand U9957 (N_9957,N_9316,N_8803);
nand U9958 (N_9958,N_9004,N_9222);
or U9959 (N_9959,N_9329,N_9067);
and U9960 (N_9960,N_9350,N_9016);
or U9961 (N_9961,N_8804,N_8800);
or U9962 (N_9962,N_8947,N_9346);
and U9963 (N_9963,N_9042,N_8981);
xor U9964 (N_9964,N_9254,N_9171);
and U9965 (N_9965,N_9332,N_9065);
nand U9966 (N_9966,N_9361,N_8782);
and U9967 (N_9967,N_9079,N_9039);
nor U9968 (N_9968,N_9055,N_9315);
xor U9969 (N_9969,N_8772,N_8921);
and U9970 (N_9970,N_9366,N_9231);
and U9971 (N_9971,N_9039,N_9121);
nand U9972 (N_9972,N_9343,N_8768);
xnor U9973 (N_9973,N_8794,N_9355);
xor U9974 (N_9974,N_9011,N_9038);
and U9975 (N_9975,N_9045,N_8957);
and U9976 (N_9976,N_8883,N_9082);
or U9977 (N_9977,N_8935,N_9167);
and U9978 (N_9978,N_9003,N_8766);
and U9979 (N_9979,N_9250,N_8984);
and U9980 (N_9980,N_9204,N_9290);
xnor U9981 (N_9981,N_9168,N_9264);
and U9982 (N_9982,N_8938,N_8770);
or U9983 (N_9983,N_9307,N_9139);
xnor U9984 (N_9984,N_8918,N_8971);
and U9985 (N_9985,N_8877,N_9112);
xor U9986 (N_9986,N_9303,N_8775);
nand U9987 (N_9987,N_9267,N_9309);
and U9988 (N_9988,N_8856,N_9336);
or U9989 (N_9989,N_9146,N_9368);
and U9990 (N_9990,N_8823,N_8864);
nand U9991 (N_9991,N_8864,N_8892);
nor U9992 (N_9992,N_8969,N_9184);
or U9993 (N_9993,N_9023,N_9333);
xnor U9994 (N_9994,N_9050,N_9334);
and U9995 (N_9995,N_8802,N_8969);
nand U9996 (N_9996,N_9126,N_8783);
and U9997 (N_9997,N_8881,N_9141);
and U9998 (N_9998,N_9182,N_8888);
nor U9999 (N_9999,N_8903,N_8966);
nand U10000 (N_10000,N_9896,N_9668);
nand U10001 (N_10001,N_9379,N_9616);
xor U10002 (N_10002,N_9509,N_9398);
nor U10003 (N_10003,N_9624,N_9642);
and U10004 (N_10004,N_9561,N_9549);
and U10005 (N_10005,N_9571,N_9590);
nor U10006 (N_10006,N_9575,N_9800);
and U10007 (N_10007,N_9512,N_9555);
and U10008 (N_10008,N_9482,N_9921);
nand U10009 (N_10009,N_9463,N_9834);
nand U10010 (N_10010,N_9399,N_9791);
nand U10011 (N_10011,N_9862,N_9598);
or U10012 (N_10012,N_9580,N_9576);
xor U10013 (N_10013,N_9637,N_9673);
and U10014 (N_10014,N_9694,N_9572);
xor U10015 (N_10015,N_9851,N_9931);
or U10016 (N_10016,N_9876,N_9559);
or U10017 (N_10017,N_9932,N_9538);
nor U10018 (N_10018,N_9454,N_9869);
xnor U10019 (N_10019,N_9383,N_9560);
and U10020 (N_10020,N_9607,N_9384);
xor U10021 (N_10021,N_9391,N_9567);
and U10022 (N_10022,N_9985,N_9669);
or U10023 (N_10023,N_9636,N_9606);
xor U10024 (N_10024,N_9734,N_9837);
xnor U10025 (N_10025,N_9836,N_9882);
or U10026 (N_10026,N_9536,N_9666);
xnor U10027 (N_10027,N_9845,N_9875);
or U10028 (N_10028,N_9486,N_9591);
and U10029 (N_10029,N_9718,N_9795);
nand U10030 (N_10030,N_9748,N_9543);
nor U10031 (N_10031,N_9641,N_9459);
xnor U10032 (N_10032,N_9422,N_9793);
and U10033 (N_10033,N_9650,N_9885);
xor U10034 (N_10034,N_9848,N_9900);
and U10035 (N_10035,N_9485,N_9674);
nor U10036 (N_10036,N_9530,N_9513);
or U10037 (N_10037,N_9424,N_9389);
or U10038 (N_10038,N_9617,N_9988);
or U10039 (N_10039,N_9393,N_9413);
or U10040 (N_10040,N_9553,N_9643);
nand U10041 (N_10041,N_9826,N_9473);
and U10042 (N_10042,N_9904,N_9649);
nor U10043 (N_10043,N_9647,N_9859);
and U10044 (N_10044,N_9770,N_9776);
and U10045 (N_10045,N_9947,N_9759);
or U10046 (N_10046,N_9442,N_9726);
or U10047 (N_10047,N_9462,N_9951);
nand U10048 (N_10048,N_9739,N_9983);
or U10049 (N_10049,N_9645,N_9550);
or U10050 (N_10050,N_9775,N_9631);
nand U10051 (N_10051,N_9919,N_9670);
nor U10052 (N_10052,N_9672,N_9764);
xor U10053 (N_10053,N_9527,N_9716);
nor U10054 (N_10054,N_9407,N_9618);
nor U10055 (N_10055,N_9972,N_9664);
xnor U10056 (N_10056,N_9994,N_9908);
xnor U10057 (N_10057,N_9853,N_9821);
and U10058 (N_10058,N_9788,N_9711);
and U10059 (N_10059,N_9426,N_9599);
xor U10060 (N_10060,N_9585,N_9749);
xor U10061 (N_10061,N_9717,N_9622);
nand U10062 (N_10062,N_9570,N_9778);
or U10063 (N_10063,N_9470,N_9743);
nand U10064 (N_10064,N_9756,N_9854);
xnor U10065 (N_10065,N_9644,N_9870);
and U10066 (N_10066,N_9843,N_9480);
and U10067 (N_10067,N_9533,N_9750);
nand U10068 (N_10068,N_9815,N_9989);
and U10069 (N_10069,N_9783,N_9547);
nor U10070 (N_10070,N_9879,N_9728);
or U10071 (N_10071,N_9472,N_9593);
or U10072 (N_10072,N_9765,N_9986);
and U10073 (N_10073,N_9600,N_9665);
nor U10074 (N_10074,N_9487,N_9823);
and U10075 (N_10075,N_9802,N_9944);
nor U10076 (N_10076,N_9754,N_9996);
nand U10077 (N_10077,N_9657,N_9918);
xor U10078 (N_10078,N_9628,N_9584);
or U10079 (N_10079,N_9496,N_9440);
xnor U10080 (N_10080,N_9762,N_9458);
or U10081 (N_10081,N_9898,N_9658);
xnor U10082 (N_10082,N_9605,N_9901);
nor U10083 (N_10083,N_9865,N_9639);
nor U10084 (N_10084,N_9774,N_9980);
xor U10085 (N_10085,N_9508,N_9707);
or U10086 (N_10086,N_9488,N_9781);
nor U10087 (N_10087,N_9796,N_9394);
nor U10088 (N_10088,N_9455,N_9970);
nor U10089 (N_10089,N_9518,N_9852);
xor U10090 (N_10090,N_9790,N_9903);
nor U10091 (N_10091,N_9629,N_9787);
nand U10092 (N_10092,N_9498,N_9648);
and U10093 (N_10093,N_9451,N_9615);
nand U10094 (N_10094,N_9706,N_9949);
xnor U10095 (N_10095,N_9577,N_9400);
or U10096 (N_10096,N_9722,N_9968);
nand U10097 (N_10097,N_9998,N_9625);
or U10098 (N_10098,N_9924,N_9514);
xor U10099 (N_10099,N_9871,N_9633);
and U10100 (N_10100,N_9652,N_9925);
nor U10101 (N_10101,N_9613,N_9840);
nor U10102 (N_10102,N_9830,N_9461);
and U10103 (N_10103,N_9943,N_9448);
xnor U10104 (N_10104,N_9727,N_9784);
xor U10105 (N_10105,N_9428,N_9566);
nor U10106 (N_10106,N_9757,N_9468);
nor U10107 (N_10107,N_9708,N_9952);
xor U10108 (N_10108,N_9376,N_9421);
xor U10109 (N_10109,N_9831,N_9506);
and U10110 (N_10110,N_9928,N_9477);
nor U10111 (N_10111,N_9945,N_9977);
or U10112 (N_10112,N_9827,N_9841);
or U10113 (N_10113,N_9655,N_9510);
or U10114 (N_10114,N_9634,N_9732);
xnor U10115 (N_10115,N_9915,N_9403);
nand U10116 (N_10116,N_9902,N_9456);
nand U10117 (N_10117,N_9752,N_9540);
nor U10118 (N_10118,N_9515,N_9965);
xnor U10119 (N_10119,N_9954,N_9948);
nor U10120 (N_10120,N_9627,N_9914);
and U10121 (N_10121,N_9844,N_9912);
and U10122 (N_10122,N_9742,N_9457);
xor U10123 (N_10123,N_9973,N_9883);
nand U10124 (N_10124,N_9683,N_9484);
nor U10125 (N_10125,N_9646,N_9856);
nor U10126 (N_10126,N_9849,N_9573);
nand U10127 (N_10127,N_9635,N_9967);
nor U10128 (N_10128,N_9934,N_9721);
and U10129 (N_10129,N_9444,N_9681);
or U10130 (N_10130,N_9773,N_9494);
and U10131 (N_10131,N_9433,N_9490);
and U10132 (N_10132,N_9659,N_9889);
xor U10133 (N_10133,N_9758,N_9528);
or U10134 (N_10134,N_9860,N_9699);
xor U10135 (N_10135,N_9493,N_9692);
xor U10136 (N_10136,N_9946,N_9897);
nor U10137 (N_10137,N_9378,N_9929);
nand U10138 (N_10138,N_9453,N_9660);
nor U10139 (N_10139,N_9464,N_9565);
nor U10140 (N_10140,N_9846,N_9736);
nor U10141 (N_10141,N_9961,N_9861);
xnor U10142 (N_10142,N_9890,N_9401);
and U10143 (N_10143,N_9704,N_9390);
or U10144 (N_10144,N_9703,N_9723);
nor U10145 (N_10145,N_9430,N_9630);
nand U10146 (N_10146,N_9663,N_9839);
or U10147 (N_10147,N_9991,N_9387);
xor U10148 (N_10148,N_9475,N_9963);
or U10149 (N_10149,N_9857,N_9735);
nor U10150 (N_10150,N_9942,N_9971);
nor U10151 (N_10151,N_9698,N_9608);
nand U10152 (N_10152,N_9385,N_9935);
nand U10153 (N_10153,N_9640,N_9632);
or U10154 (N_10154,N_9701,N_9638);
nand U10155 (N_10155,N_9911,N_9917);
xnor U10156 (N_10156,N_9738,N_9503);
nand U10157 (N_10157,N_9953,N_9812);
nor U10158 (N_10158,N_9907,N_9786);
xor U10159 (N_10159,N_9667,N_9691);
or U10160 (N_10160,N_9539,N_9810);
nand U10161 (N_10161,N_9588,N_9481);
xnor U10162 (N_10162,N_9469,N_9891);
nand U10163 (N_10163,N_9411,N_9892);
and U10164 (N_10164,N_9842,N_9868);
or U10165 (N_10165,N_9610,N_9397);
and U10166 (N_10166,N_9557,N_9386);
nor U10167 (N_10167,N_9502,N_9858);
xor U10168 (N_10168,N_9792,N_9777);
and U10169 (N_10169,N_9425,N_9979);
nor U10170 (N_10170,N_9589,N_9656);
xnor U10171 (N_10171,N_9766,N_9417);
and U10172 (N_10172,N_9677,N_9689);
or U10173 (N_10173,N_9850,N_9808);
xnor U10174 (N_10174,N_9554,N_9782);
and U10175 (N_10175,N_9761,N_9381);
and U10176 (N_10176,N_9855,N_9684);
nand U10177 (N_10177,N_9519,N_9926);
nor U10178 (N_10178,N_9495,N_9807);
and U10179 (N_10179,N_9612,N_9964);
xor U10180 (N_10180,N_9730,N_9438);
or U10181 (N_10181,N_9789,N_9930);
or U10182 (N_10182,N_9910,N_9419);
nand U10183 (N_10183,N_9937,N_9679);
xnor U10184 (N_10184,N_9872,N_9818);
nor U10185 (N_10185,N_9969,N_9603);
and U10186 (N_10186,N_9497,N_9601);
and U10187 (N_10187,N_9479,N_9466);
nand U10188 (N_10188,N_9609,N_9450);
nor U10189 (N_10189,N_9471,N_9940);
or U10190 (N_10190,N_9886,N_9895);
or U10191 (N_10191,N_9729,N_9418);
nor U10192 (N_10192,N_9753,N_9975);
nand U10193 (N_10193,N_9820,N_9751);
nand U10194 (N_10194,N_9534,N_9710);
xnor U10195 (N_10195,N_9696,N_9906);
nand U10196 (N_10196,N_9941,N_9806);
nand U10197 (N_10197,N_9956,N_9824);
or U10198 (N_10198,N_9874,N_9720);
nand U10199 (N_10199,N_9755,N_9920);
nor U10200 (N_10200,N_9744,N_9432);
and U10201 (N_10201,N_9709,N_9873);
nor U10202 (N_10202,N_9877,N_9501);
nor U10203 (N_10203,N_9564,N_9864);
nor U10204 (N_10204,N_9409,N_9913);
and U10205 (N_10205,N_9867,N_9478);
nor U10206 (N_10206,N_9825,N_9582);
and U10207 (N_10207,N_9491,N_9529);
and U10208 (N_10208,N_9548,N_9719);
or U10209 (N_10209,N_9435,N_9661);
xnor U10210 (N_10210,N_9724,N_9596);
nor U10211 (N_10211,N_9811,N_9995);
and U10212 (N_10212,N_9939,N_9653);
and U10213 (N_10213,N_9686,N_9768);
nor U10214 (N_10214,N_9887,N_9654);
and U10215 (N_10215,N_9936,N_9675);
or U10216 (N_10216,N_9705,N_9923);
or U10217 (N_10217,N_9556,N_9741);
or U10218 (N_10218,N_9521,N_9447);
nor U10219 (N_10219,N_9410,N_9552);
nor U10220 (N_10220,N_9962,N_9798);
and U10221 (N_10221,N_9767,N_9715);
nor U10222 (N_10222,N_9712,N_9938);
and U10223 (N_10223,N_9797,N_9416);
or U10224 (N_10224,N_9382,N_9687);
nand U10225 (N_10225,N_9933,N_9388);
and U10226 (N_10226,N_9429,N_9760);
nor U10227 (N_10227,N_9993,N_9747);
and U10228 (N_10228,N_9863,N_9794);
and U10229 (N_10229,N_9955,N_9779);
or U10230 (N_10230,N_9884,N_9958);
nor U10231 (N_10231,N_9982,N_9511);
and U10232 (N_10232,N_9532,N_9909);
nand U10233 (N_10233,N_9651,N_9568);
or U10234 (N_10234,N_9916,N_9922);
and U10235 (N_10235,N_9500,N_9523);
xor U10236 (N_10236,N_9813,N_9545);
xor U10237 (N_10237,N_9981,N_9733);
and U10238 (N_10238,N_9544,N_9682);
nand U10239 (N_10239,N_9434,N_9449);
and U10240 (N_10240,N_9888,N_9404);
and U10241 (N_10241,N_9678,N_9894);
and U10242 (N_10242,N_9829,N_9780);
or U10243 (N_10243,N_9396,N_9838);
xnor U10244 (N_10244,N_9423,N_9406);
nor U10245 (N_10245,N_9427,N_9412);
nand U10246 (N_10246,N_9804,N_9621);
nor U10247 (N_10247,N_9763,N_9392);
and U10248 (N_10248,N_9693,N_9586);
or U10249 (N_10249,N_9822,N_9990);
and U10250 (N_10250,N_9697,N_9563);
and U10251 (N_10251,N_9581,N_9460);
nand U10252 (N_10252,N_9662,N_9866);
nor U10253 (N_10253,N_9504,N_9602);
or U10254 (N_10254,N_9893,N_9992);
nor U10255 (N_10255,N_9524,N_9526);
xnor U10256 (N_10256,N_9769,N_9878);
nor U10257 (N_10257,N_9452,N_9620);
xor U10258 (N_10258,N_9832,N_9835);
and U10259 (N_10259,N_9695,N_9987);
xor U10260 (N_10260,N_9950,N_9405);
xnor U10261 (N_10261,N_9611,N_9772);
xor U10262 (N_10262,N_9551,N_9420);
and U10263 (N_10263,N_9999,N_9505);
xnor U10264 (N_10264,N_9492,N_9437);
nand U10265 (N_10265,N_9623,N_9467);
nor U10266 (N_10266,N_9680,N_9771);
nor U10267 (N_10267,N_9436,N_9960);
xnor U10268 (N_10268,N_9619,N_9542);
and U10269 (N_10269,N_9803,N_9997);
xnor U10270 (N_10270,N_9489,N_9959);
xor U10271 (N_10271,N_9880,N_9522);
or U10272 (N_10272,N_9562,N_9441);
nand U10273 (N_10273,N_9745,N_9688);
xor U10274 (N_10274,N_9395,N_9507);
or U10275 (N_10275,N_9966,N_9690);
xor U10276 (N_10276,N_9905,N_9685);
nor U10277 (N_10277,N_9833,N_9525);
nor U10278 (N_10278,N_9408,N_9814);
and U10279 (N_10279,N_9414,N_9558);
or U10280 (N_10280,N_9671,N_9520);
nor U10281 (N_10281,N_9537,N_9978);
nor U10282 (N_10282,N_9819,N_9574);
nand U10283 (N_10283,N_9626,N_9439);
xnor U10284 (N_10284,N_9546,N_9476);
nor U10285 (N_10285,N_9579,N_9377);
and U10286 (N_10286,N_9809,N_9592);
nand U10287 (N_10287,N_9737,N_9583);
xor U10288 (N_10288,N_9785,N_9614);
or U10289 (N_10289,N_9531,N_9740);
nand U10290 (N_10290,N_9380,N_9847);
nor U10291 (N_10291,N_9474,N_9445);
nor U10292 (N_10292,N_9597,N_9974);
xnor U10293 (N_10293,N_9899,N_9587);
nor U10294 (N_10294,N_9700,N_9927);
nand U10295 (N_10295,N_9483,N_9569);
nor U10296 (N_10296,N_9516,N_9443);
and U10297 (N_10297,N_9578,N_9881);
xnor U10298 (N_10298,N_9517,N_9957);
nor U10299 (N_10299,N_9446,N_9828);
and U10300 (N_10300,N_9676,N_9799);
xor U10301 (N_10301,N_9984,N_9801);
nand U10302 (N_10302,N_9725,N_9499);
and U10303 (N_10303,N_9746,N_9731);
or U10304 (N_10304,N_9594,N_9714);
nand U10305 (N_10305,N_9535,N_9415);
nand U10306 (N_10306,N_9702,N_9541);
nor U10307 (N_10307,N_9816,N_9402);
nand U10308 (N_10308,N_9604,N_9817);
xor U10309 (N_10309,N_9431,N_9465);
and U10310 (N_10310,N_9713,N_9375);
or U10311 (N_10311,N_9976,N_9595);
nor U10312 (N_10312,N_9805,N_9462);
xnor U10313 (N_10313,N_9655,N_9692);
or U10314 (N_10314,N_9783,N_9809);
and U10315 (N_10315,N_9801,N_9884);
and U10316 (N_10316,N_9847,N_9440);
xnor U10317 (N_10317,N_9766,N_9714);
or U10318 (N_10318,N_9781,N_9552);
nor U10319 (N_10319,N_9985,N_9670);
nand U10320 (N_10320,N_9670,N_9731);
xor U10321 (N_10321,N_9705,N_9819);
xor U10322 (N_10322,N_9485,N_9823);
xnor U10323 (N_10323,N_9744,N_9992);
nand U10324 (N_10324,N_9542,N_9496);
or U10325 (N_10325,N_9792,N_9490);
and U10326 (N_10326,N_9460,N_9787);
nor U10327 (N_10327,N_9707,N_9935);
or U10328 (N_10328,N_9383,N_9397);
nor U10329 (N_10329,N_9806,N_9872);
or U10330 (N_10330,N_9421,N_9842);
or U10331 (N_10331,N_9378,N_9708);
or U10332 (N_10332,N_9744,N_9476);
nor U10333 (N_10333,N_9617,N_9618);
or U10334 (N_10334,N_9588,N_9865);
nand U10335 (N_10335,N_9498,N_9861);
nand U10336 (N_10336,N_9915,N_9896);
nand U10337 (N_10337,N_9567,N_9752);
xor U10338 (N_10338,N_9644,N_9382);
or U10339 (N_10339,N_9757,N_9886);
or U10340 (N_10340,N_9691,N_9954);
or U10341 (N_10341,N_9411,N_9989);
and U10342 (N_10342,N_9683,N_9704);
and U10343 (N_10343,N_9878,N_9724);
nand U10344 (N_10344,N_9388,N_9919);
nor U10345 (N_10345,N_9398,N_9638);
xor U10346 (N_10346,N_9877,N_9783);
or U10347 (N_10347,N_9429,N_9569);
xnor U10348 (N_10348,N_9818,N_9715);
nand U10349 (N_10349,N_9952,N_9953);
or U10350 (N_10350,N_9640,N_9526);
or U10351 (N_10351,N_9781,N_9711);
and U10352 (N_10352,N_9880,N_9599);
and U10353 (N_10353,N_9740,N_9495);
xor U10354 (N_10354,N_9644,N_9485);
or U10355 (N_10355,N_9853,N_9763);
or U10356 (N_10356,N_9523,N_9564);
xnor U10357 (N_10357,N_9380,N_9917);
xor U10358 (N_10358,N_9789,N_9673);
nand U10359 (N_10359,N_9729,N_9644);
or U10360 (N_10360,N_9925,N_9681);
nor U10361 (N_10361,N_9593,N_9984);
or U10362 (N_10362,N_9620,N_9644);
nand U10363 (N_10363,N_9829,N_9987);
xnor U10364 (N_10364,N_9606,N_9776);
nor U10365 (N_10365,N_9378,N_9844);
or U10366 (N_10366,N_9926,N_9848);
nor U10367 (N_10367,N_9918,N_9988);
xnor U10368 (N_10368,N_9791,N_9902);
and U10369 (N_10369,N_9470,N_9457);
or U10370 (N_10370,N_9481,N_9820);
nand U10371 (N_10371,N_9418,N_9682);
nand U10372 (N_10372,N_9861,N_9765);
xor U10373 (N_10373,N_9563,N_9667);
nand U10374 (N_10374,N_9540,N_9542);
nor U10375 (N_10375,N_9741,N_9444);
and U10376 (N_10376,N_9691,N_9749);
xnor U10377 (N_10377,N_9962,N_9828);
xnor U10378 (N_10378,N_9872,N_9946);
nor U10379 (N_10379,N_9558,N_9933);
xor U10380 (N_10380,N_9841,N_9917);
and U10381 (N_10381,N_9774,N_9463);
or U10382 (N_10382,N_9608,N_9533);
or U10383 (N_10383,N_9768,N_9557);
xnor U10384 (N_10384,N_9739,N_9718);
nor U10385 (N_10385,N_9688,N_9643);
and U10386 (N_10386,N_9832,N_9739);
or U10387 (N_10387,N_9809,N_9620);
xor U10388 (N_10388,N_9645,N_9983);
nor U10389 (N_10389,N_9727,N_9950);
nand U10390 (N_10390,N_9876,N_9512);
nor U10391 (N_10391,N_9450,N_9386);
xnor U10392 (N_10392,N_9421,N_9978);
and U10393 (N_10393,N_9600,N_9431);
or U10394 (N_10394,N_9880,N_9851);
nor U10395 (N_10395,N_9663,N_9423);
nand U10396 (N_10396,N_9654,N_9740);
nor U10397 (N_10397,N_9536,N_9903);
nor U10398 (N_10398,N_9462,N_9537);
or U10399 (N_10399,N_9862,N_9767);
and U10400 (N_10400,N_9677,N_9833);
nor U10401 (N_10401,N_9787,N_9674);
nor U10402 (N_10402,N_9534,N_9963);
xor U10403 (N_10403,N_9948,N_9812);
or U10404 (N_10404,N_9595,N_9701);
xor U10405 (N_10405,N_9893,N_9716);
xnor U10406 (N_10406,N_9405,N_9627);
xor U10407 (N_10407,N_9600,N_9953);
or U10408 (N_10408,N_9641,N_9476);
nor U10409 (N_10409,N_9994,N_9852);
nor U10410 (N_10410,N_9795,N_9425);
nand U10411 (N_10411,N_9937,N_9710);
nand U10412 (N_10412,N_9923,N_9580);
nor U10413 (N_10413,N_9758,N_9444);
nand U10414 (N_10414,N_9783,N_9471);
and U10415 (N_10415,N_9663,N_9416);
xnor U10416 (N_10416,N_9618,N_9468);
xor U10417 (N_10417,N_9459,N_9802);
and U10418 (N_10418,N_9814,N_9738);
xnor U10419 (N_10419,N_9897,N_9865);
and U10420 (N_10420,N_9889,N_9938);
nor U10421 (N_10421,N_9506,N_9576);
and U10422 (N_10422,N_9409,N_9659);
xnor U10423 (N_10423,N_9960,N_9792);
nand U10424 (N_10424,N_9833,N_9756);
xnor U10425 (N_10425,N_9694,N_9987);
nor U10426 (N_10426,N_9912,N_9930);
xnor U10427 (N_10427,N_9384,N_9596);
nand U10428 (N_10428,N_9400,N_9387);
nor U10429 (N_10429,N_9484,N_9797);
nor U10430 (N_10430,N_9907,N_9808);
nand U10431 (N_10431,N_9379,N_9669);
and U10432 (N_10432,N_9920,N_9880);
nor U10433 (N_10433,N_9992,N_9715);
xor U10434 (N_10434,N_9636,N_9951);
and U10435 (N_10435,N_9890,N_9860);
and U10436 (N_10436,N_9413,N_9646);
and U10437 (N_10437,N_9463,N_9375);
nor U10438 (N_10438,N_9399,N_9469);
nand U10439 (N_10439,N_9658,N_9848);
and U10440 (N_10440,N_9726,N_9810);
or U10441 (N_10441,N_9814,N_9507);
or U10442 (N_10442,N_9734,N_9959);
nand U10443 (N_10443,N_9726,N_9438);
xor U10444 (N_10444,N_9985,N_9931);
xor U10445 (N_10445,N_9942,N_9970);
nor U10446 (N_10446,N_9892,N_9757);
or U10447 (N_10447,N_9621,N_9815);
nand U10448 (N_10448,N_9582,N_9427);
nor U10449 (N_10449,N_9790,N_9456);
or U10450 (N_10450,N_9596,N_9914);
nor U10451 (N_10451,N_9967,N_9864);
nand U10452 (N_10452,N_9524,N_9463);
nor U10453 (N_10453,N_9463,N_9694);
or U10454 (N_10454,N_9510,N_9413);
xnor U10455 (N_10455,N_9453,N_9947);
nor U10456 (N_10456,N_9769,N_9591);
nor U10457 (N_10457,N_9852,N_9752);
nand U10458 (N_10458,N_9430,N_9418);
nor U10459 (N_10459,N_9918,N_9675);
or U10460 (N_10460,N_9759,N_9499);
and U10461 (N_10461,N_9729,N_9690);
nor U10462 (N_10462,N_9697,N_9539);
xnor U10463 (N_10463,N_9997,N_9410);
nor U10464 (N_10464,N_9871,N_9899);
xnor U10465 (N_10465,N_9427,N_9819);
nand U10466 (N_10466,N_9651,N_9386);
or U10467 (N_10467,N_9767,N_9965);
nor U10468 (N_10468,N_9508,N_9556);
xor U10469 (N_10469,N_9593,N_9632);
nor U10470 (N_10470,N_9995,N_9941);
nand U10471 (N_10471,N_9600,N_9823);
xnor U10472 (N_10472,N_9586,N_9955);
and U10473 (N_10473,N_9990,N_9810);
or U10474 (N_10474,N_9402,N_9549);
or U10475 (N_10475,N_9755,N_9567);
or U10476 (N_10476,N_9490,N_9700);
and U10477 (N_10477,N_9576,N_9549);
and U10478 (N_10478,N_9883,N_9468);
xnor U10479 (N_10479,N_9426,N_9508);
or U10480 (N_10480,N_9888,N_9433);
nand U10481 (N_10481,N_9688,N_9932);
and U10482 (N_10482,N_9604,N_9957);
or U10483 (N_10483,N_9419,N_9660);
xor U10484 (N_10484,N_9689,N_9567);
nor U10485 (N_10485,N_9851,N_9955);
xor U10486 (N_10486,N_9830,N_9892);
xnor U10487 (N_10487,N_9677,N_9728);
nor U10488 (N_10488,N_9703,N_9638);
nor U10489 (N_10489,N_9461,N_9451);
or U10490 (N_10490,N_9434,N_9421);
or U10491 (N_10491,N_9920,N_9844);
nand U10492 (N_10492,N_9712,N_9385);
and U10493 (N_10493,N_9667,N_9499);
nand U10494 (N_10494,N_9901,N_9923);
nor U10495 (N_10495,N_9650,N_9503);
xnor U10496 (N_10496,N_9820,N_9666);
and U10497 (N_10497,N_9733,N_9796);
and U10498 (N_10498,N_9864,N_9712);
nor U10499 (N_10499,N_9686,N_9965);
and U10500 (N_10500,N_9723,N_9509);
nor U10501 (N_10501,N_9674,N_9574);
xor U10502 (N_10502,N_9554,N_9879);
nor U10503 (N_10503,N_9622,N_9694);
nor U10504 (N_10504,N_9887,N_9399);
nor U10505 (N_10505,N_9705,N_9873);
nor U10506 (N_10506,N_9837,N_9676);
nor U10507 (N_10507,N_9941,N_9979);
nor U10508 (N_10508,N_9584,N_9409);
or U10509 (N_10509,N_9992,N_9475);
xor U10510 (N_10510,N_9970,N_9622);
or U10511 (N_10511,N_9538,N_9955);
nor U10512 (N_10512,N_9814,N_9820);
nor U10513 (N_10513,N_9747,N_9977);
or U10514 (N_10514,N_9514,N_9511);
or U10515 (N_10515,N_9406,N_9493);
and U10516 (N_10516,N_9626,N_9841);
or U10517 (N_10517,N_9795,N_9443);
nor U10518 (N_10518,N_9562,N_9663);
or U10519 (N_10519,N_9527,N_9918);
nand U10520 (N_10520,N_9629,N_9617);
and U10521 (N_10521,N_9888,N_9737);
and U10522 (N_10522,N_9823,N_9409);
and U10523 (N_10523,N_9436,N_9675);
or U10524 (N_10524,N_9445,N_9844);
and U10525 (N_10525,N_9594,N_9608);
and U10526 (N_10526,N_9426,N_9913);
nor U10527 (N_10527,N_9734,N_9468);
nor U10528 (N_10528,N_9934,N_9981);
xnor U10529 (N_10529,N_9594,N_9784);
nor U10530 (N_10530,N_9929,N_9985);
xnor U10531 (N_10531,N_9383,N_9481);
or U10532 (N_10532,N_9628,N_9456);
nor U10533 (N_10533,N_9595,N_9506);
and U10534 (N_10534,N_9498,N_9807);
xor U10535 (N_10535,N_9759,N_9654);
or U10536 (N_10536,N_9508,N_9735);
and U10537 (N_10537,N_9848,N_9790);
nand U10538 (N_10538,N_9621,N_9578);
nor U10539 (N_10539,N_9622,N_9759);
or U10540 (N_10540,N_9459,N_9774);
nand U10541 (N_10541,N_9392,N_9593);
and U10542 (N_10542,N_9874,N_9562);
or U10543 (N_10543,N_9795,N_9851);
and U10544 (N_10544,N_9872,N_9534);
or U10545 (N_10545,N_9719,N_9653);
nand U10546 (N_10546,N_9400,N_9947);
nand U10547 (N_10547,N_9414,N_9937);
nand U10548 (N_10548,N_9933,N_9755);
nor U10549 (N_10549,N_9753,N_9790);
nor U10550 (N_10550,N_9872,N_9391);
xnor U10551 (N_10551,N_9856,N_9586);
and U10552 (N_10552,N_9822,N_9411);
and U10553 (N_10553,N_9919,N_9404);
nand U10554 (N_10554,N_9410,N_9719);
and U10555 (N_10555,N_9645,N_9969);
nand U10556 (N_10556,N_9476,N_9612);
xnor U10557 (N_10557,N_9387,N_9624);
nand U10558 (N_10558,N_9671,N_9889);
or U10559 (N_10559,N_9461,N_9430);
xnor U10560 (N_10560,N_9609,N_9582);
and U10561 (N_10561,N_9627,N_9697);
and U10562 (N_10562,N_9970,N_9956);
or U10563 (N_10563,N_9675,N_9378);
xnor U10564 (N_10564,N_9515,N_9572);
or U10565 (N_10565,N_9586,N_9656);
nand U10566 (N_10566,N_9806,N_9416);
nor U10567 (N_10567,N_9454,N_9818);
nor U10568 (N_10568,N_9808,N_9945);
and U10569 (N_10569,N_9577,N_9517);
nand U10570 (N_10570,N_9559,N_9478);
and U10571 (N_10571,N_9564,N_9854);
xnor U10572 (N_10572,N_9636,N_9968);
or U10573 (N_10573,N_9522,N_9441);
nor U10574 (N_10574,N_9390,N_9437);
nor U10575 (N_10575,N_9907,N_9677);
nor U10576 (N_10576,N_9766,N_9954);
nor U10577 (N_10577,N_9394,N_9451);
and U10578 (N_10578,N_9712,N_9631);
nand U10579 (N_10579,N_9799,N_9508);
or U10580 (N_10580,N_9767,N_9723);
or U10581 (N_10581,N_9897,N_9487);
xnor U10582 (N_10582,N_9644,N_9683);
xor U10583 (N_10583,N_9944,N_9546);
xor U10584 (N_10584,N_9675,N_9610);
nor U10585 (N_10585,N_9554,N_9816);
xnor U10586 (N_10586,N_9393,N_9983);
and U10587 (N_10587,N_9645,N_9584);
and U10588 (N_10588,N_9502,N_9687);
xnor U10589 (N_10589,N_9599,N_9392);
nand U10590 (N_10590,N_9613,N_9832);
nand U10591 (N_10591,N_9482,N_9853);
nor U10592 (N_10592,N_9899,N_9836);
xor U10593 (N_10593,N_9719,N_9880);
or U10594 (N_10594,N_9740,N_9587);
nor U10595 (N_10595,N_9664,N_9880);
nand U10596 (N_10596,N_9696,N_9580);
xor U10597 (N_10597,N_9847,N_9596);
and U10598 (N_10598,N_9615,N_9976);
xor U10599 (N_10599,N_9754,N_9768);
and U10600 (N_10600,N_9802,N_9963);
or U10601 (N_10601,N_9470,N_9477);
xor U10602 (N_10602,N_9585,N_9781);
nand U10603 (N_10603,N_9852,N_9652);
or U10604 (N_10604,N_9422,N_9555);
and U10605 (N_10605,N_9488,N_9676);
or U10606 (N_10606,N_9921,N_9966);
nand U10607 (N_10607,N_9739,N_9411);
or U10608 (N_10608,N_9622,N_9650);
nor U10609 (N_10609,N_9792,N_9935);
nand U10610 (N_10610,N_9737,N_9504);
xnor U10611 (N_10611,N_9799,N_9644);
and U10612 (N_10612,N_9718,N_9443);
or U10613 (N_10613,N_9700,N_9894);
and U10614 (N_10614,N_9781,N_9864);
nand U10615 (N_10615,N_9482,N_9591);
xnor U10616 (N_10616,N_9389,N_9806);
and U10617 (N_10617,N_9867,N_9760);
or U10618 (N_10618,N_9504,N_9533);
and U10619 (N_10619,N_9758,N_9624);
xnor U10620 (N_10620,N_9438,N_9517);
or U10621 (N_10621,N_9891,N_9814);
nor U10622 (N_10622,N_9806,N_9796);
or U10623 (N_10623,N_9749,N_9740);
or U10624 (N_10624,N_9701,N_9452);
and U10625 (N_10625,N_10527,N_10304);
nor U10626 (N_10626,N_10158,N_10481);
nor U10627 (N_10627,N_10538,N_10343);
nand U10628 (N_10628,N_10111,N_10502);
nand U10629 (N_10629,N_10194,N_10484);
xor U10630 (N_10630,N_10071,N_10623);
or U10631 (N_10631,N_10025,N_10317);
nand U10632 (N_10632,N_10178,N_10309);
nand U10633 (N_10633,N_10516,N_10499);
nand U10634 (N_10634,N_10351,N_10588);
xor U10635 (N_10635,N_10551,N_10413);
xnor U10636 (N_10636,N_10471,N_10555);
nand U10637 (N_10637,N_10344,N_10063);
nand U10638 (N_10638,N_10609,N_10357);
or U10639 (N_10639,N_10140,N_10453);
and U10640 (N_10640,N_10302,N_10314);
nor U10641 (N_10641,N_10321,N_10611);
nand U10642 (N_10642,N_10569,N_10521);
nor U10643 (N_10643,N_10531,N_10590);
nor U10644 (N_10644,N_10434,N_10168);
nor U10645 (N_10645,N_10115,N_10230);
xor U10646 (N_10646,N_10361,N_10599);
xor U10647 (N_10647,N_10188,N_10038);
nor U10648 (N_10648,N_10595,N_10187);
nor U10649 (N_10649,N_10301,N_10450);
nor U10650 (N_10650,N_10445,N_10152);
xor U10651 (N_10651,N_10478,N_10050);
nor U10652 (N_10652,N_10005,N_10269);
and U10653 (N_10653,N_10475,N_10232);
and U10654 (N_10654,N_10393,N_10617);
and U10655 (N_10655,N_10579,N_10205);
or U10656 (N_10656,N_10089,N_10616);
and U10657 (N_10657,N_10094,N_10044);
and U10658 (N_10658,N_10160,N_10104);
nor U10659 (N_10659,N_10003,N_10435);
nand U10660 (N_10660,N_10030,N_10244);
nor U10661 (N_10661,N_10219,N_10171);
and U10662 (N_10662,N_10510,N_10184);
and U10663 (N_10663,N_10008,N_10574);
and U10664 (N_10664,N_10437,N_10455);
and U10665 (N_10665,N_10325,N_10054);
nor U10666 (N_10666,N_10567,N_10525);
nor U10667 (N_10667,N_10618,N_10074);
and U10668 (N_10668,N_10007,N_10523);
xnor U10669 (N_10669,N_10572,N_10466);
or U10670 (N_10670,N_10259,N_10347);
nor U10671 (N_10671,N_10322,N_10249);
or U10672 (N_10672,N_10452,N_10355);
or U10673 (N_10673,N_10059,N_10253);
or U10674 (N_10674,N_10068,N_10203);
nand U10675 (N_10675,N_10556,N_10091);
and U10676 (N_10676,N_10405,N_10048);
nor U10677 (N_10677,N_10429,N_10065);
or U10678 (N_10678,N_10053,N_10324);
and U10679 (N_10679,N_10067,N_10486);
and U10680 (N_10680,N_10315,N_10418);
xor U10681 (N_10681,N_10487,N_10045);
nand U10682 (N_10682,N_10051,N_10542);
xnor U10683 (N_10683,N_10147,N_10124);
or U10684 (N_10684,N_10472,N_10133);
xor U10685 (N_10685,N_10083,N_10155);
nand U10686 (N_10686,N_10606,N_10423);
and U10687 (N_10687,N_10440,N_10144);
and U10688 (N_10688,N_10087,N_10143);
nor U10689 (N_10689,N_10229,N_10207);
and U10690 (N_10690,N_10526,N_10024);
and U10691 (N_10691,N_10163,N_10040);
and U10692 (N_10692,N_10585,N_10081);
xor U10693 (N_10693,N_10076,N_10305);
and U10694 (N_10694,N_10243,N_10577);
xor U10695 (N_10695,N_10443,N_10340);
and U10696 (N_10696,N_10345,N_10061);
and U10697 (N_10697,N_10278,N_10080);
nand U10698 (N_10698,N_10389,N_10075);
or U10699 (N_10699,N_10513,N_10564);
nor U10700 (N_10700,N_10239,N_10159);
nand U10701 (N_10701,N_10385,N_10032);
and U10702 (N_10702,N_10589,N_10265);
and U10703 (N_10703,N_10284,N_10494);
and U10704 (N_10704,N_10565,N_10594);
nand U10705 (N_10705,N_10198,N_10339);
and U10706 (N_10706,N_10619,N_10079);
nor U10707 (N_10707,N_10607,N_10135);
or U10708 (N_10708,N_10615,N_10404);
or U10709 (N_10709,N_10377,N_10409);
nor U10710 (N_10710,N_10245,N_10281);
and U10711 (N_10711,N_10467,N_10150);
nand U10712 (N_10712,N_10603,N_10110);
nand U10713 (N_10713,N_10495,N_10134);
or U10714 (N_10714,N_10319,N_10234);
nor U10715 (N_10715,N_10098,N_10123);
nand U10716 (N_10716,N_10575,N_10221);
or U10717 (N_10717,N_10532,N_10073);
and U10718 (N_10718,N_10493,N_10167);
nand U10719 (N_10719,N_10154,N_10388);
xnor U10720 (N_10720,N_10566,N_10557);
or U10721 (N_10721,N_10403,N_10242);
nor U10722 (N_10722,N_10176,N_10216);
xnor U10723 (N_10723,N_10046,N_10316);
nor U10724 (N_10724,N_10483,N_10199);
nor U10725 (N_10725,N_10515,N_10360);
nand U10726 (N_10726,N_10506,N_10563);
or U10727 (N_10727,N_10451,N_10534);
xnor U10728 (N_10728,N_10283,N_10420);
and U10729 (N_10729,N_10113,N_10109);
and U10730 (N_10730,N_10456,N_10069);
nand U10731 (N_10731,N_10421,N_10027);
and U10732 (N_10732,N_10224,N_10191);
or U10733 (N_10733,N_10262,N_10307);
nor U10734 (N_10734,N_10454,N_10218);
xnor U10735 (N_10735,N_10006,N_10601);
and U10736 (N_10736,N_10238,N_10255);
xor U10737 (N_10737,N_10492,N_10220);
xor U10738 (N_10738,N_10128,N_10449);
nand U10739 (N_10739,N_10227,N_10333);
xnor U10740 (N_10740,N_10479,N_10318);
and U10741 (N_10741,N_10415,N_10398);
nor U10742 (N_10742,N_10544,N_10392);
nor U10743 (N_10743,N_10182,N_10547);
and U10744 (N_10744,N_10039,N_10252);
and U10745 (N_10745,N_10596,N_10504);
and U10746 (N_10746,N_10015,N_10460);
xor U10747 (N_10747,N_10384,N_10356);
and U10748 (N_10748,N_10583,N_10272);
or U10749 (N_10749,N_10280,N_10062);
nand U10750 (N_10750,N_10179,N_10605);
and U10751 (N_10751,N_10204,N_10228);
nor U10752 (N_10752,N_10173,N_10029);
and U10753 (N_10753,N_10518,N_10349);
nand U10754 (N_10754,N_10480,N_10426);
or U10755 (N_10755,N_10086,N_10078);
xor U10756 (N_10756,N_10241,N_10608);
and U10757 (N_10757,N_10573,N_10406);
or U10758 (N_10758,N_10622,N_10041);
xnor U10759 (N_10759,N_10141,N_10267);
xor U10760 (N_10760,N_10208,N_10247);
nand U10761 (N_10761,N_10240,N_10107);
nor U10762 (N_10762,N_10522,N_10470);
nand U10763 (N_10763,N_10391,N_10335);
xor U10764 (N_10764,N_10034,N_10275);
nor U10765 (N_10765,N_10503,N_10162);
and U10766 (N_10766,N_10186,N_10164);
nor U10767 (N_10767,N_10190,N_10584);
nand U10768 (N_10768,N_10058,N_10568);
and U10769 (N_10769,N_10468,N_10130);
or U10770 (N_10770,N_10175,N_10258);
xor U10771 (N_10771,N_10047,N_10352);
nor U10772 (N_10772,N_10326,N_10271);
xnor U10773 (N_10773,N_10180,N_10019);
nor U10774 (N_10774,N_10055,N_10085);
xnor U10775 (N_10775,N_10358,N_10399);
and U10776 (N_10776,N_10233,N_10310);
xnor U10777 (N_10777,N_10016,N_10524);
xnor U10778 (N_10778,N_10461,N_10095);
xor U10779 (N_10779,N_10463,N_10490);
nor U10780 (N_10780,N_10411,N_10052);
and U10781 (N_10781,N_10174,N_10586);
and U10782 (N_10782,N_10436,N_10397);
xnor U10783 (N_10783,N_10250,N_10291);
nor U10784 (N_10784,N_10549,N_10323);
and U10785 (N_10785,N_10482,N_10552);
nor U10786 (N_10786,N_10328,N_10211);
or U10787 (N_10787,N_10402,N_10498);
xor U10788 (N_10788,N_10410,N_10013);
nor U10789 (N_10789,N_10311,N_10395);
nand U10790 (N_10790,N_10320,N_10161);
nor U10791 (N_10791,N_10373,N_10380);
and U10792 (N_10792,N_10306,N_10332);
and U10793 (N_10793,N_10587,N_10139);
or U10794 (N_10794,N_10066,N_10612);
or U10795 (N_10795,N_10541,N_10501);
nor U10796 (N_10796,N_10296,N_10096);
nand U10797 (N_10797,N_10294,N_10172);
nand U10798 (N_10798,N_10474,N_10331);
nor U10799 (N_10799,N_10313,N_10558);
nand U10800 (N_10800,N_10235,N_10394);
nand U10801 (N_10801,N_10185,N_10386);
and U10802 (N_10802,N_10485,N_10097);
and U10803 (N_10803,N_10424,N_10497);
nand U10804 (N_10804,N_10137,N_10263);
xnor U10805 (N_10805,N_10610,N_10543);
or U10806 (N_10806,N_10036,N_10289);
nand U10807 (N_10807,N_10300,N_10018);
or U10808 (N_10808,N_10042,N_10193);
nor U10809 (N_10809,N_10330,N_10375);
and U10810 (N_10810,N_10528,N_10100);
or U10811 (N_10811,N_10342,N_10469);
nand U10812 (N_10812,N_10529,N_10126);
and U10813 (N_10813,N_10299,N_10401);
xnor U10814 (N_10814,N_10446,N_10553);
or U10815 (N_10815,N_10213,N_10500);
and U10816 (N_10816,N_10517,N_10312);
or U10817 (N_10817,N_10012,N_10387);
nor U10818 (N_10818,N_10257,N_10458);
or U10819 (N_10819,N_10535,N_10582);
or U10820 (N_10820,N_10370,N_10197);
nor U10821 (N_10821,N_10004,N_10082);
nand U10822 (N_10822,N_10145,N_10441);
and U10823 (N_10823,N_10400,N_10602);
nor U10824 (N_10824,N_10488,N_10378);
and U10825 (N_10825,N_10350,N_10138);
nand U10826 (N_10826,N_10425,N_10001);
xor U10827 (N_10827,N_10181,N_10530);
or U10828 (N_10828,N_10266,N_10088);
nand U10829 (N_10829,N_10457,N_10491);
nand U10830 (N_10830,N_10009,N_10298);
or U10831 (N_10831,N_10209,N_10026);
nor U10832 (N_10832,N_10297,N_10512);
xor U10833 (N_10833,N_10214,N_10329);
xnor U10834 (N_10834,N_10279,N_10260);
nand U10835 (N_10835,N_10560,N_10105);
nor U10836 (N_10836,N_10166,N_10540);
nor U10837 (N_10837,N_10120,N_10561);
or U10838 (N_10838,N_10014,N_10362);
nor U10839 (N_10839,N_10438,N_10353);
nand U10840 (N_10840,N_10226,N_10273);
nor U10841 (N_10841,N_10576,N_10368);
or U10842 (N_10842,N_10597,N_10136);
nand U10843 (N_10843,N_10432,N_10327);
xor U10844 (N_10844,N_10427,N_10189);
and U10845 (N_10845,N_10408,N_10035);
nand U10846 (N_10846,N_10288,N_10286);
nor U10847 (N_10847,N_10334,N_10433);
xor U10848 (N_10848,N_10206,N_10442);
nand U10849 (N_10849,N_10365,N_10381);
xor U10850 (N_10850,N_10598,N_10200);
nand U10851 (N_10851,N_10090,N_10303);
nand U10852 (N_10852,N_10101,N_10505);
nand U10853 (N_10853,N_10212,N_10476);
nor U10854 (N_10854,N_10477,N_10419);
xnor U10855 (N_10855,N_10364,N_10210);
nand U10856 (N_10856,N_10002,N_10428);
and U10857 (N_10857,N_10023,N_10341);
nand U10858 (N_10858,N_10118,N_10274);
or U10859 (N_10859,N_10545,N_10519);
or U10860 (N_10860,N_10132,N_10102);
xnor U10861 (N_10861,N_10254,N_10465);
and U10862 (N_10862,N_10251,N_10020);
and U10863 (N_10863,N_10346,N_10536);
nor U10864 (N_10864,N_10570,N_10285);
and U10865 (N_10865,N_10613,N_10550);
nand U10866 (N_10866,N_10222,N_10308);
or U10867 (N_10867,N_10581,N_10022);
and U10868 (N_10868,N_10620,N_10593);
or U10869 (N_10869,N_10287,N_10183);
nand U10870 (N_10870,N_10142,N_10106);
xnor U10871 (N_10871,N_10112,N_10149);
xor U10872 (N_10872,N_10196,N_10514);
nor U10873 (N_10873,N_10156,N_10366);
and U10874 (N_10874,N_10447,N_10129);
nand U10875 (N_10875,N_10084,N_10114);
or U10876 (N_10876,N_10354,N_10407);
or U10877 (N_10877,N_10546,N_10236);
or U10878 (N_10878,N_10122,N_10416);
and U10879 (N_10879,N_10170,N_10520);
nand U10880 (N_10880,N_10056,N_10116);
nor U10881 (N_10881,N_10099,N_10290);
nor U10882 (N_10882,N_10282,N_10070);
or U10883 (N_10883,N_10464,N_10338);
nand U10884 (N_10884,N_10031,N_10037);
nand U10885 (N_10885,N_10093,N_10473);
nor U10886 (N_10886,N_10624,N_10117);
nor U10887 (N_10887,N_10383,N_10489);
or U10888 (N_10888,N_10108,N_10459);
or U10889 (N_10889,N_10376,N_10417);
xor U10890 (N_10890,N_10507,N_10430);
or U10891 (N_10891,N_10372,N_10261);
nor U10892 (N_10892,N_10604,N_10509);
and U10893 (N_10893,N_10414,N_10396);
nor U10894 (N_10894,N_10276,N_10511);
xnor U10895 (N_10895,N_10379,N_10462);
nand U10896 (N_10896,N_10439,N_10131);
nor U10897 (N_10897,N_10539,N_10359);
nand U10898 (N_10898,N_10348,N_10049);
xnor U10899 (N_10899,N_10000,N_10371);
xor U10900 (N_10900,N_10202,N_10412);
nor U10901 (N_10901,N_10121,N_10057);
or U10902 (N_10902,N_10268,N_10010);
nor U10903 (N_10903,N_10496,N_10537);
and U10904 (N_10904,N_10103,N_10336);
and U10905 (N_10905,N_10431,N_10177);
and U10906 (N_10906,N_10277,N_10559);
nor U10907 (N_10907,N_10215,N_10363);
and U10908 (N_10908,N_10367,N_10369);
or U10909 (N_10909,N_10578,N_10064);
or U10910 (N_10910,N_10337,N_10591);
xnor U10911 (N_10911,N_10270,N_10621);
nor U10912 (N_10912,N_10225,N_10562);
and U10913 (N_10913,N_10292,N_10092);
nand U10914 (N_10914,N_10169,N_10256);
and U10915 (N_10915,N_10444,N_10248);
and U10916 (N_10916,N_10508,N_10592);
nand U10917 (N_10917,N_10195,N_10011);
nor U10918 (N_10918,N_10151,N_10043);
nand U10919 (N_10919,N_10237,N_10165);
nand U10920 (N_10920,N_10153,N_10223);
or U10921 (N_10921,N_10217,N_10060);
nor U10922 (N_10922,N_10422,N_10125);
and U10923 (N_10923,N_10614,N_10554);
nor U10924 (N_10924,N_10192,N_10293);
nand U10925 (N_10925,N_10201,N_10382);
nand U10926 (N_10926,N_10580,N_10533);
and U10927 (N_10927,N_10033,N_10374);
xor U10928 (N_10928,N_10146,N_10028);
and U10929 (N_10929,N_10148,N_10571);
and U10930 (N_10930,N_10072,N_10127);
nor U10931 (N_10931,N_10264,N_10119);
and U10932 (N_10932,N_10600,N_10077);
and U10933 (N_10933,N_10390,N_10017);
xor U10934 (N_10934,N_10246,N_10295);
xnor U10935 (N_10935,N_10021,N_10231);
and U10936 (N_10936,N_10157,N_10448);
nor U10937 (N_10937,N_10548,N_10016);
or U10938 (N_10938,N_10046,N_10205);
xnor U10939 (N_10939,N_10211,N_10613);
nand U10940 (N_10940,N_10283,N_10060);
nand U10941 (N_10941,N_10157,N_10121);
xnor U10942 (N_10942,N_10500,N_10049);
xnor U10943 (N_10943,N_10514,N_10440);
nand U10944 (N_10944,N_10357,N_10051);
nor U10945 (N_10945,N_10424,N_10093);
or U10946 (N_10946,N_10239,N_10129);
nor U10947 (N_10947,N_10586,N_10183);
and U10948 (N_10948,N_10490,N_10567);
xnor U10949 (N_10949,N_10165,N_10463);
and U10950 (N_10950,N_10437,N_10182);
nor U10951 (N_10951,N_10476,N_10566);
xor U10952 (N_10952,N_10427,N_10623);
xnor U10953 (N_10953,N_10273,N_10572);
nor U10954 (N_10954,N_10041,N_10136);
and U10955 (N_10955,N_10158,N_10161);
and U10956 (N_10956,N_10255,N_10403);
or U10957 (N_10957,N_10181,N_10286);
xor U10958 (N_10958,N_10364,N_10327);
nand U10959 (N_10959,N_10064,N_10007);
or U10960 (N_10960,N_10428,N_10257);
and U10961 (N_10961,N_10372,N_10067);
or U10962 (N_10962,N_10480,N_10386);
nand U10963 (N_10963,N_10526,N_10269);
nor U10964 (N_10964,N_10232,N_10099);
or U10965 (N_10965,N_10360,N_10115);
nor U10966 (N_10966,N_10230,N_10535);
or U10967 (N_10967,N_10310,N_10205);
xnor U10968 (N_10968,N_10516,N_10138);
nor U10969 (N_10969,N_10384,N_10176);
nor U10970 (N_10970,N_10456,N_10548);
or U10971 (N_10971,N_10553,N_10159);
nand U10972 (N_10972,N_10152,N_10603);
and U10973 (N_10973,N_10589,N_10537);
nor U10974 (N_10974,N_10401,N_10523);
or U10975 (N_10975,N_10501,N_10368);
or U10976 (N_10976,N_10507,N_10333);
or U10977 (N_10977,N_10322,N_10068);
or U10978 (N_10978,N_10301,N_10451);
and U10979 (N_10979,N_10532,N_10542);
nor U10980 (N_10980,N_10220,N_10556);
and U10981 (N_10981,N_10050,N_10073);
or U10982 (N_10982,N_10461,N_10143);
or U10983 (N_10983,N_10193,N_10178);
nand U10984 (N_10984,N_10317,N_10376);
nor U10985 (N_10985,N_10147,N_10315);
nand U10986 (N_10986,N_10542,N_10234);
or U10987 (N_10987,N_10124,N_10113);
and U10988 (N_10988,N_10552,N_10381);
and U10989 (N_10989,N_10031,N_10361);
nand U10990 (N_10990,N_10228,N_10245);
xor U10991 (N_10991,N_10514,N_10067);
and U10992 (N_10992,N_10194,N_10413);
or U10993 (N_10993,N_10193,N_10571);
nand U10994 (N_10994,N_10346,N_10538);
xnor U10995 (N_10995,N_10527,N_10362);
xor U10996 (N_10996,N_10473,N_10616);
and U10997 (N_10997,N_10493,N_10464);
or U10998 (N_10998,N_10170,N_10497);
nor U10999 (N_10999,N_10405,N_10403);
or U11000 (N_11000,N_10073,N_10596);
nor U11001 (N_11001,N_10071,N_10472);
or U11002 (N_11002,N_10511,N_10598);
or U11003 (N_11003,N_10259,N_10200);
nand U11004 (N_11004,N_10581,N_10272);
xor U11005 (N_11005,N_10485,N_10113);
xnor U11006 (N_11006,N_10294,N_10134);
and U11007 (N_11007,N_10544,N_10325);
nor U11008 (N_11008,N_10516,N_10447);
and U11009 (N_11009,N_10365,N_10010);
nor U11010 (N_11010,N_10536,N_10004);
xor U11011 (N_11011,N_10075,N_10330);
or U11012 (N_11012,N_10058,N_10619);
and U11013 (N_11013,N_10607,N_10446);
xor U11014 (N_11014,N_10443,N_10038);
nand U11015 (N_11015,N_10171,N_10218);
and U11016 (N_11016,N_10621,N_10146);
xor U11017 (N_11017,N_10409,N_10083);
nand U11018 (N_11018,N_10333,N_10251);
xnor U11019 (N_11019,N_10557,N_10309);
or U11020 (N_11020,N_10464,N_10260);
and U11021 (N_11021,N_10496,N_10586);
nand U11022 (N_11022,N_10273,N_10093);
xor U11023 (N_11023,N_10014,N_10230);
nand U11024 (N_11024,N_10256,N_10489);
or U11025 (N_11025,N_10275,N_10105);
or U11026 (N_11026,N_10423,N_10060);
nand U11027 (N_11027,N_10166,N_10229);
xnor U11028 (N_11028,N_10275,N_10401);
or U11029 (N_11029,N_10216,N_10475);
nor U11030 (N_11030,N_10061,N_10173);
nand U11031 (N_11031,N_10616,N_10364);
and U11032 (N_11032,N_10154,N_10104);
xnor U11033 (N_11033,N_10227,N_10352);
nand U11034 (N_11034,N_10233,N_10109);
and U11035 (N_11035,N_10185,N_10496);
and U11036 (N_11036,N_10354,N_10140);
nor U11037 (N_11037,N_10282,N_10116);
nand U11038 (N_11038,N_10025,N_10362);
or U11039 (N_11039,N_10102,N_10447);
nor U11040 (N_11040,N_10497,N_10258);
xor U11041 (N_11041,N_10120,N_10415);
nand U11042 (N_11042,N_10293,N_10000);
nor U11043 (N_11043,N_10338,N_10247);
and U11044 (N_11044,N_10034,N_10199);
nor U11045 (N_11045,N_10613,N_10572);
nand U11046 (N_11046,N_10143,N_10202);
xor U11047 (N_11047,N_10472,N_10347);
nand U11048 (N_11048,N_10440,N_10406);
or U11049 (N_11049,N_10037,N_10318);
or U11050 (N_11050,N_10362,N_10022);
and U11051 (N_11051,N_10346,N_10231);
nor U11052 (N_11052,N_10021,N_10044);
nand U11053 (N_11053,N_10563,N_10082);
and U11054 (N_11054,N_10498,N_10470);
nand U11055 (N_11055,N_10526,N_10275);
nand U11056 (N_11056,N_10097,N_10085);
or U11057 (N_11057,N_10012,N_10428);
nor U11058 (N_11058,N_10105,N_10542);
or U11059 (N_11059,N_10398,N_10106);
nand U11060 (N_11060,N_10104,N_10131);
or U11061 (N_11061,N_10468,N_10100);
xnor U11062 (N_11062,N_10420,N_10542);
and U11063 (N_11063,N_10396,N_10388);
or U11064 (N_11064,N_10553,N_10309);
and U11065 (N_11065,N_10320,N_10132);
nor U11066 (N_11066,N_10077,N_10352);
and U11067 (N_11067,N_10448,N_10050);
and U11068 (N_11068,N_10481,N_10425);
nor U11069 (N_11069,N_10337,N_10207);
or U11070 (N_11070,N_10470,N_10499);
nor U11071 (N_11071,N_10152,N_10192);
nor U11072 (N_11072,N_10037,N_10326);
and U11073 (N_11073,N_10330,N_10469);
nand U11074 (N_11074,N_10073,N_10190);
nor U11075 (N_11075,N_10024,N_10289);
nor U11076 (N_11076,N_10267,N_10011);
and U11077 (N_11077,N_10594,N_10072);
nor U11078 (N_11078,N_10593,N_10412);
or U11079 (N_11079,N_10394,N_10443);
nor U11080 (N_11080,N_10289,N_10245);
or U11081 (N_11081,N_10279,N_10577);
or U11082 (N_11082,N_10208,N_10294);
nor U11083 (N_11083,N_10499,N_10172);
xor U11084 (N_11084,N_10281,N_10577);
nor U11085 (N_11085,N_10435,N_10057);
nor U11086 (N_11086,N_10589,N_10247);
or U11087 (N_11087,N_10524,N_10361);
xor U11088 (N_11088,N_10105,N_10155);
or U11089 (N_11089,N_10280,N_10499);
or U11090 (N_11090,N_10380,N_10389);
or U11091 (N_11091,N_10036,N_10498);
nand U11092 (N_11092,N_10087,N_10266);
or U11093 (N_11093,N_10531,N_10016);
nand U11094 (N_11094,N_10458,N_10348);
or U11095 (N_11095,N_10605,N_10394);
or U11096 (N_11096,N_10172,N_10597);
and U11097 (N_11097,N_10556,N_10080);
or U11098 (N_11098,N_10480,N_10029);
nor U11099 (N_11099,N_10013,N_10190);
nand U11100 (N_11100,N_10369,N_10081);
nand U11101 (N_11101,N_10465,N_10471);
and U11102 (N_11102,N_10074,N_10288);
and U11103 (N_11103,N_10302,N_10256);
nor U11104 (N_11104,N_10579,N_10042);
nor U11105 (N_11105,N_10309,N_10034);
nand U11106 (N_11106,N_10519,N_10550);
or U11107 (N_11107,N_10014,N_10469);
nor U11108 (N_11108,N_10612,N_10287);
nor U11109 (N_11109,N_10120,N_10585);
xor U11110 (N_11110,N_10489,N_10576);
or U11111 (N_11111,N_10423,N_10477);
nor U11112 (N_11112,N_10127,N_10472);
nand U11113 (N_11113,N_10515,N_10483);
and U11114 (N_11114,N_10565,N_10313);
nand U11115 (N_11115,N_10208,N_10275);
nor U11116 (N_11116,N_10217,N_10348);
nor U11117 (N_11117,N_10115,N_10218);
and U11118 (N_11118,N_10238,N_10248);
or U11119 (N_11119,N_10248,N_10464);
and U11120 (N_11120,N_10449,N_10602);
and U11121 (N_11121,N_10374,N_10547);
nor U11122 (N_11122,N_10142,N_10497);
and U11123 (N_11123,N_10033,N_10277);
nor U11124 (N_11124,N_10479,N_10293);
or U11125 (N_11125,N_10487,N_10276);
nand U11126 (N_11126,N_10288,N_10143);
nand U11127 (N_11127,N_10489,N_10036);
nor U11128 (N_11128,N_10372,N_10164);
nand U11129 (N_11129,N_10212,N_10067);
xor U11130 (N_11130,N_10585,N_10398);
nor U11131 (N_11131,N_10312,N_10400);
nand U11132 (N_11132,N_10269,N_10272);
and U11133 (N_11133,N_10503,N_10102);
nor U11134 (N_11134,N_10414,N_10142);
and U11135 (N_11135,N_10124,N_10335);
and U11136 (N_11136,N_10209,N_10495);
or U11137 (N_11137,N_10091,N_10105);
xnor U11138 (N_11138,N_10135,N_10225);
or U11139 (N_11139,N_10036,N_10080);
or U11140 (N_11140,N_10301,N_10181);
nand U11141 (N_11141,N_10422,N_10333);
and U11142 (N_11142,N_10231,N_10088);
xnor U11143 (N_11143,N_10043,N_10150);
or U11144 (N_11144,N_10234,N_10466);
nand U11145 (N_11145,N_10577,N_10332);
and U11146 (N_11146,N_10517,N_10240);
and U11147 (N_11147,N_10200,N_10617);
nand U11148 (N_11148,N_10307,N_10178);
nor U11149 (N_11149,N_10411,N_10128);
and U11150 (N_11150,N_10529,N_10150);
or U11151 (N_11151,N_10096,N_10331);
and U11152 (N_11152,N_10520,N_10139);
nor U11153 (N_11153,N_10548,N_10623);
xnor U11154 (N_11154,N_10601,N_10503);
nand U11155 (N_11155,N_10082,N_10565);
and U11156 (N_11156,N_10012,N_10340);
nor U11157 (N_11157,N_10418,N_10029);
xnor U11158 (N_11158,N_10202,N_10565);
xor U11159 (N_11159,N_10164,N_10382);
and U11160 (N_11160,N_10200,N_10586);
nand U11161 (N_11161,N_10578,N_10190);
nand U11162 (N_11162,N_10411,N_10405);
and U11163 (N_11163,N_10097,N_10570);
or U11164 (N_11164,N_10232,N_10519);
nor U11165 (N_11165,N_10495,N_10044);
nor U11166 (N_11166,N_10547,N_10280);
nand U11167 (N_11167,N_10413,N_10182);
or U11168 (N_11168,N_10476,N_10233);
or U11169 (N_11169,N_10078,N_10260);
or U11170 (N_11170,N_10306,N_10016);
and U11171 (N_11171,N_10397,N_10211);
nor U11172 (N_11172,N_10621,N_10367);
and U11173 (N_11173,N_10013,N_10274);
xor U11174 (N_11174,N_10434,N_10094);
xor U11175 (N_11175,N_10268,N_10297);
nand U11176 (N_11176,N_10304,N_10249);
or U11177 (N_11177,N_10289,N_10419);
nor U11178 (N_11178,N_10289,N_10167);
xor U11179 (N_11179,N_10548,N_10358);
and U11180 (N_11180,N_10076,N_10599);
nand U11181 (N_11181,N_10569,N_10211);
nor U11182 (N_11182,N_10392,N_10157);
xor U11183 (N_11183,N_10020,N_10148);
nand U11184 (N_11184,N_10360,N_10428);
xor U11185 (N_11185,N_10072,N_10035);
xor U11186 (N_11186,N_10559,N_10521);
xor U11187 (N_11187,N_10151,N_10527);
or U11188 (N_11188,N_10368,N_10391);
and U11189 (N_11189,N_10470,N_10000);
and U11190 (N_11190,N_10140,N_10304);
xnor U11191 (N_11191,N_10398,N_10520);
and U11192 (N_11192,N_10208,N_10073);
xnor U11193 (N_11193,N_10027,N_10552);
nand U11194 (N_11194,N_10278,N_10248);
xnor U11195 (N_11195,N_10407,N_10093);
or U11196 (N_11196,N_10140,N_10406);
xor U11197 (N_11197,N_10064,N_10430);
and U11198 (N_11198,N_10332,N_10418);
nand U11199 (N_11199,N_10526,N_10210);
or U11200 (N_11200,N_10462,N_10169);
and U11201 (N_11201,N_10089,N_10052);
xor U11202 (N_11202,N_10178,N_10614);
nor U11203 (N_11203,N_10238,N_10356);
nand U11204 (N_11204,N_10164,N_10282);
and U11205 (N_11205,N_10450,N_10046);
nand U11206 (N_11206,N_10087,N_10401);
nor U11207 (N_11207,N_10302,N_10002);
nand U11208 (N_11208,N_10485,N_10073);
nor U11209 (N_11209,N_10427,N_10506);
nand U11210 (N_11210,N_10564,N_10159);
and U11211 (N_11211,N_10272,N_10516);
or U11212 (N_11212,N_10149,N_10588);
or U11213 (N_11213,N_10241,N_10327);
xor U11214 (N_11214,N_10077,N_10621);
or U11215 (N_11215,N_10376,N_10546);
nor U11216 (N_11216,N_10304,N_10381);
or U11217 (N_11217,N_10280,N_10608);
xnor U11218 (N_11218,N_10622,N_10181);
xor U11219 (N_11219,N_10440,N_10101);
or U11220 (N_11220,N_10318,N_10057);
and U11221 (N_11221,N_10003,N_10082);
nor U11222 (N_11222,N_10085,N_10538);
nand U11223 (N_11223,N_10437,N_10204);
xnor U11224 (N_11224,N_10609,N_10191);
and U11225 (N_11225,N_10358,N_10060);
or U11226 (N_11226,N_10493,N_10192);
or U11227 (N_11227,N_10419,N_10511);
nand U11228 (N_11228,N_10305,N_10565);
nor U11229 (N_11229,N_10551,N_10218);
xnor U11230 (N_11230,N_10066,N_10453);
and U11231 (N_11231,N_10319,N_10553);
nand U11232 (N_11232,N_10027,N_10120);
or U11233 (N_11233,N_10085,N_10135);
nand U11234 (N_11234,N_10593,N_10067);
or U11235 (N_11235,N_10523,N_10002);
nor U11236 (N_11236,N_10156,N_10213);
and U11237 (N_11237,N_10022,N_10271);
xor U11238 (N_11238,N_10477,N_10336);
nand U11239 (N_11239,N_10336,N_10176);
and U11240 (N_11240,N_10124,N_10028);
nand U11241 (N_11241,N_10586,N_10120);
nand U11242 (N_11242,N_10234,N_10579);
nand U11243 (N_11243,N_10107,N_10561);
xnor U11244 (N_11244,N_10066,N_10006);
xnor U11245 (N_11245,N_10123,N_10172);
nor U11246 (N_11246,N_10460,N_10042);
and U11247 (N_11247,N_10494,N_10559);
xnor U11248 (N_11248,N_10619,N_10579);
xor U11249 (N_11249,N_10355,N_10325);
nor U11250 (N_11250,N_10882,N_10956);
nor U11251 (N_11251,N_10783,N_11248);
nor U11252 (N_11252,N_11145,N_10631);
and U11253 (N_11253,N_11215,N_11217);
and U11254 (N_11254,N_11247,N_10877);
or U11255 (N_11255,N_10648,N_11245);
and U11256 (N_11256,N_11119,N_11001);
nand U11257 (N_11257,N_10665,N_10975);
nand U11258 (N_11258,N_11195,N_11120);
xnor U11259 (N_11259,N_11249,N_11133);
nand U11260 (N_11260,N_10723,N_10993);
nor U11261 (N_11261,N_10827,N_10878);
nand U11262 (N_11262,N_11115,N_11040);
xor U11263 (N_11263,N_11081,N_11170);
or U11264 (N_11264,N_11136,N_10928);
and U11265 (N_11265,N_10806,N_10999);
nor U11266 (N_11266,N_10881,N_11240);
or U11267 (N_11267,N_10664,N_10946);
nand U11268 (N_11268,N_11153,N_11235);
or U11269 (N_11269,N_11039,N_11163);
or U11270 (N_11270,N_10786,N_11194);
nand U11271 (N_11271,N_11222,N_10699);
xor U11272 (N_11272,N_10867,N_10779);
or U11273 (N_11273,N_11174,N_10693);
nor U11274 (N_11274,N_11054,N_10629);
or U11275 (N_11275,N_11062,N_10793);
nand U11276 (N_11276,N_10778,N_11203);
xor U11277 (N_11277,N_11209,N_10770);
xor U11278 (N_11278,N_10897,N_10940);
xor U11279 (N_11279,N_10724,N_11078);
and U11280 (N_11280,N_10772,N_11086);
nand U11281 (N_11281,N_11157,N_11049);
xor U11282 (N_11282,N_10938,N_10791);
xor U11283 (N_11283,N_11074,N_11205);
nor U11284 (N_11284,N_11042,N_11123);
xor U11285 (N_11285,N_10874,N_11094);
xor U11286 (N_11286,N_10962,N_10990);
or U11287 (N_11287,N_10849,N_11116);
nand U11288 (N_11288,N_10932,N_10846);
or U11289 (N_11289,N_11233,N_11193);
xor U11290 (N_11290,N_11101,N_11038);
nor U11291 (N_11291,N_10773,N_11003);
nor U11292 (N_11292,N_11131,N_10769);
nor U11293 (N_11293,N_11162,N_11139);
and U11294 (N_11294,N_11018,N_10949);
or U11295 (N_11295,N_11058,N_10644);
xor U11296 (N_11296,N_10913,N_10727);
nor U11297 (N_11297,N_11085,N_10715);
xor U11298 (N_11298,N_10972,N_11009);
and U11299 (N_11299,N_10954,N_10752);
and U11300 (N_11300,N_11089,N_11099);
nor U11301 (N_11301,N_10805,N_11005);
xor U11302 (N_11302,N_11007,N_10829);
and U11303 (N_11303,N_10697,N_11188);
and U11304 (N_11304,N_11226,N_11114);
nor U11305 (N_11305,N_10689,N_10684);
or U11306 (N_11306,N_10777,N_10771);
nor U11307 (N_11307,N_10696,N_10929);
nand U11308 (N_11308,N_10994,N_10841);
nor U11309 (N_11309,N_10785,N_10804);
or U11310 (N_11310,N_11064,N_10869);
xnor U11311 (N_11311,N_10901,N_10662);
and U11312 (N_11312,N_10908,N_10981);
nor U11313 (N_11313,N_11199,N_10933);
or U11314 (N_11314,N_10987,N_10916);
nor U11315 (N_11315,N_10839,N_10930);
or U11316 (N_11316,N_11127,N_10961);
or U11317 (N_11317,N_11109,N_10904);
and U11318 (N_11318,N_11160,N_10967);
or U11319 (N_11319,N_11204,N_11095);
or U11320 (N_11320,N_10812,N_11142);
and U11321 (N_11321,N_10766,N_11105);
nor U11322 (N_11322,N_11055,N_10926);
and U11323 (N_11323,N_10982,N_10969);
nor U11324 (N_11324,N_11161,N_10645);
nand U11325 (N_11325,N_10711,N_10847);
nor U11326 (N_11326,N_10814,N_10953);
and U11327 (N_11327,N_11106,N_11167);
and U11328 (N_11328,N_10682,N_11197);
nand U11329 (N_11329,N_11056,N_10707);
or U11330 (N_11330,N_11093,N_11213);
nor U11331 (N_11331,N_10695,N_11206);
nor U11332 (N_11332,N_10730,N_10633);
and U11333 (N_11333,N_11239,N_10894);
nand U11334 (N_11334,N_11219,N_10957);
xnor U11335 (N_11335,N_10688,N_10765);
or U11336 (N_11336,N_10810,N_10870);
and U11337 (N_11337,N_10979,N_10911);
nor U11338 (N_11338,N_10927,N_10714);
nor U11339 (N_11339,N_11192,N_10892);
or U11340 (N_11340,N_11137,N_11212);
or U11341 (N_11341,N_11067,N_10641);
xor U11342 (N_11342,N_10694,N_10635);
xor U11343 (N_11343,N_10833,N_10722);
nor U11344 (N_11344,N_10815,N_11069);
nor U11345 (N_11345,N_11096,N_10922);
nor U11346 (N_11346,N_10780,N_10731);
nand U11347 (N_11347,N_11243,N_10840);
nor U11348 (N_11348,N_10658,N_11234);
xor U11349 (N_11349,N_10983,N_10835);
or U11350 (N_11350,N_10970,N_10895);
or U11351 (N_11351,N_11098,N_10676);
nor U11352 (N_11352,N_10971,N_10670);
nand U11353 (N_11353,N_11061,N_10995);
and U11354 (N_11354,N_10796,N_10755);
xor U11355 (N_11355,N_10891,N_10675);
nor U11356 (N_11356,N_10989,N_10701);
and U11357 (N_11357,N_10705,N_10753);
xor U11358 (N_11358,N_11208,N_11113);
nor U11359 (N_11359,N_11236,N_10842);
xor U11360 (N_11360,N_11237,N_10948);
nand U11361 (N_11361,N_11232,N_10817);
and U11362 (N_11362,N_10844,N_11140);
nor U11363 (N_11363,N_11190,N_10960);
nand U11364 (N_11364,N_11050,N_11057);
nand U11365 (N_11365,N_10825,N_10800);
xnor U11366 (N_11366,N_10795,N_10678);
nand U11367 (N_11367,N_10674,N_10721);
and U11368 (N_11368,N_10716,N_10743);
and U11369 (N_11369,N_11218,N_10655);
xnor U11370 (N_11370,N_10883,N_10907);
xor U11371 (N_11371,N_10725,N_11126);
xnor U11372 (N_11372,N_11238,N_10666);
xnor U11373 (N_11373,N_10855,N_11144);
or U11374 (N_11374,N_11229,N_10683);
nor U11375 (N_11375,N_10843,N_10851);
xnor U11376 (N_11376,N_10977,N_10939);
or U11377 (N_11377,N_10768,N_10638);
or U11378 (N_11378,N_10637,N_10950);
nand U11379 (N_11379,N_11191,N_11075);
or U11380 (N_11380,N_10914,N_10729);
or U11381 (N_11381,N_10710,N_10873);
nor U11382 (N_11382,N_11023,N_10738);
or U11383 (N_11383,N_10834,N_11066);
or U11384 (N_11384,N_11032,N_10642);
or U11385 (N_11385,N_10630,N_11200);
and U11386 (N_11386,N_10947,N_11117);
nor U11387 (N_11387,N_11100,N_11207);
nand U11388 (N_11388,N_10692,N_10968);
nor U11389 (N_11389,N_11189,N_10660);
nor U11390 (N_11390,N_10709,N_11181);
xnor U11391 (N_11391,N_10671,N_10634);
nor U11392 (N_11392,N_10733,N_10875);
nor U11393 (N_11393,N_11010,N_11125);
or U11394 (N_11394,N_11026,N_11172);
or U11395 (N_11395,N_11227,N_10749);
nor U11396 (N_11396,N_10708,N_10964);
and U11397 (N_11397,N_10826,N_10668);
xor U11398 (N_11398,N_10871,N_11065);
xnor U11399 (N_11399,N_11013,N_11076);
and U11400 (N_11400,N_10864,N_11068);
and U11401 (N_11401,N_10647,N_10976);
or U11402 (N_11402,N_10677,N_10736);
nand U11403 (N_11403,N_10985,N_10980);
nor U11404 (N_11404,N_11122,N_11008);
xor U11405 (N_11405,N_11045,N_10845);
nand U11406 (N_11406,N_10673,N_10718);
nand U11407 (N_11407,N_10910,N_10986);
xnor U11408 (N_11408,N_11073,N_11029);
or U11409 (N_11409,N_11108,N_11129);
nand U11410 (N_11410,N_10659,N_10737);
nand U11411 (N_11411,N_10988,N_10945);
and U11412 (N_11412,N_10650,N_10799);
nand U11413 (N_11413,N_11148,N_11090);
nor U11414 (N_11414,N_10915,N_10672);
nand U11415 (N_11415,N_11230,N_11168);
nor U11416 (N_11416,N_11110,N_11225);
or U11417 (N_11417,N_10998,N_10681);
or U11418 (N_11418,N_10703,N_10925);
and U11419 (N_11419,N_10775,N_10852);
xnor U11420 (N_11420,N_11130,N_10754);
nor U11421 (N_11421,N_11165,N_11036);
or U11422 (N_11422,N_10764,N_10717);
or U11423 (N_11423,N_10880,N_11143);
nand U11424 (N_11424,N_10746,N_11052);
nand U11425 (N_11425,N_10784,N_10811);
xor U11426 (N_11426,N_10888,N_10640);
nor U11427 (N_11427,N_10854,N_11037);
xnor U11428 (N_11428,N_10896,N_10719);
and U11429 (N_11429,N_11211,N_10757);
nand U11430 (N_11430,N_10991,N_10767);
nor U11431 (N_11431,N_11002,N_11047);
nand U11432 (N_11432,N_11201,N_11151);
and U11433 (N_11433,N_11084,N_11152);
nand U11434 (N_11434,N_10838,N_11088);
xnor U11435 (N_11435,N_11000,N_10798);
xnor U11436 (N_11436,N_11242,N_10984);
and U11437 (N_11437,N_11132,N_10959);
nor U11438 (N_11438,N_11053,N_10996);
nand U11439 (N_11439,N_10776,N_10889);
and U11440 (N_11440,N_10626,N_11185);
or U11441 (N_11441,N_10884,N_10832);
and U11442 (N_11442,N_11011,N_10763);
nor U11443 (N_11443,N_10735,N_11155);
or U11444 (N_11444,N_11231,N_10742);
and U11445 (N_11445,N_10978,N_10879);
nor U11446 (N_11446,N_11214,N_10850);
or U11447 (N_11447,N_11059,N_11080);
nor U11448 (N_11448,N_11186,N_10702);
nand U11449 (N_11449,N_10628,N_10813);
xor U11450 (N_11450,N_10905,N_10848);
and U11451 (N_11451,N_10704,N_11202);
nand U11452 (N_11452,N_11246,N_11150);
nor U11453 (N_11453,N_10906,N_10712);
xnor U11454 (N_11454,N_11027,N_10789);
nor U11455 (N_11455,N_10762,N_10781);
and U11456 (N_11456,N_10963,N_10912);
or U11457 (N_11457,N_10741,N_11012);
nor U11458 (N_11458,N_11025,N_11124);
or U11459 (N_11459,N_10822,N_11134);
xor U11460 (N_11460,N_10898,N_10790);
or U11461 (N_11461,N_11082,N_11166);
or U11462 (N_11462,N_10649,N_11118);
and U11463 (N_11463,N_11121,N_10732);
or U11464 (N_11464,N_10747,N_11224);
nor U11465 (N_11465,N_11031,N_10809);
and U11466 (N_11466,N_10820,N_11164);
and U11467 (N_11467,N_10824,N_10821);
nand U11468 (N_11468,N_10816,N_11024);
and U11469 (N_11469,N_11173,N_11028);
or U11470 (N_11470,N_11030,N_10782);
nor U11471 (N_11471,N_10687,N_10856);
nor U11472 (N_11472,N_11071,N_10974);
nor U11473 (N_11473,N_10679,N_10698);
xor U11474 (N_11474,N_11046,N_11063);
xor U11475 (N_11475,N_10934,N_11033);
or U11476 (N_11476,N_10745,N_11146);
nand U11477 (N_11477,N_10734,N_11022);
nor U11478 (N_11478,N_10652,N_11180);
and U11479 (N_11479,N_10863,N_10935);
nand U11480 (N_11480,N_10992,N_11079);
or U11481 (N_11481,N_10958,N_11244);
or U11482 (N_11482,N_10686,N_10663);
or U11483 (N_11483,N_10759,N_10876);
nor U11484 (N_11484,N_11177,N_10803);
or U11485 (N_11485,N_10691,N_10819);
nor U11486 (N_11486,N_10942,N_11017);
nor U11487 (N_11487,N_11178,N_10900);
and U11488 (N_11488,N_10627,N_10941);
nand U11489 (N_11489,N_11112,N_11210);
and U11490 (N_11490,N_11128,N_10861);
and U11491 (N_11491,N_10858,N_11141);
or U11492 (N_11492,N_11004,N_11035);
xnor U11493 (N_11493,N_10919,N_10706);
nand U11494 (N_11494,N_11149,N_11158);
or U11495 (N_11495,N_11103,N_11044);
and U11496 (N_11496,N_10973,N_10787);
or U11497 (N_11497,N_10893,N_10887);
or U11498 (N_11498,N_11169,N_11077);
nand U11499 (N_11499,N_11223,N_10920);
and U11500 (N_11500,N_10903,N_11241);
nor U11501 (N_11501,N_11159,N_10792);
and U11502 (N_11502,N_10951,N_11184);
xnor U11503 (N_11503,N_10750,N_10756);
nand U11504 (N_11504,N_11179,N_10865);
or U11505 (N_11505,N_11087,N_10760);
nand U11506 (N_11506,N_10955,N_10685);
and U11507 (N_11507,N_10936,N_10830);
nor U11508 (N_11508,N_10924,N_10944);
nor U11509 (N_11509,N_10885,N_10917);
and U11510 (N_11510,N_10868,N_11006);
nand U11511 (N_11511,N_11060,N_11092);
and U11512 (N_11512,N_10866,N_10651);
nor U11513 (N_11513,N_10952,N_10859);
xnor U11514 (N_11514,N_10831,N_11104);
nor U11515 (N_11515,N_10636,N_10857);
nand U11516 (N_11516,N_11020,N_10656);
or U11517 (N_11517,N_10890,N_10653);
nand U11518 (N_11518,N_10774,N_11070);
nor U11519 (N_11519,N_10899,N_11147);
or U11520 (N_11520,N_11016,N_11091);
xor U11521 (N_11521,N_11072,N_10909);
or U11522 (N_11522,N_10836,N_10739);
nor U11523 (N_11523,N_10801,N_11048);
or U11524 (N_11524,N_10794,N_10643);
or U11525 (N_11525,N_10740,N_11156);
or U11526 (N_11526,N_10728,N_11138);
and U11527 (N_11527,N_11187,N_11019);
xnor U11528 (N_11528,N_11175,N_10921);
or U11529 (N_11529,N_10797,N_10761);
xor U11530 (N_11530,N_10802,N_11107);
nor U11531 (N_11531,N_11198,N_10657);
and U11532 (N_11532,N_10931,N_10886);
xor U11533 (N_11533,N_10902,N_11154);
nor U11534 (N_11534,N_10828,N_10744);
or U11535 (N_11535,N_11102,N_11135);
nand U11536 (N_11536,N_10807,N_11183);
or U11537 (N_11537,N_11171,N_10632);
or U11538 (N_11538,N_11221,N_11014);
nor U11539 (N_11539,N_10818,N_10837);
nor U11540 (N_11540,N_11216,N_10667);
xor U11541 (N_11541,N_10713,N_11228);
xnor U11542 (N_11542,N_10918,N_10965);
and U11543 (N_11543,N_10625,N_10853);
nor U11544 (N_11544,N_10720,N_10808);
nor U11545 (N_11545,N_10943,N_11021);
nand U11546 (N_11546,N_11182,N_11051);
nor U11547 (N_11547,N_10680,N_10669);
nor U11548 (N_11548,N_10823,N_11196);
and U11549 (N_11549,N_10862,N_11176);
and U11550 (N_11550,N_10997,N_10751);
and U11551 (N_11551,N_10661,N_11015);
nand U11552 (N_11552,N_10748,N_10966);
or U11553 (N_11553,N_10639,N_11083);
or U11554 (N_11554,N_11043,N_11097);
and U11555 (N_11555,N_10726,N_10758);
and U11556 (N_11556,N_10860,N_10872);
and U11557 (N_11557,N_10646,N_11034);
or U11558 (N_11558,N_10937,N_10788);
nand U11559 (N_11559,N_10700,N_10923);
nand U11560 (N_11560,N_10654,N_11220);
nor U11561 (N_11561,N_10690,N_11111);
or U11562 (N_11562,N_11041,N_10868);
nand U11563 (N_11563,N_11179,N_10883);
or U11564 (N_11564,N_10719,N_11020);
and U11565 (N_11565,N_10780,N_10935);
xnor U11566 (N_11566,N_10970,N_10719);
nand U11567 (N_11567,N_10887,N_10915);
xor U11568 (N_11568,N_10749,N_11013);
nand U11569 (N_11569,N_11066,N_10736);
nor U11570 (N_11570,N_11072,N_11192);
xor U11571 (N_11571,N_10871,N_10750);
and U11572 (N_11572,N_10802,N_11039);
and U11573 (N_11573,N_10904,N_11064);
and U11574 (N_11574,N_10933,N_11026);
or U11575 (N_11575,N_10651,N_10937);
xnor U11576 (N_11576,N_10646,N_11108);
nor U11577 (N_11577,N_10883,N_10634);
xnor U11578 (N_11578,N_10785,N_10815);
nor U11579 (N_11579,N_11003,N_11070);
and U11580 (N_11580,N_10820,N_11175);
xnor U11581 (N_11581,N_10827,N_10717);
xor U11582 (N_11582,N_10871,N_10854);
xor U11583 (N_11583,N_10986,N_11211);
xor U11584 (N_11584,N_10885,N_11141);
nand U11585 (N_11585,N_10797,N_11061);
xnor U11586 (N_11586,N_10663,N_10662);
nand U11587 (N_11587,N_10947,N_11193);
nor U11588 (N_11588,N_10840,N_11136);
nand U11589 (N_11589,N_10808,N_10931);
nand U11590 (N_11590,N_10859,N_10633);
or U11591 (N_11591,N_10997,N_11028);
nor U11592 (N_11592,N_10752,N_11223);
xnor U11593 (N_11593,N_10663,N_11005);
or U11594 (N_11594,N_10883,N_10981);
nor U11595 (N_11595,N_10937,N_11078);
nand U11596 (N_11596,N_10944,N_10823);
or U11597 (N_11597,N_10705,N_10652);
xnor U11598 (N_11598,N_10777,N_10697);
xor U11599 (N_11599,N_11162,N_11180);
nand U11600 (N_11600,N_10656,N_11191);
nand U11601 (N_11601,N_10786,N_11154);
or U11602 (N_11602,N_11115,N_11108);
or U11603 (N_11603,N_11167,N_11163);
xnor U11604 (N_11604,N_10956,N_10769);
and U11605 (N_11605,N_10833,N_11117);
xnor U11606 (N_11606,N_11040,N_10817);
and U11607 (N_11607,N_11013,N_11207);
and U11608 (N_11608,N_11091,N_10910);
xor U11609 (N_11609,N_10741,N_10906);
nand U11610 (N_11610,N_11034,N_10980);
xnor U11611 (N_11611,N_10756,N_11096);
nand U11612 (N_11612,N_11069,N_10734);
xnor U11613 (N_11613,N_11168,N_11103);
or U11614 (N_11614,N_11118,N_11183);
and U11615 (N_11615,N_11107,N_10825);
xor U11616 (N_11616,N_10976,N_10785);
nand U11617 (N_11617,N_11052,N_11064);
or U11618 (N_11618,N_10696,N_11170);
and U11619 (N_11619,N_10628,N_10922);
nor U11620 (N_11620,N_10747,N_10921);
nand U11621 (N_11621,N_10957,N_11209);
nor U11622 (N_11622,N_11171,N_10858);
or U11623 (N_11623,N_10896,N_10656);
or U11624 (N_11624,N_11015,N_11239);
nor U11625 (N_11625,N_11207,N_11163);
nand U11626 (N_11626,N_10851,N_10877);
nand U11627 (N_11627,N_10961,N_11025);
nand U11628 (N_11628,N_10793,N_10668);
xor U11629 (N_11629,N_11148,N_10775);
nor U11630 (N_11630,N_10718,N_11064);
xor U11631 (N_11631,N_11131,N_11225);
nand U11632 (N_11632,N_11034,N_10843);
nand U11633 (N_11633,N_11241,N_10963);
nor U11634 (N_11634,N_11122,N_11230);
and U11635 (N_11635,N_11235,N_10919);
nand U11636 (N_11636,N_10975,N_11063);
or U11637 (N_11637,N_11116,N_10972);
xor U11638 (N_11638,N_11213,N_10746);
nand U11639 (N_11639,N_10769,N_10723);
or U11640 (N_11640,N_10976,N_10652);
and U11641 (N_11641,N_11197,N_10760);
xor U11642 (N_11642,N_10631,N_11010);
nand U11643 (N_11643,N_11137,N_11152);
nor U11644 (N_11644,N_11041,N_10905);
nand U11645 (N_11645,N_11211,N_10931);
or U11646 (N_11646,N_10911,N_10792);
and U11647 (N_11647,N_11089,N_11180);
xnor U11648 (N_11648,N_10698,N_10922);
nor U11649 (N_11649,N_10631,N_10924);
and U11650 (N_11650,N_10828,N_10681);
or U11651 (N_11651,N_10770,N_11078);
or U11652 (N_11652,N_10967,N_10677);
nor U11653 (N_11653,N_11098,N_10648);
nand U11654 (N_11654,N_10671,N_11212);
nand U11655 (N_11655,N_10940,N_10817);
or U11656 (N_11656,N_10787,N_10731);
and U11657 (N_11657,N_10644,N_10865);
nand U11658 (N_11658,N_10656,N_10667);
or U11659 (N_11659,N_11201,N_10767);
or U11660 (N_11660,N_10795,N_11112);
nand U11661 (N_11661,N_10986,N_10894);
or U11662 (N_11662,N_10659,N_10690);
or U11663 (N_11663,N_11003,N_10694);
nand U11664 (N_11664,N_11032,N_10856);
xor U11665 (N_11665,N_10948,N_10969);
xnor U11666 (N_11666,N_11214,N_10846);
nor U11667 (N_11667,N_10859,N_10684);
xnor U11668 (N_11668,N_11143,N_10710);
and U11669 (N_11669,N_10715,N_10821);
or U11670 (N_11670,N_11099,N_11193);
xnor U11671 (N_11671,N_10748,N_10915);
nand U11672 (N_11672,N_10625,N_10631);
xnor U11673 (N_11673,N_11153,N_11144);
nor U11674 (N_11674,N_11151,N_10815);
xor U11675 (N_11675,N_11091,N_11033);
nor U11676 (N_11676,N_10748,N_10901);
or U11677 (N_11677,N_11160,N_10734);
and U11678 (N_11678,N_11017,N_10966);
or U11679 (N_11679,N_10809,N_11051);
xnor U11680 (N_11680,N_10787,N_11151);
or U11681 (N_11681,N_11092,N_10631);
xnor U11682 (N_11682,N_10863,N_10873);
nand U11683 (N_11683,N_10934,N_11233);
or U11684 (N_11684,N_11065,N_11124);
xor U11685 (N_11685,N_10929,N_11112);
nand U11686 (N_11686,N_10627,N_10639);
or U11687 (N_11687,N_10691,N_11189);
xor U11688 (N_11688,N_10675,N_11090);
nor U11689 (N_11689,N_11118,N_10929);
nand U11690 (N_11690,N_11226,N_11196);
and U11691 (N_11691,N_10945,N_11066);
xnor U11692 (N_11692,N_10755,N_11036);
nor U11693 (N_11693,N_11111,N_10684);
and U11694 (N_11694,N_11249,N_10858);
or U11695 (N_11695,N_10706,N_11170);
nand U11696 (N_11696,N_11185,N_11193);
or U11697 (N_11697,N_11043,N_11102);
nor U11698 (N_11698,N_10658,N_11212);
xor U11699 (N_11699,N_10828,N_10700);
and U11700 (N_11700,N_10979,N_11115);
and U11701 (N_11701,N_11009,N_11108);
xnor U11702 (N_11702,N_10956,N_10625);
nand U11703 (N_11703,N_11005,N_10930);
nand U11704 (N_11704,N_10720,N_11236);
nor U11705 (N_11705,N_11248,N_11028);
and U11706 (N_11706,N_11179,N_10907);
and U11707 (N_11707,N_10818,N_10748);
xor U11708 (N_11708,N_10704,N_10720);
nor U11709 (N_11709,N_10695,N_11092);
nand U11710 (N_11710,N_11245,N_10725);
and U11711 (N_11711,N_10971,N_10888);
and U11712 (N_11712,N_10641,N_10873);
nor U11713 (N_11713,N_10768,N_10972);
or U11714 (N_11714,N_10659,N_10835);
or U11715 (N_11715,N_11248,N_11208);
and U11716 (N_11716,N_11245,N_10703);
nand U11717 (N_11717,N_10696,N_11146);
xor U11718 (N_11718,N_10721,N_11015);
and U11719 (N_11719,N_11207,N_11161);
nor U11720 (N_11720,N_10945,N_10889);
and U11721 (N_11721,N_10765,N_10718);
nand U11722 (N_11722,N_10925,N_11029);
and U11723 (N_11723,N_11115,N_10645);
xnor U11724 (N_11724,N_10950,N_10865);
xnor U11725 (N_11725,N_11022,N_11207);
or U11726 (N_11726,N_11013,N_10703);
and U11727 (N_11727,N_10999,N_10981);
nor U11728 (N_11728,N_10685,N_10790);
xnor U11729 (N_11729,N_10822,N_11153);
or U11730 (N_11730,N_10963,N_11046);
nor U11731 (N_11731,N_10983,N_11083);
nand U11732 (N_11732,N_11002,N_10629);
xnor U11733 (N_11733,N_11152,N_10652);
xor U11734 (N_11734,N_10875,N_11195);
or U11735 (N_11735,N_10792,N_10872);
and U11736 (N_11736,N_10909,N_10829);
and U11737 (N_11737,N_10828,N_11115);
nand U11738 (N_11738,N_11145,N_10629);
nor U11739 (N_11739,N_10915,N_10939);
and U11740 (N_11740,N_10813,N_11216);
nand U11741 (N_11741,N_10742,N_10853);
xor U11742 (N_11742,N_10829,N_10626);
nor U11743 (N_11743,N_11067,N_10726);
or U11744 (N_11744,N_11110,N_10895);
xor U11745 (N_11745,N_11035,N_10626);
xor U11746 (N_11746,N_10897,N_10649);
or U11747 (N_11747,N_10797,N_11002);
and U11748 (N_11748,N_10921,N_10812);
nand U11749 (N_11749,N_11187,N_11228);
nand U11750 (N_11750,N_11054,N_10784);
or U11751 (N_11751,N_11006,N_10805);
nand U11752 (N_11752,N_11075,N_10934);
or U11753 (N_11753,N_10845,N_11033);
nor U11754 (N_11754,N_11152,N_11138);
xnor U11755 (N_11755,N_10984,N_11132);
nor U11756 (N_11756,N_11101,N_10773);
or U11757 (N_11757,N_10950,N_10956);
xor U11758 (N_11758,N_10846,N_11166);
nand U11759 (N_11759,N_10745,N_10792);
nand U11760 (N_11760,N_10665,N_11198);
nand U11761 (N_11761,N_10664,N_10844);
nand U11762 (N_11762,N_10904,N_10684);
xnor U11763 (N_11763,N_10999,N_11127);
or U11764 (N_11764,N_11213,N_11013);
nor U11765 (N_11765,N_10641,N_10752);
nand U11766 (N_11766,N_10927,N_11182);
xnor U11767 (N_11767,N_10937,N_10715);
and U11768 (N_11768,N_10904,N_11026);
and U11769 (N_11769,N_10946,N_10978);
xor U11770 (N_11770,N_10692,N_10718);
nand U11771 (N_11771,N_10709,N_10998);
or U11772 (N_11772,N_11085,N_10667);
nand U11773 (N_11773,N_11242,N_11052);
nand U11774 (N_11774,N_10823,N_10745);
and U11775 (N_11775,N_11163,N_11236);
and U11776 (N_11776,N_11098,N_11144);
nand U11777 (N_11777,N_10646,N_10759);
xnor U11778 (N_11778,N_10691,N_11095);
nand U11779 (N_11779,N_11167,N_10876);
nor U11780 (N_11780,N_11193,N_10706);
xnor U11781 (N_11781,N_10888,N_11104);
nor U11782 (N_11782,N_10829,N_10673);
nor U11783 (N_11783,N_10883,N_10793);
or U11784 (N_11784,N_10719,N_11043);
or U11785 (N_11785,N_11015,N_11067);
or U11786 (N_11786,N_10869,N_10782);
and U11787 (N_11787,N_10878,N_10722);
or U11788 (N_11788,N_11044,N_11101);
nor U11789 (N_11789,N_11024,N_11025);
xor U11790 (N_11790,N_11078,N_11154);
or U11791 (N_11791,N_10728,N_10672);
xor U11792 (N_11792,N_11117,N_11109);
or U11793 (N_11793,N_11221,N_10776);
or U11794 (N_11794,N_10907,N_10705);
nand U11795 (N_11795,N_10689,N_11041);
nand U11796 (N_11796,N_10970,N_11081);
xnor U11797 (N_11797,N_10931,N_10734);
and U11798 (N_11798,N_10640,N_11229);
nor U11799 (N_11799,N_10726,N_10885);
or U11800 (N_11800,N_10853,N_11024);
xnor U11801 (N_11801,N_11005,N_10944);
nor U11802 (N_11802,N_10626,N_11232);
nand U11803 (N_11803,N_11242,N_10641);
nand U11804 (N_11804,N_11064,N_11179);
and U11805 (N_11805,N_10782,N_11190);
xor U11806 (N_11806,N_10730,N_11180);
nor U11807 (N_11807,N_11004,N_10953);
or U11808 (N_11808,N_10842,N_10857);
xor U11809 (N_11809,N_10655,N_10835);
and U11810 (N_11810,N_11143,N_10648);
xnor U11811 (N_11811,N_11125,N_11235);
and U11812 (N_11812,N_10973,N_11218);
and U11813 (N_11813,N_10908,N_10897);
nor U11814 (N_11814,N_10754,N_10902);
nand U11815 (N_11815,N_10633,N_10881);
nor U11816 (N_11816,N_10875,N_10648);
or U11817 (N_11817,N_10923,N_10649);
and U11818 (N_11818,N_11133,N_10685);
xor U11819 (N_11819,N_10952,N_10973);
and U11820 (N_11820,N_10763,N_11119);
nand U11821 (N_11821,N_11046,N_10843);
xor U11822 (N_11822,N_11214,N_11115);
and U11823 (N_11823,N_11238,N_11015);
nand U11824 (N_11824,N_10795,N_11247);
or U11825 (N_11825,N_11085,N_10914);
nand U11826 (N_11826,N_10960,N_11059);
nor U11827 (N_11827,N_11237,N_11061);
nand U11828 (N_11828,N_10966,N_10664);
xor U11829 (N_11829,N_11075,N_10857);
xor U11830 (N_11830,N_10982,N_11143);
xnor U11831 (N_11831,N_10759,N_11171);
nor U11832 (N_11832,N_10808,N_10928);
and U11833 (N_11833,N_10880,N_11074);
nand U11834 (N_11834,N_11001,N_11124);
nor U11835 (N_11835,N_11170,N_10727);
nand U11836 (N_11836,N_10678,N_10768);
and U11837 (N_11837,N_10784,N_11188);
nand U11838 (N_11838,N_10823,N_11115);
nand U11839 (N_11839,N_10754,N_11135);
xnor U11840 (N_11840,N_11152,N_11244);
nand U11841 (N_11841,N_11182,N_10830);
or U11842 (N_11842,N_11128,N_11154);
nor U11843 (N_11843,N_10795,N_10761);
and U11844 (N_11844,N_10839,N_11018);
and U11845 (N_11845,N_10912,N_11018);
xnor U11846 (N_11846,N_11135,N_10627);
or U11847 (N_11847,N_10955,N_10786);
nand U11848 (N_11848,N_11120,N_10759);
and U11849 (N_11849,N_11127,N_11100);
nand U11850 (N_11850,N_11166,N_10904);
xor U11851 (N_11851,N_11195,N_10820);
nor U11852 (N_11852,N_10626,N_11102);
nor U11853 (N_11853,N_10789,N_11130);
xnor U11854 (N_11854,N_11004,N_10934);
nor U11855 (N_11855,N_10861,N_11143);
xor U11856 (N_11856,N_11008,N_10900);
and U11857 (N_11857,N_11116,N_11213);
and U11858 (N_11858,N_10880,N_10706);
nand U11859 (N_11859,N_10668,N_10735);
xor U11860 (N_11860,N_10803,N_10826);
or U11861 (N_11861,N_11191,N_10720);
xor U11862 (N_11862,N_11051,N_11169);
xnor U11863 (N_11863,N_11187,N_10815);
or U11864 (N_11864,N_11171,N_11175);
nand U11865 (N_11865,N_10804,N_11079);
and U11866 (N_11866,N_10986,N_10866);
or U11867 (N_11867,N_10693,N_10678);
or U11868 (N_11868,N_10685,N_10923);
nand U11869 (N_11869,N_10712,N_10788);
or U11870 (N_11870,N_10666,N_11061);
and U11871 (N_11871,N_11124,N_10834);
or U11872 (N_11872,N_10679,N_11239);
or U11873 (N_11873,N_11202,N_11052);
or U11874 (N_11874,N_10850,N_11246);
nor U11875 (N_11875,N_11320,N_11504);
nand U11876 (N_11876,N_11479,N_11614);
nor U11877 (N_11877,N_11756,N_11720);
nand U11878 (N_11878,N_11390,N_11535);
nor U11879 (N_11879,N_11587,N_11676);
and U11880 (N_11880,N_11690,N_11509);
xor U11881 (N_11881,N_11409,N_11555);
or U11882 (N_11882,N_11495,N_11422);
nand U11883 (N_11883,N_11760,N_11499);
nand U11884 (N_11884,N_11519,N_11704);
nand U11885 (N_11885,N_11867,N_11685);
nand U11886 (N_11886,N_11385,N_11287);
nand U11887 (N_11887,N_11295,N_11682);
nor U11888 (N_11888,N_11700,N_11590);
nor U11889 (N_11889,N_11612,N_11828);
or U11890 (N_11890,N_11696,N_11799);
or U11891 (N_11891,N_11838,N_11808);
nand U11892 (N_11892,N_11692,N_11553);
nor U11893 (N_11893,N_11837,N_11669);
or U11894 (N_11894,N_11251,N_11839);
xor U11895 (N_11895,N_11402,N_11841);
and U11896 (N_11896,N_11269,N_11467);
or U11897 (N_11897,N_11259,N_11742);
xor U11898 (N_11898,N_11528,N_11683);
nand U11899 (N_11899,N_11771,N_11851);
and U11900 (N_11900,N_11842,N_11818);
and U11901 (N_11901,N_11591,N_11434);
nor U11902 (N_11902,N_11770,N_11399);
nand U11903 (N_11903,N_11373,N_11543);
and U11904 (N_11904,N_11462,N_11747);
xor U11905 (N_11905,N_11500,N_11740);
xor U11906 (N_11906,N_11581,N_11400);
or U11907 (N_11907,N_11381,N_11632);
xnor U11908 (N_11908,N_11463,N_11252);
xnor U11909 (N_11909,N_11755,N_11365);
xor U11910 (N_11910,N_11386,N_11480);
nand U11911 (N_11911,N_11477,N_11537);
or U11912 (N_11912,N_11255,N_11435);
xnor U11913 (N_11913,N_11393,N_11303);
or U11914 (N_11914,N_11860,N_11536);
and U11915 (N_11915,N_11757,N_11336);
and U11916 (N_11916,N_11677,N_11680);
or U11917 (N_11917,N_11501,N_11557);
nand U11918 (N_11918,N_11774,N_11579);
nor U11919 (N_11919,N_11453,N_11471);
nand U11920 (N_11920,N_11585,N_11331);
xnor U11921 (N_11921,N_11340,N_11468);
or U11922 (N_11922,N_11382,N_11461);
xnor U11923 (N_11923,N_11807,N_11650);
or U11924 (N_11924,N_11780,N_11298);
nor U11925 (N_11925,N_11718,N_11263);
nand U11926 (N_11926,N_11737,N_11550);
nor U11927 (N_11927,N_11337,N_11518);
or U11928 (N_11928,N_11449,N_11835);
nor U11929 (N_11929,N_11754,N_11523);
nand U11930 (N_11930,N_11710,N_11717);
nand U11931 (N_11931,N_11431,N_11634);
or U11932 (N_11932,N_11378,N_11432);
and U11933 (N_11933,N_11485,N_11670);
xnor U11934 (N_11934,N_11547,N_11641);
nor U11935 (N_11935,N_11299,N_11450);
nor U11936 (N_11936,N_11749,N_11744);
nand U11937 (N_11937,N_11443,N_11483);
xnor U11938 (N_11938,N_11711,N_11286);
nand U11939 (N_11939,N_11625,N_11761);
xor U11940 (N_11940,N_11629,N_11630);
or U11941 (N_11941,N_11530,N_11618);
and U11942 (N_11942,N_11636,N_11622);
nor U11943 (N_11943,N_11396,N_11723);
nor U11944 (N_11944,N_11486,N_11338);
xnor U11945 (N_11945,N_11638,N_11440);
xor U11946 (N_11946,N_11810,N_11308);
nand U11947 (N_11947,N_11502,N_11652);
xor U11948 (N_11948,N_11665,N_11476);
nor U11949 (N_11949,N_11640,N_11473);
nor U11950 (N_11950,N_11532,N_11408);
or U11951 (N_11951,N_11350,N_11273);
or U11952 (N_11952,N_11349,N_11376);
nor U11953 (N_11953,N_11375,N_11601);
or U11954 (N_11954,N_11291,N_11578);
nor U11955 (N_11955,N_11290,N_11297);
or U11956 (N_11956,N_11539,N_11455);
and U11957 (N_11957,N_11448,N_11369);
or U11958 (N_11958,N_11507,N_11554);
and U11959 (N_11959,N_11538,N_11441);
nand U11960 (N_11960,N_11617,N_11713);
xor U11961 (N_11961,N_11564,N_11731);
nor U11962 (N_11962,N_11663,N_11478);
nand U11963 (N_11963,N_11793,N_11459);
or U11964 (N_11964,N_11866,N_11791);
xnor U11965 (N_11965,N_11488,N_11384);
or U11966 (N_11966,N_11289,N_11417);
or U11967 (N_11967,N_11420,N_11758);
and U11968 (N_11968,N_11332,N_11442);
nor U11969 (N_11969,N_11566,N_11454);
nor U11970 (N_11970,N_11616,N_11546);
xor U11971 (N_11971,N_11412,N_11275);
and U11972 (N_11972,N_11645,N_11366);
xnor U11973 (N_11973,N_11265,N_11266);
or U11974 (N_11974,N_11796,N_11274);
or U11975 (N_11975,N_11258,N_11701);
nand U11976 (N_11976,N_11664,N_11284);
and U11977 (N_11977,N_11626,N_11869);
or U11978 (N_11978,N_11847,N_11805);
nand U11979 (N_11979,N_11458,N_11716);
and U11980 (N_11980,N_11631,N_11678);
nand U11981 (N_11981,N_11597,N_11447);
nor U11982 (N_11982,N_11773,N_11768);
xnor U11983 (N_11983,N_11753,N_11688);
or U11984 (N_11984,N_11864,N_11580);
or U11985 (N_11985,N_11611,N_11766);
nor U11986 (N_11986,N_11310,N_11671);
nor U11987 (N_11987,N_11725,N_11426);
or U11988 (N_11988,N_11620,N_11328);
nor U11989 (N_11989,N_11655,N_11673);
nand U11990 (N_11990,N_11732,N_11484);
nand U11991 (N_11991,N_11356,N_11281);
nor U11992 (N_11992,N_11806,N_11345);
and U11993 (N_11993,N_11481,N_11826);
nand U11994 (N_11994,N_11307,N_11822);
and U11995 (N_11995,N_11323,N_11668);
and U11996 (N_11996,N_11691,N_11594);
and U11997 (N_11997,N_11389,N_11750);
or U11998 (N_11998,N_11639,N_11599);
and U11999 (N_11999,N_11863,N_11293);
or U12000 (N_12000,N_11829,N_11413);
or U12001 (N_12001,N_11784,N_11868);
nor U12002 (N_12002,N_11741,N_11470);
nor U12003 (N_12003,N_11661,N_11817);
and U12004 (N_12004,N_11746,N_11445);
or U12005 (N_12005,N_11406,N_11552);
nor U12006 (N_12006,N_11407,N_11311);
xor U12007 (N_12007,N_11354,N_11637);
and U12008 (N_12008,N_11735,N_11598);
and U12009 (N_12009,N_11346,N_11823);
xor U12010 (N_12010,N_11548,N_11832);
nand U12011 (N_12011,N_11493,N_11794);
nor U12012 (N_12012,N_11268,N_11380);
xnor U12013 (N_12013,N_11658,N_11633);
nor U12014 (N_12014,N_11861,N_11526);
xor U12015 (N_12015,N_11352,N_11871);
nor U12016 (N_12016,N_11410,N_11743);
nor U12017 (N_12017,N_11306,N_11709);
nand U12018 (N_12018,N_11279,N_11474);
nand U12019 (N_12019,N_11466,N_11423);
nand U12020 (N_12020,N_11497,N_11586);
nor U12021 (N_12021,N_11475,N_11438);
or U12022 (N_12022,N_11648,N_11825);
xor U12023 (N_12023,N_11778,N_11315);
nor U12024 (N_12024,N_11790,N_11403);
xor U12025 (N_12025,N_11460,N_11524);
and U12026 (N_12026,N_11595,N_11419);
and U12027 (N_12027,N_11271,N_11421);
and U12028 (N_12028,N_11584,N_11856);
nand U12029 (N_12029,N_11785,N_11533);
nand U12030 (N_12030,N_11304,N_11635);
or U12031 (N_12031,N_11556,N_11362);
xnor U12032 (N_12032,N_11496,N_11660);
and U12033 (N_12033,N_11261,N_11583);
nor U12034 (N_12034,N_11401,N_11721);
nor U12035 (N_12035,N_11646,N_11571);
xor U12036 (N_12036,N_11656,N_11605);
nor U12037 (N_12037,N_11589,N_11264);
xor U12038 (N_12038,N_11347,N_11292);
nor U12039 (N_12039,N_11322,N_11254);
xnor U12040 (N_12040,N_11859,N_11464);
nor U12041 (N_12041,N_11674,N_11836);
nand U12042 (N_12042,N_11679,N_11510);
xor U12043 (N_12043,N_11814,N_11301);
xnor U12044 (N_12044,N_11621,N_11714);
and U12045 (N_12045,N_11873,N_11697);
xnor U12046 (N_12046,N_11831,N_11313);
nor U12047 (N_12047,N_11738,N_11703);
nor U12048 (N_12048,N_11699,N_11613);
or U12049 (N_12049,N_11573,N_11804);
nor U12050 (N_12050,N_11657,N_11514);
nor U12051 (N_12051,N_11416,N_11763);
and U12052 (N_12052,N_11736,N_11428);
xor U12053 (N_12053,N_11801,N_11772);
nand U12054 (N_12054,N_11730,N_11798);
nor U12055 (N_12055,N_11512,N_11364);
nand U12056 (N_12056,N_11803,N_11858);
nand U12057 (N_12057,N_11372,N_11374);
nand U12058 (N_12058,N_11527,N_11853);
or U12059 (N_12059,N_11394,N_11276);
nand U12060 (N_12060,N_11329,N_11250);
nor U12061 (N_12061,N_11334,N_11800);
or U12062 (N_12062,N_11494,N_11764);
nor U12063 (N_12063,N_11786,N_11872);
and U12064 (N_12064,N_11387,N_11333);
nor U12065 (N_12065,N_11371,N_11845);
and U12066 (N_12066,N_11324,N_11309);
xor U12067 (N_12067,N_11659,N_11294);
or U12068 (N_12068,N_11582,N_11686);
xnor U12069 (N_12069,N_11253,N_11545);
xnor U12070 (N_12070,N_11405,N_11698);
nor U12071 (N_12071,N_11516,N_11377);
and U12072 (N_12072,N_11865,N_11843);
or U12073 (N_12073,N_11498,N_11672);
nand U12074 (N_12074,N_11429,N_11862);
nor U12075 (N_12075,N_11812,N_11588);
nand U12076 (N_12076,N_11469,N_11642);
xnor U12077 (N_12077,N_11577,N_11813);
or U12078 (N_12078,N_11348,N_11568);
nor U12079 (N_12079,N_11318,N_11517);
xor U12080 (N_12080,N_11848,N_11596);
or U12081 (N_12081,N_11561,N_11465);
xnor U12082 (N_12082,N_11327,N_11722);
nor U12083 (N_12083,N_11726,N_11529);
or U12084 (N_12084,N_11833,N_11285);
nand U12085 (N_12085,N_11733,N_11600);
or U12086 (N_12086,N_11654,N_11855);
xnor U12087 (N_12087,N_11857,N_11451);
nor U12088 (N_12088,N_11525,N_11675);
nor U12089 (N_12089,N_11569,N_11724);
and U12090 (N_12090,N_11567,N_11344);
and U12091 (N_12091,N_11357,N_11361);
nor U12092 (N_12092,N_11715,N_11558);
nand U12093 (N_12093,N_11565,N_11358);
nor U12094 (N_12094,N_11487,N_11824);
nand U12095 (N_12095,N_11430,N_11751);
xnor U12096 (N_12096,N_11662,N_11270);
or U12097 (N_12097,N_11513,N_11752);
nand U12098 (N_12098,N_11607,N_11531);
nor U12099 (N_12099,N_11574,N_11491);
xnor U12100 (N_12100,N_11604,N_11643);
and U12101 (N_12101,N_11395,N_11830);
or U12102 (N_12102,N_11762,N_11319);
and U12103 (N_12103,N_11615,N_11572);
or U12104 (N_12104,N_11544,N_11728);
nor U12105 (N_12105,N_11666,N_11541);
xor U12106 (N_12106,N_11777,N_11489);
or U12107 (N_12107,N_11282,N_11719);
nand U12108 (N_12108,N_11379,N_11549);
nand U12109 (N_12109,N_11388,N_11262);
or U12110 (N_12110,N_11667,N_11705);
or U12111 (N_12111,N_11782,N_11300);
xor U12112 (N_12112,N_11456,N_11397);
nor U12113 (N_12113,N_11602,N_11418);
nor U12114 (N_12114,N_11424,N_11515);
xnor U12115 (N_12115,N_11444,N_11706);
or U12116 (N_12116,N_11505,N_11776);
and U12117 (N_12117,N_11606,N_11272);
xnor U12118 (N_12118,N_11288,N_11277);
or U12119 (N_12119,N_11404,N_11819);
nand U12120 (N_12120,N_11427,N_11343);
and U12121 (N_12121,N_11702,N_11849);
nor U12122 (N_12122,N_11789,N_11436);
or U12123 (N_12123,N_11425,N_11694);
and U12124 (N_12124,N_11792,N_11734);
and U12125 (N_12125,N_11852,N_11283);
and U12126 (N_12126,N_11326,N_11781);
nand U12127 (N_12127,N_11437,N_11748);
nor U12128 (N_12128,N_11593,N_11653);
and U12129 (N_12129,N_11339,N_11854);
or U12130 (N_12130,N_11844,N_11727);
nand U12131 (N_12131,N_11821,N_11840);
or U12132 (N_12132,N_11576,N_11610);
and U12133 (N_12133,N_11560,N_11712);
and U12134 (N_12134,N_11609,N_11511);
nand U12135 (N_12135,N_11452,N_11870);
and U12136 (N_12136,N_11503,N_11363);
nor U12137 (N_12137,N_11439,N_11341);
nand U12138 (N_12138,N_11522,N_11759);
xnor U12139 (N_12139,N_11797,N_11570);
xor U12140 (N_12140,N_11280,N_11472);
nand U12141 (N_12141,N_11787,N_11695);
and U12142 (N_12142,N_11342,N_11708);
nand U12143 (N_12143,N_11827,N_11351);
nand U12144 (N_12144,N_11765,N_11260);
nor U12145 (N_12145,N_11302,N_11739);
nor U12146 (N_12146,N_11411,N_11335);
nor U12147 (N_12147,N_11834,N_11359);
nor U12148 (N_12148,N_11330,N_11520);
xnor U12149 (N_12149,N_11257,N_11296);
nand U12150 (N_12150,N_11779,N_11325);
nand U12151 (N_12151,N_11534,N_11383);
nand U12152 (N_12152,N_11820,N_11769);
or U12153 (N_12153,N_11391,N_11370);
nand U12154 (N_12154,N_11767,N_11551);
and U12155 (N_12155,N_11415,N_11414);
nand U12156 (N_12156,N_11729,N_11603);
xnor U12157 (N_12157,N_11684,N_11278);
nand U12158 (N_12158,N_11317,N_11355);
nor U12159 (N_12159,N_11267,N_11809);
nand U12160 (N_12160,N_11256,N_11681);
xor U12161 (N_12161,N_11540,N_11795);
xor U12162 (N_12162,N_11563,N_11647);
or U12163 (N_12163,N_11628,N_11689);
nand U12164 (N_12164,N_11687,N_11811);
nand U12165 (N_12165,N_11562,N_11649);
or U12166 (N_12166,N_11316,N_11745);
or U12167 (N_12167,N_11398,N_11623);
nor U12168 (N_12168,N_11433,N_11592);
nor U12169 (N_12169,N_11624,N_11846);
or U12170 (N_12170,N_11368,N_11321);
xnor U12171 (N_12171,N_11312,N_11693);
or U12172 (N_12172,N_11575,N_11775);
or U12173 (N_12173,N_11521,N_11707);
or U12174 (N_12174,N_11353,N_11627);
xor U12175 (N_12175,N_11314,N_11788);
nand U12176 (N_12176,N_11457,N_11850);
nor U12177 (N_12177,N_11305,N_11360);
xor U12178 (N_12178,N_11815,N_11816);
nand U12179 (N_12179,N_11619,N_11559);
nand U12180 (N_12180,N_11482,N_11644);
nor U12181 (N_12181,N_11783,N_11608);
nand U12182 (N_12182,N_11802,N_11506);
nand U12183 (N_12183,N_11542,N_11651);
and U12184 (N_12184,N_11492,N_11446);
nand U12185 (N_12185,N_11490,N_11874);
nand U12186 (N_12186,N_11392,N_11367);
nand U12187 (N_12187,N_11508,N_11744);
or U12188 (N_12188,N_11874,N_11747);
or U12189 (N_12189,N_11768,N_11498);
and U12190 (N_12190,N_11493,N_11388);
or U12191 (N_12191,N_11785,N_11278);
xor U12192 (N_12192,N_11846,N_11418);
and U12193 (N_12193,N_11738,N_11635);
and U12194 (N_12194,N_11500,N_11537);
or U12195 (N_12195,N_11806,N_11855);
nand U12196 (N_12196,N_11568,N_11801);
xnor U12197 (N_12197,N_11510,N_11560);
xnor U12198 (N_12198,N_11532,N_11528);
nand U12199 (N_12199,N_11375,N_11763);
nor U12200 (N_12200,N_11674,N_11786);
and U12201 (N_12201,N_11447,N_11594);
nor U12202 (N_12202,N_11421,N_11331);
and U12203 (N_12203,N_11530,N_11511);
and U12204 (N_12204,N_11703,N_11798);
nor U12205 (N_12205,N_11757,N_11405);
nor U12206 (N_12206,N_11541,N_11856);
nand U12207 (N_12207,N_11753,N_11789);
nor U12208 (N_12208,N_11304,N_11751);
and U12209 (N_12209,N_11776,N_11307);
and U12210 (N_12210,N_11531,N_11815);
or U12211 (N_12211,N_11274,N_11442);
and U12212 (N_12212,N_11308,N_11578);
nor U12213 (N_12213,N_11830,N_11354);
nor U12214 (N_12214,N_11799,N_11602);
xor U12215 (N_12215,N_11737,N_11482);
and U12216 (N_12216,N_11736,N_11274);
xor U12217 (N_12217,N_11324,N_11640);
and U12218 (N_12218,N_11461,N_11437);
or U12219 (N_12219,N_11552,N_11667);
and U12220 (N_12220,N_11498,N_11540);
or U12221 (N_12221,N_11264,N_11279);
xnor U12222 (N_12222,N_11659,N_11831);
or U12223 (N_12223,N_11561,N_11861);
xnor U12224 (N_12224,N_11575,N_11655);
and U12225 (N_12225,N_11296,N_11400);
xnor U12226 (N_12226,N_11617,N_11451);
nand U12227 (N_12227,N_11634,N_11437);
xnor U12228 (N_12228,N_11346,N_11604);
and U12229 (N_12229,N_11549,N_11372);
nand U12230 (N_12230,N_11501,N_11695);
xnor U12231 (N_12231,N_11567,N_11622);
nor U12232 (N_12232,N_11575,N_11273);
xor U12233 (N_12233,N_11795,N_11665);
nand U12234 (N_12234,N_11795,N_11598);
xor U12235 (N_12235,N_11555,N_11502);
xor U12236 (N_12236,N_11266,N_11610);
xnor U12237 (N_12237,N_11637,N_11604);
nor U12238 (N_12238,N_11788,N_11406);
nor U12239 (N_12239,N_11545,N_11740);
nor U12240 (N_12240,N_11821,N_11587);
and U12241 (N_12241,N_11627,N_11403);
nor U12242 (N_12242,N_11311,N_11639);
and U12243 (N_12243,N_11497,N_11830);
nor U12244 (N_12244,N_11349,N_11486);
or U12245 (N_12245,N_11573,N_11312);
nand U12246 (N_12246,N_11388,N_11420);
and U12247 (N_12247,N_11729,N_11333);
nor U12248 (N_12248,N_11538,N_11607);
and U12249 (N_12249,N_11630,N_11759);
xor U12250 (N_12250,N_11763,N_11702);
and U12251 (N_12251,N_11579,N_11310);
xor U12252 (N_12252,N_11626,N_11646);
xor U12253 (N_12253,N_11323,N_11609);
xnor U12254 (N_12254,N_11718,N_11814);
xnor U12255 (N_12255,N_11286,N_11548);
nor U12256 (N_12256,N_11409,N_11490);
nand U12257 (N_12257,N_11594,N_11841);
xnor U12258 (N_12258,N_11677,N_11440);
xnor U12259 (N_12259,N_11749,N_11699);
and U12260 (N_12260,N_11708,N_11662);
nor U12261 (N_12261,N_11401,N_11628);
and U12262 (N_12262,N_11479,N_11525);
nand U12263 (N_12263,N_11800,N_11550);
nor U12264 (N_12264,N_11763,N_11798);
xor U12265 (N_12265,N_11260,N_11796);
nand U12266 (N_12266,N_11873,N_11432);
xnor U12267 (N_12267,N_11610,N_11465);
xnor U12268 (N_12268,N_11394,N_11630);
nand U12269 (N_12269,N_11377,N_11586);
xor U12270 (N_12270,N_11481,N_11330);
xor U12271 (N_12271,N_11539,N_11272);
and U12272 (N_12272,N_11805,N_11769);
or U12273 (N_12273,N_11766,N_11851);
and U12274 (N_12274,N_11445,N_11434);
nand U12275 (N_12275,N_11509,N_11844);
or U12276 (N_12276,N_11753,N_11435);
nand U12277 (N_12277,N_11835,N_11613);
or U12278 (N_12278,N_11739,N_11345);
and U12279 (N_12279,N_11443,N_11694);
or U12280 (N_12280,N_11699,N_11744);
or U12281 (N_12281,N_11464,N_11810);
nor U12282 (N_12282,N_11819,N_11851);
nor U12283 (N_12283,N_11699,N_11820);
nand U12284 (N_12284,N_11860,N_11824);
and U12285 (N_12285,N_11466,N_11294);
nor U12286 (N_12286,N_11386,N_11846);
xor U12287 (N_12287,N_11716,N_11708);
nand U12288 (N_12288,N_11562,N_11287);
xor U12289 (N_12289,N_11577,N_11572);
nand U12290 (N_12290,N_11753,N_11260);
nor U12291 (N_12291,N_11395,N_11475);
or U12292 (N_12292,N_11369,N_11294);
xnor U12293 (N_12293,N_11689,N_11333);
or U12294 (N_12294,N_11548,N_11337);
or U12295 (N_12295,N_11377,N_11269);
xor U12296 (N_12296,N_11306,N_11412);
and U12297 (N_12297,N_11863,N_11565);
and U12298 (N_12298,N_11256,N_11335);
or U12299 (N_12299,N_11657,N_11540);
nor U12300 (N_12300,N_11504,N_11614);
xnor U12301 (N_12301,N_11669,N_11294);
nand U12302 (N_12302,N_11507,N_11539);
or U12303 (N_12303,N_11324,N_11549);
and U12304 (N_12304,N_11671,N_11526);
nand U12305 (N_12305,N_11672,N_11466);
or U12306 (N_12306,N_11328,N_11628);
and U12307 (N_12307,N_11346,N_11442);
nand U12308 (N_12308,N_11645,N_11670);
and U12309 (N_12309,N_11603,N_11515);
or U12310 (N_12310,N_11506,N_11495);
or U12311 (N_12311,N_11325,N_11730);
xnor U12312 (N_12312,N_11814,N_11357);
nand U12313 (N_12313,N_11315,N_11264);
nand U12314 (N_12314,N_11703,N_11812);
nor U12315 (N_12315,N_11716,N_11424);
xnor U12316 (N_12316,N_11835,N_11619);
nor U12317 (N_12317,N_11411,N_11622);
nand U12318 (N_12318,N_11307,N_11330);
nor U12319 (N_12319,N_11741,N_11568);
or U12320 (N_12320,N_11293,N_11724);
and U12321 (N_12321,N_11346,N_11613);
or U12322 (N_12322,N_11278,N_11292);
or U12323 (N_12323,N_11833,N_11761);
and U12324 (N_12324,N_11695,N_11604);
and U12325 (N_12325,N_11730,N_11615);
xor U12326 (N_12326,N_11429,N_11378);
nor U12327 (N_12327,N_11755,N_11579);
nor U12328 (N_12328,N_11794,N_11337);
nand U12329 (N_12329,N_11376,N_11355);
nor U12330 (N_12330,N_11251,N_11488);
xnor U12331 (N_12331,N_11404,N_11520);
and U12332 (N_12332,N_11316,N_11286);
nand U12333 (N_12333,N_11445,N_11567);
nor U12334 (N_12334,N_11342,N_11436);
and U12335 (N_12335,N_11367,N_11818);
nor U12336 (N_12336,N_11758,N_11689);
xor U12337 (N_12337,N_11523,N_11820);
or U12338 (N_12338,N_11502,N_11675);
xor U12339 (N_12339,N_11449,N_11374);
and U12340 (N_12340,N_11801,N_11623);
nor U12341 (N_12341,N_11866,N_11338);
nand U12342 (N_12342,N_11546,N_11781);
or U12343 (N_12343,N_11528,N_11710);
and U12344 (N_12344,N_11796,N_11715);
and U12345 (N_12345,N_11736,N_11794);
xnor U12346 (N_12346,N_11857,N_11736);
or U12347 (N_12347,N_11669,N_11319);
nor U12348 (N_12348,N_11741,N_11570);
xnor U12349 (N_12349,N_11629,N_11855);
xor U12350 (N_12350,N_11446,N_11536);
nor U12351 (N_12351,N_11551,N_11399);
nor U12352 (N_12352,N_11562,N_11811);
and U12353 (N_12353,N_11662,N_11807);
nand U12354 (N_12354,N_11394,N_11355);
nor U12355 (N_12355,N_11836,N_11766);
nor U12356 (N_12356,N_11806,N_11723);
xor U12357 (N_12357,N_11543,N_11323);
or U12358 (N_12358,N_11389,N_11483);
nor U12359 (N_12359,N_11717,N_11701);
or U12360 (N_12360,N_11619,N_11272);
nand U12361 (N_12361,N_11544,N_11530);
nor U12362 (N_12362,N_11701,N_11612);
nor U12363 (N_12363,N_11375,N_11706);
nor U12364 (N_12364,N_11814,N_11617);
and U12365 (N_12365,N_11832,N_11328);
xor U12366 (N_12366,N_11265,N_11567);
or U12367 (N_12367,N_11361,N_11646);
and U12368 (N_12368,N_11717,N_11619);
and U12369 (N_12369,N_11806,N_11703);
nor U12370 (N_12370,N_11259,N_11862);
xnor U12371 (N_12371,N_11729,N_11859);
or U12372 (N_12372,N_11322,N_11580);
and U12373 (N_12373,N_11512,N_11253);
or U12374 (N_12374,N_11811,N_11873);
nand U12375 (N_12375,N_11691,N_11410);
nor U12376 (N_12376,N_11416,N_11646);
nand U12377 (N_12377,N_11407,N_11686);
and U12378 (N_12378,N_11310,N_11741);
and U12379 (N_12379,N_11839,N_11493);
xor U12380 (N_12380,N_11525,N_11262);
xor U12381 (N_12381,N_11335,N_11321);
nand U12382 (N_12382,N_11255,N_11560);
nor U12383 (N_12383,N_11534,N_11435);
nand U12384 (N_12384,N_11436,N_11515);
nor U12385 (N_12385,N_11717,N_11394);
nand U12386 (N_12386,N_11403,N_11502);
and U12387 (N_12387,N_11820,N_11819);
nand U12388 (N_12388,N_11436,N_11373);
nand U12389 (N_12389,N_11782,N_11289);
xnor U12390 (N_12390,N_11292,N_11332);
or U12391 (N_12391,N_11684,N_11422);
xnor U12392 (N_12392,N_11421,N_11395);
and U12393 (N_12393,N_11624,N_11605);
or U12394 (N_12394,N_11802,N_11650);
nor U12395 (N_12395,N_11283,N_11575);
xnor U12396 (N_12396,N_11722,N_11334);
nor U12397 (N_12397,N_11414,N_11285);
nand U12398 (N_12398,N_11347,N_11630);
nand U12399 (N_12399,N_11340,N_11409);
and U12400 (N_12400,N_11412,N_11616);
xnor U12401 (N_12401,N_11792,N_11694);
nor U12402 (N_12402,N_11760,N_11618);
or U12403 (N_12403,N_11402,N_11251);
and U12404 (N_12404,N_11613,N_11505);
or U12405 (N_12405,N_11286,N_11363);
and U12406 (N_12406,N_11457,N_11383);
or U12407 (N_12407,N_11684,N_11660);
nor U12408 (N_12408,N_11414,N_11273);
xnor U12409 (N_12409,N_11552,N_11585);
or U12410 (N_12410,N_11471,N_11871);
nand U12411 (N_12411,N_11706,N_11286);
nand U12412 (N_12412,N_11541,N_11754);
nand U12413 (N_12413,N_11656,N_11681);
and U12414 (N_12414,N_11297,N_11755);
nor U12415 (N_12415,N_11335,N_11866);
nor U12416 (N_12416,N_11681,N_11666);
nor U12417 (N_12417,N_11601,N_11360);
and U12418 (N_12418,N_11625,N_11294);
xor U12419 (N_12419,N_11545,N_11275);
or U12420 (N_12420,N_11606,N_11402);
or U12421 (N_12421,N_11525,N_11312);
nor U12422 (N_12422,N_11839,N_11564);
and U12423 (N_12423,N_11385,N_11387);
nand U12424 (N_12424,N_11681,N_11648);
and U12425 (N_12425,N_11849,N_11863);
nand U12426 (N_12426,N_11552,N_11260);
nor U12427 (N_12427,N_11658,N_11366);
or U12428 (N_12428,N_11556,N_11414);
nand U12429 (N_12429,N_11626,N_11611);
or U12430 (N_12430,N_11522,N_11504);
or U12431 (N_12431,N_11467,N_11383);
nand U12432 (N_12432,N_11471,N_11513);
or U12433 (N_12433,N_11637,N_11855);
and U12434 (N_12434,N_11352,N_11294);
xnor U12435 (N_12435,N_11699,N_11634);
nand U12436 (N_12436,N_11732,N_11740);
or U12437 (N_12437,N_11625,N_11714);
or U12438 (N_12438,N_11607,N_11632);
and U12439 (N_12439,N_11252,N_11488);
nand U12440 (N_12440,N_11481,N_11762);
and U12441 (N_12441,N_11640,N_11691);
nor U12442 (N_12442,N_11499,N_11810);
or U12443 (N_12443,N_11647,N_11789);
and U12444 (N_12444,N_11393,N_11720);
nand U12445 (N_12445,N_11297,N_11551);
xnor U12446 (N_12446,N_11452,N_11855);
nand U12447 (N_12447,N_11706,N_11317);
nand U12448 (N_12448,N_11449,N_11486);
xor U12449 (N_12449,N_11558,N_11732);
and U12450 (N_12450,N_11466,N_11867);
xor U12451 (N_12451,N_11799,N_11743);
nand U12452 (N_12452,N_11261,N_11351);
xor U12453 (N_12453,N_11772,N_11536);
nor U12454 (N_12454,N_11503,N_11619);
or U12455 (N_12455,N_11672,N_11394);
or U12456 (N_12456,N_11688,N_11404);
nand U12457 (N_12457,N_11805,N_11466);
or U12458 (N_12458,N_11261,N_11438);
and U12459 (N_12459,N_11302,N_11743);
and U12460 (N_12460,N_11579,N_11779);
xor U12461 (N_12461,N_11751,N_11463);
xnor U12462 (N_12462,N_11684,N_11336);
nor U12463 (N_12463,N_11741,N_11803);
nand U12464 (N_12464,N_11422,N_11861);
nand U12465 (N_12465,N_11586,N_11388);
nand U12466 (N_12466,N_11485,N_11405);
or U12467 (N_12467,N_11423,N_11381);
nor U12468 (N_12468,N_11713,N_11305);
nor U12469 (N_12469,N_11523,N_11840);
and U12470 (N_12470,N_11508,N_11835);
or U12471 (N_12471,N_11465,N_11382);
and U12472 (N_12472,N_11663,N_11502);
xor U12473 (N_12473,N_11457,N_11571);
or U12474 (N_12474,N_11263,N_11341);
nor U12475 (N_12475,N_11747,N_11825);
nor U12476 (N_12476,N_11332,N_11737);
and U12477 (N_12477,N_11600,N_11665);
and U12478 (N_12478,N_11768,N_11300);
and U12479 (N_12479,N_11766,N_11347);
and U12480 (N_12480,N_11666,N_11872);
nor U12481 (N_12481,N_11628,N_11666);
or U12482 (N_12482,N_11275,N_11252);
and U12483 (N_12483,N_11638,N_11329);
and U12484 (N_12484,N_11691,N_11438);
nor U12485 (N_12485,N_11816,N_11648);
nand U12486 (N_12486,N_11655,N_11727);
nand U12487 (N_12487,N_11456,N_11594);
nor U12488 (N_12488,N_11537,N_11666);
nand U12489 (N_12489,N_11376,N_11793);
nand U12490 (N_12490,N_11329,N_11528);
or U12491 (N_12491,N_11373,N_11499);
xnor U12492 (N_12492,N_11725,N_11486);
or U12493 (N_12493,N_11716,N_11797);
nor U12494 (N_12494,N_11279,N_11680);
xor U12495 (N_12495,N_11549,N_11500);
nor U12496 (N_12496,N_11413,N_11651);
or U12497 (N_12497,N_11515,N_11365);
xnor U12498 (N_12498,N_11558,N_11365);
nor U12499 (N_12499,N_11813,N_11740);
nor U12500 (N_12500,N_12000,N_12336);
xnor U12501 (N_12501,N_11887,N_12278);
xnor U12502 (N_12502,N_12457,N_12391);
xor U12503 (N_12503,N_12004,N_12006);
or U12504 (N_12504,N_12306,N_12129);
nor U12505 (N_12505,N_12413,N_12031);
and U12506 (N_12506,N_12025,N_12137);
nand U12507 (N_12507,N_12262,N_12076);
nor U12508 (N_12508,N_12140,N_11909);
xnor U12509 (N_12509,N_12467,N_11939);
nor U12510 (N_12510,N_11943,N_12444);
or U12511 (N_12511,N_11901,N_12373);
nor U12512 (N_12512,N_12052,N_12464);
nor U12513 (N_12513,N_12169,N_11989);
xnor U12514 (N_12514,N_12282,N_12481);
or U12515 (N_12515,N_12497,N_12327);
nor U12516 (N_12516,N_12427,N_11885);
or U12517 (N_12517,N_12168,N_12133);
and U12518 (N_12518,N_11950,N_12329);
or U12519 (N_12519,N_12287,N_11875);
nand U12520 (N_12520,N_12423,N_12355);
and U12521 (N_12521,N_12007,N_12390);
nand U12522 (N_12522,N_12115,N_12079);
nand U12523 (N_12523,N_12482,N_12171);
xnor U12524 (N_12524,N_12305,N_12339);
or U12525 (N_12525,N_11929,N_12178);
nor U12526 (N_12526,N_12246,N_12280);
nand U12527 (N_12527,N_12298,N_12323);
xnor U12528 (N_12528,N_11888,N_12376);
xnor U12529 (N_12529,N_12063,N_12008);
or U12530 (N_12530,N_11930,N_12107);
or U12531 (N_12531,N_12307,N_11990);
xnor U12532 (N_12532,N_12462,N_12130);
xor U12533 (N_12533,N_12114,N_11899);
xor U12534 (N_12534,N_12494,N_12225);
nand U12535 (N_12535,N_12453,N_12082);
nand U12536 (N_12536,N_12147,N_12012);
nand U12537 (N_12537,N_12197,N_12117);
nor U12538 (N_12538,N_12222,N_12402);
nand U12539 (N_12539,N_12394,N_12264);
xor U12540 (N_12540,N_12439,N_12429);
nand U12541 (N_12541,N_12220,N_11966);
and U12542 (N_12542,N_11898,N_12364);
nand U12543 (N_12543,N_12447,N_11969);
and U12544 (N_12544,N_11948,N_12466);
xnor U12545 (N_12545,N_11995,N_12293);
and U12546 (N_12546,N_12480,N_12382);
nor U12547 (N_12547,N_12002,N_12032);
nor U12548 (N_12548,N_12371,N_12363);
and U12549 (N_12549,N_12449,N_12075);
and U12550 (N_12550,N_12463,N_12037);
or U12551 (N_12551,N_12384,N_12111);
nor U12552 (N_12552,N_12426,N_12192);
and U12553 (N_12553,N_12163,N_12438);
and U12554 (N_12554,N_12217,N_11928);
nor U12555 (N_12555,N_11946,N_12119);
and U12556 (N_12556,N_12019,N_11984);
or U12557 (N_12557,N_12450,N_11920);
nor U12558 (N_12558,N_12477,N_12038);
nor U12559 (N_12559,N_11981,N_12099);
nor U12560 (N_12560,N_12150,N_11907);
xnor U12561 (N_12561,N_12370,N_11903);
nor U12562 (N_12562,N_12241,N_12036);
or U12563 (N_12563,N_12437,N_12277);
xnor U12564 (N_12564,N_11932,N_12243);
and U12565 (N_12565,N_12396,N_11983);
nand U12566 (N_12566,N_12042,N_12022);
and U12567 (N_12567,N_12242,N_11919);
nand U12568 (N_12568,N_12445,N_12026);
nor U12569 (N_12569,N_12428,N_12345);
xor U12570 (N_12570,N_12291,N_12071);
xnor U12571 (N_12571,N_12209,N_12154);
and U12572 (N_12572,N_12425,N_12128);
nand U12573 (N_12573,N_12431,N_12358);
or U12574 (N_12574,N_12380,N_12224);
and U12575 (N_12575,N_12459,N_12029);
nor U12576 (N_12576,N_12404,N_12271);
xnor U12577 (N_12577,N_12470,N_11927);
xnor U12578 (N_12578,N_11893,N_12118);
nor U12579 (N_12579,N_11979,N_12386);
and U12580 (N_12580,N_12196,N_12443);
xor U12581 (N_12581,N_12478,N_11937);
or U12582 (N_12582,N_12261,N_12283);
or U12583 (N_12583,N_11891,N_12072);
and U12584 (N_12584,N_12157,N_12145);
or U12585 (N_12585,N_12451,N_12397);
nand U12586 (N_12586,N_12043,N_11902);
or U12587 (N_12587,N_12127,N_12452);
and U12588 (N_12588,N_12434,N_12238);
nor U12589 (N_12589,N_11994,N_12260);
or U12590 (N_12590,N_12352,N_12148);
and U12591 (N_12591,N_11982,N_12263);
xor U12592 (N_12592,N_12302,N_12159);
and U12593 (N_12593,N_12347,N_12253);
or U12594 (N_12594,N_12498,N_12094);
nor U12595 (N_12595,N_12068,N_12289);
and U12596 (N_12596,N_12257,N_12274);
nand U12597 (N_12597,N_12472,N_12259);
or U12598 (N_12598,N_12389,N_12122);
and U12599 (N_12599,N_12120,N_11987);
and U12600 (N_12600,N_12448,N_11941);
nor U12601 (N_12601,N_12142,N_11997);
or U12602 (N_12602,N_12296,N_12195);
or U12603 (N_12603,N_12235,N_11960);
nor U12604 (N_12604,N_12360,N_12412);
and U12605 (N_12605,N_12184,N_12186);
nand U12606 (N_12606,N_12061,N_12285);
nor U12607 (N_12607,N_12092,N_12292);
nor U12608 (N_12608,N_12349,N_12351);
and U12609 (N_12609,N_12236,N_12149);
xor U12610 (N_12610,N_12460,N_11978);
xor U12611 (N_12611,N_12492,N_11889);
nor U12612 (N_12612,N_12177,N_12493);
nand U12613 (N_12613,N_12422,N_11878);
and U12614 (N_12614,N_12003,N_11973);
or U12615 (N_12615,N_12095,N_12183);
or U12616 (N_12616,N_12053,N_11882);
or U12617 (N_12617,N_12344,N_12106);
nor U12618 (N_12618,N_12170,N_12044);
nor U12619 (N_12619,N_12058,N_12465);
nor U12620 (N_12620,N_12294,N_12249);
and U12621 (N_12621,N_12074,N_12322);
and U12622 (N_12622,N_12488,N_11986);
nand U12623 (N_12623,N_12191,N_11958);
or U12624 (N_12624,N_12103,N_12273);
or U12625 (N_12625,N_12005,N_12180);
xnor U12626 (N_12626,N_12189,N_12164);
nand U12627 (N_12627,N_12487,N_12232);
and U12628 (N_12628,N_12419,N_11961);
or U12629 (N_12629,N_12230,N_12138);
nand U12630 (N_12630,N_11959,N_12388);
nand U12631 (N_12631,N_12317,N_12410);
nand U12632 (N_12632,N_12318,N_11947);
xor U12633 (N_12633,N_12346,N_12054);
nand U12634 (N_12634,N_12301,N_12458);
or U12635 (N_12635,N_12030,N_12226);
or U12636 (N_12636,N_12231,N_11918);
nor U12637 (N_12637,N_12288,N_11892);
or U12638 (N_12638,N_12399,N_12430);
nand U12639 (N_12639,N_12333,N_12050);
nor U12640 (N_12640,N_12039,N_11881);
xnor U12641 (N_12641,N_12237,N_12303);
nand U12642 (N_12642,N_12161,N_12014);
xor U12643 (N_12643,N_12015,N_12116);
nand U12644 (N_12644,N_11967,N_12338);
nor U12645 (N_12645,N_12272,N_12255);
and U12646 (N_12646,N_12060,N_12181);
or U12647 (N_12647,N_12420,N_12456);
xnor U12648 (N_12648,N_12250,N_12179);
or U12649 (N_12649,N_12270,N_12495);
or U12650 (N_12650,N_12350,N_12335);
or U12651 (N_12651,N_12066,N_12403);
or U12652 (N_12652,N_12299,N_11905);
nand U12653 (N_12653,N_12078,N_12165);
nor U12654 (N_12654,N_12041,N_11890);
or U12655 (N_12655,N_12134,N_11963);
or U12656 (N_12656,N_12334,N_12424);
xor U12657 (N_12657,N_12247,N_12093);
and U12658 (N_12658,N_12435,N_12319);
nor U12659 (N_12659,N_12009,N_12212);
nand U12660 (N_12660,N_12409,N_12136);
nor U12661 (N_12661,N_12300,N_12211);
xnor U12662 (N_12662,N_12240,N_12090);
nand U12663 (N_12663,N_11894,N_11936);
or U12664 (N_12664,N_12188,N_12469);
nor U12665 (N_12665,N_12342,N_12377);
or U12666 (N_12666,N_12016,N_12221);
nor U12667 (N_12667,N_12046,N_12077);
or U12668 (N_12668,N_11896,N_11968);
or U12669 (N_12669,N_11965,N_12442);
nor U12670 (N_12670,N_12141,N_12340);
xnor U12671 (N_12671,N_12112,N_12049);
and U12672 (N_12672,N_12218,N_12167);
nor U12673 (N_12673,N_12311,N_11906);
or U12674 (N_12674,N_11970,N_11993);
nor U12675 (N_12675,N_12281,N_12121);
nand U12676 (N_12676,N_11975,N_11964);
xor U12677 (N_12677,N_12055,N_12475);
or U12678 (N_12678,N_12067,N_12102);
xnor U12679 (N_12679,N_11998,N_12407);
and U12680 (N_12680,N_11972,N_12295);
or U12681 (N_12681,N_12310,N_12088);
nand U12682 (N_12682,N_12073,N_12267);
nor U12683 (N_12683,N_12208,N_11925);
and U12684 (N_12684,N_12028,N_12098);
or U12685 (N_12685,N_11900,N_12405);
nand U12686 (N_12686,N_12199,N_12353);
and U12687 (N_12687,N_12109,N_12304);
nor U12688 (N_12688,N_12104,N_12387);
or U12689 (N_12689,N_12406,N_11923);
or U12690 (N_12690,N_11933,N_12401);
or U12691 (N_12691,N_12354,N_12174);
or U12692 (N_12692,N_12372,N_12324);
nand U12693 (N_12693,N_12416,N_12328);
or U12694 (N_12694,N_12146,N_12057);
nand U12695 (N_12695,N_12040,N_12139);
nand U12696 (N_12696,N_12379,N_12124);
nor U12697 (N_12697,N_12368,N_12162);
nand U12698 (N_12698,N_12100,N_11883);
and U12699 (N_12699,N_12034,N_12479);
nor U12700 (N_12700,N_12251,N_12065);
and U12701 (N_12701,N_12244,N_11886);
and U12702 (N_12702,N_11991,N_12254);
or U12703 (N_12703,N_12474,N_12381);
nor U12704 (N_12704,N_12441,N_12290);
xnor U12705 (N_12705,N_12248,N_11913);
nor U12706 (N_12706,N_12144,N_12330);
or U12707 (N_12707,N_12010,N_12175);
xnor U12708 (N_12708,N_12275,N_12359);
nand U12709 (N_12709,N_12239,N_12160);
nor U12710 (N_12710,N_12313,N_12158);
nor U12711 (N_12711,N_11916,N_11904);
nand U12712 (N_12712,N_11944,N_12486);
nor U12713 (N_12713,N_12297,N_11876);
nand U12714 (N_12714,N_12227,N_11952);
nor U12715 (N_12715,N_12433,N_12233);
nand U12716 (N_12716,N_11917,N_12135);
xnor U12717 (N_12717,N_12193,N_12374);
or U12718 (N_12718,N_12216,N_12378);
or U12719 (N_12719,N_12446,N_12202);
nor U12720 (N_12720,N_12062,N_12200);
and U12721 (N_12721,N_12173,N_12182);
nand U12722 (N_12722,N_12045,N_11976);
nand U12723 (N_12723,N_12414,N_12468);
or U12724 (N_12724,N_12341,N_12356);
and U12725 (N_12725,N_12331,N_11996);
nor U12726 (N_12726,N_11880,N_12091);
xnor U12727 (N_12727,N_12276,N_12056);
and U12728 (N_12728,N_12337,N_12455);
nor U12729 (N_12729,N_11985,N_11974);
or U12730 (N_12730,N_12418,N_12210);
or U12731 (N_12731,N_12011,N_11921);
nand U12732 (N_12732,N_11940,N_11971);
or U12733 (N_12733,N_12070,N_12064);
nor U12734 (N_12734,N_12421,N_12018);
xnor U12735 (N_12735,N_12369,N_12153);
or U12736 (N_12736,N_12207,N_11942);
or U12737 (N_12737,N_12314,N_12383);
xnor U12738 (N_12738,N_12096,N_11949);
nand U12739 (N_12739,N_12415,N_12097);
nor U12740 (N_12740,N_11879,N_12484);
nor U12741 (N_12741,N_12223,N_12080);
nor U12742 (N_12742,N_12048,N_11953);
xor U12743 (N_12743,N_12023,N_11922);
nand U12744 (N_12744,N_12499,N_12258);
and U12745 (N_12745,N_12440,N_12190);
nand U12746 (N_12746,N_12084,N_12229);
and U12747 (N_12747,N_12013,N_12268);
or U12748 (N_12748,N_12081,N_11980);
nand U12749 (N_12749,N_11935,N_12033);
nand U12750 (N_12750,N_12234,N_12375);
or U12751 (N_12751,N_12176,N_11926);
and U12752 (N_12752,N_12131,N_12085);
or U12753 (N_12753,N_12215,N_12320);
xnor U12754 (N_12754,N_11951,N_12047);
nand U12755 (N_12755,N_12308,N_11977);
nand U12756 (N_12756,N_11934,N_12206);
nor U12757 (N_12757,N_12483,N_12214);
or U12758 (N_12758,N_11911,N_12476);
or U12759 (N_12759,N_12279,N_11914);
nor U12760 (N_12760,N_12126,N_11945);
and U12761 (N_12761,N_12366,N_12203);
xnor U12762 (N_12762,N_12108,N_12496);
nand U12763 (N_12763,N_12491,N_12385);
nand U12764 (N_12764,N_12101,N_12187);
nor U12765 (N_12765,N_12256,N_12219);
nor U12766 (N_12766,N_12252,N_12245);
and U12767 (N_12767,N_12348,N_12083);
nand U12768 (N_12768,N_12266,N_11954);
nand U12769 (N_12769,N_12172,N_12265);
or U12770 (N_12770,N_11957,N_12436);
and U12771 (N_12771,N_12059,N_12411);
and U12772 (N_12772,N_12309,N_12204);
xor U12773 (N_12773,N_11956,N_11915);
xor U12774 (N_12774,N_12473,N_12316);
and U12775 (N_12775,N_12198,N_12321);
nand U12776 (N_12776,N_12432,N_11877);
nor U12777 (N_12777,N_12489,N_12017);
or U12778 (N_12778,N_12213,N_12471);
nand U12779 (N_12779,N_12205,N_12152);
xor U12780 (N_12780,N_12185,N_11938);
and U12781 (N_12781,N_12395,N_12461);
xor U12782 (N_12782,N_12286,N_12035);
and U12783 (N_12783,N_12089,N_11931);
and U12784 (N_12784,N_12155,N_12417);
xor U12785 (N_12785,N_11955,N_12398);
xor U12786 (N_12786,N_12156,N_12110);
nand U12787 (N_12787,N_11962,N_12132);
or U12788 (N_12788,N_12326,N_12105);
or U12789 (N_12789,N_11908,N_11897);
nand U12790 (N_12790,N_12024,N_12021);
nor U12791 (N_12791,N_12087,N_11999);
xor U12792 (N_12792,N_12315,N_11988);
or U12793 (N_12793,N_12485,N_12362);
xnor U12794 (N_12794,N_12325,N_11912);
and U12795 (N_12795,N_12361,N_12194);
xor U12796 (N_12796,N_12086,N_11884);
or U12797 (N_12797,N_12166,N_12365);
or U12798 (N_12798,N_12113,N_12367);
and U12799 (N_12799,N_12027,N_12312);
and U12800 (N_12800,N_12201,N_12051);
and U12801 (N_12801,N_12343,N_11992);
nor U12802 (N_12802,N_12125,N_12392);
xor U12803 (N_12803,N_12490,N_12332);
xnor U12804 (N_12804,N_12228,N_12357);
or U12805 (N_12805,N_12269,N_12143);
and U12806 (N_12806,N_12123,N_12408);
xor U12807 (N_12807,N_11895,N_12454);
and U12808 (N_12808,N_12400,N_11910);
or U12809 (N_12809,N_12001,N_12284);
and U12810 (N_12810,N_11924,N_12151);
and U12811 (N_12811,N_12020,N_12393);
nor U12812 (N_12812,N_12069,N_12272);
or U12813 (N_12813,N_12478,N_12457);
nor U12814 (N_12814,N_12240,N_12246);
nand U12815 (N_12815,N_12020,N_12185);
nand U12816 (N_12816,N_11977,N_12475);
xnor U12817 (N_12817,N_12098,N_11908);
or U12818 (N_12818,N_12368,N_12115);
nor U12819 (N_12819,N_12024,N_12003);
nor U12820 (N_12820,N_12142,N_11922);
nand U12821 (N_12821,N_12251,N_12335);
nor U12822 (N_12822,N_12065,N_12498);
or U12823 (N_12823,N_12485,N_12081);
and U12824 (N_12824,N_12132,N_12424);
nand U12825 (N_12825,N_11958,N_11886);
nand U12826 (N_12826,N_12004,N_12415);
and U12827 (N_12827,N_12375,N_12391);
or U12828 (N_12828,N_12238,N_12393);
nand U12829 (N_12829,N_12230,N_12196);
or U12830 (N_12830,N_12084,N_11976);
and U12831 (N_12831,N_11877,N_12248);
xor U12832 (N_12832,N_12349,N_12227);
nor U12833 (N_12833,N_12239,N_12168);
nand U12834 (N_12834,N_11888,N_12117);
nor U12835 (N_12835,N_12124,N_12107);
xor U12836 (N_12836,N_12002,N_12400);
or U12837 (N_12837,N_12350,N_12366);
nor U12838 (N_12838,N_12464,N_12129);
nor U12839 (N_12839,N_12338,N_12081);
nand U12840 (N_12840,N_12293,N_12015);
and U12841 (N_12841,N_12119,N_12011);
or U12842 (N_12842,N_12437,N_12262);
nand U12843 (N_12843,N_12219,N_11940);
nor U12844 (N_12844,N_12471,N_12046);
xnor U12845 (N_12845,N_12219,N_12100);
nand U12846 (N_12846,N_12109,N_12326);
or U12847 (N_12847,N_11950,N_11978);
or U12848 (N_12848,N_11939,N_12032);
and U12849 (N_12849,N_12126,N_11898);
nand U12850 (N_12850,N_12161,N_11984);
nand U12851 (N_12851,N_12019,N_12020);
nand U12852 (N_12852,N_12095,N_11957);
or U12853 (N_12853,N_12475,N_11979);
nand U12854 (N_12854,N_11880,N_12328);
nor U12855 (N_12855,N_12177,N_12497);
nor U12856 (N_12856,N_12263,N_11895);
nor U12857 (N_12857,N_11975,N_12047);
xnor U12858 (N_12858,N_11963,N_12496);
or U12859 (N_12859,N_12353,N_11924);
xnor U12860 (N_12860,N_12498,N_12217);
nor U12861 (N_12861,N_11905,N_12080);
xnor U12862 (N_12862,N_12433,N_12474);
nor U12863 (N_12863,N_12301,N_12160);
and U12864 (N_12864,N_11990,N_12288);
nand U12865 (N_12865,N_12182,N_12096);
nand U12866 (N_12866,N_11907,N_12041);
xnor U12867 (N_12867,N_12301,N_11889);
nor U12868 (N_12868,N_12008,N_12457);
or U12869 (N_12869,N_11905,N_11962);
xnor U12870 (N_12870,N_12123,N_11927);
nand U12871 (N_12871,N_12009,N_12366);
xnor U12872 (N_12872,N_12465,N_12133);
nand U12873 (N_12873,N_12264,N_12424);
xor U12874 (N_12874,N_12356,N_12374);
nor U12875 (N_12875,N_11937,N_12340);
nand U12876 (N_12876,N_12274,N_12481);
nor U12877 (N_12877,N_12014,N_11894);
nor U12878 (N_12878,N_12028,N_12063);
and U12879 (N_12879,N_12386,N_12040);
xor U12880 (N_12880,N_12387,N_11895);
nor U12881 (N_12881,N_12358,N_11931);
nor U12882 (N_12882,N_12344,N_12351);
nand U12883 (N_12883,N_12310,N_12004);
xnor U12884 (N_12884,N_12348,N_12289);
and U12885 (N_12885,N_12298,N_12110);
or U12886 (N_12886,N_12252,N_12036);
nand U12887 (N_12887,N_11986,N_12273);
and U12888 (N_12888,N_12282,N_12248);
xor U12889 (N_12889,N_11977,N_12194);
nand U12890 (N_12890,N_11988,N_12032);
nor U12891 (N_12891,N_12142,N_12187);
or U12892 (N_12892,N_11933,N_11986);
and U12893 (N_12893,N_12132,N_12077);
nand U12894 (N_12894,N_12232,N_12320);
nand U12895 (N_12895,N_12337,N_12433);
nand U12896 (N_12896,N_11927,N_12360);
and U12897 (N_12897,N_12139,N_12430);
or U12898 (N_12898,N_12129,N_12401);
nand U12899 (N_12899,N_12254,N_12013);
xnor U12900 (N_12900,N_12317,N_11933);
nand U12901 (N_12901,N_11979,N_12025);
or U12902 (N_12902,N_12454,N_12326);
xor U12903 (N_12903,N_12445,N_12046);
and U12904 (N_12904,N_11948,N_12448);
nor U12905 (N_12905,N_11943,N_12082);
xor U12906 (N_12906,N_11972,N_12329);
nor U12907 (N_12907,N_11890,N_12269);
nand U12908 (N_12908,N_11940,N_12230);
or U12909 (N_12909,N_12018,N_12013);
nand U12910 (N_12910,N_12285,N_11893);
xnor U12911 (N_12911,N_12489,N_12048);
or U12912 (N_12912,N_12099,N_12111);
or U12913 (N_12913,N_11950,N_12054);
or U12914 (N_12914,N_12114,N_12258);
nor U12915 (N_12915,N_12150,N_12089);
nor U12916 (N_12916,N_12095,N_12151);
nand U12917 (N_12917,N_12127,N_11926);
nor U12918 (N_12918,N_11973,N_11950);
nand U12919 (N_12919,N_12030,N_12006);
nand U12920 (N_12920,N_12076,N_12327);
nand U12921 (N_12921,N_12442,N_12428);
xor U12922 (N_12922,N_11916,N_12386);
nor U12923 (N_12923,N_12392,N_12312);
or U12924 (N_12924,N_12453,N_12310);
nor U12925 (N_12925,N_12256,N_11940);
nand U12926 (N_12926,N_12196,N_12176);
and U12927 (N_12927,N_12388,N_12197);
and U12928 (N_12928,N_12208,N_12240);
and U12929 (N_12929,N_11946,N_12109);
nor U12930 (N_12930,N_11949,N_12136);
or U12931 (N_12931,N_12343,N_12178);
and U12932 (N_12932,N_11938,N_12130);
and U12933 (N_12933,N_12340,N_12092);
nand U12934 (N_12934,N_11939,N_12214);
nor U12935 (N_12935,N_11881,N_12366);
nor U12936 (N_12936,N_11968,N_12423);
nand U12937 (N_12937,N_11999,N_12066);
xor U12938 (N_12938,N_12264,N_12221);
or U12939 (N_12939,N_12390,N_12398);
nand U12940 (N_12940,N_11977,N_11934);
xnor U12941 (N_12941,N_11967,N_12461);
xnor U12942 (N_12942,N_12192,N_11987);
xnor U12943 (N_12943,N_12033,N_12009);
and U12944 (N_12944,N_12450,N_12411);
nand U12945 (N_12945,N_12177,N_12459);
nand U12946 (N_12946,N_12283,N_11881);
or U12947 (N_12947,N_12206,N_12188);
nor U12948 (N_12948,N_12375,N_12085);
xnor U12949 (N_12949,N_12090,N_11945);
and U12950 (N_12950,N_12288,N_12244);
nand U12951 (N_12951,N_12060,N_12414);
and U12952 (N_12952,N_12071,N_12407);
and U12953 (N_12953,N_12151,N_12275);
nand U12954 (N_12954,N_12140,N_12100);
and U12955 (N_12955,N_12270,N_12491);
nor U12956 (N_12956,N_12254,N_12253);
nand U12957 (N_12957,N_12362,N_12220);
xnor U12958 (N_12958,N_12196,N_12400);
nand U12959 (N_12959,N_11938,N_12072);
xnor U12960 (N_12960,N_11992,N_12359);
xor U12961 (N_12961,N_12271,N_12351);
nor U12962 (N_12962,N_11877,N_12363);
nand U12963 (N_12963,N_11972,N_12436);
or U12964 (N_12964,N_12135,N_12380);
nand U12965 (N_12965,N_12003,N_12461);
nand U12966 (N_12966,N_12202,N_11898);
nor U12967 (N_12967,N_12010,N_12343);
nand U12968 (N_12968,N_12319,N_11899);
xor U12969 (N_12969,N_12211,N_12026);
xor U12970 (N_12970,N_12159,N_12349);
nand U12971 (N_12971,N_12021,N_12444);
xor U12972 (N_12972,N_12000,N_12390);
and U12973 (N_12973,N_11944,N_12470);
nor U12974 (N_12974,N_12122,N_12480);
xor U12975 (N_12975,N_12475,N_12213);
and U12976 (N_12976,N_12284,N_12227);
or U12977 (N_12977,N_12296,N_11954);
xor U12978 (N_12978,N_12089,N_11915);
or U12979 (N_12979,N_12117,N_12435);
or U12980 (N_12980,N_12076,N_12248);
xnor U12981 (N_12981,N_12213,N_11879);
nand U12982 (N_12982,N_12259,N_12299);
nor U12983 (N_12983,N_12499,N_12213);
or U12984 (N_12984,N_12221,N_12150);
or U12985 (N_12985,N_12206,N_12418);
xnor U12986 (N_12986,N_12038,N_12353);
nor U12987 (N_12987,N_12096,N_12168);
nor U12988 (N_12988,N_12195,N_12221);
nor U12989 (N_12989,N_11988,N_12343);
nor U12990 (N_12990,N_12052,N_12463);
nand U12991 (N_12991,N_12305,N_11931);
nor U12992 (N_12992,N_12084,N_11881);
xnor U12993 (N_12993,N_12069,N_12478);
and U12994 (N_12994,N_12258,N_12152);
or U12995 (N_12995,N_12262,N_12470);
xnor U12996 (N_12996,N_11922,N_12385);
nor U12997 (N_12997,N_12394,N_12325);
or U12998 (N_12998,N_12475,N_11900);
xnor U12999 (N_12999,N_11987,N_12307);
xnor U13000 (N_13000,N_12465,N_12418);
and U13001 (N_13001,N_11949,N_12049);
xnor U13002 (N_13002,N_11926,N_12018);
nor U13003 (N_13003,N_12188,N_12078);
and U13004 (N_13004,N_12021,N_11885);
or U13005 (N_13005,N_11979,N_12138);
nor U13006 (N_13006,N_11964,N_12151);
or U13007 (N_13007,N_12297,N_12343);
and U13008 (N_13008,N_11898,N_11918);
nor U13009 (N_13009,N_12415,N_11896);
xnor U13010 (N_13010,N_12241,N_12430);
xor U13011 (N_13011,N_12331,N_12137);
nor U13012 (N_13012,N_12060,N_12075);
nor U13013 (N_13013,N_12034,N_11960);
or U13014 (N_13014,N_12238,N_12120);
nand U13015 (N_13015,N_12134,N_12283);
and U13016 (N_13016,N_12451,N_12456);
nor U13017 (N_13017,N_12304,N_12166);
and U13018 (N_13018,N_12365,N_12246);
xnor U13019 (N_13019,N_12215,N_12202);
xnor U13020 (N_13020,N_12431,N_12439);
or U13021 (N_13021,N_12061,N_12280);
and U13022 (N_13022,N_12464,N_12440);
nand U13023 (N_13023,N_12175,N_12102);
or U13024 (N_13024,N_12205,N_12304);
or U13025 (N_13025,N_12373,N_12309);
or U13026 (N_13026,N_11940,N_12106);
nand U13027 (N_13027,N_12297,N_11927);
or U13028 (N_13028,N_12313,N_12166);
and U13029 (N_13029,N_12462,N_12167);
and U13030 (N_13030,N_12076,N_12386);
nor U13031 (N_13031,N_12469,N_12363);
xnor U13032 (N_13032,N_12385,N_11959);
xnor U13033 (N_13033,N_12362,N_12264);
nand U13034 (N_13034,N_12000,N_12143);
xor U13035 (N_13035,N_11981,N_11941);
and U13036 (N_13036,N_12215,N_11948);
and U13037 (N_13037,N_11936,N_12475);
and U13038 (N_13038,N_11979,N_12321);
nor U13039 (N_13039,N_12278,N_12468);
nand U13040 (N_13040,N_12018,N_12486);
and U13041 (N_13041,N_12261,N_12131);
or U13042 (N_13042,N_12017,N_12108);
xor U13043 (N_13043,N_12084,N_11916);
xnor U13044 (N_13044,N_12437,N_12300);
and U13045 (N_13045,N_12076,N_12026);
or U13046 (N_13046,N_12127,N_11936);
xor U13047 (N_13047,N_12139,N_11931);
nand U13048 (N_13048,N_12347,N_12332);
and U13049 (N_13049,N_12023,N_12091);
nor U13050 (N_13050,N_12242,N_12217);
and U13051 (N_13051,N_12359,N_12433);
and U13052 (N_13052,N_12048,N_11894);
nand U13053 (N_13053,N_12064,N_12498);
or U13054 (N_13054,N_12397,N_12336);
or U13055 (N_13055,N_12264,N_12200);
nand U13056 (N_13056,N_12325,N_12382);
or U13057 (N_13057,N_12206,N_12085);
or U13058 (N_13058,N_12423,N_12321);
nor U13059 (N_13059,N_12278,N_12134);
xnor U13060 (N_13060,N_12134,N_12182);
xnor U13061 (N_13061,N_11883,N_12107);
and U13062 (N_13062,N_12073,N_12384);
nor U13063 (N_13063,N_12298,N_12340);
or U13064 (N_13064,N_12057,N_11896);
nor U13065 (N_13065,N_12409,N_12004);
xor U13066 (N_13066,N_11919,N_12435);
nand U13067 (N_13067,N_12487,N_12230);
xnor U13068 (N_13068,N_12316,N_12080);
nor U13069 (N_13069,N_12131,N_12205);
xor U13070 (N_13070,N_12277,N_12151);
nor U13071 (N_13071,N_12326,N_12055);
xnor U13072 (N_13072,N_12238,N_12441);
or U13073 (N_13073,N_12410,N_12426);
or U13074 (N_13074,N_12320,N_11943);
or U13075 (N_13075,N_12272,N_12084);
nand U13076 (N_13076,N_12468,N_11968);
nor U13077 (N_13077,N_12355,N_12338);
nand U13078 (N_13078,N_11979,N_12326);
or U13079 (N_13079,N_12444,N_12087);
or U13080 (N_13080,N_12172,N_11965);
and U13081 (N_13081,N_12337,N_12040);
or U13082 (N_13082,N_12377,N_12157);
xor U13083 (N_13083,N_12149,N_12257);
nand U13084 (N_13084,N_11897,N_12394);
or U13085 (N_13085,N_12388,N_11879);
nor U13086 (N_13086,N_11953,N_12377);
or U13087 (N_13087,N_11949,N_11952);
or U13088 (N_13088,N_12321,N_12007);
nor U13089 (N_13089,N_12143,N_11949);
nor U13090 (N_13090,N_12036,N_12258);
xnor U13091 (N_13091,N_11999,N_11996);
xor U13092 (N_13092,N_11943,N_12238);
nand U13093 (N_13093,N_12178,N_12148);
nor U13094 (N_13094,N_11905,N_12113);
and U13095 (N_13095,N_12312,N_12021);
xnor U13096 (N_13096,N_12004,N_12473);
or U13097 (N_13097,N_12335,N_12230);
nor U13098 (N_13098,N_12045,N_12027);
or U13099 (N_13099,N_12003,N_12464);
xor U13100 (N_13100,N_11898,N_12051);
and U13101 (N_13101,N_12487,N_11876);
or U13102 (N_13102,N_12027,N_12018);
xnor U13103 (N_13103,N_12112,N_12446);
xnor U13104 (N_13104,N_12459,N_12335);
nand U13105 (N_13105,N_12443,N_12327);
or U13106 (N_13106,N_12096,N_12129);
and U13107 (N_13107,N_12339,N_12310);
and U13108 (N_13108,N_12388,N_11940);
xor U13109 (N_13109,N_12440,N_11991);
or U13110 (N_13110,N_12326,N_12234);
xnor U13111 (N_13111,N_11979,N_11893);
nor U13112 (N_13112,N_12447,N_12445);
or U13113 (N_13113,N_11960,N_12045);
nor U13114 (N_13114,N_12023,N_12486);
nor U13115 (N_13115,N_12345,N_12264);
nor U13116 (N_13116,N_11986,N_12017);
nor U13117 (N_13117,N_11932,N_11962);
or U13118 (N_13118,N_12108,N_12104);
or U13119 (N_13119,N_12357,N_11988);
xor U13120 (N_13120,N_12137,N_12184);
nand U13121 (N_13121,N_12314,N_12053);
and U13122 (N_13122,N_12433,N_12271);
and U13123 (N_13123,N_12427,N_12436);
nor U13124 (N_13124,N_11886,N_12412);
or U13125 (N_13125,N_12762,N_12522);
and U13126 (N_13126,N_12667,N_12663);
or U13127 (N_13127,N_12846,N_12722);
xor U13128 (N_13128,N_12653,N_13097);
xnor U13129 (N_13129,N_12674,N_13018);
and U13130 (N_13130,N_12554,N_12580);
nand U13131 (N_13131,N_12710,N_12876);
nor U13132 (N_13132,N_13119,N_13056);
or U13133 (N_13133,N_13015,N_13031);
nand U13134 (N_13134,N_13027,N_13042);
and U13135 (N_13135,N_12840,N_12662);
or U13136 (N_13136,N_12808,N_12697);
nand U13137 (N_13137,N_12741,N_12953);
or U13138 (N_13138,N_12874,N_13024);
or U13139 (N_13139,N_13004,N_12806);
or U13140 (N_13140,N_13092,N_13009);
nand U13141 (N_13141,N_13005,N_12764);
or U13142 (N_13142,N_12931,N_12732);
xor U13143 (N_13143,N_12899,N_12779);
nor U13144 (N_13144,N_12929,N_13075);
and U13145 (N_13145,N_13113,N_12835);
or U13146 (N_13146,N_12628,N_13089);
and U13147 (N_13147,N_12773,N_12640);
xor U13148 (N_13148,N_13054,N_12730);
nand U13149 (N_13149,N_13094,N_12934);
or U13150 (N_13150,N_12873,N_13123);
xnor U13151 (N_13151,N_13017,N_12677);
or U13152 (N_13152,N_12603,N_12571);
xor U13153 (N_13153,N_12918,N_12803);
nand U13154 (N_13154,N_13048,N_12698);
nor U13155 (N_13155,N_12875,N_12908);
or U13156 (N_13156,N_13112,N_12557);
xnor U13157 (N_13157,N_12865,N_12688);
xnor U13158 (N_13158,N_12623,N_12532);
nand U13159 (N_13159,N_12750,N_12618);
or U13160 (N_13160,N_12924,N_12962);
xor U13161 (N_13161,N_12769,N_12827);
xnor U13162 (N_13162,N_12552,N_12699);
and U13163 (N_13163,N_12834,N_12787);
nand U13164 (N_13164,N_13105,N_12624);
nand U13165 (N_13165,N_12867,N_12968);
nor U13166 (N_13166,N_12757,N_12983);
xnor U13167 (N_13167,N_12989,N_12607);
and U13168 (N_13168,N_12724,N_12816);
and U13169 (N_13169,N_12965,N_12755);
nor U13170 (N_13170,N_13044,N_12966);
and U13171 (N_13171,N_13116,N_12939);
nand U13172 (N_13172,N_12706,N_12947);
nand U13173 (N_13173,N_12562,N_12907);
xnor U13174 (N_13174,N_12678,N_12501);
and U13175 (N_13175,N_12999,N_12782);
nand U13176 (N_13176,N_12725,N_12895);
and U13177 (N_13177,N_13003,N_12990);
nand U13178 (N_13178,N_12946,N_12525);
xor U13179 (N_13179,N_12716,N_12951);
or U13180 (N_13180,N_13036,N_12523);
or U13181 (N_13181,N_12855,N_12708);
or U13182 (N_13182,N_12957,N_12854);
nor U13183 (N_13183,N_12582,N_12701);
xor U13184 (N_13184,N_12746,N_12612);
xnor U13185 (N_13185,N_12889,N_12513);
nor U13186 (N_13186,N_12638,N_12879);
or U13187 (N_13187,N_12959,N_13006);
nand U13188 (N_13188,N_12928,N_12589);
nor U13189 (N_13189,N_12974,N_12933);
xnor U13190 (N_13190,N_13045,N_12936);
or U13191 (N_13191,N_13052,N_12941);
nor U13192 (N_13192,N_13110,N_12785);
nand U13193 (N_13193,N_12863,N_12614);
xnor U13194 (N_13194,N_12572,N_12801);
xor U13195 (N_13195,N_12853,N_12775);
nor U13196 (N_13196,N_12551,N_12717);
or U13197 (N_13197,N_12804,N_13096);
nor U13198 (N_13198,N_13071,N_13002);
nor U13199 (N_13199,N_12705,N_13019);
and U13200 (N_13200,N_12996,N_12858);
nor U13201 (N_13201,N_12903,N_13108);
nand U13202 (N_13202,N_12833,N_13060);
xor U13203 (N_13203,N_12646,N_12672);
and U13204 (N_13204,N_12950,N_12560);
nor U13205 (N_13205,N_12648,N_12765);
and U13206 (N_13206,N_12540,N_13023);
xnor U13207 (N_13207,N_13080,N_12654);
nand U13208 (N_13208,N_12770,N_12739);
xor U13209 (N_13209,N_12926,N_12505);
nand U13210 (N_13210,N_12753,N_12864);
or U13211 (N_13211,N_12594,N_12897);
nor U13212 (N_13212,N_12979,N_12862);
nor U13213 (N_13213,N_12527,N_12595);
xnor U13214 (N_13214,N_12937,N_12615);
and U13215 (N_13215,N_12866,N_13007);
and U13216 (N_13216,N_13064,N_12568);
and U13217 (N_13217,N_12963,N_13046);
nand U13218 (N_13218,N_12810,N_12689);
nand U13219 (N_13219,N_12998,N_12673);
and U13220 (N_13220,N_12791,N_12670);
xor U13221 (N_13221,N_12647,N_13051);
nand U13222 (N_13222,N_13049,N_12533);
nand U13223 (N_13223,N_12636,N_12524);
and U13224 (N_13224,N_13014,N_12780);
nand U13225 (N_13225,N_12760,N_12917);
xor U13226 (N_13226,N_12693,N_12904);
and U13227 (N_13227,N_13076,N_12519);
and U13228 (N_13228,N_13010,N_12945);
and U13229 (N_13229,N_12828,N_12839);
nor U13230 (N_13230,N_12799,N_12859);
nand U13231 (N_13231,N_12502,N_12868);
and U13232 (N_13232,N_12767,N_12598);
or U13233 (N_13233,N_13093,N_12536);
nor U13234 (N_13234,N_12606,N_12913);
or U13235 (N_13235,N_12986,N_12726);
nand U13236 (N_13236,N_13088,N_12585);
xor U13237 (N_13237,N_12652,N_13121);
nor U13238 (N_13238,N_12922,N_12970);
nor U13239 (N_13239,N_12604,N_12883);
nand U13240 (N_13240,N_12685,N_12844);
nor U13241 (N_13241,N_13030,N_12815);
xnor U13242 (N_13242,N_12586,N_12749);
xnor U13243 (N_13243,N_13011,N_13102);
nor U13244 (N_13244,N_12531,N_12581);
nor U13245 (N_13245,N_12916,N_12687);
and U13246 (N_13246,N_13041,N_12714);
and U13247 (N_13247,N_12972,N_12884);
nand U13248 (N_13248,N_12508,N_12512);
nand U13249 (N_13249,N_13039,N_13032);
and U13250 (N_13250,N_12901,N_12534);
xor U13251 (N_13251,N_12633,N_12555);
and U13252 (N_13252,N_12655,N_12644);
xnor U13253 (N_13253,N_12602,N_12664);
xnor U13254 (N_13254,N_12885,N_12831);
nand U13255 (N_13255,N_12632,N_13111);
xor U13256 (N_13256,N_12796,N_12600);
xnor U13257 (N_13257,N_12573,N_12691);
and U13258 (N_13258,N_12964,N_13095);
and U13259 (N_13259,N_13070,N_12790);
or U13260 (N_13260,N_12800,N_13124);
or U13261 (N_13261,N_13081,N_12814);
or U13262 (N_13262,N_12715,N_13029);
or U13263 (N_13263,N_13087,N_12747);
xnor U13264 (N_13264,N_12659,N_12973);
and U13265 (N_13265,N_12591,N_12807);
and U13266 (N_13266,N_12794,N_12975);
nand U13267 (N_13267,N_12980,N_12696);
or U13268 (N_13268,N_12639,N_13066);
xnor U13269 (N_13269,N_12704,N_12719);
nand U13270 (N_13270,N_13079,N_12821);
nor U13271 (N_13271,N_12583,N_13001);
or U13272 (N_13272,N_12967,N_13047);
nand U13273 (N_13273,N_12960,N_12621);
and U13274 (N_13274,N_12626,N_12823);
or U13275 (N_13275,N_13053,N_12813);
or U13276 (N_13276,N_13063,N_12976);
nand U13277 (N_13277,N_12669,N_12650);
or U13278 (N_13278,N_12993,N_13117);
nor U13279 (N_13279,N_13122,N_12981);
nor U13280 (N_13280,N_12611,N_12720);
and U13281 (N_13281,N_12656,N_12819);
xnor U13282 (N_13282,N_12894,N_12617);
nor U13283 (N_13283,N_12788,N_12507);
nor U13284 (N_13284,N_12778,N_12912);
nand U13285 (N_13285,N_13107,N_13084);
xnor U13286 (N_13286,N_12515,N_12563);
and U13287 (N_13287,N_13013,N_12902);
or U13288 (N_13288,N_12919,N_12718);
and U13289 (N_13289,N_12592,N_12878);
nor U13290 (N_13290,N_13000,N_12837);
xnor U13291 (N_13291,N_12535,N_12826);
xnor U13292 (N_13292,N_13103,N_12713);
xor U13293 (N_13293,N_12845,N_13055);
nor U13294 (N_13294,N_12786,N_13082);
nor U13295 (N_13295,N_13085,N_12943);
or U13296 (N_13296,N_12783,N_12811);
or U13297 (N_13297,N_12528,N_12756);
nor U13298 (N_13298,N_13074,N_12723);
xnor U13299 (N_13299,N_12545,N_12539);
nor U13300 (N_13300,N_12549,N_13034);
xnor U13301 (N_13301,N_13057,N_12818);
nand U13302 (N_13302,N_13037,N_12593);
or U13303 (N_13303,N_12938,N_12506);
nand U13304 (N_13304,N_12530,N_12578);
xor U13305 (N_13305,N_12570,N_12988);
xor U13306 (N_13306,N_12721,N_12590);
nor U13307 (N_13307,N_12977,N_12529);
nor U13308 (N_13308,N_12955,N_13065);
nor U13309 (N_13309,N_12751,N_12634);
nand U13310 (N_13310,N_12789,N_12860);
xnor U13311 (N_13311,N_12961,N_12822);
or U13312 (N_13312,N_12510,N_12548);
xor U13313 (N_13313,N_12759,N_12683);
or U13314 (N_13314,N_12731,N_12620);
xnor U13315 (N_13315,N_12679,N_12516);
nor U13316 (N_13316,N_12707,N_12547);
or U13317 (N_13317,N_12504,N_13100);
nand U13318 (N_13318,N_12849,N_12681);
xnor U13319 (N_13319,N_12686,N_13026);
nand U13320 (N_13320,N_12682,N_12841);
or U13321 (N_13321,N_12958,N_12608);
and U13322 (N_13322,N_12978,N_12896);
xnor U13323 (N_13323,N_12923,N_12891);
and U13324 (N_13324,N_12711,N_12748);
xor U13325 (N_13325,N_12930,N_12676);
nand U13326 (N_13326,N_12956,N_12511);
nand U13327 (N_13327,N_12574,N_12561);
xor U13328 (N_13328,N_12882,N_12579);
or U13329 (N_13329,N_12703,N_12601);
nand U13330 (N_13330,N_13059,N_12914);
nor U13331 (N_13331,N_12649,N_12635);
nor U13332 (N_13332,N_12763,N_13061);
nand U13333 (N_13333,N_12848,N_13058);
and U13334 (N_13334,N_12900,N_12949);
nand U13335 (N_13335,N_12577,N_12576);
nand U13336 (N_13336,N_13050,N_12692);
or U13337 (N_13337,N_12991,N_13101);
nor U13338 (N_13338,N_12761,N_12887);
and U13339 (N_13339,N_12736,N_12817);
and U13340 (N_13340,N_12569,N_12940);
xor U13341 (N_13341,N_12836,N_12641);
nor U13342 (N_13342,N_12599,N_12610);
and U13343 (N_13343,N_12935,N_13062);
nand U13344 (N_13344,N_12994,N_12738);
xor U13345 (N_13345,N_13077,N_13008);
nor U13346 (N_13346,N_12825,N_12772);
nand U13347 (N_13347,N_12743,N_12781);
xnor U13348 (N_13348,N_12971,N_12542);
nand U13349 (N_13349,N_12616,N_12872);
nor U13350 (N_13350,N_13086,N_12734);
xnor U13351 (N_13351,N_12565,N_12658);
nand U13352 (N_13352,N_12881,N_12666);
or U13353 (N_13353,N_12518,N_12869);
and U13354 (N_13354,N_12503,N_12852);
and U13355 (N_13355,N_12797,N_12997);
or U13356 (N_13356,N_12744,N_12671);
and U13357 (N_13357,N_12566,N_12812);
nor U13358 (N_13358,N_13090,N_13114);
and U13359 (N_13359,N_12847,N_12830);
xor U13360 (N_13360,N_13115,N_12543);
nor U13361 (N_13361,N_12932,N_12729);
xor U13362 (N_13362,N_12500,N_13022);
and U13363 (N_13363,N_13109,N_12870);
nand U13364 (N_13364,N_13104,N_12952);
or U13365 (N_13365,N_12890,N_12842);
nand U13366 (N_13366,N_12550,N_13120);
or U13367 (N_13367,N_12694,N_12798);
nand U13368 (N_13368,N_12857,N_12766);
and U13369 (N_13369,N_12909,N_12774);
xnor U13370 (N_13370,N_12927,N_12793);
xnor U13371 (N_13371,N_12643,N_12727);
nor U13372 (N_13372,N_12619,N_12630);
nor U13373 (N_13373,N_12809,N_12709);
xor U13374 (N_13374,N_12587,N_12892);
and U13375 (N_13375,N_12824,N_12661);
or U13376 (N_13376,N_13073,N_12995);
xnor U13377 (N_13377,N_12985,N_12982);
or U13378 (N_13378,N_12838,N_12712);
or U13379 (N_13379,N_12851,N_12668);
nand U13380 (N_13380,N_13033,N_12805);
nand U13381 (N_13381,N_12880,N_12893);
or U13382 (N_13382,N_12627,N_13012);
and U13383 (N_13383,N_13099,N_12657);
nor U13384 (N_13384,N_12784,N_12584);
xor U13385 (N_13385,N_12745,N_13025);
nor U13386 (N_13386,N_12915,N_12754);
xnor U13387 (N_13387,N_12920,N_13021);
nor U13388 (N_13388,N_12558,N_12861);
nor U13389 (N_13389,N_12768,N_12910);
xnor U13390 (N_13390,N_12625,N_13069);
or U13391 (N_13391,N_12905,N_12948);
or U13392 (N_13392,N_12752,N_12740);
nor U13393 (N_13393,N_12700,N_13098);
and U13394 (N_13394,N_12596,N_13028);
nor U13395 (N_13395,N_12898,N_12556);
nor U13396 (N_13396,N_12984,N_12820);
nor U13397 (N_13397,N_12521,N_12675);
nor U13398 (N_13398,N_12856,N_12771);
nor U13399 (N_13399,N_12925,N_12733);
or U13400 (N_13400,N_12629,N_12735);
or U13401 (N_13401,N_12597,N_12622);
and U13402 (N_13402,N_12538,N_13038);
nor U13403 (N_13403,N_12559,N_12509);
and U13404 (N_13404,N_12651,N_13035);
and U13405 (N_13405,N_12942,N_12921);
nor U13406 (N_13406,N_12728,N_12871);
or U13407 (N_13407,N_12564,N_12737);
nor U13408 (N_13408,N_13106,N_12526);
or U13409 (N_13409,N_12690,N_12886);
or U13410 (N_13410,N_12954,N_13091);
and U13411 (N_13411,N_12911,N_12613);
or U13412 (N_13412,N_13067,N_12877);
xor U13413 (N_13413,N_13043,N_12605);
nor U13414 (N_13414,N_12609,N_12777);
nor U13415 (N_13415,N_12758,N_12541);
nand U13416 (N_13416,N_12546,N_12802);
nor U13417 (N_13417,N_13016,N_12680);
nor U13418 (N_13418,N_12832,N_12742);
and U13419 (N_13419,N_12702,N_12567);
xnor U13420 (N_13420,N_12795,N_13040);
nor U13421 (N_13421,N_12776,N_12792);
nor U13422 (N_13422,N_12631,N_12660);
nor U13423 (N_13423,N_12520,N_13078);
nor U13424 (N_13424,N_13118,N_12969);
xnor U13425 (N_13425,N_12992,N_13072);
nand U13426 (N_13426,N_12537,N_12888);
and U13427 (N_13427,N_12944,N_12645);
nand U13428 (N_13428,N_12665,N_12906);
nor U13429 (N_13429,N_12843,N_12695);
and U13430 (N_13430,N_12684,N_12544);
or U13431 (N_13431,N_13068,N_12514);
or U13432 (N_13432,N_12637,N_12987);
or U13433 (N_13433,N_12642,N_12553);
xnor U13434 (N_13434,N_12850,N_12575);
or U13435 (N_13435,N_13020,N_12829);
and U13436 (N_13436,N_12517,N_12588);
nor U13437 (N_13437,N_13083,N_12679);
xor U13438 (N_13438,N_12667,N_13114);
xor U13439 (N_13439,N_12614,N_12747);
and U13440 (N_13440,N_12888,N_12649);
and U13441 (N_13441,N_12559,N_13027);
xnor U13442 (N_13442,N_12740,N_12594);
nand U13443 (N_13443,N_13110,N_12850);
or U13444 (N_13444,N_12792,N_13060);
or U13445 (N_13445,N_12858,N_13046);
nand U13446 (N_13446,N_12728,N_12749);
nand U13447 (N_13447,N_12646,N_12866);
xnor U13448 (N_13448,N_13038,N_12734);
and U13449 (N_13449,N_12521,N_12573);
nor U13450 (N_13450,N_12910,N_12540);
nor U13451 (N_13451,N_12989,N_12856);
nand U13452 (N_13452,N_13103,N_13049);
nand U13453 (N_13453,N_12542,N_12662);
and U13454 (N_13454,N_12954,N_12773);
and U13455 (N_13455,N_12694,N_13092);
nor U13456 (N_13456,N_12516,N_12783);
and U13457 (N_13457,N_13087,N_13105);
or U13458 (N_13458,N_12886,N_12884);
xnor U13459 (N_13459,N_12977,N_13112);
and U13460 (N_13460,N_12610,N_12614);
xnor U13461 (N_13461,N_12705,N_12673);
xnor U13462 (N_13462,N_12827,N_12626);
or U13463 (N_13463,N_12561,N_12714);
nand U13464 (N_13464,N_13116,N_12598);
nor U13465 (N_13465,N_13111,N_12676);
or U13466 (N_13466,N_13083,N_12789);
and U13467 (N_13467,N_13034,N_12802);
or U13468 (N_13468,N_12772,N_12777);
xnor U13469 (N_13469,N_12693,N_12559);
nand U13470 (N_13470,N_12647,N_12908);
xor U13471 (N_13471,N_12545,N_12859);
nand U13472 (N_13472,N_12989,N_12841);
nand U13473 (N_13473,N_13103,N_12748);
nor U13474 (N_13474,N_12572,N_13084);
and U13475 (N_13475,N_13028,N_12895);
or U13476 (N_13476,N_12944,N_12752);
and U13477 (N_13477,N_12616,N_12833);
and U13478 (N_13478,N_13053,N_12664);
or U13479 (N_13479,N_12627,N_12543);
xnor U13480 (N_13480,N_12971,N_12892);
nand U13481 (N_13481,N_12822,N_13033);
nor U13482 (N_13482,N_13096,N_12511);
or U13483 (N_13483,N_12519,N_12772);
and U13484 (N_13484,N_12724,N_12567);
nand U13485 (N_13485,N_12671,N_12635);
xor U13486 (N_13486,N_12905,N_13110);
nor U13487 (N_13487,N_12710,N_12859);
xnor U13488 (N_13488,N_12607,N_13025);
nand U13489 (N_13489,N_12652,N_12709);
nor U13490 (N_13490,N_12681,N_12839);
or U13491 (N_13491,N_12609,N_12547);
xnor U13492 (N_13492,N_12972,N_12970);
nor U13493 (N_13493,N_12954,N_12630);
nand U13494 (N_13494,N_12552,N_12832);
nor U13495 (N_13495,N_12671,N_12702);
xor U13496 (N_13496,N_12735,N_12560);
xnor U13497 (N_13497,N_12824,N_12980);
or U13498 (N_13498,N_12706,N_12502);
or U13499 (N_13499,N_12545,N_12936);
nand U13500 (N_13500,N_12923,N_12596);
nor U13501 (N_13501,N_13021,N_12877);
nor U13502 (N_13502,N_12597,N_12658);
nor U13503 (N_13503,N_12722,N_12763);
xnor U13504 (N_13504,N_12507,N_12560);
xor U13505 (N_13505,N_12605,N_12626);
xnor U13506 (N_13506,N_12888,N_12816);
nand U13507 (N_13507,N_12615,N_13014);
and U13508 (N_13508,N_12929,N_13041);
and U13509 (N_13509,N_12997,N_12925);
or U13510 (N_13510,N_12514,N_12931);
nor U13511 (N_13511,N_13074,N_12799);
nor U13512 (N_13512,N_12578,N_12522);
nor U13513 (N_13513,N_13007,N_12673);
nor U13514 (N_13514,N_12528,N_13088);
or U13515 (N_13515,N_12594,N_12535);
xor U13516 (N_13516,N_12822,N_12970);
or U13517 (N_13517,N_12872,N_12618);
and U13518 (N_13518,N_12548,N_12655);
nand U13519 (N_13519,N_13028,N_12567);
nand U13520 (N_13520,N_12997,N_12602);
and U13521 (N_13521,N_12677,N_12592);
xor U13522 (N_13522,N_12676,N_12802);
xor U13523 (N_13523,N_12661,N_13028);
or U13524 (N_13524,N_13080,N_12845);
nor U13525 (N_13525,N_12848,N_12535);
xnor U13526 (N_13526,N_12719,N_12679);
or U13527 (N_13527,N_13033,N_12738);
xor U13528 (N_13528,N_12773,N_12659);
nor U13529 (N_13529,N_12561,N_12810);
nand U13530 (N_13530,N_12946,N_12956);
nor U13531 (N_13531,N_13017,N_12778);
nand U13532 (N_13532,N_13106,N_12829);
nand U13533 (N_13533,N_12631,N_12953);
nor U13534 (N_13534,N_13079,N_12986);
and U13535 (N_13535,N_12935,N_12873);
xnor U13536 (N_13536,N_12574,N_12821);
xor U13537 (N_13537,N_12567,N_12837);
nand U13538 (N_13538,N_12746,N_12690);
xnor U13539 (N_13539,N_12866,N_13099);
nor U13540 (N_13540,N_12567,N_12734);
and U13541 (N_13541,N_12961,N_13046);
xor U13542 (N_13542,N_12558,N_13094);
and U13543 (N_13543,N_13084,N_12727);
and U13544 (N_13544,N_12942,N_12586);
xor U13545 (N_13545,N_12667,N_13085);
nand U13546 (N_13546,N_12768,N_13022);
nand U13547 (N_13547,N_13020,N_12945);
xnor U13548 (N_13548,N_12877,N_12615);
or U13549 (N_13549,N_12513,N_13061);
xor U13550 (N_13550,N_12565,N_12925);
or U13551 (N_13551,N_13115,N_12918);
nor U13552 (N_13552,N_12641,N_12969);
xor U13553 (N_13553,N_12777,N_12726);
or U13554 (N_13554,N_12823,N_12573);
nor U13555 (N_13555,N_12910,N_12812);
nand U13556 (N_13556,N_13121,N_12639);
xor U13557 (N_13557,N_13090,N_12661);
and U13558 (N_13558,N_12557,N_12783);
and U13559 (N_13559,N_12845,N_13064);
and U13560 (N_13560,N_12567,N_12712);
nand U13561 (N_13561,N_13044,N_12695);
or U13562 (N_13562,N_12978,N_12979);
or U13563 (N_13563,N_12708,N_13097);
nand U13564 (N_13564,N_12912,N_12827);
xnor U13565 (N_13565,N_12635,N_12977);
or U13566 (N_13566,N_12572,N_12576);
xnor U13567 (N_13567,N_12936,N_12514);
nor U13568 (N_13568,N_12773,N_12645);
nand U13569 (N_13569,N_12535,N_12661);
nand U13570 (N_13570,N_12830,N_13092);
or U13571 (N_13571,N_12720,N_12632);
and U13572 (N_13572,N_12755,N_12701);
nand U13573 (N_13573,N_13068,N_12830);
and U13574 (N_13574,N_12905,N_12911);
xor U13575 (N_13575,N_12748,N_12902);
and U13576 (N_13576,N_12750,N_12740);
or U13577 (N_13577,N_12619,N_12833);
or U13578 (N_13578,N_12541,N_12650);
or U13579 (N_13579,N_12786,N_12799);
and U13580 (N_13580,N_12713,N_12551);
nand U13581 (N_13581,N_13090,N_12758);
xor U13582 (N_13582,N_12722,N_12706);
and U13583 (N_13583,N_13093,N_12883);
xnor U13584 (N_13584,N_13070,N_12567);
or U13585 (N_13585,N_12695,N_12511);
or U13586 (N_13586,N_12815,N_12628);
and U13587 (N_13587,N_12540,N_12867);
xnor U13588 (N_13588,N_13115,N_12671);
or U13589 (N_13589,N_12925,N_12566);
and U13590 (N_13590,N_12686,N_12523);
xor U13591 (N_13591,N_12977,N_13018);
or U13592 (N_13592,N_12806,N_12915);
xnor U13593 (N_13593,N_12778,N_12503);
or U13594 (N_13594,N_12591,N_12667);
nor U13595 (N_13595,N_12871,N_13114);
nand U13596 (N_13596,N_13081,N_12951);
xor U13597 (N_13597,N_12539,N_12529);
or U13598 (N_13598,N_13115,N_12719);
xnor U13599 (N_13599,N_12604,N_13046);
xnor U13600 (N_13600,N_13034,N_12691);
nor U13601 (N_13601,N_13098,N_12900);
nand U13602 (N_13602,N_13071,N_12579);
xnor U13603 (N_13603,N_13118,N_12794);
and U13604 (N_13604,N_12650,N_12951);
nor U13605 (N_13605,N_13004,N_12926);
xor U13606 (N_13606,N_12653,N_12839);
nand U13607 (N_13607,N_12554,N_12979);
nor U13608 (N_13608,N_13006,N_12787);
and U13609 (N_13609,N_12539,N_13002);
or U13610 (N_13610,N_12963,N_12784);
nand U13611 (N_13611,N_12967,N_12552);
xor U13612 (N_13612,N_12997,N_13086);
nand U13613 (N_13613,N_12885,N_13082);
nand U13614 (N_13614,N_12717,N_13042);
and U13615 (N_13615,N_12685,N_13097);
and U13616 (N_13616,N_12644,N_12649);
nand U13617 (N_13617,N_12814,N_12632);
nor U13618 (N_13618,N_12600,N_13094);
and U13619 (N_13619,N_12736,N_12926);
nor U13620 (N_13620,N_12751,N_12780);
nor U13621 (N_13621,N_12963,N_12578);
nand U13622 (N_13622,N_12912,N_13089);
nor U13623 (N_13623,N_13044,N_12745);
nand U13624 (N_13624,N_12770,N_12508);
xor U13625 (N_13625,N_12527,N_12625);
nor U13626 (N_13626,N_13111,N_13085);
and U13627 (N_13627,N_12940,N_13078);
or U13628 (N_13628,N_13097,N_13086);
nand U13629 (N_13629,N_12819,N_12685);
or U13630 (N_13630,N_12916,N_12661);
and U13631 (N_13631,N_12973,N_13108);
or U13632 (N_13632,N_12866,N_12872);
nor U13633 (N_13633,N_12643,N_12962);
nor U13634 (N_13634,N_12790,N_12517);
and U13635 (N_13635,N_12887,N_13030);
xnor U13636 (N_13636,N_12889,N_12956);
nor U13637 (N_13637,N_12525,N_12684);
nand U13638 (N_13638,N_12939,N_12780);
or U13639 (N_13639,N_12939,N_12826);
or U13640 (N_13640,N_12926,N_12901);
nor U13641 (N_13641,N_12614,N_12833);
and U13642 (N_13642,N_13057,N_12875);
or U13643 (N_13643,N_12884,N_12575);
nand U13644 (N_13644,N_12804,N_12857);
nor U13645 (N_13645,N_12949,N_12613);
nor U13646 (N_13646,N_12791,N_12778);
or U13647 (N_13647,N_12823,N_13018);
nand U13648 (N_13648,N_13048,N_12542);
and U13649 (N_13649,N_12906,N_12556);
nand U13650 (N_13650,N_13077,N_12757);
nor U13651 (N_13651,N_12858,N_13122);
nor U13652 (N_13652,N_12922,N_13110);
and U13653 (N_13653,N_13014,N_12926);
nand U13654 (N_13654,N_12578,N_12688);
nor U13655 (N_13655,N_13019,N_12667);
nor U13656 (N_13656,N_12872,N_12503);
nor U13657 (N_13657,N_12884,N_12579);
nor U13658 (N_13658,N_13069,N_13035);
nor U13659 (N_13659,N_13038,N_13013);
nand U13660 (N_13660,N_12785,N_12833);
and U13661 (N_13661,N_12919,N_12996);
xnor U13662 (N_13662,N_12602,N_12774);
nand U13663 (N_13663,N_12541,N_12587);
or U13664 (N_13664,N_13075,N_12767);
or U13665 (N_13665,N_12703,N_12585);
or U13666 (N_13666,N_12703,N_12971);
xor U13667 (N_13667,N_12866,N_13038);
or U13668 (N_13668,N_12700,N_13064);
nand U13669 (N_13669,N_12782,N_13116);
or U13670 (N_13670,N_12587,N_12842);
and U13671 (N_13671,N_12733,N_12815);
nand U13672 (N_13672,N_12976,N_12605);
xnor U13673 (N_13673,N_13035,N_12866);
nand U13674 (N_13674,N_12614,N_12705);
or U13675 (N_13675,N_12603,N_12605);
xnor U13676 (N_13676,N_12808,N_12989);
nor U13677 (N_13677,N_12710,N_13031);
or U13678 (N_13678,N_12630,N_13114);
nand U13679 (N_13679,N_12533,N_12535);
nand U13680 (N_13680,N_13094,N_12852);
nand U13681 (N_13681,N_12992,N_12781);
nand U13682 (N_13682,N_12797,N_12738);
and U13683 (N_13683,N_12936,N_13117);
nand U13684 (N_13684,N_12664,N_12935);
and U13685 (N_13685,N_12648,N_12926);
nor U13686 (N_13686,N_12941,N_12606);
nand U13687 (N_13687,N_12962,N_12933);
and U13688 (N_13688,N_13042,N_12723);
and U13689 (N_13689,N_12962,N_12959);
or U13690 (N_13690,N_12789,N_13105);
or U13691 (N_13691,N_12656,N_12822);
nand U13692 (N_13692,N_13054,N_12812);
nand U13693 (N_13693,N_12834,N_12866);
or U13694 (N_13694,N_12623,N_13008);
nor U13695 (N_13695,N_13077,N_12671);
or U13696 (N_13696,N_12788,N_12984);
xnor U13697 (N_13697,N_13091,N_12842);
or U13698 (N_13698,N_12750,N_12543);
or U13699 (N_13699,N_12862,N_12585);
nand U13700 (N_13700,N_12788,N_12624);
nor U13701 (N_13701,N_12771,N_12686);
or U13702 (N_13702,N_13105,N_13035);
and U13703 (N_13703,N_12849,N_12835);
xnor U13704 (N_13704,N_12683,N_13013);
and U13705 (N_13705,N_13025,N_13040);
nand U13706 (N_13706,N_12865,N_12569);
nand U13707 (N_13707,N_12699,N_12918);
and U13708 (N_13708,N_12549,N_12647);
nor U13709 (N_13709,N_12771,N_12723);
and U13710 (N_13710,N_12523,N_12613);
xor U13711 (N_13711,N_12829,N_13110);
and U13712 (N_13712,N_12704,N_12824);
nor U13713 (N_13713,N_12747,N_12755);
or U13714 (N_13714,N_12933,N_12743);
xor U13715 (N_13715,N_12683,N_13034);
nor U13716 (N_13716,N_13111,N_12965);
and U13717 (N_13717,N_12801,N_12693);
nor U13718 (N_13718,N_12786,N_12716);
and U13719 (N_13719,N_12575,N_12664);
xnor U13720 (N_13720,N_12836,N_13119);
nand U13721 (N_13721,N_13041,N_13107);
xor U13722 (N_13722,N_12890,N_12970);
or U13723 (N_13723,N_12843,N_12728);
xnor U13724 (N_13724,N_12837,N_12810);
nand U13725 (N_13725,N_12838,N_12820);
nor U13726 (N_13726,N_12905,N_12954);
and U13727 (N_13727,N_12824,N_13074);
or U13728 (N_13728,N_13104,N_12691);
xor U13729 (N_13729,N_13081,N_12643);
or U13730 (N_13730,N_12554,N_12733);
nand U13731 (N_13731,N_12532,N_12747);
nor U13732 (N_13732,N_12743,N_12803);
and U13733 (N_13733,N_12876,N_13102);
or U13734 (N_13734,N_12790,N_12691);
and U13735 (N_13735,N_12594,N_12662);
nand U13736 (N_13736,N_13059,N_13006);
or U13737 (N_13737,N_12983,N_13070);
and U13738 (N_13738,N_12827,N_12562);
and U13739 (N_13739,N_12817,N_13070);
xor U13740 (N_13740,N_12631,N_13003);
nor U13741 (N_13741,N_12851,N_13091);
or U13742 (N_13742,N_12521,N_12797);
nand U13743 (N_13743,N_12540,N_12643);
xnor U13744 (N_13744,N_12741,N_13068);
nor U13745 (N_13745,N_12821,N_12951);
and U13746 (N_13746,N_12562,N_13000);
nor U13747 (N_13747,N_12912,N_12811);
xnor U13748 (N_13748,N_12859,N_12903);
nand U13749 (N_13749,N_12764,N_12663);
nor U13750 (N_13750,N_13578,N_13541);
nand U13751 (N_13751,N_13707,N_13691);
and U13752 (N_13752,N_13730,N_13344);
xnor U13753 (N_13753,N_13742,N_13150);
nand U13754 (N_13754,N_13470,N_13465);
and U13755 (N_13755,N_13573,N_13619);
or U13756 (N_13756,N_13645,N_13142);
and U13757 (N_13757,N_13587,N_13219);
nand U13758 (N_13758,N_13434,N_13630);
xnor U13759 (N_13759,N_13641,N_13747);
xnor U13760 (N_13760,N_13467,N_13301);
nand U13761 (N_13761,N_13611,N_13250);
nor U13762 (N_13762,N_13420,N_13677);
xnor U13763 (N_13763,N_13511,N_13409);
nor U13764 (N_13764,N_13422,N_13520);
nor U13765 (N_13765,N_13140,N_13428);
and U13766 (N_13766,N_13359,N_13287);
xor U13767 (N_13767,N_13671,N_13321);
nor U13768 (N_13768,N_13681,N_13697);
nand U13769 (N_13769,N_13205,N_13355);
and U13770 (N_13770,N_13666,N_13448);
or U13771 (N_13771,N_13188,N_13291);
or U13772 (N_13772,N_13688,N_13336);
and U13773 (N_13773,N_13550,N_13309);
or U13774 (N_13774,N_13591,N_13647);
nand U13775 (N_13775,N_13225,N_13655);
and U13776 (N_13776,N_13593,N_13684);
nor U13777 (N_13777,N_13464,N_13538);
nand U13778 (N_13778,N_13401,N_13583);
and U13779 (N_13779,N_13727,N_13518);
nand U13780 (N_13780,N_13378,N_13269);
or U13781 (N_13781,N_13594,N_13281);
and U13782 (N_13782,N_13226,N_13721);
xor U13783 (N_13783,N_13625,N_13559);
or U13784 (N_13784,N_13517,N_13168);
nor U13785 (N_13785,N_13664,N_13158);
and U13786 (N_13786,N_13329,N_13376);
and U13787 (N_13787,N_13694,N_13366);
and U13788 (N_13788,N_13739,N_13350);
and U13789 (N_13789,N_13406,N_13438);
and U13790 (N_13790,N_13689,N_13632);
xor U13791 (N_13791,N_13729,N_13624);
nand U13792 (N_13792,N_13457,N_13151);
and U13793 (N_13793,N_13155,N_13183);
or U13794 (N_13794,N_13682,N_13266);
nor U13795 (N_13795,N_13145,N_13424);
xor U13796 (N_13796,N_13516,N_13618);
and U13797 (N_13797,N_13127,N_13640);
nand U13798 (N_13798,N_13582,N_13282);
nor U13799 (N_13799,N_13455,N_13244);
nor U13800 (N_13800,N_13608,N_13508);
nand U13801 (N_13801,N_13303,N_13216);
and U13802 (N_13802,N_13567,N_13740);
and U13803 (N_13803,N_13139,N_13523);
nor U13804 (N_13804,N_13163,N_13288);
nor U13805 (N_13805,N_13462,N_13149);
and U13806 (N_13806,N_13256,N_13357);
nor U13807 (N_13807,N_13427,N_13196);
xor U13808 (N_13808,N_13502,N_13732);
nor U13809 (N_13809,N_13577,N_13481);
xnor U13810 (N_13810,N_13607,N_13135);
nand U13811 (N_13811,N_13296,N_13335);
xnor U13812 (N_13812,N_13695,N_13504);
nand U13813 (N_13813,N_13657,N_13658);
xor U13814 (N_13814,N_13514,N_13373);
nor U13815 (N_13815,N_13633,N_13408);
nand U13816 (N_13816,N_13495,N_13700);
nand U13817 (N_13817,N_13386,N_13141);
or U13818 (N_13818,N_13293,N_13643);
or U13819 (N_13819,N_13597,N_13346);
nor U13820 (N_13820,N_13543,N_13227);
or U13821 (N_13821,N_13662,N_13442);
xnor U13822 (N_13822,N_13327,N_13260);
and U13823 (N_13823,N_13445,N_13191);
and U13824 (N_13824,N_13319,N_13356);
xnor U13825 (N_13825,N_13562,N_13606);
or U13826 (N_13826,N_13546,N_13340);
and U13827 (N_13827,N_13530,N_13324);
nand U13828 (N_13828,N_13690,N_13341);
xnor U13829 (N_13829,N_13125,N_13713);
or U13830 (N_13830,N_13181,N_13230);
and U13831 (N_13831,N_13685,N_13544);
nor U13832 (N_13832,N_13274,N_13494);
nor U13833 (N_13833,N_13153,N_13236);
or U13834 (N_13834,N_13663,N_13547);
and U13835 (N_13835,N_13499,N_13268);
and U13836 (N_13836,N_13200,N_13195);
or U13837 (N_13837,N_13358,N_13369);
and U13838 (N_13838,N_13307,N_13722);
nand U13839 (N_13839,N_13642,N_13472);
or U13840 (N_13840,N_13429,N_13283);
xnor U13841 (N_13841,N_13551,N_13131);
or U13842 (N_13842,N_13352,N_13610);
and U13843 (N_13843,N_13147,N_13339);
or U13844 (N_13844,N_13733,N_13349);
nand U13845 (N_13845,N_13717,N_13699);
nor U13846 (N_13846,N_13235,N_13459);
xnor U13847 (N_13847,N_13133,N_13678);
and U13848 (N_13848,N_13414,N_13620);
xor U13849 (N_13849,N_13257,N_13672);
nor U13850 (N_13850,N_13483,N_13389);
nand U13851 (N_13851,N_13279,N_13634);
or U13852 (N_13852,N_13261,N_13186);
nor U13853 (N_13853,N_13411,N_13555);
and U13854 (N_13854,N_13390,N_13525);
and U13855 (N_13855,N_13704,N_13744);
or U13856 (N_13856,N_13454,N_13400);
nor U13857 (N_13857,N_13501,N_13271);
nor U13858 (N_13858,N_13322,N_13627);
xnor U13859 (N_13859,N_13253,N_13510);
nor U13860 (N_13860,N_13614,N_13354);
xor U13861 (N_13861,N_13696,N_13581);
and U13862 (N_13862,N_13654,N_13710);
xnor U13863 (N_13863,N_13534,N_13526);
nand U13864 (N_13864,N_13646,N_13152);
and U13865 (N_13865,N_13167,N_13580);
and U13866 (N_13866,N_13204,N_13201);
or U13867 (N_13867,N_13714,N_13749);
xnor U13868 (N_13868,N_13435,N_13206);
xor U13869 (N_13869,N_13370,N_13723);
xnor U13870 (N_13870,N_13492,N_13687);
nand U13871 (N_13871,N_13493,N_13715);
and U13872 (N_13872,N_13392,N_13217);
and U13873 (N_13873,N_13469,N_13143);
xnor U13874 (N_13874,N_13248,N_13439);
and U13875 (N_13875,N_13361,N_13192);
nand U13876 (N_13876,N_13505,N_13399);
and U13877 (N_13877,N_13426,N_13616);
nand U13878 (N_13878,N_13166,N_13323);
nand U13879 (N_13879,N_13460,N_13524);
nor U13880 (N_13880,N_13379,N_13299);
nor U13881 (N_13881,N_13576,N_13238);
and U13882 (N_13882,N_13294,N_13475);
nor U13883 (N_13883,N_13626,N_13265);
xnor U13884 (N_13884,N_13197,N_13148);
xnor U13885 (N_13885,N_13180,N_13635);
nand U13886 (N_13886,N_13639,N_13368);
nand U13887 (N_13887,N_13234,N_13665);
nand U13888 (N_13888,N_13300,N_13182);
or U13889 (N_13889,N_13285,N_13245);
xor U13890 (N_13890,N_13644,N_13566);
and U13891 (N_13891,N_13251,N_13387);
and U13892 (N_13892,N_13652,N_13239);
or U13893 (N_13893,N_13129,N_13609);
xnor U13894 (N_13894,N_13385,N_13276);
or U13895 (N_13895,N_13174,N_13337);
xor U13896 (N_13896,N_13584,N_13289);
or U13897 (N_13897,N_13474,N_13712);
and U13898 (N_13898,N_13491,N_13277);
and U13899 (N_13899,N_13193,N_13628);
xor U13900 (N_13900,N_13410,N_13212);
xor U13901 (N_13901,N_13210,N_13222);
and U13902 (N_13902,N_13160,N_13432);
nor U13903 (N_13903,N_13734,N_13456);
and U13904 (N_13904,N_13402,N_13692);
and U13905 (N_13905,N_13512,N_13348);
nor U13906 (N_13906,N_13716,N_13381);
nand U13907 (N_13907,N_13331,N_13605);
xor U13908 (N_13908,N_13421,N_13636);
xnor U13909 (N_13909,N_13130,N_13332);
or U13910 (N_13910,N_13450,N_13425);
or U13911 (N_13911,N_13683,N_13728);
nand U13912 (N_13912,N_13667,N_13668);
nand U13913 (N_13913,N_13416,N_13725);
or U13914 (N_13914,N_13709,N_13488);
or U13915 (N_13915,N_13650,N_13229);
or U13916 (N_13916,N_13603,N_13675);
nand U13917 (N_13917,N_13602,N_13476);
xnor U13918 (N_13918,N_13731,N_13487);
or U13919 (N_13919,N_13589,N_13187);
and U13920 (N_13920,N_13533,N_13506);
and U13921 (N_13921,N_13540,N_13417);
and U13922 (N_13922,N_13449,N_13480);
nand U13923 (N_13923,N_13539,N_13413);
or U13924 (N_13924,N_13209,N_13367);
nor U13925 (N_13925,N_13144,N_13231);
and U13926 (N_13926,N_13519,N_13444);
and U13927 (N_13927,N_13146,N_13586);
nand U13928 (N_13928,N_13221,N_13453);
and U13929 (N_13929,N_13372,N_13371);
nor U13930 (N_13930,N_13310,N_13484);
xor U13931 (N_13931,N_13254,N_13443);
nor U13932 (N_13932,N_13128,N_13263);
and U13933 (N_13933,N_13391,N_13554);
and U13934 (N_13934,N_13679,N_13446);
nor U13935 (N_13935,N_13553,N_13579);
nand U13936 (N_13936,N_13249,N_13264);
and U13937 (N_13937,N_13176,N_13314);
or U13938 (N_13938,N_13360,N_13441);
nor U13939 (N_13939,N_13165,N_13702);
xor U13940 (N_13940,N_13220,N_13275);
nor U13941 (N_13941,N_13637,N_13503);
and U13942 (N_13942,N_13617,N_13164);
nand U13943 (N_13943,N_13362,N_13126);
and U13944 (N_13944,N_13437,N_13393);
nand U13945 (N_13945,N_13574,N_13447);
and U13946 (N_13946,N_13568,N_13383);
xnor U13947 (N_13947,N_13179,N_13161);
nor U13948 (N_13948,N_13316,N_13592);
and U13949 (N_13949,N_13394,N_13490);
xor U13950 (N_13950,N_13433,N_13598);
xnor U13951 (N_13951,N_13527,N_13522);
nand U13952 (N_13952,N_13156,N_13178);
nand U13953 (N_13953,N_13171,N_13315);
or U13954 (N_13954,N_13500,N_13313);
nand U13955 (N_13955,N_13342,N_13375);
nand U13956 (N_13956,N_13532,N_13557);
nor U13957 (N_13957,N_13440,N_13351);
and U13958 (N_13958,N_13292,N_13267);
and U13959 (N_13959,N_13735,N_13243);
or U13960 (N_13960,N_13588,N_13564);
nand U13961 (N_13961,N_13384,N_13473);
and U13962 (N_13962,N_13738,N_13585);
xnor U13963 (N_13963,N_13173,N_13529);
nand U13964 (N_13964,N_13651,N_13136);
nand U13965 (N_13965,N_13157,N_13560);
xnor U13966 (N_13966,N_13353,N_13189);
xor U13967 (N_13967,N_13724,N_13590);
and U13968 (N_13968,N_13177,N_13537);
or U13969 (N_13969,N_13452,N_13380);
nor U13970 (N_13970,N_13482,N_13403);
and U13971 (N_13971,N_13304,N_13278);
or U13972 (N_13972,N_13240,N_13169);
nor U13973 (N_13973,N_13571,N_13302);
nand U13974 (N_13974,N_13412,N_13536);
or U13975 (N_13975,N_13218,N_13207);
nor U13976 (N_13976,N_13613,N_13228);
xor U13977 (N_13977,N_13280,N_13170);
nor U13978 (N_13978,N_13748,N_13320);
nor U13979 (N_13979,N_13515,N_13565);
nand U13980 (N_13980,N_13374,N_13737);
nand U13981 (N_13981,N_13436,N_13604);
or U13982 (N_13982,N_13134,N_13458);
and U13983 (N_13983,N_13570,N_13214);
or U13984 (N_13984,N_13270,N_13719);
xnor U13985 (N_13985,N_13398,N_13659);
and U13986 (N_13986,N_13252,N_13615);
xnor U13987 (N_13987,N_13138,N_13531);
and U13988 (N_13988,N_13132,N_13674);
or U13989 (N_13989,N_13325,N_13623);
and U13990 (N_13990,N_13159,N_13334);
xnor U13991 (N_13991,N_13345,N_13477);
or U13992 (N_13992,N_13317,N_13638);
and U13993 (N_13993,N_13698,N_13377);
xor U13994 (N_13994,N_13556,N_13693);
and U13995 (N_13995,N_13468,N_13365);
nor U13996 (N_13996,N_13545,N_13563);
nor U13997 (N_13997,N_13258,N_13552);
nand U13998 (N_13998,N_13478,N_13575);
xnor U13999 (N_13999,N_13711,N_13466);
and U14000 (N_14000,N_13363,N_13233);
nand U14001 (N_14001,N_13404,N_13298);
and U14002 (N_14002,N_13190,N_13242);
or U14003 (N_14003,N_13479,N_13471);
nand U14004 (N_14004,N_13743,N_13653);
nor U14005 (N_14005,N_13461,N_13528);
nor U14006 (N_14006,N_13415,N_13612);
or U14007 (N_14007,N_13199,N_13535);
nand U14008 (N_14008,N_13418,N_13202);
nand U14009 (N_14009,N_13621,N_13162);
xnor U14010 (N_14010,N_13232,N_13312);
nor U14011 (N_14011,N_13656,N_13396);
or U14012 (N_14012,N_13330,N_13509);
nor U14013 (N_14013,N_13572,N_13431);
xor U14014 (N_14014,N_13720,N_13549);
or U14015 (N_14015,N_13703,N_13419);
nor U14016 (N_14016,N_13463,N_13382);
and U14017 (N_14017,N_13542,N_13295);
nand U14018 (N_14018,N_13741,N_13137);
nand U14019 (N_14019,N_13649,N_13599);
or U14020 (N_14020,N_13255,N_13451);
nand U14021 (N_14021,N_13286,N_13213);
nor U14022 (N_14022,N_13548,N_13680);
and U14023 (N_14023,N_13631,N_13208);
nor U14024 (N_14024,N_13497,N_13676);
nor U14025 (N_14025,N_13622,N_13569);
nor U14026 (N_14026,N_13246,N_13669);
nor U14027 (N_14027,N_13405,N_13423);
or U14028 (N_14028,N_13318,N_13237);
and U14029 (N_14029,N_13648,N_13430);
and U14030 (N_14030,N_13272,N_13306);
xnor U14031 (N_14031,N_13259,N_13706);
or U14032 (N_14032,N_13290,N_13746);
nand U14033 (N_14033,N_13726,N_13326);
nand U14034 (N_14034,N_13558,N_13595);
and U14035 (N_14035,N_13485,N_13673);
nand U14036 (N_14036,N_13223,N_13705);
or U14037 (N_14037,N_13338,N_13561);
xnor U14038 (N_14038,N_13521,N_13211);
xnor U14039 (N_14039,N_13629,N_13215);
xnor U14040 (N_14040,N_13407,N_13224);
and U14041 (N_14041,N_13395,N_13343);
xor U14042 (N_14042,N_13596,N_13172);
nor U14043 (N_14043,N_13198,N_13600);
or U14044 (N_14044,N_13701,N_13308);
or U14045 (N_14045,N_13273,N_13347);
or U14046 (N_14046,N_13305,N_13486);
nand U14047 (N_14047,N_13718,N_13364);
nor U14048 (N_14048,N_13670,N_13241);
nor U14049 (N_14049,N_13247,N_13203);
or U14050 (N_14050,N_13297,N_13708);
or U14051 (N_14051,N_13185,N_13661);
and U14052 (N_14052,N_13284,N_13507);
nor U14053 (N_14053,N_13328,N_13489);
nand U14054 (N_14054,N_13745,N_13498);
xnor U14055 (N_14055,N_13184,N_13736);
and U14056 (N_14056,N_13601,N_13686);
xnor U14057 (N_14057,N_13333,N_13175);
nand U14058 (N_14058,N_13388,N_13154);
and U14059 (N_14059,N_13194,N_13262);
nand U14060 (N_14060,N_13311,N_13397);
and U14061 (N_14061,N_13660,N_13513);
or U14062 (N_14062,N_13496,N_13277);
and U14063 (N_14063,N_13568,N_13197);
and U14064 (N_14064,N_13237,N_13730);
and U14065 (N_14065,N_13180,N_13310);
xnor U14066 (N_14066,N_13162,N_13359);
or U14067 (N_14067,N_13425,N_13537);
nand U14068 (N_14068,N_13564,N_13482);
nand U14069 (N_14069,N_13335,N_13393);
or U14070 (N_14070,N_13216,N_13145);
nor U14071 (N_14071,N_13242,N_13686);
or U14072 (N_14072,N_13456,N_13186);
nor U14073 (N_14073,N_13433,N_13159);
nor U14074 (N_14074,N_13638,N_13585);
or U14075 (N_14075,N_13216,N_13727);
and U14076 (N_14076,N_13626,N_13228);
or U14077 (N_14077,N_13635,N_13624);
and U14078 (N_14078,N_13249,N_13272);
nand U14079 (N_14079,N_13274,N_13551);
xnor U14080 (N_14080,N_13183,N_13165);
nor U14081 (N_14081,N_13481,N_13216);
and U14082 (N_14082,N_13161,N_13211);
nand U14083 (N_14083,N_13382,N_13544);
and U14084 (N_14084,N_13129,N_13270);
nor U14085 (N_14085,N_13323,N_13724);
nor U14086 (N_14086,N_13528,N_13271);
nand U14087 (N_14087,N_13187,N_13169);
xnor U14088 (N_14088,N_13404,N_13274);
xor U14089 (N_14089,N_13632,N_13143);
nand U14090 (N_14090,N_13584,N_13532);
and U14091 (N_14091,N_13550,N_13402);
and U14092 (N_14092,N_13511,N_13550);
or U14093 (N_14093,N_13338,N_13381);
nand U14094 (N_14094,N_13395,N_13699);
and U14095 (N_14095,N_13216,N_13365);
or U14096 (N_14096,N_13697,N_13492);
nor U14097 (N_14097,N_13740,N_13636);
xor U14098 (N_14098,N_13609,N_13547);
nor U14099 (N_14099,N_13456,N_13491);
nor U14100 (N_14100,N_13407,N_13208);
xnor U14101 (N_14101,N_13621,N_13227);
nand U14102 (N_14102,N_13284,N_13508);
xor U14103 (N_14103,N_13544,N_13569);
xor U14104 (N_14104,N_13732,N_13593);
or U14105 (N_14105,N_13737,N_13408);
and U14106 (N_14106,N_13191,N_13172);
or U14107 (N_14107,N_13523,N_13279);
or U14108 (N_14108,N_13570,N_13333);
or U14109 (N_14109,N_13183,N_13270);
or U14110 (N_14110,N_13537,N_13143);
nor U14111 (N_14111,N_13340,N_13581);
nor U14112 (N_14112,N_13496,N_13297);
xor U14113 (N_14113,N_13175,N_13633);
and U14114 (N_14114,N_13305,N_13610);
nor U14115 (N_14115,N_13384,N_13511);
and U14116 (N_14116,N_13350,N_13464);
nand U14117 (N_14117,N_13347,N_13736);
or U14118 (N_14118,N_13575,N_13360);
and U14119 (N_14119,N_13434,N_13210);
nor U14120 (N_14120,N_13547,N_13440);
nand U14121 (N_14121,N_13426,N_13371);
xnor U14122 (N_14122,N_13237,N_13210);
nand U14123 (N_14123,N_13275,N_13526);
nand U14124 (N_14124,N_13626,N_13293);
nand U14125 (N_14125,N_13151,N_13526);
nor U14126 (N_14126,N_13685,N_13629);
and U14127 (N_14127,N_13684,N_13205);
nand U14128 (N_14128,N_13350,N_13456);
nand U14129 (N_14129,N_13618,N_13388);
nand U14130 (N_14130,N_13252,N_13688);
nand U14131 (N_14131,N_13483,N_13455);
nand U14132 (N_14132,N_13619,N_13330);
nor U14133 (N_14133,N_13682,N_13132);
or U14134 (N_14134,N_13735,N_13508);
nand U14135 (N_14135,N_13534,N_13609);
nand U14136 (N_14136,N_13614,N_13494);
and U14137 (N_14137,N_13657,N_13262);
nand U14138 (N_14138,N_13698,N_13746);
or U14139 (N_14139,N_13320,N_13627);
or U14140 (N_14140,N_13715,N_13288);
xnor U14141 (N_14141,N_13689,N_13380);
nor U14142 (N_14142,N_13255,N_13746);
nor U14143 (N_14143,N_13157,N_13462);
nand U14144 (N_14144,N_13549,N_13442);
and U14145 (N_14145,N_13462,N_13663);
xnor U14146 (N_14146,N_13262,N_13193);
and U14147 (N_14147,N_13224,N_13141);
xnor U14148 (N_14148,N_13520,N_13385);
nor U14149 (N_14149,N_13515,N_13170);
or U14150 (N_14150,N_13130,N_13287);
nand U14151 (N_14151,N_13503,N_13606);
and U14152 (N_14152,N_13364,N_13433);
nor U14153 (N_14153,N_13356,N_13327);
xor U14154 (N_14154,N_13749,N_13516);
nand U14155 (N_14155,N_13399,N_13428);
nor U14156 (N_14156,N_13206,N_13728);
or U14157 (N_14157,N_13392,N_13176);
xnor U14158 (N_14158,N_13185,N_13597);
and U14159 (N_14159,N_13343,N_13602);
or U14160 (N_14160,N_13329,N_13635);
nor U14161 (N_14161,N_13738,N_13587);
or U14162 (N_14162,N_13418,N_13621);
and U14163 (N_14163,N_13349,N_13419);
xor U14164 (N_14164,N_13159,N_13477);
or U14165 (N_14165,N_13212,N_13612);
nor U14166 (N_14166,N_13385,N_13212);
nand U14167 (N_14167,N_13473,N_13309);
nand U14168 (N_14168,N_13723,N_13687);
or U14169 (N_14169,N_13662,N_13466);
nor U14170 (N_14170,N_13282,N_13443);
nor U14171 (N_14171,N_13702,N_13568);
xor U14172 (N_14172,N_13172,N_13298);
xnor U14173 (N_14173,N_13419,N_13425);
nand U14174 (N_14174,N_13538,N_13690);
nor U14175 (N_14175,N_13200,N_13546);
nand U14176 (N_14176,N_13625,N_13512);
and U14177 (N_14177,N_13236,N_13417);
nor U14178 (N_14178,N_13512,N_13194);
nor U14179 (N_14179,N_13714,N_13443);
or U14180 (N_14180,N_13148,N_13240);
or U14181 (N_14181,N_13135,N_13236);
nand U14182 (N_14182,N_13568,N_13570);
xor U14183 (N_14183,N_13615,N_13642);
xnor U14184 (N_14184,N_13423,N_13635);
xnor U14185 (N_14185,N_13554,N_13563);
and U14186 (N_14186,N_13433,N_13595);
nor U14187 (N_14187,N_13642,N_13396);
xor U14188 (N_14188,N_13385,N_13300);
nand U14189 (N_14189,N_13414,N_13656);
nor U14190 (N_14190,N_13408,N_13256);
nand U14191 (N_14191,N_13150,N_13554);
nand U14192 (N_14192,N_13257,N_13677);
xnor U14193 (N_14193,N_13291,N_13387);
xnor U14194 (N_14194,N_13298,N_13675);
and U14195 (N_14195,N_13170,N_13208);
nor U14196 (N_14196,N_13264,N_13405);
nand U14197 (N_14197,N_13328,N_13498);
xor U14198 (N_14198,N_13322,N_13626);
nor U14199 (N_14199,N_13734,N_13436);
or U14200 (N_14200,N_13137,N_13191);
and U14201 (N_14201,N_13530,N_13427);
or U14202 (N_14202,N_13130,N_13664);
or U14203 (N_14203,N_13234,N_13353);
nor U14204 (N_14204,N_13212,N_13603);
nor U14205 (N_14205,N_13544,N_13662);
and U14206 (N_14206,N_13208,N_13577);
and U14207 (N_14207,N_13691,N_13511);
nand U14208 (N_14208,N_13538,N_13262);
xnor U14209 (N_14209,N_13155,N_13171);
xor U14210 (N_14210,N_13659,N_13221);
nand U14211 (N_14211,N_13235,N_13560);
nor U14212 (N_14212,N_13151,N_13493);
or U14213 (N_14213,N_13180,N_13146);
nand U14214 (N_14214,N_13427,N_13484);
or U14215 (N_14215,N_13510,N_13337);
xor U14216 (N_14216,N_13513,N_13407);
xnor U14217 (N_14217,N_13203,N_13271);
or U14218 (N_14218,N_13392,N_13198);
and U14219 (N_14219,N_13654,N_13351);
and U14220 (N_14220,N_13702,N_13237);
nand U14221 (N_14221,N_13740,N_13538);
and U14222 (N_14222,N_13317,N_13332);
or U14223 (N_14223,N_13627,N_13716);
nor U14224 (N_14224,N_13633,N_13209);
nand U14225 (N_14225,N_13663,N_13496);
xor U14226 (N_14226,N_13679,N_13149);
xor U14227 (N_14227,N_13245,N_13581);
nor U14228 (N_14228,N_13331,N_13200);
xor U14229 (N_14229,N_13290,N_13557);
and U14230 (N_14230,N_13435,N_13313);
or U14231 (N_14231,N_13443,N_13285);
nand U14232 (N_14232,N_13591,N_13559);
xor U14233 (N_14233,N_13515,N_13721);
nor U14234 (N_14234,N_13572,N_13664);
and U14235 (N_14235,N_13636,N_13654);
xnor U14236 (N_14236,N_13670,N_13546);
or U14237 (N_14237,N_13656,N_13233);
xnor U14238 (N_14238,N_13310,N_13452);
nor U14239 (N_14239,N_13371,N_13274);
nor U14240 (N_14240,N_13206,N_13374);
nand U14241 (N_14241,N_13448,N_13210);
nor U14242 (N_14242,N_13217,N_13240);
nand U14243 (N_14243,N_13606,N_13571);
or U14244 (N_14244,N_13573,N_13127);
or U14245 (N_14245,N_13621,N_13277);
and U14246 (N_14246,N_13488,N_13568);
nor U14247 (N_14247,N_13694,N_13356);
or U14248 (N_14248,N_13255,N_13441);
nand U14249 (N_14249,N_13342,N_13665);
and U14250 (N_14250,N_13619,N_13424);
nor U14251 (N_14251,N_13198,N_13388);
xnor U14252 (N_14252,N_13740,N_13145);
xor U14253 (N_14253,N_13155,N_13663);
or U14254 (N_14254,N_13691,N_13618);
xnor U14255 (N_14255,N_13169,N_13326);
or U14256 (N_14256,N_13742,N_13644);
nand U14257 (N_14257,N_13256,N_13507);
nand U14258 (N_14258,N_13499,N_13544);
xnor U14259 (N_14259,N_13517,N_13493);
and U14260 (N_14260,N_13216,N_13314);
xnor U14261 (N_14261,N_13479,N_13306);
xor U14262 (N_14262,N_13358,N_13515);
nand U14263 (N_14263,N_13717,N_13243);
nand U14264 (N_14264,N_13473,N_13617);
nand U14265 (N_14265,N_13550,N_13130);
nand U14266 (N_14266,N_13269,N_13253);
nor U14267 (N_14267,N_13668,N_13423);
or U14268 (N_14268,N_13207,N_13262);
or U14269 (N_14269,N_13174,N_13251);
xnor U14270 (N_14270,N_13571,N_13686);
and U14271 (N_14271,N_13520,N_13662);
and U14272 (N_14272,N_13652,N_13578);
and U14273 (N_14273,N_13490,N_13512);
or U14274 (N_14274,N_13549,N_13520);
and U14275 (N_14275,N_13705,N_13695);
and U14276 (N_14276,N_13134,N_13338);
or U14277 (N_14277,N_13510,N_13486);
nor U14278 (N_14278,N_13709,N_13612);
nor U14279 (N_14279,N_13725,N_13499);
and U14280 (N_14280,N_13704,N_13530);
nand U14281 (N_14281,N_13720,N_13565);
and U14282 (N_14282,N_13233,N_13276);
xnor U14283 (N_14283,N_13465,N_13499);
nand U14284 (N_14284,N_13261,N_13356);
xnor U14285 (N_14285,N_13693,N_13307);
and U14286 (N_14286,N_13202,N_13656);
nor U14287 (N_14287,N_13714,N_13305);
and U14288 (N_14288,N_13617,N_13437);
xnor U14289 (N_14289,N_13141,N_13284);
nand U14290 (N_14290,N_13631,N_13126);
and U14291 (N_14291,N_13527,N_13489);
or U14292 (N_14292,N_13743,N_13517);
xnor U14293 (N_14293,N_13171,N_13373);
nor U14294 (N_14294,N_13558,N_13436);
or U14295 (N_14295,N_13196,N_13504);
and U14296 (N_14296,N_13409,N_13280);
nor U14297 (N_14297,N_13255,N_13446);
nor U14298 (N_14298,N_13299,N_13477);
and U14299 (N_14299,N_13667,N_13581);
or U14300 (N_14300,N_13264,N_13171);
or U14301 (N_14301,N_13374,N_13598);
or U14302 (N_14302,N_13146,N_13337);
nand U14303 (N_14303,N_13567,N_13560);
and U14304 (N_14304,N_13193,N_13361);
and U14305 (N_14305,N_13284,N_13159);
nand U14306 (N_14306,N_13675,N_13611);
nand U14307 (N_14307,N_13661,N_13379);
nand U14308 (N_14308,N_13617,N_13556);
nand U14309 (N_14309,N_13480,N_13285);
nor U14310 (N_14310,N_13418,N_13727);
and U14311 (N_14311,N_13566,N_13667);
nand U14312 (N_14312,N_13495,N_13363);
nand U14313 (N_14313,N_13292,N_13206);
or U14314 (N_14314,N_13680,N_13720);
and U14315 (N_14315,N_13277,N_13390);
xnor U14316 (N_14316,N_13476,N_13316);
and U14317 (N_14317,N_13177,N_13561);
nor U14318 (N_14318,N_13457,N_13275);
xor U14319 (N_14319,N_13307,N_13562);
xnor U14320 (N_14320,N_13537,N_13217);
or U14321 (N_14321,N_13400,N_13551);
and U14322 (N_14322,N_13744,N_13521);
xnor U14323 (N_14323,N_13134,N_13294);
and U14324 (N_14324,N_13518,N_13599);
xor U14325 (N_14325,N_13223,N_13205);
nor U14326 (N_14326,N_13463,N_13377);
xor U14327 (N_14327,N_13419,N_13529);
and U14328 (N_14328,N_13453,N_13214);
nor U14329 (N_14329,N_13620,N_13380);
nand U14330 (N_14330,N_13279,N_13136);
and U14331 (N_14331,N_13609,N_13287);
nand U14332 (N_14332,N_13704,N_13731);
and U14333 (N_14333,N_13549,N_13691);
nor U14334 (N_14334,N_13558,N_13329);
nand U14335 (N_14335,N_13250,N_13289);
or U14336 (N_14336,N_13149,N_13274);
xor U14337 (N_14337,N_13502,N_13676);
nand U14338 (N_14338,N_13329,N_13243);
nand U14339 (N_14339,N_13626,N_13324);
nand U14340 (N_14340,N_13325,N_13180);
or U14341 (N_14341,N_13513,N_13710);
xor U14342 (N_14342,N_13723,N_13668);
xnor U14343 (N_14343,N_13244,N_13581);
nand U14344 (N_14344,N_13638,N_13175);
or U14345 (N_14345,N_13284,N_13322);
and U14346 (N_14346,N_13127,N_13265);
nor U14347 (N_14347,N_13166,N_13337);
xor U14348 (N_14348,N_13693,N_13597);
nor U14349 (N_14349,N_13249,N_13478);
or U14350 (N_14350,N_13537,N_13373);
nor U14351 (N_14351,N_13494,N_13609);
xor U14352 (N_14352,N_13749,N_13294);
or U14353 (N_14353,N_13745,N_13508);
nor U14354 (N_14354,N_13712,N_13351);
and U14355 (N_14355,N_13737,N_13493);
or U14356 (N_14356,N_13488,N_13691);
xor U14357 (N_14357,N_13698,N_13357);
nand U14358 (N_14358,N_13479,N_13686);
nand U14359 (N_14359,N_13546,N_13624);
nor U14360 (N_14360,N_13386,N_13719);
and U14361 (N_14361,N_13392,N_13657);
xor U14362 (N_14362,N_13613,N_13445);
nor U14363 (N_14363,N_13282,N_13216);
nor U14364 (N_14364,N_13656,N_13588);
xnor U14365 (N_14365,N_13287,N_13597);
xor U14366 (N_14366,N_13318,N_13483);
and U14367 (N_14367,N_13610,N_13735);
or U14368 (N_14368,N_13142,N_13473);
or U14369 (N_14369,N_13630,N_13252);
and U14370 (N_14370,N_13246,N_13394);
or U14371 (N_14371,N_13538,N_13596);
nor U14372 (N_14372,N_13128,N_13628);
nor U14373 (N_14373,N_13534,N_13403);
and U14374 (N_14374,N_13251,N_13722);
nand U14375 (N_14375,N_14331,N_14192);
or U14376 (N_14376,N_14338,N_13816);
nand U14377 (N_14377,N_14291,N_13967);
xor U14378 (N_14378,N_13889,N_14268);
xor U14379 (N_14379,N_14063,N_14285);
nor U14380 (N_14380,N_14178,N_13796);
nor U14381 (N_14381,N_14360,N_14145);
nand U14382 (N_14382,N_14201,N_13975);
nor U14383 (N_14383,N_13866,N_14196);
xor U14384 (N_14384,N_14177,N_14342);
xor U14385 (N_14385,N_14358,N_14209);
xnor U14386 (N_14386,N_14294,N_13873);
or U14387 (N_14387,N_14334,N_14295);
nand U14388 (N_14388,N_13973,N_14020);
and U14389 (N_14389,N_14003,N_14298);
nor U14390 (N_14390,N_14215,N_14127);
or U14391 (N_14391,N_14068,N_14310);
or U14392 (N_14392,N_14092,N_13789);
xor U14393 (N_14393,N_13867,N_13764);
nand U14394 (N_14394,N_14241,N_14278);
xor U14395 (N_14395,N_13946,N_13958);
and U14396 (N_14396,N_13872,N_14150);
nor U14397 (N_14397,N_13903,N_14151);
or U14398 (N_14398,N_14048,N_13959);
nor U14399 (N_14399,N_14040,N_14038);
or U14400 (N_14400,N_13882,N_14113);
and U14401 (N_14401,N_13979,N_14110);
nand U14402 (N_14402,N_14243,N_13910);
xor U14403 (N_14403,N_14042,N_13871);
xor U14404 (N_14404,N_14355,N_13931);
nand U14405 (N_14405,N_14045,N_14119);
xnor U14406 (N_14406,N_14115,N_14315);
nand U14407 (N_14407,N_13900,N_14262);
nor U14408 (N_14408,N_14330,N_14047);
nand U14409 (N_14409,N_13914,N_13842);
nand U14410 (N_14410,N_13806,N_14170);
or U14411 (N_14411,N_13916,N_13986);
nor U14412 (N_14412,N_13773,N_14302);
xnor U14413 (N_14413,N_14191,N_14190);
or U14414 (N_14414,N_13853,N_14299);
xnor U14415 (N_14415,N_13815,N_13972);
or U14416 (N_14416,N_14193,N_13995);
and U14417 (N_14417,N_14181,N_14146);
xnor U14418 (N_14418,N_13862,N_13854);
and U14419 (N_14419,N_13937,N_13798);
xnor U14420 (N_14420,N_13857,N_13952);
nand U14421 (N_14421,N_14025,N_13932);
nor U14422 (N_14422,N_13934,N_14004);
xnor U14423 (N_14423,N_14235,N_13938);
nand U14424 (N_14424,N_14072,N_14103);
nor U14425 (N_14425,N_13784,N_14325);
nand U14426 (N_14426,N_14129,N_13992);
or U14427 (N_14427,N_14001,N_14232);
nor U14428 (N_14428,N_14217,N_14288);
and U14429 (N_14429,N_14225,N_14261);
nand U14430 (N_14430,N_14227,N_13923);
or U14431 (N_14431,N_13943,N_14076);
and U14432 (N_14432,N_14273,N_13930);
and U14433 (N_14433,N_14208,N_13788);
xnor U14434 (N_14434,N_14237,N_14128);
or U14435 (N_14435,N_14252,N_14238);
nand U14436 (N_14436,N_14169,N_14300);
or U14437 (N_14437,N_14216,N_14030);
xor U14438 (N_14438,N_13817,N_14085);
xor U14439 (N_14439,N_14213,N_14155);
or U14440 (N_14440,N_13954,N_14000);
and U14441 (N_14441,N_14137,N_14140);
and U14442 (N_14442,N_13962,N_14319);
nand U14443 (N_14443,N_13905,N_14028);
nor U14444 (N_14444,N_13812,N_14173);
xnor U14445 (N_14445,N_13888,N_14199);
and U14446 (N_14446,N_14297,N_13845);
and U14447 (N_14447,N_13935,N_13841);
xnor U14448 (N_14448,N_14027,N_14158);
or U14449 (N_14449,N_13913,N_14323);
nand U14450 (N_14450,N_14075,N_13802);
and U14451 (N_14451,N_13790,N_14141);
or U14452 (N_14452,N_14050,N_13990);
and U14453 (N_14453,N_14182,N_14087);
or U14454 (N_14454,N_14185,N_14009);
xor U14455 (N_14455,N_13852,N_14200);
nand U14456 (N_14456,N_13980,N_14054);
or U14457 (N_14457,N_13901,N_13927);
xnor U14458 (N_14458,N_13880,N_13966);
xor U14459 (N_14459,N_14164,N_13947);
and U14460 (N_14460,N_14034,N_13826);
nand U14461 (N_14461,N_13821,N_13898);
nand U14462 (N_14462,N_14073,N_13771);
xor U14463 (N_14463,N_13890,N_14167);
and U14464 (N_14464,N_14100,N_14348);
nand U14465 (N_14465,N_14057,N_13761);
or U14466 (N_14466,N_14136,N_14174);
nor U14467 (N_14467,N_14371,N_14105);
xor U14468 (N_14468,N_13897,N_14283);
xnor U14469 (N_14469,N_14336,N_14008);
nand U14470 (N_14470,N_13831,N_14341);
or U14471 (N_14471,N_14352,N_14304);
nand U14472 (N_14472,N_14056,N_13843);
nor U14473 (N_14473,N_14257,N_14165);
xnor U14474 (N_14474,N_14359,N_13892);
nor U14475 (N_14475,N_14131,N_14039);
nand U14476 (N_14476,N_14220,N_13982);
or U14477 (N_14477,N_13860,N_14374);
nand U14478 (N_14478,N_14218,N_14249);
nor U14479 (N_14479,N_14312,N_13863);
nor U14480 (N_14480,N_14157,N_13865);
or U14481 (N_14481,N_13978,N_14077);
or U14482 (N_14482,N_13924,N_14007);
xor U14483 (N_14483,N_14154,N_14318);
and U14484 (N_14484,N_13988,N_13791);
and U14485 (N_14485,N_14244,N_13777);
or U14486 (N_14486,N_14260,N_14277);
nor U14487 (N_14487,N_14242,N_13787);
and U14488 (N_14488,N_14239,N_14287);
or U14489 (N_14489,N_13824,N_14326);
xor U14490 (N_14490,N_13908,N_14016);
nand U14491 (N_14491,N_14097,N_13752);
xnor U14492 (N_14492,N_14094,N_14067);
nor U14493 (N_14493,N_14281,N_14198);
or U14494 (N_14494,N_13756,N_13793);
nand U14495 (N_14495,N_13875,N_13754);
or U14496 (N_14496,N_14255,N_13844);
or U14497 (N_14497,N_13999,N_13835);
nor U14498 (N_14498,N_13837,N_14014);
xnor U14499 (N_14499,N_14301,N_13827);
nor U14500 (N_14500,N_14006,N_14250);
or U14501 (N_14501,N_13985,N_14161);
and U14502 (N_14502,N_14183,N_14373);
and U14503 (N_14503,N_14091,N_13770);
or U14504 (N_14504,N_14356,N_14248);
xor U14505 (N_14505,N_13762,N_13807);
nor U14506 (N_14506,N_14049,N_13885);
nand U14507 (N_14507,N_14284,N_14207);
or U14508 (N_14508,N_14274,N_14018);
xnor U14509 (N_14509,N_13769,N_13755);
nand U14510 (N_14510,N_14086,N_14149);
or U14511 (N_14511,N_14022,N_13895);
nor U14512 (N_14512,N_13783,N_14101);
xor U14513 (N_14513,N_13918,N_14187);
nor U14514 (N_14514,N_14079,N_13836);
nor U14515 (N_14515,N_13881,N_14143);
xor U14516 (N_14516,N_14132,N_14153);
xor U14517 (N_14517,N_13944,N_13981);
nor U14518 (N_14518,N_13832,N_14286);
and U14519 (N_14519,N_13922,N_14055);
nand U14520 (N_14520,N_14044,N_14052);
nor U14521 (N_14521,N_14245,N_14322);
nor U14522 (N_14522,N_13840,N_13781);
and U14523 (N_14523,N_14194,N_14060);
nand U14524 (N_14524,N_14074,N_14011);
xor U14525 (N_14525,N_14229,N_14234);
and U14526 (N_14526,N_13750,N_13948);
xor U14527 (N_14527,N_14083,N_14202);
or U14528 (N_14528,N_13998,N_14345);
nor U14529 (N_14529,N_13774,N_14353);
and U14530 (N_14530,N_13864,N_14370);
and U14531 (N_14531,N_14340,N_14139);
xor U14532 (N_14532,N_14166,N_14354);
nor U14533 (N_14533,N_13989,N_14171);
nor U14534 (N_14534,N_14362,N_14279);
and U14535 (N_14535,N_13818,N_14053);
xor U14536 (N_14536,N_13758,N_13780);
xor U14537 (N_14537,N_14184,N_14116);
or U14538 (N_14538,N_13759,N_14002);
or U14539 (N_14539,N_14095,N_13834);
nor U14540 (N_14540,N_14108,N_14046);
or U14541 (N_14541,N_14163,N_14176);
xor U14542 (N_14542,N_14061,N_14069);
xnor U14543 (N_14543,N_14264,N_13912);
nor U14544 (N_14544,N_14349,N_14320);
and U14545 (N_14545,N_14080,N_14270);
and U14546 (N_14546,N_13785,N_14346);
xor U14547 (N_14547,N_14321,N_13767);
xnor U14548 (N_14548,N_13760,N_14197);
nand U14549 (N_14549,N_13977,N_14021);
and U14550 (N_14550,N_14333,N_14082);
xnor U14551 (N_14551,N_13779,N_14147);
nand U14552 (N_14552,N_14271,N_14265);
xnor U14553 (N_14553,N_14263,N_13942);
and U14554 (N_14554,N_14316,N_14089);
nand U14555 (N_14555,N_14228,N_13951);
nor U14556 (N_14556,N_13878,N_14142);
and U14557 (N_14557,N_14123,N_14212);
and U14558 (N_14558,N_13765,N_13856);
or U14559 (N_14559,N_13768,N_13823);
and U14560 (N_14560,N_13829,N_13833);
and U14561 (N_14561,N_13949,N_14062);
nor U14562 (N_14562,N_14324,N_13820);
or U14563 (N_14563,N_14364,N_13969);
nor U14564 (N_14564,N_13955,N_13847);
xor U14565 (N_14565,N_13974,N_13961);
and U14566 (N_14566,N_13786,N_13803);
nor U14567 (N_14567,N_14081,N_14231);
xnor U14568 (N_14568,N_13772,N_13957);
nand U14569 (N_14569,N_14335,N_14272);
or U14570 (N_14570,N_13941,N_13929);
nor U14571 (N_14571,N_14107,N_13996);
or U14572 (N_14572,N_13849,N_14210);
xnor U14573 (N_14573,N_13838,N_14096);
or U14574 (N_14574,N_14357,N_14160);
nand U14575 (N_14575,N_14267,N_14180);
xnor U14576 (N_14576,N_13899,N_13921);
nand U14577 (N_14577,N_13994,N_14280);
nand U14578 (N_14578,N_14275,N_14203);
xnor U14579 (N_14579,N_13976,N_14306);
nand U14580 (N_14580,N_13907,N_14013);
or U14581 (N_14581,N_13868,N_13911);
and U14582 (N_14582,N_13876,N_13877);
xor U14583 (N_14583,N_14106,N_14204);
and U14584 (N_14584,N_13917,N_13776);
nor U14585 (N_14585,N_13984,N_14138);
and U14586 (N_14586,N_14365,N_14343);
or U14587 (N_14587,N_14254,N_14012);
and U14588 (N_14588,N_13993,N_14059);
xor U14589 (N_14589,N_14015,N_14032);
nand U14590 (N_14590,N_13808,N_13805);
or U14591 (N_14591,N_14019,N_14098);
nand U14592 (N_14592,N_13825,N_14033);
xor U14593 (N_14593,N_14292,N_13970);
nor U14594 (N_14594,N_13884,N_14226);
xnor U14595 (N_14595,N_14058,N_14120);
xor U14596 (N_14596,N_13757,N_14296);
and U14597 (N_14597,N_13983,N_14041);
or U14598 (N_14598,N_14328,N_14051);
and U14599 (N_14599,N_14367,N_14363);
or U14600 (N_14600,N_13850,N_14117);
nand U14601 (N_14601,N_14329,N_14112);
xnor U14602 (N_14602,N_14308,N_13775);
and U14603 (N_14603,N_14230,N_13902);
nor U14604 (N_14604,N_13939,N_14090);
nand U14605 (N_14605,N_14214,N_13861);
and U14606 (N_14606,N_13810,N_14369);
xnor U14607 (N_14607,N_13945,N_13940);
nor U14608 (N_14608,N_14099,N_14256);
nor U14609 (N_14609,N_13763,N_14293);
nand U14610 (N_14610,N_14188,N_14311);
and U14611 (N_14611,N_14289,N_13879);
or U14612 (N_14612,N_14347,N_14303);
and U14613 (N_14613,N_13953,N_14246);
and U14614 (N_14614,N_13830,N_14350);
nor U14615 (N_14615,N_14114,N_13920);
or U14616 (N_14616,N_14251,N_13960);
nor U14617 (N_14617,N_14031,N_13964);
nor U14618 (N_14618,N_14332,N_13887);
nand U14619 (N_14619,N_13987,N_14269);
or U14620 (N_14620,N_14071,N_14240);
or U14621 (N_14621,N_14314,N_14172);
and U14622 (N_14622,N_14253,N_14259);
nand U14623 (N_14623,N_13814,N_14327);
nor U14624 (N_14624,N_13971,N_14344);
nor U14625 (N_14625,N_14233,N_14372);
nand U14626 (N_14626,N_14064,N_13794);
or U14627 (N_14627,N_13968,N_13848);
nand U14628 (N_14628,N_13950,N_13869);
nand U14629 (N_14629,N_14189,N_13839);
nor U14630 (N_14630,N_13906,N_14043);
or U14631 (N_14631,N_13874,N_14035);
nor U14632 (N_14632,N_13804,N_14124);
nor U14633 (N_14633,N_13909,N_14339);
xnor U14634 (N_14634,N_14026,N_14084);
or U14635 (N_14635,N_14361,N_13926);
nor U14636 (N_14636,N_14118,N_14309);
xnor U14637 (N_14637,N_14266,N_14065);
nor U14638 (N_14638,N_14088,N_13799);
xnor U14639 (N_14639,N_13851,N_14305);
nor U14640 (N_14640,N_14135,N_14290);
and U14641 (N_14641,N_13919,N_14102);
nand U14642 (N_14642,N_14236,N_14125);
or U14643 (N_14643,N_14066,N_14156);
and U14644 (N_14644,N_13800,N_13828);
and U14645 (N_14645,N_13822,N_14134);
nor U14646 (N_14646,N_14206,N_14317);
nand U14647 (N_14647,N_14179,N_14104);
xor U14648 (N_14648,N_14005,N_13792);
nand U14649 (N_14649,N_14219,N_14221);
nor U14650 (N_14650,N_13855,N_14368);
nand U14651 (N_14651,N_14093,N_14313);
nor U14652 (N_14652,N_14010,N_14366);
nand U14653 (N_14653,N_13846,N_13766);
and U14654 (N_14654,N_13858,N_13859);
xor U14655 (N_14655,N_13778,N_13813);
nor U14656 (N_14656,N_13956,N_14036);
and U14657 (N_14657,N_13883,N_14111);
xor U14658 (N_14658,N_14282,N_14121);
or U14659 (N_14659,N_14023,N_13896);
nor U14660 (N_14660,N_14247,N_13894);
or U14661 (N_14661,N_13928,N_14029);
and U14662 (N_14662,N_14133,N_14152);
xnor U14663 (N_14663,N_13801,N_14307);
and U14664 (N_14664,N_14276,N_13809);
and U14665 (N_14665,N_14168,N_14126);
and U14666 (N_14666,N_14337,N_13915);
and U14667 (N_14667,N_14078,N_14037);
or U14668 (N_14668,N_14195,N_13751);
and U14669 (N_14669,N_13891,N_14175);
nor U14670 (N_14670,N_13997,N_14223);
or U14671 (N_14671,N_14130,N_14109);
or U14672 (N_14672,N_14162,N_13811);
xor U14673 (N_14673,N_14224,N_14144);
xnor U14674 (N_14674,N_13936,N_14222);
or U14675 (N_14675,N_14017,N_13870);
and U14676 (N_14676,N_14024,N_13965);
xnor U14677 (N_14677,N_14258,N_13933);
and U14678 (N_14678,N_13797,N_14211);
and U14679 (N_14679,N_13819,N_13963);
nor U14680 (N_14680,N_14159,N_13782);
xor U14681 (N_14681,N_14351,N_14205);
nor U14682 (N_14682,N_14186,N_13893);
nand U14683 (N_14683,N_13795,N_14122);
and U14684 (N_14684,N_13753,N_13886);
nor U14685 (N_14685,N_14148,N_13925);
nor U14686 (N_14686,N_13991,N_13904);
nand U14687 (N_14687,N_14070,N_14030);
nand U14688 (N_14688,N_14075,N_13989);
and U14689 (N_14689,N_13974,N_13991);
and U14690 (N_14690,N_13786,N_14313);
and U14691 (N_14691,N_13782,N_13995);
and U14692 (N_14692,N_13934,N_13949);
nand U14693 (N_14693,N_13803,N_13752);
nand U14694 (N_14694,N_13891,N_14035);
and U14695 (N_14695,N_13894,N_14257);
or U14696 (N_14696,N_13762,N_14077);
xor U14697 (N_14697,N_14067,N_13817);
xor U14698 (N_14698,N_14067,N_13836);
nor U14699 (N_14699,N_13862,N_14276);
nor U14700 (N_14700,N_13793,N_14241);
and U14701 (N_14701,N_14268,N_14057);
or U14702 (N_14702,N_14081,N_14325);
nand U14703 (N_14703,N_14362,N_13786);
and U14704 (N_14704,N_14057,N_14357);
nand U14705 (N_14705,N_13845,N_13775);
and U14706 (N_14706,N_13834,N_14092);
nand U14707 (N_14707,N_13957,N_14120);
xnor U14708 (N_14708,N_14344,N_13983);
nand U14709 (N_14709,N_14246,N_13952);
nor U14710 (N_14710,N_13813,N_14329);
nand U14711 (N_14711,N_14184,N_14143);
xor U14712 (N_14712,N_14357,N_14203);
or U14713 (N_14713,N_14151,N_14261);
and U14714 (N_14714,N_14069,N_14336);
or U14715 (N_14715,N_14116,N_13987);
and U14716 (N_14716,N_14362,N_13977);
nand U14717 (N_14717,N_14262,N_14227);
or U14718 (N_14718,N_14301,N_14179);
xnor U14719 (N_14719,N_13903,N_14227);
nor U14720 (N_14720,N_14056,N_14101);
xnor U14721 (N_14721,N_13990,N_13988);
nor U14722 (N_14722,N_13830,N_14258);
and U14723 (N_14723,N_14293,N_14142);
nor U14724 (N_14724,N_14168,N_14270);
xnor U14725 (N_14725,N_13883,N_14274);
or U14726 (N_14726,N_13826,N_13868);
nor U14727 (N_14727,N_14108,N_14352);
xnor U14728 (N_14728,N_13951,N_14058);
xnor U14729 (N_14729,N_14139,N_14213);
nor U14730 (N_14730,N_14284,N_13986);
and U14731 (N_14731,N_14142,N_13962);
or U14732 (N_14732,N_13806,N_14186);
nor U14733 (N_14733,N_14249,N_14280);
nand U14734 (N_14734,N_13817,N_14337);
and U14735 (N_14735,N_13790,N_14368);
and U14736 (N_14736,N_14265,N_14022);
and U14737 (N_14737,N_14293,N_14110);
nor U14738 (N_14738,N_14229,N_13797);
and U14739 (N_14739,N_13829,N_14117);
nand U14740 (N_14740,N_14044,N_14021);
nand U14741 (N_14741,N_14136,N_14167);
xor U14742 (N_14742,N_13908,N_13848);
or U14743 (N_14743,N_13756,N_13759);
nor U14744 (N_14744,N_13844,N_14105);
nand U14745 (N_14745,N_13807,N_14003);
xnor U14746 (N_14746,N_14153,N_14150);
xor U14747 (N_14747,N_14116,N_13964);
and U14748 (N_14748,N_14132,N_13811);
nand U14749 (N_14749,N_14199,N_14302);
nor U14750 (N_14750,N_14223,N_14294);
nand U14751 (N_14751,N_14362,N_14168);
xor U14752 (N_14752,N_13960,N_14271);
or U14753 (N_14753,N_13766,N_14245);
or U14754 (N_14754,N_14109,N_14263);
or U14755 (N_14755,N_14064,N_14170);
xnor U14756 (N_14756,N_14051,N_13909);
and U14757 (N_14757,N_13953,N_14267);
or U14758 (N_14758,N_13890,N_14098);
xnor U14759 (N_14759,N_14349,N_14242);
or U14760 (N_14760,N_14142,N_13806);
nand U14761 (N_14761,N_13854,N_13987);
nor U14762 (N_14762,N_14244,N_14053);
and U14763 (N_14763,N_13872,N_14165);
xor U14764 (N_14764,N_13895,N_13759);
xnor U14765 (N_14765,N_14356,N_13837);
nor U14766 (N_14766,N_13917,N_13943);
nor U14767 (N_14767,N_14360,N_14020);
and U14768 (N_14768,N_14280,N_14248);
xor U14769 (N_14769,N_14286,N_14173);
or U14770 (N_14770,N_13806,N_13980);
xor U14771 (N_14771,N_13882,N_14269);
nor U14772 (N_14772,N_13902,N_13773);
nor U14773 (N_14773,N_14278,N_13807);
xnor U14774 (N_14774,N_14122,N_14198);
nor U14775 (N_14775,N_14354,N_13984);
or U14776 (N_14776,N_14037,N_14212);
nor U14777 (N_14777,N_13776,N_13860);
and U14778 (N_14778,N_13929,N_14256);
nor U14779 (N_14779,N_14109,N_14234);
and U14780 (N_14780,N_13964,N_14124);
nand U14781 (N_14781,N_13792,N_13806);
and U14782 (N_14782,N_14154,N_13838);
and U14783 (N_14783,N_14238,N_14228);
or U14784 (N_14784,N_13875,N_13877);
and U14785 (N_14785,N_14241,N_14007);
xor U14786 (N_14786,N_13868,N_14027);
nand U14787 (N_14787,N_14357,N_13999);
xnor U14788 (N_14788,N_14074,N_14148);
or U14789 (N_14789,N_14267,N_13882);
nor U14790 (N_14790,N_13889,N_14065);
nor U14791 (N_14791,N_13983,N_13991);
and U14792 (N_14792,N_13808,N_14299);
nor U14793 (N_14793,N_14311,N_13927);
or U14794 (N_14794,N_13824,N_13946);
and U14795 (N_14795,N_13979,N_14252);
nand U14796 (N_14796,N_14038,N_13779);
nor U14797 (N_14797,N_13930,N_14055);
xor U14798 (N_14798,N_14056,N_14171);
or U14799 (N_14799,N_14069,N_14059);
xor U14800 (N_14800,N_13878,N_14125);
or U14801 (N_14801,N_14310,N_14326);
and U14802 (N_14802,N_13819,N_14216);
and U14803 (N_14803,N_14120,N_13801);
or U14804 (N_14804,N_13929,N_13936);
nand U14805 (N_14805,N_14348,N_14088);
and U14806 (N_14806,N_14097,N_13763);
and U14807 (N_14807,N_13891,N_14064);
nor U14808 (N_14808,N_13770,N_14256);
xnor U14809 (N_14809,N_14058,N_14322);
nor U14810 (N_14810,N_14345,N_14107);
nor U14811 (N_14811,N_13797,N_14274);
nor U14812 (N_14812,N_14009,N_14093);
nor U14813 (N_14813,N_14191,N_14311);
xor U14814 (N_14814,N_13832,N_13908);
nor U14815 (N_14815,N_13878,N_14112);
or U14816 (N_14816,N_14257,N_13840);
xor U14817 (N_14817,N_14272,N_14147);
xnor U14818 (N_14818,N_13790,N_14326);
and U14819 (N_14819,N_14085,N_13925);
nor U14820 (N_14820,N_14336,N_13781);
and U14821 (N_14821,N_14124,N_14341);
nor U14822 (N_14822,N_14227,N_13874);
or U14823 (N_14823,N_14006,N_14234);
nand U14824 (N_14824,N_14268,N_13898);
and U14825 (N_14825,N_14062,N_13953);
or U14826 (N_14826,N_14298,N_14018);
and U14827 (N_14827,N_14253,N_14330);
or U14828 (N_14828,N_14253,N_14372);
and U14829 (N_14829,N_14016,N_14280);
and U14830 (N_14830,N_14114,N_13874);
or U14831 (N_14831,N_13953,N_14084);
or U14832 (N_14832,N_13798,N_14104);
and U14833 (N_14833,N_14086,N_14232);
and U14834 (N_14834,N_13852,N_13841);
or U14835 (N_14835,N_14238,N_14348);
and U14836 (N_14836,N_14128,N_14028);
or U14837 (N_14837,N_13783,N_14001);
xnor U14838 (N_14838,N_14123,N_14096);
and U14839 (N_14839,N_13983,N_14317);
nor U14840 (N_14840,N_14221,N_14279);
nand U14841 (N_14841,N_13815,N_14039);
or U14842 (N_14842,N_13954,N_14042);
nor U14843 (N_14843,N_14050,N_14099);
nand U14844 (N_14844,N_14294,N_14056);
or U14845 (N_14845,N_14014,N_13791);
nor U14846 (N_14846,N_14151,N_14213);
and U14847 (N_14847,N_14109,N_14148);
and U14848 (N_14848,N_13906,N_13777);
and U14849 (N_14849,N_14062,N_13890);
or U14850 (N_14850,N_14264,N_13951);
and U14851 (N_14851,N_14159,N_14221);
and U14852 (N_14852,N_14197,N_14365);
nor U14853 (N_14853,N_13779,N_14141);
or U14854 (N_14854,N_14099,N_13901);
and U14855 (N_14855,N_14231,N_14053);
xnor U14856 (N_14856,N_14292,N_14049);
and U14857 (N_14857,N_14057,N_14051);
nor U14858 (N_14858,N_13824,N_14268);
xnor U14859 (N_14859,N_13833,N_14022);
nor U14860 (N_14860,N_14311,N_14102);
and U14861 (N_14861,N_14128,N_13872);
nand U14862 (N_14862,N_13851,N_13799);
nand U14863 (N_14863,N_13961,N_14221);
and U14864 (N_14864,N_13822,N_13775);
nand U14865 (N_14865,N_13881,N_14076);
and U14866 (N_14866,N_14019,N_14163);
and U14867 (N_14867,N_14240,N_13874);
nor U14868 (N_14868,N_13945,N_14039);
and U14869 (N_14869,N_14003,N_14309);
or U14870 (N_14870,N_14195,N_14298);
xnor U14871 (N_14871,N_14115,N_14011);
nand U14872 (N_14872,N_13755,N_13906);
and U14873 (N_14873,N_13910,N_13920);
nand U14874 (N_14874,N_14099,N_13777);
nor U14875 (N_14875,N_13937,N_14218);
nor U14876 (N_14876,N_14296,N_13958);
and U14877 (N_14877,N_14101,N_13833);
nor U14878 (N_14878,N_14111,N_14052);
xor U14879 (N_14879,N_13988,N_14059);
or U14880 (N_14880,N_14173,N_14030);
nor U14881 (N_14881,N_14271,N_13753);
and U14882 (N_14882,N_13796,N_14256);
or U14883 (N_14883,N_14171,N_13855);
nand U14884 (N_14884,N_13987,N_13846);
nand U14885 (N_14885,N_14210,N_14099);
and U14886 (N_14886,N_14106,N_13845);
nand U14887 (N_14887,N_14316,N_13978);
nand U14888 (N_14888,N_14144,N_13762);
and U14889 (N_14889,N_14040,N_14033);
and U14890 (N_14890,N_14073,N_13839);
xor U14891 (N_14891,N_14355,N_13806);
nor U14892 (N_14892,N_13789,N_13995);
xnor U14893 (N_14893,N_14320,N_14079);
nor U14894 (N_14894,N_13904,N_14256);
and U14895 (N_14895,N_14351,N_13807);
nor U14896 (N_14896,N_14360,N_14316);
and U14897 (N_14897,N_13777,N_14046);
and U14898 (N_14898,N_13796,N_14196);
and U14899 (N_14899,N_14002,N_14192);
nand U14900 (N_14900,N_13835,N_13924);
and U14901 (N_14901,N_14190,N_13784);
and U14902 (N_14902,N_13990,N_14166);
xor U14903 (N_14903,N_14072,N_13893);
and U14904 (N_14904,N_13783,N_14116);
nand U14905 (N_14905,N_14092,N_14016);
nand U14906 (N_14906,N_14307,N_13948);
or U14907 (N_14907,N_14309,N_14177);
xnor U14908 (N_14908,N_13774,N_14325);
xnor U14909 (N_14909,N_14031,N_14306);
and U14910 (N_14910,N_14172,N_14164);
nor U14911 (N_14911,N_14101,N_13957);
or U14912 (N_14912,N_13864,N_13847);
nor U14913 (N_14913,N_14199,N_14313);
or U14914 (N_14914,N_14132,N_13948);
or U14915 (N_14915,N_14128,N_14169);
or U14916 (N_14916,N_14095,N_14069);
xor U14917 (N_14917,N_14360,N_13762);
nand U14918 (N_14918,N_13807,N_13995);
and U14919 (N_14919,N_14073,N_14037);
nor U14920 (N_14920,N_14086,N_14301);
nor U14921 (N_14921,N_14217,N_14214);
nor U14922 (N_14922,N_14318,N_14221);
and U14923 (N_14923,N_14103,N_13798);
xnor U14924 (N_14924,N_13764,N_14307);
and U14925 (N_14925,N_14304,N_13964);
nor U14926 (N_14926,N_13825,N_14330);
or U14927 (N_14927,N_14148,N_14233);
or U14928 (N_14928,N_13851,N_14085);
xor U14929 (N_14929,N_14329,N_13943);
nand U14930 (N_14930,N_14057,N_14285);
xnor U14931 (N_14931,N_14167,N_14292);
nor U14932 (N_14932,N_13776,N_14004);
or U14933 (N_14933,N_14142,N_13991);
or U14934 (N_14934,N_14232,N_14035);
and U14935 (N_14935,N_14146,N_14318);
nand U14936 (N_14936,N_13806,N_14341);
nand U14937 (N_14937,N_14005,N_13876);
or U14938 (N_14938,N_13948,N_14028);
xor U14939 (N_14939,N_14271,N_13855);
or U14940 (N_14940,N_13846,N_14109);
xor U14941 (N_14941,N_13878,N_13818);
xor U14942 (N_14942,N_14223,N_14364);
and U14943 (N_14943,N_13915,N_13818);
xor U14944 (N_14944,N_13994,N_13950);
nor U14945 (N_14945,N_14028,N_14052);
or U14946 (N_14946,N_14055,N_14145);
nor U14947 (N_14947,N_13892,N_14305);
and U14948 (N_14948,N_13751,N_13910);
nor U14949 (N_14949,N_13792,N_14242);
and U14950 (N_14950,N_13928,N_14229);
or U14951 (N_14951,N_14110,N_14115);
nand U14952 (N_14952,N_14190,N_13768);
or U14953 (N_14953,N_13968,N_14204);
or U14954 (N_14954,N_14125,N_14170);
and U14955 (N_14955,N_13913,N_14147);
nor U14956 (N_14956,N_13985,N_14261);
or U14957 (N_14957,N_13820,N_14227);
or U14958 (N_14958,N_13969,N_14245);
or U14959 (N_14959,N_13755,N_14078);
and U14960 (N_14960,N_13917,N_13813);
xnor U14961 (N_14961,N_14277,N_14009);
xor U14962 (N_14962,N_14291,N_13878);
xor U14963 (N_14963,N_13797,N_14154);
and U14964 (N_14964,N_13857,N_14332);
xor U14965 (N_14965,N_14147,N_14031);
and U14966 (N_14966,N_14116,N_13806);
nand U14967 (N_14967,N_13771,N_14245);
xor U14968 (N_14968,N_14293,N_14044);
nand U14969 (N_14969,N_13984,N_13922);
xnor U14970 (N_14970,N_13821,N_13760);
nor U14971 (N_14971,N_13773,N_13797);
nor U14972 (N_14972,N_14212,N_14059);
xor U14973 (N_14973,N_14049,N_14040);
and U14974 (N_14974,N_13820,N_13956);
or U14975 (N_14975,N_14074,N_14062);
nand U14976 (N_14976,N_14345,N_14159);
or U14977 (N_14977,N_14121,N_14076);
xnor U14978 (N_14978,N_14143,N_13868);
or U14979 (N_14979,N_13824,N_14369);
nand U14980 (N_14980,N_14226,N_14044);
or U14981 (N_14981,N_14037,N_14338);
and U14982 (N_14982,N_13937,N_14101);
xnor U14983 (N_14983,N_13976,N_14119);
xnor U14984 (N_14984,N_13940,N_13850);
nand U14985 (N_14985,N_13764,N_14218);
nor U14986 (N_14986,N_13853,N_13861);
nand U14987 (N_14987,N_13903,N_14290);
xor U14988 (N_14988,N_13823,N_14197);
xnor U14989 (N_14989,N_14147,N_13799);
nor U14990 (N_14990,N_14350,N_13986);
nand U14991 (N_14991,N_13978,N_13827);
or U14992 (N_14992,N_13881,N_14258);
or U14993 (N_14993,N_14109,N_14289);
nand U14994 (N_14994,N_14162,N_14280);
nand U14995 (N_14995,N_14130,N_13760);
nand U14996 (N_14996,N_14261,N_14000);
or U14997 (N_14997,N_14101,N_14164);
nor U14998 (N_14998,N_14210,N_13786);
nor U14999 (N_14999,N_14032,N_14219);
nor U15000 (N_15000,N_14517,N_14912);
xor U15001 (N_15001,N_14787,N_14878);
nor U15002 (N_15002,N_14997,N_14472);
nor U15003 (N_15003,N_14768,N_14563);
nor U15004 (N_15004,N_14750,N_14614);
nand U15005 (N_15005,N_14437,N_14970);
nor U15006 (N_15006,N_14536,N_14816);
xnor U15007 (N_15007,N_14735,N_14739);
xor U15008 (N_15008,N_14705,N_14741);
nor U15009 (N_15009,N_14937,N_14594);
nor U15010 (N_15010,N_14829,N_14539);
xnor U15011 (N_15011,N_14841,N_14974);
nor U15012 (N_15012,N_14984,N_14958);
nand U15013 (N_15013,N_14480,N_14637);
or U15014 (N_15014,N_14682,N_14434);
nand U15015 (N_15015,N_14522,N_14857);
xnor U15016 (N_15016,N_14504,N_14486);
xnor U15017 (N_15017,N_14807,N_14385);
nor U15018 (N_15018,N_14846,N_14665);
xor U15019 (N_15019,N_14950,N_14773);
nor U15020 (N_15020,N_14917,N_14496);
or U15021 (N_15021,N_14985,N_14798);
nor U15022 (N_15022,N_14456,N_14626);
nand U15023 (N_15023,N_14944,N_14545);
nor U15024 (N_15024,N_14991,N_14598);
and U15025 (N_15025,N_14489,N_14929);
nand U15026 (N_15026,N_14891,N_14879);
and U15027 (N_15027,N_14964,N_14611);
xnor U15028 (N_15028,N_14689,N_14875);
nand U15029 (N_15029,N_14613,N_14534);
or U15030 (N_15030,N_14884,N_14444);
or U15031 (N_15031,N_14653,N_14723);
or U15032 (N_15032,N_14445,N_14926);
nand U15033 (N_15033,N_14392,N_14943);
and U15034 (N_15034,N_14609,N_14453);
xor U15035 (N_15035,N_14419,N_14428);
and U15036 (N_15036,N_14420,N_14721);
nand U15037 (N_15037,N_14696,N_14743);
or U15038 (N_15038,N_14572,N_14492);
nand U15039 (N_15039,N_14503,N_14400);
xor U15040 (N_15040,N_14410,N_14767);
xnor U15041 (N_15041,N_14792,N_14936);
nand U15042 (N_15042,N_14688,N_14484);
or U15043 (N_15043,N_14574,N_14691);
nor U15044 (N_15044,N_14528,N_14401);
nor U15045 (N_15045,N_14899,N_14758);
xor U15046 (N_15046,N_14999,N_14458);
and U15047 (N_15047,N_14729,N_14703);
xor U15048 (N_15048,N_14890,N_14407);
and U15049 (N_15049,N_14821,N_14905);
and U15050 (N_15050,N_14830,N_14606);
nor U15051 (N_15051,N_14479,N_14904);
and U15052 (N_15052,N_14514,N_14652);
and U15053 (N_15053,N_14789,N_14498);
nand U15054 (N_15054,N_14663,N_14780);
xnor U15055 (N_15055,N_14529,N_14477);
nand U15056 (N_15056,N_14763,N_14967);
and U15057 (N_15057,N_14892,N_14389);
xor U15058 (N_15058,N_14629,N_14955);
and U15059 (N_15059,N_14757,N_14927);
nand U15060 (N_15060,N_14465,N_14685);
or U15061 (N_15061,N_14661,N_14402);
nor U15062 (N_15062,N_14491,N_14880);
nand U15063 (N_15063,N_14573,N_14908);
or U15064 (N_15064,N_14715,N_14897);
and U15065 (N_15065,N_14725,N_14433);
xnor U15066 (N_15066,N_14840,N_14759);
nand U15067 (N_15067,N_14803,N_14508);
or U15068 (N_15068,N_14426,N_14968);
or U15069 (N_15069,N_14543,N_14646);
or U15070 (N_15070,N_14393,N_14707);
or U15071 (N_15071,N_14894,N_14555);
nand U15072 (N_15072,N_14421,N_14441);
nand U15073 (N_15073,N_14699,N_14954);
nand U15074 (N_15074,N_14923,N_14702);
xor U15075 (N_15075,N_14581,N_14435);
xnor U15076 (N_15076,N_14717,N_14404);
xor U15077 (N_15077,N_14375,N_14537);
or U15078 (N_15078,N_14980,N_14616);
and U15079 (N_15079,N_14916,N_14505);
nand U15080 (N_15080,N_14521,N_14720);
xnor U15081 (N_15081,N_14793,N_14726);
xor U15082 (N_15082,N_14818,N_14672);
nor U15083 (N_15083,N_14599,N_14542);
nand U15084 (N_15084,N_14494,N_14675);
or U15085 (N_15085,N_14893,N_14648);
nor U15086 (N_15086,N_14823,N_14815);
or U15087 (N_15087,N_14583,N_14576);
or U15088 (N_15088,N_14651,N_14742);
and U15089 (N_15089,N_14906,N_14507);
nor U15090 (N_15090,N_14495,N_14774);
or U15091 (N_15091,N_14547,N_14982);
or U15092 (N_15092,N_14799,N_14451);
and U15093 (N_15093,N_14473,N_14633);
or U15094 (N_15094,N_14518,N_14485);
xor U15095 (N_15095,N_14765,N_14832);
nor U15096 (N_15096,N_14632,N_14975);
or U15097 (N_15097,N_14783,N_14570);
nand U15098 (N_15098,N_14475,N_14378);
nand U15099 (N_15099,N_14895,N_14887);
nand U15100 (N_15100,N_14901,N_14928);
nor U15101 (N_15101,N_14949,N_14603);
and U15102 (N_15102,N_14564,N_14714);
nor U15103 (N_15103,N_14940,N_14966);
or U15104 (N_15104,N_14851,N_14585);
nand U15105 (N_15105,N_14921,N_14865);
nor U15106 (N_15106,N_14462,N_14448);
or U15107 (N_15107,N_14990,N_14744);
xnor U15108 (N_15108,N_14670,N_14946);
xor U15109 (N_15109,N_14413,N_14788);
xnor U15110 (N_15110,N_14582,N_14394);
xnor U15111 (N_15111,N_14687,N_14450);
xnor U15112 (N_15112,N_14578,N_14858);
and U15113 (N_15113,N_14838,N_14464);
xnor U15114 (N_15114,N_14595,N_14716);
and U15115 (N_15115,N_14446,N_14808);
nand U15116 (N_15116,N_14822,N_14784);
nor U15117 (N_15117,N_14403,N_14845);
nor U15118 (N_15118,N_14883,N_14515);
or U15119 (N_15119,N_14754,N_14796);
nand U15120 (N_15120,N_14551,N_14463);
or U15121 (N_15121,N_14820,N_14849);
xnor U15122 (N_15122,N_14843,N_14377);
xor U15123 (N_15123,N_14751,N_14738);
nand U15124 (N_15124,N_14761,N_14527);
nand U15125 (N_15125,N_14384,N_14532);
nand U15126 (N_15126,N_14566,N_14919);
nor U15127 (N_15127,N_14416,N_14634);
or U15128 (N_15128,N_14510,N_14449);
nor U15129 (N_15129,N_14910,N_14794);
and U15130 (N_15130,N_14658,N_14642);
and U15131 (N_15131,N_14933,N_14902);
xnor U15132 (N_15132,N_14482,N_14736);
nor U15133 (N_15133,N_14452,N_14719);
and U15134 (N_15134,N_14546,N_14429);
nor U15135 (N_15135,N_14601,N_14650);
nand U15136 (N_15136,N_14544,N_14502);
and U15137 (N_15137,N_14698,N_14431);
nor U15138 (N_15138,N_14630,N_14568);
nand U15139 (N_15139,N_14605,N_14760);
nor U15140 (N_15140,N_14981,N_14922);
xor U15141 (N_15141,N_14395,N_14959);
xnor U15142 (N_15142,N_14415,N_14524);
and U15143 (N_15143,N_14882,N_14935);
or U15144 (N_15144,N_14580,N_14994);
xor U15145 (N_15145,N_14800,N_14679);
nand U15146 (N_15146,N_14842,N_14730);
nor U15147 (N_15147,N_14628,N_14978);
or U15148 (N_15148,N_14733,N_14836);
and U15149 (N_15149,N_14483,N_14931);
or U15150 (N_15150,N_14835,N_14710);
or U15151 (N_15151,N_14971,N_14942);
nand U15152 (N_15152,N_14562,N_14864);
xnor U15153 (N_15153,N_14686,N_14938);
and U15154 (N_15154,N_14775,N_14602);
or U15155 (N_15155,N_14561,N_14681);
and U15156 (N_15156,N_14874,N_14678);
and U15157 (N_15157,N_14885,N_14749);
nor U15158 (N_15158,N_14487,N_14951);
xor U15159 (N_15159,N_14660,N_14525);
nor U15160 (N_15160,N_14376,N_14781);
and U15161 (N_15161,N_14700,N_14727);
or U15162 (N_15162,N_14918,N_14817);
and U15163 (N_15163,N_14383,N_14764);
or U15164 (N_15164,N_14693,N_14722);
and U15165 (N_15165,N_14590,N_14530);
and U15166 (N_15166,N_14618,N_14638);
or U15167 (N_15167,N_14565,N_14497);
or U15168 (N_15168,N_14855,N_14856);
and U15169 (N_15169,N_14569,N_14776);
nor U15170 (N_15170,N_14501,N_14839);
or U15171 (N_15171,N_14423,N_14621);
nand U15172 (N_15172,N_14641,N_14945);
and U15173 (N_15173,N_14493,N_14915);
nand U15174 (N_15174,N_14557,N_14947);
xnor U15175 (N_15175,N_14417,N_14844);
and U15176 (N_15176,N_14512,N_14459);
nor U15177 (N_15177,N_14554,N_14649);
xnor U15178 (N_15178,N_14996,N_14695);
xor U15179 (N_15179,N_14831,N_14668);
xnor U15180 (N_15180,N_14584,N_14674);
xnor U15181 (N_15181,N_14548,N_14506);
and U15182 (N_15182,N_14778,N_14860);
nor U15183 (N_15183,N_14397,N_14867);
or U15184 (N_15184,N_14828,N_14706);
and U15185 (N_15185,N_14834,N_14871);
nand U15186 (N_15186,N_14677,N_14430);
nand U15187 (N_15187,N_14382,N_14939);
and U15188 (N_15188,N_14694,N_14387);
and U15189 (N_15189,N_14439,N_14556);
and U15190 (N_15190,N_14523,N_14690);
nand U15191 (N_15191,N_14888,N_14934);
and U15192 (N_15192,N_14791,N_14619);
and U15193 (N_15193,N_14969,N_14913);
or U15194 (N_15194,N_14734,N_14825);
xor U15195 (N_15195,N_14627,N_14398);
xor U15196 (N_15196,N_14457,N_14511);
nor U15197 (N_15197,N_14586,N_14593);
nand U15198 (N_15198,N_14531,N_14443);
and U15199 (N_15199,N_14909,N_14617);
or U15200 (N_15200,N_14709,N_14782);
and U15201 (N_15201,N_14388,N_14639);
and U15202 (N_15202,N_14405,N_14805);
or U15203 (N_15203,N_14588,N_14802);
xnor U15204 (N_15204,N_14771,N_14610);
nand U15205 (N_15205,N_14645,N_14673);
xnor U15206 (N_15206,N_14474,N_14728);
or U15207 (N_15207,N_14655,N_14833);
or U15208 (N_15208,N_14711,N_14785);
or U15209 (N_15209,N_14809,N_14769);
or U15210 (N_15210,N_14553,N_14671);
or U15211 (N_15211,N_14797,N_14541);
nand U15212 (N_15212,N_14560,N_14806);
and U15213 (N_15213,N_14635,N_14659);
and U15214 (N_15214,N_14708,N_14914);
nor U15215 (N_15215,N_14526,N_14408);
or U15216 (N_15216,N_14516,N_14869);
and U15217 (N_15217,N_14664,N_14762);
or U15218 (N_15218,N_14684,N_14591);
nand U15219 (N_15219,N_14826,N_14697);
nor U15220 (N_15220,N_14680,N_14747);
nor U15221 (N_15221,N_14713,N_14461);
nand U15222 (N_15222,N_14795,N_14746);
nand U15223 (N_15223,N_14724,N_14881);
nor U15224 (N_15224,N_14988,N_14704);
nor U15225 (N_15225,N_14827,N_14779);
nand U15226 (N_15226,N_14889,N_14538);
and U15227 (N_15227,N_14625,N_14965);
nand U15228 (N_15228,N_14676,N_14427);
nor U15229 (N_15229,N_14752,N_14962);
or U15230 (N_15230,N_14533,N_14712);
nand U15231 (N_15231,N_14932,N_14786);
and U15232 (N_15232,N_14930,N_14737);
or U15233 (N_15233,N_14732,N_14740);
nand U15234 (N_15234,N_14812,N_14440);
and U15235 (N_15235,N_14853,N_14587);
or U15236 (N_15236,N_14748,N_14669);
xor U15237 (N_15237,N_14953,N_14549);
nand U15238 (N_15238,N_14963,N_14579);
and U15239 (N_15239,N_14592,N_14900);
nor U15240 (N_15240,N_14837,N_14575);
and U15241 (N_15241,N_14643,N_14876);
xnor U15242 (N_15242,N_14607,N_14924);
and U15243 (N_15243,N_14907,N_14386);
or U15244 (N_15244,N_14519,N_14535);
xor U15245 (N_15245,N_14972,N_14973);
nor U15246 (N_15246,N_14667,N_14868);
or U15247 (N_15247,N_14960,N_14847);
and U15248 (N_15248,N_14471,N_14468);
or U15249 (N_15249,N_14490,N_14396);
xnor U15250 (N_15250,N_14854,N_14552);
xnor U15251 (N_15251,N_14436,N_14731);
nor U15252 (N_15252,N_14500,N_14470);
xor U15253 (N_15253,N_14540,N_14425);
or U15254 (N_15254,N_14753,N_14391);
xor U15255 (N_15255,N_14432,N_14819);
nor U15256 (N_15256,N_14612,N_14872);
nand U15257 (N_15257,N_14692,N_14509);
and U15258 (N_15258,N_14801,N_14772);
and U15259 (N_15259,N_14813,N_14811);
xor U15260 (N_15260,N_14488,N_14852);
or U15261 (N_15261,N_14476,N_14898);
or U15262 (N_15262,N_14615,N_14466);
nand U15263 (N_15263,N_14409,N_14948);
xor U15264 (N_15264,N_14956,N_14756);
or U15265 (N_15265,N_14604,N_14631);
or U15266 (N_15266,N_14380,N_14447);
or U15267 (N_15267,N_14412,N_14666);
or U15268 (N_15268,N_14422,N_14640);
or U15269 (N_15269,N_14993,N_14862);
and U15270 (N_15270,N_14810,N_14877);
xor U15271 (N_15271,N_14873,N_14998);
or U15272 (N_15272,N_14636,N_14513);
nand U15273 (N_15273,N_14745,N_14469);
nor U15274 (N_15274,N_14989,N_14976);
and U15275 (N_15275,N_14454,N_14567);
xnor U15276 (N_15276,N_14824,N_14866);
nand U15277 (N_15277,N_14656,N_14920);
or U15278 (N_15278,N_14859,N_14814);
and U15279 (N_15279,N_14995,N_14790);
nand U15280 (N_15280,N_14850,N_14623);
nand U15281 (N_15281,N_14481,N_14770);
nand U15282 (N_15282,N_14571,N_14600);
nor U15283 (N_15283,N_14550,N_14379);
and U15284 (N_15284,N_14654,N_14870);
or U15285 (N_15285,N_14418,N_14755);
xnor U15286 (N_15286,N_14961,N_14622);
nand U15287 (N_15287,N_14620,N_14987);
and U15288 (N_15288,N_14478,N_14941);
nor U15289 (N_15289,N_14896,N_14577);
or U15290 (N_15290,N_14804,N_14986);
nand U15291 (N_15291,N_14766,N_14438);
nand U15292 (N_15292,N_14683,N_14925);
xor U15293 (N_15293,N_14460,N_14657);
nor U15294 (N_15294,N_14390,N_14597);
nor U15295 (N_15295,N_14979,N_14559);
xor U15296 (N_15296,N_14442,N_14777);
and U15297 (N_15297,N_14848,N_14977);
nand U15298 (N_15298,N_14499,N_14992);
nand U15299 (N_15299,N_14624,N_14863);
xnor U15300 (N_15300,N_14608,N_14589);
or U15301 (N_15301,N_14903,N_14861);
or U15302 (N_15302,N_14520,N_14647);
nor U15303 (N_15303,N_14662,N_14411);
or U15304 (N_15304,N_14406,N_14718);
nand U15305 (N_15305,N_14455,N_14911);
xnor U15306 (N_15306,N_14886,N_14596);
or U15307 (N_15307,N_14952,N_14644);
or U15308 (N_15308,N_14983,N_14701);
or U15309 (N_15309,N_14467,N_14381);
nor U15310 (N_15310,N_14424,N_14957);
nand U15311 (N_15311,N_14414,N_14558);
or U15312 (N_15312,N_14399,N_14822);
or U15313 (N_15313,N_14988,N_14677);
or U15314 (N_15314,N_14432,N_14403);
and U15315 (N_15315,N_14849,N_14639);
or U15316 (N_15316,N_14385,N_14654);
xor U15317 (N_15317,N_14502,N_14856);
nand U15318 (N_15318,N_14831,N_14777);
or U15319 (N_15319,N_14945,N_14933);
nand U15320 (N_15320,N_14648,N_14562);
and U15321 (N_15321,N_14910,N_14474);
nand U15322 (N_15322,N_14423,N_14722);
or U15323 (N_15323,N_14726,N_14964);
and U15324 (N_15324,N_14404,N_14468);
or U15325 (N_15325,N_14901,N_14806);
or U15326 (N_15326,N_14879,N_14398);
xor U15327 (N_15327,N_14883,N_14490);
and U15328 (N_15328,N_14501,N_14968);
nand U15329 (N_15329,N_14510,N_14969);
or U15330 (N_15330,N_14616,N_14872);
nor U15331 (N_15331,N_14996,N_14789);
nor U15332 (N_15332,N_14383,N_14887);
nor U15333 (N_15333,N_14804,N_14746);
or U15334 (N_15334,N_14989,N_14830);
nand U15335 (N_15335,N_14843,N_14923);
and U15336 (N_15336,N_14997,N_14917);
and U15337 (N_15337,N_14911,N_14476);
nand U15338 (N_15338,N_14785,N_14461);
nand U15339 (N_15339,N_14764,N_14379);
and U15340 (N_15340,N_14881,N_14501);
xnor U15341 (N_15341,N_14519,N_14438);
nor U15342 (N_15342,N_14837,N_14665);
xor U15343 (N_15343,N_14952,N_14984);
and U15344 (N_15344,N_14604,N_14501);
and U15345 (N_15345,N_14591,N_14845);
nor U15346 (N_15346,N_14617,N_14388);
xnor U15347 (N_15347,N_14941,N_14643);
or U15348 (N_15348,N_14491,N_14816);
nor U15349 (N_15349,N_14482,N_14519);
and U15350 (N_15350,N_14536,N_14668);
nor U15351 (N_15351,N_14984,N_14539);
xor U15352 (N_15352,N_14794,N_14742);
nand U15353 (N_15353,N_14671,N_14555);
or U15354 (N_15354,N_14844,N_14423);
nor U15355 (N_15355,N_14749,N_14675);
or U15356 (N_15356,N_14983,N_14824);
xnor U15357 (N_15357,N_14925,N_14850);
and U15358 (N_15358,N_14540,N_14852);
or U15359 (N_15359,N_14784,N_14835);
nor U15360 (N_15360,N_14944,N_14433);
nand U15361 (N_15361,N_14506,N_14955);
and U15362 (N_15362,N_14941,N_14437);
xnor U15363 (N_15363,N_14775,N_14987);
and U15364 (N_15364,N_14575,N_14793);
nand U15365 (N_15365,N_14851,N_14578);
xnor U15366 (N_15366,N_14697,N_14860);
nand U15367 (N_15367,N_14633,N_14639);
nor U15368 (N_15368,N_14506,N_14472);
or U15369 (N_15369,N_14848,N_14383);
nand U15370 (N_15370,N_14889,N_14603);
nor U15371 (N_15371,N_14528,N_14444);
nor U15372 (N_15372,N_14452,N_14883);
nand U15373 (N_15373,N_14392,N_14742);
and U15374 (N_15374,N_14922,N_14719);
nand U15375 (N_15375,N_14869,N_14490);
xnor U15376 (N_15376,N_14399,N_14742);
nor U15377 (N_15377,N_14454,N_14422);
and U15378 (N_15378,N_14966,N_14477);
or U15379 (N_15379,N_14470,N_14571);
xnor U15380 (N_15380,N_14955,N_14878);
xor U15381 (N_15381,N_14474,N_14862);
nand U15382 (N_15382,N_14772,N_14612);
xor U15383 (N_15383,N_14506,N_14820);
nor U15384 (N_15384,N_14974,N_14730);
xor U15385 (N_15385,N_14812,N_14668);
xnor U15386 (N_15386,N_14385,N_14569);
nor U15387 (N_15387,N_14532,N_14959);
and U15388 (N_15388,N_14764,N_14759);
and U15389 (N_15389,N_14513,N_14630);
nor U15390 (N_15390,N_14616,N_14779);
xnor U15391 (N_15391,N_14887,N_14664);
xnor U15392 (N_15392,N_14644,N_14422);
nand U15393 (N_15393,N_14836,N_14400);
nor U15394 (N_15394,N_14596,N_14923);
and U15395 (N_15395,N_14931,N_14766);
xor U15396 (N_15396,N_14982,N_14517);
and U15397 (N_15397,N_14562,N_14630);
or U15398 (N_15398,N_14848,N_14481);
or U15399 (N_15399,N_14650,N_14981);
and U15400 (N_15400,N_14918,N_14810);
or U15401 (N_15401,N_14550,N_14678);
nand U15402 (N_15402,N_14938,N_14929);
or U15403 (N_15403,N_14696,N_14950);
and U15404 (N_15404,N_14692,N_14980);
nand U15405 (N_15405,N_14574,N_14389);
nand U15406 (N_15406,N_14613,N_14887);
xor U15407 (N_15407,N_14549,N_14642);
nor U15408 (N_15408,N_14733,N_14830);
or U15409 (N_15409,N_14692,N_14596);
or U15410 (N_15410,N_14587,N_14782);
nor U15411 (N_15411,N_14618,N_14383);
xnor U15412 (N_15412,N_14791,N_14718);
nand U15413 (N_15413,N_14434,N_14823);
nor U15414 (N_15414,N_14670,N_14922);
nand U15415 (N_15415,N_14973,N_14631);
and U15416 (N_15416,N_14917,N_14505);
and U15417 (N_15417,N_14817,N_14956);
nor U15418 (N_15418,N_14915,N_14426);
nor U15419 (N_15419,N_14971,N_14573);
or U15420 (N_15420,N_14448,N_14458);
xor U15421 (N_15421,N_14920,N_14909);
or U15422 (N_15422,N_14905,N_14861);
xor U15423 (N_15423,N_14807,N_14473);
xor U15424 (N_15424,N_14778,N_14981);
or U15425 (N_15425,N_14780,N_14622);
nor U15426 (N_15426,N_14569,N_14632);
and U15427 (N_15427,N_14796,N_14448);
nor U15428 (N_15428,N_14685,N_14512);
nor U15429 (N_15429,N_14565,N_14579);
nand U15430 (N_15430,N_14508,N_14734);
xor U15431 (N_15431,N_14751,N_14770);
xor U15432 (N_15432,N_14542,N_14555);
nor U15433 (N_15433,N_14378,N_14498);
nand U15434 (N_15434,N_14683,N_14745);
nor U15435 (N_15435,N_14976,N_14739);
xnor U15436 (N_15436,N_14443,N_14991);
and U15437 (N_15437,N_14376,N_14722);
nor U15438 (N_15438,N_14828,N_14720);
or U15439 (N_15439,N_14634,N_14947);
or U15440 (N_15440,N_14988,N_14904);
xnor U15441 (N_15441,N_14597,N_14516);
and U15442 (N_15442,N_14686,N_14950);
and U15443 (N_15443,N_14881,N_14716);
nor U15444 (N_15444,N_14947,N_14829);
xor U15445 (N_15445,N_14621,N_14853);
nor U15446 (N_15446,N_14707,N_14608);
or U15447 (N_15447,N_14790,N_14864);
nand U15448 (N_15448,N_14645,N_14422);
nand U15449 (N_15449,N_14513,N_14995);
nor U15450 (N_15450,N_14719,N_14681);
nand U15451 (N_15451,N_14461,N_14559);
nor U15452 (N_15452,N_14776,N_14745);
xor U15453 (N_15453,N_14774,N_14624);
xnor U15454 (N_15454,N_14535,N_14895);
nand U15455 (N_15455,N_14533,N_14970);
nor U15456 (N_15456,N_14905,N_14567);
xnor U15457 (N_15457,N_14593,N_14471);
nor U15458 (N_15458,N_14471,N_14839);
and U15459 (N_15459,N_14543,N_14588);
nor U15460 (N_15460,N_14813,N_14991);
and U15461 (N_15461,N_14417,N_14465);
or U15462 (N_15462,N_14462,N_14385);
and U15463 (N_15463,N_14987,N_14425);
nor U15464 (N_15464,N_14452,N_14951);
nand U15465 (N_15465,N_14941,N_14809);
nor U15466 (N_15466,N_14824,N_14512);
xnor U15467 (N_15467,N_14627,N_14610);
nand U15468 (N_15468,N_14644,N_14720);
or U15469 (N_15469,N_14663,N_14623);
nor U15470 (N_15470,N_14667,N_14503);
xnor U15471 (N_15471,N_14673,N_14382);
xor U15472 (N_15472,N_14704,N_14801);
nand U15473 (N_15473,N_14838,N_14787);
xnor U15474 (N_15474,N_14426,N_14619);
and U15475 (N_15475,N_14728,N_14645);
xor U15476 (N_15476,N_14516,N_14660);
xnor U15477 (N_15477,N_14534,N_14851);
or U15478 (N_15478,N_14448,N_14765);
nand U15479 (N_15479,N_14396,N_14784);
or U15480 (N_15480,N_14752,N_14412);
or U15481 (N_15481,N_14828,N_14663);
nand U15482 (N_15482,N_14381,N_14736);
nand U15483 (N_15483,N_14642,N_14858);
nor U15484 (N_15484,N_14697,N_14985);
or U15485 (N_15485,N_14742,N_14383);
nor U15486 (N_15486,N_14545,N_14786);
nor U15487 (N_15487,N_14936,N_14639);
nand U15488 (N_15488,N_14812,N_14645);
and U15489 (N_15489,N_14708,N_14882);
or U15490 (N_15490,N_14694,N_14504);
or U15491 (N_15491,N_14482,N_14729);
or U15492 (N_15492,N_14729,N_14791);
or U15493 (N_15493,N_14973,N_14913);
nand U15494 (N_15494,N_14524,N_14847);
nand U15495 (N_15495,N_14937,N_14453);
and U15496 (N_15496,N_14817,N_14896);
nand U15497 (N_15497,N_14734,N_14640);
and U15498 (N_15498,N_14961,N_14591);
nand U15499 (N_15499,N_14941,N_14783);
nor U15500 (N_15500,N_14504,N_14890);
xor U15501 (N_15501,N_14551,N_14462);
xnor U15502 (N_15502,N_14765,N_14639);
nor U15503 (N_15503,N_14665,N_14623);
nand U15504 (N_15504,N_14845,N_14982);
nor U15505 (N_15505,N_14544,N_14609);
or U15506 (N_15506,N_14612,N_14558);
nand U15507 (N_15507,N_14806,N_14537);
and U15508 (N_15508,N_14393,N_14586);
or U15509 (N_15509,N_14758,N_14715);
nand U15510 (N_15510,N_14929,N_14829);
and U15511 (N_15511,N_14901,N_14984);
or U15512 (N_15512,N_14402,N_14580);
xor U15513 (N_15513,N_14659,N_14712);
and U15514 (N_15514,N_14697,N_14520);
nand U15515 (N_15515,N_14938,N_14759);
nand U15516 (N_15516,N_14872,N_14520);
or U15517 (N_15517,N_14610,N_14772);
or U15518 (N_15518,N_14550,N_14856);
nor U15519 (N_15519,N_14502,N_14492);
nand U15520 (N_15520,N_14639,N_14586);
and U15521 (N_15521,N_14819,N_14548);
or U15522 (N_15522,N_14985,N_14904);
nand U15523 (N_15523,N_14632,N_14855);
xor U15524 (N_15524,N_14759,N_14989);
nand U15525 (N_15525,N_14457,N_14975);
and U15526 (N_15526,N_14391,N_14778);
nand U15527 (N_15527,N_14768,N_14662);
nor U15528 (N_15528,N_14861,N_14634);
xnor U15529 (N_15529,N_14635,N_14585);
nor U15530 (N_15530,N_14960,N_14840);
xor U15531 (N_15531,N_14524,N_14702);
and U15532 (N_15532,N_14792,N_14546);
nand U15533 (N_15533,N_14556,N_14959);
nand U15534 (N_15534,N_14972,N_14900);
and U15535 (N_15535,N_14815,N_14489);
and U15536 (N_15536,N_14870,N_14572);
nand U15537 (N_15537,N_14893,N_14557);
or U15538 (N_15538,N_14631,N_14985);
nand U15539 (N_15539,N_14730,N_14556);
nand U15540 (N_15540,N_14583,N_14550);
or U15541 (N_15541,N_14971,N_14440);
xor U15542 (N_15542,N_14626,N_14845);
xnor U15543 (N_15543,N_14795,N_14675);
or U15544 (N_15544,N_14561,N_14772);
xor U15545 (N_15545,N_14660,N_14979);
or U15546 (N_15546,N_14699,N_14669);
or U15547 (N_15547,N_14394,N_14666);
xor U15548 (N_15548,N_14403,N_14610);
nand U15549 (N_15549,N_14635,N_14942);
xor U15550 (N_15550,N_14446,N_14634);
and U15551 (N_15551,N_14682,N_14595);
or U15552 (N_15552,N_14619,N_14959);
nand U15553 (N_15553,N_14801,N_14451);
nor U15554 (N_15554,N_14829,N_14533);
nor U15555 (N_15555,N_14713,N_14450);
nand U15556 (N_15556,N_14737,N_14697);
or U15557 (N_15557,N_14872,N_14783);
and U15558 (N_15558,N_14575,N_14842);
and U15559 (N_15559,N_14994,N_14392);
and U15560 (N_15560,N_14546,N_14629);
and U15561 (N_15561,N_14612,N_14834);
xor U15562 (N_15562,N_14392,N_14685);
nand U15563 (N_15563,N_14649,N_14654);
and U15564 (N_15564,N_14997,N_14613);
nand U15565 (N_15565,N_14705,N_14559);
and U15566 (N_15566,N_14825,N_14831);
and U15567 (N_15567,N_14818,N_14609);
nand U15568 (N_15568,N_14593,N_14405);
or U15569 (N_15569,N_14712,N_14889);
xor U15570 (N_15570,N_14512,N_14667);
nand U15571 (N_15571,N_14968,N_14627);
or U15572 (N_15572,N_14896,N_14481);
nor U15573 (N_15573,N_14924,N_14703);
xnor U15574 (N_15574,N_14435,N_14451);
nor U15575 (N_15575,N_14702,N_14999);
and U15576 (N_15576,N_14491,N_14679);
xor U15577 (N_15577,N_14919,N_14773);
or U15578 (N_15578,N_14933,N_14655);
nand U15579 (N_15579,N_14999,N_14692);
xor U15580 (N_15580,N_14543,N_14428);
or U15581 (N_15581,N_14633,N_14402);
nor U15582 (N_15582,N_14415,N_14390);
or U15583 (N_15583,N_14797,N_14422);
xor U15584 (N_15584,N_14679,N_14956);
nand U15585 (N_15585,N_14871,N_14794);
nor U15586 (N_15586,N_14803,N_14637);
and U15587 (N_15587,N_14781,N_14600);
xnor U15588 (N_15588,N_14532,N_14808);
or U15589 (N_15589,N_14983,N_14692);
nand U15590 (N_15590,N_14907,N_14749);
nor U15591 (N_15591,N_14933,N_14457);
or U15592 (N_15592,N_14937,N_14396);
xor U15593 (N_15593,N_14624,N_14830);
nor U15594 (N_15594,N_14554,N_14827);
nor U15595 (N_15595,N_14937,N_14624);
nor U15596 (N_15596,N_14882,N_14700);
xor U15597 (N_15597,N_14478,N_14570);
nor U15598 (N_15598,N_14417,N_14672);
or U15599 (N_15599,N_14499,N_14732);
nand U15600 (N_15600,N_14534,N_14773);
nor U15601 (N_15601,N_14842,N_14553);
and U15602 (N_15602,N_14747,N_14992);
or U15603 (N_15603,N_14568,N_14664);
xor U15604 (N_15604,N_14500,N_14456);
and U15605 (N_15605,N_14649,N_14462);
xnor U15606 (N_15606,N_14877,N_14666);
xnor U15607 (N_15607,N_14497,N_14754);
and U15608 (N_15608,N_14771,N_14757);
xor U15609 (N_15609,N_14682,N_14503);
nor U15610 (N_15610,N_14485,N_14683);
xor U15611 (N_15611,N_14465,N_14404);
nand U15612 (N_15612,N_14632,N_14553);
xor U15613 (N_15613,N_14828,N_14943);
nor U15614 (N_15614,N_14947,N_14946);
and U15615 (N_15615,N_14404,N_14687);
nor U15616 (N_15616,N_14836,N_14870);
and U15617 (N_15617,N_14669,N_14694);
xnor U15618 (N_15618,N_14448,N_14473);
xnor U15619 (N_15619,N_14676,N_14565);
nor U15620 (N_15620,N_14525,N_14994);
and U15621 (N_15621,N_14541,N_14490);
xor U15622 (N_15622,N_14442,N_14917);
xnor U15623 (N_15623,N_14928,N_14513);
or U15624 (N_15624,N_14667,N_14945);
or U15625 (N_15625,N_15606,N_15205);
nand U15626 (N_15626,N_15623,N_15446);
nor U15627 (N_15627,N_15176,N_15448);
xor U15628 (N_15628,N_15159,N_15400);
nand U15629 (N_15629,N_15452,N_15476);
xnor U15630 (N_15630,N_15390,N_15428);
xnor U15631 (N_15631,N_15086,N_15032);
nand U15632 (N_15632,N_15076,N_15341);
nor U15633 (N_15633,N_15152,N_15099);
xnor U15634 (N_15634,N_15318,N_15153);
nor U15635 (N_15635,N_15046,N_15060);
nor U15636 (N_15636,N_15305,N_15059);
nor U15637 (N_15637,N_15325,N_15409);
nand U15638 (N_15638,N_15352,N_15173);
and U15639 (N_15639,N_15149,N_15609);
nor U15640 (N_15640,N_15396,N_15431);
nor U15641 (N_15641,N_15168,N_15054);
nand U15642 (N_15642,N_15199,N_15284);
or U15643 (N_15643,N_15276,N_15299);
nand U15644 (N_15644,N_15279,N_15272);
and U15645 (N_15645,N_15610,N_15415);
nand U15646 (N_15646,N_15391,N_15235);
or U15647 (N_15647,N_15438,N_15355);
xnor U15648 (N_15648,N_15566,N_15483);
or U15649 (N_15649,N_15124,N_15374);
xnor U15650 (N_15650,N_15463,N_15586);
and U15651 (N_15651,N_15209,N_15023);
or U15652 (N_15652,N_15293,N_15494);
nand U15653 (N_15653,N_15552,N_15201);
nand U15654 (N_15654,N_15560,N_15128);
and U15655 (N_15655,N_15557,N_15257);
and U15656 (N_15656,N_15114,N_15102);
nand U15657 (N_15657,N_15150,N_15321);
or U15658 (N_15658,N_15356,N_15323);
nor U15659 (N_15659,N_15090,N_15616);
nor U15660 (N_15660,N_15269,N_15345);
xor U15661 (N_15661,N_15118,N_15392);
xnor U15662 (N_15662,N_15229,N_15270);
xor U15663 (N_15663,N_15389,N_15061);
xor U15664 (N_15664,N_15237,N_15291);
or U15665 (N_15665,N_15327,N_15074);
and U15666 (N_15666,N_15250,N_15185);
xnor U15667 (N_15667,N_15144,N_15581);
xnor U15668 (N_15668,N_15600,N_15047);
or U15669 (N_15669,N_15550,N_15624);
xor U15670 (N_15670,N_15154,N_15454);
nand U15671 (N_15671,N_15614,N_15466);
xor U15672 (N_15672,N_15009,N_15363);
nor U15673 (N_15673,N_15435,N_15445);
xnor U15674 (N_15674,N_15125,N_15013);
nor U15675 (N_15675,N_15522,N_15079);
nor U15676 (N_15676,N_15018,N_15183);
nand U15677 (N_15677,N_15597,N_15535);
or U15678 (N_15678,N_15178,N_15576);
and U15679 (N_15679,N_15200,N_15069);
nand U15680 (N_15680,N_15174,N_15077);
or U15681 (N_15681,N_15575,N_15555);
xor U15682 (N_15682,N_15070,N_15603);
or U15683 (N_15683,N_15005,N_15155);
and U15684 (N_15684,N_15110,N_15437);
xnor U15685 (N_15685,N_15567,N_15207);
or U15686 (N_15686,N_15472,N_15222);
xnor U15687 (N_15687,N_15167,N_15097);
xnor U15688 (N_15688,N_15608,N_15334);
nor U15689 (N_15689,N_15596,N_15529);
or U15690 (N_15690,N_15386,N_15073);
nor U15691 (N_15691,N_15314,N_15198);
xor U15692 (N_15692,N_15584,N_15292);
xor U15693 (N_15693,N_15211,N_15516);
or U15694 (N_15694,N_15251,N_15213);
and U15695 (N_15695,N_15406,N_15460);
nand U15696 (N_15696,N_15265,N_15430);
or U15697 (N_15697,N_15326,N_15338);
nand U15698 (N_15698,N_15108,N_15471);
or U15699 (N_15699,N_15485,N_15242);
xnor U15700 (N_15700,N_15563,N_15337);
nor U15701 (N_15701,N_15620,N_15311);
nor U15702 (N_15702,N_15263,N_15619);
nor U15703 (N_15703,N_15157,N_15231);
xnor U15704 (N_15704,N_15324,N_15006);
xor U15705 (N_15705,N_15481,N_15210);
and U15706 (N_15706,N_15611,N_15387);
nor U15707 (N_15707,N_15598,N_15024);
nor U15708 (N_15708,N_15336,N_15310);
and U15709 (N_15709,N_15495,N_15513);
nor U15710 (N_15710,N_15426,N_15408);
xor U15711 (N_15711,N_15008,N_15546);
nand U15712 (N_15712,N_15177,N_15524);
nand U15713 (N_15713,N_15453,N_15595);
nor U15714 (N_15714,N_15376,N_15458);
or U15715 (N_15715,N_15421,N_15062);
nand U15716 (N_15716,N_15085,N_15056);
xnor U15717 (N_15717,N_15244,N_15568);
or U15718 (N_15718,N_15122,N_15506);
xor U15719 (N_15719,N_15562,N_15119);
nand U15720 (N_15720,N_15112,N_15302);
nor U15721 (N_15721,N_15249,N_15350);
or U15722 (N_15722,N_15289,N_15353);
and U15723 (N_15723,N_15480,N_15540);
nand U15724 (N_15724,N_15378,N_15503);
xnor U15725 (N_15725,N_15021,N_15343);
nand U15726 (N_15726,N_15105,N_15239);
or U15727 (N_15727,N_15515,N_15256);
or U15728 (N_15728,N_15601,N_15440);
and U15729 (N_15729,N_15206,N_15161);
nand U15730 (N_15730,N_15233,N_15354);
nor U15731 (N_15731,N_15156,N_15593);
nand U15732 (N_15732,N_15227,N_15084);
nand U15733 (N_15733,N_15285,N_15160);
or U15734 (N_15734,N_15377,N_15312);
and U15735 (N_15735,N_15017,N_15115);
xnor U15736 (N_15736,N_15038,N_15232);
xnor U15737 (N_15737,N_15219,N_15425);
nand U15738 (N_15738,N_15208,N_15351);
or U15739 (N_15739,N_15175,N_15297);
or U15740 (N_15740,N_15439,N_15604);
and U15741 (N_15741,N_15340,N_15322);
and U15742 (N_15742,N_15587,N_15166);
or U15743 (N_15743,N_15578,N_15298);
and U15744 (N_15744,N_15026,N_15477);
nor U15745 (N_15745,N_15103,N_15382);
or U15746 (N_15746,N_15228,N_15014);
and U15747 (N_15747,N_15190,N_15246);
or U15748 (N_15748,N_15591,N_15470);
or U15749 (N_15749,N_15308,N_15573);
or U15750 (N_15750,N_15277,N_15364);
or U15751 (N_15751,N_15525,N_15333);
nand U15752 (N_15752,N_15011,N_15545);
nand U15753 (N_15753,N_15055,N_15398);
nor U15754 (N_15754,N_15347,N_15148);
or U15755 (N_15755,N_15050,N_15262);
xor U15756 (N_15756,N_15045,N_15413);
and U15757 (N_15757,N_15004,N_15007);
or U15758 (N_15758,N_15127,N_15582);
nand U15759 (N_15759,N_15275,N_15489);
xor U15760 (N_15760,N_15320,N_15258);
and U15761 (N_15761,N_15511,N_15344);
xnor U15762 (N_15762,N_15295,N_15574);
xnor U15763 (N_15763,N_15189,N_15100);
and U15764 (N_15764,N_15532,N_15399);
xnor U15765 (N_15765,N_15375,N_15420);
or U15766 (N_15766,N_15003,N_15255);
nand U15767 (N_15767,N_15083,N_15622);
or U15768 (N_15768,N_15501,N_15362);
and U15769 (N_15769,N_15225,N_15081);
nor U15770 (N_15770,N_15106,N_15134);
nand U15771 (N_15771,N_15057,N_15309);
nor U15772 (N_15772,N_15181,N_15123);
nor U15773 (N_15773,N_15380,N_15510);
and U15774 (N_15774,N_15456,N_15131);
nor U15775 (N_15775,N_15319,N_15137);
nor U15776 (N_15776,N_15037,N_15520);
and U15777 (N_15777,N_15607,N_15163);
nand U15778 (N_15778,N_15514,N_15414);
xnor U15779 (N_15779,N_15332,N_15087);
nor U15780 (N_15780,N_15412,N_15465);
nand U15781 (N_15781,N_15182,N_15368);
or U15782 (N_15782,N_15381,N_15397);
nand U15783 (N_15783,N_15585,N_15192);
nor U15784 (N_15784,N_15195,N_15294);
or U15785 (N_15785,N_15335,N_15496);
or U15786 (N_15786,N_15290,N_15098);
nor U15787 (N_15787,N_15570,N_15360);
nor U15788 (N_15788,N_15474,N_15469);
and U15789 (N_15789,N_15526,N_15259);
nor U15790 (N_15790,N_15245,N_15618);
xor U15791 (N_15791,N_15170,N_15221);
nor U15792 (N_15792,N_15569,N_15551);
and U15793 (N_15793,N_15444,N_15104);
and U15794 (N_15794,N_15488,N_15410);
and U15795 (N_15795,N_15039,N_15533);
xnor U15796 (N_15796,N_15313,N_15530);
or U15797 (N_15797,N_15145,N_15080);
xnor U15798 (N_15798,N_15214,N_15180);
and U15799 (N_15799,N_15143,N_15253);
and U15800 (N_15800,N_15349,N_15130);
nand U15801 (N_15801,N_15405,N_15063);
and U15802 (N_15802,N_15162,N_15527);
xnor U15803 (N_15803,N_15034,N_15486);
nand U15804 (N_15804,N_15478,N_15001);
nand U15805 (N_15805,N_15531,N_15049);
nor U15806 (N_15806,N_15508,N_15191);
nor U15807 (N_15807,N_15095,N_15434);
nand U15808 (N_15808,N_15543,N_15395);
or U15809 (N_15809,N_15141,N_15539);
xor U15810 (N_15810,N_15432,N_15388);
and U15811 (N_15811,N_15184,N_15218);
or U15812 (N_15812,N_15558,N_15371);
nand U15813 (N_15813,N_15497,N_15553);
xnor U15814 (N_15814,N_15241,N_15126);
and U15815 (N_15815,N_15113,N_15212);
and U15816 (N_15816,N_15065,N_15042);
or U15817 (N_15817,N_15164,N_15462);
xor U15818 (N_15818,N_15359,N_15519);
xnor U15819 (N_15819,N_15147,N_15223);
and U15820 (N_15820,N_15120,N_15554);
nand U15821 (N_15821,N_15043,N_15082);
nor U15822 (N_15822,N_15136,N_15549);
nor U15823 (N_15823,N_15129,N_15548);
or U15824 (N_15824,N_15169,N_15407);
xor U15825 (N_15825,N_15484,N_15194);
and U15826 (N_15826,N_15101,N_15594);
and U15827 (N_15827,N_15093,N_15599);
or U15828 (N_15828,N_15538,N_15040);
and U15829 (N_15829,N_15547,N_15328);
nand U15830 (N_15830,N_15357,N_15138);
and U15831 (N_15831,N_15066,N_15367);
nor U15832 (N_15832,N_15556,N_15030);
xnor U15833 (N_15833,N_15092,N_15117);
or U15834 (N_15834,N_15304,N_15450);
nand U15835 (N_15835,N_15507,N_15579);
nor U15836 (N_15836,N_15427,N_15058);
and U15837 (N_15837,N_15204,N_15559);
or U15838 (N_15838,N_15491,N_15036);
nand U15839 (N_15839,N_15215,N_15565);
and U15840 (N_15840,N_15287,N_15536);
and U15841 (N_15841,N_15248,N_15278);
nand U15842 (N_15842,N_15505,N_15234);
and U15843 (N_15843,N_15361,N_15442);
nand U15844 (N_15844,N_15016,N_15500);
nand U15845 (N_15845,N_15067,N_15365);
nor U15846 (N_15846,N_15064,N_15089);
xor U15847 (N_15847,N_15588,N_15142);
and U15848 (N_15848,N_15369,N_15296);
nor U15849 (N_15849,N_15271,N_15401);
nand U15850 (N_15850,N_15385,N_15028);
nand U15851 (N_15851,N_15171,N_15286);
or U15852 (N_15852,N_15133,N_15331);
or U15853 (N_15853,N_15504,N_15226);
nand U15854 (N_15854,N_15188,N_15419);
nor U15855 (N_15855,N_15346,N_15424);
xnor U15856 (N_15856,N_15482,N_15025);
nand U15857 (N_15857,N_15523,N_15457);
nand U15858 (N_15858,N_15317,N_15542);
nor U15859 (N_15859,N_15202,N_15288);
and U15860 (N_15860,N_15455,N_15422);
nand U15861 (N_15861,N_15139,N_15267);
or U15862 (N_15862,N_15473,N_15281);
and U15863 (N_15863,N_15306,N_15193);
xor U15864 (N_15864,N_15197,N_15274);
nand U15865 (N_15865,N_15260,N_15094);
xnor U15866 (N_15866,N_15053,N_15052);
nor U15867 (N_15867,N_15372,N_15404);
xnor U15868 (N_15868,N_15468,N_15041);
nor U15869 (N_15869,N_15273,N_15612);
or U15870 (N_15870,N_15078,N_15528);
and U15871 (N_15871,N_15561,N_15577);
xnor U15872 (N_15872,N_15592,N_15475);
nand U15873 (N_15873,N_15339,N_15048);
and U15874 (N_15874,N_15012,N_15402);
or U15875 (N_15875,N_15348,N_15264);
xnor U15876 (N_15876,N_15534,N_15383);
and U15877 (N_15877,N_15224,N_15140);
xnor U15878 (N_15878,N_15019,N_15280);
nand U15879 (N_15879,N_15203,N_15358);
and U15880 (N_15880,N_15379,N_15151);
xnor U15881 (N_15881,N_15107,N_15394);
or U15882 (N_15882,N_15502,N_15590);
xnor U15883 (N_15883,N_15370,N_15467);
xor U15884 (N_15884,N_15315,N_15418);
nor U15885 (N_15885,N_15490,N_15564);
or U15886 (N_15886,N_15411,N_15512);
or U15887 (N_15887,N_15261,N_15051);
and U15888 (N_15888,N_15132,N_15583);
nor U15889 (N_15889,N_15499,N_15423);
xnor U15890 (N_15890,N_15429,N_15517);
or U15891 (N_15891,N_15373,N_15088);
and U15892 (N_15892,N_15072,N_15165);
nor U15893 (N_15893,N_15135,N_15236);
xor U15894 (N_15894,N_15416,N_15303);
and U15895 (N_15895,N_15498,N_15330);
or U15896 (N_15896,N_15451,N_15307);
or U15897 (N_15897,N_15493,N_15096);
or U15898 (N_15898,N_15572,N_15449);
or U15899 (N_15899,N_15254,N_15247);
nor U15900 (N_15900,N_15436,N_15033);
nor U15901 (N_15901,N_15179,N_15417);
xnor U15902 (N_15902,N_15464,N_15443);
nor U15903 (N_15903,N_15544,N_15329);
nand U15904 (N_15904,N_15252,N_15230);
or U15905 (N_15905,N_15000,N_15111);
nand U15906 (N_15906,N_15240,N_15020);
nand U15907 (N_15907,N_15518,N_15403);
nand U15908 (N_15908,N_15342,N_15187);
nand U15909 (N_15909,N_15479,N_15282);
nand U15910 (N_15910,N_15121,N_15071);
and U15911 (N_15911,N_15268,N_15172);
or U15912 (N_15912,N_15447,N_15602);
nand U15913 (N_15913,N_15509,N_15196);
and U15914 (N_15914,N_15589,N_15571);
nor U15915 (N_15915,N_15441,N_15243);
nor U15916 (N_15916,N_15116,N_15015);
nand U15917 (N_15917,N_15029,N_15091);
and U15918 (N_15918,N_15580,N_15146);
nor U15919 (N_15919,N_15301,N_15537);
nand U15920 (N_15920,N_15615,N_15487);
nand U15921 (N_15921,N_15266,N_15541);
or U15922 (N_15922,N_15002,N_15068);
and U15923 (N_15923,N_15384,N_15492);
nor U15924 (N_15924,N_15027,N_15217);
xor U15925 (N_15925,N_15283,N_15010);
nor U15926 (N_15926,N_15075,N_15216);
xnor U15927 (N_15927,N_15621,N_15461);
nor U15928 (N_15928,N_15220,N_15605);
nand U15929 (N_15929,N_15238,N_15031);
nor U15930 (N_15930,N_15035,N_15617);
xor U15931 (N_15931,N_15044,N_15521);
nand U15932 (N_15932,N_15366,N_15186);
xnor U15933 (N_15933,N_15300,N_15022);
xor U15934 (N_15934,N_15109,N_15158);
and U15935 (N_15935,N_15393,N_15433);
xnor U15936 (N_15936,N_15459,N_15613);
and U15937 (N_15937,N_15316,N_15075);
nor U15938 (N_15938,N_15160,N_15078);
nor U15939 (N_15939,N_15312,N_15116);
xnor U15940 (N_15940,N_15208,N_15353);
and U15941 (N_15941,N_15495,N_15487);
and U15942 (N_15942,N_15097,N_15409);
and U15943 (N_15943,N_15609,N_15327);
xor U15944 (N_15944,N_15339,N_15513);
or U15945 (N_15945,N_15408,N_15427);
or U15946 (N_15946,N_15417,N_15373);
nand U15947 (N_15947,N_15590,N_15474);
nand U15948 (N_15948,N_15356,N_15282);
nand U15949 (N_15949,N_15042,N_15148);
nand U15950 (N_15950,N_15321,N_15088);
nand U15951 (N_15951,N_15030,N_15066);
and U15952 (N_15952,N_15530,N_15352);
nand U15953 (N_15953,N_15330,N_15601);
and U15954 (N_15954,N_15499,N_15072);
xor U15955 (N_15955,N_15166,N_15553);
and U15956 (N_15956,N_15439,N_15066);
or U15957 (N_15957,N_15078,N_15423);
or U15958 (N_15958,N_15149,N_15304);
nand U15959 (N_15959,N_15368,N_15163);
and U15960 (N_15960,N_15156,N_15193);
nand U15961 (N_15961,N_15125,N_15461);
xor U15962 (N_15962,N_15419,N_15401);
xnor U15963 (N_15963,N_15241,N_15484);
nor U15964 (N_15964,N_15216,N_15168);
xor U15965 (N_15965,N_15616,N_15229);
nand U15966 (N_15966,N_15086,N_15073);
and U15967 (N_15967,N_15381,N_15090);
nand U15968 (N_15968,N_15608,N_15197);
and U15969 (N_15969,N_15622,N_15121);
or U15970 (N_15970,N_15366,N_15459);
or U15971 (N_15971,N_15039,N_15374);
or U15972 (N_15972,N_15170,N_15042);
nor U15973 (N_15973,N_15416,N_15260);
and U15974 (N_15974,N_15449,N_15129);
or U15975 (N_15975,N_15406,N_15216);
and U15976 (N_15976,N_15534,N_15219);
xor U15977 (N_15977,N_15068,N_15083);
nor U15978 (N_15978,N_15605,N_15415);
xnor U15979 (N_15979,N_15545,N_15379);
and U15980 (N_15980,N_15328,N_15063);
xnor U15981 (N_15981,N_15052,N_15391);
nor U15982 (N_15982,N_15435,N_15489);
or U15983 (N_15983,N_15334,N_15414);
nor U15984 (N_15984,N_15584,N_15206);
xor U15985 (N_15985,N_15597,N_15432);
nor U15986 (N_15986,N_15375,N_15028);
or U15987 (N_15987,N_15571,N_15336);
or U15988 (N_15988,N_15363,N_15044);
xor U15989 (N_15989,N_15215,N_15531);
or U15990 (N_15990,N_15008,N_15139);
xor U15991 (N_15991,N_15063,N_15388);
and U15992 (N_15992,N_15503,N_15454);
nor U15993 (N_15993,N_15600,N_15216);
xor U15994 (N_15994,N_15344,N_15115);
xnor U15995 (N_15995,N_15432,N_15053);
nand U15996 (N_15996,N_15172,N_15297);
xor U15997 (N_15997,N_15573,N_15490);
nand U15998 (N_15998,N_15225,N_15155);
nor U15999 (N_15999,N_15183,N_15126);
and U16000 (N_16000,N_15529,N_15178);
xor U16001 (N_16001,N_15567,N_15218);
or U16002 (N_16002,N_15441,N_15339);
and U16003 (N_16003,N_15016,N_15364);
or U16004 (N_16004,N_15108,N_15621);
nor U16005 (N_16005,N_15355,N_15142);
xnor U16006 (N_16006,N_15380,N_15408);
and U16007 (N_16007,N_15278,N_15351);
xor U16008 (N_16008,N_15495,N_15156);
xor U16009 (N_16009,N_15566,N_15548);
and U16010 (N_16010,N_15239,N_15481);
or U16011 (N_16011,N_15487,N_15071);
and U16012 (N_16012,N_15329,N_15618);
and U16013 (N_16013,N_15153,N_15398);
and U16014 (N_16014,N_15573,N_15207);
and U16015 (N_16015,N_15104,N_15554);
nand U16016 (N_16016,N_15073,N_15321);
nand U16017 (N_16017,N_15374,N_15016);
nand U16018 (N_16018,N_15416,N_15515);
nor U16019 (N_16019,N_15176,N_15569);
nand U16020 (N_16020,N_15505,N_15323);
and U16021 (N_16021,N_15458,N_15284);
nor U16022 (N_16022,N_15222,N_15220);
xnor U16023 (N_16023,N_15345,N_15524);
xnor U16024 (N_16024,N_15104,N_15085);
xor U16025 (N_16025,N_15592,N_15375);
and U16026 (N_16026,N_15111,N_15451);
or U16027 (N_16027,N_15151,N_15486);
xnor U16028 (N_16028,N_15322,N_15367);
and U16029 (N_16029,N_15149,N_15222);
xor U16030 (N_16030,N_15354,N_15144);
and U16031 (N_16031,N_15089,N_15498);
or U16032 (N_16032,N_15526,N_15237);
and U16033 (N_16033,N_15414,N_15611);
and U16034 (N_16034,N_15092,N_15400);
or U16035 (N_16035,N_15614,N_15526);
and U16036 (N_16036,N_15117,N_15010);
nand U16037 (N_16037,N_15175,N_15087);
or U16038 (N_16038,N_15090,N_15358);
nor U16039 (N_16039,N_15200,N_15421);
and U16040 (N_16040,N_15054,N_15101);
xor U16041 (N_16041,N_15052,N_15119);
xor U16042 (N_16042,N_15391,N_15553);
and U16043 (N_16043,N_15454,N_15510);
or U16044 (N_16044,N_15080,N_15453);
or U16045 (N_16045,N_15527,N_15243);
xor U16046 (N_16046,N_15614,N_15145);
nor U16047 (N_16047,N_15577,N_15331);
nor U16048 (N_16048,N_15377,N_15374);
nand U16049 (N_16049,N_15381,N_15405);
xor U16050 (N_16050,N_15528,N_15209);
nor U16051 (N_16051,N_15191,N_15593);
xor U16052 (N_16052,N_15137,N_15468);
nor U16053 (N_16053,N_15063,N_15059);
nor U16054 (N_16054,N_15377,N_15296);
and U16055 (N_16055,N_15499,N_15586);
xnor U16056 (N_16056,N_15273,N_15555);
and U16057 (N_16057,N_15112,N_15453);
and U16058 (N_16058,N_15369,N_15361);
xnor U16059 (N_16059,N_15610,N_15448);
or U16060 (N_16060,N_15391,N_15149);
or U16061 (N_16061,N_15527,N_15545);
and U16062 (N_16062,N_15175,N_15411);
nor U16063 (N_16063,N_15610,N_15189);
and U16064 (N_16064,N_15437,N_15253);
nand U16065 (N_16065,N_15502,N_15001);
or U16066 (N_16066,N_15525,N_15108);
xor U16067 (N_16067,N_15284,N_15427);
or U16068 (N_16068,N_15059,N_15544);
nor U16069 (N_16069,N_15438,N_15405);
nor U16070 (N_16070,N_15071,N_15529);
xor U16071 (N_16071,N_15623,N_15006);
and U16072 (N_16072,N_15368,N_15037);
nor U16073 (N_16073,N_15105,N_15082);
or U16074 (N_16074,N_15245,N_15546);
nand U16075 (N_16075,N_15440,N_15605);
and U16076 (N_16076,N_15413,N_15471);
nand U16077 (N_16077,N_15352,N_15159);
nand U16078 (N_16078,N_15356,N_15403);
or U16079 (N_16079,N_15496,N_15328);
and U16080 (N_16080,N_15157,N_15086);
nor U16081 (N_16081,N_15399,N_15490);
nand U16082 (N_16082,N_15403,N_15385);
or U16083 (N_16083,N_15530,N_15503);
and U16084 (N_16084,N_15214,N_15581);
nor U16085 (N_16085,N_15074,N_15350);
and U16086 (N_16086,N_15141,N_15579);
or U16087 (N_16087,N_15262,N_15311);
and U16088 (N_16088,N_15283,N_15500);
xnor U16089 (N_16089,N_15545,N_15329);
or U16090 (N_16090,N_15437,N_15502);
or U16091 (N_16091,N_15319,N_15222);
or U16092 (N_16092,N_15612,N_15256);
nor U16093 (N_16093,N_15564,N_15476);
and U16094 (N_16094,N_15012,N_15035);
xnor U16095 (N_16095,N_15373,N_15388);
or U16096 (N_16096,N_15262,N_15561);
nand U16097 (N_16097,N_15344,N_15196);
or U16098 (N_16098,N_15274,N_15234);
nand U16099 (N_16099,N_15079,N_15434);
and U16100 (N_16100,N_15196,N_15590);
xnor U16101 (N_16101,N_15206,N_15125);
xnor U16102 (N_16102,N_15376,N_15307);
or U16103 (N_16103,N_15388,N_15266);
nor U16104 (N_16104,N_15019,N_15163);
and U16105 (N_16105,N_15383,N_15264);
nor U16106 (N_16106,N_15147,N_15171);
xnor U16107 (N_16107,N_15535,N_15079);
xor U16108 (N_16108,N_15034,N_15610);
nor U16109 (N_16109,N_15323,N_15119);
nor U16110 (N_16110,N_15234,N_15396);
xnor U16111 (N_16111,N_15377,N_15005);
nor U16112 (N_16112,N_15065,N_15499);
nor U16113 (N_16113,N_15312,N_15464);
and U16114 (N_16114,N_15522,N_15611);
and U16115 (N_16115,N_15151,N_15457);
and U16116 (N_16116,N_15446,N_15507);
nor U16117 (N_16117,N_15472,N_15170);
xor U16118 (N_16118,N_15565,N_15399);
or U16119 (N_16119,N_15501,N_15521);
and U16120 (N_16120,N_15181,N_15435);
xor U16121 (N_16121,N_15181,N_15377);
and U16122 (N_16122,N_15179,N_15046);
or U16123 (N_16123,N_15430,N_15438);
nand U16124 (N_16124,N_15262,N_15616);
nor U16125 (N_16125,N_15214,N_15073);
nor U16126 (N_16126,N_15541,N_15305);
or U16127 (N_16127,N_15037,N_15616);
nor U16128 (N_16128,N_15059,N_15532);
xnor U16129 (N_16129,N_15335,N_15038);
nand U16130 (N_16130,N_15068,N_15237);
xor U16131 (N_16131,N_15381,N_15419);
nor U16132 (N_16132,N_15567,N_15433);
xor U16133 (N_16133,N_15391,N_15321);
nor U16134 (N_16134,N_15273,N_15301);
or U16135 (N_16135,N_15004,N_15362);
and U16136 (N_16136,N_15132,N_15221);
and U16137 (N_16137,N_15623,N_15530);
or U16138 (N_16138,N_15211,N_15479);
xor U16139 (N_16139,N_15053,N_15524);
nand U16140 (N_16140,N_15360,N_15475);
and U16141 (N_16141,N_15236,N_15583);
nor U16142 (N_16142,N_15483,N_15018);
xnor U16143 (N_16143,N_15019,N_15141);
nor U16144 (N_16144,N_15172,N_15178);
and U16145 (N_16145,N_15589,N_15303);
or U16146 (N_16146,N_15131,N_15074);
xor U16147 (N_16147,N_15237,N_15067);
or U16148 (N_16148,N_15471,N_15139);
or U16149 (N_16149,N_15105,N_15408);
nand U16150 (N_16150,N_15613,N_15592);
or U16151 (N_16151,N_15134,N_15566);
nand U16152 (N_16152,N_15576,N_15314);
or U16153 (N_16153,N_15293,N_15220);
nor U16154 (N_16154,N_15527,N_15164);
nand U16155 (N_16155,N_15042,N_15043);
nor U16156 (N_16156,N_15278,N_15510);
nor U16157 (N_16157,N_15248,N_15091);
xor U16158 (N_16158,N_15064,N_15223);
or U16159 (N_16159,N_15520,N_15605);
xor U16160 (N_16160,N_15191,N_15012);
nor U16161 (N_16161,N_15352,N_15052);
xnor U16162 (N_16162,N_15610,N_15380);
nor U16163 (N_16163,N_15572,N_15341);
and U16164 (N_16164,N_15460,N_15253);
xor U16165 (N_16165,N_15520,N_15612);
or U16166 (N_16166,N_15021,N_15234);
xor U16167 (N_16167,N_15199,N_15526);
xnor U16168 (N_16168,N_15459,N_15113);
and U16169 (N_16169,N_15014,N_15471);
nand U16170 (N_16170,N_15126,N_15589);
nor U16171 (N_16171,N_15519,N_15290);
nor U16172 (N_16172,N_15090,N_15567);
nor U16173 (N_16173,N_15014,N_15272);
xor U16174 (N_16174,N_15299,N_15569);
nand U16175 (N_16175,N_15619,N_15119);
or U16176 (N_16176,N_15135,N_15413);
xnor U16177 (N_16177,N_15302,N_15071);
and U16178 (N_16178,N_15488,N_15210);
xor U16179 (N_16179,N_15120,N_15175);
and U16180 (N_16180,N_15467,N_15416);
nand U16181 (N_16181,N_15058,N_15392);
and U16182 (N_16182,N_15588,N_15100);
xnor U16183 (N_16183,N_15225,N_15031);
nor U16184 (N_16184,N_15306,N_15578);
and U16185 (N_16185,N_15354,N_15502);
or U16186 (N_16186,N_15082,N_15469);
nor U16187 (N_16187,N_15169,N_15062);
xor U16188 (N_16188,N_15517,N_15591);
or U16189 (N_16189,N_15347,N_15262);
or U16190 (N_16190,N_15010,N_15504);
xnor U16191 (N_16191,N_15178,N_15340);
nor U16192 (N_16192,N_15545,N_15249);
nand U16193 (N_16193,N_15616,N_15233);
nor U16194 (N_16194,N_15547,N_15000);
nand U16195 (N_16195,N_15360,N_15386);
xnor U16196 (N_16196,N_15580,N_15520);
and U16197 (N_16197,N_15014,N_15291);
xor U16198 (N_16198,N_15440,N_15186);
nand U16199 (N_16199,N_15263,N_15096);
or U16200 (N_16200,N_15195,N_15461);
xnor U16201 (N_16201,N_15594,N_15436);
or U16202 (N_16202,N_15624,N_15350);
nor U16203 (N_16203,N_15433,N_15152);
nor U16204 (N_16204,N_15291,N_15243);
or U16205 (N_16205,N_15016,N_15167);
nor U16206 (N_16206,N_15281,N_15080);
nor U16207 (N_16207,N_15284,N_15492);
nand U16208 (N_16208,N_15076,N_15311);
nor U16209 (N_16209,N_15608,N_15477);
or U16210 (N_16210,N_15007,N_15615);
and U16211 (N_16211,N_15497,N_15504);
or U16212 (N_16212,N_15366,N_15097);
and U16213 (N_16213,N_15560,N_15018);
nor U16214 (N_16214,N_15542,N_15432);
or U16215 (N_16215,N_15175,N_15093);
nor U16216 (N_16216,N_15316,N_15461);
xor U16217 (N_16217,N_15463,N_15015);
and U16218 (N_16218,N_15040,N_15354);
or U16219 (N_16219,N_15478,N_15270);
and U16220 (N_16220,N_15470,N_15230);
or U16221 (N_16221,N_15046,N_15018);
or U16222 (N_16222,N_15101,N_15371);
and U16223 (N_16223,N_15385,N_15423);
nand U16224 (N_16224,N_15419,N_15504);
xor U16225 (N_16225,N_15140,N_15387);
and U16226 (N_16226,N_15211,N_15167);
nor U16227 (N_16227,N_15160,N_15046);
xnor U16228 (N_16228,N_15050,N_15621);
or U16229 (N_16229,N_15156,N_15424);
nand U16230 (N_16230,N_15210,N_15524);
nand U16231 (N_16231,N_15374,N_15436);
nand U16232 (N_16232,N_15504,N_15298);
or U16233 (N_16233,N_15217,N_15157);
nor U16234 (N_16234,N_15612,N_15333);
nor U16235 (N_16235,N_15081,N_15022);
xor U16236 (N_16236,N_15605,N_15238);
xor U16237 (N_16237,N_15415,N_15504);
xnor U16238 (N_16238,N_15554,N_15037);
or U16239 (N_16239,N_15209,N_15103);
and U16240 (N_16240,N_15147,N_15162);
xor U16241 (N_16241,N_15216,N_15568);
nor U16242 (N_16242,N_15128,N_15068);
or U16243 (N_16243,N_15516,N_15604);
and U16244 (N_16244,N_15309,N_15221);
xor U16245 (N_16245,N_15609,N_15059);
xor U16246 (N_16246,N_15586,N_15173);
xnor U16247 (N_16247,N_15443,N_15463);
nor U16248 (N_16248,N_15473,N_15445);
xnor U16249 (N_16249,N_15038,N_15316);
nand U16250 (N_16250,N_15736,N_15746);
and U16251 (N_16251,N_15639,N_15855);
nor U16252 (N_16252,N_16075,N_15885);
nand U16253 (N_16253,N_15716,N_15936);
or U16254 (N_16254,N_16236,N_15793);
nand U16255 (N_16255,N_16234,N_15672);
nor U16256 (N_16256,N_15897,N_16119);
or U16257 (N_16257,N_16194,N_15912);
and U16258 (N_16258,N_16036,N_15808);
nor U16259 (N_16259,N_15939,N_15934);
xnor U16260 (N_16260,N_16177,N_15747);
xor U16261 (N_16261,N_15698,N_16191);
nand U16262 (N_16262,N_16089,N_15911);
nand U16263 (N_16263,N_16240,N_15880);
xnor U16264 (N_16264,N_15967,N_15663);
nand U16265 (N_16265,N_15711,N_15688);
or U16266 (N_16266,N_16027,N_15728);
nor U16267 (N_16267,N_15893,N_16193);
or U16268 (N_16268,N_15948,N_16121);
nor U16269 (N_16269,N_15817,N_16144);
nand U16270 (N_16270,N_16043,N_16167);
nand U16271 (N_16271,N_15684,N_15866);
nand U16272 (N_16272,N_15838,N_15729);
xnor U16273 (N_16273,N_15992,N_15661);
nand U16274 (N_16274,N_15914,N_15771);
nand U16275 (N_16275,N_16059,N_16171);
and U16276 (N_16276,N_16047,N_16046);
or U16277 (N_16277,N_15676,N_16107);
nor U16278 (N_16278,N_16019,N_15803);
or U16279 (N_16279,N_16081,N_16136);
xnor U16280 (N_16280,N_15785,N_16198);
xnor U16281 (N_16281,N_16220,N_15642);
or U16282 (N_16282,N_16230,N_15677);
xnor U16283 (N_16283,N_16017,N_15935);
or U16284 (N_16284,N_15840,N_16025);
and U16285 (N_16285,N_15730,N_16020);
and U16286 (N_16286,N_15882,N_15789);
nor U16287 (N_16287,N_15997,N_15768);
nor U16288 (N_16288,N_15726,N_16073);
xor U16289 (N_16289,N_15990,N_16050);
and U16290 (N_16290,N_15778,N_15998);
nand U16291 (N_16291,N_15976,N_15918);
or U16292 (N_16292,N_15647,N_15950);
nor U16293 (N_16293,N_15937,N_16080);
or U16294 (N_16294,N_15909,N_16207);
nor U16295 (N_16295,N_15818,N_15791);
and U16296 (N_16296,N_16164,N_16183);
and U16297 (N_16297,N_15902,N_16238);
xor U16298 (N_16298,N_16201,N_15883);
or U16299 (N_16299,N_15843,N_16233);
nand U16300 (N_16300,N_15712,N_16231);
or U16301 (N_16301,N_15938,N_16071);
nor U16302 (N_16302,N_16060,N_15714);
nor U16303 (N_16303,N_16056,N_15851);
and U16304 (N_16304,N_15634,N_16096);
xnor U16305 (N_16305,N_15847,N_15995);
and U16306 (N_16306,N_16221,N_15784);
xor U16307 (N_16307,N_15812,N_16108);
xor U16308 (N_16308,N_15969,N_15750);
or U16309 (N_16309,N_15655,N_16052);
and U16310 (N_16310,N_15870,N_15919);
nor U16311 (N_16311,N_16094,N_16217);
nor U16312 (N_16312,N_15830,N_15899);
nor U16313 (N_16313,N_15983,N_16133);
xnor U16314 (N_16314,N_16162,N_15761);
nand U16315 (N_16315,N_15790,N_15862);
nor U16316 (N_16316,N_15942,N_15890);
nand U16317 (N_16317,N_15701,N_15766);
or U16318 (N_16318,N_16099,N_16166);
nor U16319 (N_16319,N_15668,N_16186);
and U16320 (N_16320,N_15953,N_16249);
xnor U16321 (N_16321,N_15713,N_15955);
or U16322 (N_16322,N_15806,N_15649);
xnor U16323 (N_16323,N_16208,N_15993);
xor U16324 (N_16324,N_15929,N_15987);
nand U16325 (N_16325,N_16004,N_15654);
or U16326 (N_16326,N_16148,N_16012);
xnor U16327 (N_16327,N_16216,N_16091);
or U16328 (N_16328,N_15896,N_15986);
nor U16329 (N_16329,N_15756,N_16113);
nor U16330 (N_16330,N_16082,N_16172);
nor U16331 (N_16331,N_16032,N_15844);
or U16332 (N_16332,N_15631,N_15693);
and U16333 (N_16333,N_16190,N_16045);
nor U16334 (N_16334,N_16070,N_15719);
nand U16335 (N_16335,N_16154,N_16226);
and U16336 (N_16336,N_15779,N_15679);
nand U16337 (N_16337,N_15645,N_16007);
nor U16338 (N_16338,N_16102,N_15906);
nand U16339 (N_16339,N_15651,N_15833);
nor U16340 (N_16340,N_15895,N_16041);
and U16341 (N_16341,N_16158,N_15872);
nand U16342 (N_16342,N_16222,N_16212);
nor U16343 (N_16343,N_15717,N_15968);
nand U16344 (N_16344,N_15674,N_15744);
xnor U16345 (N_16345,N_15792,N_16112);
and U16346 (N_16346,N_15845,N_15748);
nand U16347 (N_16347,N_15877,N_16124);
nand U16348 (N_16348,N_15798,N_15832);
xnor U16349 (N_16349,N_16176,N_15641);
and U16350 (N_16350,N_16127,N_15947);
and U16351 (N_16351,N_16078,N_16142);
and U16352 (N_16352,N_15894,N_15821);
or U16353 (N_16353,N_15694,N_15664);
or U16354 (N_16354,N_15762,N_15900);
nor U16355 (N_16355,N_16165,N_15898);
or U16356 (N_16356,N_16155,N_16131);
nor U16357 (N_16357,N_16084,N_15765);
or U16358 (N_16358,N_15921,N_15873);
xor U16359 (N_16359,N_16040,N_15743);
nor U16360 (N_16360,N_16140,N_15846);
or U16361 (N_16361,N_15920,N_15959);
xnor U16362 (N_16362,N_15783,N_15853);
nand U16363 (N_16363,N_16024,N_15985);
or U16364 (N_16364,N_16151,N_16197);
or U16365 (N_16365,N_15773,N_15741);
xor U16366 (N_16366,N_15974,N_15656);
and U16367 (N_16367,N_15648,N_15977);
and U16368 (N_16368,N_15800,N_15715);
or U16369 (N_16369,N_15695,N_15738);
xor U16370 (N_16370,N_15966,N_15770);
xnor U16371 (N_16371,N_15829,N_16211);
or U16372 (N_16372,N_15700,N_15644);
nand U16373 (N_16373,N_16031,N_16120);
xnor U16374 (N_16374,N_16209,N_15665);
or U16375 (N_16375,N_16072,N_16063);
nand U16376 (N_16376,N_16068,N_16141);
xnor U16377 (N_16377,N_15629,N_16175);
nand U16378 (N_16378,N_16247,N_15834);
and U16379 (N_16379,N_15903,N_16067);
nor U16380 (N_16380,N_16122,N_15856);
nand U16381 (N_16381,N_15813,N_16092);
xnor U16382 (N_16382,N_16095,N_15731);
nor U16383 (N_16383,N_15822,N_15922);
nor U16384 (N_16384,N_16015,N_16110);
nor U16385 (N_16385,N_16066,N_15901);
and U16386 (N_16386,N_16022,N_16214);
nor U16387 (N_16387,N_16196,N_16069);
xor U16388 (N_16388,N_16077,N_15923);
and U16389 (N_16389,N_16138,N_15879);
xor U16390 (N_16390,N_15857,N_15697);
or U16391 (N_16391,N_15915,N_16180);
nand U16392 (N_16392,N_15708,N_16173);
nand U16393 (N_16393,N_15742,N_15907);
nor U16394 (N_16394,N_15994,N_15940);
or U16395 (N_16395,N_16029,N_15957);
and U16396 (N_16396,N_15943,N_15703);
or U16397 (N_16397,N_15867,N_15706);
xnor U16398 (N_16398,N_15981,N_15777);
nand U16399 (N_16399,N_15763,N_16241);
nand U16400 (N_16400,N_15827,N_16129);
xor U16401 (N_16401,N_15795,N_16076);
and U16402 (N_16402,N_16009,N_15787);
and U16403 (N_16403,N_15973,N_15875);
nand U16404 (N_16404,N_16218,N_16181);
or U16405 (N_16405,N_16192,N_16023);
nor U16406 (N_16406,N_16044,N_16168);
and U16407 (N_16407,N_16106,N_15797);
nand U16408 (N_16408,N_15849,N_16039);
nor U16409 (N_16409,N_16239,N_16011);
nand U16410 (N_16410,N_16083,N_15764);
nand U16411 (N_16411,N_15687,N_16088);
nor U16412 (N_16412,N_16243,N_16195);
xor U16413 (N_16413,N_15626,N_16058);
xor U16414 (N_16414,N_15632,N_16123);
xnor U16415 (N_16415,N_15657,N_16202);
or U16416 (N_16416,N_16188,N_15886);
nor U16417 (N_16417,N_15905,N_16161);
nor U16418 (N_16418,N_15751,N_16090);
xnor U16419 (N_16419,N_15666,N_15961);
nand U16420 (N_16420,N_16206,N_15759);
nor U16421 (N_16421,N_16054,N_15908);
or U16422 (N_16422,N_15686,N_15802);
xor U16423 (N_16423,N_15889,N_15637);
and U16424 (N_16424,N_15718,N_16210);
xor U16425 (N_16425,N_16157,N_16055);
nand U16426 (N_16426,N_16185,N_16097);
or U16427 (N_16427,N_16246,N_15740);
nand U16428 (N_16428,N_15944,N_15754);
xor U16429 (N_16429,N_15868,N_15927);
xnor U16430 (N_16430,N_16104,N_16100);
nand U16431 (N_16431,N_16018,N_15678);
or U16432 (N_16432,N_15917,N_16126);
or U16433 (N_16433,N_15991,N_15627);
xnor U16434 (N_16434,N_16085,N_16049);
and U16435 (N_16435,N_15650,N_15681);
xor U16436 (N_16436,N_15788,N_15635);
nor U16437 (N_16437,N_15815,N_15824);
nand U16438 (N_16438,N_16228,N_15887);
xor U16439 (N_16439,N_15956,N_15752);
nand U16440 (N_16440,N_15774,N_16160);
or U16441 (N_16441,N_15858,N_15660);
nor U16442 (N_16442,N_15702,N_16021);
nand U16443 (N_16443,N_15996,N_15772);
nor U16444 (N_16444,N_16115,N_15720);
nand U16445 (N_16445,N_15941,N_15630);
nand U16446 (N_16446,N_15760,N_15757);
and U16447 (N_16447,N_16143,N_16135);
or U16448 (N_16448,N_16184,N_16153);
or U16449 (N_16449,N_15932,N_15837);
nand U16450 (N_16450,N_16232,N_15958);
nand U16451 (N_16451,N_16223,N_15662);
and U16452 (N_16452,N_16098,N_16169);
and U16453 (N_16453,N_15689,N_15733);
and U16454 (N_16454,N_15928,N_15675);
nand U16455 (N_16455,N_15680,N_15864);
nand U16456 (N_16456,N_15916,N_16003);
xor U16457 (N_16457,N_15850,N_15781);
or U16458 (N_16458,N_15904,N_15696);
nand U16459 (N_16459,N_16026,N_15735);
nor U16460 (N_16460,N_15739,N_16000);
nor U16461 (N_16461,N_16087,N_16150);
nand U16462 (N_16462,N_15636,N_16132);
or U16463 (N_16463,N_15972,N_15839);
or U16464 (N_16464,N_16002,N_16203);
xor U16465 (N_16465,N_15732,N_15848);
and U16466 (N_16466,N_15769,N_15705);
nand U16467 (N_16467,N_15876,N_15749);
or U16468 (N_16468,N_16146,N_16053);
nor U16469 (N_16469,N_16174,N_15874);
xor U16470 (N_16470,N_15999,N_15805);
and U16471 (N_16471,N_15737,N_15975);
nand U16472 (N_16472,N_15962,N_15925);
or U16473 (N_16473,N_15807,N_16001);
nand U16474 (N_16474,N_15669,N_15682);
nand U16475 (N_16475,N_15799,N_16204);
nor U16476 (N_16476,N_16074,N_15725);
xnor U16477 (N_16477,N_15745,N_16187);
xnor U16478 (N_16478,N_16118,N_15704);
nor U16479 (N_16479,N_16179,N_15685);
xnor U16480 (N_16480,N_15640,N_15933);
nand U16481 (N_16481,N_15721,N_15724);
xnor U16482 (N_16482,N_15653,N_15796);
nand U16483 (N_16483,N_15710,N_15691);
nand U16484 (N_16484,N_15828,N_15825);
xor U16485 (N_16485,N_15891,N_15633);
or U16486 (N_16486,N_16038,N_15804);
xor U16487 (N_16487,N_16152,N_16033);
or U16488 (N_16488,N_15810,N_15671);
xor U16489 (N_16489,N_16242,N_15811);
nor U16490 (N_16490,N_15884,N_16145);
and U16491 (N_16491,N_15988,N_16064);
xor U16492 (N_16492,N_15707,N_15926);
or U16493 (N_16493,N_15690,N_15775);
nand U16494 (N_16494,N_15964,N_16147);
xnor U16495 (N_16495,N_15692,N_16013);
xor U16496 (N_16496,N_16079,N_15816);
nor U16497 (N_16497,N_15831,N_15722);
and U16498 (N_16498,N_15869,N_15819);
nand U16499 (N_16499,N_16219,N_15951);
or U16500 (N_16500,N_15755,N_15863);
nand U16501 (N_16501,N_16215,N_15826);
or U16502 (N_16502,N_15970,N_16010);
nand U16503 (N_16503,N_15931,N_16229);
nand U16504 (N_16504,N_16093,N_15980);
xor U16505 (N_16505,N_15979,N_15652);
and U16506 (N_16506,N_16248,N_15628);
and U16507 (N_16507,N_15952,N_15861);
xor U16508 (N_16508,N_15658,N_16086);
xor U16509 (N_16509,N_15780,N_15965);
nor U16510 (N_16510,N_15982,N_15758);
xor U16511 (N_16511,N_15801,N_16109);
nand U16512 (N_16512,N_16244,N_15945);
xnor U16513 (N_16513,N_16130,N_15809);
nand U16514 (N_16514,N_15673,N_15865);
nand U16515 (N_16515,N_15727,N_16030);
nand U16516 (N_16516,N_16037,N_15625);
xnor U16517 (N_16517,N_16156,N_15989);
and U16518 (N_16518,N_15786,N_15913);
xnor U16519 (N_16519,N_15734,N_15978);
nor U16520 (N_16520,N_16235,N_15835);
and U16521 (N_16521,N_16006,N_15723);
nand U16522 (N_16522,N_15638,N_15823);
or U16523 (N_16523,N_16117,N_15946);
nor U16524 (N_16524,N_16134,N_15852);
nor U16525 (N_16525,N_16182,N_15878);
and U16526 (N_16526,N_16224,N_16178);
nor U16527 (N_16527,N_15854,N_15930);
nor U16528 (N_16528,N_16159,N_16213);
nor U16529 (N_16529,N_15860,N_15709);
or U16530 (N_16530,N_15859,N_15753);
and U16531 (N_16531,N_16103,N_15820);
and U16532 (N_16532,N_15963,N_15984);
nand U16533 (N_16533,N_16114,N_15841);
nand U16534 (N_16534,N_16227,N_16137);
nand U16535 (N_16535,N_16005,N_15646);
or U16536 (N_16536,N_15683,N_16237);
or U16537 (N_16537,N_16016,N_16163);
and U16538 (N_16538,N_16061,N_16051);
or U16539 (N_16539,N_16065,N_15871);
nand U16540 (N_16540,N_15782,N_16189);
nand U16541 (N_16541,N_16057,N_16048);
nand U16542 (N_16542,N_15842,N_15924);
nor U16543 (N_16543,N_15776,N_16028);
and U16544 (N_16544,N_16105,N_16062);
nand U16545 (N_16545,N_16116,N_16034);
nor U16546 (N_16546,N_16200,N_16125);
nand U16547 (N_16547,N_15949,N_15794);
or U16548 (N_16548,N_15643,N_15670);
or U16549 (N_16549,N_15659,N_16042);
xnor U16550 (N_16550,N_16170,N_15892);
or U16551 (N_16551,N_15881,N_16101);
nand U16552 (N_16552,N_15667,N_15699);
xor U16553 (N_16553,N_15767,N_15888);
and U16554 (N_16554,N_16139,N_16225);
nand U16555 (N_16555,N_16111,N_15836);
or U16556 (N_16556,N_16199,N_15971);
or U16557 (N_16557,N_16128,N_16205);
nor U16558 (N_16558,N_15954,N_16035);
nor U16559 (N_16559,N_15960,N_16245);
or U16560 (N_16560,N_16149,N_16008);
and U16561 (N_16561,N_15814,N_15910);
or U16562 (N_16562,N_16014,N_16035);
or U16563 (N_16563,N_15776,N_16081);
xor U16564 (N_16564,N_15780,N_15720);
nand U16565 (N_16565,N_16208,N_15996);
nor U16566 (N_16566,N_16044,N_15738);
and U16567 (N_16567,N_16106,N_15801);
xnor U16568 (N_16568,N_16063,N_15673);
nand U16569 (N_16569,N_16082,N_15980);
nand U16570 (N_16570,N_15703,N_16172);
or U16571 (N_16571,N_15732,N_16193);
nor U16572 (N_16572,N_16199,N_15893);
nor U16573 (N_16573,N_16152,N_15657);
and U16574 (N_16574,N_16064,N_15807);
or U16575 (N_16575,N_16182,N_16060);
or U16576 (N_16576,N_15642,N_15627);
and U16577 (N_16577,N_15638,N_16127);
or U16578 (N_16578,N_16044,N_15628);
and U16579 (N_16579,N_15792,N_16096);
xnor U16580 (N_16580,N_15959,N_15757);
or U16581 (N_16581,N_16204,N_15835);
xnor U16582 (N_16582,N_16232,N_15759);
and U16583 (N_16583,N_16071,N_15648);
and U16584 (N_16584,N_15847,N_15770);
and U16585 (N_16585,N_16167,N_16191);
or U16586 (N_16586,N_16040,N_15641);
xor U16587 (N_16587,N_15697,N_16210);
nand U16588 (N_16588,N_15810,N_16116);
and U16589 (N_16589,N_16166,N_15711);
xnor U16590 (N_16590,N_15933,N_16087);
and U16591 (N_16591,N_16216,N_15760);
xnor U16592 (N_16592,N_16147,N_15667);
nand U16593 (N_16593,N_16019,N_15697);
or U16594 (N_16594,N_15944,N_15935);
or U16595 (N_16595,N_15658,N_16157);
nand U16596 (N_16596,N_15914,N_15706);
nor U16597 (N_16597,N_15948,N_15817);
nor U16598 (N_16598,N_15996,N_15910);
xor U16599 (N_16599,N_16048,N_15915);
nand U16600 (N_16600,N_15788,N_15662);
and U16601 (N_16601,N_15669,N_16181);
and U16602 (N_16602,N_16048,N_16239);
nand U16603 (N_16603,N_16061,N_15862);
nor U16604 (N_16604,N_16013,N_15937);
and U16605 (N_16605,N_15670,N_16068);
xnor U16606 (N_16606,N_15947,N_16099);
xor U16607 (N_16607,N_16009,N_15676);
and U16608 (N_16608,N_16245,N_15873);
nand U16609 (N_16609,N_15908,N_15829);
nand U16610 (N_16610,N_15797,N_15968);
or U16611 (N_16611,N_16031,N_16140);
nand U16612 (N_16612,N_16148,N_15991);
xnor U16613 (N_16613,N_16036,N_16102);
or U16614 (N_16614,N_15704,N_15912);
nor U16615 (N_16615,N_16023,N_16064);
nand U16616 (N_16616,N_15676,N_15645);
nand U16617 (N_16617,N_15745,N_16044);
or U16618 (N_16618,N_15736,N_16156);
xnor U16619 (N_16619,N_15871,N_15882);
nand U16620 (N_16620,N_16089,N_16163);
xnor U16621 (N_16621,N_16052,N_16077);
nand U16622 (N_16622,N_16041,N_16089);
nand U16623 (N_16623,N_15803,N_15742);
or U16624 (N_16624,N_15999,N_15772);
and U16625 (N_16625,N_15736,N_15949);
and U16626 (N_16626,N_15853,N_15838);
or U16627 (N_16627,N_16127,N_15749);
nor U16628 (N_16628,N_16015,N_15707);
xnor U16629 (N_16629,N_15942,N_15834);
and U16630 (N_16630,N_15971,N_15749);
nor U16631 (N_16631,N_15923,N_16226);
nor U16632 (N_16632,N_15931,N_15869);
and U16633 (N_16633,N_16244,N_15766);
or U16634 (N_16634,N_15697,N_16224);
and U16635 (N_16635,N_15640,N_15747);
or U16636 (N_16636,N_16217,N_16236);
and U16637 (N_16637,N_15756,N_15839);
nor U16638 (N_16638,N_15881,N_16088);
xnor U16639 (N_16639,N_15872,N_15945);
and U16640 (N_16640,N_15971,N_15647);
and U16641 (N_16641,N_16240,N_16058);
nand U16642 (N_16642,N_15975,N_16055);
or U16643 (N_16643,N_15640,N_16159);
xor U16644 (N_16644,N_15807,N_15933);
and U16645 (N_16645,N_16207,N_16008);
nand U16646 (N_16646,N_16235,N_16114);
or U16647 (N_16647,N_16068,N_15856);
xor U16648 (N_16648,N_15763,N_15710);
or U16649 (N_16649,N_16243,N_16102);
and U16650 (N_16650,N_15753,N_15943);
or U16651 (N_16651,N_15899,N_16007);
xnor U16652 (N_16652,N_15882,N_15729);
nor U16653 (N_16653,N_15642,N_16027);
or U16654 (N_16654,N_16243,N_16152);
and U16655 (N_16655,N_15677,N_15800);
nand U16656 (N_16656,N_15683,N_15631);
nor U16657 (N_16657,N_15803,N_16013);
xor U16658 (N_16658,N_16248,N_16245);
nand U16659 (N_16659,N_16211,N_16039);
nand U16660 (N_16660,N_15672,N_15643);
nor U16661 (N_16661,N_16018,N_16228);
xor U16662 (N_16662,N_16198,N_15851);
nor U16663 (N_16663,N_15811,N_15663);
and U16664 (N_16664,N_15721,N_15727);
nand U16665 (N_16665,N_15899,N_16129);
and U16666 (N_16666,N_16195,N_16082);
nor U16667 (N_16667,N_16181,N_15779);
nor U16668 (N_16668,N_15904,N_15735);
nor U16669 (N_16669,N_15839,N_16113);
and U16670 (N_16670,N_15883,N_15790);
and U16671 (N_16671,N_16070,N_15799);
nand U16672 (N_16672,N_15700,N_15879);
or U16673 (N_16673,N_15794,N_16114);
xor U16674 (N_16674,N_15703,N_15709);
or U16675 (N_16675,N_16153,N_16155);
nand U16676 (N_16676,N_15994,N_16249);
nor U16677 (N_16677,N_15904,N_15685);
and U16678 (N_16678,N_16083,N_15953);
and U16679 (N_16679,N_15847,N_16209);
nor U16680 (N_16680,N_15759,N_16143);
xnor U16681 (N_16681,N_15760,N_15625);
and U16682 (N_16682,N_16096,N_16052);
xor U16683 (N_16683,N_15747,N_16096);
nor U16684 (N_16684,N_15694,N_15978);
nand U16685 (N_16685,N_15881,N_16130);
and U16686 (N_16686,N_15930,N_16104);
and U16687 (N_16687,N_15802,N_15669);
xnor U16688 (N_16688,N_16176,N_16198);
and U16689 (N_16689,N_16200,N_16003);
nand U16690 (N_16690,N_16193,N_15724);
nand U16691 (N_16691,N_15983,N_16190);
xor U16692 (N_16692,N_16067,N_15809);
xnor U16693 (N_16693,N_15896,N_16158);
and U16694 (N_16694,N_15639,N_15940);
xor U16695 (N_16695,N_16240,N_16000);
xor U16696 (N_16696,N_15886,N_15896);
and U16697 (N_16697,N_15938,N_15822);
xnor U16698 (N_16698,N_16027,N_15675);
nor U16699 (N_16699,N_15771,N_15965);
nand U16700 (N_16700,N_16152,N_15767);
nand U16701 (N_16701,N_15652,N_16209);
xnor U16702 (N_16702,N_15805,N_15895);
and U16703 (N_16703,N_16005,N_15864);
or U16704 (N_16704,N_15745,N_15864);
xnor U16705 (N_16705,N_16011,N_15877);
or U16706 (N_16706,N_16047,N_15923);
nand U16707 (N_16707,N_15769,N_15741);
nand U16708 (N_16708,N_15840,N_15802);
nand U16709 (N_16709,N_16169,N_16086);
or U16710 (N_16710,N_16145,N_15711);
or U16711 (N_16711,N_16131,N_16169);
and U16712 (N_16712,N_15640,N_15971);
nand U16713 (N_16713,N_16148,N_15835);
nand U16714 (N_16714,N_16011,N_15774);
nor U16715 (N_16715,N_16080,N_16051);
nand U16716 (N_16716,N_15797,N_16224);
nand U16717 (N_16717,N_15885,N_15965);
and U16718 (N_16718,N_15902,N_15625);
nor U16719 (N_16719,N_15676,N_16174);
xnor U16720 (N_16720,N_16169,N_15643);
xnor U16721 (N_16721,N_15858,N_15750);
or U16722 (N_16722,N_16045,N_15690);
nor U16723 (N_16723,N_15901,N_15765);
nand U16724 (N_16724,N_16008,N_16079);
nand U16725 (N_16725,N_15953,N_15855);
or U16726 (N_16726,N_15811,N_15890);
nand U16727 (N_16727,N_15630,N_15946);
nor U16728 (N_16728,N_16012,N_16198);
or U16729 (N_16729,N_15923,N_15908);
nand U16730 (N_16730,N_15697,N_15921);
nand U16731 (N_16731,N_15781,N_16039);
nand U16732 (N_16732,N_15716,N_15907);
nand U16733 (N_16733,N_15956,N_15897);
xnor U16734 (N_16734,N_16053,N_15678);
nor U16735 (N_16735,N_16091,N_15706);
nand U16736 (N_16736,N_16152,N_16247);
xnor U16737 (N_16737,N_16198,N_16249);
and U16738 (N_16738,N_16138,N_15966);
xnor U16739 (N_16739,N_15849,N_16234);
or U16740 (N_16740,N_15866,N_16173);
and U16741 (N_16741,N_16208,N_16161);
xor U16742 (N_16742,N_15785,N_15879);
nor U16743 (N_16743,N_16151,N_16020);
or U16744 (N_16744,N_15983,N_15834);
nor U16745 (N_16745,N_15896,N_15844);
xor U16746 (N_16746,N_15874,N_16118);
or U16747 (N_16747,N_16184,N_16046);
nand U16748 (N_16748,N_15944,N_16221);
xor U16749 (N_16749,N_15799,N_15720);
and U16750 (N_16750,N_15773,N_15883);
nor U16751 (N_16751,N_16022,N_15991);
nand U16752 (N_16752,N_15895,N_15870);
nand U16753 (N_16753,N_15765,N_16123);
nor U16754 (N_16754,N_15672,N_16041);
and U16755 (N_16755,N_15805,N_16007);
nor U16756 (N_16756,N_16010,N_15861);
xnor U16757 (N_16757,N_15999,N_15881);
and U16758 (N_16758,N_15734,N_16168);
xnor U16759 (N_16759,N_15820,N_15815);
nor U16760 (N_16760,N_15762,N_16048);
nand U16761 (N_16761,N_16001,N_15636);
nor U16762 (N_16762,N_15986,N_16050);
and U16763 (N_16763,N_16104,N_16062);
or U16764 (N_16764,N_15642,N_15947);
nand U16765 (N_16765,N_16065,N_15668);
and U16766 (N_16766,N_15696,N_16034);
or U16767 (N_16767,N_16216,N_15816);
or U16768 (N_16768,N_16046,N_16073);
nor U16769 (N_16769,N_15659,N_15769);
nand U16770 (N_16770,N_15820,N_16057);
and U16771 (N_16771,N_16190,N_15651);
or U16772 (N_16772,N_16165,N_15663);
nand U16773 (N_16773,N_16235,N_15651);
xor U16774 (N_16774,N_15704,N_16071);
or U16775 (N_16775,N_15926,N_15679);
and U16776 (N_16776,N_16044,N_16191);
nand U16777 (N_16777,N_16212,N_15863);
and U16778 (N_16778,N_16081,N_15638);
xor U16779 (N_16779,N_16218,N_15736);
nor U16780 (N_16780,N_15635,N_15907);
or U16781 (N_16781,N_15993,N_15960);
xnor U16782 (N_16782,N_15980,N_15785);
or U16783 (N_16783,N_16131,N_15809);
xnor U16784 (N_16784,N_16005,N_16169);
and U16785 (N_16785,N_16164,N_15915);
xnor U16786 (N_16786,N_16125,N_16012);
nor U16787 (N_16787,N_16076,N_15692);
nand U16788 (N_16788,N_16136,N_15957);
xnor U16789 (N_16789,N_16204,N_16233);
xor U16790 (N_16790,N_16243,N_15811);
xnor U16791 (N_16791,N_16224,N_15737);
or U16792 (N_16792,N_16018,N_15957);
nand U16793 (N_16793,N_16158,N_15674);
or U16794 (N_16794,N_16144,N_16235);
and U16795 (N_16795,N_15997,N_15926);
and U16796 (N_16796,N_15807,N_15974);
nor U16797 (N_16797,N_15826,N_16236);
nor U16798 (N_16798,N_16096,N_15834);
nor U16799 (N_16799,N_16190,N_15855);
and U16800 (N_16800,N_16205,N_15965);
and U16801 (N_16801,N_15926,N_15637);
xor U16802 (N_16802,N_15742,N_15827);
nor U16803 (N_16803,N_16000,N_16181);
xor U16804 (N_16804,N_15679,N_16046);
nor U16805 (N_16805,N_15683,N_15691);
xor U16806 (N_16806,N_16176,N_15761);
or U16807 (N_16807,N_16093,N_15940);
or U16808 (N_16808,N_15937,N_16182);
or U16809 (N_16809,N_15850,N_16236);
nor U16810 (N_16810,N_15641,N_15930);
or U16811 (N_16811,N_15889,N_15683);
nor U16812 (N_16812,N_15667,N_15761);
or U16813 (N_16813,N_16074,N_15796);
xor U16814 (N_16814,N_16167,N_16203);
nor U16815 (N_16815,N_16084,N_15841);
or U16816 (N_16816,N_16150,N_16148);
and U16817 (N_16817,N_16155,N_15955);
nor U16818 (N_16818,N_15987,N_15975);
xor U16819 (N_16819,N_16107,N_15948);
nor U16820 (N_16820,N_15690,N_16097);
or U16821 (N_16821,N_15784,N_15959);
and U16822 (N_16822,N_15698,N_15682);
nor U16823 (N_16823,N_16215,N_16208);
nor U16824 (N_16824,N_15897,N_16049);
nand U16825 (N_16825,N_16203,N_16215);
xor U16826 (N_16826,N_15895,N_15834);
nor U16827 (N_16827,N_16156,N_16217);
xor U16828 (N_16828,N_16138,N_15790);
and U16829 (N_16829,N_15746,N_16235);
and U16830 (N_16830,N_15706,N_16057);
xor U16831 (N_16831,N_15628,N_16047);
nor U16832 (N_16832,N_16025,N_16124);
or U16833 (N_16833,N_16116,N_15684);
and U16834 (N_16834,N_16157,N_15668);
and U16835 (N_16835,N_15796,N_16170);
and U16836 (N_16836,N_15725,N_15807);
nand U16837 (N_16837,N_16058,N_15784);
or U16838 (N_16838,N_16034,N_16063);
or U16839 (N_16839,N_15835,N_16015);
nand U16840 (N_16840,N_15632,N_15830);
nor U16841 (N_16841,N_15685,N_15669);
nor U16842 (N_16842,N_16053,N_16159);
and U16843 (N_16843,N_16069,N_15942);
nand U16844 (N_16844,N_15990,N_16238);
xnor U16845 (N_16845,N_15679,N_15718);
nor U16846 (N_16846,N_16170,N_16048);
or U16847 (N_16847,N_15956,N_16039);
nand U16848 (N_16848,N_15886,N_15869);
nor U16849 (N_16849,N_16169,N_16110);
nand U16850 (N_16850,N_15701,N_15802);
and U16851 (N_16851,N_16064,N_15774);
xnor U16852 (N_16852,N_16225,N_16073);
or U16853 (N_16853,N_15810,N_15901);
xor U16854 (N_16854,N_15908,N_16091);
nand U16855 (N_16855,N_15818,N_15819);
or U16856 (N_16856,N_16104,N_16031);
xor U16857 (N_16857,N_15714,N_15664);
nor U16858 (N_16858,N_15914,N_16062);
nand U16859 (N_16859,N_15902,N_16093);
xor U16860 (N_16860,N_16249,N_15954);
and U16861 (N_16861,N_16081,N_16202);
and U16862 (N_16862,N_16025,N_15935);
nand U16863 (N_16863,N_16230,N_15636);
xnor U16864 (N_16864,N_15839,N_15854);
nor U16865 (N_16865,N_15737,N_16198);
or U16866 (N_16866,N_15921,N_16035);
nand U16867 (N_16867,N_16016,N_16195);
and U16868 (N_16868,N_16151,N_16048);
nand U16869 (N_16869,N_16036,N_15740);
and U16870 (N_16870,N_15998,N_16230);
xnor U16871 (N_16871,N_15691,N_15945);
xor U16872 (N_16872,N_15813,N_15900);
and U16873 (N_16873,N_15722,N_16221);
and U16874 (N_16874,N_15778,N_16201);
or U16875 (N_16875,N_16599,N_16434);
and U16876 (N_16876,N_16749,N_16631);
nand U16877 (N_16877,N_16283,N_16873);
xnor U16878 (N_16878,N_16588,N_16484);
or U16879 (N_16879,N_16784,N_16767);
or U16880 (N_16880,N_16681,N_16662);
nor U16881 (N_16881,N_16268,N_16627);
nand U16882 (N_16882,N_16794,N_16281);
or U16883 (N_16883,N_16630,N_16814);
or U16884 (N_16884,N_16423,N_16428);
or U16885 (N_16885,N_16715,N_16388);
and U16886 (N_16886,N_16723,N_16467);
and U16887 (N_16887,N_16389,N_16514);
nand U16888 (N_16888,N_16653,N_16813);
xnor U16889 (N_16889,N_16259,N_16506);
xnor U16890 (N_16890,N_16387,N_16580);
and U16891 (N_16891,N_16337,N_16610);
and U16892 (N_16892,N_16604,N_16343);
nand U16893 (N_16893,N_16673,N_16785);
xnor U16894 (N_16894,N_16545,N_16503);
or U16895 (N_16895,N_16350,N_16362);
or U16896 (N_16896,N_16755,N_16534);
and U16897 (N_16897,N_16596,N_16846);
nor U16898 (N_16898,N_16451,N_16318);
nand U16899 (N_16899,N_16776,N_16658);
or U16900 (N_16900,N_16479,N_16316);
xor U16901 (N_16901,N_16393,N_16517);
nand U16902 (N_16902,N_16802,N_16296);
and U16903 (N_16903,N_16402,N_16555);
or U16904 (N_16904,N_16450,N_16668);
or U16905 (N_16905,N_16553,N_16375);
nand U16906 (N_16906,N_16691,N_16772);
nor U16907 (N_16907,N_16633,N_16427);
and U16908 (N_16908,N_16460,N_16406);
and U16909 (N_16909,N_16314,N_16556);
nor U16910 (N_16910,N_16410,N_16733);
nor U16911 (N_16911,N_16826,N_16509);
xor U16912 (N_16912,N_16649,N_16367);
and U16913 (N_16913,N_16600,N_16525);
and U16914 (N_16914,N_16251,N_16686);
xnor U16915 (N_16915,N_16601,N_16657);
and U16916 (N_16916,N_16414,N_16605);
nor U16917 (N_16917,N_16824,N_16618);
nor U16918 (N_16918,N_16488,N_16510);
and U16919 (N_16919,N_16300,N_16677);
and U16920 (N_16920,N_16523,N_16266);
nor U16921 (N_16921,N_16522,N_16408);
nor U16922 (N_16922,N_16758,N_16313);
or U16923 (N_16923,N_16319,N_16850);
nor U16924 (N_16924,N_16789,N_16355);
nor U16925 (N_16925,N_16378,N_16843);
xor U16926 (N_16926,N_16377,N_16255);
xnor U16927 (N_16927,N_16796,N_16575);
and U16928 (N_16928,N_16663,N_16445);
nor U16929 (N_16929,N_16271,N_16409);
nand U16930 (N_16930,N_16589,N_16728);
nand U16931 (N_16931,N_16780,N_16819);
nand U16932 (N_16932,N_16822,N_16628);
nand U16933 (N_16933,N_16828,N_16487);
nor U16934 (N_16934,N_16443,N_16284);
and U16935 (N_16935,N_16262,N_16611);
nor U16936 (N_16936,N_16299,N_16512);
nor U16937 (N_16937,N_16264,N_16579);
nor U16938 (N_16938,N_16727,N_16400);
and U16939 (N_16939,N_16647,N_16521);
and U16940 (N_16940,N_16874,N_16440);
nor U16941 (N_16941,N_16404,N_16646);
xor U16942 (N_16942,N_16497,N_16261);
and U16943 (N_16943,N_16498,N_16621);
xnor U16944 (N_16944,N_16547,N_16698);
nor U16945 (N_16945,N_16357,N_16680);
and U16946 (N_16946,N_16616,N_16861);
or U16947 (N_16947,N_16608,N_16321);
nand U16948 (N_16948,N_16660,N_16379);
nand U16949 (N_16949,N_16469,N_16474);
xor U16950 (N_16950,N_16369,N_16598);
and U16951 (N_16951,N_16690,N_16650);
xor U16952 (N_16952,N_16753,N_16446);
xor U16953 (N_16953,N_16415,N_16865);
or U16954 (N_16954,N_16501,N_16396);
nor U16955 (N_16955,N_16540,N_16371);
nand U16956 (N_16956,N_16679,N_16380);
and U16957 (N_16957,N_16326,N_16320);
or U16958 (N_16958,N_16654,N_16461);
or U16959 (N_16959,N_16513,N_16490);
or U16960 (N_16960,N_16349,N_16549);
or U16961 (N_16961,N_16855,N_16322);
nand U16962 (N_16962,N_16421,N_16529);
nand U16963 (N_16963,N_16615,N_16481);
nand U16964 (N_16964,N_16693,N_16643);
xor U16965 (N_16965,N_16834,N_16459);
and U16966 (N_16966,N_16412,N_16325);
nor U16967 (N_16967,N_16527,N_16291);
nor U16968 (N_16968,N_16815,N_16516);
or U16969 (N_16969,N_16807,N_16724);
xnor U16970 (N_16970,N_16661,N_16609);
and U16971 (N_16971,N_16636,N_16825);
or U16972 (N_16972,N_16572,N_16818);
nor U16973 (N_16973,N_16416,N_16821);
nor U16974 (N_16974,N_16612,N_16842);
nand U16975 (N_16975,N_16436,N_16713);
or U16976 (N_16976,N_16413,N_16442);
nor U16977 (N_16977,N_16839,N_16801);
or U16978 (N_16978,N_16561,N_16260);
nor U16979 (N_16979,N_16703,N_16868);
and U16980 (N_16980,N_16398,N_16366);
nor U16981 (N_16981,N_16429,N_16456);
nand U16982 (N_16982,N_16606,N_16507);
or U16983 (N_16983,N_16324,N_16701);
nand U16984 (N_16984,N_16315,N_16641);
nand U16985 (N_16985,N_16613,N_16564);
or U16986 (N_16986,N_16747,N_16483);
nor U16987 (N_16987,N_16695,N_16614);
and U16988 (N_16988,N_16504,N_16417);
and U16989 (N_16989,N_16265,N_16519);
nand U16990 (N_16990,N_16769,N_16797);
nor U16991 (N_16991,N_16625,N_16629);
and U16992 (N_16992,N_16699,N_16346);
and U16993 (N_16993,N_16358,N_16392);
or U16994 (N_16994,N_16750,N_16752);
nor U16995 (N_16995,N_16515,N_16478);
nor U16996 (N_16996,N_16333,N_16538);
and U16997 (N_16997,N_16759,N_16746);
xnor U16998 (N_16998,N_16433,N_16803);
xnor U16999 (N_16999,N_16526,N_16341);
xnor U17000 (N_17000,N_16340,N_16293);
nor U17001 (N_17001,N_16448,N_16697);
xor U17002 (N_17002,N_16872,N_16773);
nand U17003 (N_17003,N_16642,N_16499);
nand U17004 (N_17004,N_16301,N_16317);
or U17005 (N_17005,N_16859,N_16401);
nand U17006 (N_17006,N_16528,N_16505);
nand U17007 (N_17007,N_16591,N_16840);
and U17008 (N_17008,N_16269,N_16275);
xnor U17009 (N_17009,N_16684,N_16458);
nor U17010 (N_17010,N_16786,N_16774);
nand U17011 (N_17011,N_16383,N_16576);
or U17012 (N_17012,N_16287,N_16637);
xor U17013 (N_17013,N_16360,N_16390);
or U17014 (N_17014,N_16544,N_16634);
xnor U17015 (N_17015,N_16732,N_16473);
xnor U17016 (N_17016,N_16430,N_16573);
xnor U17017 (N_17017,N_16672,N_16730);
nand U17018 (N_17018,N_16811,N_16832);
and U17019 (N_17019,N_16280,N_16419);
nand U17020 (N_17020,N_16585,N_16737);
nand U17021 (N_17021,N_16263,N_16667);
and U17022 (N_17022,N_16309,N_16353);
and U17023 (N_17023,N_16620,N_16258);
nor U17024 (N_17024,N_16708,N_16775);
or U17025 (N_17025,N_16711,N_16381);
or U17026 (N_17026,N_16439,N_16761);
nand U17027 (N_17027,N_16619,N_16793);
nand U17028 (N_17028,N_16756,N_16726);
xnor U17029 (N_17029,N_16531,N_16339);
and U17030 (N_17030,N_16477,N_16804);
nor U17031 (N_17031,N_16305,N_16480);
nor U17032 (N_17032,N_16565,N_16705);
nor U17033 (N_17033,N_16462,N_16838);
or U17034 (N_17034,N_16670,N_16739);
or U17035 (N_17035,N_16721,N_16472);
or U17036 (N_17036,N_16454,N_16577);
nor U17037 (N_17037,N_16568,N_16827);
xor U17038 (N_17038,N_16787,N_16762);
nand U17039 (N_17039,N_16652,N_16548);
or U17040 (N_17040,N_16716,N_16338);
nand U17041 (N_17041,N_16869,N_16745);
nor U17042 (N_17042,N_16788,N_16295);
or U17043 (N_17043,N_16252,N_16552);
nor U17044 (N_17044,N_16744,N_16465);
or U17045 (N_17045,N_16279,N_16331);
nand U17046 (N_17046,N_16536,N_16671);
nand U17047 (N_17047,N_16607,N_16345);
nand U17048 (N_17048,N_16494,N_16664);
and U17049 (N_17049,N_16623,N_16566);
and U17050 (N_17050,N_16812,N_16347);
nor U17051 (N_17051,N_16790,N_16849);
nor U17052 (N_17052,N_16656,N_16655);
nor U17053 (N_17053,N_16741,N_16841);
or U17054 (N_17054,N_16276,N_16791);
and U17055 (N_17055,N_16256,N_16282);
nand U17056 (N_17056,N_16783,N_16782);
or U17057 (N_17057,N_16645,N_16253);
and U17058 (N_17058,N_16518,N_16798);
nor U17059 (N_17059,N_16254,N_16535);
and U17060 (N_17060,N_16274,N_16809);
or U17061 (N_17061,N_16622,N_16468);
nor U17062 (N_17062,N_16332,N_16298);
nor U17063 (N_17063,N_16688,N_16725);
xnor U17064 (N_17064,N_16635,N_16453);
nand U17065 (N_17065,N_16867,N_16836);
or U17066 (N_17066,N_16289,N_16471);
or U17067 (N_17067,N_16530,N_16748);
and U17068 (N_17068,N_16718,N_16593);
nand U17069 (N_17069,N_16336,N_16738);
xnor U17070 (N_17070,N_16675,N_16297);
or U17071 (N_17071,N_16704,N_16648);
or U17072 (N_17072,N_16851,N_16560);
nor U17073 (N_17073,N_16624,N_16444);
nand U17074 (N_17074,N_16403,N_16689);
nand U17075 (N_17075,N_16397,N_16763);
nand U17076 (N_17076,N_16386,N_16592);
nor U17077 (N_17077,N_16569,N_16632);
nand U17078 (N_17078,N_16702,N_16511);
and U17079 (N_17079,N_16823,N_16356);
nor U17080 (N_17080,N_16502,N_16543);
xor U17081 (N_17081,N_16278,N_16370);
nor U17082 (N_17082,N_16581,N_16651);
or U17083 (N_17083,N_16270,N_16368);
or U17084 (N_17084,N_16476,N_16848);
and U17085 (N_17085,N_16420,N_16372);
nor U17086 (N_17086,N_16563,N_16617);
nand U17087 (N_17087,N_16640,N_16312);
and U17088 (N_17088,N_16682,N_16496);
nand U17089 (N_17089,N_16795,N_16644);
xor U17090 (N_17090,N_16700,N_16853);
or U17091 (N_17091,N_16344,N_16768);
nand U17092 (N_17092,N_16712,N_16447);
and U17093 (N_17093,N_16342,N_16734);
and U17094 (N_17094,N_16463,N_16659);
nand U17095 (N_17095,N_16754,N_16595);
and U17096 (N_17096,N_16665,N_16683);
or U17097 (N_17097,N_16714,N_16364);
and U17098 (N_17098,N_16335,N_16435);
or U17099 (N_17099,N_16495,N_16457);
nor U17100 (N_17100,N_16764,N_16272);
nand U17101 (N_17101,N_16485,N_16524);
xor U17102 (N_17102,N_16666,N_16292);
nor U17103 (N_17103,N_16597,N_16602);
and U17104 (N_17104,N_16860,N_16866);
and U17105 (N_17105,N_16710,N_16719);
or U17106 (N_17106,N_16348,N_16405);
nand U17107 (N_17107,N_16307,N_16351);
nand U17108 (N_17108,N_16707,N_16489);
xnor U17109 (N_17109,N_16399,N_16720);
xor U17110 (N_17110,N_16328,N_16582);
xnor U17111 (N_17111,N_16559,N_16845);
nor U17112 (N_17112,N_16323,N_16810);
nand U17113 (N_17113,N_16422,N_16740);
xor U17114 (N_17114,N_16831,N_16742);
xnor U17115 (N_17115,N_16692,N_16722);
or U17116 (N_17116,N_16781,N_16603);
xor U17117 (N_17117,N_16303,N_16546);
nand U17118 (N_17118,N_16709,N_16584);
nor U17119 (N_17119,N_16583,N_16407);
or U17120 (N_17120,N_16586,N_16431);
nor U17121 (N_17121,N_16578,N_16574);
xor U17122 (N_17122,N_16449,N_16854);
and U17123 (N_17123,N_16533,N_16327);
nor U17124 (N_17124,N_16441,N_16491);
nand U17125 (N_17125,N_16771,N_16777);
xor U17126 (N_17126,N_16302,N_16792);
nand U17127 (N_17127,N_16395,N_16829);
or U17128 (N_17128,N_16587,N_16466);
xor U17129 (N_17129,N_16354,N_16508);
nand U17130 (N_17130,N_16562,N_16492);
or U17131 (N_17131,N_16844,N_16374);
or U17132 (N_17132,N_16806,N_16833);
nor U17133 (N_17133,N_16816,N_16852);
nand U17134 (N_17134,N_16385,N_16557);
and U17135 (N_17135,N_16455,N_16482);
and U17136 (N_17136,N_16669,N_16594);
or U17137 (N_17137,N_16359,N_16418);
or U17138 (N_17138,N_16550,N_16365);
nor U17139 (N_17139,N_16500,N_16542);
nand U17140 (N_17140,N_16856,N_16539);
or U17141 (N_17141,N_16743,N_16330);
nor U17142 (N_17142,N_16567,N_16382);
xnor U17143 (N_17143,N_16800,N_16862);
nor U17144 (N_17144,N_16778,N_16308);
or U17145 (N_17145,N_16257,N_16765);
nand U17146 (N_17146,N_16678,N_16871);
and U17147 (N_17147,N_16639,N_16857);
or U17148 (N_17148,N_16532,N_16558);
nand U17149 (N_17149,N_16696,N_16685);
or U17150 (N_17150,N_16424,N_16570);
or U17151 (N_17151,N_16304,N_16858);
xnor U17152 (N_17152,N_16376,N_16464);
xor U17153 (N_17153,N_16250,N_16361);
xnor U17154 (N_17154,N_16306,N_16551);
xor U17155 (N_17155,N_16537,N_16805);
and U17156 (N_17156,N_16286,N_16273);
nand U17157 (N_17157,N_16486,N_16438);
nand U17158 (N_17158,N_16310,N_16432);
or U17159 (N_17159,N_16779,N_16554);
xor U17160 (N_17160,N_16373,N_16452);
and U17161 (N_17161,N_16837,N_16329);
nor U17162 (N_17162,N_16285,N_16290);
or U17163 (N_17163,N_16475,N_16817);
nand U17164 (N_17164,N_16847,N_16425);
nand U17165 (N_17165,N_16835,N_16470);
nor U17166 (N_17166,N_16735,N_16760);
and U17167 (N_17167,N_16520,N_16493);
or U17168 (N_17168,N_16751,N_16820);
xnor U17169 (N_17169,N_16736,N_16694);
or U17170 (N_17170,N_16541,N_16571);
nor U17171 (N_17171,N_16799,N_16863);
xnor U17172 (N_17172,N_16687,N_16870);
and U17173 (N_17173,N_16808,N_16267);
and U17174 (N_17174,N_16590,N_16352);
xnor U17175 (N_17175,N_16384,N_16437);
and U17176 (N_17176,N_16729,N_16294);
and U17177 (N_17177,N_16288,N_16766);
nand U17178 (N_17178,N_16394,N_16830);
nand U17179 (N_17179,N_16676,N_16770);
nor U17180 (N_17180,N_16757,N_16706);
nor U17181 (N_17181,N_16311,N_16411);
and U17182 (N_17182,N_16731,N_16864);
xor U17183 (N_17183,N_16717,N_16277);
and U17184 (N_17184,N_16363,N_16426);
xnor U17185 (N_17185,N_16638,N_16674);
nor U17186 (N_17186,N_16391,N_16334);
nor U17187 (N_17187,N_16626,N_16512);
or U17188 (N_17188,N_16425,N_16673);
or U17189 (N_17189,N_16796,N_16298);
nor U17190 (N_17190,N_16501,N_16395);
nand U17191 (N_17191,N_16286,N_16309);
xor U17192 (N_17192,N_16555,N_16582);
nor U17193 (N_17193,N_16255,N_16421);
nand U17194 (N_17194,N_16582,N_16788);
nand U17195 (N_17195,N_16821,N_16646);
or U17196 (N_17196,N_16795,N_16585);
xor U17197 (N_17197,N_16442,N_16494);
or U17198 (N_17198,N_16477,N_16844);
and U17199 (N_17199,N_16510,N_16501);
nor U17200 (N_17200,N_16808,N_16290);
or U17201 (N_17201,N_16373,N_16700);
and U17202 (N_17202,N_16826,N_16581);
and U17203 (N_17203,N_16864,N_16646);
xnor U17204 (N_17204,N_16851,N_16814);
or U17205 (N_17205,N_16829,N_16737);
xor U17206 (N_17206,N_16485,N_16390);
nand U17207 (N_17207,N_16721,N_16594);
or U17208 (N_17208,N_16800,N_16748);
xnor U17209 (N_17209,N_16764,N_16627);
nor U17210 (N_17210,N_16600,N_16287);
or U17211 (N_17211,N_16453,N_16537);
xor U17212 (N_17212,N_16466,N_16589);
and U17213 (N_17213,N_16365,N_16287);
nor U17214 (N_17214,N_16450,N_16690);
nor U17215 (N_17215,N_16702,N_16270);
nor U17216 (N_17216,N_16761,N_16719);
and U17217 (N_17217,N_16859,N_16627);
and U17218 (N_17218,N_16369,N_16568);
xor U17219 (N_17219,N_16569,N_16747);
xnor U17220 (N_17220,N_16341,N_16859);
or U17221 (N_17221,N_16256,N_16438);
or U17222 (N_17222,N_16365,N_16616);
or U17223 (N_17223,N_16846,N_16454);
nor U17224 (N_17224,N_16434,N_16797);
nand U17225 (N_17225,N_16831,N_16488);
nand U17226 (N_17226,N_16606,N_16374);
nor U17227 (N_17227,N_16517,N_16836);
nor U17228 (N_17228,N_16554,N_16811);
nor U17229 (N_17229,N_16319,N_16772);
nand U17230 (N_17230,N_16830,N_16256);
xor U17231 (N_17231,N_16489,N_16820);
nor U17232 (N_17232,N_16736,N_16770);
and U17233 (N_17233,N_16358,N_16819);
nand U17234 (N_17234,N_16723,N_16530);
xor U17235 (N_17235,N_16322,N_16281);
or U17236 (N_17236,N_16760,N_16528);
xor U17237 (N_17237,N_16384,N_16366);
and U17238 (N_17238,N_16329,N_16638);
or U17239 (N_17239,N_16351,N_16441);
and U17240 (N_17240,N_16313,N_16594);
nor U17241 (N_17241,N_16525,N_16527);
nor U17242 (N_17242,N_16516,N_16640);
xor U17243 (N_17243,N_16762,N_16343);
nand U17244 (N_17244,N_16676,N_16621);
xnor U17245 (N_17245,N_16438,N_16464);
and U17246 (N_17246,N_16845,N_16321);
or U17247 (N_17247,N_16817,N_16480);
or U17248 (N_17248,N_16746,N_16348);
nor U17249 (N_17249,N_16387,N_16428);
nand U17250 (N_17250,N_16830,N_16869);
and U17251 (N_17251,N_16618,N_16374);
or U17252 (N_17252,N_16714,N_16517);
nand U17253 (N_17253,N_16591,N_16464);
nand U17254 (N_17254,N_16610,N_16780);
and U17255 (N_17255,N_16618,N_16686);
and U17256 (N_17256,N_16376,N_16349);
and U17257 (N_17257,N_16514,N_16835);
nor U17258 (N_17258,N_16705,N_16624);
and U17259 (N_17259,N_16761,N_16303);
nor U17260 (N_17260,N_16765,N_16596);
and U17261 (N_17261,N_16387,N_16538);
nand U17262 (N_17262,N_16272,N_16527);
or U17263 (N_17263,N_16845,N_16411);
nand U17264 (N_17264,N_16555,N_16537);
or U17265 (N_17265,N_16658,N_16452);
or U17266 (N_17266,N_16643,N_16611);
or U17267 (N_17267,N_16598,N_16741);
nor U17268 (N_17268,N_16764,N_16784);
nand U17269 (N_17269,N_16613,N_16512);
or U17270 (N_17270,N_16707,N_16549);
and U17271 (N_17271,N_16800,N_16718);
nand U17272 (N_17272,N_16629,N_16801);
and U17273 (N_17273,N_16576,N_16719);
nor U17274 (N_17274,N_16650,N_16384);
or U17275 (N_17275,N_16569,N_16416);
nor U17276 (N_17276,N_16341,N_16603);
or U17277 (N_17277,N_16271,N_16551);
nand U17278 (N_17278,N_16370,N_16856);
nand U17279 (N_17279,N_16816,N_16781);
xor U17280 (N_17280,N_16304,N_16407);
nand U17281 (N_17281,N_16573,N_16782);
or U17282 (N_17282,N_16374,N_16508);
nor U17283 (N_17283,N_16650,N_16591);
nor U17284 (N_17284,N_16513,N_16407);
nand U17285 (N_17285,N_16268,N_16443);
and U17286 (N_17286,N_16709,N_16738);
and U17287 (N_17287,N_16379,N_16274);
or U17288 (N_17288,N_16493,N_16508);
nor U17289 (N_17289,N_16823,N_16521);
xor U17290 (N_17290,N_16329,N_16551);
xnor U17291 (N_17291,N_16473,N_16505);
and U17292 (N_17292,N_16819,N_16733);
nor U17293 (N_17293,N_16681,N_16838);
and U17294 (N_17294,N_16792,N_16789);
nor U17295 (N_17295,N_16709,N_16837);
nor U17296 (N_17296,N_16579,N_16856);
and U17297 (N_17297,N_16623,N_16593);
nand U17298 (N_17298,N_16288,N_16861);
and U17299 (N_17299,N_16846,N_16752);
and U17300 (N_17300,N_16691,N_16371);
or U17301 (N_17301,N_16482,N_16539);
xor U17302 (N_17302,N_16774,N_16268);
and U17303 (N_17303,N_16274,N_16671);
xnor U17304 (N_17304,N_16812,N_16838);
or U17305 (N_17305,N_16663,N_16334);
or U17306 (N_17306,N_16672,N_16615);
nor U17307 (N_17307,N_16355,N_16840);
and U17308 (N_17308,N_16585,N_16788);
xnor U17309 (N_17309,N_16356,N_16557);
nand U17310 (N_17310,N_16318,N_16361);
nor U17311 (N_17311,N_16325,N_16402);
and U17312 (N_17312,N_16352,N_16372);
nor U17313 (N_17313,N_16513,N_16744);
nand U17314 (N_17314,N_16568,N_16464);
and U17315 (N_17315,N_16674,N_16866);
nand U17316 (N_17316,N_16388,N_16421);
xor U17317 (N_17317,N_16294,N_16498);
nor U17318 (N_17318,N_16534,N_16698);
nor U17319 (N_17319,N_16581,N_16830);
nor U17320 (N_17320,N_16708,N_16723);
nand U17321 (N_17321,N_16287,N_16869);
or U17322 (N_17322,N_16355,N_16583);
xor U17323 (N_17323,N_16338,N_16706);
nor U17324 (N_17324,N_16772,N_16719);
nand U17325 (N_17325,N_16316,N_16766);
nand U17326 (N_17326,N_16790,N_16628);
nor U17327 (N_17327,N_16847,N_16295);
and U17328 (N_17328,N_16872,N_16460);
nor U17329 (N_17329,N_16760,N_16362);
nor U17330 (N_17330,N_16821,N_16596);
nor U17331 (N_17331,N_16597,N_16610);
or U17332 (N_17332,N_16556,N_16555);
xor U17333 (N_17333,N_16598,N_16847);
nor U17334 (N_17334,N_16796,N_16399);
nor U17335 (N_17335,N_16638,N_16782);
xor U17336 (N_17336,N_16846,N_16829);
nand U17337 (N_17337,N_16628,N_16455);
nor U17338 (N_17338,N_16448,N_16835);
or U17339 (N_17339,N_16714,N_16843);
or U17340 (N_17340,N_16746,N_16811);
nand U17341 (N_17341,N_16615,N_16519);
and U17342 (N_17342,N_16543,N_16815);
and U17343 (N_17343,N_16375,N_16724);
nor U17344 (N_17344,N_16800,N_16608);
or U17345 (N_17345,N_16432,N_16553);
nor U17346 (N_17346,N_16541,N_16441);
nand U17347 (N_17347,N_16831,N_16749);
nor U17348 (N_17348,N_16631,N_16332);
xnor U17349 (N_17349,N_16376,N_16814);
nand U17350 (N_17350,N_16772,N_16537);
nand U17351 (N_17351,N_16552,N_16272);
nand U17352 (N_17352,N_16455,N_16282);
or U17353 (N_17353,N_16781,N_16430);
xor U17354 (N_17354,N_16361,N_16432);
and U17355 (N_17355,N_16426,N_16534);
xor U17356 (N_17356,N_16755,N_16745);
xnor U17357 (N_17357,N_16845,N_16251);
and U17358 (N_17358,N_16417,N_16593);
xor U17359 (N_17359,N_16367,N_16863);
and U17360 (N_17360,N_16779,N_16328);
nor U17361 (N_17361,N_16818,N_16383);
nor U17362 (N_17362,N_16384,N_16542);
xor U17363 (N_17363,N_16653,N_16864);
and U17364 (N_17364,N_16492,N_16637);
xor U17365 (N_17365,N_16337,N_16474);
xnor U17366 (N_17366,N_16354,N_16832);
nor U17367 (N_17367,N_16341,N_16376);
nor U17368 (N_17368,N_16821,N_16373);
nand U17369 (N_17369,N_16800,N_16752);
or U17370 (N_17370,N_16692,N_16760);
nor U17371 (N_17371,N_16544,N_16853);
xor U17372 (N_17372,N_16452,N_16639);
nand U17373 (N_17373,N_16652,N_16363);
nor U17374 (N_17374,N_16329,N_16519);
or U17375 (N_17375,N_16699,N_16537);
xnor U17376 (N_17376,N_16779,N_16296);
nor U17377 (N_17377,N_16863,N_16818);
and U17378 (N_17378,N_16644,N_16784);
or U17379 (N_17379,N_16692,N_16482);
nand U17380 (N_17380,N_16660,N_16518);
and U17381 (N_17381,N_16492,N_16331);
nand U17382 (N_17382,N_16604,N_16613);
xor U17383 (N_17383,N_16310,N_16817);
nor U17384 (N_17384,N_16765,N_16658);
or U17385 (N_17385,N_16699,N_16424);
or U17386 (N_17386,N_16261,N_16582);
nand U17387 (N_17387,N_16827,N_16638);
and U17388 (N_17388,N_16620,N_16785);
nor U17389 (N_17389,N_16350,N_16412);
nor U17390 (N_17390,N_16589,N_16834);
or U17391 (N_17391,N_16442,N_16706);
and U17392 (N_17392,N_16484,N_16852);
nand U17393 (N_17393,N_16868,N_16845);
or U17394 (N_17394,N_16561,N_16317);
nand U17395 (N_17395,N_16257,N_16645);
and U17396 (N_17396,N_16476,N_16608);
and U17397 (N_17397,N_16363,N_16270);
and U17398 (N_17398,N_16874,N_16781);
nor U17399 (N_17399,N_16585,N_16309);
and U17400 (N_17400,N_16778,N_16257);
xnor U17401 (N_17401,N_16421,N_16675);
nor U17402 (N_17402,N_16516,N_16805);
or U17403 (N_17403,N_16471,N_16764);
nand U17404 (N_17404,N_16297,N_16499);
nand U17405 (N_17405,N_16707,N_16713);
xor U17406 (N_17406,N_16385,N_16290);
nor U17407 (N_17407,N_16282,N_16634);
nand U17408 (N_17408,N_16737,N_16806);
and U17409 (N_17409,N_16281,N_16345);
or U17410 (N_17410,N_16253,N_16481);
nor U17411 (N_17411,N_16680,N_16617);
xor U17412 (N_17412,N_16868,N_16619);
nand U17413 (N_17413,N_16557,N_16669);
nand U17414 (N_17414,N_16702,N_16577);
nor U17415 (N_17415,N_16337,N_16661);
xor U17416 (N_17416,N_16804,N_16511);
and U17417 (N_17417,N_16296,N_16311);
or U17418 (N_17418,N_16382,N_16701);
nand U17419 (N_17419,N_16426,N_16824);
xnor U17420 (N_17420,N_16840,N_16531);
xnor U17421 (N_17421,N_16461,N_16539);
xnor U17422 (N_17422,N_16463,N_16356);
and U17423 (N_17423,N_16593,N_16648);
xor U17424 (N_17424,N_16430,N_16523);
or U17425 (N_17425,N_16418,N_16862);
xnor U17426 (N_17426,N_16610,N_16613);
or U17427 (N_17427,N_16604,N_16848);
nand U17428 (N_17428,N_16539,N_16684);
or U17429 (N_17429,N_16380,N_16388);
nand U17430 (N_17430,N_16593,N_16691);
and U17431 (N_17431,N_16381,N_16610);
nand U17432 (N_17432,N_16809,N_16312);
or U17433 (N_17433,N_16798,N_16807);
xnor U17434 (N_17434,N_16745,N_16585);
nor U17435 (N_17435,N_16666,N_16865);
nor U17436 (N_17436,N_16693,N_16323);
xnor U17437 (N_17437,N_16422,N_16582);
and U17438 (N_17438,N_16444,N_16657);
xnor U17439 (N_17439,N_16553,N_16626);
xnor U17440 (N_17440,N_16573,N_16594);
nand U17441 (N_17441,N_16431,N_16424);
nor U17442 (N_17442,N_16583,N_16714);
nor U17443 (N_17443,N_16374,N_16429);
and U17444 (N_17444,N_16812,N_16544);
or U17445 (N_17445,N_16292,N_16524);
and U17446 (N_17446,N_16393,N_16342);
nor U17447 (N_17447,N_16421,N_16798);
nand U17448 (N_17448,N_16294,N_16589);
or U17449 (N_17449,N_16606,N_16713);
nand U17450 (N_17450,N_16554,N_16296);
nor U17451 (N_17451,N_16507,N_16452);
nand U17452 (N_17452,N_16525,N_16684);
and U17453 (N_17453,N_16832,N_16423);
nor U17454 (N_17454,N_16462,N_16545);
nor U17455 (N_17455,N_16684,N_16322);
and U17456 (N_17456,N_16294,N_16573);
nor U17457 (N_17457,N_16862,N_16296);
nor U17458 (N_17458,N_16323,N_16354);
nor U17459 (N_17459,N_16445,N_16316);
and U17460 (N_17460,N_16465,N_16725);
xor U17461 (N_17461,N_16816,N_16421);
nor U17462 (N_17462,N_16766,N_16614);
and U17463 (N_17463,N_16292,N_16348);
nor U17464 (N_17464,N_16268,N_16586);
nor U17465 (N_17465,N_16720,N_16830);
and U17466 (N_17466,N_16764,N_16573);
and U17467 (N_17467,N_16468,N_16740);
and U17468 (N_17468,N_16729,N_16749);
and U17469 (N_17469,N_16477,N_16850);
nand U17470 (N_17470,N_16830,N_16793);
nor U17471 (N_17471,N_16582,N_16286);
nor U17472 (N_17472,N_16854,N_16376);
nand U17473 (N_17473,N_16313,N_16451);
nand U17474 (N_17474,N_16764,N_16666);
and U17475 (N_17475,N_16625,N_16760);
or U17476 (N_17476,N_16563,N_16853);
or U17477 (N_17477,N_16832,N_16429);
xor U17478 (N_17478,N_16451,N_16752);
nor U17479 (N_17479,N_16409,N_16291);
and U17480 (N_17480,N_16324,N_16716);
and U17481 (N_17481,N_16709,N_16387);
and U17482 (N_17482,N_16531,N_16322);
xnor U17483 (N_17483,N_16620,N_16529);
nor U17484 (N_17484,N_16374,N_16271);
nor U17485 (N_17485,N_16300,N_16309);
or U17486 (N_17486,N_16669,N_16757);
nand U17487 (N_17487,N_16260,N_16415);
xor U17488 (N_17488,N_16855,N_16424);
nand U17489 (N_17489,N_16508,N_16649);
nand U17490 (N_17490,N_16494,N_16843);
and U17491 (N_17491,N_16665,N_16783);
xor U17492 (N_17492,N_16481,N_16302);
nor U17493 (N_17493,N_16460,N_16719);
and U17494 (N_17494,N_16516,N_16521);
nor U17495 (N_17495,N_16340,N_16688);
xnor U17496 (N_17496,N_16859,N_16536);
nand U17497 (N_17497,N_16452,N_16409);
nor U17498 (N_17498,N_16521,N_16373);
nand U17499 (N_17499,N_16793,N_16359);
xor U17500 (N_17500,N_17481,N_17347);
nor U17501 (N_17501,N_16973,N_17260);
xor U17502 (N_17502,N_17438,N_17114);
and U17503 (N_17503,N_17423,N_17368);
xnor U17504 (N_17504,N_17035,N_17119);
and U17505 (N_17505,N_17101,N_17098);
or U17506 (N_17506,N_17470,N_17181);
or U17507 (N_17507,N_17175,N_17443);
xor U17508 (N_17508,N_17441,N_17070);
nand U17509 (N_17509,N_16915,N_17212);
or U17510 (N_17510,N_17432,N_17128);
xor U17511 (N_17511,N_17028,N_17229);
or U17512 (N_17512,N_17308,N_17293);
nor U17513 (N_17513,N_17310,N_17233);
nor U17514 (N_17514,N_17311,N_17295);
or U17515 (N_17515,N_17485,N_17077);
or U17516 (N_17516,N_16987,N_17091);
nand U17517 (N_17517,N_17292,N_17069);
nand U17518 (N_17518,N_17173,N_17477);
or U17519 (N_17519,N_17284,N_17376);
nor U17520 (N_17520,N_17219,N_17297);
xnor U17521 (N_17521,N_17476,N_16925);
nor U17522 (N_17522,N_17375,N_17123);
nand U17523 (N_17523,N_17268,N_17457);
nand U17524 (N_17524,N_17436,N_16888);
nor U17525 (N_17525,N_17388,N_16953);
or U17526 (N_17526,N_17362,N_16956);
nand U17527 (N_17527,N_16905,N_17027);
xnor U17528 (N_17528,N_16940,N_17294);
nor U17529 (N_17529,N_17170,N_17176);
or U17530 (N_17530,N_17277,N_17187);
and U17531 (N_17531,N_17287,N_17495);
or U17532 (N_17532,N_17235,N_17163);
xor U17533 (N_17533,N_17274,N_17102);
and U17534 (N_17534,N_17052,N_17357);
xor U17535 (N_17535,N_17285,N_16913);
nor U17536 (N_17536,N_16961,N_17019);
and U17537 (N_17537,N_17304,N_17248);
xnor U17538 (N_17538,N_16957,N_16991);
and U17539 (N_17539,N_17036,N_17334);
or U17540 (N_17540,N_17026,N_17456);
and U17541 (N_17541,N_17409,N_17426);
nand U17542 (N_17542,N_17048,N_16970);
nor U17543 (N_17543,N_17254,N_17356);
xnor U17544 (N_17544,N_17029,N_17392);
or U17545 (N_17545,N_17144,N_17309);
and U17546 (N_17546,N_17373,N_17122);
or U17547 (N_17547,N_16974,N_17404);
or U17548 (N_17548,N_17059,N_17461);
and U17549 (N_17549,N_17251,N_17132);
and U17550 (N_17550,N_17116,N_17321);
or U17551 (N_17551,N_17004,N_17113);
and U17552 (N_17552,N_17330,N_17261);
and U17553 (N_17553,N_17156,N_16881);
and U17554 (N_17554,N_17191,N_17097);
xor U17555 (N_17555,N_17136,N_17068);
nand U17556 (N_17556,N_17395,N_17449);
nand U17557 (N_17557,N_17482,N_17224);
and U17558 (N_17558,N_16930,N_17088);
xor U17559 (N_17559,N_17230,N_17290);
nand U17560 (N_17560,N_17315,N_16929);
nor U17561 (N_17561,N_17110,N_16896);
and U17562 (N_17562,N_17333,N_17343);
and U17563 (N_17563,N_17275,N_17360);
nor U17564 (N_17564,N_17281,N_17008);
or U17565 (N_17565,N_17227,N_17090);
nand U17566 (N_17566,N_16943,N_17272);
and U17567 (N_17567,N_17418,N_17021);
nor U17568 (N_17568,N_17165,N_16918);
and U17569 (N_17569,N_17263,N_17468);
or U17570 (N_17570,N_17329,N_16971);
xor U17571 (N_17571,N_17312,N_17053);
nand U17572 (N_17572,N_17016,N_17013);
nand U17573 (N_17573,N_16897,N_17015);
nand U17574 (N_17574,N_16902,N_17139);
nand U17575 (N_17575,N_17168,N_17147);
or U17576 (N_17576,N_17462,N_17446);
nand U17577 (N_17577,N_17313,N_17475);
xor U17578 (N_17578,N_17345,N_16919);
nand U17579 (N_17579,N_16922,N_16995);
or U17580 (N_17580,N_16955,N_17190);
and U17581 (N_17581,N_16931,N_17497);
and U17582 (N_17582,N_17370,N_16997);
nand U17583 (N_17583,N_17141,N_17269);
nor U17584 (N_17584,N_17197,N_17403);
xnor U17585 (N_17585,N_17124,N_17369);
nor U17586 (N_17586,N_17283,N_16920);
and U17587 (N_17587,N_17332,N_17397);
xnor U17588 (N_17588,N_17352,N_17422);
and U17589 (N_17589,N_17483,N_17039);
nor U17590 (N_17590,N_17444,N_17066);
nand U17591 (N_17591,N_16948,N_16951);
nand U17592 (N_17592,N_17379,N_16972);
or U17593 (N_17593,N_16937,N_16993);
nor U17594 (N_17594,N_17428,N_17194);
and U17595 (N_17595,N_17301,N_17220);
nor U17596 (N_17596,N_17217,N_16923);
nor U17597 (N_17597,N_17009,N_16959);
and U17598 (N_17598,N_17431,N_17244);
nor U17599 (N_17599,N_16910,N_17323);
nand U17600 (N_17600,N_17253,N_17084);
xor U17601 (N_17601,N_17266,N_17276);
or U17602 (N_17602,N_17078,N_17002);
or U17603 (N_17603,N_16939,N_17377);
nand U17604 (N_17604,N_17046,N_16946);
xor U17605 (N_17605,N_17151,N_17023);
nor U17606 (N_17606,N_17458,N_17020);
nor U17607 (N_17607,N_17092,N_16983);
nor U17608 (N_17608,N_17089,N_17363);
nand U17609 (N_17609,N_17391,N_17307);
nand U17610 (N_17610,N_17240,N_17051);
nand U17611 (N_17611,N_17467,N_16932);
and U17612 (N_17612,N_17188,N_17299);
nor U17613 (N_17613,N_17282,N_17152);
and U17614 (N_17614,N_17365,N_17396);
nor U17615 (N_17615,N_17095,N_17419);
and U17616 (N_17616,N_16924,N_17206);
nor U17617 (N_17617,N_16884,N_17288);
or U17618 (N_17618,N_16942,N_17385);
nor U17619 (N_17619,N_17427,N_17160);
nand U17620 (N_17620,N_17417,N_17382);
xor U17621 (N_17621,N_17127,N_16962);
nor U17622 (N_17622,N_17082,N_16889);
nand U17623 (N_17623,N_16989,N_17350);
or U17624 (N_17624,N_17496,N_17169);
or U17625 (N_17625,N_17264,N_17390);
nor U17626 (N_17626,N_16911,N_17087);
nand U17627 (N_17627,N_17489,N_17162);
and U17628 (N_17628,N_16958,N_16945);
xor U17629 (N_17629,N_16994,N_17111);
nand U17630 (N_17630,N_16933,N_17085);
or U17631 (N_17631,N_17262,N_17246);
and U17632 (N_17632,N_17414,N_17305);
and U17633 (N_17633,N_16965,N_16944);
or U17634 (N_17634,N_17351,N_17228);
xor U17635 (N_17635,N_17234,N_17161);
nand U17636 (N_17636,N_16886,N_17171);
nand U17637 (N_17637,N_17179,N_17083);
and U17638 (N_17638,N_17259,N_17241);
nand U17639 (N_17639,N_17093,N_16921);
or U17640 (N_17640,N_16941,N_17384);
nor U17641 (N_17641,N_17204,N_17335);
or U17642 (N_17642,N_17058,N_17226);
nor U17643 (N_17643,N_16899,N_17189);
nor U17644 (N_17644,N_17231,N_17022);
and U17645 (N_17645,N_17402,N_17215);
nor U17646 (N_17646,N_17056,N_17183);
or U17647 (N_17647,N_17131,N_17112);
and U17648 (N_17648,N_17065,N_17355);
xor U17649 (N_17649,N_17353,N_17478);
and U17650 (N_17650,N_17211,N_17367);
or U17651 (N_17651,N_17216,N_16895);
nand U17652 (N_17652,N_17416,N_16934);
or U17653 (N_17653,N_17177,N_17079);
or U17654 (N_17654,N_17439,N_17317);
or U17655 (N_17655,N_17214,N_17205);
nor U17656 (N_17656,N_17000,N_17001);
or U17657 (N_17657,N_17464,N_17209);
and U17658 (N_17658,N_17080,N_16947);
nand U17659 (N_17659,N_17279,N_16908);
or U17660 (N_17660,N_17412,N_17420);
nand U17661 (N_17661,N_17401,N_16875);
nand U17662 (N_17662,N_17232,N_17225);
nand U17663 (N_17663,N_16883,N_17349);
nand U17664 (N_17664,N_16927,N_17474);
and U17665 (N_17665,N_16952,N_17106);
and U17666 (N_17666,N_17034,N_17492);
or U17667 (N_17667,N_17129,N_16882);
or U17668 (N_17668,N_17435,N_17180);
nor U17669 (N_17669,N_17440,N_17198);
nand U17670 (N_17670,N_16976,N_16954);
nor U17671 (N_17671,N_17314,N_17207);
xnor U17672 (N_17672,N_17354,N_17239);
xor U17673 (N_17673,N_17459,N_17167);
xnor U17674 (N_17674,N_17371,N_17054);
xor U17675 (N_17675,N_17045,N_17463);
and U17676 (N_17676,N_17302,N_17223);
nor U17677 (N_17677,N_17252,N_17146);
and U17678 (N_17678,N_17405,N_17201);
and U17679 (N_17679,N_16904,N_17073);
xor U17680 (N_17680,N_17149,N_17071);
nand U17681 (N_17681,N_17258,N_17319);
xnor U17682 (N_17682,N_16990,N_17452);
and U17683 (N_17683,N_17471,N_17433);
or U17684 (N_17684,N_17142,N_17324);
and U17685 (N_17685,N_17493,N_17378);
and U17686 (N_17686,N_17243,N_17108);
nor U17687 (N_17687,N_17399,N_16998);
nor U17688 (N_17688,N_16876,N_17429);
and U17689 (N_17689,N_17407,N_17256);
nor U17690 (N_17690,N_17094,N_17273);
and U17691 (N_17691,N_17327,N_17267);
or U17692 (N_17692,N_16969,N_17050);
or U17693 (N_17693,N_17242,N_17487);
and U17694 (N_17694,N_16950,N_17118);
and U17695 (N_17695,N_17460,N_17099);
nor U17696 (N_17696,N_17133,N_16936);
nor U17697 (N_17697,N_16916,N_17451);
or U17698 (N_17698,N_17140,N_17041);
nor U17699 (N_17699,N_17072,N_17364);
nand U17700 (N_17700,N_17030,N_17255);
nor U17701 (N_17701,N_16975,N_16906);
nand U17702 (N_17702,N_17040,N_17424);
or U17703 (N_17703,N_17208,N_17380);
or U17704 (N_17704,N_17096,N_16985);
and U17705 (N_17705,N_17306,N_17195);
or U17706 (N_17706,N_17130,N_17010);
nand U17707 (N_17707,N_16900,N_17331);
or U17708 (N_17708,N_17265,N_17383);
xor U17709 (N_17709,N_17421,N_17044);
nand U17710 (N_17710,N_17320,N_17011);
and U17711 (N_17711,N_16885,N_17076);
xnor U17712 (N_17712,N_16966,N_17488);
xor U17713 (N_17713,N_17017,N_17137);
nand U17714 (N_17714,N_16980,N_17042);
or U17715 (N_17715,N_17491,N_17166);
nand U17716 (N_17716,N_17164,N_17086);
nor U17717 (N_17717,N_17328,N_17105);
or U17718 (N_17718,N_17245,N_17055);
nor U17719 (N_17719,N_17291,N_17155);
xor U17720 (N_17720,N_17237,N_17326);
nor U17721 (N_17721,N_17120,N_16909);
or U17722 (N_17722,N_16935,N_17494);
and U17723 (N_17723,N_17006,N_16890);
or U17724 (N_17724,N_17143,N_17469);
xnor U17725 (N_17725,N_17145,N_16968);
or U17726 (N_17726,N_17289,N_17341);
nor U17727 (N_17727,N_17466,N_17037);
and U17728 (N_17728,N_17061,N_17174);
xor U17729 (N_17729,N_17186,N_17024);
xor U17730 (N_17730,N_17398,N_17003);
nand U17731 (N_17731,N_17430,N_17340);
and U17732 (N_17732,N_17296,N_17005);
xnor U17733 (N_17733,N_16963,N_17150);
nor U17734 (N_17734,N_17411,N_17337);
nand U17735 (N_17735,N_17012,N_16977);
or U17736 (N_17736,N_17032,N_17318);
or U17737 (N_17737,N_17450,N_17192);
or U17738 (N_17738,N_16887,N_17154);
nor U17739 (N_17739,N_17406,N_17067);
nor U17740 (N_17740,N_17257,N_17210);
xor U17741 (N_17741,N_17322,N_17081);
nand U17742 (N_17742,N_17358,N_17203);
and U17743 (N_17743,N_17338,N_17453);
xor U17744 (N_17744,N_17342,N_16893);
nor U17745 (N_17745,N_17387,N_17238);
nand U17746 (N_17746,N_16986,N_16878);
nor U17747 (N_17747,N_17300,N_17400);
or U17748 (N_17748,N_17184,N_16960);
and U17749 (N_17749,N_16892,N_17104);
nor U17750 (N_17750,N_17158,N_17107);
xnor U17751 (N_17751,N_17063,N_17316);
xor U17752 (N_17752,N_17425,N_17202);
and U17753 (N_17753,N_17064,N_16981);
and U17754 (N_17754,N_17408,N_17182);
and U17755 (N_17755,N_17007,N_17100);
nor U17756 (N_17756,N_17121,N_17125);
nand U17757 (N_17757,N_17454,N_17445);
and U17758 (N_17758,N_17303,N_17361);
nor U17759 (N_17759,N_17336,N_16949);
and U17760 (N_17760,N_16928,N_16984);
xor U17761 (N_17761,N_16891,N_17060);
nor U17762 (N_17762,N_17193,N_16996);
or U17763 (N_17763,N_17447,N_16880);
or U17764 (N_17764,N_17394,N_17014);
nor U17765 (N_17765,N_17025,N_16914);
nand U17766 (N_17766,N_17280,N_16907);
or U17767 (N_17767,N_17410,N_17172);
or U17768 (N_17768,N_17126,N_17148);
and U17769 (N_17769,N_17486,N_17134);
nand U17770 (N_17770,N_17413,N_17344);
nand U17771 (N_17771,N_17222,N_17031);
or U17772 (N_17772,N_17221,N_16894);
and U17773 (N_17773,N_17490,N_16877);
nand U17774 (N_17774,N_17359,N_17442);
xor U17775 (N_17775,N_17448,N_16926);
nor U17776 (N_17776,N_17138,N_17386);
and U17777 (N_17777,N_16898,N_17339);
and U17778 (N_17778,N_17199,N_16917);
xnor U17779 (N_17779,N_17075,N_17473);
nor U17780 (N_17780,N_16979,N_17437);
nor U17781 (N_17781,N_17218,N_17381);
xor U17782 (N_17782,N_17109,N_16988);
xnor U17783 (N_17783,N_17117,N_16978);
and U17784 (N_17784,N_17455,N_16999);
or U17785 (N_17785,N_17278,N_17062);
and U17786 (N_17786,N_17047,N_17038);
nand U17787 (N_17787,N_17346,N_17103);
nand U17788 (N_17788,N_17480,N_17374);
or U17789 (N_17789,N_16912,N_17159);
nand U17790 (N_17790,N_17196,N_17249);
and U17791 (N_17791,N_16982,N_17157);
nor U17792 (N_17792,N_17213,N_17270);
nor U17793 (N_17793,N_17153,N_17200);
and U17794 (N_17794,N_17348,N_17185);
or U17795 (N_17795,N_17178,N_17434);
nand U17796 (N_17796,N_17389,N_17415);
and U17797 (N_17797,N_17049,N_17484);
nor U17798 (N_17798,N_17250,N_17472);
nand U17799 (N_17799,N_17074,N_16967);
nor U17800 (N_17800,N_16992,N_17247);
nor U17801 (N_17801,N_17043,N_17286);
nand U17802 (N_17802,N_17372,N_17018);
nand U17803 (N_17803,N_16879,N_17298);
or U17804 (N_17804,N_17033,N_17115);
or U17805 (N_17805,N_17325,N_17479);
nand U17806 (N_17806,N_17498,N_16964);
nand U17807 (N_17807,N_17465,N_17499);
or U17808 (N_17808,N_16901,N_16938);
and U17809 (N_17809,N_16903,N_17057);
and U17810 (N_17810,N_17271,N_17393);
or U17811 (N_17811,N_17236,N_17366);
or U17812 (N_17812,N_17135,N_16968);
or U17813 (N_17813,N_17089,N_16940);
nand U17814 (N_17814,N_17140,N_17313);
nor U17815 (N_17815,N_17256,N_17010);
nand U17816 (N_17816,N_17319,N_17282);
nor U17817 (N_17817,N_17126,N_17461);
nor U17818 (N_17818,N_17490,N_16948);
or U17819 (N_17819,N_17481,N_17096);
nor U17820 (N_17820,N_17287,N_17258);
nand U17821 (N_17821,N_17251,N_16942);
or U17822 (N_17822,N_17146,N_17240);
xor U17823 (N_17823,N_17373,N_17386);
and U17824 (N_17824,N_17199,N_17353);
or U17825 (N_17825,N_17372,N_17480);
nand U17826 (N_17826,N_17406,N_16920);
xnor U17827 (N_17827,N_17407,N_17446);
nor U17828 (N_17828,N_17100,N_17498);
or U17829 (N_17829,N_17384,N_17049);
nor U17830 (N_17830,N_17101,N_17129);
xor U17831 (N_17831,N_16949,N_16994);
or U17832 (N_17832,N_17327,N_16930);
and U17833 (N_17833,N_17024,N_17187);
and U17834 (N_17834,N_16960,N_17257);
nand U17835 (N_17835,N_17124,N_17495);
and U17836 (N_17836,N_17439,N_17457);
or U17837 (N_17837,N_16934,N_17468);
nor U17838 (N_17838,N_16895,N_17370);
nor U17839 (N_17839,N_16953,N_16973);
and U17840 (N_17840,N_17359,N_17453);
nor U17841 (N_17841,N_17014,N_17107);
and U17842 (N_17842,N_17097,N_16908);
nor U17843 (N_17843,N_17363,N_17386);
or U17844 (N_17844,N_17033,N_17412);
and U17845 (N_17845,N_17174,N_17433);
nor U17846 (N_17846,N_17130,N_17111);
xor U17847 (N_17847,N_17200,N_17493);
and U17848 (N_17848,N_17291,N_16887);
and U17849 (N_17849,N_17054,N_17033);
and U17850 (N_17850,N_16922,N_17391);
and U17851 (N_17851,N_17318,N_17000);
xnor U17852 (N_17852,N_17285,N_16898);
and U17853 (N_17853,N_16895,N_17265);
and U17854 (N_17854,N_17435,N_17462);
or U17855 (N_17855,N_17040,N_17392);
or U17856 (N_17856,N_17476,N_17070);
xnor U17857 (N_17857,N_17076,N_16896);
xnor U17858 (N_17858,N_16890,N_16994);
and U17859 (N_17859,N_17294,N_16953);
nor U17860 (N_17860,N_17027,N_17408);
nand U17861 (N_17861,N_17097,N_16989);
xor U17862 (N_17862,N_17433,N_17150);
nor U17863 (N_17863,N_17140,N_17430);
nor U17864 (N_17864,N_17276,N_17218);
xnor U17865 (N_17865,N_17482,N_17398);
nand U17866 (N_17866,N_17064,N_17144);
or U17867 (N_17867,N_17230,N_17145);
and U17868 (N_17868,N_17054,N_17221);
nor U17869 (N_17869,N_17414,N_17062);
nand U17870 (N_17870,N_16940,N_17337);
or U17871 (N_17871,N_17026,N_17028);
xor U17872 (N_17872,N_17066,N_16919);
nand U17873 (N_17873,N_16908,N_17088);
nand U17874 (N_17874,N_17029,N_17224);
xor U17875 (N_17875,N_17220,N_16954);
xor U17876 (N_17876,N_17254,N_17440);
xnor U17877 (N_17877,N_17241,N_17363);
nand U17878 (N_17878,N_16905,N_17267);
and U17879 (N_17879,N_17151,N_17013);
and U17880 (N_17880,N_17201,N_17492);
and U17881 (N_17881,N_17009,N_17379);
or U17882 (N_17882,N_16998,N_17173);
nand U17883 (N_17883,N_17005,N_17127);
xnor U17884 (N_17884,N_17349,N_17396);
nand U17885 (N_17885,N_17133,N_17470);
or U17886 (N_17886,N_17008,N_17180);
or U17887 (N_17887,N_17331,N_17379);
nand U17888 (N_17888,N_17433,N_17480);
xor U17889 (N_17889,N_17034,N_17180);
and U17890 (N_17890,N_17389,N_16991);
xor U17891 (N_17891,N_17164,N_17209);
nand U17892 (N_17892,N_17328,N_17242);
or U17893 (N_17893,N_17257,N_17403);
or U17894 (N_17894,N_17187,N_17164);
and U17895 (N_17895,N_16962,N_17237);
xor U17896 (N_17896,N_17077,N_16936);
or U17897 (N_17897,N_17260,N_16960);
or U17898 (N_17898,N_16921,N_16958);
and U17899 (N_17899,N_17295,N_17091);
xnor U17900 (N_17900,N_17240,N_17346);
and U17901 (N_17901,N_17151,N_17322);
and U17902 (N_17902,N_17481,N_17287);
or U17903 (N_17903,N_16999,N_17099);
or U17904 (N_17904,N_17407,N_17395);
and U17905 (N_17905,N_17449,N_17493);
nor U17906 (N_17906,N_17036,N_17442);
xor U17907 (N_17907,N_17103,N_16977);
xnor U17908 (N_17908,N_17071,N_16957);
nand U17909 (N_17909,N_17132,N_17034);
xor U17910 (N_17910,N_17103,N_16888);
nor U17911 (N_17911,N_17146,N_17123);
and U17912 (N_17912,N_17467,N_17315);
or U17913 (N_17913,N_17412,N_17374);
xnor U17914 (N_17914,N_17001,N_17055);
nand U17915 (N_17915,N_16950,N_17314);
xnor U17916 (N_17916,N_17336,N_17333);
nor U17917 (N_17917,N_17429,N_16964);
xnor U17918 (N_17918,N_17134,N_17386);
nand U17919 (N_17919,N_17498,N_17120);
nor U17920 (N_17920,N_17300,N_17384);
and U17921 (N_17921,N_16982,N_17472);
nand U17922 (N_17922,N_17024,N_17188);
nor U17923 (N_17923,N_17253,N_16988);
and U17924 (N_17924,N_17306,N_16983);
nand U17925 (N_17925,N_17432,N_17238);
nand U17926 (N_17926,N_17429,N_17316);
xnor U17927 (N_17927,N_17125,N_17313);
and U17928 (N_17928,N_17052,N_17043);
nand U17929 (N_17929,N_17210,N_17446);
nand U17930 (N_17930,N_17350,N_16970);
and U17931 (N_17931,N_16931,N_17252);
nor U17932 (N_17932,N_17285,N_17251);
nand U17933 (N_17933,N_17146,N_16928);
nand U17934 (N_17934,N_17461,N_16928);
xnor U17935 (N_17935,N_17190,N_17455);
xor U17936 (N_17936,N_17063,N_17233);
nor U17937 (N_17937,N_17328,N_17301);
and U17938 (N_17938,N_17480,N_16995);
xor U17939 (N_17939,N_16967,N_16943);
or U17940 (N_17940,N_17405,N_16899);
xnor U17941 (N_17941,N_17388,N_17204);
nand U17942 (N_17942,N_17377,N_17215);
xnor U17943 (N_17943,N_16932,N_17010);
nor U17944 (N_17944,N_17427,N_16968);
and U17945 (N_17945,N_17240,N_17050);
nand U17946 (N_17946,N_16887,N_17060);
and U17947 (N_17947,N_17069,N_16975);
or U17948 (N_17948,N_16957,N_17427);
xnor U17949 (N_17949,N_17257,N_16991);
xnor U17950 (N_17950,N_17217,N_17052);
nand U17951 (N_17951,N_17368,N_17127);
or U17952 (N_17952,N_17361,N_17452);
nand U17953 (N_17953,N_17152,N_16988);
nor U17954 (N_17954,N_17469,N_17449);
nor U17955 (N_17955,N_17286,N_17046);
xnor U17956 (N_17956,N_17476,N_17147);
and U17957 (N_17957,N_17271,N_17281);
xnor U17958 (N_17958,N_17368,N_17410);
and U17959 (N_17959,N_16900,N_17381);
and U17960 (N_17960,N_16917,N_17001);
xor U17961 (N_17961,N_16924,N_16962);
or U17962 (N_17962,N_17195,N_17373);
xnor U17963 (N_17963,N_17106,N_17466);
nor U17964 (N_17964,N_17179,N_17259);
nor U17965 (N_17965,N_17072,N_17049);
and U17966 (N_17966,N_17187,N_16983);
xnor U17967 (N_17967,N_17150,N_17344);
and U17968 (N_17968,N_17332,N_17107);
nor U17969 (N_17969,N_17019,N_17068);
xnor U17970 (N_17970,N_17051,N_17414);
and U17971 (N_17971,N_17445,N_16991);
or U17972 (N_17972,N_17140,N_16934);
xor U17973 (N_17973,N_17239,N_17283);
nand U17974 (N_17974,N_16894,N_17324);
xnor U17975 (N_17975,N_17446,N_16883);
or U17976 (N_17976,N_17449,N_17173);
nor U17977 (N_17977,N_17060,N_17153);
or U17978 (N_17978,N_17364,N_17078);
xor U17979 (N_17979,N_17093,N_17407);
xor U17980 (N_17980,N_17170,N_17437);
or U17981 (N_17981,N_17474,N_17260);
or U17982 (N_17982,N_17354,N_17377);
nand U17983 (N_17983,N_17237,N_16976);
and U17984 (N_17984,N_17209,N_17381);
and U17985 (N_17985,N_17209,N_17450);
nand U17986 (N_17986,N_17356,N_17163);
xor U17987 (N_17987,N_17248,N_17147);
xnor U17988 (N_17988,N_17313,N_16907);
or U17989 (N_17989,N_17309,N_17055);
nor U17990 (N_17990,N_17366,N_17407);
nand U17991 (N_17991,N_17032,N_16967);
or U17992 (N_17992,N_17475,N_16891);
nand U17993 (N_17993,N_16978,N_17021);
nor U17994 (N_17994,N_17374,N_17134);
nand U17995 (N_17995,N_17423,N_16997);
or U17996 (N_17996,N_17098,N_17498);
nand U17997 (N_17997,N_17429,N_17314);
nand U17998 (N_17998,N_17266,N_17230);
nor U17999 (N_17999,N_17321,N_17495);
nand U18000 (N_18000,N_17447,N_17049);
or U18001 (N_18001,N_17372,N_16951);
xor U18002 (N_18002,N_17405,N_17203);
nand U18003 (N_18003,N_17340,N_17277);
and U18004 (N_18004,N_17440,N_17239);
or U18005 (N_18005,N_17418,N_16982);
and U18006 (N_18006,N_17235,N_17344);
or U18007 (N_18007,N_17450,N_16971);
or U18008 (N_18008,N_17041,N_16955);
and U18009 (N_18009,N_16980,N_17342);
nor U18010 (N_18010,N_17471,N_17005);
or U18011 (N_18011,N_17106,N_17450);
nor U18012 (N_18012,N_17200,N_17110);
and U18013 (N_18013,N_17463,N_16934);
nor U18014 (N_18014,N_17309,N_17419);
or U18015 (N_18015,N_17439,N_17266);
nand U18016 (N_18016,N_16982,N_17128);
or U18017 (N_18017,N_16922,N_17461);
xnor U18018 (N_18018,N_17378,N_17076);
nor U18019 (N_18019,N_17330,N_17034);
nor U18020 (N_18020,N_17331,N_17347);
nand U18021 (N_18021,N_17024,N_17234);
nor U18022 (N_18022,N_17017,N_17014);
and U18023 (N_18023,N_17179,N_17396);
nand U18024 (N_18024,N_17154,N_16944);
xor U18025 (N_18025,N_17022,N_17432);
xnor U18026 (N_18026,N_17265,N_17443);
nor U18027 (N_18027,N_17154,N_17469);
xnor U18028 (N_18028,N_17390,N_17313);
or U18029 (N_18029,N_16890,N_17228);
xnor U18030 (N_18030,N_17172,N_17080);
and U18031 (N_18031,N_17478,N_17177);
or U18032 (N_18032,N_17210,N_17269);
nor U18033 (N_18033,N_17091,N_16938);
xor U18034 (N_18034,N_17185,N_17182);
nand U18035 (N_18035,N_17351,N_16895);
and U18036 (N_18036,N_17151,N_17443);
or U18037 (N_18037,N_17054,N_17166);
nand U18038 (N_18038,N_17091,N_17066);
nor U18039 (N_18039,N_17212,N_17043);
nor U18040 (N_18040,N_17431,N_16900);
xnor U18041 (N_18041,N_17420,N_17233);
or U18042 (N_18042,N_17206,N_16909);
or U18043 (N_18043,N_17245,N_17336);
xnor U18044 (N_18044,N_17273,N_17084);
nor U18045 (N_18045,N_17306,N_17291);
nand U18046 (N_18046,N_17461,N_17032);
or U18047 (N_18047,N_17028,N_17085);
nand U18048 (N_18048,N_17079,N_17373);
or U18049 (N_18049,N_16893,N_17249);
and U18050 (N_18050,N_17090,N_17126);
nor U18051 (N_18051,N_17267,N_16932);
nor U18052 (N_18052,N_17301,N_17410);
and U18053 (N_18053,N_17341,N_17307);
or U18054 (N_18054,N_17164,N_17293);
nand U18055 (N_18055,N_17213,N_16943);
and U18056 (N_18056,N_17066,N_16988);
nand U18057 (N_18057,N_17276,N_16924);
or U18058 (N_18058,N_17157,N_17126);
or U18059 (N_18059,N_16885,N_17444);
and U18060 (N_18060,N_17383,N_17443);
or U18061 (N_18061,N_17403,N_17266);
nor U18062 (N_18062,N_17432,N_17378);
xor U18063 (N_18063,N_17344,N_17323);
and U18064 (N_18064,N_16944,N_17047);
xnor U18065 (N_18065,N_17086,N_17172);
or U18066 (N_18066,N_17333,N_17217);
xor U18067 (N_18067,N_17030,N_17494);
nand U18068 (N_18068,N_17431,N_16997);
or U18069 (N_18069,N_17441,N_17272);
or U18070 (N_18070,N_17067,N_16902);
xnor U18071 (N_18071,N_17123,N_17128);
or U18072 (N_18072,N_16960,N_16928);
and U18073 (N_18073,N_16993,N_17441);
nand U18074 (N_18074,N_17151,N_17465);
or U18075 (N_18075,N_17233,N_17086);
or U18076 (N_18076,N_17191,N_17189);
xnor U18077 (N_18077,N_17429,N_17299);
and U18078 (N_18078,N_16990,N_16877);
xor U18079 (N_18079,N_17200,N_17064);
and U18080 (N_18080,N_16937,N_16909);
or U18081 (N_18081,N_17049,N_16952);
nor U18082 (N_18082,N_17041,N_17113);
nor U18083 (N_18083,N_16881,N_17139);
or U18084 (N_18084,N_17208,N_16995);
or U18085 (N_18085,N_17158,N_17238);
and U18086 (N_18086,N_17007,N_17105);
nand U18087 (N_18087,N_16924,N_17466);
nor U18088 (N_18088,N_17396,N_17415);
xor U18089 (N_18089,N_17331,N_17306);
nor U18090 (N_18090,N_16942,N_17423);
or U18091 (N_18091,N_17362,N_17044);
nor U18092 (N_18092,N_17376,N_17372);
nand U18093 (N_18093,N_17185,N_16908);
nor U18094 (N_18094,N_17144,N_17386);
and U18095 (N_18095,N_17424,N_17263);
xnor U18096 (N_18096,N_17110,N_17344);
nand U18097 (N_18097,N_17360,N_17179);
or U18098 (N_18098,N_17380,N_16933);
xor U18099 (N_18099,N_17244,N_16971);
and U18100 (N_18100,N_17316,N_17202);
or U18101 (N_18101,N_17389,N_17162);
xor U18102 (N_18102,N_17177,N_17492);
or U18103 (N_18103,N_17358,N_17028);
nor U18104 (N_18104,N_17151,N_16976);
nand U18105 (N_18105,N_17078,N_16980);
and U18106 (N_18106,N_17248,N_17229);
and U18107 (N_18107,N_17367,N_17264);
and U18108 (N_18108,N_17092,N_17064);
or U18109 (N_18109,N_17260,N_17286);
and U18110 (N_18110,N_17408,N_17349);
xor U18111 (N_18111,N_17191,N_17281);
or U18112 (N_18112,N_16914,N_16968);
nor U18113 (N_18113,N_17371,N_17392);
nor U18114 (N_18114,N_16996,N_16890);
nor U18115 (N_18115,N_17458,N_17333);
nor U18116 (N_18116,N_16893,N_17168);
nor U18117 (N_18117,N_17357,N_17471);
nand U18118 (N_18118,N_17062,N_16877);
nand U18119 (N_18119,N_16927,N_17234);
xor U18120 (N_18120,N_17323,N_17281);
nor U18121 (N_18121,N_17452,N_17303);
xnor U18122 (N_18122,N_17009,N_16898);
and U18123 (N_18123,N_17391,N_17088);
nand U18124 (N_18124,N_17100,N_17460);
xnor U18125 (N_18125,N_17899,N_17782);
or U18126 (N_18126,N_17988,N_18104);
nor U18127 (N_18127,N_17944,N_17941);
xnor U18128 (N_18128,N_17893,N_17815);
xor U18129 (N_18129,N_17993,N_17875);
or U18130 (N_18130,N_18022,N_17938);
and U18131 (N_18131,N_17780,N_17730);
xnor U18132 (N_18132,N_17967,N_17719);
or U18133 (N_18133,N_17904,N_18051);
xnor U18134 (N_18134,N_17720,N_17871);
xnor U18135 (N_18135,N_17610,N_17616);
or U18136 (N_18136,N_17992,N_17521);
and U18137 (N_18137,N_17796,N_17697);
and U18138 (N_18138,N_17999,N_17688);
and U18139 (N_18139,N_17791,N_17576);
nor U18140 (N_18140,N_18105,N_17885);
or U18141 (N_18141,N_17593,N_18078);
nor U18142 (N_18142,N_17703,N_17590);
and U18143 (N_18143,N_17627,N_17809);
nor U18144 (N_18144,N_18048,N_18119);
nor U18145 (N_18145,N_17802,N_17755);
or U18146 (N_18146,N_17770,N_17951);
or U18147 (N_18147,N_17766,N_17784);
nor U18148 (N_18148,N_17563,N_17997);
or U18149 (N_18149,N_17526,N_17538);
xnor U18150 (N_18150,N_17775,N_18116);
and U18151 (N_18151,N_17693,N_18049);
or U18152 (N_18152,N_18080,N_17920);
or U18153 (N_18153,N_17671,N_18054);
and U18154 (N_18154,N_18031,N_17581);
or U18155 (N_18155,N_17772,N_17767);
nand U18156 (N_18156,N_18082,N_17573);
nor U18157 (N_18157,N_17669,N_18075);
nand U18158 (N_18158,N_17710,N_17965);
xor U18159 (N_18159,N_17761,N_17540);
or U18160 (N_18160,N_17886,N_17586);
nor U18161 (N_18161,N_17636,N_17624);
and U18162 (N_18162,N_17986,N_18065);
and U18163 (N_18163,N_18035,N_18053);
nand U18164 (N_18164,N_17634,N_17855);
xor U18165 (N_18165,N_17884,N_17783);
nand U18166 (N_18166,N_17959,N_18006);
nand U18167 (N_18167,N_18076,N_17830);
xor U18168 (N_18168,N_17918,N_17608);
nand U18169 (N_18169,N_17858,N_18044);
and U18170 (N_18170,N_17870,N_17571);
or U18171 (N_18171,N_17691,N_17905);
or U18172 (N_18172,N_17749,N_17942);
and U18173 (N_18173,N_17652,N_17642);
or U18174 (N_18174,N_17950,N_18028);
nor U18175 (N_18175,N_17917,N_17829);
nand U18176 (N_18176,N_17823,N_18036);
nor U18177 (N_18177,N_17790,N_17838);
xor U18178 (N_18178,N_17511,N_18072);
nand U18179 (N_18179,N_17923,N_18074);
nor U18180 (N_18180,N_17928,N_17776);
or U18181 (N_18181,N_18101,N_17851);
xnor U18182 (N_18182,N_18115,N_17699);
nand U18183 (N_18183,N_18000,N_18029);
nor U18184 (N_18184,N_17867,N_17759);
or U18185 (N_18185,N_17792,N_17544);
nand U18186 (N_18186,N_17512,N_17515);
nand U18187 (N_18187,N_17701,N_17713);
nand U18188 (N_18188,N_18045,N_17507);
xor U18189 (N_18189,N_18086,N_17737);
xnor U18190 (N_18190,N_17648,N_18109);
or U18191 (N_18191,N_17717,N_17700);
and U18192 (N_18192,N_17910,N_17975);
and U18193 (N_18193,N_17738,N_17556);
and U18194 (N_18194,N_17981,N_18114);
nor U18195 (N_18195,N_18093,N_17622);
nor U18196 (N_18196,N_17862,N_17650);
nor U18197 (N_18197,N_17668,N_17606);
or U18198 (N_18198,N_18061,N_18012);
xnor U18199 (N_18199,N_17646,N_17837);
and U18200 (N_18200,N_17712,N_17752);
or U18201 (N_18201,N_17629,N_17531);
nor U18202 (N_18202,N_18100,N_17872);
nand U18203 (N_18203,N_17553,N_17908);
nand U18204 (N_18204,N_17528,N_17747);
or U18205 (N_18205,N_17825,N_17869);
nand U18206 (N_18206,N_18071,N_18026);
xor U18207 (N_18207,N_17760,N_17618);
or U18208 (N_18208,N_17902,N_17647);
and U18209 (N_18209,N_17554,N_17534);
nor U18210 (N_18210,N_17572,N_17548);
nor U18211 (N_18211,N_17524,N_17961);
nand U18212 (N_18212,N_18102,N_17612);
and U18213 (N_18213,N_17504,N_17958);
nand U18214 (N_18214,N_18020,N_17503);
or U18215 (N_18215,N_18112,N_18039);
and U18216 (N_18216,N_17960,N_17707);
and U18217 (N_18217,N_17968,N_17810);
nor U18218 (N_18218,N_17841,N_17644);
xnor U18219 (N_18219,N_17694,N_17845);
nor U18220 (N_18220,N_17705,N_17501);
nor U18221 (N_18221,N_17532,N_18085);
nand U18222 (N_18222,N_18095,N_18097);
xnor U18223 (N_18223,N_17681,N_17769);
nand U18224 (N_18224,N_17682,N_17779);
or U18225 (N_18225,N_17660,N_17991);
and U18226 (N_18226,N_17550,N_18013);
xor U18227 (N_18227,N_17623,N_17639);
and U18228 (N_18228,N_18091,N_17708);
nor U18229 (N_18229,N_17580,N_17729);
nor U18230 (N_18230,N_18014,N_17846);
nand U18231 (N_18231,N_17926,N_17685);
nor U18232 (N_18232,N_17736,N_17709);
xor U18233 (N_18233,N_18034,N_18042);
or U18234 (N_18234,N_17847,N_17804);
or U18235 (N_18235,N_18041,N_17551);
xnor U18236 (N_18236,N_17848,N_17637);
xor U18237 (N_18237,N_17953,N_17964);
nand U18238 (N_18238,N_17843,N_18059);
nor U18239 (N_18239,N_17764,N_17750);
nor U18240 (N_18240,N_17666,N_17995);
or U18241 (N_18241,N_18001,N_17733);
and U18242 (N_18242,N_17596,N_17724);
xnor U18243 (N_18243,N_17814,N_17892);
nor U18244 (N_18244,N_18008,N_18010);
nor U18245 (N_18245,N_17781,N_17600);
nand U18246 (N_18246,N_17582,N_17541);
xnor U18247 (N_18247,N_17907,N_17665);
nor U18248 (N_18248,N_17765,N_17704);
and U18249 (N_18249,N_17990,N_17946);
nor U18250 (N_18250,N_17604,N_17773);
nand U18251 (N_18251,N_18098,N_17849);
or U18252 (N_18252,N_17741,N_17569);
nor U18253 (N_18253,N_17966,N_17913);
nor U18254 (N_18254,N_17661,N_17686);
nand U18255 (N_18255,N_17803,N_17527);
and U18256 (N_18256,N_17901,N_17565);
or U18257 (N_18257,N_17577,N_17891);
nor U18258 (N_18258,N_17833,N_17678);
nand U18259 (N_18259,N_17954,N_17864);
nand U18260 (N_18260,N_17989,N_17878);
nor U18261 (N_18261,N_18021,N_18124);
xor U18262 (N_18262,N_17840,N_17949);
xor U18263 (N_18263,N_17836,N_17529);
nor U18264 (N_18264,N_17732,N_17806);
nand U18265 (N_18265,N_17957,N_17900);
nor U18266 (N_18266,N_17785,N_18087);
nand U18267 (N_18267,N_17795,N_17692);
nor U18268 (N_18268,N_17638,N_17683);
xor U18269 (N_18269,N_17976,N_17658);
or U18270 (N_18270,N_17930,N_17500);
and U18271 (N_18271,N_17579,N_18073);
nor U18272 (N_18272,N_18062,N_17919);
nand U18273 (N_18273,N_18047,N_17863);
and U18274 (N_18274,N_18056,N_18108);
nand U18275 (N_18275,N_17695,N_17943);
or U18276 (N_18276,N_17906,N_17625);
nor U18277 (N_18277,N_18060,N_17522);
nor U18278 (N_18278,N_18079,N_17559);
nand U18279 (N_18279,N_18077,N_18122);
nor U18280 (N_18280,N_17832,N_18011);
xor U18281 (N_18281,N_17860,N_17630);
and U18282 (N_18282,N_17801,N_17628);
or U18283 (N_18283,N_17613,N_17757);
nor U18284 (N_18284,N_17876,N_17687);
nand U18285 (N_18285,N_17877,N_17653);
xnor U18286 (N_18286,N_17980,N_18024);
or U18287 (N_18287,N_17824,N_18052);
or U18288 (N_18288,N_17649,N_17510);
xor U18289 (N_18289,N_17994,N_17530);
nor U18290 (N_18290,N_17799,N_17711);
nor U18291 (N_18291,N_18019,N_17505);
nor U18292 (N_18292,N_17927,N_17952);
or U18293 (N_18293,N_17812,N_17599);
nand U18294 (N_18294,N_17575,N_17754);
nor U18295 (N_18295,N_17974,N_17727);
xnor U18296 (N_18296,N_17853,N_18017);
and U18297 (N_18297,N_17818,N_17977);
nor U18298 (N_18298,N_17535,N_17857);
nand U18299 (N_18299,N_17866,N_17543);
nand U18300 (N_18300,N_18007,N_17674);
or U18301 (N_18301,N_17735,N_17971);
or U18302 (N_18302,N_17798,N_17819);
and U18303 (N_18303,N_17520,N_17696);
and U18304 (N_18304,N_17962,N_17721);
xnor U18305 (N_18305,N_17585,N_17894);
or U18306 (N_18306,N_17880,N_17873);
nor U18307 (N_18307,N_18057,N_17523);
or U18308 (N_18308,N_17739,N_17898);
and U18309 (N_18309,N_17786,N_17982);
xnor U18310 (N_18310,N_17842,N_17537);
xor U18311 (N_18311,N_17929,N_17821);
xnor U18312 (N_18312,N_17883,N_17787);
xnor U18313 (N_18313,N_17595,N_17684);
xor U18314 (N_18314,N_17662,N_17984);
xnor U18315 (N_18315,N_18120,N_17656);
and U18316 (N_18316,N_17865,N_17698);
xnor U18317 (N_18317,N_17635,N_17558);
or U18318 (N_18318,N_17817,N_18009);
xnor U18319 (N_18319,N_17731,N_17879);
nor U18320 (N_18320,N_18058,N_17562);
nand U18321 (N_18321,N_17615,N_17714);
and U18322 (N_18322,N_18092,N_17777);
nor U18323 (N_18323,N_17690,N_17808);
or U18324 (N_18324,N_18003,N_17987);
xor U18325 (N_18325,N_17936,N_17723);
xor U18326 (N_18326,N_17746,N_17664);
nor U18327 (N_18327,N_17852,N_17659);
or U18328 (N_18328,N_17850,N_17722);
and U18329 (N_18329,N_17611,N_18096);
nand U18330 (N_18330,N_17956,N_18094);
and U18331 (N_18331,N_18121,N_17728);
nand U18332 (N_18332,N_18046,N_17868);
and U18333 (N_18333,N_18117,N_17516);
xnor U18334 (N_18334,N_17614,N_17542);
and U18335 (N_18335,N_18088,N_18016);
xnor U18336 (N_18336,N_17560,N_17859);
nand U18337 (N_18337,N_17602,N_17633);
nand U18338 (N_18338,N_17509,N_17589);
nor U18339 (N_18339,N_17963,N_17856);
xor U18340 (N_18340,N_17985,N_17831);
and U18341 (N_18341,N_17584,N_17771);
and U18342 (N_18342,N_18068,N_18015);
and U18343 (N_18343,N_17567,N_17932);
nor U18344 (N_18344,N_18123,N_17854);
and U18345 (N_18345,N_17566,N_17667);
nor U18346 (N_18346,N_18043,N_18025);
nor U18347 (N_18347,N_17948,N_17525);
nor U18348 (N_18348,N_17547,N_17912);
and U18349 (N_18349,N_17587,N_17725);
and U18350 (N_18350,N_18050,N_18113);
nand U18351 (N_18351,N_17751,N_17740);
nor U18352 (N_18352,N_17983,N_17549);
or U18353 (N_18353,N_17508,N_17621);
or U18354 (N_18354,N_18081,N_17679);
xor U18355 (N_18355,N_17839,N_17706);
or U18356 (N_18356,N_17574,N_17788);
xnor U18357 (N_18357,N_17916,N_17689);
xor U18358 (N_18358,N_18111,N_18118);
or U18359 (N_18359,N_18055,N_17670);
and U18360 (N_18360,N_17597,N_17887);
and U18361 (N_18361,N_17915,N_17677);
xor U18362 (N_18362,N_17718,N_17763);
or U18363 (N_18363,N_17546,N_17655);
or U18364 (N_18364,N_17758,N_17924);
and U18365 (N_18365,N_17591,N_17672);
nor U18366 (N_18366,N_17643,N_18038);
or U18367 (N_18367,N_17807,N_18083);
xor U18368 (N_18368,N_17617,N_17861);
and U18369 (N_18369,N_17895,N_17947);
xor U18370 (N_18370,N_17513,N_18084);
and U18371 (N_18371,N_17568,N_17619);
nor U18372 (N_18372,N_17970,N_17588);
nor U18373 (N_18373,N_18032,N_17925);
nand U18374 (N_18374,N_17756,N_17874);
nand U18375 (N_18375,N_17998,N_17518);
xor U18376 (N_18376,N_17794,N_17673);
nand U18377 (N_18377,N_17914,N_18004);
nand U18378 (N_18378,N_18002,N_17889);
nand U18379 (N_18379,N_17564,N_17502);
nor U18380 (N_18380,N_17545,N_17969);
nor U18381 (N_18381,N_18033,N_17578);
or U18382 (N_18382,N_17657,N_17654);
and U18383 (N_18383,N_17903,N_17922);
nor U18384 (N_18384,N_17937,N_17557);
or U18385 (N_18385,N_17607,N_17506);
nand U18386 (N_18386,N_17921,N_17774);
or U18387 (N_18387,N_17598,N_18107);
nor U18388 (N_18388,N_17882,N_17931);
nand U18389 (N_18389,N_17640,N_17805);
nor U18390 (N_18390,N_18103,N_17844);
or U18391 (N_18391,N_17539,N_17835);
nor U18392 (N_18392,N_17680,N_18018);
xnor U18393 (N_18393,N_17828,N_17603);
xnor U18394 (N_18394,N_17955,N_17519);
and U18395 (N_18395,N_17702,N_17797);
or U18396 (N_18396,N_17826,N_17514);
nand U18397 (N_18397,N_17676,N_17827);
or U18398 (N_18398,N_17978,N_17651);
nand U18399 (N_18399,N_17940,N_17813);
xor U18400 (N_18400,N_17973,N_17726);
or U18401 (N_18401,N_17609,N_17896);
and U18402 (N_18402,N_17793,N_17935);
xor U18403 (N_18403,N_17561,N_18064);
and U18404 (N_18404,N_18066,N_17536);
nand U18405 (N_18405,N_17555,N_17753);
xnor U18406 (N_18406,N_17645,N_17979);
and U18407 (N_18407,N_17768,N_17945);
and U18408 (N_18408,N_17601,N_18106);
and U18409 (N_18409,N_17552,N_17620);
and U18410 (N_18410,N_17939,N_17811);
nand U18411 (N_18411,N_17631,N_17816);
and U18412 (N_18412,N_17778,N_17734);
and U18413 (N_18413,N_17933,N_17583);
or U18414 (N_18414,N_17715,N_18005);
nand U18415 (N_18415,N_17934,N_17909);
nand U18416 (N_18416,N_17890,N_17605);
nor U18417 (N_18417,N_17744,N_17716);
and U18418 (N_18418,N_17570,N_17800);
nand U18419 (N_18419,N_18040,N_18110);
nor U18420 (N_18420,N_18037,N_17663);
nand U18421 (N_18421,N_17897,N_18069);
and U18422 (N_18422,N_18023,N_18030);
or U18423 (N_18423,N_17742,N_17972);
and U18424 (N_18424,N_18089,N_18027);
nand U18425 (N_18425,N_17675,N_17888);
and U18426 (N_18426,N_18067,N_18063);
or U18427 (N_18427,N_18090,N_17911);
xnor U18428 (N_18428,N_17632,N_18070);
xor U18429 (N_18429,N_17743,N_17594);
nand U18430 (N_18430,N_17762,N_17789);
nor U18431 (N_18431,N_17820,N_17881);
xnor U18432 (N_18432,N_17834,N_17517);
xnor U18433 (N_18433,N_17748,N_17745);
nand U18434 (N_18434,N_17641,N_18099);
xnor U18435 (N_18435,N_17592,N_17996);
xnor U18436 (N_18436,N_17533,N_17626);
nor U18437 (N_18437,N_17822,N_17850);
xnor U18438 (N_18438,N_17976,N_17684);
or U18439 (N_18439,N_17594,N_17520);
nor U18440 (N_18440,N_17772,N_18058);
nand U18441 (N_18441,N_17787,N_17540);
nand U18442 (N_18442,N_17624,N_17675);
nor U18443 (N_18443,N_18021,N_17545);
or U18444 (N_18444,N_17526,N_17724);
xnor U18445 (N_18445,N_18001,N_17952);
xor U18446 (N_18446,N_17848,N_18066);
nand U18447 (N_18447,N_17832,N_17701);
xnor U18448 (N_18448,N_17622,N_17723);
nor U18449 (N_18449,N_17513,N_18068);
and U18450 (N_18450,N_18108,N_18011);
or U18451 (N_18451,N_18053,N_18107);
nor U18452 (N_18452,N_17854,N_17936);
or U18453 (N_18453,N_17649,N_17542);
xnor U18454 (N_18454,N_18082,N_17884);
nor U18455 (N_18455,N_17575,N_17782);
xor U18456 (N_18456,N_17603,N_18071);
or U18457 (N_18457,N_17663,N_17588);
and U18458 (N_18458,N_17944,N_17946);
nand U18459 (N_18459,N_17827,N_17802);
xnor U18460 (N_18460,N_17596,N_17650);
and U18461 (N_18461,N_17765,N_17846);
or U18462 (N_18462,N_17604,N_17706);
xor U18463 (N_18463,N_17786,N_18113);
nor U18464 (N_18464,N_17579,N_17735);
nand U18465 (N_18465,N_17931,N_17813);
nand U18466 (N_18466,N_17900,N_17828);
nand U18467 (N_18467,N_18056,N_17835);
xnor U18468 (N_18468,N_17693,N_17825);
and U18469 (N_18469,N_17831,N_17920);
nor U18470 (N_18470,N_17913,N_17758);
nor U18471 (N_18471,N_17641,N_17650);
or U18472 (N_18472,N_17789,N_18110);
or U18473 (N_18473,N_17921,N_17659);
and U18474 (N_18474,N_17554,N_17836);
and U18475 (N_18475,N_18097,N_17902);
xor U18476 (N_18476,N_17749,N_17839);
or U18477 (N_18477,N_17842,N_17800);
or U18478 (N_18478,N_17980,N_17988);
xor U18479 (N_18479,N_17916,N_17664);
and U18480 (N_18480,N_18047,N_17857);
xor U18481 (N_18481,N_17880,N_18072);
or U18482 (N_18482,N_17956,N_17936);
nor U18483 (N_18483,N_17866,N_17724);
nand U18484 (N_18484,N_17854,N_17656);
nor U18485 (N_18485,N_17647,N_18056);
nor U18486 (N_18486,N_17740,N_18119);
or U18487 (N_18487,N_17552,N_17693);
nand U18488 (N_18488,N_17703,N_18108);
xnor U18489 (N_18489,N_17538,N_17622);
nor U18490 (N_18490,N_17706,N_18082);
xnor U18491 (N_18491,N_17776,N_17833);
or U18492 (N_18492,N_17803,N_18060);
and U18493 (N_18493,N_17531,N_18076);
and U18494 (N_18494,N_17878,N_17949);
nor U18495 (N_18495,N_17996,N_17650);
nand U18496 (N_18496,N_18061,N_18050);
nor U18497 (N_18497,N_17921,N_17741);
or U18498 (N_18498,N_17662,N_17574);
or U18499 (N_18499,N_18118,N_17563);
or U18500 (N_18500,N_17563,N_17531);
nand U18501 (N_18501,N_17593,N_17888);
and U18502 (N_18502,N_17852,N_18068);
nor U18503 (N_18503,N_18117,N_17847);
xor U18504 (N_18504,N_18054,N_17783);
nor U18505 (N_18505,N_17534,N_17958);
nor U18506 (N_18506,N_17890,N_17734);
nor U18507 (N_18507,N_17629,N_18049);
or U18508 (N_18508,N_17940,N_17545);
nor U18509 (N_18509,N_17613,N_17948);
xnor U18510 (N_18510,N_17852,N_17990);
or U18511 (N_18511,N_17928,N_17672);
nand U18512 (N_18512,N_18069,N_17552);
and U18513 (N_18513,N_18074,N_17952);
nand U18514 (N_18514,N_17810,N_17560);
and U18515 (N_18515,N_17995,N_17826);
or U18516 (N_18516,N_17784,N_17820);
nor U18517 (N_18517,N_17575,N_17632);
and U18518 (N_18518,N_17888,N_17954);
nand U18519 (N_18519,N_17951,N_18111);
xnor U18520 (N_18520,N_17956,N_17749);
and U18521 (N_18521,N_17960,N_17654);
nand U18522 (N_18522,N_17702,N_17717);
nor U18523 (N_18523,N_18066,N_17513);
nor U18524 (N_18524,N_17903,N_17871);
nor U18525 (N_18525,N_17921,N_17598);
xor U18526 (N_18526,N_17617,N_17677);
or U18527 (N_18527,N_17685,N_17654);
or U18528 (N_18528,N_18104,N_18001);
nor U18529 (N_18529,N_17833,N_17513);
or U18530 (N_18530,N_17960,N_17829);
and U18531 (N_18531,N_17881,N_18108);
nor U18532 (N_18532,N_17815,N_17648);
and U18533 (N_18533,N_18052,N_17600);
nand U18534 (N_18534,N_17900,N_17667);
nand U18535 (N_18535,N_18043,N_17558);
nand U18536 (N_18536,N_18071,N_17622);
nor U18537 (N_18537,N_17956,N_18052);
or U18538 (N_18538,N_18052,N_17688);
xor U18539 (N_18539,N_17988,N_17555);
nor U18540 (N_18540,N_17698,N_17708);
and U18541 (N_18541,N_17999,N_17664);
nor U18542 (N_18542,N_18021,N_17857);
xnor U18543 (N_18543,N_17887,N_17684);
xnor U18544 (N_18544,N_17522,N_17535);
nor U18545 (N_18545,N_17560,N_17951);
xnor U18546 (N_18546,N_17909,N_17970);
or U18547 (N_18547,N_17894,N_18112);
xor U18548 (N_18548,N_18103,N_17686);
and U18549 (N_18549,N_17714,N_17530);
and U18550 (N_18550,N_17984,N_17915);
xnor U18551 (N_18551,N_17924,N_17945);
nand U18552 (N_18552,N_17728,N_17889);
or U18553 (N_18553,N_18004,N_17975);
nand U18554 (N_18554,N_17509,N_17524);
and U18555 (N_18555,N_17510,N_18071);
nand U18556 (N_18556,N_17961,N_17563);
xnor U18557 (N_18557,N_17851,N_17699);
and U18558 (N_18558,N_18014,N_17590);
or U18559 (N_18559,N_18079,N_17705);
nor U18560 (N_18560,N_17571,N_17562);
nand U18561 (N_18561,N_18055,N_17983);
and U18562 (N_18562,N_17998,N_18097);
nand U18563 (N_18563,N_17891,N_17910);
or U18564 (N_18564,N_17885,N_17990);
xor U18565 (N_18565,N_17545,N_17505);
xnor U18566 (N_18566,N_18032,N_17848);
nand U18567 (N_18567,N_18086,N_17663);
and U18568 (N_18568,N_18098,N_17804);
nand U18569 (N_18569,N_17656,N_17795);
xor U18570 (N_18570,N_17860,N_17949);
and U18571 (N_18571,N_18020,N_17964);
nor U18572 (N_18572,N_17629,N_18073);
or U18573 (N_18573,N_17568,N_17988);
and U18574 (N_18574,N_17999,N_17950);
xor U18575 (N_18575,N_17726,N_17668);
and U18576 (N_18576,N_17769,N_17796);
and U18577 (N_18577,N_17743,N_17933);
or U18578 (N_18578,N_17894,N_18070);
nor U18579 (N_18579,N_17879,N_17522);
nor U18580 (N_18580,N_17720,N_17752);
and U18581 (N_18581,N_17725,N_18089);
xnor U18582 (N_18582,N_17551,N_17802);
and U18583 (N_18583,N_17913,N_17728);
nand U18584 (N_18584,N_17535,N_17873);
xor U18585 (N_18585,N_18093,N_18025);
xnor U18586 (N_18586,N_17837,N_17513);
nor U18587 (N_18587,N_17810,N_17730);
xor U18588 (N_18588,N_17929,N_17755);
and U18589 (N_18589,N_17681,N_17679);
xnor U18590 (N_18590,N_18016,N_17557);
nor U18591 (N_18591,N_17787,N_17621);
nand U18592 (N_18592,N_17878,N_17850);
nor U18593 (N_18593,N_17737,N_17592);
nand U18594 (N_18594,N_17505,N_17504);
and U18595 (N_18595,N_17715,N_18090);
nor U18596 (N_18596,N_17793,N_17815);
xnor U18597 (N_18597,N_17664,N_17826);
or U18598 (N_18598,N_18029,N_17696);
or U18599 (N_18599,N_17571,N_17658);
and U18600 (N_18600,N_17819,N_18112);
and U18601 (N_18601,N_18087,N_17827);
xor U18602 (N_18602,N_17564,N_18086);
or U18603 (N_18603,N_17961,N_17900);
or U18604 (N_18604,N_17590,N_17672);
nand U18605 (N_18605,N_17717,N_17730);
and U18606 (N_18606,N_18027,N_18072);
nor U18607 (N_18607,N_17899,N_17625);
and U18608 (N_18608,N_17904,N_17774);
or U18609 (N_18609,N_18090,N_17898);
and U18610 (N_18610,N_17794,N_17577);
nand U18611 (N_18611,N_17735,N_18015);
xor U18612 (N_18612,N_18037,N_17636);
nor U18613 (N_18613,N_17877,N_17610);
and U18614 (N_18614,N_17576,N_17881);
nor U18615 (N_18615,N_17933,N_17619);
nand U18616 (N_18616,N_18082,N_17609);
and U18617 (N_18617,N_18030,N_17873);
or U18618 (N_18618,N_17871,N_17591);
nor U18619 (N_18619,N_17807,N_17505);
and U18620 (N_18620,N_17751,N_17586);
or U18621 (N_18621,N_17710,N_17758);
and U18622 (N_18622,N_17834,N_17975);
or U18623 (N_18623,N_17829,N_18106);
or U18624 (N_18624,N_17786,N_18097);
and U18625 (N_18625,N_17991,N_17979);
xor U18626 (N_18626,N_17858,N_17892);
or U18627 (N_18627,N_17615,N_17786);
xnor U18628 (N_18628,N_17847,N_18107);
nor U18629 (N_18629,N_18079,N_17663);
xnor U18630 (N_18630,N_17923,N_17927);
and U18631 (N_18631,N_17782,N_18042);
or U18632 (N_18632,N_17505,N_18015);
xnor U18633 (N_18633,N_17792,N_17782);
or U18634 (N_18634,N_17544,N_18059);
or U18635 (N_18635,N_18061,N_18085);
or U18636 (N_18636,N_17867,N_18000);
or U18637 (N_18637,N_17835,N_17942);
or U18638 (N_18638,N_17965,N_17747);
nand U18639 (N_18639,N_17818,N_17980);
nand U18640 (N_18640,N_17562,N_17537);
xor U18641 (N_18641,N_18083,N_17744);
or U18642 (N_18642,N_17824,N_17984);
and U18643 (N_18643,N_17568,N_17532);
nor U18644 (N_18644,N_18106,N_17795);
nand U18645 (N_18645,N_18026,N_17530);
and U18646 (N_18646,N_17590,N_17805);
nor U18647 (N_18647,N_17932,N_17659);
nand U18648 (N_18648,N_17530,N_17918);
or U18649 (N_18649,N_17768,N_17993);
xor U18650 (N_18650,N_18083,N_18027);
nor U18651 (N_18651,N_17553,N_18086);
nand U18652 (N_18652,N_17929,N_17700);
xnor U18653 (N_18653,N_17900,N_17950);
nor U18654 (N_18654,N_17799,N_17744);
or U18655 (N_18655,N_17925,N_18117);
or U18656 (N_18656,N_17741,N_17837);
or U18657 (N_18657,N_17700,N_17751);
nand U18658 (N_18658,N_17723,N_17721);
and U18659 (N_18659,N_17543,N_17894);
nor U18660 (N_18660,N_17827,N_17656);
and U18661 (N_18661,N_17995,N_17729);
xnor U18662 (N_18662,N_17775,N_17954);
nor U18663 (N_18663,N_17846,N_17854);
xnor U18664 (N_18664,N_18084,N_18020);
nor U18665 (N_18665,N_17716,N_17698);
nor U18666 (N_18666,N_17668,N_17981);
and U18667 (N_18667,N_17746,N_17503);
nor U18668 (N_18668,N_17671,N_17707);
or U18669 (N_18669,N_17600,N_17971);
xor U18670 (N_18670,N_18121,N_18076);
nand U18671 (N_18671,N_18084,N_17680);
nand U18672 (N_18672,N_17765,N_17503);
and U18673 (N_18673,N_17886,N_17909);
nand U18674 (N_18674,N_17942,N_17764);
nand U18675 (N_18675,N_17645,N_17938);
and U18676 (N_18676,N_17820,N_17958);
nand U18677 (N_18677,N_17841,N_17811);
nor U18678 (N_18678,N_17609,N_18084);
or U18679 (N_18679,N_17770,N_17695);
or U18680 (N_18680,N_17992,N_17911);
xnor U18681 (N_18681,N_17789,N_17865);
xnor U18682 (N_18682,N_18073,N_18031);
xor U18683 (N_18683,N_17772,N_17632);
xnor U18684 (N_18684,N_18089,N_17911);
and U18685 (N_18685,N_17534,N_18001);
xnor U18686 (N_18686,N_18099,N_17610);
nand U18687 (N_18687,N_17551,N_17756);
nor U18688 (N_18688,N_17654,N_17983);
nand U18689 (N_18689,N_18068,N_17554);
nor U18690 (N_18690,N_18107,N_17981);
nand U18691 (N_18691,N_17818,N_17726);
xnor U18692 (N_18692,N_17987,N_17750);
and U18693 (N_18693,N_17810,N_18117);
or U18694 (N_18694,N_17777,N_18003);
xnor U18695 (N_18695,N_18009,N_17803);
nor U18696 (N_18696,N_17665,N_18057);
xnor U18697 (N_18697,N_17627,N_17723);
nand U18698 (N_18698,N_17861,N_17828);
nand U18699 (N_18699,N_17641,N_17672);
and U18700 (N_18700,N_17687,N_17741);
nand U18701 (N_18701,N_17675,N_17822);
nand U18702 (N_18702,N_17677,N_17935);
and U18703 (N_18703,N_17630,N_18109);
nor U18704 (N_18704,N_17754,N_17804);
or U18705 (N_18705,N_17852,N_17778);
nor U18706 (N_18706,N_17978,N_18044);
nand U18707 (N_18707,N_17570,N_17572);
and U18708 (N_18708,N_17921,N_17780);
nor U18709 (N_18709,N_17611,N_17841);
or U18710 (N_18710,N_17597,N_17567);
nor U18711 (N_18711,N_17722,N_17790);
nand U18712 (N_18712,N_17679,N_17844);
or U18713 (N_18713,N_17739,N_17930);
and U18714 (N_18714,N_17608,N_17695);
nand U18715 (N_18715,N_18038,N_17816);
xor U18716 (N_18716,N_17591,N_17622);
or U18717 (N_18717,N_17938,N_17866);
nor U18718 (N_18718,N_18041,N_17597);
xnor U18719 (N_18719,N_18013,N_18024);
or U18720 (N_18720,N_17701,N_17664);
nor U18721 (N_18721,N_17513,N_18085);
xnor U18722 (N_18722,N_18017,N_17851);
nor U18723 (N_18723,N_17734,N_18059);
and U18724 (N_18724,N_18043,N_18056);
or U18725 (N_18725,N_17824,N_17579);
and U18726 (N_18726,N_17574,N_17720);
or U18727 (N_18727,N_17940,N_17797);
or U18728 (N_18728,N_17849,N_17550);
and U18729 (N_18729,N_17835,N_17922);
nand U18730 (N_18730,N_18061,N_17606);
or U18731 (N_18731,N_17582,N_17918);
nand U18732 (N_18732,N_17697,N_17914);
nor U18733 (N_18733,N_18105,N_18119);
and U18734 (N_18734,N_17875,N_17561);
and U18735 (N_18735,N_18102,N_18039);
nor U18736 (N_18736,N_17822,N_18065);
and U18737 (N_18737,N_17860,N_17675);
xnor U18738 (N_18738,N_17644,N_17817);
or U18739 (N_18739,N_18094,N_18082);
xnor U18740 (N_18740,N_17612,N_17994);
nand U18741 (N_18741,N_17901,N_18040);
xnor U18742 (N_18742,N_18051,N_17903);
or U18743 (N_18743,N_17584,N_17630);
or U18744 (N_18744,N_18084,N_17707);
nor U18745 (N_18745,N_17546,N_17680);
and U18746 (N_18746,N_18010,N_18066);
or U18747 (N_18747,N_17735,N_17537);
nand U18748 (N_18748,N_17706,N_17507);
and U18749 (N_18749,N_18017,N_17667);
xnor U18750 (N_18750,N_18560,N_18544);
nor U18751 (N_18751,N_18281,N_18173);
and U18752 (N_18752,N_18688,N_18710);
or U18753 (N_18753,N_18714,N_18335);
or U18754 (N_18754,N_18383,N_18210);
and U18755 (N_18755,N_18378,N_18271);
nor U18756 (N_18756,N_18564,N_18324);
and U18757 (N_18757,N_18503,N_18429);
and U18758 (N_18758,N_18589,N_18581);
nor U18759 (N_18759,N_18627,N_18336);
nand U18760 (N_18760,N_18571,N_18616);
or U18761 (N_18761,N_18224,N_18229);
nor U18762 (N_18762,N_18657,N_18708);
xnor U18763 (N_18763,N_18275,N_18142);
nand U18764 (N_18764,N_18143,N_18456);
xnor U18765 (N_18765,N_18370,N_18240);
xnor U18766 (N_18766,N_18339,N_18608);
nor U18767 (N_18767,N_18220,N_18660);
or U18768 (N_18768,N_18158,N_18464);
and U18769 (N_18769,N_18128,N_18368);
nor U18770 (N_18770,N_18527,N_18215);
xor U18771 (N_18771,N_18524,N_18314);
xor U18772 (N_18772,N_18737,N_18591);
and U18773 (N_18773,N_18323,N_18572);
and U18774 (N_18774,N_18167,N_18685);
nand U18775 (N_18775,N_18172,N_18310);
xnor U18776 (N_18776,N_18605,N_18562);
xor U18777 (N_18777,N_18146,N_18397);
nor U18778 (N_18778,N_18197,N_18595);
and U18779 (N_18779,N_18318,N_18648);
or U18780 (N_18780,N_18625,N_18175);
nand U18781 (N_18781,N_18325,N_18157);
nand U18782 (N_18782,N_18398,N_18443);
nor U18783 (N_18783,N_18460,N_18408);
or U18784 (N_18784,N_18668,N_18635);
nor U18785 (N_18785,N_18301,N_18206);
and U18786 (N_18786,N_18150,N_18534);
or U18787 (N_18787,N_18593,N_18191);
and U18788 (N_18788,N_18289,N_18435);
nand U18789 (N_18789,N_18252,N_18543);
and U18790 (N_18790,N_18662,N_18586);
nand U18791 (N_18791,N_18386,N_18154);
xnor U18792 (N_18792,N_18419,N_18396);
nand U18793 (N_18793,N_18288,N_18343);
nand U18794 (N_18794,N_18719,N_18187);
and U18795 (N_18795,N_18319,N_18259);
and U18796 (N_18796,N_18156,N_18748);
and U18797 (N_18797,N_18451,N_18497);
nand U18798 (N_18798,N_18476,N_18282);
nand U18799 (N_18799,N_18365,N_18274);
nand U18800 (N_18800,N_18516,N_18701);
xnor U18801 (N_18801,N_18494,N_18413);
and U18802 (N_18802,N_18739,N_18705);
xor U18803 (N_18803,N_18184,N_18717);
xnor U18804 (N_18804,N_18269,N_18461);
and U18805 (N_18805,N_18514,N_18328);
and U18806 (N_18806,N_18345,N_18607);
xnor U18807 (N_18807,N_18392,N_18499);
nand U18808 (N_18808,N_18257,N_18663);
nand U18809 (N_18809,N_18350,N_18638);
xor U18810 (N_18810,N_18471,N_18576);
nand U18811 (N_18811,N_18330,N_18528);
or U18812 (N_18812,N_18641,N_18412);
nand U18813 (N_18813,N_18130,N_18377);
xor U18814 (N_18814,N_18478,N_18284);
xor U18815 (N_18815,N_18311,N_18263);
and U18816 (N_18816,N_18691,N_18632);
or U18817 (N_18817,N_18587,N_18148);
xnor U18818 (N_18818,N_18504,N_18305);
or U18819 (N_18819,N_18585,N_18568);
xnor U18820 (N_18820,N_18747,N_18420);
nor U18821 (N_18821,N_18555,N_18556);
nor U18822 (N_18822,N_18549,N_18293);
nand U18823 (N_18823,N_18236,N_18518);
xor U18824 (N_18824,N_18487,N_18457);
and U18825 (N_18825,N_18453,N_18597);
nor U18826 (N_18826,N_18447,N_18351);
or U18827 (N_18827,N_18127,N_18380);
nor U18828 (N_18828,N_18250,N_18715);
xnor U18829 (N_18829,N_18190,N_18394);
xnor U18830 (N_18830,N_18431,N_18302);
or U18831 (N_18831,N_18432,N_18683);
nand U18832 (N_18832,N_18165,N_18481);
nand U18833 (N_18833,N_18132,N_18211);
or U18834 (N_18834,N_18465,N_18410);
or U18835 (N_18835,N_18619,N_18277);
or U18836 (N_18836,N_18601,N_18170);
xor U18837 (N_18837,N_18505,N_18131);
nor U18838 (N_18838,N_18462,N_18709);
nand U18839 (N_18839,N_18234,N_18452);
and U18840 (N_18840,N_18455,N_18653);
or U18841 (N_18841,N_18634,N_18253);
xor U18842 (N_18842,N_18295,N_18508);
and U18843 (N_18843,N_18574,N_18696);
nand U18844 (N_18844,N_18369,N_18539);
nor U18845 (N_18845,N_18602,N_18569);
xor U18846 (N_18846,N_18567,N_18164);
nand U18847 (N_18847,N_18332,N_18260);
xnor U18848 (N_18848,N_18686,N_18376);
or U18849 (N_18849,N_18270,N_18306);
nor U18850 (N_18850,N_18375,N_18561);
nor U18851 (N_18851,N_18160,N_18525);
or U18852 (N_18852,N_18553,N_18590);
nor U18853 (N_18853,N_18440,N_18340);
or U18854 (N_18854,N_18326,N_18520);
or U18855 (N_18855,N_18312,N_18613);
nand U18856 (N_18856,N_18303,N_18235);
nor U18857 (N_18857,N_18353,N_18268);
nor U18858 (N_18858,N_18584,N_18149);
nor U18859 (N_18859,N_18171,N_18205);
nor U18860 (N_18860,N_18519,N_18321);
nor U18861 (N_18861,N_18427,N_18675);
nor U18862 (N_18862,N_18139,N_18741);
or U18863 (N_18863,N_18283,N_18680);
nor U18864 (N_18864,N_18484,N_18218);
or U18865 (N_18865,N_18728,N_18198);
xor U18866 (N_18866,N_18145,N_18551);
or U18867 (N_18867,N_18612,N_18459);
nor U18868 (N_18868,N_18298,N_18473);
or U18869 (N_18869,N_18698,N_18722);
and U18870 (N_18870,N_18249,N_18266);
or U18871 (N_18871,N_18533,N_18406);
nor U18872 (N_18872,N_18529,N_18384);
or U18873 (N_18873,N_18687,N_18322);
nand U18874 (N_18874,N_18341,N_18292);
and U18875 (N_18875,N_18162,N_18600);
nand U18876 (N_18876,N_18645,N_18547);
nand U18877 (N_18877,N_18189,N_18407);
nor U18878 (N_18878,N_18690,N_18573);
nor U18879 (N_18879,N_18347,N_18617);
xnor U18880 (N_18880,N_18671,N_18530);
nand U18881 (N_18881,N_18209,N_18570);
nor U18882 (N_18882,N_18542,N_18193);
and U18883 (N_18883,N_18490,N_18517);
and U18884 (N_18884,N_18689,N_18214);
or U18885 (N_18885,N_18241,N_18446);
and U18886 (N_18886,N_18161,N_18618);
or U18887 (N_18887,N_18649,N_18466);
and U18888 (N_18888,N_18624,N_18694);
or U18889 (N_18889,N_18180,N_18444);
and U18890 (N_18890,N_18201,N_18577);
xnor U18891 (N_18891,N_18434,N_18422);
nand U18892 (N_18892,N_18475,N_18230);
nand U18893 (N_18893,N_18313,N_18418);
nor U18894 (N_18894,N_18196,N_18672);
or U18895 (N_18895,N_18639,N_18513);
or U18896 (N_18896,N_18631,N_18223);
or U18897 (N_18897,N_18450,N_18448);
nor U18898 (N_18898,N_18381,N_18136);
and U18899 (N_18899,N_18592,N_18192);
and U18900 (N_18900,N_18548,N_18507);
xnor U18901 (N_18901,N_18238,N_18644);
or U18902 (N_18902,N_18633,N_18417);
or U18903 (N_18903,N_18509,N_18256);
and U18904 (N_18904,N_18628,N_18362);
and U18905 (N_18905,N_18134,N_18399);
and U18906 (N_18906,N_18402,N_18267);
or U18907 (N_18907,N_18183,N_18174);
xnor U18908 (N_18908,N_18338,N_18656);
nor U18909 (N_18909,N_18512,N_18379);
and U18910 (N_18910,N_18329,N_18285);
xor U18911 (N_18911,N_18225,N_18575);
and U18912 (N_18912,N_18536,N_18711);
nand U18913 (N_18913,N_18299,N_18538);
or U18914 (N_18914,N_18439,N_18674);
nor U18915 (N_18915,N_18185,N_18188);
xnor U18916 (N_18916,N_18501,N_18309);
and U18917 (N_18917,N_18203,N_18231);
nor U18918 (N_18918,N_18526,N_18469);
nor U18919 (N_18919,N_18428,N_18470);
nand U18920 (N_18920,N_18337,N_18578);
and U18921 (N_18921,N_18491,N_18153);
xor U18922 (N_18922,N_18678,N_18565);
nor U18923 (N_18923,N_18409,N_18178);
nor U18924 (N_18924,N_18580,N_18272);
nand U18925 (N_18925,N_18726,N_18673);
nand U18926 (N_18926,N_18506,N_18261);
and U18927 (N_18927,N_18721,N_18364);
or U18928 (N_18928,N_18498,N_18354);
xnor U18929 (N_18929,N_18712,N_18411);
xor U18930 (N_18930,N_18194,N_18489);
or U18931 (N_18931,N_18738,N_18403);
nor U18932 (N_18932,N_18242,N_18135);
nand U18933 (N_18933,N_18125,N_18226);
nand U18934 (N_18934,N_18287,N_18286);
or U18935 (N_18935,N_18598,N_18342);
nor U18936 (N_18936,N_18221,N_18488);
and U18937 (N_18937,N_18290,N_18233);
nand U18938 (N_18938,N_18692,N_18137);
xnor U18939 (N_18939,N_18730,N_18317);
nor U18940 (N_18940,N_18308,N_18623);
and U18941 (N_18941,N_18344,N_18316);
nand U18942 (N_18942,N_18636,N_18141);
xor U18943 (N_18943,N_18749,N_18733);
and U18944 (N_18944,N_18596,N_18546);
or U18945 (N_18945,N_18151,N_18248);
nand U18946 (N_18946,N_18258,N_18480);
nand U18947 (N_18947,N_18449,N_18155);
nand U18948 (N_18948,N_18729,N_18199);
nand U18949 (N_18949,N_18346,N_18725);
xor U18950 (N_18950,N_18495,N_18640);
and U18951 (N_18951,N_18693,N_18247);
nor U18952 (N_18952,N_18670,N_18723);
xnor U18953 (N_18953,N_18176,N_18716);
nand U18954 (N_18954,N_18361,N_18442);
xor U18955 (N_18955,N_18642,N_18445);
nand U18956 (N_18956,N_18382,N_18219);
nand U18957 (N_18957,N_18352,N_18621);
or U18958 (N_18958,N_18264,N_18280);
nand U18959 (N_18959,N_18666,N_18742);
and U18960 (N_18960,N_18731,N_18604);
nor U18961 (N_18961,N_18637,N_18493);
nand U18962 (N_18962,N_18706,N_18727);
or U18963 (N_18963,N_18676,N_18679);
nor U18964 (N_18964,N_18239,N_18232);
xor U18965 (N_18965,N_18357,N_18331);
or U18966 (N_18966,N_18646,N_18647);
and U18967 (N_18967,N_18208,N_18168);
or U18968 (N_18968,N_18179,N_18744);
and U18969 (N_18969,N_18521,N_18579);
nor U18970 (N_18970,N_18182,N_18366);
or U18971 (N_18971,N_18677,N_18129);
nand U18972 (N_18972,N_18522,N_18421);
or U18973 (N_18973,N_18404,N_18159);
and U18974 (N_18974,N_18485,N_18273);
nand U18975 (N_18975,N_18294,N_18279);
nor U18976 (N_18976,N_18395,N_18416);
and U18977 (N_18977,N_18320,N_18724);
nand U18978 (N_18978,N_18745,N_18486);
xor U18979 (N_18979,N_18603,N_18643);
xor U18980 (N_18980,N_18550,N_18177);
nand U18981 (N_18981,N_18746,N_18393);
nand U18982 (N_18982,N_18474,N_18140);
nor U18983 (N_18983,N_18371,N_18734);
and U18984 (N_18984,N_18246,N_18265);
and U18985 (N_18985,N_18718,N_18307);
xnor U18986 (N_18986,N_18667,N_18207);
and U18987 (N_18987,N_18222,N_18212);
nand U18988 (N_18988,N_18515,N_18463);
xnor U18989 (N_18989,N_18611,N_18372);
xnor U18990 (N_18990,N_18620,N_18610);
or U18991 (N_18991,N_18669,N_18554);
and U18992 (N_18992,N_18682,N_18437);
or U18993 (N_18993,N_18588,N_18699);
or U18994 (N_18994,N_18483,N_18540);
or U18995 (N_18995,N_18359,N_18583);
and U18996 (N_18996,N_18424,N_18296);
nor U18997 (N_18997,N_18423,N_18626);
and U18998 (N_18998,N_18144,N_18472);
xnor U18999 (N_18999,N_18438,N_18531);
and U19000 (N_19000,N_18496,N_18532);
and U19001 (N_19001,N_18251,N_18652);
xor U19002 (N_19002,N_18700,N_18436);
nor U19003 (N_19003,N_18622,N_18736);
nor U19004 (N_19004,N_18401,N_18358);
nor U19005 (N_19005,N_18743,N_18213);
nor U19006 (N_19006,N_18441,N_18390);
or U19007 (N_19007,N_18228,N_18126);
and U19008 (N_19008,N_18426,N_18433);
and U19009 (N_19009,N_18245,N_18454);
and U19010 (N_19010,N_18732,N_18348);
nand U19011 (N_19011,N_18181,N_18511);
and U19012 (N_19012,N_18166,N_18629);
and U19013 (N_19013,N_18237,N_18684);
xor U19014 (N_19014,N_18650,N_18468);
nand U19015 (N_19015,N_18255,N_18606);
xnor U19016 (N_19016,N_18415,N_18186);
xnor U19017 (N_19017,N_18510,N_18664);
and U19018 (N_19018,N_18467,N_18300);
nand U19019 (N_19019,N_18388,N_18492);
or U19020 (N_19020,N_18349,N_18557);
xor U19021 (N_19021,N_18374,N_18630);
nand U19022 (N_19022,N_18704,N_18363);
xor U19023 (N_19023,N_18661,N_18315);
or U19024 (N_19024,N_18367,N_18425);
xnor U19025 (N_19025,N_18535,N_18615);
nor U19026 (N_19026,N_18740,N_18477);
or U19027 (N_19027,N_18216,N_18243);
and U19028 (N_19028,N_18655,N_18720);
or U19029 (N_19029,N_18482,N_18334);
xnor U19030 (N_19030,N_18502,N_18360);
or U19031 (N_19031,N_18244,N_18703);
or U19032 (N_19032,N_18195,N_18387);
nor U19033 (N_19033,N_18566,N_18479);
or U19034 (N_19034,N_18697,N_18658);
nor U19035 (N_19035,N_18659,N_18707);
nand U19036 (N_19036,N_18202,N_18389);
nand U19037 (N_19037,N_18430,N_18541);
or U19038 (N_19038,N_18291,N_18563);
nand U19039 (N_19039,N_18254,N_18278);
nor U19040 (N_19040,N_18400,N_18169);
xnor U19041 (N_19041,N_18414,N_18385);
nand U19042 (N_19042,N_18333,N_18594);
nor U19043 (N_19043,N_18405,N_18276);
xnor U19044 (N_19044,N_18138,N_18500);
and U19045 (N_19045,N_18163,N_18552);
and U19046 (N_19046,N_18262,N_18559);
nor U19047 (N_19047,N_18558,N_18599);
and U19048 (N_19048,N_18651,N_18204);
or U19049 (N_19049,N_18152,N_18297);
or U19050 (N_19050,N_18537,N_18355);
nor U19051 (N_19051,N_18200,N_18654);
or U19052 (N_19052,N_18695,N_18304);
or U19053 (N_19053,N_18458,N_18523);
and U19054 (N_19054,N_18665,N_18614);
nor U19055 (N_19055,N_18681,N_18227);
or U19056 (N_19056,N_18217,N_18391);
or U19057 (N_19057,N_18373,N_18582);
or U19058 (N_19058,N_18609,N_18702);
nor U19059 (N_19059,N_18735,N_18356);
or U19060 (N_19060,N_18545,N_18147);
nor U19061 (N_19061,N_18713,N_18133);
xor U19062 (N_19062,N_18327,N_18336);
xnor U19063 (N_19063,N_18228,N_18217);
or U19064 (N_19064,N_18143,N_18555);
nand U19065 (N_19065,N_18362,N_18635);
nor U19066 (N_19066,N_18730,N_18681);
or U19067 (N_19067,N_18522,N_18501);
or U19068 (N_19068,N_18477,N_18470);
and U19069 (N_19069,N_18222,N_18229);
or U19070 (N_19070,N_18334,N_18710);
or U19071 (N_19071,N_18169,N_18135);
nor U19072 (N_19072,N_18253,N_18349);
and U19073 (N_19073,N_18727,N_18523);
and U19074 (N_19074,N_18159,N_18515);
nand U19075 (N_19075,N_18505,N_18520);
xnor U19076 (N_19076,N_18367,N_18531);
nand U19077 (N_19077,N_18608,N_18630);
nor U19078 (N_19078,N_18328,N_18599);
nor U19079 (N_19079,N_18524,N_18487);
or U19080 (N_19080,N_18274,N_18589);
nand U19081 (N_19081,N_18165,N_18497);
xor U19082 (N_19082,N_18643,N_18450);
xnor U19083 (N_19083,N_18304,N_18369);
nor U19084 (N_19084,N_18229,N_18733);
xor U19085 (N_19085,N_18672,N_18628);
nor U19086 (N_19086,N_18401,N_18428);
or U19087 (N_19087,N_18672,N_18480);
nor U19088 (N_19088,N_18357,N_18341);
nor U19089 (N_19089,N_18678,N_18379);
xnor U19090 (N_19090,N_18232,N_18202);
or U19091 (N_19091,N_18555,N_18584);
or U19092 (N_19092,N_18292,N_18390);
nor U19093 (N_19093,N_18336,N_18304);
and U19094 (N_19094,N_18605,N_18464);
nand U19095 (N_19095,N_18338,N_18254);
xor U19096 (N_19096,N_18165,N_18187);
nand U19097 (N_19097,N_18389,N_18512);
nand U19098 (N_19098,N_18132,N_18634);
and U19099 (N_19099,N_18151,N_18264);
and U19100 (N_19100,N_18373,N_18284);
xor U19101 (N_19101,N_18357,N_18622);
or U19102 (N_19102,N_18409,N_18679);
or U19103 (N_19103,N_18468,N_18207);
and U19104 (N_19104,N_18294,N_18354);
or U19105 (N_19105,N_18687,N_18580);
xor U19106 (N_19106,N_18720,N_18195);
nand U19107 (N_19107,N_18726,N_18308);
nand U19108 (N_19108,N_18364,N_18156);
nor U19109 (N_19109,N_18291,N_18155);
or U19110 (N_19110,N_18485,N_18140);
xor U19111 (N_19111,N_18631,N_18149);
nand U19112 (N_19112,N_18444,N_18250);
and U19113 (N_19113,N_18308,N_18263);
or U19114 (N_19114,N_18329,N_18747);
or U19115 (N_19115,N_18275,N_18194);
xnor U19116 (N_19116,N_18343,N_18560);
xor U19117 (N_19117,N_18326,N_18592);
or U19118 (N_19118,N_18476,N_18210);
nor U19119 (N_19119,N_18373,N_18712);
and U19120 (N_19120,N_18446,N_18266);
xnor U19121 (N_19121,N_18199,N_18373);
or U19122 (N_19122,N_18355,N_18729);
xor U19123 (N_19123,N_18612,N_18317);
or U19124 (N_19124,N_18241,N_18360);
nor U19125 (N_19125,N_18158,N_18135);
or U19126 (N_19126,N_18706,N_18407);
nor U19127 (N_19127,N_18225,N_18374);
xor U19128 (N_19128,N_18211,N_18640);
nor U19129 (N_19129,N_18283,N_18534);
or U19130 (N_19130,N_18198,N_18398);
nor U19131 (N_19131,N_18506,N_18237);
xnor U19132 (N_19132,N_18633,N_18248);
and U19133 (N_19133,N_18331,N_18704);
nand U19134 (N_19134,N_18188,N_18700);
and U19135 (N_19135,N_18623,N_18525);
and U19136 (N_19136,N_18662,N_18465);
or U19137 (N_19137,N_18593,N_18355);
and U19138 (N_19138,N_18210,N_18146);
nand U19139 (N_19139,N_18165,N_18548);
xnor U19140 (N_19140,N_18137,N_18719);
nand U19141 (N_19141,N_18688,N_18247);
and U19142 (N_19142,N_18722,N_18359);
nand U19143 (N_19143,N_18407,N_18364);
nand U19144 (N_19144,N_18544,N_18709);
and U19145 (N_19145,N_18515,N_18402);
nor U19146 (N_19146,N_18668,N_18461);
nand U19147 (N_19147,N_18277,N_18696);
and U19148 (N_19148,N_18364,N_18422);
and U19149 (N_19149,N_18483,N_18329);
nor U19150 (N_19150,N_18555,N_18672);
nor U19151 (N_19151,N_18595,N_18719);
nand U19152 (N_19152,N_18288,N_18269);
or U19153 (N_19153,N_18452,N_18229);
xnor U19154 (N_19154,N_18409,N_18172);
nand U19155 (N_19155,N_18692,N_18267);
nor U19156 (N_19156,N_18607,N_18539);
xnor U19157 (N_19157,N_18605,N_18594);
or U19158 (N_19158,N_18688,N_18690);
or U19159 (N_19159,N_18624,N_18267);
nor U19160 (N_19160,N_18275,N_18200);
xor U19161 (N_19161,N_18410,N_18732);
or U19162 (N_19162,N_18451,N_18568);
or U19163 (N_19163,N_18485,N_18639);
nor U19164 (N_19164,N_18366,N_18536);
nor U19165 (N_19165,N_18670,N_18379);
nand U19166 (N_19166,N_18581,N_18575);
nand U19167 (N_19167,N_18237,N_18140);
xor U19168 (N_19168,N_18159,N_18385);
or U19169 (N_19169,N_18503,N_18469);
or U19170 (N_19170,N_18385,N_18300);
nand U19171 (N_19171,N_18627,N_18693);
xor U19172 (N_19172,N_18551,N_18271);
xnor U19173 (N_19173,N_18673,N_18565);
and U19174 (N_19174,N_18444,N_18295);
or U19175 (N_19175,N_18412,N_18451);
or U19176 (N_19176,N_18354,N_18617);
xnor U19177 (N_19177,N_18676,N_18557);
xnor U19178 (N_19178,N_18359,N_18370);
and U19179 (N_19179,N_18555,N_18273);
nand U19180 (N_19180,N_18316,N_18622);
nor U19181 (N_19181,N_18540,N_18647);
or U19182 (N_19182,N_18315,N_18600);
nor U19183 (N_19183,N_18727,N_18215);
nor U19184 (N_19184,N_18615,N_18450);
xnor U19185 (N_19185,N_18463,N_18157);
nand U19186 (N_19186,N_18642,N_18585);
nand U19187 (N_19187,N_18472,N_18372);
nor U19188 (N_19188,N_18358,N_18292);
xnor U19189 (N_19189,N_18342,N_18559);
nor U19190 (N_19190,N_18226,N_18725);
nand U19191 (N_19191,N_18128,N_18184);
and U19192 (N_19192,N_18714,N_18520);
nor U19193 (N_19193,N_18322,N_18711);
nand U19194 (N_19194,N_18142,N_18402);
and U19195 (N_19195,N_18719,N_18184);
nand U19196 (N_19196,N_18469,N_18694);
or U19197 (N_19197,N_18596,N_18701);
xnor U19198 (N_19198,N_18403,N_18304);
xor U19199 (N_19199,N_18159,N_18249);
xnor U19200 (N_19200,N_18740,N_18242);
xnor U19201 (N_19201,N_18399,N_18512);
nand U19202 (N_19202,N_18472,N_18432);
or U19203 (N_19203,N_18251,N_18686);
nor U19204 (N_19204,N_18387,N_18225);
nor U19205 (N_19205,N_18206,N_18669);
nor U19206 (N_19206,N_18557,N_18137);
or U19207 (N_19207,N_18253,N_18208);
nand U19208 (N_19208,N_18362,N_18279);
or U19209 (N_19209,N_18201,N_18532);
nor U19210 (N_19210,N_18378,N_18171);
xor U19211 (N_19211,N_18569,N_18434);
or U19212 (N_19212,N_18264,N_18681);
nand U19213 (N_19213,N_18542,N_18575);
nor U19214 (N_19214,N_18131,N_18327);
nand U19215 (N_19215,N_18243,N_18512);
and U19216 (N_19216,N_18370,N_18386);
nor U19217 (N_19217,N_18546,N_18669);
xor U19218 (N_19218,N_18691,N_18163);
and U19219 (N_19219,N_18602,N_18468);
and U19220 (N_19220,N_18356,N_18629);
xor U19221 (N_19221,N_18421,N_18614);
and U19222 (N_19222,N_18611,N_18374);
or U19223 (N_19223,N_18319,N_18633);
or U19224 (N_19224,N_18577,N_18198);
nor U19225 (N_19225,N_18385,N_18157);
nor U19226 (N_19226,N_18624,N_18312);
or U19227 (N_19227,N_18738,N_18647);
xnor U19228 (N_19228,N_18139,N_18725);
and U19229 (N_19229,N_18436,N_18284);
or U19230 (N_19230,N_18312,N_18156);
nor U19231 (N_19231,N_18250,N_18435);
nand U19232 (N_19232,N_18477,N_18356);
nand U19233 (N_19233,N_18167,N_18302);
nor U19234 (N_19234,N_18581,N_18386);
nand U19235 (N_19235,N_18678,N_18181);
and U19236 (N_19236,N_18391,N_18510);
xnor U19237 (N_19237,N_18728,N_18492);
or U19238 (N_19238,N_18255,N_18621);
and U19239 (N_19239,N_18207,N_18445);
nor U19240 (N_19240,N_18492,N_18156);
and U19241 (N_19241,N_18358,N_18175);
nor U19242 (N_19242,N_18421,N_18406);
nand U19243 (N_19243,N_18263,N_18184);
or U19244 (N_19244,N_18427,N_18398);
xnor U19245 (N_19245,N_18187,N_18637);
and U19246 (N_19246,N_18386,N_18518);
nor U19247 (N_19247,N_18330,N_18711);
xnor U19248 (N_19248,N_18191,N_18277);
nor U19249 (N_19249,N_18748,N_18456);
or U19250 (N_19250,N_18188,N_18403);
and U19251 (N_19251,N_18492,N_18418);
nor U19252 (N_19252,N_18399,N_18157);
or U19253 (N_19253,N_18483,N_18199);
nand U19254 (N_19254,N_18207,N_18683);
and U19255 (N_19255,N_18147,N_18745);
or U19256 (N_19256,N_18399,N_18644);
or U19257 (N_19257,N_18436,N_18282);
and U19258 (N_19258,N_18162,N_18211);
nand U19259 (N_19259,N_18655,N_18552);
or U19260 (N_19260,N_18685,N_18260);
and U19261 (N_19261,N_18191,N_18664);
xor U19262 (N_19262,N_18682,N_18510);
xor U19263 (N_19263,N_18719,N_18664);
nor U19264 (N_19264,N_18552,N_18708);
xnor U19265 (N_19265,N_18464,N_18280);
or U19266 (N_19266,N_18281,N_18452);
nor U19267 (N_19267,N_18746,N_18138);
and U19268 (N_19268,N_18387,N_18424);
and U19269 (N_19269,N_18380,N_18665);
nor U19270 (N_19270,N_18376,N_18210);
xor U19271 (N_19271,N_18139,N_18321);
xor U19272 (N_19272,N_18548,N_18699);
nor U19273 (N_19273,N_18453,N_18222);
or U19274 (N_19274,N_18350,N_18409);
and U19275 (N_19275,N_18274,N_18306);
nand U19276 (N_19276,N_18487,N_18350);
and U19277 (N_19277,N_18529,N_18715);
or U19278 (N_19278,N_18585,N_18492);
and U19279 (N_19279,N_18649,N_18310);
or U19280 (N_19280,N_18480,N_18382);
or U19281 (N_19281,N_18496,N_18684);
xor U19282 (N_19282,N_18669,N_18353);
xnor U19283 (N_19283,N_18608,N_18594);
nor U19284 (N_19284,N_18188,N_18361);
xnor U19285 (N_19285,N_18582,N_18541);
or U19286 (N_19286,N_18261,N_18296);
nor U19287 (N_19287,N_18626,N_18146);
xor U19288 (N_19288,N_18260,N_18646);
and U19289 (N_19289,N_18438,N_18743);
or U19290 (N_19290,N_18226,N_18351);
or U19291 (N_19291,N_18601,N_18334);
or U19292 (N_19292,N_18268,N_18143);
xor U19293 (N_19293,N_18139,N_18689);
xor U19294 (N_19294,N_18344,N_18644);
nand U19295 (N_19295,N_18241,N_18696);
nand U19296 (N_19296,N_18229,N_18332);
and U19297 (N_19297,N_18267,N_18644);
nor U19298 (N_19298,N_18233,N_18545);
or U19299 (N_19299,N_18265,N_18135);
nand U19300 (N_19300,N_18163,N_18417);
and U19301 (N_19301,N_18181,N_18661);
and U19302 (N_19302,N_18517,N_18723);
and U19303 (N_19303,N_18558,N_18665);
and U19304 (N_19304,N_18217,N_18153);
xnor U19305 (N_19305,N_18319,N_18738);
nand U19306 (N_19306,N_18242,N_18163);
or U19307 (N_19307,N_18672,N_18151);
and U19308 (N_19308,N_18505,N_18391);
and U19309 (N_19309,N_18552,N_18416);
and U19310 (N_19310,N_18574,N_18434);
nor U19311 (N_19311,N_18281,N_18219);
and U19312 (N_19312,N_18741,N_18679);
nand U19313 (N_19313,N_18370,N_18409);
or U19314 (N_19314,N_18560,N_18567);
nor U19315 (N_19315,N_18351,N_18374);
xnor U19316 (N_19316,N_18259,N_18471);
and U19317 (N_19317,N_18237,N_18150);
nand U19318 (N_19318,N_18569,N_18252);
nand U19319 (N_19319,N_18173,N_18627);
xnor U19320 (N_19320,N_18167,N_18304);
xnor U19321 (N_19321,N_18731,N_18556);
nor U19322 (N_19322,N_18493,N_18486);
or U19323 (N_19323,N_18201,N_18503);
and U19324 (N_19324,N_18283,N_18671);
or U19325 (N_19325,N_18488,N_18317);
nand U19326 (N_19326,N_18243,N_18133);
nand U19327 (N_19327,N_18282,N_18568);
xnor U19328 (N_19328,N_18273,N_18606);
and U19329 (N_19329,N_18151,N_18665);
or U19330 (N_19330,N_18138,N_18287);
nor U19331 (N_19331,N_18284,N_18248);
or U19332 (N_19332,N_18677,N_18538);
or U19333 (N_19333,N_18514,N_18164);
or U19334 (N_19334,N_18517,N_18679);
or U19335 (N_19335,N_18633,N_18623);
nor U19336 (N_19336,N_18642,N_18314);
nor U19337 (N_19337,N_18266,N_18382);
nor U19338 (N_19338,N_18570,N_18376);
xor U19339 (N_19339,N_18180,N_18160);
nand U19340 (N_19340,N_18655,N_18396);
nand U19341 (N_19341,N_18395,N_18235);
xnor U19342 (N_19342,N_18389,N_18729);
or U19343 (N_19343,N_18381,N_18202);
xor U19344 (N_19344,N_18612,N_18749);
and U19345 (N_19345,N_18392,N_18617);
nor U19346 (N_19346,N_18718,N_18507);
or U19347 (N_19347,N_18711,N_18380);
and U19348 (N_19348,N_18225,N_18375);
and U19349 (N_19349,N_18144,N_18506);
and U19350 (N_19350,N_18273,N_18439);
xnor U19351 (N_19351,N_18141,N_18620);
or U19352 (N_19352,N_18621,N_18692);
or U19353 (N_19353,N_18132,N_18373);
or U19354 (N_19354,N_18177,N_18694);
nor U19355 (N_19355,N_18246,N_18648);
nand U19356 (N_19356,N_18391,N_18169);
or U19357 (N_19357,N_18126,N_18180);
nand U19358 (N_19358,N_18489,N_18726);
and U19359 (N_19359,N_18575,N_18199);
xor U19360 (N_19360,N_18233,N_18449);
nand U19361 (N_19361,N_18399,N_18265);
nor U19362 (N_19362,N_18706,N_18658);
xnor U19363 (N_19363,N_18171,N_18571);
and U19364 (N_19364,N_18195,N_18558);
xnor U19365 (N_19365,N_18476,N_18592);
nand U19366 (N_19366,N_18399,N_18152);
and U19367 (N_19367,N_18276,N_18193);
and U19368 (N_19368,N_18398,N_18400);
xor U19369 (N_19369,N_18386,N_18708);
nand U19370 (N_19370,N_18611,N_18636);
and U19371 (N_19371,N_18339,N_18468);
nand U19372 (N_19372,N_18749,N_18146);
and U19373 (N_19373,N_18326,N_18259);
or U19374 (N_19374,N_18351,N_18146);
xnor U19375 (N_19375,N_18915,N_19162);
and U19376 (N_19376,N_18838,N_18911);
xnor U19377 (N_19377,N_19097,N_19102);
nand U19378 (N_19378,N_18951,N_19183);
and U19379 (N_19379,N_19363,N_18789);
or U19380 (N_19380,N_18875,N_18824);
nor U19381 (N_19381,N_19154,N_19141);
nand U19382 (N_19382,N_19130,N_19021);
nand U19383 (N_19383,N_18968,N_18899);
and U19384 (N_19384,N_19266,N_19319);
xnor U19385 (N_19385,N_19028,N_19082);
nor U19386 (N_19386,N_19370,N_18934);
xor U19387 (N_19387,N_19084,N_19253);
nand U19388 (N_19388,N_19177,N_19030);
nor U19389 (N_19389,N_19263,N_18914);
nor U19390 (N_19390,N_19094,N_19346);
nor U19391 (N_19391,N_19205,N_19220);
nand U19392 (N_19392,N_19295,N_18800);
nand U19393 (N_19393,N_19280,N_19077);
nor U19394 (N_19394,N_18909,N_18971);
or U19395 (N_19395,N_19005,N_19190);
nand U19396 (N_19396,N_19039,N_18794);
and U19397 (N_19397,N_19219,N_18771);
xnor U19398 (N_19398,N_19074,N_19336);
xnor U19399 (N_19399,N_19085,N_19257);
and U19400 (N_19400,N_18872,N_18760);
nand U19401 (N_19401,N_18844,N_19080);
nand U19402 (N_19402,N_18969,N_19095);
nand U19403 (N_19403,N_19222,N_19287);
xnor U19404 (N_19404,N_18990,N_18873);
or U19405 (N_19405,N_19309,N_19156);
nor U19406 (N_19406,N_19216,N_18846);
nor U19407 (N_19407,N_18837,N_18750);
xnor U19408 (N_19408,N_19264,N_18821);
or U19409 (N_19409,N_18945,N_19184);
xor U19410 (N_19410,N_19187,N_18881);
nor U19411 (N_19411,N_19099,N_19078);
and U19412 (N_19412,N_18754,N_18799);
nor U19413 (N_19413,N_18977,N_18974);
nand U19414 (N_19414,N_19349,N_18952);
or U19415 (N_19415,N_19040,N_18777);
and U19416 (N_19416,N_18988,N_18765);
and U19417 (N_19417,N_19125,N_19252);
xor U19418 (N_19418,N_19091,N_19152);
or U19419 (N_19419,N_19001,N_18852);
xor U19420 (N_19420,N_19176,N_18785);
nor U19421 (N_19421,N_19246,N_18978);
xor U19422 (N_19422,N_19301,N_18987);
xor U19423 (N_19423,N_18946,N_19019);
or U19424 (N_19424,N_18774,N_19208);
xor U19425 (N_19425,N_18888,N_19150);
xnor U19426 (N_19426,N_18757,N_19004);
nor U19427 (N_19427,N_19120,N_19015);
nand U19428 (N_19428,N_19278,N_19058);
or U19429 (N_19429,N_19075,N_18880);
nor U19430 (N_19430,N_19139,N_19116);
and U19431 (N_19431,N_19013,N_18902);
nor U19432 (N_19432,N_19124,N_19364);
xor U19433 (N_19433,N_19047,N_18903);
nand U19434 (N_19434,N_18885,N_18912);
and U19435 (N_19435,N_18819,N_18829);
xor U19436 (N_19436,N_18869,N_19088);
nor U19437 (N_19437,N_19062,N_19193);
or U19438 (N_19438,N_19274,N_18877);
and U19439 (N_19439,N_18924,N_19332);
or U19440 (N_19440,N_18790,N_18815);
nand U19441 (N_19441,N_19338,N_19329);
nand U19442 (N_19442,N_19248,N_18897);
nand U19443 (N_19443,N_18953,N_18989);
and U19444 (N_19444,N_19344,N_19159);
nand U19445 (N_19445,N_18926,N_19008);
and U19446 (N_19446,N_18857,N_18890);
xnor U19447 (N_19447,N_19136,N_19144);
nor U19448 (N_19448,N_19113,N_18905);
xor U19449 (N_19449,N_18938,N_18893);
xor U19450 (N_19450,N_19290,N_19305);
nor U19451 (N_19451,N_18916,N_18887);
and U19452 (N_19452,N_18768,N_18894);
nand U19453 (N_19453,N_19191,N_19024);
and U19454 (N_19454,N_19054,N_19299);
xor U19455 (N_19455,N_18848,N_18787);
xnor U19456 (N_19456,N_19284,N_18986);
nand U19457 (N_19457,N_19052,N_18830);
and U19458 (N_19458,N_18940,N_18967);
xor U19459 (N_19459,N_19064,N_18854);
or U19460 (N_19460,N_19371,N_19225);
nor U19461 (N_19461,N_19142,N_19237);
and U19462 (N_19462,N_19151,N_18860);
or U19463 (N_19463,N_18878,N_19131);
and U19464 (N_19464,N_18923,N_19149);
nand U19465 (N_19465,N_18944,N_19112);
or U19466 (N_19466,N_19317,N_19166);
xor U19467 (N_19467,N_19209,N_19175);
nor U19468 (N_19468,N_19354,N_19218);
nand U19469 (N_19469,N_19341,N_18751);
nand U19470 (N_19470,N_19111,N_19081);
and U19471 (N_19471,N_19160,N_19357);
nand U19472 (N_19472,N_18983,N_18861);
nor U19473 (N_19473,N_19161,N_19228);
nand U19474 (N_19474,N_18836,N_19022);
xnor U19475 (N_19475,N_19200,N_18845);
nand U19476 (N_19476,N_18985,N_19065);
nand U19477 (N_19477,N_18862,N_18801);
nand U19478 (N_19478,N_19276,N_19206);
xnor U19479 (N_19479,N_19070,N_18831);
nor U19480 (N_19480,N_18866,N_18853);
nand U19481 (N_19481,N_19326,N_19126);
and U19482 (N_19482,N_18805,N_18808);
nand U19483 (N_19483,N_19330,N_19087);
and U19484 (N_19484,N_19163,N_19242);
xor U19485 (N_19485,N_18939,N_19198);
nor U19486 (N_19486,N_19288,N_19251);
and U19487 (N_19487,N_18975,N_18847);
nor U19488 (N_19488,N_18895,N_18889);
and U19489 (N_19489,N_19038,N_18908);
nor U19490 (N_19490,N_19292,N_18965);
xor U19491 (N_19491,N_18904,N_19217);
or U19492 (N_19492,N_18858,N_18758);
nor U19493 (N_19493,N_19259,N_19037);
nor U19494 (N_19494,N_18930,N_19195);
and U19495 (N_19495,N_19034,N_19270);
xor U19496 (N_19496,N_18792,N_19098);
or U19497 (N_19497,N_19173,N_19308);
xor U19498 (N_19498,N_19221,N_19245);
xnor U19499 (N_19499,N_19369,N_19304);
xnor U19500 (N_19500,N_18841,N_18898);
nor U19501 (N_19501,N_19179,N_19289);
nor U19502 (N_19502,N_18892,N_18850);
xnor U19503 (N_19503,N_19046,N_19254);
and U19504 (N_19504,N_19135,N_19048);
or U19505 (N_19505,N_18835,N_19339);
or U19506 (N_19506,N_19045,N_18913);
nor U19507 (N_19507,N_18943,N_19282);
or U19508 (N_19508,N_19026,N_19044);
and U19509 (N_19509,N_18918,N_18851);
xor U19510 (N_19510,N_18999,N_18922);
and U19511 (N_19511,N_19106,N_19324);
and U19512 (N_19512,N_18901,N_19239);
xnor U19513 (N_19513,N_19050,N_18963);
nand U19514 (N_19514,N_19128,N_18991);
nor U19515 (N_19515,N_18883,N_18783);
nor U19516 (N_19516,N_19172,N_18992);
nor U19517 (N_19517,N_19360,N_19114);
nand U19518 (N_19518,N_19223,N_19079);
and U19519 (N_19519,N_19262,N_18871);
nand U19520 (N_19520,N_19189,N_19066);
nand U19521 (N_19521,N_19041,N_18772);
nor U19522 (N_19522,N_19236,N_18752);
and U19523 (N_19523,N_19240,N_19291);
nor U19524 (N_19524,N_19235,N_19132);
xor U19525 (N_19525,N_18766,N_19256);
nand U19526 (N_19526,N_19201,N_18896);
nand U19527 (N_19527,N_19213,N_19063);
and U19528 (N_19528,N_19090,N_19170);
nor U19529 (N_19529,N_19212,N_19303);
or U19530 (N_19530,N_19140,N_19231);
nand U19531 (N_19531,N_19298,N_19232);
and U19532 (N_19532,N_19117,N_19020);
xor U19533 (N_19533,N_19322,N_19007);
and U19534 (N_19534,N_19076,N_18804);
nand U19535 (N_19535,N_19355,N_19023);
xor U19536 (N_19536,N_18755,N_19321);
and U19537 (N_19537,N_18906,N_19277);
and U19538 (N_19538,N_18947,N_19027);
and U19539 (N_19539,N_19169,N_19343);
nor U19540 (N_19540,N_18795,N_18784);
nand U19541 (N_19541,N_18884,N_19096);
xor U19542 (N_19542,N_19347,N_18996);
or U19543 (N_19543,N_18798,N_18811);
nand U19544 (N_19544,N_19294,N_19334);
and U19545 (N_19545,N_19086,N_19153);
and U19546 (N_19546,N_18870,N_18941);
nand U19547 (N_19547,N_18810,N_18782);
nor U19548 (N_19548,N_19059,N_19250);
or U19549 (N_19549,N_19268,N_19311);
and U19550 (N_19550,N_18973,N_19226);
nand U19551 (N_19551,N_19325,N_18833);
xnor U19552 (N_19552,N_19337,N_18959);
and U19553 (N_19553,N_19035,N_18840);
xnor U19554 (N_19554,N_19108,N_19271);
nor U19555 (N_19555,N_19122,N_19313);
or U19556 (N_19556,N_18886,N_19164);
nand U19557 (N_19557,N_18948,N_18781);
nor U19558 (N_19558,N_18865,N_19061);
nor U19559 (N_19559,N_18956,N_18842);
nand U19560 (N_19560,N_18961,N_18917);
and U19561 (N_19561,N_19197,N_19186);
nand U19562 (N_19562,N_19158,N_18976);
nor U19563 (N_19563,N_19211,N_18767);
nor U19564 (N_19564,N_19167,N_18927);
nor U19565 (N_19565,N_19283,N_19127);
nor U19566 (N_19566,N_18809,N_19042);
and U19567 (N_19567,N_19067,N_19143);
or U19568 (N_19568,N_18960,N_18776);
and U19569 (N_19569,N_19243,N_18775);
nand U19570 (N_19570,N_18773,N_19286);
nor U19571 (N_19571,N_19204,N_18962);
and U19572 (N_19572,N_19109,N_18763);
xor U19573 (N_19573,N_19134,N_19014);
and U19574 (N_19574,N_19315,N_18910);
nand U19575 (N_19575,N_19361,N_19255);
nand U19576 (N_19576,N_18882,N_19053);
nor U19577 (N_19577,N_19016,N_18966);
and U19578 (N_19578,N_18957,N_18891);
and U19579 (N_19579,N_19306,N_19003);
nand U19580 (N_19580,N_19351,N_19331);
and U19581 (N_19581,N_19133,N_19168);
xnor U19582 (N_19582,N_19258,N_18788);
nor U19583 (N_19583,N_19055,N_18839);
and U19584 (N_19584,N_19178,N_18949);
nand U19585 (N_19585,N_18753,N_18859);
nor U19586 (N_19586,N_18982,N_18843);
xnor U19587 (N_19587,N_19194,N_18907);
nor U19588 (N_19588,N_18761,N_19210);
nor U19589 (N_19589,N_19146,N_19000);
nand U19590 (N_19590,N_19032,N_18814);
or U19591 (N_19591,N_18812,N_19310);
and U19592 (N_19592,N_19068,N_19374);
xnor U19593 (N_19593,N_19297,N_19368);
xnor U19594 (N_19594,N_18964,N_18867);
and U19595 (N_19595,N_19029,N_18817);
or U19596 (N_19596,N_18942,N_18834);
nor U19597 (N_19597,N_19241,N_18806);
nor U19598 (N_19598,N_19137,N_19018);
xnor U19599 (N_19599,N_18826,N_19275);
xor U19600 (N_19600,N_18925,N_19269);
nor U19601 (N_19601,N_19089,N_18856);
xnor U19602 (N_19602,N_19373,N_18876);
xnor U19603 (N_19603,N_18997,N_19107);
and U19604 (N_19604,N_19011,N_19300);
or U19605 (N_19605,N_19318,N_18769);
or U19606 (N_19606,N_19335,N_18828);
nand U19607 (N_19607,N_18998,N_18984);
or U19608 (N_19608,N_18931,N_18950);
nor U19609 (N_19609,N_19345,N_19267);
nor U19610 (N_19610,N_18921,N_19069);
nor U19611 (N_19611,N_19352,N_19043);
nor U19612 (N_19612,N_18919,N_19006);
nand U19613 (N_19613,N_19157,N_19072);
and U19614 (N_19614,N_19051,N_19350);
xnor U19615 (N_19615,N_19207,N_18900);
xor U19616 (N_19616,N_19180,N_19333);
xor U19617 (N_19617,N_18970,N_19199);
and U19618 (N_19618,N_18929,N_19010);
or U19619 (N_19619,N_18827,N_19312);
or U19620 (N_19620,N_19060,N_19174);
nor U19621 (N_19621,N_19234,N_19049);
xor U19622 (N_19622,N_19323,N_18779);
nand U19623 (N_19623,N_19147,N_18832);
xnor U19624 (N_19624,N_18822,N_18855);
xnor U19625 (N_19625,N_18972,N_18937);
nor U19626 (N_19626,N_19118,N_18823);
and U19627 (N_19627,N_19249,N_19202);
and U19628 (N_19628,N_18994,N_19233);
and U19629 (N_19629,N_19307,N_18825);
nand U19630 (N_19630,N_18879,N_18756);
nand U19631 (N_19631,N_19073,N_19293);
and U19632 (N_19632,N_19009,N_19367);
nor U19633 (N_19633,N_19265,N_19372);
nor U19634 (N_19634,N_19340,N_19012);
nand U19635 (N_19635,N_19229,N_19123);
nand U19636 (N_19636,N_18863,N_19273);
nand U19637 (N_19637,N_18935,N_18802);
xnor U19638 (N_19638,N_18980,N_19171);
or U19639 (N_19639,N_18770,N_19002);
nor U19640 (N_19640,N_18813,N_19031);
and U19641 (N_19641,N_19115,N_18849);
nor U19642 (N_19642,N_19181,N_18796);
nand U19643 (N_19643,N_19272,N_19327);
xor U19644 (N_19644,N_18780,N_19296);
nand U19645 (N_19645,N_18874,N_19025);
nor U19646 (N_19646,N_18762,N_18920);
nor U19647 (N_19647,N_19342,N_18981);
and U19648 (N_19648,N_19056,N_19105);
or U19649 (N_19649,N_18979,N_18868);
nor U19650 (N_19650,N_19036,N_18928);
or U19651 (N_19651,N_19071,N_18793);
nor U19652 (N_19652,N_19185,N_18807);
xnor U19653 (N_19653,N_19366,N_19188);
and U19654 (N_19654,N_19358,N_19033);
nor U19655 (N_19655,N_18820,N_18818);
or U19656 (N_19656,N_18995,N_19328);
nand U19657 (N_19657,N_19314,N_19203);
nor U19658 (N_19658,N_19302,N_19119);
and U19659 (N_19659,N_18958,N_19017);
xnor U19660 (N_19660,N_19148,N_19182);
nor U19661 (N_19661,N_19356,N_18954);
nor U19662 (N_19662,N_19230,N_19103);
nand U19663 (N_19663,N_19238,N_19083);
and U19664 (N_19664,N_19247,N_18816);
xnor U19665 (N_19665,N_18797,N_19165);
nand U19666 (N_19666,N_19281,N_19214);
nand U19667 (N_19667,N_19261,N_19359);
nand U19668 (N_19668,N_18803,N_18764);
or U19669 (N_19669,N_19155,N_19362);
nor U19670 (N_19670,N_18791,N_19353);
nand U19671 (N_19671,N_19320,N_19093);
or U19672 (N_19672,N_19215,N_19196);
nor U19673 (N_19673,N_19192,N_19244);
nand U19674 (N_19674,N_19129,N_18933);
or U19675 (N_19675,N_19145,N_19057);
or U19676 (N_19676,N_18936,N_18993);
and U19677 (N_19677,N_19279,N_19100);
and U19678 (N_19678,N_19104,N_19224);
and U19679 (N_19679,N_18955,N_19121);
and U19680 (N_19680,N_19260,N_18759);
nand U19681 (N_19681,N_19348,N_19227);
and U19682 (N_19682,N_19285,N_19101);
or U19683 (N_19683,N_18786,N_19316);
xnor U19684 (N_19684,N_19138,N_18932);
xor U19685 (N_19685,N_18778,N_19365);
nand U19686 (N_19686,N_19110,N_19092);
or U19687 (N_19687,N_18864,N_18862);
nand U19688 (N_19688,N_19194,N_19330);
nor U19689 (N_19689,N_19185,N_19041);
or U19690 (N_19690,N_19292,N_18780);
nor U19691 (N_19691,N_19331,N_18888);
and U19692 (N_19692,N_18950,N_19191);
nor U19693 (N_19693,N_19084,N_19060);
nand U19694 (N_19694,N_19022,N_19128);
or U19695 (N_19695,N_19279,N_19060);
nor U19696 (N_19696,N_18873,N_19204);
nand U19697 (N_19697,N_19166,N_19327);
nand U19698 (N_19698,N_18791,N_18871);
and U19699 (N_19699,N_19249,N_18750);
and U19700 (N_19700,N_18827,N_18869);
xnor U19701 (N_19701,N_19135,N_19200);
or U19702 (N_19702,N_18893,N_19295);
nand U19703 (N_19703,N_18780,N_19114);
or U19704 (N_19704,N_19082,N_19356);
or U19705 (N_19705,N_19301,N_19077);
or U19706 (N_19706,N_19144,N_18982);
or U19707 (N_19707,N_18765,N_18801);
nand U19708 (N_19708,N_19249,N_18850);
nand U19709 (N_19709,N_19293,N_19106);
nand U19710 (N_19710,N_18771,N_19132);
nand U19711 (N_19711,N_18928,N_19051);
or U19712 (N_19712,N_19369,N_19013);
and U19713 (N_19713,N_19230,N_18981);
or U19714 (N_19714,N_19116,N_18815);
xnor U19715 (N_19715,N_18806,N_19065);
nand U19716 (N_19716,N_19298,N_19216);
and U19717 (N_19717,N_18905,N_18803);
and U19718 (N_19718,N_19319,N_19057);
nor U19719 (N_19719,N_19036,N_19008);
or U19720 (N_19720,N_18812,N_19187);
xnor U19721 (N_19721,N_19036,N_18991);
or U19722 (N_19722,N_19152,N_19315);
nand U19723 (N_19723,N_19092,N_18786);
xnor U19724 (N_19724,N_19094,N_18869);
or U19725 (N_19725,N_19277,N_18788);
xnor U19726 (N_19726,N_19231,N_18758);
xor U19727 (N_19727,N_19098,N_19133);
nor U19728 (N_19728,N_18939,N_18893);
xnor U19729 (N_19729,N_19278,N_18875);
nand U19730 (N_19730,N_19181,N_18941);
nand U19731 (N_19731,N_18986,N_19277);
nor U19732 (N_19732,N_19057,N_18789);
nand U19733 (N_19733,N_19330,N_18967);
nor U19734 (N_19734,N_19355,N_19162);
or U19735 (N_19735,N_19192,N_19084);
or U19736 (N_19736,N_18875,N_18914);
nor U19737 (N_19737,N_18865,N_19213);
nor U19738 (N_19738,N_19210,N_18883);
nand U19739 (N_19739,N_19271,N_18911);
nand U19740 (N_19740,N_19298,N_18956);
nor U19741 (N_19741,N_19071,N_19341);
or U19742 (N_19742,N_19312,N_19342);
xor U19743 (N_19743,N_18985,N_18755);
xor U19744 (N_19744,N_19112,N_18996);
nand U19745 (N_19745,N_18873,N_19078);
xor U19746 (N_19746,N_18868,N_18927);
and U19747 (N_19747,N_18879,N_18991);
xnor U19748 (N_19748,N_19287,N_19343);
and U19749 (N_19749,N_19371,N_19071);
or U19750 (N_19750,N_18754,N_18942);
nor U19751 (N_19751,N_19123,N_18898);
nor U19752 (N_19752,N_19218,N_18758);
nand U19753 (N_19753,N_19060,N_19078);
nand U19754 (N_19754,N_19195,N_19033);
xnor U19755 (N_19755,N_18980,N_18947);
or U19756 (N_19756,N_19253,N_19254);
or U19757 (N_19757,N_18837,N_18855);
nor U19758 (N_19758,N_19343,N_19173);
xnor U19759 (N_19759,N_19222,N_19353);
or U19760 (N_19760,N_18835,N_18876);
and U19761 (N_19761,N_18945,N_18944);
nor U19762 (N_19762,N_19232,N_19188);
or U19763 (N_19763,N_19060,N_19241);
nand U19764 (N_19764,N_19253,N_18990);
xor U19765 (N_19765,N_19237,N_18796);
xnor U19766 (N_19766,N_18840,N_19106);
nor U19767 (N_19767,N_19203,N_18810);
or U19768 (N_19768,N_19359,N_18815);
or U19769 (N_19769,N_19107,N_18914);
or U19770 (N_19770,N_19200,N_19349);
xor U19771 (N_19771,N_19357,N_18970);
and U19772 (N_19772,N_18901,N_18863);
and U19773 (N_19773,N_18836,N_18887);
or U19774 (N_19774,N_18987,N_19242);
and U19775 (N_19775,N_19252,N_19016);
xor U19776 (N_19776,N_18792,N_19156);
nor U19777 (N_19777,N_19320,N_19078);
xor U19778 (N_19778,N_19331,N_19356);
or U19779 (N_19779,N_18955,N_18929);
and U19780 (N_19780,N_18803,N_19180);
and U19781 (N_19781,N_18910,N_19281);
or U19782 (N_19782,N_18838,N_19001);
or U19783 (N_19783,N_18997,N_18947);
nor U19784 (N_19784,N_19219,N_19022);
nor U19785 (N_19785,N_19305,N_19058);
nand U19786 (N_19786,N_18933,N_19163);
and U19787 (N_19787,N_19120,N_19064);
nor U19788 (N_19788,N_19037,N_19324);
and U19789 (N_19789,N_19360,N_19280);
nand U19790 (N_19790,N_19118,N_19169);
nand U19791 (N_19791,N_19355,N_18756);
nand U19792 (N_19792,N_19238,N_19040);
nor U19793 (N_19793,N_19187,N_19200);
xor U19794 (N_19794,N_19150,N_18854);
nor U19795 (N_19795,N_19348,N_19366);
and U19796 (N_19796,N_19083,N_19188);
xnor U19797 (N_19797,N_18943,N_19162);
xnor U19798 (N_19798,N_19315,N_18944);
and U19799 (N_19799,N_19162,N_19124);
or U19800 (N_19800,N_19063,N_18878);
nor U19801 (N_19801,N_18785,N_19081);
nand U19802 (N_19802,N_19306,N_19222);
nor U19803 (N_19803,N_19349,N_18989);
xnor U19804 (N_19804,N_18885,N_19251);
nor U19805 (N_19805,N_19338,N_19090);
xor U19806 (N_19806,N_19055,N_19241);
nor U19807 (N_19807,N_19066,N_19040);
xor U19808 (N_19808,N_18910,N_19134);
nor U19809 (N_19809,N_19130,N_18830);
or U19810 (N_19810,N_18841,N_18882);
nand U19811 (N_19811,N_18781,N_19271);
and U19812 (N_19812,N_18815,N_19282);
xnor U19813 (N_19813,N_19025,N_19196);
nor U19814 (N_19814,N_19235,N_19149);
and U19815 (N_19815,N_18878,N_19044);
nand U19816 (N_19816,N_19159,N_19234);
xnor U19817 (N_19817,N_18780,N_18831);
nor U19818 (N_19818,N_18875,N_19296);
nand U19819 (N_19819,N_19275,N_19104);
or U19820 (N_19820,N_19136,N_19032);
nand U19821 (N_19821,N_19099,N_18750);
and U19822 (N_19822,N_19098,N_19264);
nor U19823 (N_19823,N_19260,N_19096);
nand U19824 (N_19824,N_19105,N_19118);
nor U19825 (N_19825,N_19245,N_19234);
nand U19826 (N_19826,N_18997,N_19198);
or U19827 (N_19827,N_19246,N_18836);
nand U19828 (N_19828,N_19305,N_19060);
and U19829 (N_19829,N_18777,N_19074);
xnor U19830 (N_19830,N_19093,N_18750);
nand U19831 (N_19831,N_19366,N_18840);
xnor U19832 (N_19832,N_19277,N_18843);
nand U19833 (N_19833,N_18842,N_19189);
nand U19834 (N_19834,N_19072,N_19096);
and U19835 (N_19835,N_18775,N_18955);
nor U19836 (N_19836,N_18854,N_19037);
and U19837 (N_19837,N_19041,N_19362);
or U19838 (N_19838,N_18901,N_19129);
or U19839 (N_19839,N_19035,N_19284);
nor U19840 (N_19840,N_18855,N_18782);
and U19841 (N_19841,N_19203,N_18924);
xor U19842 (N_19842,N_19069,N_19001);
or U19843 (N_19843,N_19212,N_19369);
nor U19844 (N_19844,N_19344,N_19235);
xor U19845 (N_19845,N_18960,N_18865);
nand U19846 (N_19846,N_19245,N_19179);
or U19847 (N_19847,N_19324,N_19165);
xnor U19848 (N_19848,N_18941,N_19098);
or U19849 (N_19849,N_18832,N_19008);
nor U19850 (N_19850,N_18800,N_18813);
nor U19851 (N_19851,N_19077,N_19017);
or U19852 (N_19852,N_19184,N_18957);
or U19853 (N_19853,N_19314,N_18796);
xnor U19854 (N_19854,N_18799,N_18969);
or U19855 (N_19855,N_19094,N_18938);
and U19856 (N_19856,N_18997,N_19209);
or U19857 (N_19857,N_19018,N_19356);
xnor U19858 (N_19858,N_19101,N_18848);
xnor U19859 (N_19859,N_18956,N_19040);
xnor U19860 (N_19860,N_18936,N_18916);
nand U19861 (N_19861,N_19133,N_18909);
nand U19862 (N_19862,N_19289,N_18980);
nor U19863 (N_19863,N_18981,N_19256);
and U19864 (N_19864,N_19236,N_18954);
or U19865 (N_19865,N_19340,N_19371);
nor U19866 (N_19866,N_18938,N_18927);
or U19867 (N_19867,N_19288,N_18801);
xor U19868 (N_19868,N_19343,N_18976);
or U19869 (N_19869,N_18843,N_18864);
nand U19870 (N_19870,N_19289,N_19251);
nand U19871 (N_19871,N_18964,N_19212);
xnor U19872 (N_19872,N_18970,N_19295);
and U19873 (N_19873,N_18860,N_19309);
or U19874 (N_19874,N_18930,N_19189);
and U19875 (N_19875,N_19331,N_19277);
xnor U19876 (N_19876,N_19304,N_18957);
nor U19877 (N_19877,N_18789,N_18944);
or U19878 (N_19878,N_19095,N_18847);
and U19879 (N_19879,N_19311,N_18966);
xor U19880 (N_19880,N_19253,N_19270);
nand U19881 (N_19881,N_19337,N_19186);
nand U19882 (N_19882,N_19328,N_18984);
nor U19883 (N_19883,N_19176,N_19301);
nand U19884 (N_19884,N_19289,N_19032);
nor U19885 (N_19885,N_19350,N_19064);
or U19886 (N_19886,N_19021,N_18979);
nor U19887 (N_19887,N_18883,N_19021);
xor U19888 (N_19888,N_19353,N_19304);
nor U19889 (N_19889,N_18857,N_19195);
and U19890 (N_19890,N_19095,N_19148);
nor U19891 (N_19891,N_19126,N_18821);
and U19892 (N_19892,N_19177,N_19245);
nor U19893 (N_19893,N_19296,N_19286);
xnor U19894 (N_19894,N_19004,N_19289);
nand U19895 (N_19895,N_19161,N_19160);
nand U19896 (N_19896,N_19347,N_19131);
xnor U19897 (N_19897,N_19274,N_19236);
nor U19898 (N_19898,N_18963,N_19002);
or U19899 (N_19899,N_18838,N_19249);
nor U19900 (N_19900,N_18780,N_18795);
nor U19901 (N_19901,N_19124,N_18989);
xor U19902 (N_19902,N_19257,N_19154);
nor U19903 (N_19903,N_19272,N_19357);
or U19904 (N_19904,N_19051,N_19183);
xor U19905 (N_19905,N_19354,N_19099);
nor U19906 (N_19906,N_19305,N_19130);
nand U19907 (N_19907,N_19095,N_19314);
nand U19908 (N_19908,N_19221,N_19192);
and U19909 (N_19909,N_18975,N_19204);
xnor U19910 (N_19910,N_19128,N_19155);
nand U19911 (N_19911,N_19098,N_19007);
and U19912 (N_19912,N_18839,N_18872);
or U19913 (N_19913,N_19020,N_18851);
xor U19914 (N_19914,N_19021,N_18976);
xor U19915 (N_19915,N_19074,N_19258);
and U19916 (N_19916,N_19165,N_18966);
and U19917 (N_19917,N_19016,N_19286);
nor U19918 (N_19918,N_18973,N_19037);
and U19919 (N_19919,N_19200,N_18837);
nor U19920 (N_19920,N_19047,N_19230);
and U19921 (N_19921,N_18991,N_18820);
nor U19922 (N_19922,N_19085,N_19328);
and U19923 (N_19923,N_18877,N_18996);
nor U19924 (N_19924,N_18769,N_19103);
xor U19925 (N_19925,N_19108,N_19010);
or U19926 (N_19926,N_18861,N_18844);
nand U19927 (N_19927,N_19351,N_19173);
xor U19928 (N_19928,N_18790,N_18943);
xnor U19929 (N_19929,N_18756,N_19042);
and U19930 (N_19930,N_19288,N_19020);
or U19931 (N_19931,N_19223,N_18932);
or U19932 (N_19932,N_19004,N_19023);
xor U19933 (N_19933,N_19303,N_18757);
and U19934 (N_19934,N_19060,N_19301);
and U19935 (N_19935,N_19006,N_19063);
and U19936 (N_19936,N_18893,N_19272);
nor U19937 (N_19937,N_18807,N_19016);
xor U19938 (N_19938,N_19044,N_18893);
xor U19939 (N_19939,N_18836,N_18877);
xnor U19940 (N_19940,N_19309,N_19088);
xnor U19941 (N_19941,N_19123,N_19114);
xor U19942 (N_19942,N_18753,N_19079);
nand U19943 (N_19943,N_19151,N_18989);
xnor U19944 (N_19944,N_19276,N_19021);
nor U19945 (N_19945,N_18767,N_19075);
nand U19946 (N_19946,N_19124,N_19046);
and U19947 (N_19947,N_18777,N_19316);
nand U19948 (N_19948,N_18755,N_19086);
nor U19949 (N_19949,N_19147,N_18935);
nor U19950 (N_19950,N_18890,N_19162);
xor U19951 (N_19951,N_18917,N_19185);
xnor U19952 (N_19952,N_19097,N_19255);
xnor U19953 (N_19953,N_19009,N_19136);
nor U19954 (N_19954,N_18823,N_19217);
xnor U19955 (N_19955,N_18971,N_18950);
and U19956 (N_19956,N_18992,N_19202);
nand U19957 (N_19957,N_19085,N_18926);
nor U19958 (N_19958,N_19273,N_18881);
xor U19959 (N_19959,N_19347,N_18918);
nand U19960 (N_19960,N_19022,N_19020);
and U19961 (N_19961,N_18825,N_19090);
nor U19962 (N_19962,N_19247,N_19084);
nand U19963 (N_19963,N_18865,N_18853);
or U19964 (N_19964,N_19043,N_19308);
or U19965 (N_19965,N_18924,N_19026);
nand U19966 (N_19966,N_19282,N_19004);
nand U19967 (N_19967,N_18793,N_18812);
or U19968 (N_19968,N_19289,N_19197);
nor U19969 (N_19969,N_19345,N_18811);
xnor U19970 (N_19970,N_19098,N_19010);
or U19971 (N_19971,N_19058,N_18904);
and U19972 (N_19972,N_18925,N_19146);
nand U19973 (N_19973,N_19297,N_19281);
and U19974 (N_19974,N_19246,N_19005);
nand U19975 (N_19975,N_18888,N_19113);
nor U19976 (N_19976,N_19105,N_19239);
xnor U19977 (N_19977,N_18970,N_18861);
xor U19978 (N_19978,N_19110,N_19252);
nand U19979 (N_19979,N_18850,N_19221);
nand U19980 (N_19980,N_18969,N_18811);
xnor U19981 (N_19981,N_18947,N_19055);
nand U19982 (N_19982,N_18785,N_18861);
and U19983 (N_19983,N_18797,N_18828);
xnor U19984 (N_19984,N_19116,N_19066);
or U19985 (N_19985,N_18983,N_18809);
nand U19986 (N_19986,N_18941,N_19359);
nor U19987 (N_19987,N_19270,N_19071);
xor U19988 (N_19988,N_18870,N_18937);
nor U19989 (N_19989,N_19155,N_18948);
nor U19990 (N_19990,N_18756,N_19119);
or U19991 (N_19991,N_19041,N_19299);
or U19992 (N_19992,N_19130,N_18850);
xor U19993 (N_19993,N_18826,N_18837);
or U19994 (N_19994,N_19040,N_18958);
nand U19995 (N_19995,N_18978,N_19057);
nor U19996 (N_19996,N_18767,N_18954);
xnor U19997 (N_19997,N_19350,N_18878);
nand U19998 (N_19998,N_19042,N_18785);
nand U19999 (N_19999,N_19293,N_18790);
and U20000 (N_20000,N_19749,N_19621);
and U20001 (N_20001,N_19495,N_19993);
and U20002 (N_20002,N_19706,N_19766);
nand U20003 (N_20003,N_19574,N_19813);
nand U20004 (N_20004,N_19840,N_19432);
nor U20005 (N_20005,N_19822,N_19549);
and U20006 (N_20006,N_19435,N_19675);
and U20007 (N_20007,N_19577,N_19454);
or U20008 (N_20008,N_19963,N_19415);
nor U20009 (N_20009,N_19836,N_19828);
nand U20010 (N_20010,N_19704,N_19763);
and U20011 (N_20011,N_19928,N_19613);
and U20012 (N_20012,N_19851,N_19666);
nand U20013 (N_20013,N_19392,N_19565);
nor U20014 (N_20014,N_19412,N_19870);
nor U20015 (N_20015,N_19859,N_19992);
nor U20016 (N_20016,N_19714,N_19848);
and U20017 (N_20017,N_19852,N_19531);
xor U20018 (N_20018,N_19806,N_19391);
and U20019 (N_20019,N_19664,N_19610);
and U20020 (N_20020,N_19665,N_19383);
nor U20021 (N_20021,N_19409,N_19983);
nor U20022 (N_20022,N_19834,N_19541);
nand U20023 (N_20023,N_19602,N_19820);
xnor U20024 (N_20024,N_19878,N_19910);
xnor U20025 (N_20025,N_19723,N_19999);
xor U20026 (N_20026,N_19566,N_19635);
and U20027 (N_20027,N_19518,N_19452);
xor U20028 (N_20028,N_19601,N_19396);
xor U20029 (N_20029,N_19428,N_19490);
or U20030 (N_20030,N_19973,N_19379);
xnor U20031 (N_20031,N_19690,N_19743);
and U20032 (N_20032,N_19960,N_19485);
and U20033 (N_20033,N_19819,N_19673);
nand U20034 (N_20034,N_19867,N_19948);
xnor U20035 (N_20035,N_19789,N_19833);
xor U20036 (N_20036,N_19896,N_19536);
or U20037 (N_20037,N_19684,N_19744);
nand U20038 (N_20038,N_19529,N_19865);
and U20039 (N_20039,N_19825,N_19900);
or U20040 (N_20040,N_19886,N_19762);
nor U20041 (N_20041,N_19569,N_19829);
and U20042 (N_20042,N_19755,N_19500);
xnor U20043 (N_20043,N_19423,N_19578);
nor U20044 (N_20044,N_19926,N_19542);
nor U20045 (N_20045,N_19464,N_19547);
nor U20046 (N_20046,N_19861,N_19471);
nor U20047 (N_20047,N_19933,N_19949);
xnor U20048 (N_20048,N_19699,N_19850);
nor U20049 (N_20049,N_19742,N_19639);
nor U20050 (N_20050,N_19571,N_19731);
nor U20051 (N_20051,N_19390,N_19959);
xor U20052 (N_20052,N_19545,N_19971);
or U20053 (N_20053,N_19670,N_19404);
and U20054 (N_20054,N_19652,N_19650);
nor U20055 (N_20055,N_19871,N_19687);
nor U20056 (N_20056,N_19802,N_19539);
nand U20057 (N_20057,N_19440,N_19898);
and U20058 (N_20058,N_19853,N_19698);
nor U20059 (N_20059,N_19930,N_19872);
xor U20060 (N_20060,N_19676,N_19425);
and U20061 (N_20061,N_19672,N_19380);
and U20062 (N_20062,N_19589,N_19663);
or U20063 (N_20063,N_19644,N_19625);
nand U20064 (N_20064,N_19997,N_19645);
nand U20065 (N_20065,N_19551,N_19800);
and U20066 (N_20066,N_19831,N_19609);
nor U20067 (N_20067,N_19512,N_19597);
and U20068 (N_20068,N_19453,N_19430);
or U20069 (N_20069,N_19641,N_19510);
xnor U20070 (N_20070,N_19908,N_19513);
xor U20071 (N_20071,N_19969,N_19702);
nand U20072 (N_20072,N_19481,N_19517);
or U20073 (N_20073,N_19446,N_19901);
or U20074 (N_20074,N_19527,N_19709);
or U20075 (N_20075,N_19592,N_19920);
nor U20076 (N_20076,N_19739,N_19581);
xor U20077 (N_20077,N_19895,N_19932);
and U20078 (N_20078,N_19897,N_19923);
nor U20079 (N_20079,N_19594,N_19951);
or U20080 (N_20080,N_19433,N_19669);
xor U20081 (N_20081,N_19975,N_19907);
and U20082 (N_20082,N_19799,N_19449);
nand U20083 (N_20083,N_19795,N_19462);
nand U20084 (N_20084,N_19942,N_19436);
xnor U20085 (N_20085,N_19576,N_19546);
and U20086 (N_20086,N_19860,N_19842);
nor U20087 (N_20087,N_19407,N_19441);
and U20088 (N_20088,N_19768,N_19747);
or U20089 (N_20089,N_19659,N_19889);
nand U20090 (N_20090,N_19656,N_19382);
nand U20091 (N_20091,N_19522,N_19798);
xor U20092 (N_20092,N_19801,N_19535);
xnor U20093 (N_20093,N_19587,N_19520);
nor U20094 (N_20094,N_19680,N_19816);
and U20095 (N_20095,N_19771,N_19781);
or U20096 (N_20096,N_19695,N_19980);
or U20097 (N_20097,N_19525,N_19403);
xor U20098 (N_20098,N_19721,N_19729);
nand U20099 (N_20099,N_19604,N_19387);
and U20100 (N_20100,N_19437,N_19761);
or U20101 (N_20101,N_19572,N_19470);
and U20102 (N_20102,N_19855,N_19996);
nand U20103 (N_20103,N_19735,N_19679);
nor U20104 (N_20104,N_19655,N_19552);
nand U20105 (N_20105,N_19398,N_19465);
and U20106 (N_20106,N_19710,N_19455);
xnor U20107 (N_20107,N_19778,N_19791);
xnor U20108 (N_20108,N_19994,N_19523);
nor U20109 (N_20109,N_19752,N_19805);
nand U20110 (N_20110,N_19413,N_19906);
nor U20111 (N_20111,N_19422,N_19788);
or U20112 (N_20112,N_19925,N_19748);
nor U20113 (N_20113,N_19628,N_19562);
or U20114 (N_20114,N_19492,N_19692);
and U20115 (N_20115,N_19854,N_19693);
and U20116 (N_20116,N_19651,N_19775);
nand U20117 (N_20117,N_19660,N_19890);
xor U20118 (N_20118,N_19640,N_19899);
nand U20119 (N_20119,N_19489,N_19875);
nor U20120 (N_20120,N_19984,N_19429);
nand U20121 (N_20121,N_19629,N_19620);
nor U20122 (N_20122,N_19649,N_19919);
and U20123 (N_20123,N_19982,N_19796);
xor U20124 (N_20124,N_19480,N_19944);
or U20125 (N_20125,N_19599,N_19705);
or U20126 (N_20126,N_19420,N_19627);
xnor U20127 (N_20127,N_19499,N_19807);
xnor U20128 (N_20128,N_19733,N_19503);
or U20129 (N_20129,N_19892,N_19862);
and U20130 (N_20130,N_19902,N_19881);
xnor U20131 (N_20131,N_19674,N_19956);
xnor U20132 (N_20132,N_19779,N_19866);
xnor U20133 (N_20133,N_19904,N_19616);
xor U20134 (N_20134,N_19397,N_19504);
xor U20135 (N_20135,N_19938,N_19882);
or U20136 (N_20136,N_19548,N_19654);
nand U20137 (N_20137,N_19506,N_19691);
and U20138 (N_20138,N_19626,N_19486);
and U20139 (N_20139,N_19515,N_19786);
or U20140 (N_20140,N_19488,N_19401);
xor U20141 (N_20141,N_19737,N_19814);
nor U20142 (N_20142,N_19792,N_19745);
and U20143 (N_20143,N_19421,N_19939);
or U20144 (N_20144,N_19668,N_19978);
nand U20145 (N_20145,N_19377,N_19718);
nor U20146 (N_20146,N_19957,N_19468);
nand U20147 (N_20147,N_19880,N_19482);
xnor U20148 (N_20148,N_19824,N_19979);
xor U20149 (N_20149,N_19491,N_19917);
or U20150 (N_20150,N_19533,N_19568);
nor U20151 (N_20151,N_19634,N_19911);
nand U20152 (N_20152,N_19456,N_19858);
xor U20153 (N_20153,N_19451,N_19385);
or U20154 (N_20154,N_19757,N_19877);
or U20155 (N_20155,N_19774,N_19765);
or U20156 (N_20156,N_19722,N_19927);
nor U20157 (N_20157,N_19438,N_19484);
nor U20158 (N_20158,N_19958,N_19519);
nand U20159 (N_20159,N_19934,N_19473);
and U20160 (N_20160,N_19740,N_19563);
nand U20161 (N_20161,N_19444,N_19719);
nand U20162 (N_20162,N_19450,N_19399);
xor U20163 (N_20163,N_19493,N_19564);
nand U20164 (N_20164,N_19794,N_19918);
nor U20165 (N_20165,N_19427,N_19479);
nor U20166 (N_20166,N_19402,N_19653);
and U20167 (N_20167,N_19558,N_19947);
or U20168 (N_20168,N_19685,N_19395);
nor U20169 (N_20169,N_19717,N_19914);
and U20170 (N_20170,N_19727,N_19595);
and U20171 (N_20171,N_19478,N_19955);
or U20172 (N_20172,N_19913,N_19746);
nand U20173 (N_20173,N_19393,N_19888);
nor U20174 (N_20174,N_19400,N_19458);
xor U20175 (N_20175,N_19561,N_19724);
or U20176 (N_20176,N_19732,N_19411);
xor U20177 (N_20177,N_19497,N_19476);
nand U20178 (N_20178,N_19869,N_19624);
nor U20179 (N_20179,N_19414,N_19924);
nand U20180 (N_20180,N_19844,N_19553);
nor U20181 (N_20181,N_19784,N_19753);
xor U20182 (N_20182,N_19826,N_19937);
or U20183 (N_20183,N_19758,N_19534);
xor U20184 (N_20184,N_19688,N_19388);
xor U20185 (N_20185,N_19847,N_19637);
or U20186 (N_20186,N_19968,N_19474);
xnor U20187 (N_20187,N_19728,N_19868);
nand U20188 (N_20188,N_19579,N_19459);
and U20189 (N_20189,N_19528,N_19560);
or U20190 (N_20190,N_19642,N_19885);
and U20191 (N_20191,N_19405,N_19600);
or U20192 (N_20192,N_19448,N_19985);
and U20193 (N_20193,N_19821,N_19443);
nor U20194 (N_20194,N_19593,N_19683);
nor U20195 (N_20195,N_19508,N_19950);
and U20196 (N_20196,N_19697,N_19804);
or U20197 (N_20197,N_19583,N_19720);
xor U20198 (N_20198,N_19922,N_19953);
and U20199 (N_20199,N_19661,N_19410);
xnor U20200 (N_20200,N_19418,N_19803);
or U20201 (N_20201,N_19460,N_19416);
or U20202 (N_20202,N_19961,N_19883);
and U20203 (N_20203,N_19967,N_19505);
nor U20204 (N_20204,N_19730,N_19770);
nor U20205 (N_20205,N_19573,N_19823);
xor U20206 (N_20206,N_19544,N_19394);
or U20207 (N_20207,N_19483,N_19894);
xnor U20208 (N_20208,N_19475,N_19671);
and U20209 (N_20209,N_19445,N_19736);
and U20210 (N_20210,N_19667,N_19590);
nand U20211 (N_20211,N_19682,N_19630);
or U20212 (N_20212,N_19707,N_19631);
and U20213 (N_20213,N_19686,N_19694);
or U20214 (N_20214,N_19511,N_19759);
and U20215 (N_20215,N_19972,N_19384);
nor U20216 (N_20216,N_19703,N_19965);
or U20217 (N_20217,N_19431,N_19469);
nand U20218 (N_20218,N_19389,N_19463);
nand U20219 (N_20219,N_19678,N_19606);
nor U20220 (N_20220,N_19905,N_19808);
or U20221 (N_20221,N_19843,N_19550);
and U20222 (N_20222,N_19532,N_19750);
and U20223 (N_20223,N_19810,N_19989);
nand U20224 (N_20224,N_19375,N_19526);
xnor U20225 (N_20225,N_19530,N_19472);
and U20226 (N_20226,N_19509,N_19845);
or U20227 (N_20227,N_19540,N_19677);
or U20228 (N_20228,N_19618,N_19608);
xnor U20229 (N_20229,N_19605,N_19838);
or U20230 (N_20230,N_19945,N_19891);
or U20231 (N_20231,N_19738,N_19514);
nor U20232 (N_20232,N_19818,N_19632);
or U20233 (N_20233,N_19696,N_19507);
nor U20234 (N_20234,N_19700,N_19584);
and U20235 (N_20235,N_19648,N_19936);
and U20236 (N_20236,N_19582,N_19543);
nor U20237 (N_20237,N_19426,N_19619);
nand U20238 (N_20238,N_19931,N_19557);
or U20239 (N_20239,N_19419,N_19811);
nand U20240 (N_20240,N_19466,N_19643);
and U20241 (N_20241,N_19408,N_19974);
and U20242 (N_20242,N_19783,N_19417);
or U20243 (N_20243,N_19596,N_19767);
and U20244 (N_20244,N_19498,N_19467);
xnor U20245 (N_20245,N_19636,N_19494);
or U20246 (N_20246,N_19764,N_19998);
xor U20247 (N_20247,N_19725,N_19785);
or U20248 (N_20248,N_19782,N_19772);
and U20249 (N_20249,N_19903,N_19754);
nand U20250 (N_20250,N_19943,N_19386);
and U20251 (N_20251,N_19457,N_19787);
and U20252 (N_20252,N_19952,N_19991);
nor U20253 (N_20253,N_19777,N_19734);
and U20254 (N_20254,N_19516,N_19887);
and U20255 (N_20255,N_19713,N_19559);
and U20256 (N_20256,N_19567,N_19760);
nor U20257 (N_20257,N_19521,N_19935);
or U20258 (N_20258,N_19555,N_19376);
or U20259 (N_20259,N_19647,N_19580);
nor U20260 (N_20260,N_19585,N_19442);
xor U20261 (N_20261,N_19614,N_19909);
xor U20262 (N_20262,N_19812,N_19815);
xor U20263 (N_20263,N_19929,N_19835);
nand U20264 (N_20264,N_19434,N_19726);
or U20265 (N_20265,N_19538,N_19611);
and U20266 (N_20266,N_19873,N_19406);
and U20267 (N_20267,N_19962,N_19477);
nand U20268 (N_20268,N_19591,N_19708);
and U20269 (N_20269,N_19623,N_19874);
nor U20270 (N_20270,N_19977,N_19741);
xnor U20271 (N_20271,N_19986,N_19837);
and U20272 (N_20272,N_19646,N_19921);
nand U20273 (N_20273,N_19780,N_19612);
or U20274 (N_20274,N_19570,N_19658);
or U20275 (N_20275,N_19940,N_19776);
or U20276 (N_20276,N_19487,N_19439);
or U20277 (N_20277,N_19756,N_19916);
and U20278 (N_20278,N_19424,N_19701);
nand U20279 (N_20279,N_19846,N_19841);
and U20280 (N_20280,N_19378,N_19893);
nand U20281 (N_20281,N_19856,N_19617);
nor U20282 (N_20282,N_19981,N_19751);
nor U20283 (N_20283,N_19461,N_19827);
or U20284 (N_20284,N_19501,N_19502);
and U20285 (N_20285,N_19638,N_19715);
xnor U20286 (N_20286,N_19830,N_19711);
and U20287 (N_20287,N_19954,N_19987);
xor U20288 (N_20288,N_19879,N_19790);
and U20289 (N_20289,N_19716,N_19863);
nand U20290 (N_20290,N_19809,N_19915);
nor U20291 (N_20291,N_19884,N_19615);
or U20292 (N_20292,N_19941,N_19849);
nand U20293 (N_20293,N_19970,N_19817);
or U20294 (N_20294,N_19554,N_19537);
nor U20295 (N_20295,N_19447,N_19598);
nor U20296 (N_20296,N_19496,N_19797);
xor U20297 (N_20297,N_19995,N_19912);
or U20298 (N_20298,N_19681,N_19633);
and U20299 (N_20299,N_19839,N_19657);
or U20300 (N_20300,N_19793,N_19712);
and U20301 (N_20301,N_19662,N_19769);
xnor U20302 (N_20302,N_19556,N_19864);
nor U20303 (N_20303,N_19381,N_19990);
or U20304 (N_20304,N_19575,N_19964);
xor U20305 (N_20305,N_19773,N_19607);
nand U20306 (N_20306,N_19603,N_19857);
or U20307 (N_20307,N_19622,N_19988);
or U20308 (N_20308,N_19976,N_19689);
or U20309 (N_20309,N_19946,N_19832);
and U20310 (N_20310,N_19966,N_19876);
or U20311 (N_20311,N_19588,N_19524);
xor U20312 (N_20312,N_19586,N_19614);
and U20313 (N_20313,N_19668,N_19489);
or U20314 (N_20314,N_19849,N_19406);
xor U20315 (N_20315,N_19767,N_19659);
nor U20316 (N_20316,N_19448,N_19387);
and U20317 (N_20317,N_19732,N_19447);
xnor U20318 (N_20318,N_19668,N_19633);
or U20319 (N_20319,N_19795,N_19415);
nand U20320 (N_20320,N_19766,N_19732);
nand U20321 (N_20321,N_19495,N_19445);
and U20322 (N_20322,N_19984,N_19445);
xnor U20323 (N_20323,N_19586,N_19735);
and U20324 (N_20324,N_19791,N_19735);
nand U20325 (N_20325,N_19858,N_19774);
nor U20326 (N_20326,N_19595,N_19570);
nand U20327 (N_20327,N_19568,N_19567);
xnor U20328 (N_20328,N_19773,N_19674);
nor U20329 (N_20329,N_19599,N_19499);
nor U20330 (N_20330,N_19901,N_19676);
and U20331 (N_20331,N_19951,N_19574);
nor U20332 (N_20332,N_19979,N_19625);
nor U20333 (N_20333,N_19407,N_19513);
or U20334 (N_20334,N_19688,N_19576);
and U20335 (N_20335,N_19802,N_19463);
nand U20336 (N_20336,N_19811,N_19412);
nand U20337 (N_20337,N_19924,N_19969);
nand U20338 (N_20338,N_19780,N_19721);
nor U20339 (N_20339,N_19817,N_19392);
or U20340 (N_20340,N_19420,N_19424);
and U20341 (N_20341,N_19918,N_19382);
and U20342 (N_20342,N_19947,N_19615);
nor U20343 (N_20343,N_19541,N_19931);
and U20344 (N_20344,N_19793,N_19486);
and U20345 (N_20345,N_19729,N_19924);
and U20346 (N_20346,N_19437,N_19681);
xnor U20347 (N_20347,N_19917,N_19881);
nand U20348 (N_20348,N_19707,N_19595);
and U20349 (N_20349,N_19819,N_19801);
nand U20350 (N_20350,N_19512,N_19916);
nor U20351 (N_20351,N_19598,N_19605);
and U20352 (N_20352,N_19918,N_19923);
and U20353 (N_20353,N_19770,N_19715);
nor U20354 (N_20354,N_19924,N_19984);
xnor U20355 (N_20355,N_19754,N_19955);
nand U20356 (N_20356,N_19498,N_19563);
nor U20357 (N_20357,N_19512,N_19579);
xnor U20358 (N_20358,N_19859,N_19655);
xor U20359 (N_20359,N_19951,N_19571);
and U20360 (N_20360,N_19500,N_19932);
and U20361 (N_20361,N_19429,N_19403);
or U20362 (N_20362,N_19658,N_19765);
or U20363 (N_20363,N_19853,N_19908);
and U20364 (N_20364,N_19869,N_19626);
nor U20365 (N_20365,N_19406,N_19973);
xor U20366 (N_20366,N_19658,N_19752);
nand U20367 (N_20367,N_19680,N_19670);
or U20368 (N_20368,N_19589,N_19877);
or U20369 (N_20369,N_19402,N_19511);
xor U20370 (N_20370,N_19490,N_19654);
and U20371 (N_20371,N_19563,N_19807);
nor U20372 (N_20372,N_19889,N_19549);
or U20373 (N_20373,N_19920,N_19864);
nand U20374 (N_20374,N_19844,N_19463);
nand U20375 (N_20375,N_19874,N_19468);
nor U20376 (N_20376,N_19567,N_19660);
nor U20377 (N_20377,N_19379,N_19723);
nor U20378 (N_20378,N_19424,N_19569);
xnor U20379 (N_20379,N_19478,N_19380);
nand U20380 (N_20380,N_19792,N_19615);
xnor U20381 (N_20381,N_19806,N_19781);
or U20382 (N_20382,N_19494,N_19531);
xor U20383 (N_20383,N_19993,N_19695);
or U20384 (N_20384,N_19385,N_19799);
and U20385 (N_20385,N_19520,N_19607);
and U20386 (N_20386,N_19918,N_19606);
and U20387 (N_20387,N_19903,N_19724);
and U20388 (N_20388,N_19693,N_19668);
or U20389 (N_20389,N_19963,N_19881);
xor U20390 (N_20390,N_19486,N_19380);
nor U20391 (N_20391,N_19393,N_19635);
nand U20392 (N_20392,N_19731,N_19660);
nor U20393 (N_20393,N_19900,N_19947);
and U20394 (N_20394,N_19797,N_19400);
or U20395 (N_20395,N_19579,N_19568);
and U20396 (N_20396,N_19456,N_19752);
xnor U20397 (N_20397,N_19477,N_19644);
nand U20398 (N_20398,N_19516,N_19861);
nor U20399 (N_20399,N_19418,N_19511);
nand U20400 (N_20400,N_19412,N_19693);
nand U20401 (N_20401,N_19710,N_19752);
and U20402 (N_20402,N_19602,N_19549);
xnor U20403 (N_20403,N_19610,N_19407);
nor U20404 (N_20404,N_19420,N_19611);
nand U20405 (N_20405,N_19641,N_19923);
nand U20406 (N_20406,N_19520,N_19525);
xor U20407 (N_20407,N_19711,N_19818);
xnor U20408 (N_20408,N_19405,N_19633);
and U20409 (N_20409,N_19829,N_19624);
xor U20410 (N_20410,N_19379,N_19436);
and U20411 (N_20411,N_19569,N_19784);
nor U20412 (N_20412,N_19798,N_19823);
or U20413 (N_20413,N_19706,N_19953);
or U20414 (N_20414,N_19385,N_19855);
xnor U20415 (N_20415,N_19736,N_19641);
and U20416 (N_20416,N_19796,N_19571);
and U20417 (N_20417,N_19376,N_19379);
and U20418 (N_20418,N_19422,N_19892);
nand U20419 (N_20419,N_19717,N_19960);
and U20420 (N_20420,N_19807,N_19591);
nand U20421 (N_20421,N_19707,N_19693);
nor U20422 (N_20422,N_19983,N_19822);
or U20423 (N_20423,N_19416,N_19698);
nor U20424 (N_20424,N_19933,N_19753);
nor U20425 (N_20425,N_19560,N_19376);
nand U20426 (N_20426,N_19917,N_19420);
or U20427 (N_20427,N_19961,N_19375);
and U20428 (N_20428,N_19629,N_19662);
or U20429 (N_20429,N_19889,N_19393);
nand U20430 (N_20430,N_19739,N_19834);
nor U20431 (N_20431,N_19843,N_19393);
xor U20432 (N_20432,N_19779,N_19870);
nand U20433 (N_20433,N_19880,N_19543);
xnor U20434 (N_20434,N_19597,N_19481);
xnor U20435 (N_20435,N_19907,N_19821);
xnor U20436 (N_20436,N_19893,N_19975);
or U20437 (N_20437,N_19815,N_19859);
nand U20438 (N_20438,N_19982,N_19410);
or U20439 (N_20439,N_19733,N_19795);
or U20440 (N_20440,N_19501,N_19544);
and U20441 (N_20441,N_19722,N_19417);
nand U20442 (N_20442,N_19543,N_19851);
nor U20443 (N_20443,N_19706,N_19585);
nand U20444 (N_20444,N_19695,N_19702);
and U20445 (N_20445,N_19708,N_19896);
nand U20446 (N_20446,N_19479,N_19905);
or U20447 (N_20447,N_19673,N_19726);
nand U20448 (N_20448,N_19470,N_19564);
or U20449 (N_20449,N_19661,N_19663);
and U20450 (N_20450,N_19919,N_19749);
and U20451 (N_20451,N_19787,N_19590);
nor U20452 (N_20452,N_19661,N_19759);
and U20453 (N_20453,N_19657,N_19785);
nor U20454 (N_20454,N_19467,N_19524);
or U20455 (N_20455,N_19563,N_19856);
nand U20456 (N_20456,N_19724,N_19501);
nand U20457 (N_20457,N_19671,N_19497);
nor U20458 (N_20458,N_19390,N_19397);
xnor U20459 (N_20459,N_19421,N_19478);
nor U20460 (N_20460,N_19631,N_19792);
nand U20461 (N_20461,N_19563,N_19434);
nor U20462 (N_20462,N_19712,N_19587);
or U20463 (N_20463,N_19995,N_19595);
and U20464 (N_20464,N_19782,N_19548);
and U20465 (N_20465,N_19767,N_19870);
and U20466 (N_20466,N_19433,N_19559);
xnor U20467 (N_20467,N_19577,N_19497);
nor U20468 (N_20468,N_19501,N_19535);
nor U20469 (N_20469,N_19554,N_19876);
xnor U20470 (N_20470,N_19411,N_19947);
xor U20471 (N_20471,N_19705,N_19631);
or U20472 (N_20472,N_19745,N_19630);
nor U20473 (N_20473,N_19787,N_19562);
nand U20474 (N_20474,N_19739,N_19511);
or U20475 (N_20475,N_19523,N_19693);
xor U20476 (N_20476,N_19533,N_19809);
xnor U20477 (N_20477,N_19611,N_19941);
or U20478 (N_20478,N_19866,N_19983);
and U20479 (N_20479,N_19649,N_19686);
nand U20480 (N_20480,N_19592,N_19934);
nand U20481 (N_20481,N_19989,N_19674);
nand U20482 (N_20482,N_19758,N_19847);
xnor U20483 (N_20483,N_19543,N_19611);
xnor U20484 (N_20484,N_19950,N_19670);
or U20485 (N_20485,N_19588,N_19887);
and U20486 (N_20486,N_19793,N_19960);
and U20487 (N_20487,N_19381,N_19766);
nor U20488 (N_20488,N_19627,N_19501);
nand U20489 (N_20489,N_19469,N_19939);
and U20490 (N_20490,N_19942,N_19632);
nand U20491 (N_20491,N_19629,N_19967);
or U20492 (N_20492,N_19866,N_19412);
nand U20493 (N_20493,N_19563,N_19379);
nor U20494 (N_20494,N_19464,N_19920);
or U20495 (N_20495,N_19396,N_19801);
nand U20496 (N_20496,N_19611,N_19749);
nor U20497 (N_20497,N_19604,N_19818);
nor U20498 (N_20498,N_19853,N_19494);
nand U20499 (N_20499,N_19940,N_19793);
and U20500 (N_20500,N_19499,N_19669);
nor U20501 (N_20501,N_19820,N_19827);
nand U20502 (N_20502,N_19827,N_19736);
nor U20503 (N_20503,N_19955,N_19463);
nor U20504 (N_20504,N_19608,N_19541);
nand U20505 (N_20505,N_19833,N_19980);
nand U20506 (N_20506,N_19925,N_19382);
nor U20507 (N_20507,N_19893,N_19648);
and U20508 (N_20508,N_19401,N_19420);
or U20509 (N_20509,N_19834,N_19561);
and U20510 (N_20510,N_19612,N_19624);
or U20511 (N_20511,N_19935,N_19786);
xnor U20512 (N_20512,N_19914,N_19425);
xnor U20513 (N_20513,N_19646,N_19990);
nor U20514 (N_20514,N_19634,N_19713);
or U20515 (N_20515,N_19816,N_19826);
and U20516 (N_20516,N_19778,N_19886);
nor U20517 (N_20517,N_19609,N_19406);
nor U20518 (N_20518,N_19926,N_19467);
or U20519 (N_20519,N_19763,N_19648);
or U20520 (N_20520,N_19586,N_19548);
nand U20521 (N_20521,N_19790,N_19758);
nand U20522 (N_20522,N_19837,N_19916);
xnor U20523 (N_20523,N_19524,N_19683);
nor U20524 (N_20524,N_19446,N_19537);
and U20525 (N_20525,N_19439,N_19842);
or U20526 (N_20526,N_19386,N_19408);
nor U20527 (N_20527,N_19416,N_19666);
xor U20528 (N_20528,N_19686,N_19437);
nand U20529 (N_20529,N_19386,N_19429);
nor U20530 (N_20530,N_19621,N_19686);
nand U20531 (N_20531,N_19942,N_19780);
and U20532 (N_20532,N_19589,N_19781);
and U20533 (N_20533,N_19910,N_19987);
xor U20534 (N_20534,N_19665,N_19596);
nand U20535 (N_20535,N_19559,N_19933);
nand U20536 (N_20536,N_19804,N_19928);
nand U20537 (N_20537,N_19660,N_19424);
nand U20538 (N_20538,N_19801,N_19964);
nor U20539 (N_20539,N_19732,N_19875);
xnor U20540 (N_20540,N_19593,N_19442);
xnor U20541 (N_20541,N_19794,N_19855);
or U20542 (N_20542,N_19806,N_19379);
and U20543 (N_20543,N_19881,N_19827);
or U20544 (N_20544,N_19605,N_19616);
or U20545 (N_20545,N_19754,N_19929);
or U20546 (N_20546,N_19459,N_19928);
or U20547 (N_20547,N_19836,N_19580);
nor U20548 (N_20548,N_19465,N_19803);
or U20549 (N_20549,N_19896,N_19943);
and U20550 (N_20550,N_19886,N_19777);
nor U20551 (N_20551,N_19455,N_19979);
nand U20552 (N_20552,N_19969,N_19833);
nand U20553 (N_20553,N_19931,N_19768);
and U20554 (N_20554,N_19505,N_19587);
or U20555 (N_20555,N_19518,N_19650);
nor U20556 (N_20556,N_19931,N_19503);
and U20557 (N_20557,N_19607,N_19584);
nor U20558 (N_20558,N_19430,N_19693);
and U20559 (N_20559,N_19425,N_19550);
and U20560 (N_20560,N_19522,N_19917);
and U20561 (N_20561,N_19775,N_19824);
and U20562 (N_20562,N_19468,N_19912);
nand U20563 (N_20563,N_19535,N_19377);
and U20564 (N_20564,N_19383,N_19942);
and U20565 (N_20565,N_19848,N_19707);
nor U20566 (N_20566,N_19410,N_19850);
or U20567 (N_20567,N_19438,N_19500);
xor U20568 (N_20568,N_19512,N_19639);
xnor U20569 (N_20569,N_19965,N_19888);
nor U20570 (N_20570,N_19484,N_19791);
nor U20571 (N_20571,N_19659,N_19636);
or U20572 (N_20572,N_19483,N_19575);
and U20573 (N_20573,N_19751,N_19945);
nor U20574 (N_20574,N_19984,N_19553);
and U20575 (N_20575,N_19618,N_19570);
nor U20576 (N_20576,N_19676,N_19423);
and U20577 (N_20577,N_19824,N_19833);
and U20578 (N_20578,N_19865,N_19692);
nor U20579 (N_20579,N_19895,N_19944);
xor U20580 (N_20580,N_19936,N_19625);
and U20581 (N_20581,N_19656,N_19669);
nor U20582 (N_20582,N_19922,N_19507);
nor U20583 (N_20583,N_19609,N_19453);
nor U20584 (N_20584,N_19995,N_19611);
and U20585 (N_20585,N_19407,N_19704);
or U20586 (N_20586,N_19586,N_19978);
xor U20587 (N_20587,N_19930,N_19733);
xnor U20588 (N_20588,N_19861,N_19971);
xnor U20589 (N_20589,N_19500,N_19688);
or U20590 (N_20590,N_19527,N_19712);
xnor U20591 (N_20591,N_19752,N_19811);
xor U20592 (N_20592,N_19923,N_19665);
or U20593 (N_20593,N_19879,N_19815);
and U20594 (N_20594,N_19896,N_19546);
and U20595 (N_20595,N_19589,N_19800);
xnor U20596 (N_20596,N_19494,N_19992);
nor U20597 (N_20597,N_19844,N_19513);
xor U20598 (N_20598,N_19952,N_19550);
or U20599 (N_20599,N_19716,N_19912);
nand U20600 (N_20600,N_19386,N_19498);
nand U20601 (N_20601,N_19953,N_19382);
or U20602 (N_20602,N_19564,N_19376);
nand U20603 (N_20603,N_19923,N_19567);
nand U20604 (N_20604,N_19477,N_19871);
nor U20605 (N_20605,N_19631,N_19855);
or U20606 (N_20606,N_19665,N_19578);
nand U20607 (N_20607,N_19949,N_19854);
nor U20608 (N_20608,N_19879,N_19407);
xnor U20609 (N_20609,N_19984,N_19513);
and U20610 (N_20610,N_19908,N_19382);
xor U20611 (N_20611,N_19743,N_19711);
xnor U20612 (N_20612,N_19848,N_19932);
xnor U20613 (N_20613,N_19927,N_19486);
xor U20614 (N_20614,N_19613,N_19628);
nand U20615 (N_20615,N_19895,N_19409);
nor U20616 (N_20616,N_19666,N_19893);
nor U20617 (N_20617,N_19700,N_19548);
nor U20618 (N_20618,N_19612,N_19420);
xor U20619 (N_20619,N_19805,N_19509);
or U20620 (N_20620,N_19484,N_19565);
xor U20621 (N_20621,N_19872,N_19599);
xor U20622 (N_20622,N_19542,N_19532);
xor U20623 (N_20623,N_19675,N_19819);
nand U20624 (N_20624,N_19652,N_19958);
and U20625 (N_20625,N_20565,N_20623);
or U20626 (N_20626,N_20279,N_20314);
and U20627 (N_20627,N_20494,N_20492);
and U20628 (N_20628,N_20035,N_20557);
xnor U20629 (N_20629,N_20382,N_20520);
and U20630 (N_20630,N_20386,N_20496);
and U20631 (N_20631,N_20242,N_20562);
nand U20632 (N_20632,N_20000,N_20147);
xnor U20633 (N_20633,N_20060,N_20078);
nor U20634 (N_20634,N_20488,N_20402);
or U20635 (N_20635,N_20568,N_20048);
nand U20636 (N_20636,N_20381,N_20175);
and U20637 (N_20637,N_20469,N_20309);
or U20638 (N_20638,N_20094,N_20390);
xor U20639 (N_20639,N_20030,N_20505);
nor U20640 (N_20640,N_20289,N_20512);
nor U20641 (N_20641,N_20401,N_20235);
nand U20642 (N_20642,N_20613,N_20589);
nor U20643 (N_20643,N_20597,N_20383);
or U20644 (N_20644,N_20617,N_20564);
or U20645 (N_20645,N_20145,N_20215);
xnor U20646 (N_20646,N_20362,N_20421);
nand U20647 (N_20647,N_20211,N_20157);
nand U20648 (N_20648,N_20270,N_20409);
xnor U20649 (N_20649,N_20224,N_20546);
xnor U20650 (N_20650,N_20076,N_20218);
xor U20651 (N_20651,N_20277,N_20422);
nand U20652 (N_20652,N_20561,N_20275);
nor U20653 (N_20653,N_20538,N_20184);
xnor U20654 (N_20654,N_20083,N_20418);
and U20655 (N_20655,N_20302,N_20349);
and U20656 (N_20656,N_20149,N_20027);
nand U20657 (N_20657,N_20013,N_20025);
nand U20658 (N_20658,N_20282,N_20273);
nand U20659 (N_20659,N_20438,N_20487);
and U20660 (N_20660,N_20037,N_20519);
or U20661 (N_20661,N_20377,N_20466);
and U20662 (N_20662,N_20011,N_20034);
and U20663 (N_20663,N_20023,N_20042);
and U20664 (N_20664,N_20266,N_20353);
nand U20665 (N_20665,N_20411,N_20357);
xor U20666 (N_20666,N_20222,N_20615);
xor U20667 (N_20667,N_20190,N_20529);
nand U20668 (N_20668,N_20081,N_20572);
nand U20669 (N_20669,N_20533,N_20256);
xnor U20670 (N_20670,N_20513,N_20344);
and U20671 (N_20671,N_20303,N_20293);
xor U20672 (N_20672,N_20053,N_20442);
nor U20673 (N_20673,N_20280,N_20281);
xor U20674 (N_20674,N_20372,N_20603);
nand U20675 (N_20675,N_20290,N_20598);
nand U20676 (N_20676,N_20294,N_20047);
xnor U20677 (N_20677,N_20050,N_20006);
or U20678 (N_20678,N_20130,N_20062);
and U20679 (N_20679,N_20406,N_20521);
xor U20680 (N_20680,N_20111,N_20611);
and U20681 (N_20681,N_20182,N_20503);
or U20682 (N_20682,N_20250,N_20459);
nand U20683 (N_20683,N_20312,N_20549);
nand U20684 (N_20684,N_20423,N_20579);
and U20685 (N_20685,N_20255,N_20236);
xnor U20686 (N_20686,N_20456,N_20345);
xor U20687 (N_20687,N_20371,N_20536);
and U20688 (N_20688,N_20257,N_20246);
xor U20689 (N_20689,N_20159,N_20142);
xor U20690 (N_20690,N_20040,N_20168);
or U20691 (N_20691,N_20074,N_20299);
and U20692 (N_20692,N_20511,N_20051);
nand U20693 (N_20693,N_20419,N_20311);
nand U20694 (N_20694,N_20583,N_20514);
xnor U20695 (N_20695,N_20272,N_20284);
and U20696 (N_20696,N_20465,N_20497);
xor U20697 (N_20697,N_20563,N_20115);
or U20698 (N_20698,N_20096,N_20458);
or U20699 (N_20699,N_20265,N_20249);
and U20700 (N_20700,N_20123,N_20193);
nor U20701 (N_20701,N_20286,N_20378);
nor U20702 (N_20702,N_20283,N_20334);
and U20703 (N_20703,N_20531,N_20443);
xor U20704 (N_20704,N_20140,N_20194);
nand U20705 (N_20705,N_20073,N_20331);
and U20706 (N_20706,N_20204,N_20189);
and U20707 (N_20707,N_20210,N_20535);
and U20708 (N_20708,N_20365,N_20486);
xnor U20709 (N_20709,N_20374,N_20495);
nor U20710 (N_20710,N_20435,N_20044);
nor U20711 (N_20711,N_20305,N_20616);
xnor U20712 (N_20712,N_20354,N_20560);
nor U20713 (N_20713,N_20103,N_20376);
nor U20714 (N_20714,N_20241,N_20446);
or U20715 (N_20715,N_20101,N_20476);
nor U20716 (N_20716,N_20434,N_20315);
nor U20717 (N_20717,N_20306,N_20567);
or U20718 (N_20718,N_20327,N_20346);
xnor U20719 (N_20719,N_20395,N_20231);
xnor U20720 (N_20720,N_20120,N_20069);
nor U20721 (N_20721,N_20500,N_20274);
xor U20722 (N_20722,N_20198,N_20399);
nor U20723 (N_20723,N_20291,N_20018);
xor U20724 (N_20724,N_20163,N_20188);
nand U20725 (N_20725,N_20169,N_20239);
or U20726 (N_20726,N_20424,N_20186);
or U20727 (N_20727,N_20219,N_20439);
and U20728 (N_20728,N_20417,N_20114);
nor U20729 (N_20729,N_20473,N_20475);
nor U20730 (N_20730,N_20226,N_20229);
and U20731 (N_20731,N_20098,N_20252);
and U20732 (N_20732,N_20366,N_20498);
nand U20733 (N_20733,N_20251,N_20178);
nand U20734 (N_20734,N_20179,N_20271);
nand U20735 (N_20735,N_20172,N_20092);
nand U20736 (N_20736,N_20043,N_20574);
xnor U20737 (N_20737,N_20232,N_20367);
nand U20738 (N_20738,N_20126,N_20326);
xnor U20739 (N_20739,N_20217,N_20379);
xnor U20740 (N_20740,N_20065,N_20407);
nor U20741 (N_20741,N_20622,N_20138);
or U20742 (N_20742,N_20287,N_20400);
or U20743 (N_20743,N_20522,N_20079);
and U20744 (N_20744,N_20196,N_20174);
or U20745 (N_20745,N_20032,N_20359);
or U20746 (N_20746,N_20595,N_20405);
and U20747 (N_20747,N_20484,N_20524);
or U20748 (N_20748,N_20454,N_20244);
xnor U20749 (N_20749,N_20097,N_20045);
and U20750 (N_20750,N_20122,N_20223);
xor U20751 (N_20751,N_20152,N_20610);
xor U20752 (N_20752,N_20554,N_20333);
or U20753 (N_20753,N_20391,N_20012);
or U20754 (N_20754,N_20195,N_20398);
or U20755 (N_20755,N_20119,N_20267);
and U20756 (N_20756,N_20599,N_20005);
nor U20757 (N_20757,N_20584,N_20298);
nor U20758 (N_20758,N_20009,N_20516);
or U20759 (N_20759,N_20243,N_20506);
nor U20760 (N_20760,N_20136,N_20363);
or U20761 (N_20761,N_20426,N_20124);
nand U20762 (N_20762,N_20368,N_20033);
nor U20763 (N_20763,N_20090,N_20385);
and U20764 (N_20764,N_20165,N_20001);
xor U20765 (N_20765,N_20141,N_20491);
nand U20766 (N_20766,N_20370,N_20602);
or U20767 (N_20767,N_20324,N_20089);
xnor U20768 (N_20768,N_20453,N_20340);
nand U20769 (N_20769,N_20518,N_20206);
xnor U20770 (N_20770,N_20148,N_20228);
nor U20771 (N_20771,N_20348,N_20343);
nand U20772 (N_20772,N_20416,N_20071);
and U20773 (N_20773,N_20181,N_20620);
nor U20774 (N_20774,N_20430,N_20014);
xnor U20775 (N_20775,N_20067,N_20029);
and U20776 (N_20776,N_20039,N_20091);
nor U20777 (N_20777,N_20003,N_20007);
nor U20778 (N_20778,N_20341,N_20117);
and U20779 (N_20779,N_20307,N_20601);
or U20780 (N_20780,N_20262,N_20133);
and U20781 (N_20781,N_20428,N_20173);
nand U20782 (N_20782,N_20397,N_20555);
nand U20783 (N_20783,N_20057,N_20444);
xnor U20784 (N_20784,N_20110,N_20300);
xnor U20785 (N_20785,N_20461,N_20154);
and U20786 (N_20786,N_20261,N_20104);
nand U20787 (N_20787,N_20143,N_20134);
xnor U20788 (N_20788,N_20537,N_20452);
or U20789 (N_20789,N_20288,N_20156);
nor U20790 (N_20790,N_20129,N_20176);
and U20791 (N_20791,N_20591,N_20054);
nand U20792 (N_20792,N_20216,N_20441);
or U20793 (N_20793,N_20026,N_20509);
and U20794 (N_20794,N_20170,N_20480);
xnor U20795 (N_20795,N_20209,N_20082);
or U20796 (N_20796,N_20541,N_20268);
nor U20797 (N_20797,N_20508,N_20197);
and U20798 (N_20798,N_20118,N_20325);
xnor U20799 (N_20799,N_20607,N_20539);
nor U20800 (N_20800,N_20396,N_20201);
xnor U20801 (N_20801,N_20121,N_20502);
nor U20802 (N_20802,N_20046,N_20455);
nand U20803 (N_20803,N_20301,N_20609);
nand U20804 (N_20804,N_20404,N_20336);
and U20805 (N_20805,N_20478,N_20105);
or U20806 (N_20806,N_20463,N_20113);
xor U20807 (N_20807,N_20087,N_20575);
or U20808 (N_20808,N_20116,N_20576);
xnor U20809 (N_20809,N_20551,N_20493);
xnor U20810 (N_20810,N_20022,N_20167);
and U20811 (N_20811,N_20445,N_20171);
xor U20812 (N_20812,N_20080,N_20304);
xnor U20813 (N_20813,N_20019,N_20581);
and U20814 (N_20814,N_20548,N_20059);
or U20815 (N_20815,N_20479,N_20166);
or U20816 (N_20816,N_20146,N_20127);
nor U20817 (N_20817,N_20225,N_20394);
and U20818 (N_20818,N_20036,N_20319);
or U20819 (N_20819,N_20342,N_20403);
and U20820 (N_20820,N_20483,N_20297);
or U20821 (N_20821,N_20450,N_20004);
xor U20822 (N_20822,N_20112,N_20332);
or U20823 (N_20823,N_20542,N_20618);
nand U20824 (N_20824,N_20544,N_20467);
and U20825 (N_20825,N_20472,N_20164);
or U20826 (N_20826,N_20093,N_20318);
xnor U20827 (N_20827,N_20477,N_20269);
xor U20828 (N_20828,N_20553,N_20585);
or U20829 (N_20829,N_20373,N_20107);
and U20830 (N_20830,N_20144,N_20501);
and U20831 (N_20831,N_20412,N_20109);
or U20832 (N_20832,N_20462,N_20614);
nand U20833 (N_20833,N_20202,N_20180);
nand U20834 (N_20834,N_20214,N_20571);
or U20835 (N_20835,N_20070,N_20183);
nand U20836 (N_20836,N_20350,N_20199);
and U20837 (N_20837,N_20203,N_20056);
nand U20838 (N_20838,N_20260,N_20517);
nand U20839 (N_20839,N_20160,N_20594);
xor U20840 (N_20840,N_20328,N_20532);
xnor U20841 (N_20841,N_20322,N_20507);
and U20842 (N_20842,N_20612,N_20296);
xnor U20843 (N_20843,N_20155,N_20320);
nand U20844 (N_20844,N_20245,N_20052);
and U20845 (N_20845,N_20408,N_20310);
nand U20846 (N_20846,N_20460,N_20570);
and U20847 (N_20847,N_20323,N_20085);
and U20848 (N_20848,N_20084,N_20008);
nand U20849 (N_20849,N_20102,N_20361);
xnor U20850 (N_20850,N_20150,N_20552);
and U20851 (N_20851,N_20375,N_20545);
nand U20852 (N_20852,N_20021,N_20436);
or U20853 (N_20853,N_20464,N_20582);
xnor U20854 (N_20854,N_20528,N_20077);
and U20855 (N_20855,N_20308,N_20414);
nand U20856 (N_20856,N_20125,N_20237);
and U20857 (N_20857,N_20276,N_20578);
nor U20858 (N_20858,N_20468,N_20431);
xor U20859 (N_20859,N_20068,N_20388);
or U20860 (N_20860,N_20471,N_20457);
xnor U20861 (N_20861,N_20410,N_20504);
nand U20862 (N_20862,N_20220,N_20432);
nor U20863 (N_20863,N_20041,N_20187);
and U20864 (N_20864,N_20447,N_20259);
nor U20865 (N_20865,N_20015,N_20017);
or U20866 (N_20866,N_20002,N_20413);
and U20867 (N_20867,N_20254,N_20020);
and U20868 (N_20868,N_20337,N_20534);
or U20869 (N_20869,N_20556,N_20221);
nand U20870 (N_20870,N_20064,N_20470);
or U20871 (N_20871,N_20525,N_20429);
nand U20872 (N_20872,N_20580,N_20352);
nor U20873 (N_20873,N_20619,N_20010);
and U20874 (N_20874,N_20200,N_20527);
or U20875 (N_20875,N_20240,N_20106);
nor U20876 (N_20876,N_20606,N_20285);
nand U20877 (N_20877,N_20387,N_20031);
and U20878 (N_20878,N_20151,N_20449);
nor U20879 (N_20879,N_20347,N_20192);
xor U20880 (N_20880,N_20024,N_20088);
xor U20881 (N_20881,N_20016,N_20061);
nor U20882 (N_20882,N_20356,N_20566);
nand U20883 (N_20883,N_20351,N_20329);
nand U20884 (N_20884,N_20389,N_20437);
and U20885 (N_20885,N_20086,N_20415);
nor U20886 (N_20886,N_20358,N_20588);
nor U20887 (N_20887,N_20230,N_20339);
nand U20888 (N_20888,N_20558,N_20600);
xor U20889 (N_20889,N_20208,N_20392);
nor U20890 (N_20890,N_20569,N_20135);
or U20891 (N_20891,N_20295,N_20063);
or U20892 (N_20892,N_20608,N_20380);
xor U20893 (N_20893,N_20510,N_20132);
nor U20894 (N_20894,N_20604,N_20515);
nand U20895 (N_20895,N_20540,N_20247);
nor U20896 (N_20896,N_20213,N_20605);
or U20897 (N_20897,N_20177,N_20384);
and U20898 (N_20898,N_20587,N_20058);
xnor U20899 (N_20899,N_20253,N_20258);
nor U20900 (N_20900,N_20233,N_20066);
and U20901 (N_20901,N_20212,N_20028);
nand U20902 (N_20902,N_20448,N_20278);
or U20903 (N_20903,N_20590,N_20205);
or U20904 (N_20904,N_20137,N_20523);
nor U20905 (N_20905,N_20543,N_20128);
nand U20906 (N_20906,N_20108,N_20420);
nor U20907 (N_20907,N_20158,N_20248);
xor U20908 (N_20908,N_20313,N_20038);
nor U20909 (N_20909,N_20139,N_20481);
or U20910 (N_20910,N_20234,N_20055);
xnor U20911 (N_20911,N_20474,N_20451);
and U20912 (N_20912,N_20238,N_20049);
and U20913 (N_20913,N_20099,N_20321);
xnor U20914 (N_20914,N_20596,N_20573);
or U20915 (N_20915,N_20316,N_20621);
nor U20916 (N_20916,N_20207,N_20433);
nor U20917 (N_20917,N_20364,N_20162);
xnor U20918 (N_20918,N_20592,N_20369);
nor U20919 (N_20919,N_20292,N_20263);
nor U20920 (N_20920,N_20586,N_20317);
nor U20921 (N_20921,N_20577,N_20355);
and U20922 (N_20922,N_20530,N_20264);
or U20923 (N_20923,N_20338,N_20499);
or U20924 (N_20924,N_20161,N_20335);
or U20925 (N_20925,N_20131,N_20440);
or U20926 (N_20926,N_20559,N_20485);
xor U20927 (N_20927,N_20075,N_20547);
nor U20928 (N_20928,N_20185,N_20095);
xnor U20929 (N_20929,N_20550,N_20624);
nor U20930 (N_20930,N_20490,N_20100);
or U20931 (N_20931,N_20482,N_20526);
xnor U20932 (N_20932,N_20330,N_20360);
and U20933 (N_20933,N_20427,N_20191);
nor U20934 (N_20934,N_20072,N_20489);
and U20935 (N_20935,N_20153,N_20227);
nand U20936 (N_20936,N_20393,N_20425);
nor U20937 (N_20937,N_20593,N_20123);
and U20938 (N_20938,N_20032,N_20241);
nand U20939 (N_20939,N_20376,N_20475);
nor U20940 (N_20940,N_20140,N_20125);
or U20941 (N_20941,N_20365,N_20425);
nand U20942 (N_20942,N_20281,N_20222);
nand U20943 (N_20943,N_20054,N_20490);
or U20944 (N_20944,N_20138,N_20339);
and U20945 (N_20945,N_20210,N_20522);
and U20946 (N_20946,N_20415,N_20576);
xor U20947 (N_20947,N_20104,N_20140);
nor U20948 (N_20948,N_20001,N_20164);
and U20949 (N_20949,N_20524,N_20485);
nor U20950 (N_20950,N_20533,N_20189);
xnor U20951 (N_20951,N_20388,N_20139);
nor U20952 (N_20952,N_20526,N_20575);
or U20953 (N_20953,N_20398,N_20217);
nand U20954 (N_20954,N_20400,N_20525);
nand U20955 (N_20955,N_20444,N_20377);
xnor U20956 (N_20956,N_20479,N_20543);
and U20957 (N_20957,N_20436,N_20530);
and U20958 (N_20958,N_20107,N_20338);
and U20959 (N_20959,N_20457,N_20240);
nand U20960 (N_20960,N_20305,N_20142);
nand U20961 (N_20961,N_20497,N_20070);
xor U20962 (N_20962,N_20166,N_20088);
xor U20963 (N_20963,N_20183,N_20191);
or U20964 (N_20964,N_20503,N_20554);
or U20965 (N_20965,N_20545,N_20423);
and U20966 (N_20966,N_20532,N_20217);
nor U20967 (N_20967,N_20546,N_20171);
xnor U20968 (N_20968,N_20022,N_20079);
xnor U20969 (N_20969,N_20323,N_20269);
and U20970 (N_20970,N_20258,N_20363);
and U20971 (N_20971,N_20277,N_20494);
xnor U20972 (N_20972,N_20119,N_20154);
nor U20973 (N_20973,N_20414,N_20354);
or U20974 (N_20974,N_20096,N_20503);
xor U20975 (N_20975,N_20442,N_20090);
or U20976 (N_20976,N_20449,N_20030);
xnor U20977 (N_20977,N_20516,N_20095);
or U20978 (N_20978,N_20152,N_20483);
nor U20979 (N_20979,N_20046,N_20483);
or U20980 (N_20980,N_20576,N_20374);
or U20981 (N_20981,N_20168,N_20322);
or U20982 (N_20982,N_20185,N_20465);
and U20983 (N_20983,N_20186,N_20003);
nor U20984 (N_20984,N_20368,N_20349);
nand U20985 (N_20985,N_20349,N_20252);
and U20986 (N_20986,N_20119,N_20140);
or U20987 (N_20987,N_20330,N_20320);
nor U20988 (N_20988,N_20120,N_20307);
or U20989 (N_20989,N_20200,N_20019);
nor U20990 (N_20990,N_20462,N_20495);
xnor U20991 (N_20991,N_20428,N_20487);
and U20992 (N_20992,N_20222,N_20216);
xor U20993 (N_20993,N_20323,N_20236);
or U20994 (N_20994,N_20129,N_20016);
and U20995 (N_20995,N_20232,N_20192);
nor U20996 (N_20996,N_20204,N_20070);
or U20997 (N_20997,N_20394,N_20490);
nor U20998 (N_20998,N_20008,N_20372);
xor U20999 (N_20999,N_20178,N_20441);
xor U21000 (N_21000,N_20614,N_20621);
or U21001 (N_21001,N_20420,N_20045);
xnor U21002 (N_21002,N_20227,N_20457);
and U21003 (N_21003,N_20232,N_20187);
nand U21004 (N_21004,N_20039,N_20498);
nand U21005 (N_21005,N_20398,N_20001);
or U21006 (N_21006,N_20296,N_20400);
xor U21007 (N_21007,N_20088,N_20448);
or U21008 (N_21008,N_20571,N_20415);
and U21009 (N_21009,N_20604,N_20467);
nand U21010 (N_21010,N_20227,N_20400);
xor U21011 (N_21011,N_20109,N_20528);
nor U21012 (N_21012,N_20205,N_20394);
nand U21013 (N_21013,N_20332,N_20257);
or U21014 (N_21014,N_20460,N_20018);
nor U21015 (N_21015,N_20132,N_20178);
nand U21016 (N_21016,N_20603,N_20511);
nor U21017 (N_21017,N_20520,N_20559);
xor U21018 (N_21018,N_20478,N_20303);
and U21019 (N_21019,N_20390,N_20097);
xor U21020 (N_21020,N_20213,N_20139);
xor U21021 (N_21021,N_20246,N_20364);
or U21022 (N_21022,N_20404,N_20369);
nor U21023 (N_21023,N_20556,N_20545);
xor U21024 (N_21024,N_20106,N_20562);
nor U21025 (N_21025,N_20381,N_20060);
nand U21026 (N_21026,N_20377,N_20186);
and U21027 (N_21027,N_20058,N_20334);
nor U21028 (N_21028,N_20392,N_20366);
xnor U21029 (N_21029,N_20054,N_20539);
and U21030 (N_21030,N_20421,N_20482);
nor U21031 (N_21031,N_20491,N_20427);
xnor U21032 (N_21032,N_20430,N_20619);
or U21033 (N_21033,N_20579,N_20450);
or U21034 (N_21034,N_20052,N_20419);
or U21035 (N_21035,N_20091,N_20199);
xnor U21036 (N_21036,N_20049,N_20364);
nor U21037 (N_21037,N_20281,N_20438);
xnor U21038 (N_21038,N_20532,N_20401);
nor U21039 (N_21039,N_20415,N_20005);
nand U21040 (N_21040,N_20392,N_20118);
xor U21041 (N_21041,N_20257,N_20548);
nor U21042 (N_21042,N_20506,N_20561);
and U21043 (N_21043,N_20353,N_20309);
nand U21044 (N_21044,N_20620,N_20057);
nand U21045 (N_21045,N_20100,N_20205);
and U21046 (N_21046,N_20260,N_20238);
nand U21047 (N_21047,N_20510,N_20379);
xnor U21048 (N_21048,N_20463,N_20145);
and U21049 (N_21049,N_20539,N_20247);
and U21050 (N_21050,N_20220,N_20407);
nand U21051 (N_21051,N_20614,N_20053);
nand U21052 (N_21052,N_20182,N_20155);
nor U21053 (N_21053,N_20113,N_20470);
nand U21054 (N_21054,N_20194,N_20072);
or U21055 (N_21055,N_20584,N_20193);
or U21056 (N_21056,N_20104,N_20254);
nor U21057 (N_21057,N_20308,N_20606);
nand U21058 (N_21058,N_20624,N_20428);
or U21059 (N_21059,N_20092,N_20162);
and U21060 (N_21060,N_20111,N_20315);
xnor U21061 (N_21061,N_20488,N_20095);
nand U21062 (N_21062,N_20517,N_20581);
nand U21063 (N_21063,N_20320,N_20321);
nor U21064 (N_21064,N_20614,N_20289);
and U21065 (N_21065,N_20469,N_20036);
and U21066 (N_21066,N_20093,N_20495);
and U21067 (N_21067,N_20018,N_20506);
or U21068 (N_21068,N_20463,N_20337);
xor U21069 (N_21069,N_20196,N_20403);
or U21070 (N_21070,N_20555,N_20174);
nor U21071 (N_21071,N_20021,N_20607);
or U21072 (N_21072,N_20233,N_20474);
and U21073 (N_21073,N_20568,N_20533);
xor U21074 (N_21074,N_20084,N_20616);
and U21075 (N_21075,N_20040,N_20039);
nand U21076 (N_21076,N_20170,N_20373);
nor U21077 (N_21077,N_20405,N_20307);
nor U21078 (N_21078,N_20134,N_20114);
xnor U21079 (N_21079,N_20318,N_20326);
and U21080 (N_21080,N_20343,N_20449);
and U21081 (N_21081,N_20116,N_20398);
nor U21082 (N_21082,N_20220,N_20466);
xor U21083 (N_21083,N_20291,N_20470);
and U21084 (N_21084,N_20604,N_20053);
nand U21085 (N_21085,N_20568,N_20303);
nand U21086 (N_21086,N_20093,N_20242);
nor U21087 (N_21087,N_20575,N_20386);
or U21088 (N_21088,N_20303,N_20503);
nand U21089 (N_21089,N_20356,N_20572);
and U21090 (N_21090,N_20464,N_20573);
or U21091 (N_21091,N_20222,N_20165);
and U21092 (N_21092,N_20002,N_20379);
nand U21093 (N_21093,N_20041,N_20368);
or U21094 (N_21094,N_20132,N_20514);
and U21095 (N_21095,N_20607,N_20587);
or U21096 (N_21096,N_20613,N_20263);
and U21097 (N_21097,N_20330,N_20541);
and U21098 (N_21098,N_20610,N_20428);
xnor U21099 (N_21099,N_20188,N_20454);
xor U21100 (N_21100,N_20009,N_20087);
xor U21101 (N_21101,N_20572,N_20327);
and U21102 (N_21102,N_20417,N_20265);
nor U21103 (N_21103,N_20268,N_20107);
or U21104 (N_21104,N_20175,N_20590);
nand U21105 (N_21105,N_20275,N_20463);
xnor U21106 (N_21106,N_20486,N_20229);
nor U21107 (N_21107,N_20157,N_20397);
nor U21108 (N_21108,N_20369,N_20277);
xnor U21109 (N_21109,N_20571,N_20411);
nand U21110 (N_21110,N_20204,N_20581);
xor U21111 (N_21111,N_20498,N_20561);
or U21112 (N_21112,N_20449,N_20559);
or U21113 (N_21113,N_20180,N_20334);
xnor U21114 (N_21114,N_20503,N_20402);
and U21115 (N_21115,N_20219,N_20313);
and U21116 (N_21116,N_20027,N_20474);
nand U21117 (N_21117,N_20589,N_20585);
or U21118 (N_21118,N_20577,N_20108);
xor U21119 (N_21119,N_20596,N_20145);
or U21120 (N_21120,N_20180,N_20384);
nor U21121 (N_21121,N_20111,N_20132);
or U21122 (N_21122,N_20042,N_20594);
nand U21123 (N_21123,N_20358,N_20469);
or U21124 (N_21124,N_20455,N_20227);
nor U21125 (N_21125,N_20433,N_20398);
nor U21126 (N_21126,N_20198,N_20252);
nor U21127 (N_21127,N_20374,N_20472);
nand U21128 (N_21128,N_20445,N_20288);
and U21129 (N_21129,N_20249,N_20474);
nand U21130 (N_21130,N_20276,N_20424);
or U21131 (N_21131,N_20479,N_20183);
and U21132 (N_21132,N_20305,N_20313);
nand U21133 (N_21133,N_20372,N_20112);
or U21134 (N_21134,N_20439,N_20129);
nor U21135 (N_21135,N_20005,N_20397);
or U21136 (N_21136,N_20124,N_20367);
or U21137 (N_21137,N_20277,N_20133);
and U21138 (N_21138,N_20450,N_20390);
nor U21139 (N_21139,N_20516,N_20415);
and U21140 (N_21140,N_20505,N_20594);
or U21141 (N_21141,N_20179,N_20030);
nor U21142 (N_21142,N_20132,N_20528);
and U21143 (N_21143,N_20121,N_20240);
and U21144 (N_21144,N_20285,N_20240);
nand U21145 (N_21145,N_20264,N_20344);
nand U21146 (N_21146,N_20001,N_20307);
and U21147 (N_21147,N_20010,N_20026);
nand U21148 (N_21148,N_20623,N_20562);
or U21149 (N_21149,N_20132,N_20623);
nand U21150 (N_21150,N_20510,N_20453);
or U21151 (N_21151,N_20033,N_20377);
and U21152 (N_21152,N_20218,N_20591);
and U21153 (N_21153,N_20617,N_20582);
or U21154 (N_21154,N_20521,N_20340);
or U21155 (N_21155,N_20406,N_20344);
or U21156 (N_21156,N_20595,N_20502);
or U21157 (N_21157,N_20227,N_20141);
nor U21158 (N_21158,N_20217,N_20593);
xor U21159 (N_21159,N_20390,N_20507);
xnor U21160 (N_21160,N_20177,N_20530);
nor U21161 (N_21161,N_20280,N_20340);
xnor U21162 (N_21162,N_20080,N_20263);
nor U21163 (N_21163,N_20010,N_20055);
or U21164 (N_21164,N_20545,N_20615);
and U21165 (N_21165,N_20204,N_20569);
nor U21166 (N_21166,N_20159,N_20608);
or U21167 (N_21167,N_20328,N_20312);
and U21168 (N_21168,N_20165,N_20139);
xnor U21169 (N_21169,N_20376,N_20026);
xnor U21170 (N_21170,N_20484,N_20612);
or U21171 (N_21171,N_20303,N_20576);
nor U21172 (N_21172,N_20396,N_20001);
xnor U21173 (N_21173,N_20345,N_20415);
and U21174 (N_21174,N_20322,N_20084);
and U21175 (N_21175,N_20606,N_20181);
nand U21176 (N_21176,N_20147,N_20287);
xor U21177 (N_21177,N_20211,N_20505);
or U21178 (N_21178,N_20469,N_20062);
and U21179 (N_21179,N_20202,N_20110);
xnor U21180 (N_21180,N_20060,N_20240);
and U21181 (N_21181,N_20213,N_20495);
nand U21182 (N_21182,N_20354,N_20068);
or U21183 (N_21183,N_20045,N_20022);
or U21184 (N_21184,N_20029,N_20527);
nand U21185 (N_21185,N_20060,N_20135);
xnor U21186 (N_21186,N_20248,N_20121);
or U21187 (N_21187,N_20541,N_20304);
and U21188 (N_21188,N_20437,N_20289);
xnor U21189 (N_21189,N_20240,N_20263);
nand U21190 (N_21190,N_20491,N_20158);
nand U21191 (N_21191,N_20257,N_20091);
and U21192 (N_21192,N_20219,N_20120);
or U21193 (N_21193,N_20226,N_20169);
and U21194 (N_21194,N_20168,N_20109);
nand U21195 (N_21195,N_20229,N_20343);
xor U21196 (N_21196,N_20483,N_20400);
xnor U21197 (N_21197,N_20169,N_20111);
xnor U21198 (N_21198,N_20491,N_20619);
or U21199 (N_21199,N_20103,N_20475);
or U21200 (N_21200,N_20242,N_20380);
and U21201 (N_21201,N_20033,N_20303);
nand U21202 (N_21202,N_20461,N_20495);
and U21203 (N_21203,N_20151,N_20326);
or U21204 (N_21204,N_20573,N_20298);
and U21205 (N_21205,N_20363,N_20133);
and U21206 (N_21206,N_20010,N_20348);
nor U21207 (N_21207,N_20582,N_20564);
xor U21208 (N_21208,N_20338,N_20091);
and U21209 (N_21209,N_20411,N_20399);
nor U21210 (N_21210,N_20411,N_20054);
nand U21211 (N_21211,N_20379,N_20436);
and U21212 (N_21212,N_20417,N_20009);
nor U21213 (N_21213,N_20572,N_20035);
nor U21214 (N_21214,N_20511,N_20418);
xor U21215 (N_21215,N_20620,N_20161);
and U21216 (N_21216,N_20080,N_20029);
nand U21217 (N_21217,N_20136,N_20273);
xnor U21218 (N_21218,N_20124,N_20196);
xor U21219 (N_21219,N_20165,N_20358);
or U21220 (N_21220,N_20319,N_20108);
or U21221 (N_21221,N_20586,N_20557);
xnor U21222 (N_21222,N_20176,N_20291);
xor U21223 (N_21223,N_20622,N_20072);
or U21224 (N_21224,N_20047,N_20477);
xor U21225 (N_21225,N_20347,N_20266);
or U21226 (N_21226,N_20215,N_20388);
and U21227 (N_21227,N_20099,N_20597);
or U21228 (N_21228,N_20533,N_20169);
or U21229 (N_21229,N_20204,N_20618);
nor U21230 (N_21230,N_20415,N_20021);
nor U21231 (N_21231,N_20614,N_20452);
or U21232 (N_21232,N_20369,N_20407);
nand U21233 (N_21233,N_20112,N_20384);
nor U21234 (N_21234,N_20320,N_20553);
xor U21235 (N_21235,N_20089,N_20139);
and U21236 (N_21236,N_20031,N_20140);
nand U21237 (N_21237,N_20168,N_20562);
or U21238 (N_21238,N_20113,N_20102);
and U21239 (N_21239,N_20282,N_20544);
nand U21240 (N_21240,N_20220,N_20043);
xor U21241 (N_21241,N_20153,N_20072);
xor U21242 (N_21242,N_20318,N_20331);
xor U21243 (N_21243,N_20307,N_20280);
nand U21244 (N_21244,N_20250,N_20288);
and U21245 (N_21245,N_20328,N_20001);
nor U21246 (N_21246,N_20103,N_20223);
xnor U21247 (N_21247,N_20017,N_20547);
nand U21248 (N_21248,N_20343,N_20039);
nand U21249 (N_21249,N_20131,N_20139);
or U21250 (N_21250,N_21159,N_21125);
xor U21251 (N_21251,N_20768,N_20826);
nand U21252 (N_21252,N_21141,N_21153);
nor U21253 (N_21253,N_20808,N_21007);
nor U21254 (N_21254,N_21170,N_21012);
nand U21255 (N_21255,N_21149,N_20916);
and U21256 (N_21256,N_20807,N_20968);
or U21257 (N_21257,N_20760,N_20770);
xor U21258 (N_21258,N_21167,N_21232);
and U21259 (N_21259,N_21095,N_20701);
xor U21260 (N_21260,N_21106,N_21092);
nand U21261 (N_21261,N_20816,N_21046);
xor U21262 (N_21262,N_20709,N_20664);
xnor U21263 (N_21263,N_21230,N_20758);
or U21264 (N_21264,N_20980,N_20902);
xnor U21265 (N_21265,N_21113,N_20628);
or U21266 (N_21266,N_20663,N_20836);
and U21267 (N_21267,N_20651,N_20736);
nand U21268 (N_21268,N_20898,N_21104);
and U21269 (N_21269,N_20831,N_20793);
or U21270 (N_21270,N_20756,N_21119);
xnor U21271 (N_21271,N_20914,N_20781);
xor U21272 (N_21272,N_20962,N_20657);
nand U21273 (N_21273,N_21193,N_21004);
xor U21274 (N_21274,N_20650,N_20821);
xor U21275 (N_21275,N_20918,N_21073);
nor U21276 (N_21276,N_20975,N_20994);
and U21277 (N_21277,N_21094,N_21084);
or U21278 (N_21278,N_20668,N_20921);
nand U21279 (N_21279,N_21160,N_21054);
and U21280 (N_21280,N_21057,N_20870);
or U21281 (N_21281,N_21089,N_21195);
and U21282 (N_21282,N_20656,N_21215);
nor U21283 (N_21283,N_20744,N_20800);
nand U21284 (N_21284,N_21152,N_21086);
or U21285 (N_21285,N_20928,N_21174);
nor U21286 (N_21286,N_20762,N_20894);
xnor U21287 (N_21287,N_21117,N_21143);
and U21288 (N_21288,N_21060,N_21044);
nor U21289 (N_21289,N_20697,N_21108);
nand U21290 (N_21290,N_20678,N_20704);
xor U21291 (N_21291,N_21175,N_20645);
or U21292 (N_21292,N_21079,N_20794);
or U21293 (N_21293,N_20765,N_21098);
nor U21294 (N_21294,N_21158,N_20636);
nor U21295 (N_21295,N_21024,N_20661);
nor U21296 (N_21296,N_21136,N_21068);
and U21297 (N_21297,N_21135,N_20630);
nand U21298 (N_21298,N_20908,N_21103);
nor U21299 (N_21299,N_20949,N_20647);
or U21300 (N_21300,N_21243,N_20967);
nand U21301 (N_21301,N_20752,N_20899);
nand U21302 (N_21302,N_20690,N_20728);
xnor U21303 (N_21303,N_20738,N_20990);
nor U21304 (N_21304,N_20845,N_20839);
and U21305 (N_21305,N_20764,N_21091);
xnor U21306 (N_21306,N_21052,N_20635);
xnor U21307 (N_21307,N_20979,N_20820);
xor U21308 (N_21308,N_21006,N_21192);
and U21309 (N_21309,N_20689,N_20667);
and U21310 (N_21310,N_20907,N_21048);
xor U21311 (N_21311,N_21029,N_21178);
xnor U21312 (N_21312,N_20951,N_21019);
xnor U21313 (N_21313,N_21242,N_20776);
or U21314 (N_21314,N_21115,N_21214);
and U21315 (N_21315,N_21154,N_21142);
or U21316 (N_21316,N_21134,N_20833);
or U21317 (N_21317,N_20873,N_21222);
xor U21318 (N_21318,N_21082,N_20988);
xnor U21319 (N_21319,N_21122,N_20745);
nand U21320 (N_21320,N_20790,N_20723);
nand U21321 (N_21321,N_20766,N_21190);
nor U21322 (N_21322,N_20740,N_21072);
nor U21323 (N_21323,N_21055,N_20632);
and U21324 (N_21324,N_20725,N_21123);
xor U21325 (N_21325,N_20885,N_21010);
nor U21326 (N_21326,N_20785,N_21067);
and U21327 (N_21327,N_20981,N_20824);
xor U21328 (N_21328,N_20940,N_21188);
xnor U21329 (N_21329,N_20639,N_21023);
or U21330 (N_21330,N_20755,N_20796);
and U21331 (N_21331,N_21062,N_21191);
xor U21332 (N_21332,N_21241,N_20864);
and U21333 (N_21333,N_21201,N_20933);
xor U21334 (N_21334,N_21020,N_20685);
xnor U21335 (N_21335,N_20695,N_20976);
nand U21336 (N_21336,N_20754,N_20943);
nor U21337 (N_21337,N_21231,N_20669);
nand U21338 (N_21338,N_20901,N_21164);
or U21339 (N_21339,N_20903,N_20735);
nor U21340 (N_21340,N_21220,N_20900);
nor U21341 (N_21341,N_20855,N_20835);
nor U21342 (N_21342,N_20642,N_20978);
or U21343 (N_21343,N_20970,N_20662);
and U21344 (N_21344,N_21051,N_20658);
and U21345 (N_21345,N_20998,N_21172);
nand U21346 (N_21346,N_20782,N_21083);
and U21347 (N_21347,N_20818,N_20799);
nor U21348 (N_21348,N_20684,N_20959);
nand U21349 (N_21349,N_20761,N_20784);
nand U21350 (N_21350,N_20640,N_20786);
xnor U21351 (N_21351,N_20787,N_20643);
xor U21352 (N_21352,N_20986,N_20737);
nand U21353 (N_21353,N_21173,N_20625);
nor U21354 (N_21354,N_20960,N_20847);
or U21355 (N_21355,N_21041,N_20763);
xnor U21356 (N_21356,N_20806,N_20712);
nor U21357 (N_21357,N_20869,N_20671);
or U21358 (N_21358,N_20665,N_20673);
or U21359 (N_21359,N_21026,N_20983);
nand U21360 (N_21360,N_20846,N_20891);
or U21361 (N_21361,N_20823,N_21209);
nand U21362 (N_21362,N_20925,N_21197);
nand U21363 (N_21363,N_20681,N_20795);
xor U21364 (N_21364,N_21144,N_20773);
nor U21365 (N_21365,N_21075,N_20931);
nor U21366 (N_21366,N_20880,N_20775);
nor U21367 (N_21367,N_20742,N_21227);
and U21368 (N_21368,N_21003,N_21226);
and U21369 (N_21369,N_20841,N_20734);
and U21370 (N_21370,N_20827,N_21116);
nor U21371 (N_21371,N_20686,N_21240);
nand U21372 (N_21372,N_21169,N_21070);
nor U21373 (N_21373,N_20683,N_20759);
nor U21374 (N_21374,N_21049,N_21210);
nand U21375 (N_21375,N_20927,N_21182);
nor U21376 (N_21376,N_21071,N_20797);
and U21377 (N_21377,N_20739,N_21247);
or U21378 (N_21378,N_20929,N_21080);
xor U21379 (N_21379,N_21147,N_21000);
nand U21380 (N_21380,N_20666,N_21223);
or U21381 (N_21381,N_21235,N_21196);
or U21382 (N_21382,N_20741,N_20874);
xor U21383 (N_21383,N_21107,N_20857);
xnor U21384 (N_21384,N_21217,N_21176);
xor U21385 (N_21385,N_20655,N_20912);
xor U21386 (N_21386,N_20850,N_20714);
or U21387 (N_21387,N_20953,N_20715);
and U21388 (N_21388,N_20868,N_21179);
xor U21389 (N_21389,N_21030,N_20886);
and U21390 (N_21390,N_21138,N_21034);
and U21391 (N_21391,N_20811,N_20915);
xor U21392 (N_21392,N_20746,N_21213);
nand U21393 (N_21393,N_20682,N_21148);
xor U21394 (N_21394,N_20644,N_20677);
xor U21395 (N_21395,N_21180,N_20838);
or U21396 (N_21396,N_20629,N_21132);
xor U21397 (N_21397,N_21001,N_20822);
or U21398 (N_21398,N_20649,N_21245);
xor U21399 (N_21399,N_20828,N_20863);
nand U21400 (N_21400,N_20637,N_20711);
and U21401 (N_21401,N_21163,N_20906);
or U21402 (N_21402,N_21037,N_20798);
nor U21403 (N_21403,N_21111,N_20948);
nor U21404 (N_21404,N_21014,N_21165);
xnor U21405 (N_21405,N_20930,N_20946);
nand U21406 (N_21406,N_21043,N_21090);
xnor U21407 (N_21407,N_20887,N_20965);
nor U21408 (N_21408,N_20952,N_21109);
nand U21409 (N_21409,N_21121,N_20893);
nand U21410 (N_21410,N_20923,N_21127);
nor U21411 (N_21411,N_20802,N_20654);
nor U21412 (N_21412,N_21047,N_20634);
nor U21413 (N_21413,N_21225,N_21204);
and U21414 (N_21414,N_21038,N_21033);
and U21415 (N_21415,N_20939,N_20913);
xnor U21416 (N_21416,N_21237,N_21088);
xnor U21417 (N_21417,N_20837,N_21128);
or U21418 (N_21418,N_21234,N_21015);
nand U21419 (N_21419,N_21099,N_20973);
nor U21420 (N_21420,N_21157,N_20638);
nand U21421 (N_21421,N_20692,N_20890);
xnor U21422 (N_21422,N_20883,N_21228);
and U21423 (N_21423,N_21236,N_21074);
and U21424 (N_21424,N_20733,N_20710);
nand U21425 (N_21425,N_20767,N_21040);
or U21426 (N_21426,N_20964,N_20875);
nor U21427 (N_21427,N_21207,N_20920);
or U21428 (N_21428,N_21077,N_21112);
or U21429 (N_21429,N_21124,N_21239);
nor U21430 (N_21430,N_20693,N_20865);
nand U21431 (N_21431,N_20722,N_20956);
nand U21432 (N_21432,N_20972,N_20878);
nand U21433 (N_21433,N_21065,N_20653);
and U21434 (N_21434,N_20945,N_21181);
and U21435 (N_21435,N_20926,N_21013);
xor U21436 (N_21436,N_21168,N_21246);
or U21437 (N_21437,N_21059,N_20985);
or U21438 (N_21438,N_21200,N_20788);
nand U21439 (N_21439,N_21146,N_20705);
and U21440 (N_21440,N_21221,N_21139);
xnor U21441 (N_21441,N_20852,N_21161);
and U21442 (N_21442,N_20702,N_20969);
or U21443 (N_21443,N_20717,N_20932);
and U21444 (N_21444,N_20812,N_20860);
xor U21445 (N_21445,N_21058,N_21177);
nor U21446 (N_21446,N_20955,N_21025);
xnor U21447 (N_21447,N_20996,N_20938);
nand U21448 (N_21448,N_20861,N_21205);
nor U21449 (N_21449,N_20732,N_20958);
and U21450 (N_21450,N_20751,N_20957);
or U21451 (N_21451,N_21027,N_21150);
nor U21452 (N_21452,N_20849,N_21118);
xor U21453 (N_21453,N_20687,N_20753);
and U21454 (N_21454,N_21005,N_20747);
nor U21455 (N_21455,N_20844,N_20699);
xor U21456 (N_21456,N_21017,N_21224);
nor U21457 (N_21457,N_21145,N_21216);
or U21458 (N_21458,N_20774,N_21249);
xnor U21459 (N_21459,N_20631,N_20727);
or U21460 (N_21460,N_20905,N_21096);
xor U21461 (N_21461,N_20748,N_20924);
nand U21462 (N_21462,N_20783,N_20789);
nor U21463 (N_21463,N_20877,N_20721);
or U21464 (N_21464,N_20867,N_20809);
or U21465 (N_21465,N_21140,N_20743);
nand U21466 (N_21466,N_21061,N_21032);
nand U21467 (N_21467,N_20935,N_20872);
nor U21468 (N_21468,N_20713,N_21035);
nand U21469 (N_21469,N_20676,N_20659);
nor U21470 (N_21470,N_20853,N_20791);
nand U21471 (N_21471,N_20862,N_20729);
xnor U21472 (N_21472,N_20724,N_20750);
or U21473 (N_21473,N_20817,N_20904);
and U21474 (N_21474,N_21187,N_21101);
nor U21475 (N_21475,N_20819,N_21211);
xor U21476 (N_21476,N_20660,N_21248);
nand U21477 (N_21477,N_20897,N_21039);
and U21478 (N_21478,N_20779,N_21053);
nor U21479 (N_21479,N_20999,N_20749);
xor U21480 (N_21480,N_21100,N_21130);
nor U21481 (N_21481,N_21137,N_21042);
nor U21482 (N_21482,N_20730,N_21131);
and U21483 (N_21483,N_20830,N_20731);
or U21484 (N_21484,N_20672,N_20936);
and U21485 (N_21485,N_20881,N_20834);
or U21486 (N_21486,N_20706,N_20718);
nor U21487 (N_21487,N_20832,N_20719);
xor U21488 (N_21488,N_20984,N_21156);
xnor U21489 (N_21489,N_20700,N_20679);
xnor U21490 (N_21490,N_21120,N_21208);
and U21491 (N_21491,N_20696,N_20792);
or U21492 (N_21492,N_20648,N_20757);
xnor U21493 (N_21493,N_21036,N_20895);
nor U21494 (N_21494,N_21206,N_21097);
or U21495 (N_21495,N_20982,N_20726);
nor U21496 (N_21496,N_20910,N_20825);
xnor U21497 (N_21497,N_20934,N_21218);
nand U21498 (N_21498,N_20829,N_20974);
nand U21499 (N_21499,N_20771,N_21009);
nor U21500 (N_21500,N_21110,N_20871);
nor U21501 (N_21501,N_21028,N_21008);
and U21502 (N_21502,N_20892,N_21114);
and U21503 (N_21503,N_20843,N_20815);
xor U21504 (N_21504,N_20992,N_20889);
nor U21505 (N_21505,N_20641,N_20987);
nand U21506 (N_21506,N_21078,N_21018);
nand U21507 (N_21507,N_21063,N_20778);
and U21508 (N_21508,N_21244,N_20777);
nor U21509 (N_21509,N_20993,N_20882);
xor U21510 (N_21510,N_20810,N_20944);
or U21511 (N_21511,N_21021,N_21087);
nor U21512 (N_21512,N_20626,N_20694);
or U21513 (N_21513,N_20814,N_20674);
nor U21514 (N_21514,N_20848,N_20698);
xor U21515 (N_21515,N_21011,N_21186);
nor U21516 (N_21516,N_20801,N_20971);
nand U21517 (N_21517,N_21064,N_20896);
xor U21518 (N_21518,N_20917,N_20627);
or U21519 (N_21519,N_21155,N_21002);
xor U21520 (N_21520,N_20937,N_20888);
or U21521 (N_21521,N_20991,N_21050);
nor U21522 (N_21522,N_21162,N_20966);
and U21523 (N_21523,N_21133,N_21229);
nor U21524 (N_21524,N_21102,N_20652);
xor U21525 (N_21525,N_20909,N_20911);
xor U21526 (N_21526,N_20997,N_21238);
xor U21527 (N_21527,N_20805,N_20720);
nand U21528 (N_21528,N_20977,N_21184);
xnor U21529 (N_21529,N_21056,N_20942);
or U21530 (N_21530,N_20842,N_20866);
xor U21531 (N_21531,N_20859,N_20840);
nor U21532 (N_21532,N_21129,N_20961);
or U21533 (N_21533,N_20633,N_20803);
xor U21534 (N_21534,N_20922,N_20769);
and U21535 (N_21535,N_21203,N_20691);
nand U21536 (N_21536,N_20646,N_20675);
or U21537 (N_21537,N_21045,N_21151);
xnor U21538 (N_21538,N_20879,N_21031);
xor U21539 (N_21539,N_20919,N_21022);
or U21540 (N_21540,N_20950,N_21171);
xor U21541 (N_21541,N_21198,N_21066);
or U21542 (N_21542,N_21166,N_20851);
or U21543 (N_21543,N_20941,N_21126);
and U21544 (N_21544,N_21016,N_20884);
nand U21545 (N_21545,N_21076,N_20813);
nor U21546 (N_21546,N_21081,N_20772);
or U21547 (N_21547,N_20780,N_20708);
or U21548 (N_21548,N_20670,N_20954);
nand U21549 (N_21549,N_21212,N_20703);
xnor U21550 (N_21550,N_20854,N_20989);
nor U21551 (N_21551,N_20856,N_20680);
and U21552 (N_21552,N_21105,N_21219);
or U21553 (N_21553,N_20947,N_20688);
or U21554 (N_21554,N_21185,N_21233);
or U21555 (N_21555,N_20963,N_21085);
xor U21556 (N_21556,N_20876,N_20995);
nor U21557 (N_21557,N_20804,N_21199);
xor U21558 (N_21558,N_21093,N_21202);
or U21559 (N_21559,N_21189,N_20707);
nor U21560 (N_21560,N_21183,N_21069);
xnor U21561 (N_21561,N_20716,N_20858);
nor U21562 (N_21562,N_21194,N_21126);
and U21563 (N_21563,N_21140,N_21043);
nand U21564 (N_21564,N_20692,N_21059);
nor U21565 (N_21565,N_20720,N_21211);
xnor U21566 (N_21566,N_21022,N_21237);
and U21567 (N_21567,N_21220,N_20857);
or U21568 (N_21568,N_21147,N_20832);
or U21569 (N_21569,N_21108,N_20626);
and U21570 (N_21570,N_21086,N_20655);
xnor U21571 (N_21571,N_21165,N_20713);
xnor U21572 (N_21572,N_21157,N_21122);
nor U21573 (N_21573,N_20758,N_20855);
nor U21574 (N_21574,N_21194,N_20953);
xnor U21575 (N_21575,N_20781,N_21113);
nor U21576 (N_21576,N_20660,N_20874);
nor U21577 (N_21577,N_20868,N_20653);
or U21578 (N_21578,N_20870,N_20853);
or U21579 (N_21579,N_21085,N_20818);
nand U21580 (N_21580,N_21028,N_21079);
and U21581 (N_21581,N_20750,N_21072);
nor U21582 (N_21582,N_20776,N_20873);
or U21583 (N_21583,N_21094,N_21134);
xnor U21584 (N_21584,N_20789,N_21152);
or U21585 (N_21585,N_20792,N_20732);
nor U21586 (N_21586,N_21033,N_21084);
or U21587 (N_21587,N_20998,N_20749);
xor U21588 (N_21588,N_21187,N_21040);
nand U21589 (N_21589,N_20996,N_21047);
xor U21590 (N_21590,N_21221,N_20909);
or U21591 (N_21591,N_20691,N_20827);
xor U21592 (N_21592,N_20938,N_20811);
or U21593 (N_21593,N_21034,N_20661);
xnor U21594 (N_21594,N_21031,N_20842);
nand U21595 (N_21595,N_20913,N_20994);
nand U21596 (N_21596,N_20953,N_20977);
xor U21597 (N_21597,N_20897,N_20681);
nor U21598 (N_21598,N_20840,N_20829);
nand U21599 (N_21599,N_20656,N_20752);
and U21600 (N_21600,N_21196,N_21009);
nor U21601 (N_21601,N_21167,N_20803);
or U21602 (N_21602,N_21042,N_20625);
and U21603 (N_21603,N_21010,N_20759);
and U21604 (N_21604,N_20705,N_20839);
and U21605 (N_21605,N_21230,N_21147);
nand U21606 (N_21606,N_20790,N_21221);
and U21607 (N_21607,N_21067,N_20724);
nor U21608 (N_21608,N_20679,N_20772);
xor U21609 (N_21609,N_20840,N_20753);
and U21610 (N_21610,N_20673,N_21205);
xor U21611 (N_21611,N_20888,N_20732);
nor U21612 (N_21612,N_21137,N_20891);
xor U21613 (N_21613,N_20731,N_20709);
nor U21614 (N_21614,N_20899,N_20941);
and U21615 (N_21615,N_21189,N_21079);
and U21616 (N_21616,N_20881,N_20759);
xor U21617 (N_21617,N_20987,N_21117);
nand U21618 (N_21618,N_20834,N_21131);
or U21619 (N_21619,N_20700,N_20739);
or U21620 (N_21620,N_20708,N_21048);
nand U21621 (N_21621,N_20833,N_20835);
xnor U21622 (N_21622,N_20769,N_20904);
or U21623 (N_21623,N_20749,N_20896);
nor U21624 (N_21624,N_20693,N_20732);
or U21625 (N_21625,N_21091,N_21166);
xor U21626 (N_21626,N_21048,N_21116);
nor U21627 (N_21627,N_20818,N_20732);
nand U21628 (N_21628,N_21103,N_20905);
nor U21629 (N_21629,N_20806,N_21171);
nor U21630 (N_21630,N_20783,N_20722);
and U21631 (N_21631,N_20896,N_21042);
and U21632 (N_21632,N_20628,N_20690);
xnor U21633 (N_21633,N_21236,N_21094);
xor U21634 (N_21634,N_20836,N_21023);
xnor U21635 (N_21635,N_21202,N_20971);
and U21636 (N_21636,N_20995,N_20959);
nor U21637 (N_21637,N_20693,N_20909);
nor U21638 (N_21638,N_21150,N_20907);
and U21639 (N_21639,N_21077,N_21006);
nand U21640 (N_21640,N_21175,N_20644);
and U21641 (N_21641,N_21173,N_20749);
or U21642 (N_21642,N_20985,N_21043);
nor U21643 (N_21643,N_20654,N_20702);
or U21644 (N_21644,N_21120,N_20708);
nor U21645 (N_21645,N_21156,N_20929);
xor U21646 (N_21646,N_20972,N_21015);
or U21647 (N_21647,N_21000,N_20688);
nand U21648 (N_21648,N_21198,N_20672);
nor U21649 (N_21649,N_20995,N_20764);
nor U21650 (N_21650,N_21025,N_20968);
and U21651 (N_21651,N_21234,N_20793);
or U21652 (N_21652,N_21011,N_21188);
nand U21653 (N_21653,N_21121,N_20999);
xor U21654 (N_21654,N_21007,N_20916);
xor U21655 (N_21655,N_21148,N_20818);
xor U21656 (N_21656,N_21140,N_20928);
or U21657 (N_21657,N_20954,N_20686);
xor U21658 (N_21658,N_20716,N_20916);
and U21659 (N_21659,N_20791,N_21162);
nor U21660 (N_21660,N_20992,N_21248);
or U21661 (N_21661,N_20880,N_20709);
nand U21662 (N_21662,N_21033,N_21081);
or U21663 (N_21663,N_20970,N_20692);
nand U21664 (N_21664,N_21025,N_20668);
nor U21665 (N_21665,N_21197,N_21019);
and U21666 (N_21666,N_21214,N_20933);
xnor U21667 (N_21667,N_20676,N_20989);
nor U21668 (N_21668,N_21223,N_21082);
nor U21669 (N_21669,N_20710,N_21111);
and U21670 (N_21670,N_20958,N_20863);
xor U21671 (N_21671,N_20982,N_21137);
nor U21672 (N_21672,N_20800,N_21234);
nor U21673 (N_21673,N_20894,N_20766);
nand U21674 (N_21674,N_21107,N_20740);
and U21675 (N_21675,N_20927,N_20763);
xnor U21676 (N_21676,N_20788,N_20638);
nand U21677 (N_21677,N_21111,N_21225);
or U21678 (N_21678,N_21171,N_21054);
or U21679 (N_21679,N_21148,N_20901);
nor U21680 (N_21680,N_20772,N_21073);
or U21681 (N_21681,N_20894,N_21094);
and U21682 (N_21682,N_21113,N_20726);
xnor U21683 (N_21683,N_20828,N_20967);
nor U21684 (N_21684,N_21000,N_21012);
xor U21685 (N_21685,N_20834,N_20890);
and U21686 (N_21686,N_20883,N_20697);
nor U21687 (N_21687,N_20851,N_21156);
xor U21688 (N_21688,N_21033,N_20863);
or U21689 (N_21689,N_21107,N_21085);
nand U21690 (N_21690,N_21136,N_21003);
nand U21691 (N_21691,N_21162,N_20935);
or U21692 (N_21692,N_20894,N_20909);
xor U21693 (N_21693,N_20944,N_21044);
and U21694 (N_21694,N_20723,N_20740);
nor U21695 (N_21695,N_20709,N_20722);
xor U21696 (N_21696,N_20713,N_21064);
and U21697 (N_21697,N_21147,N_20957);
or U21698 (N_21698,N_20938,N_20743);
nand U21699 (N_21699,N_20708,N_20943);
xor U21700 (N_21700,N_20699,N_20788);
or U21701 (N_21701,N_20812,N_21205);
xnor U21702 (N_21702,N_21058,N_20649);
xor U21703 (N_21703,N_20950,N_20803);
and U21704 (N_21704,N_20657,N_21227);
or U21705 (N_21705,N_21203,N_20698);
or U21706 (N_21706,N_20933,N_21011);
xnor U21707 (N_21707,N_20737,N_20761);
nand U21708 (N_21708,N_21017,N_20680);
and U21709 (N_21709,N_20839,N_20736);
nand U21710 (N_21710,N_20637,N_20826);
xnor U21711 (N_21711,N_21078,N_21047);
nor U21712 (N_21712,N_20921,N_21017);
nor U21713 (N_21713,N_20787,N_21227);
and U21714 (N_21714,N_21055,N_21212);
and U21715 (N_21715,N_20934,N_21134);
xnor U21716 (N_21716,N_20652,N_21122);
xnor U21717 (N_21717,N_21236,N_21111);
and U21718 (N_21718,N_20706,N_21165);
nor U21719 (N_21719,N_20774,N_21218);
or U21720 (N_21720,N_20908,N_21197);
xnor U21721 (N_21721,N_20961,N_21216);
nor U21722 (N_21722,N_20626,N_21065);
nand U21723 (N_21723,N_21154,N_21208);
or U21724 (N_21724,N_20767,N_20819);
xor U21725 (N_21725,N_20939,N_20760);
nand U21726 (N_21726,N_21019,N_20680);
and U21727 (N_21727,N_21067,N_20812);
nor U21728 (N_21728,N_21073,N_20811);
nor U21729 (N_21729,N_20744,N_21070);
xor U21730 (N_21730,N_21205,N_20718);
xnor U21731 (N_21731,N_20863,N_20940);
or U21732 (N_21732,N_21050,N_20635);
and U21733 (N_21733,N_20797,N_21190);
nor U21734 (N_21734,N_20762,N_20691);
nand U21735 (N_21735,N_20878,N_21182);
xor U21736 (N_21736,N_21234,N_20830);
nor U21737 (N_21737,N_21239,N_21174);
nand U21738 (N_21738,N_20747,N_20866);
and U21739 (N_21739,N_21104,N_20726);
or U21740 (N_21740,N_20993,N_21209);
nor U21741 (N_21741,N_20796,N_20926);
or U21742 (N_21742,N_21202,N_21098);
nand U21743 (N_21743,N_20905,N_20963);
xor U21744 (N_21744,N_21083,N_21075);
nor U21745 (N_21745,N_20704,N_20665);
xnor U21746 (N_21746,N_21202,N_21017);
nor U21747 (N_21747,N_20861,N_20978);
nor U21748 (N_21748,N_20801,N_21182);
nand U21749 (N_21749,N_20937,N_20628);
nand U21750 (N_21750,N_21234,N_20779);
nand U21751 (N_21751,N_21237,N_20881);
xnor U21752 (N_21752,N_20706,N_20755);
nor U21753 (N_21753,N_21090,N_21180);
or U21754 (N_21754,N_20691,N_20752);
nor U21755 (N_21755,N_21115,N_20768);
xnor U21756 (N_21756,N_20683,N_20633);
or U21757 (N_21757,N_21025,N_20689);
or U21758 (N_21758,N_20893,N_21231);
and U21759 (N_21759,N_21235,N_20773);
and U21760 (N_21760,N_20736,N_20809);
and U21761 (N_21761,N_20856,N_20630);
nor U21762 (N_21762,N_20814,N_20779);
nand U21763 (N_21763,N_21118,N_20972);
and U21764 (N_21764,N_21136,N_21174);
and U21765 (N_21765,N_20665,N_20747);
nand U21766 (N_21766,N_21190,N_20631);
nand U21767 (N_21767,N_20722,N_21080);
nor U21768 (N_21768,N_20783,N_20847);
nand U21769 (N_21769,N_21068,N_21041);
or U21770 (N_21770,N_21195,N_20982);
nor U21771 (N_21771,N_21221,N_20664);
xnor U21772 (N_21772,N_20686,N_20961);
or U21773 (N_21773,N_20944,N_21042);
and U21774 (N_21774,N_21114,N_20690);
nand U21775 (N_21775,N_21138,N_20645);
nor U21776 (N_21776,N_21039,N_21187);
and U21777 (N_21777,N_20911,N_20801);
nand U21778 (N_21778,N_21034,N_20923);
and U21779 (N_21779,N_20980,N_21037);
nand U21780 (N_21780,N_20979,N_21165);
and U21781 (N_21781,N_20843,N_21228);
or U21782 (N_21782,N_20907,N_21068);
nand U21783 (N_21783,N_21194,N_20627);
nand U21784 (N_21784,N_21006,N_20647);
nor U21785 (N_21785,N_20664,N_20663);
nor U21786 (N_21786,N_20936,N_20883);
xnor U21787 (N_21787,N_20741,N_20648);
nor U21788 (N_21788,N_21112,N_21045);
xor U21789 (N_21789,N_20916,N_20796);
nand U21790 (N_21790,N_21218,N_20894);
or U21791 (N_21791,N_20657,N_20655);
xnor U21792 (N_21792,N_20712,N_20807);
nor U21793 (N_21793,N_21139,N_21079);
or U21794 (N_21794,N_21136,N_20948);
or U21795 (N_21795,N_20863,N_21025);
and U21796 (N_21796,N_21189,N_21092);
nor U21797 (N_21797,N_20871,N_20827);
nor U21798 (N_21798,N_21133,N_21063);
xor U21799 (N_21799,N_20706,N_20931);
nor U21800 (N_21800,N_20848,N_21104);
nor U21801 (N_21801,N_21151,N_21065);
xor U21802 (N_21802,N_20911,N_20913);
nor U21803 (N_21803,N_20693,N_20761);
and U21804 (N_21804,N_20953,N_20692);
xor U21805 (N_21805,N_21063,N_20974);
xor U21806 (N_21806,N_20911,N_20899);
or U21807 (N_21807,N_20660,N_21157);
and U21808 (N_21808,N_21094,N_20639);
or U21809 (N_21809,N_20934,N_21247);
or U21810 (N_21810,N_20772,N_20682);
and U21811 (N_21811,N_21014,N_20987);
nor U21812 (N_21812,N_21223,N_21080);
nand U21813 (N_21813,N_20721,N_21055);
and U21814 (N_21814,N_21211,N_20884);
or U21815 (N_21815,N_20700,N_20901);
and U21816 (N_21816,N_20900,N_21040);
and U21817 (N_21817,N_20693,N_20679);
xor U21818 (N_21818,N_20977,N_20773);
or U21819 (N_21819,N_20930,N_21211);
and U21820 (N_21820,N_21041,N_20871);
nor U21821 (N_21821,N_20912,N_20736);
nand U21822 (N_21822,N_20949,N_20727);
nor U21823 (N_21823,N_21151,N_20651);
nand U21824 (N_21824,N_20859,N_20780);
nand U21825 (N_21825,N_21159,N_21086);
and U21826 (N_21826,N_20807,N_20794);
xor U21827 (N_21827,N_20706,N_20868);
and U21828 (N_21828,N_21019,N_20855);
or U21829 (N_21829,N_21055,N_20757);
and U21830 (N_21830,N_20757,N_20661);
or U21831 (N_21831,N_20700,N_21048);
nor U21832 (N_21832,N_20883,N_21012);
or U21833 (N_21833,N_20762,N_21179);
xor U21834 (N_21834,N_21118,N_21027);
nor U21835 (N_21835,N_20979,N_20777);
nor U21836 (N_21836,N_20907,N_20809);
nor U21837 (N_21837,N_21023,N_20642);
nand U21838 (N_21838,N_20793,N_21086);
nor U21839 (N_21839,N_21115,N_20909);
and U21840 (N_21840,N_20756,N_20977);
xor U21841 (N_21841,N_20889,N_21122);
and U21842 (N_21842,N_20757,N_20940);
or U21843 (N_21843,N_20885,N_21199);
nand U21844 (N_21844,N_21076,N_20646);
nand U21845 (N_21845,N_21102,N_20884);
xor U21846 (N_21846,N_20858,N_20663);
and U21847 (N_21847,N_21004,N_21195);
and U21848 (N_21848,N_21160,N_20770);
xor U21849 (N_21849,N_21071,N_20794);
nor U21850 (N_21850,N_21076,N_21029);
xor U21851 (N_21851,N_21185,N_20655);
nand U21852 (N_21852,N_20903,N_20724);
and U21853 (N_21853,N_21126,N_20868);
and U21854 (N_21854,N_21118,N_21222);
or U21855 (N_21855,N_20639,N_20794);
or U21856 (N_21856,N_21071,N_21032);
nor U21857 (N_21857,N_21155,N_21187);
and U21858 (N_21858,N_20787,N_21228);
and U21859 (N_21859,N_20632,N_20835);
nor U21860 (N_21860,N_21153,N_20718);
or U21861 (N_21861,N_21218,N_21130);
and U21862 (N_21862,N_21011,N_21035);
xnor U21863 (N_21863,N_20643,N_20691);
and U21864 (N_21864,N_20656,N_21168);
xnor U21865 (N_21865,N_21033,N_20815);
and U21866 (N_21866,N_20837,N_20770);
and U21867 (N_21867,N_20817,N_20954);
and U21868 (N_21868,N_21202,N_20961);
and U21869 (N_21869,N_21038,N_21154);
or U21870 (N_21870,N_21024,N_20857);
nor U21871 (N_21871,N_21161,N_21185);
and U21872 (N_21872,N_20641,N_20896);
xor U21873 (N_21873,N_21019,N_21227);
nand U21874 (N_21874,N_20784,N_21241);
nor U21875 (N_21875,N_21790,N_21383);
nor U21876 (N_21876,N_21621,N_21452);
and U21877 (N_21877,N_21727,N_21746);
or U21878 (N_21878,N_21289,N_21367);
and U21879 (N_21879,N_21281,N_21374);
nand U21880 (N_21880,N_21486,N_21574);
and U21881 (N_21881,N_21445,N_21840);
nand U21882 (N_21882,N_21769,N_21555);
nand U21883 (N_21883,N_21552,N_21647);
nand U21884 (N_21884,N_21791,N_21829);
xor U21885 (N_21885,N_21314,N_21601);
nor U21886 (N_21886,N_21300,N_21804);
nand U21887 (N_21887,N_21515,N_21352);
nor U21888 (N_21888,N_21873,N_21558);
or U21889 (N_21889,N_21807,N_21378);
xor U21890 (N_21890,N_21866,N_21660);
nand U21891 (N_21891,N_21571,N_21475);
and U21892 (N_21892,N_21382,N_21424);
nand U21893 (N_21893,N_21604,N_21573);
or U21894 (N_21894,N_21322,N_21526);
nand U21895 (N_21895,N_21666,N_21407);
xor U21896 (N_21896,N_21413,N_21419);
nor U21897 (N_21897,N_21271,N_21462);
and U21898 (N_21898,N_21653,N_21345);
and U21899 (N_21899,N_21737,N_21635);
xor U21900 (N_21900,N_21631,N_21576);
nor U21901 (N_21901,N_21533,N_21273);
and U21902 (N_21902,N_21312,N_21388);
nand U21903 (N_21903,N_21588,N_21390);
and U21904 (N_21904,N_21251,N_21614);
nand U21905 (N_21905,N_21285,N_21639);
and U21906 (N_21906,N_21584,N_21747);
nand U21907 (N_21907,N_21557,N_21793);
and U21908 (N_21908,N_21669,N_21288);
and U21909 (N_21909,N_21609,N_21753);
or U21910 (N_21910,N_21250,N_21270);
xnor U21911 (N_21911,N_21633,N_21376);
xor U21912 (N_21912,N_21551,N_21550);
nand U21913 (N_21913,N_21869,N_21538);
nand U21914 (N_21914,N_21825,N_21777);
nor U21915 (N_21915,N_21366,N_21658);
and U21916 (N_21916,N_21556,N_21703);
or U21917 (N_21917,N_21547,N_21763);
or U21918 (N_21918,N_21835,N_21774);
and U21919 (N_21919,N_21872,N_21582);
and U21920 (N_21920,N_21827,N_21710);
and U21921 (N_21921,N_21623,N_21491);
xor U21922 (N_21922,N_21781,N_21401);
or U21923 (N_21923,N_21455,N_21267);
xnor U21924 (N_21924,N_21411,N_21615);
nand U21925 (N_21925,N_21393,N_21854);
nand U21926 (N_21926,N_21570,N_21684);
nor U21927 (N_21927,N_21524,N_21649);
nand U21928 (N_21928,N_21467,N_21287);
and U21929 (N_21929,N_21479,N_21853);
and U21930 (N_21930,N_21762,N_21437);
nand U21931 (N_21931,N_21333,N_21328);
xor U21932 (N_21932,N_21778,N_21788);
nand U21933 (N_21933,N_21792,N_21372);
and U21934 (N_21934,N_21798,N_21838);
or U21935 (N_21935,N_21801,N_21664);
xnor U21936 (N_21936,N_21643,N_21338);
nor U21937 (N_21937,N_21448,N_21339);
xor U21938 (N_21938,N_21433,N_21868);
and U21939 (N_21939,N_21266,N_21818);
nor U21940 (N_21940,N_21704,N_21566);
nor U21941 (N_21941,N_21325,N_21430);
or U21942 (N_21942,N_21600,N_21292);
nor U21943 (N_21943,N_21644,N_21849);
nor U21944 (N_21944,N_21662,N_21484);
or U21945 (N_21945,N_21408,N_21326);
and U21946 (N_21946,N_21867,N_21636);
xor U21947 (N_21947,N_21841,N_21559);
nor U21948 (N_21948,N_21745,N_21441);
xnor U21949 (N_21949,N_21307,N_21375);
nor U21950 (N_21950,N_21725,N_21805);
nand U21951 (N_21951,N_21482,N_21799);
xor U21952 (N_21952,N_21264,N_21523);
nor U21953 (N_21953,N_21688,N_21539);
or U21954 (N_21954,N_21580,N_21506);
nor U21955 (N_21955,N_21504,N_21820);
nor U21956 (N_21956,N_21443,N_21412);
and U21957 (N_21957,N_21404,N_21565);
and U21958 (N_21958,N_21837,N_21630);
nor U21959 (N_21959,N_21634,N_21530);
nand U21960 (N_21960,N_21641,N_21396);
or U21961 (N_21961,N_21739,N_21817);
nor U21962 (N_21962,N_21864,N_21668);
nor U21963 (N_21963,N_21808,N_21765);
or U21964 (N_21964,N_21597,N_21712);
or U21965 (N_21965,N_21714,N_21253);
nor U21966 (N_21966,N_21436,N_21358);
xor U21967 (N_21967,N_21269,N_21625);
nand U21968 (N_21968,N_21719,N_21537);
xnor U21969 (N_21969,N_21613,N_21650);
nor U21970 (N_21970,N_21832,N_21489);
and U21971 (N_21971,N_21286,N_21473);
nor U21972 (N_21972,N_21834,N_21816);
nor U21973 (N_21973,N_21729,N_21255);
nor U21974 (N_21974,N_21276,N_21735);
and U21975 (N_21975,N_21562,N_21324);
and U21976 (N_21976,N_21478,N_21359);
nand U21977 (N_21977,N_21371,N_21463);
xnor U21978 (N_21978,N_21357,N_21744);
and U21979 (N_21979,N_21685,N_21284);
and U21980 (N_21980,N_21477,N_21593);
nand U21981 (N_21981,N_21458,N_21402);
or U21982 (N_21982,N_21370,N_21498);
or U21983 (N_21983,N_21709,N_21579);
and U21984 (N_21984,N_21858,N_21447);
nor U21985 (N_21985,N_21654,N_21564);
nor U21986 (N_21986,N_21466,N_21606);
and U21987 (N_21987,N_21331,N_21617);
nor U21988 (N_21988,N_21410,N_21568);
nor U21989 (N_21989,N_21356,N_21545);
xnor U21990 (N_21990,N_21578,N_21546);
and U21991 (N_21991,N_21715,N_21569);
xnor U21992 (N_21992,N_21616,N_21656);
xnor U21993 (N_21993,N_21377,N_21561);
or U21994 (N_21994,N_21700,N_21845);
and U21995 (N_21995,N_21379,N_21741);
nand U21996 (N_21996,N_21503,N_21456);
or U21997 (N_21997,N_21335,N_21696);
or U21998 (N_21998,N_21296,N_21529);
or U21999 (N_21999,N_21342,N_21416);
or U22000 (N_22000,N_21469,N_21786);
nor U22001 (N_22001,N_21351,N_21549);
xnor U22002 (N_22002,N_21518,N_21680);
and U22003 (N_22003,N_21317,N_21585);
or U22004 (N_22004,N_21787,N_21398);
nor U22005 (N_22005,N_21295,N_21797);
or U22006 (N_22006,N_21290,N_21732);
nand U22007 (N_22007,N_21364,N_21567);
nor U22008 (N_22008,N_21676,N_21507);
or U22009 (N_22009,N_21646,N_21803);
or U22010 (N_22010,N_21389,N_21303);
nor U22011 (N_22011,N_21420,N_21502);
and U22012 (N_22012,N_21794,N_21387);
xnor U22013 (N_22013,N_21397,N_21505);
nand U22014 (N_22014,N_21789,N_21319);
or U22015 (N_22015,N_21422,N_21861);
or U22016 (N_22016,N_21439,N_21348);
or U22017 (N_22017,N_21464,N_21305);
nand U22018 (N_22018,N_21771,N_21612);
nor U22019 (N_22019,N_21723,N_21687);
nor U22020 (N_22020,N_21446,N_21627);
nand U22021 (N_22021,N_21531,N_21310);
nor U22022 (N_22022,N_21427,N_21842);
and U22023 (N_22023,N_21671,N_21707);
xnor U22024 (N_22024,N_21721,N_21428);
and U22025 (N_22025,N_21252,N_21423);
nor U22026 (N_22026,N_21409,N_21283);
and U22027 (N_22027,N_21855,N_21444);
or U22028 (N_22028,N_21773,N_21716);
or U22029 (N_22029,N_21583,N_21435);
xor U22030 (N_22030,N_21485,N_21536);
xor U22031 (N_22031,N_21850,N_21831);
xor U22032 (N_22032,N_21670,N_21481);
and U22033 (N_22033,N_21690,N_21532);
nand U22034 (N_22034,N_21418,N_21293);
and U22035 (N_22035,N_21577,N_21736);
and U22036 (N_22036,N_21581,N_21492);
or U22037 (N_22037,N_21391,N_21760);
nor U22038 (N_22038,N_21839,N_21749);
or U22039 (N_22039,N_21767,N_21496);
nor U22040 (N_22040,N_21618,N_21318);
xor U22041 (N_22041,N_21628,N_21860);
nand U22042 (N_22042,N_21513,N_21501);
xnor U22043 (N_22043,N_21764,N_21701);
and U22044 (N_22044,N_21655,N_21663);
nor U22045 (N_22045,N_21493,N_21302);
or U22046 (N_22046,N_21355,N_21697);
and U22047 (N_22047,N_21728,N_21373);
nor U22048 (N_22048,N_21857,N_21472);
or U22049 (N_22049,N_21598,N_21748);
nor U22050 (N_22050,N_21519,N_21674);
nand U22051 (N_22051,N_21752,N_21677);
nand U22052 (N_22052,N_21278,N_21432);
and U22053 (N_22053,N_21711,N_21731);
nor U22054 (N_22054,N_21354,N_21806);
or U22055 (N_22055,N_21535,N_21488);
or U22056 (N_22056,N_21695,N_21306);
or U22057 (N_22057,N_21821,N_21626);
or U22058 (N_22058,N_21599,N_21282);
and U22059 (N_22059,N_21415,N_21470);
and U22060 (N_22060,N_21694,N_21844);
nor U22061 (N_22061,N_21812,N_21785);
and U22062 (N_22062,N_21607,N_21349);
xnor U22063 (N_22063,N_21309,N_21595);
xnor U22064 (N_22064,N_21642,N_21361);
xnor U22065 (N_22065,N_21843,N_21661);
and U22066 (N_22066,N_21483,N_21534);
or U22067 (N_22067,N_21454,N_21648);
nand U22068 (N_22068,N_21421,N_21717);
and U22069 (N_22069,N_21321,N_21657);
nor U22070 (N_22070,N_21743,N_21261);
and U22071 (N_22071,N_21605,N_21724);
or U22072 (N_22072,N_21499,N_21759);
nand U22073 (N_22073,N_21259,N_21543);
and U22074 (N_22074,N_21602,N_21332);
nor U22075 (N_22075,N_21770,N_21809);
xnor U22076 (N_22076,N_21802,N_21330);
and U22077 (N_22077,N_21541,N_21299);
nand U22078 (N_22078,N_21343,N_21863);
xnor U22079 (N_22079,N_21638,N_21368);
nand U22080 (N_22080,N_21722,N_21603);
and U22081 (N_22081,N_21308,N_21386);
nor U22082 (N_22082,N_21414,N_21851);
and U22083 (N_22083,N_21672,N_21750);
or U22084 (N_22084,N_21692,N_21651);
nor U22085 (N_22085,N_21399,N_21346);
nand U22086 (N_22086,N_21874,N_21311);
or U22087 (N_22087,N_21652,N_21275);
xor U22088 (N_22088,N_21590,N_21337);
or U22089 (N_22089,N_21780,N_21673);
xor U22090 (N_22090,N_21540,N_21836);
nand U22091 (N_22091,N_21406,N_21822);
and U22092 (N_22092,N_21796,N_21608);
xor U22093 (N_22093,N_21553,N_21675);
nand U22094 (N_22094,N_21682,N_21340);
and U22095 (N_22095,N_21800,N_21548);
nand U22096 (N_22096,N_21563,N_21544);
nand U22097 (N_22097,N_21783,N_21334);
xnor U22098 (N_22098,N_21510,N_21596);
or U22099 (N_22099,N_21527,N_21450);
nor U22100 (N_22100,N_21329,N_21279);
or U22101 (N_22101,N_21811,N_21591);
nand U22102 (N_22102,N_21733,N_21575);
or U22103 (N_22103,N_21678,N_21495);
and U22104 (N_22104,N_21718,N_21681);
and U22105 (N_22105,N_21830,N_21742);
xor U22106 (N_22106,N_21619,N_21637);
nand U22107 (N_22107,N_21517,N_21708);
nor U22108 (N_22108,N_21826,N_21665);
or U22109 (N_22109,N_21726,N_21341);
nor U22110 (N_22110,N_21686,N_21611);
nor U22111 (N_22111,N_21586,N_21350);
nor U22112 (N_22112,N_21620,N_21395);
and U22113 (N_22113,N_21693,N_21813);
and U22114 (N_22114,N_21405,N_21667);
and U22115 (N_22115,N_21698,N_21865);
nor U22116 (N_22116,N_21766,N_21320);
nor U22117 (N_22117,N_21756,N_21468);
nand U22118 (N_22118,N_21344,N_21438);
and U22119 (N_22119,N_21757,N_21699);
or U22120 (N_22120,N_21852,N_21316);
xnor U22121 (N_22121,N_21294,N_21500);
nand U22122 (N_22122,N_21683,N_21272);
or U22123 (N_22123,N_21847,N_21828);
xnor U22124 (N_22124,N_21775,N_21521);
or U22125 (N_22125,N_21417,N_21347);
and U22126 (N_22126,N_21610,N_21560);
nor U22127 (N_22127,N_21740,N_21297);
nor U22128 (N_22128,N_21480,N_21870);
or U22129 (N_22129,N_21385,N_21460);
nand U22130 (N_22130,N_21810,N_21449);
xor U22131 (N_22131,N_21327,N_21819);
and U22132 (N_22132,N_21795,N_21512);
xnor U22133 (N_22133,N_21516,N_21862);
nor U22134 (N_22134,N_21824,N_21301);
or U22135 (N_22135,N_21465,N_21514);
nand U22136 (N_22136,N_21440,N_21542);
nand U22137 (N_22137,N_21846,N_21362);
nor U22138 (N_22138,N_21772,N_21280);
xnor U22139 (N_22139,N_21257,N_21476);
xnor U22140 (N_22140,N_21525,N_21429);
xor U22141 (N_22141,N_21426,N_21365);
xor U22142 (N_22142,N_21451,N_21823);
or U22143 (N_22143,N_21291,N_21833);
or U22144 (N_22144,N_21702,N_21814);
nor U22145 (N_22145,N_21640,N_21730);
nor U22146 (N_22146,N_21323,N_21490);
and U22147 (N_22147,N_21629,N_21848);
or U22148 (N_22148,N_21442,N_21400);
nor U22149 (N_22149,N_21751,N_21254);
nand U22150 (N_22150,N_21520,N_21632);
and U22151 (N_22151,N_21815,N_21494);
xor U22152 (N_22152,N_21784,N_21782);
nand U22153 (N_22153,N_21256,N_21758);
and U22154 (N_22154,N_21511,N_21645);
and U22155 (N_22155,N_21554,N_21471);
nor U22156 (N_22156,N_21497,N_21720);
or U22157 (N_22157,N_21755,N_21260);
xnor U22158 (N_22158,N_21457,N_21509);
and U22159 (N_22159,N_21353,N_21689);
and U22160 (N_22160,N_21474,N_21381);
xor U22161 (N_22161,N_21734,N_21392);
nor U22162 (N_22162,N_21336,N_21434);
or U22163 (N_22163,N_21369,N_21268);
xor U22164 (N_22164,N_21659,N_21713);
and U22165 (N_22165,N_21360,N_21738);
nand U22166 (N_22166,N_21691,N_21315);
nor U22167 (N_22167,N_21754,N_21508);
xnor U22168 (N_22168,N_21461,N_21587);
or U22169 (N_22169,N_21425,N_21594);
or U22170 (N_22170,N_21776,N_21313);
and U22171 (N_22171,N_21856,N_21262);
nand U22172 (N_22172,N_21768,N_21705);
xor U22173 (N_22173,N_21871,N_21622);
and U22174 (N_22174,N_21453,N_21403);
xor U22175 (N_22175,N_21363,N_21522);
nor U22176 (N_22176,N_21528,N_21592);
or U22177 (N_22177,N_21572,N_21624);
or U22178 (N_22178,N_21380,N_21258);
nor U22179 (N_22179,N_21431,N_21761);
xnor U22180 (N_22180,N_21589,N_21394);
nand U22181 (N_22181,N_21265,N_21263);
nor U22182 (N_22182,N_21679,N_21487);
and U22183 (N_22183,N_21779,N_21277);
and U22184 (N_22184,N_21859,N_21304);
nand U22185 (N_22185,N_21298,N_21274);
xor U22186 (N_22186,N_21459,N_21706);
xor U22187 (N_22187,N_21384,N_21454);
nor U22188 (N_22188,N_21817,N_21395);
and U22189 (N_22189,N_21716,N_21668);
nand U22190 (N_22190,N_21604,N_21713);
nor U22191 (N_22191,N_21318,N_21534);
and U22192 (N_22192,N_21718,N_21498);
and U22193 (N_22193,N_21509,N_21551);
nand U22194 (N_22194,N_21809,N_21581);
nand U22195 (N_22195,N_21397,N_21704);
and U22196 (N_22196,N_21763,N_21773);
xor U22197 (N_22197,N_21455,N_21665);
and U22198 (N_22198,N_21363,N_21712);
and U22199 (N_22199,N_21569,N_21684);
xor U22200 (N_22200,N_21596,N_21409);
and U22201 (N_22201,N_21856,N_21685);
xor U22202 (N_22202,N_21480,N_21358);
nor U22203 (N_22203,N_21553,N_21454);
xnor U22204 (N_22204,N_21275,N_21533);
or U22205 (N_22205,N_21564,N_21831);
nor U22206 (N_22206,N_21576,N_21547);
nand U22207 (N_22207,N_21671,N_21605);
nor U22208 (N_22208,N_21399,N_21598);
and U22209 (N_22209,N_21428,N_21534);
nor U22210 (N_22210,N_21662,N_21696);
nand U22211 (N_22211,N_21776,N_21384);
or U22212 (N_22212,N_21541,N_21349);
nand U22213 (N_22213,N_21742,N_21869);
nor U22214 (N_22214,N_21487,N_21540);
and U22215 (N_22215,N_21663,N_21688);
xnor U22216 (N_22216,N_21530,N_21667);
or U22217 (N_22217,N_21513,N_21496);
nand U22218 (N_22218,N_21664,N_21484);
and U22219 (N_22219,N_21759,N_21764);
and U22220 (N_22220,N_21811,N_21314);
nand U22221 (N_22221,N_21543,N_21793);
and U22222 (N_22222,N_21588,N_21385);
nor U22223 (N_22223,N_21447,N_21309);
or U22224 (N_22224,N_21794,N_21850);
xnor U22225 (N_22225,N_21268,N_21459);
or U22226 (N_22226,N_21627,N_21706);
and U22227 (N_22227,N_21714,N_21546);
nor U22228 (N_22228,N_21590,N_21346);
and U22229 (N_22229,N_21643,N_21780);
or U22230 (N_22230,N_21348,N_21784);
xor U22231 (N_22231,N_21804,N_21779);
nand U22232 (N_22232,N_21297,N_21519);
nor U22233 (N_22233,N_21678,N_21707);
and U22234 (N_22234,N_21502,N_21737);
and U22235 (N_22235,N_21865,N_21296);
and U22236 (N_22236,N_21662,N_21552);
xnor U22237 (N_22237,N_21627,N_21829);
and U22238 (N_22238,N_21696,N_21562);
or U22239 (N_22239,N_21819,N_21700);
xnor U22240 (N_22240,N_21600,N_21344);
nand U22241 (N_22241,N_21767,N_21713);
nor U22242 (N_22242,N_21817,N_21800);
xor U22243 (N_22243,N_21723,N_21478);
xor U22244 (N_22244,N_21515,N_21735);
nor U22245 (N_22245,N_21586,N_21684);
nand U22246 (N_22246,N_21489,N_21292);
and U22247 (N_22247,N_21312,N_21475);
nor U22248 (N_22248,N_21826,N_21855);
or U22249 (N_22249,N_21632,N_21318);
and U22250 (N_22250,N_21721,N_21584);
nor U22251 (N_22251,N_21620,N_21261);
xor U22252 (N_22252,N_21807,N_21409);
or U22253 (N_22253,N_21387,N_21541);
or U22254 (N_22254,N_21378,N_21418);
or U22255 (N_22255,N_21357,N_21613);
nand U22256 (N_22256,N_21448,N_21860);
nand U22257 (N_22257,N_21443,N_21653);
xor U22258 (N_22258,N_21393,N_21400);
nand U22259 (N_22259,N_21663,N_21504);
or U22260 (N_22260,N_21342,N_21816);
nor U22261 (N_22261,N_21332,N_21673);
nor U22262 (N_22262,N_21267,N_21500);
nand U22263 (N_22263,N_21701,N_21456);
nand U22264 (N_22264,N_21447,N_21688);
nand U22265 (N_22265,N_21252,N_21659);
or U22266 (N_22266,N_21679,N_21610);
nor U22267 (N_22267,N_21494,N_21701);
nor U22268 (N_22268,N_21295,N_21326);
and U22269 (N_22269,N_21484,N_21512);
and U22270 (N_22270,N_21605,N_21731);
xnor U22271 (N_22271,N_21328,N_21460);
nor U22272 (N_22272,N_21277,N_21576);
or U22273 (N_22273,N_21736,N_21395);
or U22274 (N_22274,N_21348,N_21252);
and U22275 (N_22275,N_21680,N_21757);
or U22276 (N_22276,N_21733,N_21697);
xor U22277 (N_22277,N_21760,N_21654);
nand U22278 (N_22278,N_21295,N_21253);
xnor U22279 (N_22279,N_21829,N_21283);
and U22280 (N_22280,N_21718,N_21506);
xnor U22281 (N_22281,N_21501,N_21262);
or U22282 (N_22282,N_21792,N_21718);
nand U22283 (N_22283,N_21778,N_21342);
nand U22284 (N_22284,N_21605,N_21670);
xor U22285 (N_22285,N_21608,N_21635);
xnor U22286 (N_22286,N_21604,N_21812);
or U22287 (N_22287,N_21495,N_21390);
xnor U22288 (N_22288,N_21819,N_21270);
xnor U22289 (N_22289,N_21693,N_21375);
or U22290 (N_22290,N_21787,N_21397);
xor U22291 (N_22291,N_21486,N_21863);
xnor U22292 (N_22292,N_21684,N_21553);
and U22293 (N_22293,N_21722,N_21799);
nand U22294 (N_22294,N_21671,N_21744);
or U22295 (N_22295,N_21766,N_21368);
or U22296 (N_22296,N_21337,N_21757);
nor U22297 (N_22297,N_21854,N_21314);
and U22298 (N_22298,N_21784,N_21465);
nand U22299 (N_22299,N_21524,N_21386);
nand U22300 (N_22300,N_21793,N_21639);
and U22301 (N_22301,N_21653,N_21804);
or U22302 (N_22302,N_21568,N_21277);
nor U22303 (N_22303,N_21807,N_21872);
nor U22304 (N_22304,N_21440,N_21795);
or U22305 (N_22305,N_21271,N_21440);
nor U22306 (N_22306,N_21703,N_21325);
nor U22307 (N_22307,N_21739,N_21391);
and U22308 (N_22308,N_21535,N_21388);
and U22309 (N_22309,N_21789,N_21560);
xnor U22310 (N_22310,N_21756,N_21469);
nor U22311 (N_22311,N_21443,N_21558);
nor U22312 (N_22312,N_21810,N_21823);
xor U22313 (N_22313,N_21654,N_21425);
xor U22314 (N_22314,N_21618,N_21559);
xnor U22315 (N_22315,N_21847,N_21570);
nand U22316 (N_22316,N_21424,N_21648);
xor U22317 (N_22317,N_21427,N_21272);
xor U22318 (N_22318,N_21492,N_21530);
or U22319 (N_22319,N_21555,N_21714);
nor U22320 (N_22320,N_21680,N_21698);
and U22321 (N_22321,N_21538,N_21773);
nor U22322 (N_22322,N_21654,N_21449);
xor U22323 (N_22323,N_21462,N_21316);
xnor U22324 (N_22324,N_21391,N_21665);
or U22325 (N_22325,N_21311,N_21648);
nand U22326 (N_22326,N_21356,N_21436);
nor U22327 (N_22327,N_21862,N_21376);
nor U22328 (N_22328,N_21531,N_21429);
and U22329 (N_22329,N_21382,N_21442);
or U22330 (N_22330,N_21776,N_21680);
or U22331 (N_22331,N_21656,N_21797);
nor U22332 (N_22332,N_21475,N_21442);
nand U22333 (N_22333,N_21714,N_21668);
nand U22334 (N_22334,N_21287,N_21757);
nor U22335 (N_22335,N_21594,N_21849);
xnor U22336 (N_22336,N_21843,N_21805);
or U22337 (N_22337,N_21543,N_21492);
and U22338 (N_22338,N_21507,N_21599);
nand U22339 (N_22339,N_21755,N_21478);
xnor U22340 (N_22340,N_21408,N_21456);
xor U22341 (N_22341,N_21860,N_21316);
xnor U22342 (N_22342,N_21707,N_21561);
nor U22343 (N_22343,N_21775,N_21350);
or U22344 (N_22344,N_21256,N_21592);
or U22345 (N_22345,N_21547,N_21293);
and U22346 (N_22346,N_21567,N_21302);
nand U22347 (N_22347,N_21363,N_21867);
nor U22348 (N_22348,N_21633,N_21562);
nand U22349 (N_22349,N_21591,N_21528);
nor U22350 (N_22350,N_21782,N_21738);
and U22351 (N_22351,N_21256,N_21796);
nand U22352 (N_22352,N_21676,N_21646);
or U22353 (N_22353,N_21451,N_21763);
and U22354 (N_22354,N_21549,N_21410);
nor U22355 (N_22355,N_21730,N_21347);
nand U22356 (N_22356,N_21503,N_21742);
or U22357 (N_22357,N_21254,N_21267);
or U22358 (N_22358,N_21292,N_21714);
nor U22359 (N_22359,N_21699,N_21626);
xnor U22360 (N_22360,N_21260,N_21534);
and U22361 (N_22361,N_21643,N_21810);
or U22362 (N_22362,N_21816,N_21323);
nand U22363 (N_22363,N_21777,N_21540);
xnor U22364 (N_22364,N_21839,N_21727);
nor U22365 (N_22365,N_21350,N_21389);
nand U22366 (N_22366,N_21629,N_21601);
and U22367 (N_22367,N_21345,N_21366);
xnor U22368 (N_22368,N_21718,N_21423);
nor U22369 (N_22369,N_21546,N_21560);
nor U22370 (N_22370,N_21792,N_21623);
nand U22371 (N_22371,N_21401,N_21303);
or U22372 (N_22372,N_21307,N_21818);
xnor U22373 (N_22373,N_21604,N_21410);
nor U22374 (N_22374,N_21292,N_21839);
nor U22375 (N_22375,N_21346,N_21257);
xor U22376 (N_22376,N_21854,N_21411);
or U22377 (N_22377,N_21852,N_21547);
and U22378 (N_22378,N_21561,N_21753);
nor U22379 (N_22379,N_21522,N_21738);
and U22380 (N_22380,N_21750,N_21475);
and U22381 (N_22381,N_21654,N_21842);
or U22382 (N_22382,N_21759,N_21278);
xor U22383 (N_22383,N_21694,N_21264);
nor U22384 (N_22384,N_21409,N_21509);
xor U22385 (N_22385,N_21576,N_21837);
xor U22386 (N_22386,N_21841,N_21403);
xor U22387 (N_22387,N_21807,N_21718);
nand U22388 (N_22388,N_21424,N_21583);
nor U22389 (N_22389,N_21650,N_21344);
nor U22390 (N_22390,N_21473,N_21761);
and U22391 (N_22391,N_21624,N_21412);
and U22392 (N_22392,N_21469,N_21837);
or U22393 (N_22393,N_21601,N_21332);
xor U22394 (N_22394,N_21464,N_21699);
nor U22395 (N_22395,N_21395,N_21635);
or U22396 (N_22396,N_21431,N_21821);
or U22397 (N_22397,N_21665,N_21673);
nand U22398 (N_22398,N_21782,N_21278);
nor U22399 (N_22399,N_21576,N_21368);
xor U22400 (N_22400,N_21558,N_21494);
or U22401 (N_22401,N_21288,N_21793);
nor U22402 (N_22402,N_21648,N_21866);
nor U22403 (N_22403,N_21559,N_21713);
nand U22404 (N_22404,N_21834,N_21425);
nand U22405 (N_22405,N_21575,N_21752);
nor U22406 (N_22406,N_21710,N_21347);
and U22407 (N_22407,N_21525,N_21546);
nand U22408 (N_22408,N_21438,N_21527);
and U22409 (N_22409,N_21383,N_21825);
or U22410 (N_22410,N_21262,N_21796);
xor U22411 (N_22411,N_21269,N_21763);
nor U22412 (N_22412,N_21465,N_21758);
or U22413 (N_22413,N_21669,N_21441);
nand U22414 (N_22414,N_21293,N_21519);
or U22415 (N_22415,N_21848,N_21795);
and U22416 (N_22416,N_21818,N_21672);
xor U22417 (N_22417,N_21750,N_21576);
or U22418 (N_22418,N_21376,N_21377);
nand U22419 (N_22419,N_21762,N_21303);
xnor U22420 (N_22420,N_21790,N_21504);
nand U22421 (N_22421,N_21563,N_21327);
xnor U22422 (N_22422,N_21699,N_21308);
xor U22423 (N_22423,N_21330,N_21337);
nand U22424 (N_22424,N_21450,N_21427);
and U22425 (N_22425,N_21693,N_21859);
and U22426 (N_22426,N_21686,N_21653);
nand U22427 (N_22427,N_21254,N_21522);
or U22428 (N_22428,N_21755,N_21540);
nand U22429 (N_22429,N_21389,N_21276);
nor U22430 (N_22430,N_21683,N_21314);
or U22431 (N_22431,N_21828,N_21642);
and U22432 (N_22432,N_21327,N_21370);
nand U22433 (N_22433,N_21499,N_21348);
nor U22434 (N_22434,N_21301,N_21828);
and U22435 (N_22435,N_21659,N_21479);
and U22436 (N_22436,N_21587,N_21588);
and U22437 (N_22437,N_21847,N_21551);
nand U22438 (N_22438,N_21786,N_21556);
nand U22439 (N_22439,N_21776,N_21867);
or U22440 (N_22440,N_21284,N_21374);
or U22441 (N_22441,N_21361,N_21427);
xor U22442 (N_22442,N_21796,N_21690);
and U22443 (N_22443,N_21626,N_21373);
nand U22444 (N_22444,N_21572,N_21868);
nand U22445 (N_22445,N_21579,N_21845);
or U22446 (N_22446,N_21577,N_21464);
or U22447 (N_22447,N_21579,N_21706);
nor U22448 (N_22448,N_21313,N_21359);
nand U22449 (N_22449,N_21508,N_21640);
or U22450 (N_22450,N_21670,N_21696);
or U22451 (N_22451,N_21755,N_21784);
nor U22452 (N_22452,N_21654,N_21506);
xnor U22453 (N_22453,N_21373,N_21454);
nor U22454 (N_22454,N_21626,N_21616);
nor U22455 (N_22455,N_21533,N_21756);
nand U22456 (N_22456,N_21291,N_21336);
or U22457 (N_22457,N_21455,N_21782);
nor U22458 (N_22458,N_21765,N_21422);
xor U22459 (N_22459,N_21426,N_21474);
and U22460 (N_22460,N_21439,N_21448);
nand U22461 (N_22461,N_21697,N_21322);
nand U22462 (N_22462,N_21552,N_21328);
nand U22463 (N_22463,N_21262,N_21575);
nand U22464 (N_22464,N_21527,N_21687);
nor U22465 (N_22465,N_21416,N_21280);
or U22466 (N_22466,N_21747,N_21796);
nand U22467 (N_22467,N_21699,N_21568);
xnor U22468 (N_22468,N_21594,N_21328);
nor U22469 (N_22469,N_21678,N_21614);
or U22470 (N_22470,N_21550,N_21300);
or U22471 (N_22471,N_21489,N_21769);
nand U22472 (N_22472,N_21265,N_21732);
xor U22473 (N_22473,N_21560,N_21615);
nand U22474 (N_22474,N_21803,N_21288);
or U22475 (N_22475,N_21759,N_21287);
and U22476 (N_22476,N_21687,N_21487);
xor U22477 (N_22477,N_21744,N_21639);
nor U22478 (N_22478,N_21757,N_21658);
or U22479 (N_22479,N_21427,N_21315);
xnor U22480 (N_22480,N_21459,N_21794);
nand U22481 (N_22481,N_21296,N_21663);
nor U22482 (N_22482,N_21464,N_21636);
nand U22483 (N_22483,N_21521,N_21398);
and U22484 (N_22484,N_21453,N_21455);
or U22485 (N_22485,N_21586,N_21669);
nand U22486 (N_22486,N_21706,N_21400);
nor U22487 (N_22487,N_21374,N_21252);
xnor U22488 (N_22488,N_21766,N_21701);
nor U22489 (N_22489,N_21367,N_21368);
or U22490 (N_22490,N_21485,N_21686);
and U22491 (N_22491,N_21618,N_21744);
xor U22492 (N_22492,N_21551,N_21740);
and U22493 (N_22493,N_21783,N_21282);
xor U22494 (N_22494,N_21467,N_21401);
and U22495 (N_22495,N_21638,N_21797);
nand U22496 (N_22496,N_21527,N_21845);
and U22497 (N_22497,N_21678,N_21752);
and U22498 (N_22498,N_21394,N_21293);
or U22499 (N_22499,N_21623,N_21776);
nand U22500 (N_22500,N_21903,N_22186);
or U22501 (N_22501,N_22072,N_22332);
nand U22502 (N_22502,N_22259,N_22406);
or U22503 (N_22503,N_22303,N_22291);
xnor U22504 (N_22504,N_21983,N_22223);
nor U22505 (N_22505,N_22044,N_22434);
nor U22506 (N_22506,N_22251,N_22198);
nand U22507 (N_22507,N_22344,N_21897);
nand U22508 (N_22508,N_21995,N_22420);
or U22509 (N_22509,N_22067,N_22338);
and U22510 (N_22510,N_21881,N_21909);
xor U22511 (N_22511,N_22146,N_22260);
nor U22512 (N_22512,N_22034,N_22196);
and U22513 (N_22513,N_22159,N_22378);
nor U22514 (N_22514,N_21939,N_22158);
and U22515 (N_22515,N_21933,N_22097);
or U22516 (N_22516,N_22239,N_22137);
or U22517 (N_22517,N_22087,N_22334);
and U22518 (N_22518,N_22219,N_22032);
nor U22519 (N_22519,N_22481,N_22400);
and U22520 (N_22520,N_22084,N_22021);
or U22521 (N_22521,N_22240,N_22285);
or U22522 (N_22522,N_22323,N_21892);
and U22523 (N_22523,N_22255,N_22184);
nor U22524 (N_22524,N_22248,N_21911);
and U22525 (N_22525,N_22404,N_22283);
nand U22526 (N_22526,N_22357,N_22363);
xor U22527 (N_22527,N_22138,N_22000);
and U22528 (N_22528,N_22007,N_22041);
nand U22529 (N_22529,N_22276,N_22010);
nand U22530 (N_22530,N_22225,N_22413);
xnor U22531 (N_22531,N_21955,N_21895);
nor U22532 (N_22532,N_21887,N_22215);
and U22533 (N_22533,N_22218,N_22485);
nor U22534 (N_22534,N_22499,N_22222);
nor U22535 (N_22535,N_21922,N_22487);
xor U22536 (N_22536,N_22473,N_22391);
xnor U22537 (N_22537,N_21919,N_22373);
nand U22538 (N_22538,N_22235,N_22377);
or U22539 (N_22539,N_21988,N_22091);
or U22540 (N_22540,N_22178,N_22359);
and U22541 (N_22541,N_22463,N_22236);
nand U22542 (N_22542,N_22289,N_22452);
or U22543 (N_22543,N_22011,N_22267);
or U22544 (N_22544,N_22179,N_22453);
and U22545 (N_22545,N_22203,N_22419);
nor U22546 (N_22546,N_22144,N_22100);
nor U22547 (N_22547,N_22086,N_22284);
or U22548 (N_22548,N_22350,N_21885);
or U22549 (N_22549,N_21958,N_22266);
xnor U22550 (N_22550,N_21968,N_22015);
and U22551 (N_22551,N_22166,N_21945);
xor U22552 (N_22552,N_22120,N_22183);
xor U22553 (N_22553,N_22057,N_22279);
nand U22554 (N_22554,N_22245,N_22282);
xor U22555 (N_22555,N_22448,N_22017);
and U22556 (N_22556,N_22125,N_22148);
xor U22557 (N_22557,N_22022,N_21879);
xor U22558 (N_22558,N_22168,N_22117);
and U22559 (N_22559,N_22135,N_22293);
and U22560 (N_22560,N_22066,N_22190);
xnor U22561 (N_22561,N_22016,N_22442);
nor U22562 (N_22562,N_22263,N_21970);
or U22563 (N_22563,N_22437,N_22033);
or U22564 (N_22564,N_22055,N_22409);
xor U22565 (N_22565,N_22206,N_22471);
xor U22566 (N_22566,N_22108,N_21984);
nor U22567 (N_22567,N_22336,N_22224);
nor U22568 (N_22568,N_21972,N_22256);
nand U22569 (N_22569,N_22035,N_22474);
and U22570 (N_22570,N_22164,N_22046);
and U22571 (N_22571,N_21891,N_22172);
or U22572 (N_22572,N_22369,N_22412);
nand U22573 (N_22573,N_22354,N_21947);
xor U22574 (N_22574,N_22227,N_22064);
and U22575 (N_22575,N_22189,N_22243);
nand U22576 (N_22576,N_22162,N_22229);
nor U22577 (N_22577,N_22286,N_22079);
or U22578 (N_22578,N_22273,N_22207);
nand U22579 (N_22579,N_22375,N_22492);
or U22580 (N_22580,N_22073,N_22360);
and U22581 (N_22581,N_21921,N_22423);
nand U22582 (N_22582,N_22053,N_22265);
and U22583 (N_22583,N_22109,N_22074);
nor U22584 (N_22584,N_21898,N_22362);
xor U22585 (N_22585,N_22193,N_22132);
nand U22586 (N_22586,N_22083,N_21925);
nor U22587 (N_22587,N_22330,N_21977);
nor U22588 (N_22588,N_22313,N_22005);
or U22589 (N_22589,N_21930,N_22416);
nand U22590 (N_22590,N_21913,N_22317);
and U22591 (N_22591,N_22187,N_22201);
nor U22592 (N_22592,N_22292,N_22069);
or U22593 (N_22593,N_22287,N_22226);
or U22594 (N_22594,N_21959,N_21979);
xnor U22595 (N_22595,N_22173,N_22107);
and U22596 (N_22596,N_22358,N_22361);
xor U22597 (N_22597,N_22060,N_22092);
xor U22598 (N_22598,N_22068,N_22479);
and U22599 (N_22599,N_22451,N_22456);
nand U22600 (N_22600,N_22040,N_21996);
nor U22601 (N_22601,N_22331,N_22401);
or U22602 (N_22602,N_22270,N_21993);
and U22603 (N_22603,N_22105,N_21893);
nand U22604 (N_22604,N_22150,N_22116);
and U22605 (N_22605,N_22315,N_22395);
and U22606 (N_22606,N_22444,N_21976);
nor U22607 (N_22607,N_22037,N_22488);
xor U22608 (N_22608,N_22290,N_22200);
nand U22609 (N_22609,N_22381,N_22392);
nand U22610 (N_22610,N_21875,N_22441);
nor U22611 (N_22611,N_22121,N_22050);
nand U22612 (N_22612,N_22333,N_21907);
or U22613 (N_22613,N_22128,N_22249);
xor U22614 (N_22614,N_22337,N_21936);
nor U22615 (N_22615,N_22341,N_22418);
nand U22616 (N_22616,N_21935,N_22408);
nand U22617 (N_22617,N_22304,N_22433);
nor U22618 (N_22618,N_22212,N_22071);
xnor U22619 (N_22619,N_22296,N_21908);
and U22620 (N_22620,N_22197,N_22177);
and U22621 (N_22621,N_21923,N_22280);
xnor U22622 (N_22622,N_22281,N_22153);
xnor U22623 (N_22623,N_21929,N_21927);
or U22624 (N_22624,N_22003,N_22352);
or U22625 (N_22625,N_21989,N_21987);
nor U22626 (N_22626,N_21950,N_22415);
and U22627 (N_22627,N_22062,N_22209);
and U22628 (N_22628,N_21997,N_22470);
or U22629 (N_22629,N_22300,N_22461);
and U22630 (N_22630,N_22482,N_21986);
and U22631 (N_22631,N_22440,N_21980);
nor U22632 (N_22632,N_21938,N_22048);
xor U22633 (N_22633,N_21949,N_21926);
nor U22634 (N_22634,N_22477,N_22047);
and U22635 (N_22635,N_22101,N_22013);
nor U22636 (N_22636,N_22340,N_22102);
nor U22637 (N_22637,N_21946,N_22320);
xnor U22638 (N_22638,N_22329,N_21912);
or U22639 (N_22639,N_22385,N_22090);
or U22640 (N_22640,N_21994,N_22242);
and U22641 (N_22641,N_21941,N_22335);
xor U22642 (N_22642,N_22043,N_21966);
and U22643 (N_22643,N_21937,N_22387);
nand U22644 (N_22644,N_22498,N_22151);
or U22645 (N_22645,N_22110,N_21905);
and U22646 (N_22646,N_22221,N_22009);
xor U22647 (N_22647,N_22491,N_22112);
xor U22648 (N_22648,N_22113,N_22371);
nor U22649 (N_22649,N_22462,N_22364);
nor U22650 (N_22650,N_22230,N_22428);
and U22651 (N_22651,N_22126,N_22347);
nor U22652 (N_22652,N_22233,N_21961);
xnor U22653 (N_22653,N_22081,N_21975);
xnor U22654 (N_22654,N_22351,N_22308);
nor U22655 (N_22655,N_22088,N_22051);
nor U22656 (N_22656,N_21904,N_21971);
nand U22657 (N_22657,N_22123,N_21878);
or U22658 (N_22658,N_22322,N_22275);
nor U22659 (N_22659,N_22185,N_22438);
nand U22660 (N_22660,N_22326,N_22250);
or U22661 (N_22661,N_22188,N_21954);
or U22662 (N_22662,N_22370,N_21981);
nor U22663 (N_22663,N_22211,N_22228);
or U22664 (N_22664,N_22001,N_22460);
and U22665 (N_22665,N_22169,N_21969);
nand U22666 (N_22666,N_22403,N_22075);
or U22667 (N_22667,N_22268,N_22214);
xor U22668 (N_22668,N_22455,N_22042);
or U22669 (N_22669,N_22136,N_22254);
nand U22670 (N_22670,N_21900,N_22099);
or U22671 (N_22671,N_22143,N_21880);
nand U22672 (N_22672,N_22008,N_22124);
xor U22673 (N_22673,N_22096,N_22494);
nand U22674 (N_22674,N_21992,N_21899);
or U22675 (N_22675,N_21951,N_22439);
xor U22676 (N_22676,N_22443,N_22195);
and U22677 (N_22677,N_22157,N_22390);
xor U22678 (N_22678,N_22339,N_22237);
nor U22679 (N_22679,N_22495,N_22277);
xnor U22680 (N_22680,N_22253,N_22383);
and U22681 (N_22681,N_21963,N_22122);
xnor U22682 (N_22682,N_22141,N_22054);
nand U22683 (N_22683,N_22305,N_22098);
xor U22684 (N_22684,N_22059,N_22468);
xor U22685 (N_22685,N_22382,N_22376);
xor U22686 (N_22686,N_22103,N_22213);
and U22687 (N_22687,N_22307,N_22111);
and U22688 (N_22688,N_22171,N_21882);
nand U22689 (N_22689,N_22131,N_22104);
nor U22690 (N_22690,N_22476,N_21974);
or U22691 (N_22691,N_22127,N_22147);
nor U22692 (N_22692,N_22119,N_22346);
or U22693 (N_22693,N_22061,N_22274);
and U22694 (N_22694,N_21931,N_22410);
and U22695 (N_22695,N_22244,N_21985);
nand U22696 (N_22696,N_22134,N_21894);
xnor U22697 (N_22697,N_22085,N_22310);
or U22698 (N_22698,N_22258,N_21999);
xor U22699 (N_22699,N_22130,N_21973);
nand U22700 (N_22700,N_21960,N_22324);
and U22701 (N_22701,N_21914,N_22149);
and U22702 (N_22702,N_22058,N_22167);
nand U22703 (N_22703,N_22036,N_21952);
nor U22704 (N_22704,N_22002,N_22379);
and U22705 (N_22705,N_22398,N_21886);
nand U22706 (N_22706,N_22238,N_21940);
or U22707 (N_22707,N_22095,N_22252);
xnor U22708 (N_22708,N_22264,N_22205);
and U22709 (N_22709,N_22247,N_21915);
xnor U22710 (N_22710,N_22430,N_22397);
nor U22711 (N_22711,N_21901,N_21998);
xor U22712 (N_22712,N_21890,N_22368);
nand U22713 (N_22713,N_22489,N_22045);
nand U22714 (N_22714,N_22165,N_22140);
or U22715 (N_22715,N_22160,N_22393);
nor U22716 (N_22716,N_21889,N_22475);
or U22717 (N_22717,N_21896,N_22319);
nor U22718 (N_22718,N_22272,N_22464);
and U22719 (N_22719,N_22139,N_22161);
xor U22720 (N_22720,N_22269,N_21876);
and U22721 (N_22721,N_22306,N_22199);
and U22722 (N_22722,N_22380,N_21957);
nor U22723 (N_22723,N_21944,N_22309);
xor U22724 (N_22724,N_22325,N_22316);
nor U22725 (N_22725,N_22114,N_22450);
or U22726 (N_22726,N_22082,N_21943);
nand U22727 (N_22727,N_21934,N_22429);
xnor U22728 (N_22728,N_22342,N_22155);
nand U22729 (N_22729,N_22065,N_22278);
or U22730 (N_22730,N_22175,N_22421);
and U22731 (N_22731,N_22449,N_22145);
and U22732 (N_22732,N_22445,N_22356);
nor U22733 (N_22733,N_22355,N_21978);
nand U22734 (N_22734,N_22049,N_22469);
or U22735 (N_22735,N_22029,N_21991);
nor U22736 (N_22736,N_22093,N_21888);
nor U22737 (N_22737,N_22407,N_22204);
nand U22738 (N_22738,N_22388,N_22394);
nor U22739 (N_22739,N_22129,N_22194);
xnor U22740 (N_22740,N_22241,N_22056);
nand U22741 (N_22741,N_22353,N_22070);
nor U22742 (N_22742,N_22202,N_22454);
and U22743 (N_22743,N_22374,N_22025);
nand U22744 (N_22744,N_22026,N_22435);
xor U22745 (N_22745,N_22295,N_22457);
xnor U22746 (N_22746,N_22318,N_22483);
nand U22747 (N_22747,N_22302,N_21877);
xnor U22748 (N_22748,N_22447,N_21902);
nor U22749 (N_22749,N_21982,N_21942);
or U22750 (N_22750,N_22031,N_21924);
nor U22751 (N_22751,N_22163,N_22261);
nand U22752 (N_22752,N_22367,N_22343);
nor U22753 (N_22753,N_22301,N_22180);
nor U22754 (N_22754,N_22038,N_21928);
nor U22755 (N_22755,N_22411,N_22389);
nor U22756 (N_22756,N_21990,N_22484);
or U22757 (N_22757,N_22432,N_22118);
xor U22758 (N_22758,N_22297,N_22349);
xnor U22759 (N_22759,N_22497,N_22019);
xnor U22760 (N_22760,N_22312,N_21967);
and U22761 (N_22761,N_22446,N_22076);
xor U22762 (N_22762,N_22386,N_22142);
nand U22763 (N_22763,N_22262,N_22217);
and U22764 (N_22764,N_22399,N_22094);
or U22765 (N_22765,N_22472,N_22314);
and U22766 (N_22766,N_22458,N_22366);
xnor U22767 (N_22767,N_22288,N_22004);
or U22768 (N_22768,N_22311,N_22181);
and U22769 (N_22769,N_21956,N_21920);
nor U22770 (N_22770,N_22208,N_22372);
nand U22771 (N_22771,N_22176,N_22012);
or U22772 (N_22772,N_22170,N_22467);
or U22773 (N_22773,N_22246,N_22478);
nor U22774 (N_22774,N_22425,N_22384);
nor U22775 (N_22775,N_22271,N_22365);
nand U22776 (N_22776,N_22321,N_22152);
or U22777 (N_22777,N_22182,N_22257);
xor U22778 (N_22778,N_22298,N_22327);
and U22779 (N_22779,N_22028,N_21964);
nand U22780 (N_22780,N_22345,N_22466);
and U22781 (N_22781,N_21910,N_22089);
and U22782 (N_22782,N_22052,N_22431);
nand U22783 (N_22783,N_21948,N_22422);
or U22784 (N_22784,N_22133,N_22014);
and U22785 (N_22785,N_22232,N_21918);
or U22786 (N_22786,N_22027,N_22490);
and U22787 (N_22787,N_22174,N_22424);
or U22788 (N_22788,N_21953,N_22459);
nor U22789 (N_22789,N_22493,N_22191);
xor U22790 (N_22790,N_22023,N_22024);
and U22791 (N_22791,N_22299,N_22436);
nand U22792 (N_22792,N_22020,N_22192);
xor U22793 (N_22793,N_22063,N_22115);
xnor U22794 (N_22794,N_22402,N_22080);
nor U22795 (N_22795,N_22348,N_22234);
xnor U22796 (N_22796,N_22405,N_22220);
nand U22797 (N_22797,N_21965,N_21962);
nand U22798 (N_22798,N_22216,N_22156);
nand U22799 (N_22799,N_22006,N_22231);
nand U22800 (N_22800,N_22078,N_22077);
nor U22801 (N_22801,N_22480,N_21884);
or U22802 (N_22802,N_22210,N_22106);
or U22803 (N_22803,N_21916,N_22396);
nand U22804 (N_22804,N_21906,N_22039);
nand U22805 (N_22805,N_21883,N_22018);
nand U22806 (N_22806,N_22294,N_22426);
nor U22807 (N_22807,N_22496,N_22030);
nand U22808 (N_22808,N_22154,N_22486);
or U22809 (N_22809,N_21932,N_22328);
nand U22810 (N_22810,N_22465,N_22417);
or U22811 (N_22811,N_22414,N_22427);
xnor U22812 (N_22812,N_21917,N_22190);
nand U22813 (N_22813,N_22201,N_22284);
xnor U22814 (N_22814,N_22313,N_22449);
nand U22815 (N_22815,N_22270,N_21940);
or U22816 (N_22816,N_22010,N_22360);
nand U22817 (N_22817,N_21895,N_22279);
or U22818 (N_22818,N_22170,N_22386);
nor U22819 (N_22819,N_22385,N_22495);
nand U22820 (N_22820,N_22249,N_22304);
and U22821 (N_22821,N_22021,N_21899);
or U22822 (N_22822,N_22215,N_22006);
or U22823 (N_22823,N_22454,N_22050);
nor U22824 (N_22824,N_22430,N_22316);
nor U22825 (N_22825,N_22386,N_22211);
and U22826 (N_22826,N_22466,N_22347);
or U22827 (N_22827,N_22081,N_22299);
nand U22828 (N_22828,N_22429,N_21977);
and U22829 (N_22829,N_22350,N_22211);
nand U22830 (N_22830,N_22411,N_22175);
or U22831 (N_22831,N_22364,N_22069);
or U22832 (N_22832,N_22488,N_22493);
nor U22833 (N_22833,N_22227,N_22315);
xor U22834 (N_22834,N_22309,N_22214);
xnor U22835 (N_22835,N_22143,N_22356);
or U22836 (N_22836,N_21909,N_22401);
and U22837 (N_22837,N_22323,N_22159);
xnor U22838 (N_22838,N_22068,N_22409);
xor U22839 (N_22839,N_21938,N_22161);
nor U22840 (N_22840,N_22069,N_22050);
nor U22841 (N_22841,N_22113,N_22155);
and U22842 (N_22842,N_22371,N_22298);
or U22843 (N_22843,N_22204,N_22110);
or U22844 (N_22844,N_21965,N_22046);
and U22845 (N_22845,N_22499,N_22029);
nand U22846 (N_22846,N_22186,N_22400);
nand U22847 (N_22847,N_22063,N_22049);
xnor U22848 (N_22848,N_22407,N_21924);
nor U22849 (N_22849,N_22244,N_22023);
xnor U22850 (N_22850,N_21934,N_21933);
xnor U22851 (N_22851,N_22341,N_22463);
xor U22852 (N_22852,N_22498,N_22349);
xnor U22853 (N_22853,N_21930,N_21990);
and U22854 (N_22854,N_22322,N_22303);
and U22855 (N_22855,N_22163,N_22325);
and U22856 (N_22856,N_22434,N_22226);
and U22857 (N_22857,N_22412,N_22148);
xor U22858 (N_22858,N_22014,N_22322);
and U22859 (N_22859,N_22354,N_22046);
xnor U22860 (N_22860,N_22227,N_22464);
or U22861 (N_22861,N_22010,N_22165);
nand U22862 (N_22862,N_22373,N_22152);
and U22863 (N_22863,N_22141,N_22206);
nor U22864 (N_22864,N_22037,N_22458);
nor U22865 (N_22865,N_22447,N_22261);
or U22866 (N_22866,N_21906,N_21951);
and U22867 (N_22867,N_22111,N_22399);
xnor U22868 (N_22868,N_22397,N_22171);
nand U22869 (N_22869,N_22390,N_22424);
and U22870 (N_22870,N_22447,N_22380);
nand U22871 (N_22871,N_22062,N_22488);
xor U22872 (N_22872,N_22166,N_22144);
or U22873 (N_22873,N_22117,N_21914);
and U22874 (N_22874,N_22096,N_22152);
nand U22875 (N_22875,N_22005,N_22111);
nand U22876 (N_22876,N_22002,N_21984);
xor U22877 (N_22877,N_22153,N_21996);
nor U22878 (N_22878,N_22080,N_22194);
xor U22879 (N_22879,N_22017,N_21885);
and U22880 (N_22880,N_22082,N_22129);
xor U22881 (N_22881,N_22271,N_22066);
and U22882 (N_22882,N_22437,N_22068);
or U22883 (N_22883,N_22432,N_22379);
or U22884 (N_22884,N_21977,N_21991);
and U22885 (N_22885,N_22056,N_22206);
xor U22886 (N_22886,N_22468,N_22199);
xnor U22887 (N_22887,N_22131,N_21926);
or U22888 (N_22888,N_22481,N_22023);
nor U22889 (N_22889,N_22201,N_22451);
xor U22890 (N_22890,N_22202,N_22491);
and U22891 (N_22891,N_22000,N_21927);
nor U22892 (N_22892,N_22152,N_22240);
or U22893 (N_22893,N_21920,N_22348);
and U22894 (N_22894,N_22313,N_22048);
or U22895 (N_22895,N_22309,N_22075);
and U22896 (N_22896,N_22107,N_22062);
xor U22897 (N_22897,N_22220,N_22015);
and U22898 (N_22898,N_22287,N_21900);
xor U22899 (N_22899,N_22055,N_22291);
nand U22900 (N_22900,N_21959,N_22001);
nor U22901 (N_22901,N_21890,N_22491);
or U22902 (N_22902,N_21911,N_22281);
xor U22903 (N_22903,N_22400,N_22409);
nor U22904 (N_22904,N_22236,N_21951);
or U22905 (N_22905,N_22333,N_22016);
xnor U22906 (N_22906,N_21979,N_21976);
and U22907 (N_22907,N_22436,N_22210);
xor U22908 (N_22908,N_22324,N_22207);
and U22909 (N_22909,N_22236,N_22325);
nand U22910 (N_22910,N_21876,N_22314);
nor U22911 (N_22911,N_22139,N_22003);
and U22912 (N_22912,N_22455,N_22203);
nand U22913 (N_22913,N_22031,N_22071);
nand U22914 (N_22914,N_22305,N_22025);
nand U22915 (N_22915,N_22494,N_22243);
nand U22916 (N_22916,N_21896,N_22427);
nor U22917 (N_22917,N_22405,N_22376);
xor U22918 (N_22918,N_21880,N_22251);
xnor U22919 (N_22919,N_22317,N_21927);
nor U22920 (N_22920,N_22220,N_22414);
nand U22921 (N_22921,N_22179,N_22123);
or U22922 (N_22922,N_22097,N_22026);
and U22923 (N_22923,N_22173,N_22282);
and U22924 (N_22924,N_22270,N_21915);
nand U22925 (N_22925,N_22117,N_22439);
xor U22926 (N_22926,N_22462,N_21978);
nand U22927 (N_22927,N_21992,N_22379);
nand U22928 (N_22928,N_22476,N_22059);
nor U22929 (N_22929,N_22162,N_21969);
or U22930 (N_22930,N_22366,N_22475);
nand U22931 (N_22931,N_22199,N_22121);
nor U22932 (N_22932,N_22225,N_22063);
nor U22933 (N_22933,N_22150,N_22425);
nor U22934 (N_22934,N_22449,N_22332);
or U22935 (N_22935,N_22249,N_22324);
nor U22936 (N_22936,N_22490,N_22190);
and U22937 (N_22937,N_22393,N_22426);
or U22938 (N_22938,N_22170,N_22164);
and U22939 (N_22939,N_22434,N_22224);
xor U22940 (N_22940,N_22397,N_22149);
nand U22941 (N_22941,N_22133,N_22391);
nor U22942 (N_22942,N_22117,N_22088);
xor U22943 (N_22943,N_22400,N_22381);
nor U22944 (N_22944,N_22040,N_22319);
or U22945 (N_22945,N_22462,N_22151);
xor U22946 (N_22946,N_22428,N_22287);
nor U22947 (N_22947,N_22222,N_22093);
nor U22948 (N_22948,N_22385,N_22125);
xor U22949 (N_22949,N_21939,N_22301);
and U22950 (N_22950,N_22441,N_22220);
xor U22951 (N_22951,N_21964,N_21991);
nor U22952 (N_22952,N_22404,N_22285);
nor U22953 (N_22953,N_21908,N_22081);
and U22954 (N_22954,N_22189,N_22055);
nor U22955 (N_22955,N_22373,N_22320);
nor U22956 (N_22956,N_22469,N_21922);
or U22957 (N_22957,N_21977,N_22110);
nand U22958 (N_22958,N_21909,N_21904);
nor U22959 (N_22959,N_22416,N_21959);
nand U22960 (N_22960,N_22339,N_21976);
or U22961 (N_22961,N_22045,N_22265);
and U22962 (N_22962,N_22170,N_22378);
nor U22963 (N_22963,N_22253,N_22365);
or U22964 (N_22964,N_22161,N_22121);
or U22965 (N_22965,N_22448,N_21887);
nor U22966 (N_22966,N_22481,N_22391);
xor U22967 (N_22967,N_22295,N_22053);
or U22968 (N_22968,N_22465,N_22234);
and U22969 (N_22969,N_22024,N_22169);
and U22970 (N_22970,N_22325,N_21908);
nand U22971 (N_22971,N_22153,N_22043);
or U22972 (N_22972,N_22095,N_22479);
and U22973 (N_22973,N_22209,N_22291);
and U22974 (N_22974,N_22448,N_22067);
or U22975 (N_22975,N_21915,N_22407);
and U22976 (N_22976,N_22036,N_21968);
nand U22977 (N_22977,N_21991,N_22338);
xnor U22978 (N_22978,N_22359,N_21976);
xor U22979 (N_22979,N_22327,N_21959);
nand U22980 (N_22980,N_22132,N_22413);
xnor U22981 (N_22981,N_22004,N_22423);
xnor U22982 (N_22982,N_22435,N_22469);
nand U22983 (N_22983,N_22280,N_22215);
xnor U22984 (N_22984,N_22111,N_22418);
nand U22985 (N_22985,N_22287,N_21998);
and U22986 (N_22986,N_22006,N_22211);
and U22987 (N_22987,N_22102,N_22167);
xor U22988 (N_22988,N_22273,N_22401);
and U22989 (N_22989,N_21904,N_21948);
or U22990 (N_22990,N_22470,N_22042);
xor U22991 (N_22991,N_22477,N_22181);
nand U22992 (N_22992,N_22058,N_22072);
or U22993 (N_22993,N_22293,N_22127);
nor U22994 (N_22994,N_22160,N_22245);
nor U22995 (N_22995,N_22261,N_22149);
nor U22996 (N_22996,N_22211,N_22465);
xor U22997 (N_22997,N_22224,N_22433);
xor U22998 (N_22998,N_22001,N_21913);
nor U22999 (N_22999,N_22086,N_22392);
xor U23000 (N_23000,N_22077,N_22337);
nor U23001 (N_23001,N_22111,N_21937);
nand U23002 (N_23002,N_22286,N_22224);
and U23003 (N_23003,N_22289,N_22121);
nor U23004 (N_23004,N_22008,N_22247);
nand U23005 (N_23005,N_22457,N_22111);
xnor U23006 (N_23006,N_22410,N_22063);
nor U23007 (N_23007,N_22170,N_22114);
nor U23008 (N_23008,N_21960,N_21907);
xnor U23009 (N_23009,N_22210,N_22469);
nor U23010 (N_23010,N_22166,N_22347);
nor U23011 (N_23011,N_22438,N_21963);
nor U23012 (N_23012,N_22356,N_21974);
nor U23013 (N_23013,N_22214,N_22112);
or U23014 (N_23014,N_22036,N_22070);
or U23015 (N_23015,N_21920,N_22430);
and U23016 (N_23016,N_22115,N_22360);
or U23017 (N_23017,N_22272,N_22042);
or U23018 (N_23018,N_21967,N_22410);
xor U23019 (N_23019,N_22073,N_22004);
nor U23020 (N_23020,N_22423,N_21914);
nand U23021 (N_23021,N_21945,N_22459);
nand U23022 (N_23022,N_22244,N_21930);
or U23023 (N_23023,N_21883,N_22129);
nor U23024 (N_23024,N_22007,N_22361);
nand U23025 (N_23025,N_21993,N_21970);
xor U23026 (N_23026,N_22200,N_21911);
xnor U23027 (N_23027,N_22418,N_21891);
nand U23028 (N_23028,N_22271,N_22077);
or U23029 (N_23029,N_22082,N_22381);
xnor U23030 (N_23030,N_22276,N_22139);
and U23031 (N_23031,N_22485,N_22162);
or U23032 (N_23032,N_22294,N_22063);
nand U23033 (N_23033,N_22096,N_21899);
or U23034 (N_23034,N_22392,N_22162);
or U23035 (N_23035,N_22347,N_22460);
nor U23036 (N_23036,N_22235,N_21998);
or U23037 (N_23037,N_22425,N_22049);
or U23038 (N_23038,N_22010,N_21995);
nand U23039 (N_23039,N_21880,N_22050);
nand U23040 (N_23040,N_21959,N_22469);
and U23041 (N_23041,N_22497,N_22270);
nand U23042 (N_23042,N_22010,N_22068);
nand U23043 (N_23043,N_21881,N_22199);
xnor U23044 (N_23044,N_22472,N_21883);
nand U23045 (N_23045,N_22408,N_21950);
xnor U23046 (N_23046,N_22284,N_21974);
nor U23047 (N_23047,N_22485,N_22450);
and U23048 (N_23048,N_21993,N_22117);
xnor U23049 (N_23049,N_22338,N_22399);
and U23050 (N_23050,N_22125,N_22232);
or U23051 (N_23051,N_22156,N_22445);
and U23052 (N_23052,N_22235,N_22254);
and U23053 (N_23053,N_21878,N_22070);
and U23054 (N_23054,N_21918,N_21987);
nor U23055 (N_23055,N_22445,N_22331);
and U23056 (N_23056,N_22479,N_22088);
xnor U23057 (N_23057,N_22095,N_22265);
and U23058 (N_23058,N_22243,N_22014);
or U23059 (N_23059,N_22228,N_22374);
xnor U23060 (N_23060,N_22470,N_22291);
xnor U23061 (N_23061,N_22199,N_21992);
nor U23062 (N_23062,N_22178,N_22291);
nor U23063 (N_23063,N_22373,N_21877);
nor U23064 (N_23064,N_22268,N_21875);
nand U23065 (N_23065,N_21960,N_22225);
nand U23066 (N_23066,N_22351,N_22265);
xor U23067 (N_23067,N_22325,N_22176);
and U23068 (N_23068,N_22123,N_22339);
nand U23069 (N_23069,N_22071,N_22437);
xnor U23070 (N_23070,N_22489,N_22074);
and U23071 (N_23071,N_22108,N_22146);
nand U23072 (N_23072,N_22473,N_22176);
or U23073 (N_23073,N_21938,N_21991);
or U23074 (N_23074,N_22131,N_22122);
and U23075 (N_23075,N_22072,N_22317);
and U23076 (N_23076,N_21901,N_22324);
nand U23077 (N_23077,N_22442,N_22443);
nor U23078 (N_23078,N_22220,N_22021);
nand U23079 (N_23079,N_22483,N_22175);
and U23080 (N_23080,N_22042,N_22180);
xor U23081 (N_23081,N_22331,N_22181);
or U23082 (N_23082,N_22123,N_22131);
xnor U23083 (N_23083,N_22308,N_22266);
nand U23084 (N_23084,N_21920,N_21915);
xor U23085 (N_23085,N_22430,N_22265);
and U23086 (N_23086,N_22053,N_22037);
or U23087 (N_23087,N_22300,N_22421);
or U23088 (N_23088,N_22091,N_22417);
nor U23089 (N_23089,N_22311,N_22211);
or U23090 (N_23090,N_21952,N_22372);
or U23091 (N_23091,N_22337,N_22050);
nand U23092 (N_23092,N_22120,N_21952);
nor U23093 (N_23093,N_22429,N_22498);
and U23094 (N_23094,N_21945,N_22012);
and U23095 (N_23095,N_22256,N_22142);
nand U23096 (N_23096,N_22049,N_21972);
or U23097 (N_23097,N_22322,N_22294);
or U23098 (N_23098,N_22470,N_22414);
xor U23099 (N_23099,N_22132,N_22143);
nor U23100 (N_23100,N_22182,N_21928);
or U23101 (N_23101,N_21947,N_22237);
or U23102 (N_23102,N_22396,N_22013);
nor U23103 (N_23103,N_22431,N_22185);
nor U23104 (N_23104,N_22113,N_22297);
or U23105 (N_23105,N_21906,N_22020);
nor U23106 (N_23106,N_22385,N_22414);
nand U23107 (N_23107,N_22044,N_22414);
nor U23108 (N_23108,N_22013,N_22403);
nor U23109 (N_23109,N_21933,N_22393);
xor U23110 (N_23110,N_22273,N_22175);
nor U23111 (N_23111,N_22254,N_22161);
nand U23112 (N_23112,N_22334,N_21912);
or U23113 (N_23113,N_22214,N_22043);
nand U23114 (N_23114,N_22028,N_22088);
nand U23115 (N_23115,N_22424,N_22066);
nor U23116 (N_23116,N_22256,N_22287);
nand U23117 (N_23117,N_22490,N_21991);
or U23118 (N_23118,N_22422,N_21957);
nand U23119 (N_23119,N_22019,N_22474);
xnor U23120 (N_23120,N_22242,N_22197);
xnor U23121 (N_23121,N_22094,N_22305);
nand U23122 (N_23122,N_22226,N_22362);
nor U23123 (N_23123,N_22274,N_22270);
or U23124 (N_23124,N_21881,N_22375);
xor U23125 (N_23125,N_22673,N_22732);
and U23126 (N_23126,N_22517,N_22640);
and U23127 (N_23127,N_22511,N_22837);
xnor U23128 (N_23128,N_23008,N_22576);
and U23129 (N_23129,N_23052,N_22868);
or U23130 (N_23130,N_22674,N_22928);
nand U23131 (N_23131,N_22643,N_22892);
and U23132 (N_23132,N_22555,N_22735);
nor U23133 (N_23133,N_22636,N_23030);
and U23134 (N_23134,N_22639,N_22951);
nand U23135 (N_23135,N_22687,N_23070);
nor U23136 (N_23136,N_22904,N_22948);
xnor U23137 (N_23137,N_22574,N_22535);
xnor U23138 (N_23138,N_22572,N_23087);
nor U23139 (N_23139,N_22608,N_23000);
nand U23140 (N_23140,N_23073,N_22693);
xor U23141 (N_23141,N_22896,N_23090);
nand U23142 (N_23142,N_22558,N_22692);
nand U23143 (N_23143,N_22884,N_22723);
or U23144 (N_23144,N_22831,N_22520);
and U23145 (N_23145,N_23033,N_23044);
nand U23146 (N_23146,N_22568,N_22798);
and U23147 (N_23147,N_23049,N_22720);
nand U23148 (N_23148,N_23025,N_22669);
and U23149 (N_23149,N_23048,N_22654);
nand U23150 (N_23150,N_22626,N_23115);
and U23151 (N_23151,N_23078,N_22695);
xor U23152 (N_23152,N_23014,N_23076);
and U23153 (N_23153,N_23060,N_22995);
nand U23154 (N_23154,N_22706,N_23036);
and U23155 (N_23155,N_22953,N_22502);
nand U23156 (N_23156,N_22570,N_23081);
xnor U23157 (N_23157,N_22908,N_22856);
xnor U23158 (N_23158,N_22834,N_22738);
and U23159 (N_23159,N_22665,N_22997);
and U23160 (N_23160,N_22657,N_22745);
nand U23161 (N_23161,N_23040,N_22854);
and U23162 (N_23162,N_22623,N_23056);
xnor U23163 (N_23163,N_22552,N_22905);
nor U23164 (N_23164,N_22697,N_23028);
nor U23165 (N_23165,N_22785,N_22685);
nor U23166 (N_23166,N_22596,N_22719);
and U23167 (N_23167,N_22542,N_22755);
and U23168 (N_23168,N_22569,N_22959);
xnor U23169 (N_23169,N_22726,N_23019);
or U23170 (N_23170,N_22603,N_22514);
or U23171 (N_23171,N_22763,N_22510);
nor U23172 (N_23172,N_22847,N_22686);
xor U23173 (N_23173,N_23006,N_22938);
or U23174 (N_23174,N_22939,N_22593);
xnor U23175 (N_23175,N_22714,N_22614);
nand U23176 (N_23176,N_22747,N_22800);
and U23177 (N_23177,N_22507,N_23102);
xor U23178 (N_23178,N_22897,N_23041);
and U23179 (N_23179,N_23082,N_22870);
xnor U23180 (N_23180,N_22950,N_23086);
or U23181 (N_23181,N_22586,N_22575);
and U23182 (N_23182,N_22887,N_22820);
nand U23183 (N_23183,N_22590,N_23035);
or U23184 (N_23184,N_22671,N_22838);
and U23185 (N_23185,N_22547,N_22979);
and U23186 (N_23186,N_22795,N_22606);
nor U23187 (N_23187,N_22543,N_22787);
or U23188 (N_23188,N_22935,N_22779);
nor U23189 (N_23189,N_22810,N_23106);
and U23190 (N_23190,N_22923,N_22754);
nand U23191 (N_23191,N_22956,N_22961);
xor U23192 (N_23192,N_22528,N_23047);
or U23193 (N_23193,N_22728,N_22529);
nor U23194 (N_23194,N_22781,N_22925);
xnor U23195 (N_23195,N_22522,N_22663);
and U23196 (N_23196,N_23109,N_22912);
and U23197 (N_23197,N_22610,N_23095);
nor U23198 (N_23198,N_22734,N_23072);
or U23199 (N_23199,N_22545,N_22962);
nand U23200 (N_23200,N_22906,N_22767);
or U23201 (N_23201,N_22599,N_22913);
nand U23202 (N_23202,N_22773,N_22981);
nand U23203 (N_23203,N_22984,N_22952);
and U23204 (N_23204,N_22790,N_22611);
nor U23205 (N_23205,N_23009,N_22698);
nand U23206 (N_23206,N_22597,N_22613);
or U23207 (N_23207,N_22667,N_22982);
nand U23208 (N_23208,N_22716,N_22818);
nor U23209 (N_23209,N_22877,N_22554);
or U23210 (N_23210,N_22889,N_22929);
nand U23211 (N_23211,N_22607,N_22677);
or U23212 (N_23212,N_23005,N_22565);
nor U23213 (N_23213,N_23007,N_22624);
nor U23214 (N_23214,N_22777,N_22770);
nor U23215 (N_23215,N_22827,N_22993);
nor U23216 (N_23216,N_22646,N_22530);
nand U23217 (N_23217,N_22976,N_22942);
nand U23218 (N_23218,N_22805,N_22855);
xnor U23219 (N_23219,N_22524,N_22821);
or U23220 (N_23220,N_22762,N_22516);
nor U23221 (N_23221,N_23031,N_22653);
nand U23222 (N_23222,N_22825,N_22650);
or U23223 (N_23223,N_22937,N_22883);
xor U23224 (N_23224,N_22644,N_22869);
nand U23225 (N_23225,N_22743,N_23004);
and U23226 (N_23226,N_23020,N_22722);
or U23227 (N_23227,N_22562,N_22771);
and U23228 (N_23228,N_22751,N_22915);
and U23229 (N_23229,N_22927,N_22512);
nor U23230 (N_23230,N_23043,N_22843);
nor U23231 (N_23231,N_22591,N_22801);
or U23232 (N_23232,N_23037,N_23021);
nand U23233 (N_23233,N_22642,N_23124);
and U23234 (N_23234,N_22954,N_23069);
nor U23235 (N_23235,N_22721,N_22679);
xnor U23236 (N_23236,N_23108,N_22595);
and U23237 (N_23237,N_22753,N_22963);
or U23238 (N_23238,N_23023,N_22811);
nand U23239 (N_23239,N_22957,N_22660);
and U23240 (N_23240,N_22824,N_23061);
or U23241 (N_23241,N_22534,N_22578);
and U23242 (N_23242,N_23075,N_23071);
and U23243 (N_23243,N_22668,N_22794);
xnor U23244 (N_23244,N_22849,N_22983);
nand U23245 (N_23245,N_22619,N_22740);
xor U23246 (N_23246,N_22598,N_22560);
nor U23247 (N_23247,N_22876,N_22713);
nand U23248 (N_23248,N_22901,N_23114);
nor U23249 (N_23249,N_22826,N_22500);
or U23250 (N_23250,N_22752,N_23015);
or U23251 (N_23251,N_22622,N_23107);
and U23252 (N_23252,N_23074,N_22823);
xnor U23253 (N_23253,N_22866,N_22549);
or U23254 (N_23254,N_22909,N_22916);
or U23255 (N_23255,N_22756,N_23013);
nor U23256 (N_23256,N_22830,N_22631);
and U23257 (N_23257,N_23116,N_22689);
or U23258 (N_23258,N_22617,N_22947);
nand U23259 (N_23259,N_22899,N_22969);
and U23260 (N_23260,N_23120,N_22509);
or U23261 (N_23261,N_22550,N_22975);
and U23262 (N_23262,N_23017,N_22583);
or U23263 (N_23263,N_22691,N_22998);
nor U23264 (N_23264,N_23010,N_22731);
nor U23265 (N_23265,N_22955,N_23066);
and U23266 (N_23266,N_23022,N_22638);
and U23267 (N_23267,N_22637,N_22532);
xnor U23268 (N_23268,N_22835,N_22605);
or U23269 (N_23269,N_22725,N_22661);
nor U23270 (N_23270,N_22531,N_22612);
nor U23271 (N_23271,N_22807,N_22885);
and U23272 (N_23272,N_22793,N_22840);
nor U23273 (N_23273,N_22678,N_22737);
xnor U23274 (N_23274,N_22965,N_22662);
nor U23275 (N_23275,N_22609,N_22933);
nand U23276 (N_23276,N_22898,N_22601);
nand U23277 (N_23277,N_22921,N_22633);
nand U23278 (N_23278,N_23117,N_22635);
nand U23279 (N_23279,N_23092,N_22527);
or U23280 (N_23280,N_22733,N_22804);
nor U23281 (N_23281,N_22513,N_23059);
or U23282 (N_23282,N_22924,N_22776);
and U23283 (N_23283,N_22836,N_22708);
and U23284 (N_23284,N_22778,N_22974);
nand U23285 (N_23285,N_23085,N_22658);
or U23286 (N_23286,N_22567,N_22628);
and U23287 (N_23287,N_22627,N_22594);
or U23288 (N_23288,N_22880,N_22920);
xor U23289 (N_23289,N_23026,N_23012);
nor U23290 (N_23290,N_22703,N_22931);
nand U23291 (N_23291,N_22645,N_22602);
nor U23292 (N_23292,N_22649,N_22544);
and U23293 (N_23293,N_22707,N_22515);
or U23294 (N_23294,N_22682,N_22537);
xor U23295 (N_23295,N_22799,N_22985);
nand U23296 (N_23296,N_22676,N_22651);
and U23297 (N_23297,N_23062,N_23110);
and U23298 (N_23298,N_22742,N_22988);
and U23299 (N_23299,N_22540,N_22964);
and U23300 (N_23300,N_22729,N_22848);
nor U23301 (N_23301,N_22859,N_22875);
xnor U23302 (N_23302,N_22618,N_22699);
and U23303 (N_23303,N_22978,N_22566);
and U23304 (N_23304,N_22715,N_22630);
or U23305 (N_23305,N_22766,N_22894);
xor U23306 (N_23306,N_23118,N_22992);
nor U23307 (N_23307,N_22744,N_22816);
nor U23308 (N_23308,N_22914,N_22621);
nor U23309 (N_23309,N_22863,N_22629);
nand U23310 (N_23310,N_22541,N_23084);
nor U23311 (N_23311,N_22521,N_22930);
nand U23312 (N_23312,N_22919,N_22768);
and U23313 (N_23313,N_22700,N_22705);
nor U23314 (N_23314,N_22775,N_23089);
and U23315 (N_23315,N_22760,N_22796);
nand U23316 (N_23316,N_22881,N_23098);
nand U23317 (N_23317,N_22943,N_22806);
nand U23318 (N_23318,N_22553,N_22783);
xor U23319 (N_23319,N_22519,N_22862);
and U23320 (N_23320,N_22846,N_22970);
nor U23321 (N_23321,N_22971,N_23053);
xor U23322 (N_23322,N_22815,N_22926);
xor U23323 (N_23323,N_22579,N_22585);
nor U23324 (N_23324,N_23101,N_22758);
nand U23325 (N_23325,N_22791,N_22874);
or U23326 (N_23326,N_22886,N_22973);
nand U23327 (N_23327,N_23080,N_23119);
nor U23328 (N_23328,N_22803,N_23051);
or U23329 (N_23329,N_22844,N_22523);
and U23330 (N_23330,N_22890,N_22994);
nand U23331 (N_23331,N_22587,N_22871);
and U23332 (N_23332,N_22584,N_22556);
or U23333 (N_23333,N_22563,N_22538);
and U23334 (N_23334,N_22533,N_23046);
xnor U23335 (N_23335,N_22911,N_22839);
or U23336 (N_23336,N_22893,N_22809);
xnor U23337 (N_23337,N_22941,N_22864);
xor U23338 (N_23338,N_23094,N_23097);
xor U23339 (N_23339,N_22501,N_22526);
or U23340 (N_23340,N_22967,N_22694);
and U23341 (N_23341,N_23122,N_23003);
and U23342 (N_23342,N_22832,N_22504);
or U23343 (N_23343,N_22548,N_23029);
or U23344 (N_23344,N_23100,N_22666);
nor U23345 (N_23345,N_22784,N_22764);
and U23346 (N_23346,N_22891,N_22940);
or U23347 (N_23347,N_22739,N_22882);
xor U23348 (N_23348,N_22902,N_23039);
or U23349 (N_23349,N_22748,N_22918);
xor U23350 (N_23350,N_22684,N_22681);
nor U23351 (N_23351,N_22680,N_23016);
or U23352 (N_23352,N_22865,N_22505);
nand U23353 (N_23353,N_22960,N_22972);
xnor U23354 (N_23354,N_22711,N_23091);
and U23355 (N_23355,N_22712,N_22852);
xnor U23356 (N_23356,N_23055,N_23032);
and U23357 (N_23357,N_22945,N_22620);
xnor U23358 (N_23358,N_23042,N_22616);
nand U23359 (N_23359,N_23105,N_22503);
nand U23360 (N_23360,N_22564,N_22727);
nand U23361 (N_23361,N_22656,N_23099);
xnor U23362 (N_23362,N_22808,N_23093);
nor U23363 (N_23363,N_22996,N_22858);
or U23364 (N_23364,N_22861,N_22750);
or U23365 (N_23365,N_22842,N_22857);
or U23366 (N_23366,N_22683,N_23123);
nand U23367 (N_23367,N_23018,N_22625);
or U23368 (N_23368,N_22772,N_23096);
nand U23369 (N_23369,N_22670,N_22652);
nand U23370 (N_23370,N_22573,N_23027);
nor U23371 (N_23371,N_22710,N_23104);
nor U23372 (N_23372,N_22990,N_22724);
nand U23373 (N_23373,N_22508,N_22592);
xnor U23374 (N_23374,N_22581,N_22910);
nand U23375 (N_23375,N_22802,N_23067);
nor U23376 (N_23376,N_22765,N_22934);
and U23377 (N_23377,N_23054,N_22814);
nor U23378 (N_23378,N_22786,N_22717);
nand U23379 (N_23379,N_22949,N_22632);
or U23380 (N_23380,N_22518,N_22819);
nand U23381 (N_23381,N_23079,N_22980);
and U23382 (N_23382,N_22966,N_22917);
nor U23383 (N_23383,N_22696,N_22944);
and U23384 (N_23384,N_23083,N_22506);
or U23385 (N_23385,N_22539,N_22853);
and U23386 (N_23386,N_22780,N_22741);
and U23387 (N_23387,N_22664,N_22690);
or U23388 (N_23388,N_22648,N_23050);
nor U23389 (N_23389,N_22907,N_23045);
or U23390 (N_23390,N_22672,N_22888);
or U23391 (N_23391,N_22525,N_22789);
and U23392 (N_23392,N_22936,N_22987);
nand U23393 (N_23393,N_22873,N_23002);
and U23394 (N_23394,N_22851,N_23063);
nor U23395 (N_23395,N_23111,N_22577);
nor U23396 (N_23396,N_23077,N_22932);
nand U23397 (N_23397,N_22788,N_22561);
xor U23398 (N_23398,N_22647,N_22817);
or U23399 (N_23399,N_22782,N_22958);
and U23400 (N_23400,N_22774,N_22655);
or U23401 (N_23401,N_23011,N_22641);
and U23402 (N_23402,N_22833,N_22536);
nor U23403 (N_23403,N_23057,N_22588);
and U23404 (N_23404,N_23113,N_22850);
and U23405 (N_23405,N_22895,N_22769);
or U23406 (N_23406,N_22559,N_22999);
xnor U23407 (N_23407,N_22709,N_22986);
nor U23408 (N_23408,N_22659,N_22946);
nand U23409 (N_23409,N_23065,N_22977);
nand U23410 (N_23410,N_22600,N_22792);
xor U23411 (N_23411,N_22878,N_22604);
nor U23412 (N_23412,N_22730,N_22812);
nor U23413 (N_23413,N_22828,N_23121);
and U23414 (N_23414,N_22867,N_22872);
nor U23415 (N_23415,N_22841,N_22702);
nor U23416 (N_23416,N_22991,N_22582);
xnor U23417 (N_23417,N_22845,N_22900);
or U23418 (N_23418,N_23024,N_22989);
and U23419 (N_23419,N_23038,N_22571);
nand U23420 (N_23420,N_22615,N_22589);
xnor U23421 (N_23421,N_23058,N_23034);
nor U23422 (N_23422,N_22718,N_22546);
nor U23423 (N_23423,N_22879,N_22903);
nor U23424 (N_23424,N_22736,N_22675);
nor U23425 (N_23425,N_22704,N_23064);
and U23426 (N_23426,N_23001,N_22749);
and U23427 (N_23427,N_22813,N_22759);
or U23428 (N_23428,N_22701,N_22797);
or U23429 (N_23429,N_22968,N_22922);
and U23430 (N_23430,N_22757,N_22761);
nand U23431 (N_23431,N_22829,N_22634);
and U23432 (N_23432,N_22860,N_23103);
nor U23433 (N_23433,N_22580,N_23068);
nand U23434 (N_23434,N_22746,N_22822);
or U23435 (N_23435,N_22557,N_23112);
nand U23436 (N_23436,N_22688,N_22551);
xor U23437 (N_23437,N_23088,N_23115);
nor U23438 (N_23438,N_23074,N_22587);
xor U23439 (N_23439,N_22690,N_22863);
nand U23440 (N_23440,N_22882,N_22968);
or U23441 (N_23441,N_22539,N_23109);
and U23442 (N_23442,N_23049,N_22887);
nor U23443 (N_23443,N_22727,N_22534);
and U23444 (N_23444,N_22900,N_22698);
or U23445 (N_23445,N_22988,N_22832);
xnor U23446 (N_23446,N_22809,N_22930);
xor U23447 (N_23447,N_22782,N_22898);
or U23448 (N_23448,N_23010,N_22533);
nor U23449 (N_23449,N_23123,N_22634);
nor U23450 (N_23450,N_22723,N_22977);
nor U23451 (N_23451,N_22684,N_22996);
or U23452 (N_23452,N_22909,N_23027);
nor U23453 (N_23453,N_23110,N_23042);
xnor U23454 (N_23454,N_22709,N_22973);
nand U23455 (N_23455,N_22902,N_22908);
and U23456 (N_23456,N_22724,N_22968);
nor U23457 (N_23457,N_22859,N_22516);
and U23458 (N_23458,N_22745,N_22623);
or U23459 (N_23459,N_23091,N_23013);
nor U23460 (N_23460,N_22670,N_22865);
xor U23461 (N_23461,N_22954,N_22613);
nand U23462 (N_23462,N_22510,N_23105);
nand U23463 (N_23463,N_22757,N_23093);
xor U23464 (N_23464,N_22653,N_22912);
nor U23465 (N_23465,N_22656,N_22937);
xnor U23466 (N_23466,N_22568,N_22522);
and U23467 (N_23467,N_22852,N_22798);
nor U23468 (N_23468,N_23002,N_22556);
nor U23469 (N_23469,N_23078,N_22950);
and U23470 (N_23470,N_23037,N_22651);
and U23471 (N_23471,N_23061,N_22796);
and U23472 (N_23472,N_22820,N_22712);
or U23473 (N_23473,N_22535,N_22615);
nor U23474 (N_23474,N_22537,N_22508);
nor U23475 (N_23475,N_22578,N_22802);
nor U23476 (N_23476,N_22698,N_22873);
and U23477 (N_23477,N_22785,N_22953);
xor U23478 (N_23478,N_22587,N_22900);
or U23479 (N_23479,N_22768,N_23103);
nor U23480 (N_23480,N_23009,N_23034);
or U23481 (N_23481,N_22951,N_22914);
or U23482 (N_23482,N_22725,N_22693);
and U23483 (N_23483,N_22942,N_22800);
nand U23484 (N_23484,N_23085,N_22685);
nand U23485 (N_23485,N_22670,N_22626);
and U23486 (N_23486,N_22685,N_22933);
or U23487 (N_23487,N_22725,N_22720);
and U23488 (N_23488,N_22769,N_22521);
nor U23489 (N_23489,N_22523,N_22605);
or U23490 (N_23490,N_22676,N_22885);
nand U23491 (N_23491,N_22586,N_22527);
nor U23492 (N_23492,N_22684,N_22712);
nand U23493 (N_23493,N_22978,N_22571);
nor U23494 (N_23494,N_22721,N_22601);
nor U23495 (N_23495,N_22708,N_22585);
or U23496 (N_23496,N_22841,N_23043);
and U23497 (N_23497,N_22518,N_22561);
xor U23498 (N_23498,N_22660,N_23048);
or U23499 (N_23499,N_23022,N_22814);
nand U23500 (N_23500,N_23005,N_22822);
nand U23501 (N_23501,N_22667,N_22783);
nor U23502 (N_23502,N_23052,N_22979);
xnor U23503 (N_23503,N_22848,N_23033);
and U23504 (N_23504,N_23021,N_22958);
nor U23505 (N_23505,N_22796,N_22698);
nand U23506 (N_23506,N_22508,N_22824);
and U23507 (N_23507,N_23085,N_22892);
nand U23508 (N_23508,N_22515,N_22640);
nand U23509 (N_23509,N_22628,N_22995);
nand U23510 (N_23510,N_22857,N_23103);
nor U23511 (N_23511,N_22690,N_23009);
xor U23512 (N_23512,N_22814,N_22558);
xnor U23513 (N_23513,N_22851,N_22898);
xnor U23514 (N_23514,N_23124,N_23025);
and U23515 (N_23515,N_22725,N_22953);
and U23516 (N_23516,N_22994,N_22766);
nand U23517 (N_23517,N_23005,N_22885);
and U23518 (N_23518,N_23085,N_22618);
nand U23519 (N_23519,N_22524,N_22755);
or U23520 (N_23520,N_23065,N_23096);
nand U23521 (N_23521,N_23047,N_22686);
and U23522 (N_23522,N_22992,N_22503);
or U23523 (N_23523,N_22933,N_22832);
nor U23524 (N_23524,N_22529,N_22646);
nor U23525 (N_23525,N_22817,N_22890);
nor U23526 (N_23526,N_22781,N_22718);
or U23527 (N_23527,N_23082,N_22970);
nand U23528 (N_23528,N_22805,N_22596);
and U23529 (N_23529,N_22852,N_22607);
nand U23530 (N_23530,N_22961,N_22593);
nand U23531 (N_23531,N_22974,N_22786);
and U23532 (N_23532,N_22700,N_23102);
nor U23533 (N_23533,N_22531,N_22924);
nand U23534 (N_23534,N_22968,N_22584);
and U23535 (N_23535,N_22601,N_22823);
nand U23536 (N_23536,N_23051,N_23041);
nor U23537 (N_23537,N_22583,N_22584);
nor U23538 (N_23538,N_22643,N_22628);
and U23539 (N_23539,N_22656,N_22508);
xor U23540 (N_23540,N_22872,N_22865);
or U23541 (N_23541,N_22537,N_22670);
nor U23542 (N_23542,N_23023,N_22775);
and U23543 (N_23543,N_23031,N_22555);
or U23544 (N_23544,N_23056,N_22528);
or U23545 (N_23545,N_22974,N_22699);
and U23546 (N_23546,N_22554,N_22881);
nand U23547 (N_23547,N_22963,N_22569);
and U23548 (N_23548,N_22740,N_22734);
or U23549 (N_23549,N_22897,N_22875);
or U23550 (N_23550,N_22770,N_22790);
nor U23551 (N_23551,N_22565,N_22766);
or U23552 (N_23552,N_22587,N_22995);
nand U23553 (N_23553,N_23034,N_22922);
xnor U23554 (N_23554,N_23103,N_22909);
xnor U23555 (N_23555,N_22737,N_23091);
and U23556 (N_23556,N_22712,N_22830);
nor U23557 (N_23557,N_22778,N_22978);
and U23558 (N_23558,N_22668,N_22717);
xor U23559 (N_23559,N_22826,N_22607);
nand U23560 (N_23560,N_22920,N_22738);
nor U23561 (N_23561,N_23104,N_22934);
nand U23562 (N_23562,N_22907,N_23015);
nand U23563 (N_23563,N_22633,N_23003);
nor U23564 (N_23564,N_22647,N_22829);
or U23565 (N_23565,N_23028,N_22561);
or U23566 (N_23566,N_22578,N_22671);
and U23567 (N_23567,N_22792,N_22817);
or U23568 (N_23568,N_22933,N_23044);
nor U23569 (N_23569,N_22834,N_22687);
or U23570 (N_23570,N_22622,N_22950);
or U23571 (N_23571,N_22830,N_23001);
or U23572 (N_23572,N_22638,N_22662);
nor U23573 (N_23573,N_22539,N_22564);
nand U23574 (N_23574,N_22817,N_22829);
nor U23575 (N_23575,N_23066,N_23097);
nor U23576 (N_23576,N_22962,N_22579);
or U23577 (N_23577,N_22536,N_22963);
nor U23578 (N_23578,N_22752,N_23054);
nand U23579 (N_23579,N_23009,N_22884);
xnor U23580 (N_23580,N_22939,N_23102);
nor U23581 (N_23581,N_23124,N_22884);
or U23582 (N_23582,N_22764,N_22881);
or U23583 (N_23583,N_22922,N_23116);
xnor U23584 (N_23584,N_22733,N_23092);
nand U23585 (N_23585,N_22524,N_22939);
nand U23586 (N_23586,N_23086,N_22681);
and U23587 (N_23587,N_23093,N_22695);
nor U23588 (N_23588,N_22966,N_22585);
xor U23589 (N_23589,N_22638,N_22969);
or U23590 (N_23590,N_22626,N_23013);
nor U23591 (N_23591,N_23071,N_23121);
and U23592 (N_23592,N_22857,N_22568);
nor U23593 (N_23593,N_22533,N_22528);
and U23594 (N_23594,N_22704,N_22864);
nor U23595 (N_23595,N_23054,N_22599);
xnor U23596 (N_23596,N_22744,N_22903);
and U23597 (N_23597,N_22765,N_22906);
or U23598 (N_23598,N_22585,N_22752);
nor U23599 (N_23599,N_22714,N_22766);
nand U23600 (N_23600,N_22732,N_22966);
and U23601 (N_23601,N_22961,N_22509);
nand U23602 (N_23602,N_22560,N_23039);
and U23603 (N_23603,N_22684,N_23011);
nor U23604 (N_23604,N_23083,N_22836);
xor U23605 (N_23605,N_22890,N_22979);
nor U23606 (N_23606,N_22965,N_22664);
or U23607 (N_23607,N_22609,N_22611);
nor U23608 (N_23608,N_22551,N_22763);
nand U23609 (N_23609,N_22612,N_22924);
nand U23610 (N_23610,N_23051,N_22617);
nand U23611 (N_23611,N_22824,N_22628);
and U23612 (N_23612,N_22949,N_22705);
nor U23613 (N_23613,N_23018,N_22582);
xor U23614 (N_23614,N_22954,N_22748);
or U23615 (N_23615,N_22575,N_22911);
nor U23616 (N_23616,N_23014,N_22652);
xnor U23617 (N_23617,N_22765,N_22584);
xor U23618 (N_23618,N_22914,N_23024);
xor U23619 (N_23619,N_22902,N_22895);
xor U23620 (N_23620,N_22616,N_22585);
and U23621 (N_23621,N_22544,N_23097);
or U23622 (N_23622,N_23112,N_23008);
and U23623 (N_23623,N_23064,N_22718);
nor U23624 (N_23624,N_22999,N_23059);
xnor U23625 (N_23625,N_22732,N_22584);
or U23626 (N_23626,N_23007,N_23015);
and U23627 (N_23627,N_22930,N_22886);
and U23628 (N_23628,N_22834,N_22920);
or U23629 (N_23629,N_23039,N_22608);
xnor U23630 (N_23630,N_22588,N_22713);
xor U23631 (N_23631,N_22999,N_22692);
or U23632 (N_23632,N_22864,N_22723);
or U23633 (N_23633,N_22685,N_22802);
xnor U23634 (N_23634,N_22877,N_23121);
and U23635 (N_23635,N_23094,N_22868);
nand U23636 (N_23636,N_22629,N_22507);
and U23637 (N_23637,N_22927,N_22887);
nor U23638 (N_23638,N_22949,N_22924);
or U23639 (N_23639,N_23014,N_22861);
xor U23640 (N_23640,N_22661,N_23091);
and U23641 (N_23641,N_22996,N_22973);
nand U23642 (N_23642,N_23080,N_22726);
nor U23643 (N_23643,N_22637,N_22515);
nor U23644 (N_23644,N_22734,N_22613);
or U23645 (N_23645,N_22690,N_22931);
nor U23646 (N_23646,N_22954,N_22736);
and U23647 (N_23647,N_22919,N_22748);
nand U23648 (N_23648,N_22881,N_22997);
and U23649 (N_23649,N_22886,N_22965);
or U23650 (N_23650,N_22772,N_22581);
nor U23651 (N_23651,N_23002,N_22803);
or U23652 (N_23652,N_22725,N_22858);
xor U23653 (N_23653,N_23057,N_22670);
nand U23654 (N_23654,N_22655,N_22798);
and U23655 (N_23655,N_22926,N_22708);
nand U23656 (N_23656,N_22952,N_22672);
nand U23657 (N_23657,N_23102,N_22512);
and U23658 (N_23658,N_22797,N_22688);
xnor U23659 (N_23659,N_22895,N_22738);
or U23660 (N_23660,N_22651,N_22956);
xnor U23661 (N_23661,N_22769,N_22944);
or U23662 (N_23662,N_22656,N_22533);
xnor U23663 (N_23663,N_22912,N_22810);
nor U23664 (N_23664,N_22882,N_22896);
or U23665 (N_23665,N_23071,N_22910);
nor U23666 (N_23666,N_22850,N_22813);
nor U23667 (N_23667,N_22933,N_22998);
nor U23668 (N_23668,N_22962,N_22665);
nand U23669 (N_23669,N_22726,N_22730);
nand U23670 (N_23670,N_22622,N_22945);
nor U23671 (N_23671,N_22944,N_22908);
xor U23672 (N_23672,N_22966,N_22972);
or U23673 (N_23673,N_22600,N_22807);
nand U23674 (N_23674,N_22849,N_22818);
nand U23675 (N_23675,N_23065,N_23103);
xnor U23676 (N_23676,N_22854,N_22544);
and U23677 (N_23677,N_22510,N_22775);
nand U23678 (N_23678,N_23001,N_22751);
or U23679 (N_23679,N_22695,N_23051);
nor U23680 (N_23680,N_22629,N_22792);
xnor U23681 (N_23681,N_22869,N_22940);
and U23682 (N_23682,N_23122,N_22945);
nand U23683 (N_23683,N_22823,N_22684);
nand U23684 (N_23684,N_22806,N_22780);
nand U23685 (N_23685,N_22636,N_22926);
nand U23686 (N_23686,N_22679,N_22920);
and U23687 (N_23687,N_22701,N_22500);
or U23688 (N_23688,N_23028,N_22623);
nand U23689 (N_23689,N_22828,N_22911);
xor U23690 (N_23690,N_23122,N_22828);
and U23691 (N_23691,N_23086,N_22695);
and U23692 (N_23692,N_22649,N_22993);
and U23693 (N_23693,N_22665,N_22989);
nor U23694 (N_23694,N_22803,N_22770);
and U23695 (N_23695,N_22759,N_22935);
nor U23696 (N_23696,N_22630,N_22866);
nand U23697 (N_23697,N_23056,N_22773);
or U23698 (N_23698,N_22869,N_22654);
xor U23699 (N_23699,N_22895,N_22882);
or U23700 (N_23700,N_23053,N_22554);
or U23701 (N_23701,N_22912,N_22648);
and U23702 (N_23702,N_22980,N_22558);
nand U23703 (N_23703,N_23069,N_22952);
or U23704 (N_23704,N_23022,N_22568);
or U23705 (N_23705,N_22550,N_22627);
nor U23706 (N_23706,N_22992,N_22597);
and U23707 (N_23707,N_22741,N_22878);
or U23708 (N_23708,N_23124,N_22817);
nand U23709 (N_23709,N_22551,N_22848);
nor U23710 (N_23710,N_22708,N_22713);
and U23711 (N_23711,N_22923,N_23022);
nor U23712 (N_23712,N_23024,N_22529);
xor U23713 (N_23713,N_22985,N_22573);
or U23714 (N_23714,N_22705,N_22643);
xor U23715 (N_23715,N_22638,N_22706);
nor U23716 (N_23716,N_22826,N_22735);
xnor U23717 (N_23717,N_22788,N_22785);
nor U23718 (N_23718,N_22530,N_23005);
xnor U23719 (N_23719,N_22545,N_23021);
or U23720 (N_23720,N_22895,N_22889);
nand U23721 (N_23721,N_22865,N_22577);
nor U23722 (N_23722,N_23002,N_23005);
nor U23723 (N_23723,N_22685,N_22623);
nor U23724 (N_23724,N_23111,N_22613);
or U23725 (N_23725,N_23014,N_22553);
nand U23726 (N_23726,N_22567,N_22671);
nand U23727 (N_23727,N_22514,N_22874);
and U23728 (N_23728,N_22828,N_22694);
or U23729 (N_23729,N_22893,N_22927);
xor U23730 (N_23730,N_22591,N_22523);
nor U23731 (N_23731,N_22771,N_22844);
or U23732 (N_23732,N_22641,N_23088);
or U23733 (N_23733,N_22979,N_23092);
and U23734 (N_23734,N_22532,N_22947);
xor U23735 (N_23735,N_22950,N_22921);
or U23736 (N_23736,N_22930,N_22953);
nor U23737 (N_23737,N_22660,N_22662);
xnor U23738 (N_23738,N_22750,N_22962);
and U23739 (N_23739,N_23053,N_22504);
nand U23740 (N_23740,N_22520,N_23027);
and U23741 (N_23741,N_22943,N_22884);
nand U23742 (N_23742,N_23045,N_22996);
xor U23743 (N_23743,N_22977,N_23071);
or U23744 (N_23744,N_22826,N_22935);
and U23745 (N_23745,N_22751,N_22649);
or U23746 (N_23746,N_22999,N_22763);
and U23747 (N_23747,N_22656,N_22810);
or U23748 (N_23748,N_22803,N_22936);
nor U23749 (N_23749,N_22717,N_23048);
xor U23750 (N_23750,N_23160,N_23282);
nand U23751 (N_23751,N_23157,N_23129);
and U23752 (N_23752,N_23605,N_23274);
nor U23753 (N_23753,N_23668,N_23465);
and U23754 (N_23754,N_23429,N_23587);
nand U23755 (N_23755,N_23232,N_23151);
or U23756 (N_23756,N_23171,N_23264);
or U23757 (N_23757,N_23502,N_23571);
xnor U23758 (N_23758,N_23165,N_23213);
and U23759 (N_23759,N_23442,N_23545);
xor U23760 (N_23760,N_23435,N_23714);
xor U23761 (N_23761,N_23309,N_23567);
and U23762 (N_23762,N_23632,N_23402);
or U23763 (N_23763,N_23494,N_23734);
xor U23764 (N_23764,N_23425,N_23622);
nand U23765 (N_23765,N_23644,N_23542);
or U23766 (N_23766,N_23691,N_23531);
or U23767 (N_23767,N_23392,N_23307);
nor U23768 (N_23768,N_23496,N_23711);
xnor U23769 (N_23769,N_23369,N_23619);
or U23770 (N_23770,N_23743,N_23246);
and U23771 (N_23771,N_23315,N_23651);
nand U23772 (N_23772,N_23235,N_23658);
or U23773 (N_23773,N_23710,N_23158);
xor U23774 (N_23774,N_23700,N_23546);
nand U23775 (N_23775,N_23516,N_23188);
xor U23776 (N_23776,N_23287,N_23503);
and U23777 (N_23777,N_23280,N_23154);
nand U23778 (N_23778,N_23702,N_23589);
or U23779 (N_23779,N_23138,N_23732);
and U23780 (N_23780,N_23519,N_23306);
nand U23781 (N_23781,N_23437,N_23703);
xor U23782 (N_23782,N_23329,N_23436);
xor U23783 (N_23783,N_23548,N_23736);
xor U23784 (N_23784,N_23247,N_23665);
nand U23785 (N_23785,N_23370,N_23467);
nor U23786 (N_23786,N_23493,N_23471);
nand U23787 (N_23787,N_23145,N_23662);
or U23788 (N_23788,N_23476,N_23621);
or U23789 (N_23789,N_23628,N_23230);
or U23790 (N_23790,N_23483,N_23741);
nor U23791 (N_23791,N_23196,N_23387);
nand U23792 (N_23792,N_23506,N_23341);
and U23793 (N_23793,N_23608,N_23418);
nor U23794 (N_23794,N_23352,N_23221);
and U23795 (N_23795,N_23408,N_23223);
nor U23796 (N_23796,N_23505,N_23458);
nand U23797 (N_23797,N_23217,N_23434);
xor U23798 (N_23798,N_23300,N_23739);
nor U23799 (N_23799,N_23149,N_23378);
or U23800 (N_23800,N_23731,N_23231);
xor U23801 (N_23801,N_23459,N_23322);
nor U23802 (N_23802,N_23504,N_23616);
nand U23803 (N_23803,N_23219,N_23648);
nand U23804 (N_23804,N_23432,N_23699);
xor U23805 (N_23805,N_23128,N_23414);
or U23806 (N_23806,N_23438,N_23253);
xnor U23807 (N_23807,N_23272,N_23278);
nor U23808 (N_23808,N_23177,N_23368);
nand U23809 (N_23809,N_23570,N_23299);
nand U23810 (N_23810,N_23705,N_23245);
and U23811 (N_23811,N_23540,N_23321);
nor U23812 (N_23812,N_23286,N_23681);
nor U23813 (N_23813,N_23355,N_23332);
nor U23814 (N_23814,N_23331,N_23529);
xnor U23815 (N_23815,N_23720,N_23412);
xor U23816 (N_23816,N_23281,N_23746);
nor U23817 (N_23817,N_23569,N_23684);
nor U23818 (N_23818,N_23533,N_23228);
and U23819 (N_23819,N_23450,N_23285);
xnor U23820 (N_23820,N_23379,N_23359);
or U23821 (N_23821,N_23690,N_23389);
xor U23822 (N_23822,N_23348,N_23682);
or U23823 (N_23823,N_23233,N_23468);
and U23824 (N_23824,N_23222,N_23553);
or U23825 (N_23825,N_23683,N_23187);
and U23826 (N_23826,N_23664,N_23740);
or U23827 (N_23827,N_23515,N_23183);
or U23828 (N_23828,N_23715,N_23475);
and U23829 (N_23829,N_23501,N_23537);
nand U23830 (N_23830,N_23381,N_23634);
and U23831 (N_23831,N_23641,N_23688);
or U23832 (N_23832,N_23376,N_23524);
xor U23833 (N_23833,N_23159,N_23422);
nand U23834 (N_23834,N_23627,N_23335);
xnor U23835 (N_23835,N_23197,N_23561);
nor U23836 (N_23836,N_23513,N_23581);
nand U23837 (N_23837,N_23696,N_23637);
or U23838 (N_23838,N_23595,N_23510);
and U23839 (N_23839,N_23319,N_23443);
and U23840 (N_23840,N_23125,N_23562);
xor U23841 (N_23841,N_23292,N_23265);
or U23842 (N_23842,N_23488,N_23350);
xor U23843 (N_23843,N_23206,N_23706);
nand U23844 (N_23844,N_23345,N_23630);
nand U23845 (N_23845,N_23185,N_23534);
or U23846 (N_23846,N_23168,N_23400);
and U23847 (N_23847,N_23251,N_23574);
or U23848 (N_23848,N_23176,N_23631);
or U23849 (N_23849,N_23304,N_23426);
nand U23850 (N_23850,N_23744,N_23357);
nand U23851 (N_23851,N_23127,N_23656);
nand U23852 (N_23852,N_23270,N_23729);
nor U23853 (N_23853,N_23749,N_23719);
or U23854 (N_23854,N_23579,N_23236);
xnor U23855 (N_23855,N_23727,N_23298);
nor U23856 (N_23856,N_23733,N_23267);
nor U23857 (N_23857,N_23486,N_23184);
or U23858 (N_23858,N_23709,N_23130);
xor U23859 (N_23859,N_23224,N_23216);
xor U23860 (N_23860,N_23137,N_23491);
or U23861 (N_23861,N_23153,N_23255);
or U23862 (N_23862,N_23191,N_23591);
and U23863 (N_23863,N_23615,N_23411);
nand U23864 (N_23864,N_23257,N_23593);
nand U23865 (N_23865,N_23209,N_23606);
nor U23866 (N_23866,N_23742,N_23337);
xor U23867 (N_23867,N_23661,N_23268);
nor U23868 (N_23868,N_23156,N_23576);
or U23869 (N_23869,N_23473,N_23351);
nor U23870 (N_23870,N_23240,N_23340);
nand U23871 (N_23871,N_23239,N_23404);
xnor U23872 (N_23872,N_23364,N_23334);
or U23873 (N_23873,N_23347,N_23472);
nand U23874 (N_23874,N_23655,N_23611);
and U23875 (N_23875,N_23126,N_23324);
nand U23876 (N_23876,N_23417,N_23617);
nor U23877 (N_23877,N_23445,N_23193);
nor U23878 (N_23878,N_23419,N_23618);
nor U23879 (N_23879,N_23164,N_23523);
and U23880 (N_23880,N_23312,N_23673);
or U23881 (N_23881,N_23250,N_23205);
xor U23882 (N_23882,N_23557,N_23363);
nor U23883 (N_23883,N_23202,N_23693);
and U23884 (N_23884,N_23313,N_23512);
or U23885 (N_23885,N_23406,N_23344);
or U23886 (N_23886,N_23600,N_23578);
or U23887 (N_23887,N_23479,N_23713);
or U23888 (N_23888,N_23712,N_23447);
and U23889 (N_23889,N_23132,N_23624);
and U23890 (N_23890,N_23291,N_23423);
nand U23891 (N_23891,N_23199,N_23717);
xnor U23892 (N_23892,N_23262,N_23674);
and U23893 (N_23893,N_23249,N_23290);
nand U23894 (N_23894,N_23566,N_23416);
xor U23895 (N_23895,N_23410,N_23528);
or U23896 (N_23896,N_23462,N_23413);
nand U23897 (N_23897,N_23716,N_23666);
nand U23898 (N_23898,N_23441,N_23480);
and U23899 (N_23899,N_23207,N_23358);
xor U23900 (N_23900,N_23572,N_23390);
and U23901 (N_23901,N_23195,N_23660);
or U23902 (N_23902,N_23603,N_23718);
nor U23903 (N_23903,N_23497,N_23421);
nor U23904 (N_23904,N_23254,N_23403);
or U23905 (N_23905,N_23427,N_23747);
nor U23906 (N_23906,N_23730,N_23178);
or U23907 (N_23907,N_23590,N_23643);
nor U23908 (N_23908,N_23568,N_23607);
or U23909 (N_23909,N_23330,N_23584);
or U23910 (N_23910,N_23234,N_23194);
or U23911 (N_23911,N_23377,N_23398);
xnor U23912 (N_23912,N_23386,N_23511);
xnor U23913 (N_23913,N_23293,N_23580);
and U23914 (N_23914,N_23653,N_23675);
and U23915 (N_23915,N_23614,N_23563);
nand U23916 (N_23916,N_23198,N_23499);
or U23917 (N_23917,N_23173,N_23170);
and U23918 (N_23918,N_23204,N_23564);
xor U23919 (N_23919,N_23144,N_23181);
nor U23920 (N_23920,N_23671,N_23526);
or U23921 (N_23921,N_23180,N_23484);
and U23922 (N_23922,N_23252,N_23565);
nand U23923 (N_23923,N_23200,N_23261);
nor U23924 (N_23924,N_23517,N_23449);
and U23925 (N_23925,N_23647,N_23162);
or U23926 (N_23926,N_23271,N_23288);
nand U23927 (N_23927,N_23596,N_23679);
xnor U23928 (N_23928,N_23316,N_23509);
or U23929 (N_23929,N_23657,N_23147);
or U23930 (N_23930,N_23361,N_23310);
xnor U23931 (N_23931,N_23672,N_23444);
and U23932 (N_23932,N_23670,N_23244);
or U23933 (N_23933,N_23396,N_23308);
or U23934 (N_23934,N_23210,N_23559);
nand U23935 (N_23935,N_23169,N_23609);
nor U23936 (N_23936,N_23133,N_23725);
xnor U23937 (N_23937,N_23136,N_23678);
and U23938 (N_23938,N_23555,N_23325);
or U23939 (N_23939,N_23586,N_23346);
nand U23940 (N_23940,N_23735,N_23260);
xor U23941 (N_23941,N_23652,N_23463);
nor U23942 (N_23942,N_23201,N_23726);
xor U23943 (N_23943,N_23558,N_23338);
and U23944 (N_23944,N_23650,N_23374);
xor U23945 (N_23945,N_23382,N_23520);
xnor U23946 (N_23946,N_23311,N_23259);
or U23947 (N_23947,N_23326,N_23539);
nand U23948 (N_23948,N_23461,N_23284);
xor U23949 (N_23949,N_23294,N_23192);
or U23950 (N_23950,N_23141,N_23535);
xor U23951 (N_23951,N_23482,N_23544);
nand U23952 (N_23952,N_23166,N_23277);
xor U23953 (N_23953,N_23646,N_23380);
or U23954 (N_23954,N_23645,N_23372);
nor U23955 (N_23955,N_23214,N_23582);
nor U23956 (N_23956,N_23454,N_23556);
nor U23957 (N_23957,N_23415,N_23135);
nand U23958 (N_23958,N_23687,N_23393);
xor U23959 (N_23959,N_23139,N_23226);
nor U23960 (N_23960,N_23466,N_23456);
and U23961 (N_23961,N_23375,N_23266);
xor U23962 (N_23962,N_23638,N_23161);
or U23963 (N_23963,N_23635,N_23242);
xnor U23964 (N_23964,N_23623,N_23685);
nand U23965 (N_23965,N_23433,N_23440);
nor U23966 (N_23966,N_23521,N_23323);
xnor U23967 (N_23967,N_23723,N_23680);
nand U23968 (N_23968,N_23490,N_23498);
nand U23969 (N_23969,N_23669,N_23186);
nor U23970 (N_23970,N_23543,N_23667);
xor U23971 (N_23971,N_23279,N_23227);
xor U23972 (N_23972,N_23612,N_23577);
xnor U23973 (N_23973,N_23554,N_23318);
nand U23974 (N_23974,N_23405,N_23424);
or U23975 (N_23975,N_23560,N_23677);
nand U23976 (N_23976,N_23722,N_23708);
nand U23977 (N_23977,N_23163,N_23273);
and U23978 (N_23978,N_23547,N_23659);
nor U23979 (N_23979,N_23431,N_23384);
nor U23980 (N_23980,N_23407,N_23317);
xnor U23981 (N_23981,N_23167,N_23238);
nor U23982 (N_23982,N_23388,N_23301);
nor U23983 (N_23983,N_23697,N_23707);
nor U23984 (N_23984,N_23551,N_23453);
or U23985 (N_23985,N_23243,N_23446);
nor U23986 (N_23986,N_23457,N_23269);
nor U23987 (N_23987,N_23140,N_23460);
or U23988 (N_23988,N_23625,N_23514);
nor U23989 (N_23989,N_23549,N_23508);
nor U23990 (N_23990,N_23212,N_23399);
xor U23991 (N_23991,N_23143,N_23371);
xor U23992 (N_23992,N_23724,N_23642);
nand U23993 (N_23993,N_23583,N_23314);
and U23994 (N_23994,N_23302,N_23492);
and U23995 (N_23995,N_23489,N_23604);
xnor U23996 (N_23996,N_23366,N_23686);
nand U23997 (N_23997,N_23694,N_23328);
nor U23998 (N_23998,N_23189,N_23704);
and U23999 (N_23999,N_23692,N_23391);
nor U24000 (N_24000,N_23203,N_23530);
nor U24001 (N_24001,N_23220,N_23430);
or U24002 (N_24002,N_23594,N_23575);
nor U24003 (N_24003,N_23320,N_23525);
and U24004 (N_24004,N_23155,N_23737);
or U24005 (N_24005,N_23538,N_23728);
nand U24006 (N_24006,N_23640,N_23146);
nand U24007 (N_24007,N_23283,N_23409);
and U24008 (N_24008,N_23385,N_23738);
or U24009 (N_24009,N_23474,N_23597);
or U24010 (N_24010,N_23598,N_23439);
xnor U24011 (N_24011,N_23541,N_23367);
or U24012 (N_24012,N_23485,N_23373);
xor U24013 (N_24013,N_23175,N_23536);
or U24014 (N_24014,N_23481,N_23601);
xnor U24015 (N_24015,N_23518,N_23428);
and U24016 (N_24016,N_23532,N_23343);
or U24017 (N_24017,N_23552,N_23342);
or U24018 (N_24018,N_23451,N_23225);
or U24019 (N_24019,N_23150,N_23383);
xnor U24020 (N_24020,N_23295,N_23237);
nand U24021 (N_24021,N_23349,N_23639);
xor U24022 (N_24022,N_23550,N_23592);
nor U24023 (N_24023,N_23585,N_23477);
and U24024 (N_24024,N_23613,N_23636);
xnor U24025 (N_24025,N_23172,N_23649);
nand U24026 (N_24026,N_23229,N_23487);
or U24027 (N_24027,N_23211,N_23296);
nand U24028 (N_24028,N_23626,N_23297);
xnor U24029 (N_24029,N_23327,N_23362);
or U24030 (N_24030,N_23303,N_23470);
nand U24031 (N_24031,N_23573,N_23633);
nor U24032 (N_24032,N_23339,N_23452);
nand U24033 (N_24033,N_23745,N_23248);
nor U24034 (N_24034,N_23241,N_23263);
nor U24035 (N_24035,N_23721,N_23289);
or U24036 (N_24036,N_23333,N_23353);
and U24037 (N_24037,N_23689,N_23478);
nand U24038 (N_24038,N_23190,N_23275);
and U24039 (N_24039,N_23620,N_23701);
and U24040 (N_24040,N_23397,N_23174);
nand U24041 (N_24041,N_23148,N_23131);
or U24042 (N_24042,N_23256,N_23629);
nor U24043 (N_24043,N_23464,N_23395);
nand U24044 (N_24044,N_23179,N_23469);
xor U24045 (N_24045,N_23401,N_23507);
xor U24046 (N_24046,N_23455,N_23495);
nor U24047 (N_24047,N_23420,N_23360);
or U24048 (N_24048,N_23215,N_23522);
or U24049 (N_24049,N_23208,N_23676);
and U24050 (N_24050,N_23354,N_23695);
xor U24051 (N_24051,N_23142,N_23394);
and U24052 (N_24052,N_23276,N_23588);
or U24053 (N_24053,N_23602,N_23448);
or U24054 (N_24054,N_23356,N_23336);
nor U24055 (N_24055,N_23305,N_23218);
xor U24056 (N_24056,N_23527,N_23663);
and U24057 (N_24057,N_23182,N_23365);
xnor U24058 (N_24058,N_23654,N_23500);
or U24059 (N_24059,N_23610,N_23599);
xor U24060 (N_24060,N_23748,N_23152);
nor U24061 (N_24061,N_23258,N_23698);
nand U24062 (N_24062,N_23134,N_23349);
or U24063 (N_24063,N_23723,N_23641);
or U24064 (N_24064,N_23283,N_23471);
and U24065 (N_24065,N_23239,N_23624);
nor U24066 (N_24066,N_23547,N_23218);
or U24067 (N_24067,N_23250,N_23619);
xnor U24068 (N_24068,N_23515,N_23453);
or U24069 (N_24069,N_23663,N_23722);
and U24070 (N_24070,N_23666,N_23474);
nor U24071 (N_24071,N_23199,N_23306);
xor U24072 (N_24072,N_23318,N_23188);
and U24073 (N_24073,N_23302,N_23590);
nor U24074 (N_24074,N_23192,N_23324);
nor U24075 (N_24075,N_23712,N_23513);
and U24076 (N_24076,N_23621,N_23668);
or U24077 (N_24077,N_23501,N_23327);
nand U24078 (N_24078,N_23138,N_23135);
or U24079 (N_24079,N_23473,N_23156);
and U24080 (N_24080,N_23566,N_23508);
xnor U24081 (N_24081,N_23643,N_23351);
and U24082 (N_24082,N_23259,N_23317);
nor U24083 (N_24083,N_23226,N_23732);
nand U24084 (N_24084,N_23353,N_23390);
and U24085 (N_24085,N_23403,N_23495);
or U24086 (N_24086,N_23152,N_23214);
and U24087 (N_24087,N_23255,N_23129);
and U24088 (N_24088,N_23201,N_23582);
xnor U24089 (N_24089,N_23196,N_23487);
xnor U24090 (N_24090,N_23168,N_23289);
and U24091 (N_24091,N_23674,N_23449);
nor U24092 (N_24092,N_23699,N_23599);
nand U24093 (N_24093,N_23283,N_23642);
nand U24094 (N_24094,N_23179,N_23346);
nand U24095 (N_24095,N_23320,N_23713);
or U24096 (N_24096,N_23365,N_23329);
xor U24097 (N_24097,N_23707,N_23166);
xor U24098 (N_24098,N_23182,N_23343);
nor U24099 (N_24099,N_23350,N_23313);
nor U24100 (N_24100,N_23557,N_23746);
nand U24101 (N_24101,N_23491,N_23632);
xor U24102 (N_24102,N_23324,N_23176);
or U24103 (N_24103,N_23394,N_23323);
nor U24104 (N_24104,N_23488,N_23359);
nor U24105 (N_24105,N_23620,N_23464);
nand U24106 (N_24106,N_23313,N_23227);
xnor U24107 (N_24107,N_23739,N_23627);
nand U24108 (N_24108,N_23376,N_23532);
or U24109 (N_24109,N_23606,N_23369);
or U24110 (N_24110,N_23135,N_23725);
nand U24111 (N_24111,N_23687,N_23282);
or U24112 (N_24112,N_23210,N_23552);
or U24113 (N_24113,N_23544,N_23706);
nor U24114 (N_24114,N_23497,N_23620);
nand U24115 (N_24115,N_23349,N_23744);
xor U24116 (N_24116,N_23675,N_23702);
and U24117 (N_24117,N_23662,N_23504);
and U24118 (N_24118,N_23335,N_23390);
nor U24119 (N_24119,N_23342,N_23259);
nand U24120 (N_24120,N_23197,N_23505);
xnor U24121 (N_24121,N_23241,N_23748);
nor U24122 (N_24122,N_23287,N_23721);
or U24123 (N_24123,N_23230,N_23252);
or U24124 (N_24124,N_23135,N_23463);
nand U24125 (N_24125,N_23384,N_23262);
xor U24126 (N_24126,N_23625,N_23246);
nand U24127 (N_24127,N_23246,N_23445);
or U24128 (N_24128,N_23245,N_23682);
xor U24129 (N_24129,N_23711,N_23317);
and U24130 (N_24130,N_23693,N_23306);
nand U24131 (N_24131,N_23574,N_23685);
xnor U24132 (N_24132,N_23323,N_23288);
and U24133 (N_24133,N_23220,N_23401);
nand U24134 (N_24134,N_23605,N_23258);
nand U24135 (N_24135,N_23566,N_23578);
xnor U24136 (N_24136,N_23672,N_23581);
nand U24137 (N_24137,N_23713,N_23492);
nand U24138 (N_24138,N_23469,N_23515);
nor U24139 (N_24139,N_23315,N_23482);
and U24140 (N_24140,N_23428,N_23171);
and U24141 (N_24141,N_23617,N_23745);
and U24142 (N_24142,N_23266,N_23189);
or U24143 (N_24143,N_23463,N_23516);
nand U24144 (N_24144,N_23716,N_23504);
nor U24145 (N_24145,N_23717,N_23235);
and U24146 (N_24146,N_23605,N_23604);
and U24147 (N_24147,N_23426,N_23710);
or U24148 (N_24148,N_23569,N_23343);
nor U24149 (N_24149,N_23421,N_23320);
and U24150 (N_24150,N_23429,N_23682);
xnor U24151 (N_24151,N_23222,N_23276);
and U24152 (N_24152,N_23723,N_23214);
and U24153 (N_24153,N_23158,N_23439);
nand U24154 (N_24154,N_23397,N_23706);
and U24155 (N_24155,N_23260,N_23507);
and U24156 (N_24156,N_23581,N_23238);
nor U24157 (N_24157,N_23684,N_23534);
xnor U24158 (N_24158,N_23686,N_23424);
nor U24159 (N_24159,N_23417,N_23221);
xor U24160 (N_24160,N_23647,N_23289);
nand U24161 (N_24161,N_23412,N_23196);
nand U24162 (N_24162,N_23147,N_23746);
and U24163 (N_24163,N_23537,N_23745);
nand U24164 (N_24164,N_23567,N_23659);
and U24165 (N_24165,N_23544,N_23611);
nand U24166 (N_24166,N_23354,N_23154);
xor U24167 (N_24167,N_23485,N_23129);
nor U24168 (N_24168,N_23291,N_23344);
xor U24169 (N_24169,N_23545,N_23457);
xnor U24170 (N_24170,N_23539,N_23127);
or U24171 (N_24171,N_23212,N_23695);
nor U24172 (N_24172,N_23171,N_23619);
and U24173 (N_24173,N_23710,N_23354);
or U24174 (N_24174,N_23675,N_23535);
xor U24175 (N_24175,N_23668,N_23452);
nand U24176 (N_24176,N_23127,N_23649);
or U24177 (N_24177,N_23260,N_23249);
or U24178 (N_24178,N_23253,N_23308);
or U24179 (N_24179,N_23326,N_23615);
or U24180 (N_24180,N_23260,N_23479);
and U24181 (N_24181,N_23215,N_23151);
or U24182 (N_24182,N_23594,N_23170);
or U24183 (N_24183,N_23196,N_23194);
or U24184 (N_24184,N_23638,N_23557);
nor U24185 (N_24185,N_23703,N_23520);
nand U24186 (N_24186,N_23577,N_23144);
and U24187 (N_24187,N_23222,N_23499);
xnor U24188 (N_24188,N_23699,N_23717);
or U24189 (N_24189,N_23263,N_23556);
nor U24190 (N_24190,N_23692,N_23665);
or U24191 (N_24191,N_23247,N_23653);
and U24192 (N_24192,N_23131,N_23433);
xor U24193 (N_24193,N_23687,N_23603);
or U24194 (N_24194,N_23229,N_23551);
xnor U24195 (N_24195,N_23147,N_23658);
or U24196 (N_24196,N_23476,N_23337);
and U24197 (N_24197,N_23404,N_23133);
and U24198 (N_24198,N_23297,N_23510);
xor U24199 (N_24199,N_23693,N_23423);
or U24200 (N_24200,N_23640,N_23681);
and U24201 (N_24201,N_23669,N_23481);
nor U24202 (N_24202,N_23458,N_23533);
or U24203 (N_24203,N_23724,N_23194);
nor U24204 (N_24204,N_23725,N_23470);
or U24205 (N_24205,N_23528,N_23443);
or U24206 (N_24206,N_23462,N_23540);
nor U24207 (N_24207,N_23482,N_23625);
nand U24208 (N_24208,N_23231,N_23342);
and U24209 (N_24209,N_23304,N_23555);
nand U24210 (N_24210,N_23313,N_23510);
nand U24211 (N_24211,N_23415,N_23394);
nor U24212 (N_24212,N_23131,N_23235);
nand U24213 (N_24213,N_23415,N_23641);
nand U24214 (N_24214,N_23493,N_23732);
nor U24215 (N_24215,N_23343,N_23682);
xor U24216 (N_24216,N_23144,N_23397);
nand U24217 (N_24217,N_23231,N_23539);
or U24218 (N_24218,N_23653,N_23360);
nor U24219 (N_24219,N_23300,N_23187);
nand U24220 (N_24220,N_23585,N_23132);
nand U24221 (N_24221,N_23384,N_23323);
nor U24222 (N_24222,N_23497,N_23447);
xor U24223 (N_24223,N_23672,N_23472);
or U24224 (N_24224,N_23146,N_23430);
or U24225 (N_24225,N_23365,N_23225);
xnor U24226 (N_24226,N_23590,N_23571);
xor U24227 (N_24227,N_23437,N_23538);
or U24228 (N_24228,N_23669,N_23356);
nand U24229 (N_24229,N_23654,N_23186);
nor U24230 (N_24230,N_23257,N_23225);
or U24231 (N_24231,N_23270,N_23742);
nand U24232 (N_24232,N_23136,N_23491);
or U24233 (N_24233,N_23452,N_23227);
nor U24234 (N_24234,N_23330,N_23253);
xnor U24235 (N_24235,N_23678,N_23308);
nand U24236 (N_24236,N_23471,N_23727);
xnor U24237 (N_24237,N_23713,N_23497);
nor U24238 (N_24238,N_23331,N_23283);
xor U24239 (N_24239,N_23251,N_23727);
nand U24240 (N_24240,N_23437,N_23614);
or U24241 (N_24241,N_23632,N_23293);
and U24242 (N_24242,N_23622,N_23733);
and U24243 (N_24243,N_23218,N_23443);
or U24244 (N_24244,N_23670,N_23426);
nor U24245 (N_24245,N_23211,N_23671);
and U24246 (N_24246,N_23271,N_23268);
or U24247 (N_24247,N_23224,N_23556);
xor U24248 (N_24248,N_23651,N_23263);
nand U24249 (N_24249,N_23509,N_23738);
nand U24250 (N_24250,N_23425,N_23259);
and U24251 (N_24251,N_23665,N_23612);
nor U24252 (N_24252,N_23308,N_23672);
xnor U24253 (N_24253,N_23481,N_23574);
or U24254 (N_24254,N_23418,N_23230);
or U24255 (N_24255,N_23375,N_23696);
and U24256 (N_24256,N_23518,N_23410);
and U24257 (N_24257,N_23608,N_23744);
nor U24258 (N_24258,N_23280,N_23477);
xor U24259 (N_24259,N_23305,N_23250);
and U24260 (N_24260,N_23131,N_23187);
or U24261 (N_24261,N_23735,N_23614);
nand U24262 (N_24262,N_23727,N_23728);
and U24263 (N_24263,N_23241,N_23414);
nand U24264 (N_24264,N_23319,N_23571);
nand U24265 (N_24265,N_23480,N_23519);
nor U24266 (N_24266,N_23602,N_23309);
nor U24267 (N_24267,N_23541,N_23308);
xnor U24268 (N_24268,N_23250,N_23480);
or U24269 (N_24269,N_23533,N_23321);
xor U24270 (N_24270,N_23200,N_23363);
xnor U24271 (N_24271,N_23361,N_23695);
and U24272 (N_24272,N_23675,N_23328);
or U24273 (N_24273,N_23538,N_23496);
and U24274 (N_24274,N_23170,N_23706);
nand U24275 (N_24275,N_23286,N_23595);
and U24276 (N_24276,N_23180,N_23604);
nor U24277 (N_24277,N_23214,N_23456);
xnor U24278 (N_24278,N_23745,N_23691);
xnor U24279 (N_24279,N_23715,N_23202);
xnor U24280 (N_24280,N_23401,N_23189);
xnor U24281 (N_24281,N_23505,N_23529);
or U24282 (N_24282,N_23662,N_23280);
and U24283 (N_24283,N_23577,N_23213);
nor U24284 (N_24284,N_23394,N_23372);
nor U24285 (N_24285,N_23448,N_23562);
and U24286 (N_24286,N_23378,N_23231);
and U24287 (N_24287,N_23181,N_23520);
or U24288 (N_24288,N_23323,N_23627);
nand U24289 (N_24289,N_23212,N_23361);
and U24290 (N_24290,N_23387,N_23142);
and U24291 (N_24291,N_23562,N_23529);
nand U24292 (N_24292,N_23427,N_23216);
and U24293 (N_24293,N_23622,N_23389);
nor U24294 (N_24294,N_23738,N_23236);
nand U24295 (N_24295,N_23484,N_23471);
and U24296 (N_24296,N_23511,N_23674);
nand U24297 (N_24297,N_23721,N_23473);
xnor U24298 (N_24298,N_23665,N_23465);
and U24299 (N_24299,N_23259,N_23320);
nor U24300 (N_24300,N_23705,N_23332);
or U24301 (N_24301,N_23305,N_23646);
and U24302 (N_24302,N_23554,N_23179);
and U24303 (N_24303,N_23250,N_23226);
xnor U24304 (N_24304,N_23572,N_23167);
nand U24305 (N_24305,N_23438,N_23223);
nor U24306 (N_24306,N_23379,N_23161);
or U24307 (N_24307,N_23225,N_23735);
or U24308 (N_24308,N_23703,N_23428);
nand U24309 (N_24309,N_23724,N_23564);
or U24310 (N_24310,N_23234,N_23621);
nand U24311 (N_24311,N_23394,N_23598);
nand U24312 (N_24312,N_23356,N_23540);
nor U24313 (N_24313,N_23224,N_23455);
xnor U24314 (N_24314,N_23534,N_23668);
nand U24315 (N_24315,N_23478,N_23663);
nor U24316 (N_24316,N_23201,N_23518);
nor U24317 (N_24317,N_23145,N_23147);
nand U24318 (N_24318,N_23299,N_23663);
xnor U24319 (N_24319,N_23552,N_23280);
nand U24320 (N_24320,N_23271,N_23683);
and U24321 (N_24321,N_23345,N_23371);
nor U24322 (N_24322,N_23656,N_23588);
nor U24323 (N_24323,N_23459,N_23488);
or U24324 (N_24324,N_23359,N_23240);
nor U24325 (N_24325,N_23480,N_23713);
nand U24326 (N_24326,N_23442,N_23445);
nor U24327 (N_24327,N_23157,N_23204);
or U24328 (N_24328,N_23351,N_23546);
nor U24329 (N_24329,N_23748,N_23422);
xnor U24330 (N_24330,N_23604,N_23600);
nand U24331 (N_24331,N_23214,N_23249);
and U24332 (N_24332,N_23395,N_23229);
or U24333 (N_24333,N_23502,N_23264);
and U24334 (N_24334,N_23538,N_23399);
and U24335 (N_24335,N_23678,N_23406);
nor U24336 (N_24336,N_23547,N_23569);
nand U24337 (N_24337,N_23710,N_23684);
and U24338 (N_24338,N_23352,N_23548);
nand U24339 (N_24339,N_23371,N_23265);
xor U24340 (N_24340,N_23609,N_23674);
and U24341 (N_24341,N_23356,N_23266);
nand U24342 (N_24342,N_23282,N_23411);
and U24343 (N_24343,N_23149,N_23608);
nor U24344 (N_24344,N_23739,N_23424);
xnor U24345 (N_24345,N_23381,N_23153);
and U24346 (N_24346,N_23467,N_23392);
or U24347 (N_24347,N_23596,N_23627);
and U24348 (N_24348,N_23510,N_23532);
xnor U24349 (N_24349,N_23704,N_23488);
nor U24350 (N_24350,N_23323,N_23493);
nor U24351 (N_24351,N_23645,N_23484);
and U24352 (N_24352,N_23524,N_23247);
nand U24353 (N_24353,N_23188,N_23324);
xnor U24354 (N_24354,N_23370,N_23256);
and U24355 (N_24355,N_23174,N_23542);
and U24356 (N_24356,N_23454,N_23512);
nand U24357 (N_24357,N_23600,N_23450);
or U24358 (N_24358,N_23418,N_23610);
xor U24359 (N_24359,N_23515,N_23279);
nor U24360 (N_24360,N_23195,N_23631);
and U24361 (N_24361,N_23196,N_23299);
and U24362 (N_24362,N_23148,N_23591);
nor U24363 (N_24363,N_23691,N_23156);
or U24364 (N_24364,N_23742,N_23721);
nand U24365 (N_24365,N_23669,N_23424);
or U24366 (N_24366,N_23383,N_23547);
and U24367 (N_24367,N_23331,N_23333);
and U24368 (N_24368,N_23166,N_23268);
nor U24369 (N_24369,N_23690,N_23273);
nand U24370 (N_24370,N_23256,N_23334);
and U24371 (N_24371,N_23307,N_23660);
nor U24372 (N_24372,N_23626,N_23522);
and U24373 (N_24373,N_23484,N_23155);
nor U24374 (N_24374,N_23216,N_23714);
xor U24375 (N_24375,N_24133,N_23949);
and U24376 (N_24376,N_24186,N_23892);
xnor U24377 (N_24377,N_24337,N_24180);
xnor U24378 (N_24378,N_24045,N_23982);
nand U24379 (N_24379,N_24087,N_24101);
nor U24380 (N_24380,N_24373,N_23973);
nand U24381 (N_24381,N_24030,N_24077);
nor U24382 (N_24382,N_23937,N_23946);
nor U24383 (N_24383,N_24216,N_24312);
or U24384 (N_24384,N_23789,N_23986);
nand U24385 (N_24385,N_23880,N_24081);
and U24386 (N_24386,N_24232,N_24158);
or U24387 (N_24387,N_23885,N_24119);
xor U24388 (N_24388,N_23984,N_24126);
nand U24389 (N_24389,N_24224,N_23894);
and U24390 (N_24390,N_23807,N_24089);
nor U24391 (N_24391,N_24141,N_24091);
xnor U24392 (N_24392,N_24292,N_23914);
or U24393 (N_24393,N_24291,N_23839);
xnor U24394 (N_24394,N_24155,N_24169);
and U24395 (N_24395,N_23996,N_23833);
xor U24396 (N_24396,N_23907,N_24098);
nand U24397 (N_24397,N_24238,N_23778);
or U24398 (N_24398,N_23875,N_24111);
and U24399 (N_24399,N_23795,N_23969);
or U24400 (N_24400,N_24107,N_23995);
nand U24401 (N_24401,N_23815,N_23947);
xor U24402 (N_24402,N_24104,N_24191);
nand U24403 (N_24403,N_23757,N_24202);
nand U24404 (N_24404,N_23906,N_23966);
or U24405 (N_24405,N_23932,N_23896);
xor U24406 (N_24406,N_23941,N_24157);
nand U24407 (N_24407,N_24192,N_24143);
or U24408 (N_24408,N_24340,N_23766);
xnor U24409 (N_24409,N_23988,N_23888);
and U24410 (N_24410,N_24173,N_24042);
or U24411 (N_24411,N_23989,N_23769);
nor U24412 (N_24412,N_24288,N_24055);
nor U24413 (N_24413,N_24175,N_24294);
nand U24414 (N_24414,N_24132,N_24116);
nand U24415 (N_24415,N_24115,N_24165);
nand U24416 (N_24416,N_24039,N_23876);
xor U24417 (N_24417,N_23871,N_24122);
nand U24418 (N_24418,N_23879,N_23884);
nor U24419 (N_24419,N_23849,N_23828);
or U24420 (N_24420,N_24050,N_24334);
nor U24421 (N_24421,N_24052,N_24043);
and U24422 (N_24422,N_24240,N_24059);
nand U24423 (N_24423,N_24250,N_23926);
nand U24424 (N_24424,N_23813,N_23878);
or U24425 (N_24425,N_24276,N_23983);
and U24426 (N_24426,N_24219,N_23905);
or U24427 (N_24427,N_23809,N_23868);
or U24428 (N_24428,N_24067,N_24363);
and U24429 (N_24429,N_24233,N_24073);
and U24430 (N_24430,N_23832,N_24053);
nor U24431 (N_24431,N_24128,N_24011);
and U24432 (N_24432,N_23862,N_24283);
and U24433 (N_24433,N_24237,N_23797);
nand U24434 (N_24434,N_23760,N_23758);
nor U24435 (N_24435,N_24106,N_24351);
nand U24436 (N_24436,N_24035,N_24287);
or U24437 (N_24437,N_24172,N_24293);
nor U24438 (N_24438,N_24002,N_23812);
nor U24439 (N_24439,N_24003,N_24093);
xor U24440 (N_24440,N_24307,N_23843);
xnor U24441 (N_24441,N_23854,N_23818);
nand U24442 (N_24442,N_24020,N_23931);
or U24443 (N_24443,N_24282,N_24153);
and U24444 (N_24444,N_24356,N_23800);
or U24445 (N_24445,N_24161,N_24201);
or U24446 (N_24446,N_23831,N_24222);
or U24447 (N_24447,N_24114,N_24362);
nand U24448 (N_24448,N_24195,N_24321);
and U24449 (N_24449,N_24206,N_24062);
nor U24450 (N_24450,N_24350,N_24308);
and U24451 (N_24451,N_23985,N_23951);
nand U24452 (N_24452,N_23837,N_23955);
nand U24453 (N_24453,N_23847,N_24085);
or U24454 (N_24454,N_23957,N_24121);
xnor U24455 (N_24455,N_24084,N_23846);
nor U24456 (N_24456,N_23997,N_24313);
and U24457 (N_24457,N_23979,N_24159);
xor U24458 (N_24458,N_23981,N_24215);
nand U24459 (N_24459,N_24160,N_24264);
nor U24460 (N_24460,N_24247,N_23762);
and U24461 (N_24461,N_24295,N_24148);
xnor U24462 (N_24462,N_24317,N_24174);
or U24463 (N_24463,N_23883,N_24086);
or U24464 (N_24464,N_23841,N_24253);
xor U24465 (N_24465,N_24124,N_24271);
or U24466 (N_24466,N_23943,N_23808);
and U24467 (N_24467,N_24017,N_24070);
or U24468 (N_24468,N_23919,N_23882);
nor U24469 (N_24469,N_24349,N_24127);
or U24470 (N_24470,N_23819,N_24024);
xor U24471 (N_24471,N_24280,N_24210);
and U24472 (N_24472,N_24069,N_24185);
or U24473 (N_24473,N_24140,N_24171);
or U24474 (N_24474,N_24008,N_23793);
xor U24475 (N_24475,N_23781,N_24197);
xor U24476 (N_24476,N_23835,N_24080);
nand U24477 (N_24477,N_24142,N_24242);
or U24478 (N_24478,N_24023,N_24044);
xnor U24479 (N_24479,N_23825,N_23791);
xnor U24480 (N_24480,N_23796,N_24095);
nand U24481 (N_24481,N_24096,N_24156);
nand U24482 (N_24482,N_23820,N_24259);
nand U24483 (N_24483,N_24103,N_24322);
xor U24484 (N_24484,N_24167,N_24040);
xnor U24485 (N_24485,N_23804,N_24117);
nor U24486 (N_24486,N_24061,N_23844);
nor U24487 (N_24487,N_24331,N_24014);
nand U24488 (N_24488,N_23848,N_23802);
nand U24489 (N_24489,N_24251,N_23889);
nand U24490 (N_24490,N_24269,N_23806);
xor U24491 (N_24491,N_23962,N_23805);
nand U24492 (N_24492,N_24088,N_23952);
or U24493 (N_24493,N_24353,N_23920);
nor U24494 (N_24494,N_23759,N_23908);
or U24495 (N_24495,N_23790,N_24068);
xor U24496 (N_24496,N_24268,N_24208);
and U24497 (N_24497,N_23913,N_24105);
or U24498 (N_24498,N_24299,N_24248);
xnor U24499 (N_24499,N_24138,N_24012);
nor U24500 (N_24500,N_24004,N_23799);
xnor U24501 (N_24501,N_23754,N_24342);
xnor U24502 (N_24502,N_24236,N_24041);
nor U24503 (N_24503,N_24267,N_24252);
xnor U24504 (N_24504,N_23823,N_24209);
or U24505 (N_24505,N_24212,N_24179);
or U24506 (N_24506,N_24365,N_24223);
nor U24507 (N_24507,N_24245,N_23788);
and U24508 (N_24508,N_24314,N_24108);
and U24509 (N_24509,N_24125,N_24190);
nor U24510 (N_24510,N_23827,N_24225);
or U24511 (N_24511,N_23936,N_24151);
xnor U24512 (N_24512,N_23770,N_23923);
nand U24513 (N_24513,N_23874,N_23777);
or U24514 (N_24514,N_23953,N_23910);
nand U24515 (N_24515,N_23856,N_24304);
nor U24516 (N_24516,N_24135,N_23773);
or U24517 (N_24517,N_24200,N_23980);
and U24518 (N_24518,N_24181,N_24131);
nor U24519 (N_24519,N_24320,N_24094);
and U24520 (N_24520,N_24338,N_24277);
and U24521 (N_24521,N_24249,N_23909);
nor U24522 (N_24522,N_23929,N_24255);
xnor U24523 (N_24523,N_23930,N_23824);
nand U24524 (N_24524,N_24332,N_24170);
xor U24525 (N_24525,N_23954,N_23842);
or U24526 (N_24526,N_24246,N_23959);
and U24527 (N_24527,N_24099,N_24120);
xor U24528 (N_24528,N_23971,N_24305);
nor U24529 (N_24529,N_24203,N_24330);
and U24530 (N_24530,N_23893,N_24336);
or U24531 (N_24531,N_23897,N_24051);
or U24532 (N_24532,N_24164,N_24278);
and U24533 (N_24533,N_24037,N_24207);
xnor U24534 (N_24534,N_23921,N_24266);
and U24535 (N_24535,N_24046,N_24359);
nand U24536 (N_24536,N_24297,N_23976);
nand U24537 (N_24537,N_23934,N_24129);
and U24538 (N_24538,N_23821,N_24234);
xnor U24539 (N_24539,N_24047,N_24025);
nand U24540 (N_24540,N_23785,N_24256);
xnor U24541 (N_24541,N_23903,N_24281);
or U24542 (N_24542,N_24066,N_24031);
or U24543 (N_24543,N_24354,N_24265);
nor U24544 (N_24544,N_23869,N_24072);
xor U24545 (N_24545,N_24021,N_24372);
xor U24546 (N_24546,N_23834,N_23990);
nor U24547 (N_24547,N_23775,N_24341);
and U24548 (N_24548,N_23840,N_23960);
or U24549 (N_24549,N_24056,N_24065);
nand U24550 (N_24550,N_24235,N_23977);
and U24551 (N_24551,N_24007,N_24227);
nand U24552 (N_24552,N_24316,N_24286);
nand U24553 (N_24553,N_24213,N_23851);
xnor U24554 (N_24554,N_24346,N_23863);
and U24555 (N_24555,N_23916,N_23928);
and U24556 (N_24556,N_23956,N_24188);
nand U24557 (N_24557,N_24029,N_23752);
or U24558 (N_24558,N_24149,N_24000);
xnor U24559 (N_24559,N_24364,N_23776);
and U24560 (N_24560,N_24327,N_24090);
nand U24561 (N_24561,N_24198,N_24339);
and U24562 (N_24562,N_23810,N_24315);
or U24563 (N_24563,N_24345,N_24118);
or U24564 (N_24564,N_23751,N_23940);
nand U24565 (N_24565,N_24071,N_24303);
or U24566 (N_24566,N_23991,N_24054);
and U24567 (N_24567,N_24183,N_24205);
and U24568 (N_24568,N_23784,N_23826);
and U24569 (N_24569,N_24296,N_23899);
nand U24570 (N_24570,N_23873,N_24184);
and U24571 (N_24571,N_24163,N_24344);
nor U24572 (N_24572,N_23803,N_23881);
xnor U24573 (N_24573,N_24019,N_23912);
xnor U24574 (N_24574,N_23968,N_24368);
xnor U24575 (N_24575,N_24326,N_23902);
nand U24576 (N_24576,N_24009,N_24371);
nor U24577 (N_24577,N_24302,N_23755);
nor U24578 (N_24578,N_23898,N_24074);
xor U24579 (N_24579,N_24319,N_23786);
nand U24580 (N_24580,N_24136,N_23938);
nor U24581 (N_24581,N_23877,N_24328);
nor U24582 (N_24582,N_24150,N_24300);
xnor U24583 (N_24583,N_24262,N_24145);
nand U24584 (N_24584,N_24366,N_24178);
nor U24585 (N_24585,N_24123,N_23867);
xor U24586 (N_24586,N_24358,N_24199);
xor U24587 (N_24587,N_24102,N_24005);
or U24588 (N_24588,N_24284,N_23922);
nand U24589 (N_24589,N_23964,N_24063);
or U24590 (N_24590,N_23763,N_24311);
or U24591 (N_24591,N_23782,N_23970);
or U24592 (N_24592,N_24194,N_24082);
nor U24593 (N_24593,N_24367,N_23974);
and U24594 (N_24594,N_23787,N_23994);
nand U24595 (N_24595,N_24285,N_24301);
and U24596 (N_24596,N_23895,N_23935);
or U24597 (N_24597,N_23865,N_23948);
and U24598 (N_24598,N_23857,N_23838);
xor U24599 (N_24599,N_23860,N_23891);
nand U24600 (N_24600,N_24026,N_23829);
and U24601 (N_24601,N_23939,N_24083);
nor U24602 (N_24602,N_24130,N_24360);
xnor U24603 (N_24603,N_24275,N_24347);
nand U24604 (N_24604,N_23925,N_24289);
and U24605 (N_24605,N_24369,N_24261);
nand U24606 (N_24606,N_23767,N_23992);
nand U24607 (N_24607,N_24076,N_23887);
and U24608 (N_24608,N_23942,N_23999);
or U24609 (N_24609,N_23780,N_24187);
nor U24610 (N_24610,N_24147,N_23772);
nor U24611 (N_24611,N_23963,N_23918);
or U24612 (N_24612,N_24176,N_23978);
or U24613 (N_24613,N_24211,N_24038);
and U24614 (N_24614,N_23817,N_24109);
xnor U24615 (N_24615,N_24168,N_23779);
or U24616 (N_24616,N_24323,N_23822);
or U24617 (N_24617,N_24060,N_24258);
nor U24618 (N_24618,N_24204,N_23904);
nor U24619 (N_24619,N_24058,N_24309);
xnor U24620 (N_24620,N_23859,N_24162);
or U24621 (N_24621,N_23792,N_23987);
xor U24622 (N_24622,N_23972,N_24243);
or U24623 (N_24623,N_23886,N_24231);
and U24624 (N_24624,N_23811,N_23794);
nor U24625 (N_24625,N_24214,N_24310);
nand U24626 (N_24626,N_24048,N_23764);
or U24627 (N_24627,N_24022,N_23771);
nand U24628 (N_24628,N_24335,N_24097);
nor U24629 (N_24629,N_24306,N_23830);
and U24630 (N_24630,N_24177,N_23998);
xor U24631 (N_24631,N_24329,N_23933);
nand U24632 (N_24632,N_24348,N_24027);
xor U24633 (N_24633,N_24374,N_23944);
xnor U24634 (N_24634,N_23750,N_24032);
or U24635 (N_24635,N_23901,N_24146);
and U24636 (N_24636,N_24220,N_23924);
or U24637 (N_24637,N_24196,N_24013);
nand U24638 (N_24638,N_24370,N_24272);
or U24639 (N_24639,N_23774,N_24006);
and U24640 (N_24640,N_23993,N_23756);
xor U24641 (N_24641,N_24033,N_24218);
and U24642 (N_24642,N_23836,N_24137);
or U24643 (N_24643,N_23927,N_23801);
nor U24644 (N_24644,N_24092,N_23768);
xor U24645 (N_24645,N_24112,N_24263);
or U24646 (N_24646,N_24134,N_24270);
nand U24647 (N_24647,N_24290,N_23945);
and U24648 (N_24648,N_23798,N_24057);
nand U24649 (N_24649,N_24049,N_24217);
nor U24650 (N_24650,N_23961,N_24154);
nor U24651 (N_24651,N_24257,N_24193);
or U24652 (N_24652,N_24343,N_24113);
nor U24653 (N_24653,N_23761,N_24144);
nand U24654 (N_24654,N_24036,N_24016);
and U24655 (N_24655,N_24274,N_23965);
xor U24656 (N_24656,N_24100,N_24079);
nor U24657 (N_24657,N_24324,N_24189);
and U24658 (N_24658,N_23958,N_24152);
xnor U24659 (N_24659,N_24333,N_24166);
or U24660 (N_24660,N_24229,N_23853);
or U24661 (N_24661,N_24182,N_23845);
nor U24662 (N_24662,N_24075,N_24001);
or U24663 (N_24663,N_23858,N_24078);
and U24664 (N_24664,N_23967,N_24273);
and U24665 (N_24665,N_24352,N_23890);
nand U24666 (N_24666,N_24064,N_24241);
xor U24667 (N_24667,N_24355,N_24034);
and U24668 (N_24668,N_24110,N_24298);
and U24669 (N_24669,N_23872,N_23816);
nand U24670 (N_24670,N_23870,N_24279);
and U24671 (N_24671,N_23866,N_23861);
nor U24672 (N_24672,N_23852,N_24325);
nand U24673 (N_24673,N_23855,N_24228);
or U24674 (N_24674,N_23917,N_24318);
or U24675 (N_24675,N_24361,N_24254);
nor U24676 (N_24676,N_23814,N_24230);
xor U24677 (N_24677,N_23900,N_24010);
nor U24678 (N_24678,N_24028,N_24260);
or U24679 (N_24679,N_23850,N_24357);
nor U24680 (N_24680,N_24015,N_23950);
nor U24681 (N_24681,N_24239,N_23753);
or U24682 (N_24682,N_23783,N_23765);
nand U24683 (N_24683,N_23915,N_24018);
or U24684 (N_24684,N_24139,N_24226);
nor U24685 (N_24685,N_24244,N_23911);
and U24686 (N_24686,N_23864,N_23975);
nand U24687 (N_24687,N_24221,N_23912);
nor U24688 (N_24688,N_23859,N_24253);
and U24689 (N_24689,N_24274,N_24156);
and U24690 (N_24690,N_24134,N_24233);
nor U24691 (N_24691,N_23973,N_23750);
nand U24692 (N_24692,N_23850,N_24044);
nor U24693 (N_24693,N_23990,N_24119);
or U24694 (N_24694,N_24046,N_23942);
xnor U24695 (N_24695,N_24266,N_24175);
nand U24696 (N_24696,N_23949,N_23904);
or U24697 (N_24697,N_24074,N_23891);
nor U24698 (N_24698,N_24066,N_23873);
or U24699 (N_24699,N_24258,N_24127);
nor U24700 (N_24700,N_24328,N_24267);
and U24701 (N_24701,N_24055,N_24219);
and U24702 (N_24702,N_24215,N_23774);
nor U24703 (N_24703,N_23988,N_23968);
and U24704 (N_24704,N_24179,N_23985);
nor U24705 (N_24705,N_24044,N_24230);
nand U24706 (N_24706,N_24174,N_23760);
xnor U24707 (N_24707,N_23940,N_24141);
nand U24708 (N_24708,N_24182,N_24135);
nor U24709 (N_24709,N_24275,N_23981);
and U24710 (N_24710,N_24062,N_24359);
nand U24711 (N_24711,N_23984,N_23774);
nor U24712 (N_24712,N_24291,N_24228);
or U24713 (N_24713,N_24034,N_24182);
xnor U24714 (N_24714,N_24066,N_23893);
nand U24715 (N_24715,N_23861,N_24343);
nor U24716 (N_24716,N_23803,N_24039);
or U24717 (N_24717,N_23867,N_24067);
nand U24718 (N_24718,N_23934,N_24130);
nor U24719 (N_24719,N_23912,N_24257);
and U24720 (N_24720,N_23834,N_24121);
nand U24721 (N_24721,N_23776,N_24095);
nor U24722 (N_24722,N_23832,N_24010);
or U24723 (N_24723,N_23821,N_24160);
or U24724 (N_24724,N_24318,N_24065);
nand U24725 (N_24725,N_23910,N_24024);
nand U24726 (N_24726,N_24223,N_23844);
nand U24727 (N_24727,N_24221,N_23922);
or U24728 (N_24728,N_24178,N_24145);
nand U24729 (N_24729,N_24185,N_24301);
and U24730 (N_24730,N_24310,N_23797);
xor U24731 (N_24731,N_24337,N_23955);
or U24732 (N_24732,N_23867,N_24037);
and U24733 (N_24733,N_24123,N_24286);
xnor U24734 (N_24734,N_24039,N_24142);
nor U24735 (N_24735,N_24332,N_24242);
or U24736 (N_24736,N_24008,N_24100);
and U24737 (N_24737,N_24268,N_24312);
nor U24738 (N_24738,N_24275,N_24356);
or U24739 (N_24739,N_23760,N_24047);
nor U24740 (N_24740,N_24325,N_24368);
and U24741 (N_24741,N_23968,N_23918);
nand U24742 (N_24742,N_23971,N_24309);
xnor U24743 (N_24743,N_23869,N_23807);
or U24744 (N_24744,N_24169,N_23776);
nor U24745 (N_24745,N_24338,N_23931);
nand U24746 (N_24746,N_23773,N_23838);
nor U24747 (N_24747,N_24040,N_24255);
xor U24748 (N_24748,N_24359,N_24283);
nor U24749 (N_24749,N_24318,N_23765);
nor U24750 (N_24750,N_23830,N_24062);
and U24751 (N_24751,N_23899,N_24101);
nand U24752 (N_24752,N_24049,N_24260);
nand U24753 (N_24753,N_24225,N_24281);
nor U24754 (N_24754,N_24268,N_24370);
nand U24755 (N_24755,N_24176,N_24342);
and U24756 (N_24756,N_23773,N_24309);
or U24757 (N_24757,N_24112,N_23893);
nand U24758 (N_24758,N_23766,N_24064);
xor U24759 (N_24759,N_24035,N_24065);
or U24760 (N_24760,N_24101,N_24203);
nand U24761 (N_24761,N_24353,N_24059);
and U24762 (N_24762,N_24128,N_24026);
and U24763 (N_24763,N_23796,N_24148);
nor U24764 (N_24764,N_23864,N_24253);
nand U24765 (N_24765,N_24278,N_24087);
nand U24766 (N_24766,N_23936,N_23814);
and U24767 (N_24767,N_24037,N_24088);
and U24768 (N_24768,N_24004,N_23948);
or U24769 (N_24769,N_23790,N_23993);
nor U24770 (N_24770,N_24071,N_24194);
and U24771 (N_24771,N_23817,N_23762);
and U24772 (N_24772,N_24165,N_24246);
xnor U24773 (N_24773,N_24244,N_23877);
or U24774 (N_24774,N_24150,N_24309);
xor U24775 (N_24775,N_24107,N_24022);
xor U24776 (N_24776,N_24116,N_23992);
xnor U24777 (N_24777,N_23876,N_24142);
nor U24778 (N_24778,N_23992,N_24168);
nor U24779 (N_24779,N_23958,N_24208);
nand U24780 (N_24780,N_24271,N_24152);
nand U24781 (N_24781,N_24167,N_23956);
xor U24782 (N_24782,N_24294,N_24185);
xor U24783 (N_24783,N_23973,N_24087);
nand U24784 (N_24784,N_24012,N_24140);
and U24785 (N_24785,N_23760,N_24049);
xor U24786 (N_24786,N_24153,N_24360);
and U24787 (N_24787,N_24161,N_23850);
and U24788 (N_24788,N_24114,N_24318);
nor U24789 (N_24789,N_23769,N_23974);
or U24790 (N_24790,N_24320,N_24012);
nand U24791 (N_24791,N_24244,N_24117);
xor U24792 (N_24792,N_24188,N_23766);
and U24793 (N_24793,N_24337,N_23877);
nand U24794 (N_24794,N_24250,N_23789);
and U24795 (N_24795,N_23915,N_24373);
and U24796 (N_24796,N_24143,N_24275);
nor U24797 (N_24797,N_24319,N_24051);
or U24798 (N_24798,N_24293,N_24307);
nor U24799 (N_24799,N_23981,N_24193);
and U24800 (N_24800,N_24342,N_24238);
nor U24801 (N_24801,N_24030,N_24356);
xor U24802 (N_24802,N_24210,N_23918);
and U24803 (N_24803,N_23805,N_23786);
nand U24804 (N_24804,N_24125,N_23927);
nand U24805 (N_24805,N_23814,N_23944);
nor U24806 (N_24806,N_23868,N_24333);
nor U24807 (N_24807,N_24000,N_24247);
xor U24808 (N_24808,N_24109,N_24212);
or U24809 (N_24809,N_23860,N_24157);
or U24810 (N_24810,N_23817,N_23979);
nand U24811 (N_24811,N_23934,N_23840);
and U24812 (N_24812,N_24270,N_24014);
or U24813 (N_24813,N_24091,N_24113);
xor U24814 (N_24814,N_24050,N_23783);
and U24815 (N_24815,N_23769,N_24236);
or U24816 (N_24816,N_24109,N_23897);
and U24817 (N_24817,N_23862,N_23858);
xor U24818 (N_24818,N_24131,N_23898);
or U24819 (N_24819,N_24005,N_24026);
xnor U24820 (N_24820,N_24154,N_24195);
nand U24821 (N_24821,N_24051,N_24121);
nand U24822 (N_24822,N_24264,N_24363);
nand U24823 (N_24823,N_24102,N_24019);
nand U24824 (N_24824,N_23772,N_24106);
or U24825 (N_24825,N_23855,N_23984);
xor U24826 (N_24826,N_24183,N_23978);
or U24827 (N_24827,N_23964,N_23922);
xor U24828 (N_24828,N_23997,N_24243);
nor U24829 (N_24829,N_23779,N_24339);
xor U24830 (N_24830,N_23902,N_23972);
or U24831 (N_24831,N_24010,N_24144);
nand U24832 (N_24832,N_23967,N_23919);
nor U24833 (N_24833,N_23910,N_23955);
nor U24834 (N_24834,N_24361,N_24286);
nand U24835 (N_24835,N_24101,N_23959);
nand U24836 (N_24836,N_23820,N_24039);
xor U24837 (N_24837,N_24033,N_23805);
nand U24838 (N_24838,N_24300,N_24044);
and U24839 (N_24839,N_24348,N_24031);
and U24840 (N_24840,N_24136,N_24014);
and U24841 (N_24841,N_24138,N_23871);
nor U24842 (N_24842,N_23915,N_23962);
or U24843 (N_24843,N_23982,N_24137);
and U24844 (N_24844,N_24288,N_24285);
or U24845 (N_24845,N_23998,N_23803);
nor U24846 (N_24846,N_23904,N_24315);
or U24847 (N_24847,N_23767,N_24155);
nor U24848 (N_24848,N_24226,N_23820);
nand U24849 (N_24849,N_23786,N_24255);
or U24850 (N_24850,N_24175,N_24049);
nand U24851 (N_24851,N_24093,N_24154);
or U24852 (N_24852,N_24227,N_23990);
xnor U24853 (N_24853,N_23852,N_24279);
nand U24854 (N_24854,N_24347,N_24244);
xor U24855 (N_24855,N_24142,N_24305);
nor U24856 (N_24856,N_24139,N_24175);
nand U24857 (N_24857,N_23765,N_23767);
and U24858 (N_24858,N_24209,N_23976);
nor U24859 (N_24859,N_23800,N_23910);
or U24860 (N_24860,N_24043,N_24295);
nand U24861 (N_24861,N_24085,N_24030);
nand U24862 (N_24862,N_24017,N_23837);
and U24863 (N_24863,N_24089,N_24110);
or U24864 (N_24864,N_24374,N_24355);
nand U24865 (N_24865,N_24229,N_23796);
nand U24866 (N_24866,N_24170,N_24222);
or U24867 (N_24867,N_24339,N_24353);
and U24868 (N_24868,N_23844,N_23865);
nor U24869 (N_24869,N_23861,N_24021);
nor U24870 (N_24870,N_23862,N_23962);
xor U24871 (N_24871,N_23960,N_24312);
nand U24872 (N_24872,N_24032,N_24350);
or U24873 (N_24873,N_23832,N_24082);
nand U24874 (N_24874,N_23760,N_24374);
xor U24875 (N_24875,N_24325,N_24164);
xnor U24876 (N_24876,N_24096,N_23878);
and U24877 (N_24877,N_23964,N_24371);
nor U24878 (N_24878,N_24228,N_23871);
or U24879 (N_24879,N_24222,N_23955);
nand U24880 (N_24880,N_23936,N_24062);
and U24881 (N_24881,N_24324,N_24195);
and U24882 (N_24882,N_23809,N_24281);
and U24883 (N_24883,N_24292,N_23804);
or U24884 (N_24884,N_23783,N_24323);
xnor U24885 (N_24885,N_24053,N_23918);
xor U24886 (N_24886,N_24007,N_24229);
xor U24887 (N_24887,N_24109,N_23760);
and U24888 (N_24888,N_24283,N_23846);
nor U24889 (N_24889,N_24113,N_23843);
nand U24890 (N_24890,N_24174,N_24204);
and U24891 (N_24891,N_23802,N_24374);
nand U24892 (N_24892,N_24060,N_24261);
nor U24893 (N_24893,N_24102,N_23836);
and U24894 (N_24894,N_24104,N_24251);
or U24895 (N_24895,N_23954,N_23853);
and U24896 (N_24896,N_23889,N_24365);
xor U24897 (N_24897,N_24002,N_23935);
or U24898 (N_24898,N_24115,N_24349);
xnor U24899 (N_24899,N_24106,N_24092);
and U24900 (N_24900,N_24104,N_24241);
xnor U24901 (N_24901,N_23841,N_23981);
nor U24902 (N_24902,N_23920,N_23959);
or U24903 (N_24903,N_23771,N_23868);
xor U24904 (N_24904,N_24356,N_24177);
and U24905 (N_24905,N_23955,N_24365);
nand U24906 (N_24906,N_24139,N_24191);
or U24907 (N_24907,N_24269,N_23873);
or U24908 (N_24908,N_23910,N_24049);
xnor U24909 (N_24909,N_23965,N_23972);
nand U24910 (N_24910,N_23947,N_23850);
xor U24911 (N_24911,N_24111,N_23848);
and U24912 (N_24912,N_24003,N_24329);
nand U24913 (N_24913,N_23841,N_23994);
nand U24914 (N_24914,N_23825,N_23956);
or U24915 (N_24915,N_24120,N_24008);
or U24916 (N_24916,N_23981,N_24052);
xor U24917 (N_24917,N_23940,N_24024);
and U24918 (N_24918,N_24212,N_23825);
nor U24919 (N_24919,N_24248,N_24110);
xnor U24920 (N_24920,N_24241,N_24235);
and U24921 (N_24921,N_23757,N_23844);
and U24922 (N_24922,N_24336,N_24072);
and U24923 (N_24923,N_24290,N_23783);
or U24924 (N_24924,N_24175,N_24135);
nand U24925 (N_24925,N_23921,N_24141);
nand U24926 (N_24926,N_23771,N_24102);
xnor U24927 (N_24927,N_24294,N_24359);
nor U24928 (N_24928,N_23919,N_24283);
and U24929 (N_24929,N_24005,N_24222);
nor U24930 (N_24930,N_23982,N_23826);
nand U24931 (N_24931,N_24363,N_23951);
and U24932 (N_24932,N_24349,N_24007);
xnor U24933 (N_24933,N_23897,N_23782);
or U24934 (N_24934,N_23757,N_24276);
nand U24935 (N_24935,N_24268,N_24036);
or U24936 (N_24936,N_24314,N_24184);
nand U24937 (N_24937,N_23960,N_24327);
nor U24938 (N_24938,N_24029,N_24009);
xnor U24939 (N_24939,N_24264,N_23898);
xnor U24940 (N_24940,N_24042,N_23991);
and U24941 (N_24941,N_23956,N_24209);
xnor U24942 (N_24942,N_24332,N_23778);
and U24943 (N_24943,N_23805,N_23931);
or U24944 (N_24944,N_24162,N_24143);
xnor U24945 (N_24945,N_24320,N_24241);
or U24946 (N_24946,N_24024,N_24221);
nand U24947 (N_24947,N_24281,N_23917);
xnor U24948 (N_24948,N_23862,N_24356);
and U24949 (N_24949,N_23887,N_23881);
xor U24950 (N_24950,N_24328,N_23976);
nor U24951 (N_24951,N_24012,N_24158);
nor U24952 (N_24952,N_23901,N_24097);
xor U24953 (N_24953,N_24008,N_23798);
nor U24954 (N_24954,N_24004,N_24239);
and U24955 (N_24955,N_24107,N_24253);
nand U24956 (N_24956,N_24332,N_24167);
and U24957 (N_24957,N_23754,N_24029);
and U24958 (N_24958,N_23858,N_24040);
xnor U24959 (N_24959,N_24361,N_24009);
nand U24960 (N_24960,N_24350,N_24158);
nand U24961 (N_24961,N_24180,N_23907);
xnor U24962 (N_24962,N_24000,N_23777);
nor U24963 (N_24963,N_23944,N_24122);
nand U24964 (N_24964,N_24114,N_23822);
nor U24965 (N_24965,N_24066,N_24103);
nor U24966 (N_24966,N_24271,N_23779);
nor U24967 (N_24967,N_23751,N_23893);
or U24968 (N_24968,N_24363,N_24091);
nand U24969 (N_24969,N_23996,N_24006);
nand U24970 (N_24970,N_24221,N_23839);
nor U24971 (N_24971,N_24183,N_23846);
and U24972 (N_24972,N_23949,N_24038);
nor U24973 (N_24973,N_24247,N_24150);
xnor U24974 (N_24974,N_23975,N_24207);
xor U24975 (N_24975,N_24318,N_24245);
and U24976 (N_24976,N_23938,N_23833);
or U24977 (N_24977,N_23804,N_23917);
nor U24978 (N_24978,N_24134,N_24037);
nand U24979 (N_24979,N_24030,N_24041);
nor U24980 (N_24980,N_23980,N_24330);
xor U24981 (N_24981,N_23955,N_23938);
nand U24982 (N_24982,N_24025,N_24311);
xnor U24983 (N_24983,N_24265,N_24122);
nand U24984 (N_24984,N_24100,N_24088);
and U24985 (N_24985,N_24207,N_23793);
nand U24986 (N_24986,N_24108,N_23836);
or U24987 (N_24987,N_23754,N_23923);
and U24988 (N_24988,N_23859,N_23845);
nor U24989 (N_24989,N_23865,N_24032);
and U24990 (N_24990,N_24235,N_23844);
or U24991 (N_24991,N_24020,N_23866);
nor U24992 (N_24992,N_24339,N_24070);
xnor U24993 (N_24993,N_24268,N_24324);
nor U24994 (N_24994,N_24351,N_24356);
nor U24995 (N_24995,N_24195,N_23998);
nand U24996 (N_24996,N_23932,N_24101);
or U24997 (N_24997,N_24133,N_24119);
xnor U24998 (N_24998,N_23896,N_24354);
xor U24999 (N_24999,N_23820,N_23788);
nand UO_0 (O_0,N_24947,N_24593);
nor UO_1 (O_1,N_24908,N_24629);
or UO_2 (O_2,N_24594,N_24873);
nor UO_3 (O_3,N_24484,N_24399);
or UO_4 (O_4,N_24450,N_24770);
or UO_5 (O_5,N_24497,N_24452);
xor UO_6 (O_6,N_24479,N_24971);
nor UO_7 (O_7,N_24750,N_24694);
and UO_8 (O_8,N_24702,N_24490);
nor UO_9 (O_9,N_24521,N_24481);
nand UO_10 (O_10,N_24863,N_24790);
or UO_11 (O_11,N_24981,N_24675);
xnor UO_12 (O_12,N_24499,N_24639);
and UO_13 (O_13,N_24482,N_24568);
or UO_14 (O_14,N_24422,N_24591);
and UO_15 (O_15,N_24772,N_24793);
and UO_16 (O_16,N_24526,N_24607);
xnor UO_17 (O_17,N_24620,N_24931);
or UO_18 (O_18,N_24692,N_24710);
and UO_19 (O_19,N_24673,N_24705);
nor UO_20 (O_20,N_24932,N_24378);
nor UO_21 (O_21,N_24744,N_24385);
or UO_22 (O_22,N_24718,N_24666);
or UO_23 (O_23,N_24796,N_24418);
or UO_24 (O_24,N_24530,N_24782);
nand UO_25 (O_25,N_24831,N_24432);
or UO_26 (O_26,N_24738,N_24457);
nand UO_27 (O_27,N_24560,N_24676);
and UO_28 (O_28,N_24876,N_24819);
nor UO_29 (O_29,N_24402,N_24655);
nand UO_30 (O_30,N_24522,N_24935);
nor UO_31 (O_31,N_24431,N_24816);
or UO_32 (O_32,N_24534,N_24421);
nand UO_33 (O_33,N_24492,N_24466);
or UO_34 (O_34,N_24989,N_24445);
xnor UO_35 (O_35,N_24566,N_24756);
xnor UO_36 (O_36,N_24850,N_24608);
and UO_37 (O_37,N_24415,N_24952);
and UO_38 (O_38,N_24780,N_24392);
xor UO_39 (O_39,N_24730,N_24754);
nand UO_40 (O_40,N_24965,N_24985);
nor UO_41 (O_41,N_24945,N_24476);
xor UO_42 (O_42,N_24766,N_24471);
xnor UO_43 (O_43,N_24635,N_24458);
or UO_44 (O_44,N_24752,N_24595);
and UO_45 (O_45,N_24486,N_24511);
nor UO_46 (O_46,N_24740,N_24646);
or UO_47 (O_47,N_24428,N_24659);
and UO_48 (O_48,N_24930,N_24872);
nor UO_49 (O_49,N_24685,N_24441);
nor UO_50 (O_50,N_24893,N_24825);
and UO_51 (O_51,N_24890,N_24680);
nor UO_52 (O_52,N_24464,N_24609);
and UO_53 (O_53,N_24383,N_24777);
and UO_54 (O_54,N_24824,N_24689);
or UO_55 (O_55,N_24483,N_24964);
xnor UO_56 (O_56,N_24860,N_24543);
nor UO_57 (O_57,N_24882,N_24443);
xnor UO_58 (O_58,N_24943,N_24540);
xor UO_59 (O_59,N_24552,N_24918);
nor UO_60 (O_60,N_24570,N_24454);
nand UO_61 (O_61,N_24628,N_24670);
nand UO_62 (O_62,N_24884,N_24849);
nor UO_63 (O_63,N_24983,N_24791);
nand UO_64 (O_64,N_24455,N_24838);
nand UO_65 (O_65,N_24425,N_24644);
xor UO_66 (O_66,N_24697,N_24924);
nand UO_67 (O_67,N_24956,N_24732);
nand UO_68 (O_68,N_24539,N_24914);
or UO_69 (O_69,N_24827,N_24888);
or UO_70 (O_70,N_24404,N_24742);
or UO_71 (O_71,N_24653,N_24435);
and UO_72 (O_72,N_24645,N_24864);
xor UO_73 (O_73,N_24624,N_24743);
and UO_74 (O_74,N_24671,N_24892);
xor UO_75 (O_75,N_24986,N_24869);
nor UO_76 (O_76,N_24447,N_24792);
nor UO_77 (O_77,N_24800,N_24672);
nor UO_78 (O_78,N_24913,N_24717);
nor UO_79 (O_79,N_24597,N_24917);
and UO_80 (O_80,N_24919,N_24708);
and UO_81 (O_81,N_24508,N_24396);
nor UO_82 (O_82,N_24668,N_24934);
xor UO_83 (O_83,N_24895,N_24788);
or UO_84 (O_84,N_24758,N_24830);
xnor UO_85 (O_85,N_24720,N_24787);
xnor UO_86 (O_86,N_24563,N_24871);
or UO_87 (O_87,N_24386,N_24991);
nor UO_88 (O_88,N_24938,N_24546);
and UO_89 (O_89,N_24648,N_24569);
or UO_90 (O_90,N_24489,N_24974);
and UO_91 (O_91,N_24498,N_24714);
and UO_92 (O_92,N_24493,N_24683);
nor UO_93 (O_93,N_24998,N_24516);
nor UO_94 (O_94,N_24394,N_24496);
xor UO_95 (O_95,N_24937,N_24505);
nand UO_96 (O_96,N_24901,N_24783);
and UO_97 (O_97,N_24598,N_24398);
and UO_98 (O_98,N_24701,N_24604);
and UO_99 (O_99,N_24815,N_24590);
or UO_100 (O_100,N_24384,N_24564);
nor UO_101 (O_101,N_24376,N_24829);
xnor UO_102 (O_102,N_24573,N_24741);
and UO_103 (O_103,N_24746,N_24433);
or UO_104 (O_104,N_24706,N_24407);
nor UO_105 (O_105,N_24762,N_24693);
xnor UO_106 (O_106,N_24948,N_24865);
xor UO_107 (O_107,N_24465,N_24390);
xor UO_108 (O_108,N_24381,N_24536);
nor UO_109 (O_109,N_24857,N_24760);
or UO_110 (O_110,N_24468,N_24640);
nand UO_111 (O_111,N_24669,N_24870);
or UO_112 (O_112,N_24520,N_24695);
or UO_113 (O_113,N_24423,N_24518);
or UO_114 (O_114,N_24627,N_24388);
nor UO_115 (O_115,N_24529,N_24707);
xor UO_116 (O_116,N_24663,N_24515);
and UO_117 (O_117,N_24904,N_24618);
and UO_118 (O_118,N_24665,N_24773);
and UO_119 (O_119,N_24549,N_24592);
or UO_120 (O_120,N_24656,N_24583);
nand UO_121 (O_121,N_24649,N_24400);
or UO_122 (O_122,N_24711,N_24678);
and UO_123 (O_123,N_24774,N_24939);
or UO_124 (O_124,N_24531,N_24726);
xnor UO_125 (O_125,N_24467,N_24963);
and UO_126 (O_126,N_24703,N_24719);
nor UO_127 (O_127,N_24581,N_24996);
or UO_128 (O_128,N_24734,N_24619);
nor UO_129 (O_129,N_24761,N_24387);
nand UO_130 (O_130,N_24621,N_24833);
and UO_131 (O_131,N_24571,N_24941);
nand UO_132 (O_132,N_24453,N_24973);
nor UO_133 (O_133,N_24554,N_24839);
nand UO_134 (O_134,N_24537,N_24955);
and UO_135 (O_135,N_24915,N_24843);
and UO_136 (O_136,N_24379,N_24419);
nand UO_137 (O_137,N_24958,N_24690);
xnor UO_138 (O_138,N_24451,N_24854);
xor UO_139 (O_139,N_24514,N_24555);
or UO_140 (O_140,N_24954,N_24634);
or UO_141 (O_141,N_24551,N_24686);
and UO_142 (O_142,N_24507,N_24887);
or UO_143 (O_143,N_24840,N_24562);
xnor UO_144 (O_144,N_24699,N_24764);
or UO_145 (O_145,N_24512,N_24897);
nand UO_146 (O_146,N_24970,N_24812);
xor UO_147 (O_147,N_24959,N_24643);
nand UO_148 (O_148,N_24894,N_24736);
or UO_149 (O_149,N_24667,N_24900);
or UO_150 (O_150,N_24929,N_24962);
or UO_151 (O_151,N_24709,N_24821);
or UO_152 (O_152,N_24927,N_24802);
xnor UO_153 (O_153,N_24920,N_24757);
and UO_154 (O_154,N_24911,N_24978);
nand UO_155 (O_155,N_24995,N_24704);
xnor UO_156 (O_156,N_24579,N_24382);
and UO_157 (O_157,N_24747,N_24698);
or UO_158 (O_158,N_24818,N_24679);
nor UO_159 (O_159,N_24949,N_24556);
nand UO_160 (O_160,N_24874,N_24784);
nor UO_161 (O_161,N_24377,N_24632);
or UO_162 (O_162,N_24565,N_24687);
or UO_163 (O_163,N_24866,N_24462);
nand UO_164 (O_164,N_24406,N_24605);
nor UO_165 (O_165,N_24999,N_24763);
nand UO_166 (O_166,N_24807,N_24828);
nor UO_167 (O_167,N_24391,N_24826);
or UO_168 (O_168,N_24994,N_24416);
and UO_169 (O_169,N_24889,N_24805);
and UO_170 (O_170,N_24688,N_24622);
and UO_171 (O_171,N_24808,N_24885);
nor UO_172 (O_172,N_24841,N_24380);
xor UO_173 (O_173,N_24735,N_24724);
or UO_174 (O_174,N_24559,N_24944);
nor UO_175 (O_175,N_24868,N_24879);
xor UO_176 (O_176,N_24633,N_24681);
or UO_177 (O_177,N_24910,N_24631);
or UO_178 (O_178,N_24501,N_24960);
xnor UO_179 (O_179,N_24519,N_24528);
and UO_180 (O_180,N_24982,N_24584);
or UO_181 (O_181,N_24713,N_24523);
or UO_182 (O_182,N_24405,N_24538);
xor UO_183 (O_183,N_24611,N_24936);
and UO_184 (O_184,N_24651,N_24532);
nand UO_185 (O_185,N_24961,N_24811);
or UO_186 (O_186,N_24424,N_24438);
xnor UO_187 (O_187,N_24980,N_24737);
nand UO_188 (O_188,N_24596,N_24755);
nand UO_189 (O_189,N_24733,N_24923);
xnor UO_190 (O_190,N_24775,N_24728);
nor UO_191 (O_191,N_24798,N_24420);
and UO_192 (O_192,N_24636,N_24469);
nor UO_193 (O_193,N_24968,N_24558);
nand UO_194 (O_194,N_24846,N_24485);
and UO_195 (O_195,N_24925,N_24660);
nor UO_196 (O_196,N_24436,N_24557);
xnor UO_197 (O_197,N_24801,N_24967);
nand UO_198 (O_198,N_24535,N_24842);
nor UO_199 (O_199,N_24395,N_24448);
and UO_200 (O_200,N_24542,N_24567);
and UO_201 (O_201,N_24411,N_24822);
or UO_202 (O_202,N_24778,N_24856);
nor UO_203 (O_203,N_24753,N_24969);
and UO_204 (O_204,N_24461,N_24647);
or UO_205 (O_205,N_24427,N_24606);
or UO_206 (O_206,N_24577,N_24806);
or UO_207 (O_207,N_24617,N_24550);
nor UO_208 (O_208,N_24859,N_24661);
or UO_209 (O_209,N_24921,N_24877);
or UO_210 (O_210,N_24545,N_24823);
xnor UO_211 (O_211,N_24899,N_24853);
and UO_212 (O_212,N_24510,N_24613);
nor UO_213 (O_213,N_24883,N_24771);
nor UO_214 (O_214,N_24898,N_24803);
or UO_215 (O_215,N_24674,N_24861);
xnor UO_216 (O_216,N_24582,N_24623);
and UO_217 (O_217,N_24615,N_24933);
and UO_218 (O_218,N_24979,N_24765);
nor UO_219 (O_219,N_24804,N_24642);
or UO_220 (O_220,N_24503,N_24797);
nor UO_221 (O_221,N_24715,N_24767);
nand UO_222 (O_222,N_24928,N_24414);
xor UO_223 (O_223,N_24727,N_24723);
or UO_224 (O_224,N_24602,N_24813);
and UO_225 (O_225,N_24957,N_24662);
xnor UO_226 (O_226,N_24942,N_24814);
and UO_227 (O_227,N_24657,N_24578);
nand UO_228 (O_228,N_24972,N_24525);
and UO_229 (O_229,N_24886,N_24691);
and UO_230 (O_230,N_24652,N_24601);
nand UO_231 (O_231,N_24459,N_24474);
or UO_232 (O_232,N_24940,N_24553);
xor UO_233 (O_233,N_24739,N_24906);
nor UO_234 (O_234,N_24412,N_24463);
nor UO_235 (O_235,N_24729,N_24951);
nor UO_236 (O_236,N_24878,N_24475);
nor UO_237 (O_237,N_24907,N_24835);
xor UO_238 (O_238,N_24544,N_24408);
nand UO_239 (O_239,N_24988,N_24527);
xnor UO_240 (O_240,N_24851,N_24480);
and UO_241 (O_241,N_24781,N_24891);
or UO_242 (O_242,N_24905,N_24587);
or UO_243 (O_243,N_24682,N_24575);
and UO_244 (O_244,N_24820,N_24614);
and UO_245 (O_245,N_24588,N_24446);
or UO_246 (O_246,N_24426,N_24848);
xor UO_247 (O_247,N_24413,N_24610);
and UO_248 (O_248,N_24456,N_24700);
nand UO_249 (O_249,N_24776,N_24844);
nor UO_250 (O_250,N_24903,N_24616);
xnor UO_251 (O_251,N_24799,N_24795);
and UO_252 (O_252,N_24576,N_24997);
xor UO_253 (O_253,N_24902,N_24495);
or UO_254 (O_254,N_24855,N_24502);
nand UO_255 (O_255,N_24880,N_24789);
nor UO_256 (O_256,N_24442,N_24867);
nor UO_257 (O_257,N_24984,N_24430);
xor UO_258 (O_258,N_24975,N_24524);
xnor UO_259 (O_259,N_24990,N_24832);
nand UO_260 (O_260,N_24429,N_24712);
nor UO_261 (O_261,N_24417,N_24722);
nand UO_262 (O_262,N_24494,N_24513);
and UO_263 (O_263,N_24836,N_24547);
nor UO_264 (O_264,N_24768,N_24460);
or UO_265 (O_265,N_24946,N_24637);
nand UO_266 (O_266,N_24779,N_24858);
or UO_267 (O_267,N_24852,N_24477);
nand UO_268 (O_268,N_24664,N_24487);
nand UO_269 (O_269,N_24916,N_24731);
xor UO_270 (O_270,N_24834,N_24769);
xnor UO_271 (O_271,N_24600,N_24574);
or UO_272 (O_272,N_24389,N_24572);
xor UO_273 (O_273,N_24953,N_24794);
nor UO_274 (O_274,N_24725,N_24397);
nor UO_275 (O_275,N_24875,N_24992);
and UO_276 (O_276,N_24401,N_24654);
nand UO_277 (O_277,N_24410,N_24817);
and UO_278 (O_278,N_24548,N_24603);
nor UO_279 (O_279,N_24478,N_24409);
nand UO_280 (O_280,N_24439,N_24589);
and UO_281 (O_281,N_24950,N_24977);
and UO_282 (O_282,N_24403,N_24626);
nor UO_283 (O_283,N_24922,N_24745);
xor UO_284 (O_284,N_24912,N_24966);
nand UO_285 (O_285,N_24437,N_24785);
xnor UO_286 (O_286,N_24500,N_24580);
and UO_287 (O_287,N_24881,N_24488);
nand UO_288 (O_288,N_24585,N_24491);
nand UO_289 (O_289,N_24759,N_24896);
nor UO_290 (O_290,N_24625,N_24976);
or UO_291 (O_291,N_24641,N_24586);
or UO_292 (O_292,N_24749,N_24449);
and UO_293 (O_293,N_24517,N_24599);
nand UO_294 (O_294,N_24440,N_24638);
and UO_295 (O_295,N_24473,N_24716);
and UO_296 (O_296,N_24472,N_24444);
nand UO_297 (O_297,N_24393,N_24926);
nand UO_298 (O_298,N_24470,N_24786);
and UO_299 (O_299,N_24509,N_24810);
nor UO_300 (O_300,N_24751,N_24862);
xnor UO_301 (O_301,N_24847,N_24809);
and UO_302 (O_302,N_24677,N_24612);
nor UO_303 (O_303,N_24541,N_24748);
nor UO_304 (O_304,N_24658,N_24375);
nand UO_305 (O_305,N_24987,N_24696);
xor UO_306 (O_306,N_24533,N_24561);
and UO_307 (O_307,N_24504,N_24684);
nand UO_308 (O_308,N_24650,N_24434);
nor UO_309 (O_309,N_24506,N_24837);
or UO_310 (O_310,N_24845,N_24721);
xnor UO_311 (O_311,N_24909,N_24630);
nand UO_312 (O_312,N_24993,N_24753);
xor UO_313 (O_313,N_24901,N_24706);
and UO_314 (O_314,N_24934,N_24688);
or UO_315 (O_315,N_24924,N_24810);
xor UO_316 (O_316,N_24759,N_24466);
xor UO_317 (O_317,N_24819,N_24969);
xnor UO_318 (O_318,N_24921,N_24475);
and UO_319 (O_319,N_24633,N_24830);
nand UO_320 (O_320,N_24888,N_24700);
nor UO_321 (O_321,N_24769,N_24727);
or UO_322 (O_322,N_24803,N_24598);
nor UO_323 (O_323,N_24561,N_24438);
xor UO_324 (O_324,N_24932,N_24961);
xnor UO_325 (O_325,N_24389,N_24430);
xnor UO_326 (O_326,N_24636,N_24749);
xnor UO_327 (O_327,N_24433,N_24584);
xor UO_328 (O_328,N_24690,N_24695);
xnor UO_329 (O_329,N_24780,N_24685);
nand UO_330 (O_330,N_24725,N_24514);
xor UO_331 (O_331,N_24655,N_24612);
nand UO_332 (O_332,N_24539,N_24416);
and UO_333 (O_333,N_24972,N_24612);
xnor UO_334 (O_334,N_24901,N_24815);
nor UO_335 (O_335,N_24887,N_24963);
and UO_336 (O_336,N_24572,N_24758);
or UO_337 (O_337,N_24773,N_24730);
and UO_338 (O_338,N_24418,N_24900);
xnor UO_339 (O_339,N_24459,N_24513);
xnor UO_340 (O_340,N_24493,N_24650);
nor UO_341 (O_341,N_24845,N_24834);
or UO_342 (O_342,N_24865,N_24694);
and UO_343 (O_343,N_24814,N_24442);
nor UO_344 (O_344,N_24701,N_24430);
and UO_345 (O_345,N_24895,N_24912);
or UO_346 (O_346,N_24969,N_24974);
nand UO_347 (O_347,N_24592,N_24981);
nand UO_348 (O_348,N_24891,N_24416);
xnor UO_349 (O_349,N_24823,N_24514);
and UO_350 (O_350,N_24905,N_24470);
nand UO_351 (O_351,N_24593,N_24537);
nor UO_352 (O_352,N_24554,N_24994);
and UO_353 (O_353,N_24985,N_24706);
and UO_354 (O_354,N_24755,N_24881);
nand UO_355 (O_355,N_24595,N_24679);
xnor UO_356 (O_356,N_24444,N_24411);
xnor UO_357 (O_357,N_24843,N_24534);
nand UO_358 (O_358,N_24981,N_24797);
and UO_359 (O_359,N_24730,N_24786);
nand UO_360 (O_360,N_24546,N_24660);
nor UO_361 (O_361,N_24390,N_24955);
or UO_362 (O_362,N_24819,N_24604);
and UO_363 (O_363,N_24975,N_24544);
and UO_364 (O_364,N_24541,N_24465);
nand UO_365 (O_365,N_24738,N_24420);
xor UO_366 (O_366,N_24686,N_24940);
xnor UO_367 (O_367,N_24794,N_24435);
nor UO_368 (O_368,N_24826,N_24980);
nor UO_369 (O_369,N_24402,N_24485);
nand UO_370 (O_370,N_24924,N_24601);
xnor UO_371 (O_371,N_24888,N_24607);
or UO_372 (O_372,N_24858,N_24810);
nand UO_373 (O_373,N_24619,N_24391);
nand UO_374 (O_374,N_24763,N_24672);
or UO_375 (O_375,N_24999,N_24375);
or UO_376 (O_376,N_24997,N_24475);
or UO_377 (O_377,N_24627,N_24941);
xnor UO_378 (O_378,N_24482,N_24691);
nand UO_379 (O_379,N_24500,N_24527);
nand UO_380 (O_380,N_24390,N_24876);
nand UO_381 (O_381,N_24832,N_24661);
or UO_382 (O_382,N_24719,N_24849);
xnor UO_383 (O_383,N_24923,N_24793);
or UO_384 (O_384,N_24405,N_24758);
or UO_385 (O_385,N_24705,N_24980);
nand UO_386 (O_386,N_24427,N_24970);
xor UO_387 (O_387,N_24663,N_24435);
and UO_388 (O_388,N_24520,N_24467);
nor UO_389 (O_389,N_24390,N_24681);
or UO_390 (O_390,N_24801,N_24559);
xor UO_391 (O_391,N_24827,N_24553);
nand UO_392 (O_392,N_24680,N_24868);
or UO_393 (O_393,N_24625,N_24893);
and UO_394 (O_394,N_24375,N_24468);
xnor UO_395 (O_395,N_24433,N_24853);
xor UO_396 (O_396,N_24432,N_24552);
and UO_397 (O_397,N_24556,N_24970);
xnor UO_398 (O_398,N_24844,N_24710);
xor UO_399 (O_399,N_24713,N_24803);
and UO_400 (O_400,N_24428,N_24831);
nor UO_401 (O_401,N_24519,N_24850);
xnor UO_402 (O_402,N_24898,N_24745);
or UO_403 (O_403,N_24914,N_24990);
and UO_404 (O_404,N_24676,N_24535);
or UO_405 (O_405,N_24414,N_24722);
and UO_406 (O_406,N_24826,N_24851);
xor UO_407 (O_407,N_24575,N_24964);
or UO_408 (O_408,N_24522,N_24745);
xnor UO_409 (O_409,N_24405,N_24749);
or UO_410 (O_410,N_24863,N_24477);
nand UO_411 (O_411,N_24417,N_24665);
nand UO_412 (O_412,N_24562,N_24507);
or UO_413 (O_413,N_24759,N_24379);
nor UO_414 (O_414,N_24940,N_24769);
and UO_415 (O_415,N_24925,N_24544);
or UO_416 (O_416,N_24501,N_24538);
or UO_417 (O_417,N_24731,N_24849);
and UO_418 (O_418,N_24849,N_24625);
or UO_419 (O_419,N_24976,N_24698);
and UO_420 (O_420,N_24810,N_24692);
nor UO_421 (O_421,N_24940,N_24562);
nor UO_422 (O_422,N_24872,N_24839);
nor UO_423 (O_423,N_24445,N_24440);
xor UO_424 (O_424,N_24562,N_24402);
xor UO_425 (O_425,N_24740,N_24827);
and UO_426 (O_426,N_24439,N_24744);
nor UO_427 (O_427,N_24553,N_24963);
and UO_428 (O_428,N_24804,N_24620);
nor UO_429 (O_429,N_24867,N_24875);
or UO_430 (O_430,N_24823,N_24834);
nand UO_431 (O_431,N_24391,N_24521);
nor UO_432 (O_432,N_24504,N_24390);
or UO_433 (O_433,N_24395,N_24811);
or UO_434 (O_434,N_24735,N_24469);
nand UO_435 (O_435,N_24761,N_24537);
or UO_436 (O_436,N_24979,N_24432);
nor UO_437 (O_437,N_24423,N_24404);
and UO_438 (O_438,N_24950,N_24875);
nand UO_439 (O_439,N_24755,N_24387);
or UO_440 (O_440,N_24574,N_24914);
nor UO_441 (O_441,N_24591,N_24533);
xor UO_442 (O_442,N_24833,N_24817);
or UO_443 (O_443,N_24603,N_24503);
and UO_444 (O_444,N_24878,N_24474);
xor UO_445 (O_445,N_24987,N_24536);
and UO_446 (O_446,N_24459,N_24793);
nor UO_447 (O_447,N_24871,N_24462);
or UO_448 (O_448,N_24380,N_24739);
and UO_449 (O_449,N_24541,N_24487);
nor UO_450 (O_450,N_24705,N_24635);
xnor UO_451 (O_451,N_24379,N_24602);
and UO_452 (O_452,N_24814,N_24959);
xnor UO_453 (O_453,N_24605,N_24760);
xnor UO_454 (O_454,N_24894,N_24956);
nor UO_455 (O_455,N_24436,N_24432);
nand UO_456 (O_456,N_24661,N_24589);
nand UO_457 (O_457,N_24583,N_24398);
and UO_458 (O_458,N_24898,N_24379);
nand UO_459 (O_459,N_24588,N_24683);
and UO_460 (O_460,N_24677,N_24731);
nor UO_461 (O_461,N_24520,N_24988);
or UO_462 (O_462,N_24782,N_24550);
nand UO_463 (O_463,N_24564,N_24702);
and UO_464 (O_464,N_24758,N_24818);
xor UO_465 (O_465,N_24430,N_24938);
and UO_466 (O_466,N_24915,N_24802);
xor UO_467 (O_467,N_24888,N_24871);
and UO_468 (O_468,N_24694,N_24706);
nor UO_469 (O_469,N_24711,N_24809);
and UO_470 (O_470,N_24879,N_24445);
and UO_471 (O_471,N_24930,N_24742);
and UO_472 (O_472,N_24400,N_24570);
nor UO_473 (O_473,N_24426,N_24989);
nor UO_474 (O_474,N_24625,N_24970);
nand UO_475 (O_475,N_24729,N_24836);
nor UO_476 (O_476,N_24857,N_24989);
nand UO_477 (O_477,N_24415,N_24948);
and UO_478 (O_478,N_24541,N_24635);
nor UO_479 (O_479,N_24390,N_24748);
xor UO_480 (O_480,N_24561,N_24485);
and UO_481 (O_481,N_24530,N_24998);
xnor UO_482 (O_482,N_24724,N_24828);
nand UO_483 (O_483,N_24398,N_24496);
xor UO_484 (O_484,N_24998,N_24625);
and UO_485 (O_485,N_24764,N_24467);
nor UO_486 (O_486,N_24476,N_24533);
nand UO_487 (O_487,N_24862,N_24379);
nand UO_488 (O_488,N_24583,N_24406);
nor UO_489 (O_489,N_24393,N_24693);
and UO_490 (O_490,N_24726,N_24699);
xor UO_491 (O_491,N_24851,N_24707);
and UO_492 (O_492,N_24899,N_24712);
xor UO_493 (O_493,N_24680,N_24878);
xnor UO_494 (O_494,N_24378,N_24819);
nor UO_495 (O_495,N_24427,N_24918);
or UO_496 (O_496,N_24708,N_24863);
nor UO_497 (O_497,N_24450,N_24418);
or UO_498 (O_498,N_24514,N_24466);
nor UO_499 (O_499,N_24477,N_24590);
or UO_500 (O_500,N_24598,N_24557);
nor UO_501 (O_501,N_24575,N_24392);
and UO_502 (O_502,N_24671,N_24945);
or UO_503 (O_503,N_24698,N_24446);
or UO_504 (O_504,N_24861,N_24497);
nor UO_505 (O_505,N_24868,N_24713);
nor UO_506 (O_506,N_24846,N_24458);
and UO_507 (O_507,N_24975,N_24610);
nand UO_508 (O_508,N_24453,N_24450);
and UO_509 (O_509,N_24661,N_24856);
and UO_510 (O_510,N_24911,N_24816);
nor UO_511 (O_511,N_24899,N_24644);
and UO_512 (O_512,N_24877,N_24920);
nand UO_513 (O_513,N_24864,N_24460);
xnor UO_514 (O_514,N_24802,N_24826);
nand UO_515 (O_515,N_24762,N_24621);
nor UO_516 (O_516,N_24454,N_24829);
or UO_517 (O_517,N_24749,N_24404);
nor UO_518 (O_518,N_24754,N_24662);
xnor UO_519 (O_519,N_24757,N_24423);
nor UO_520 (O_520,N_24785,N_24588);
xor UO_521 (O_521,N_24787,N_24723);
nand UO_522 (O_522,N_24603,N_24400);
and UO_523 (O_523,N_24593,N_24743);
nand UO_524 (O_524,N_24967,N_24825);
and UO_525 (O_525,N_24629,N_24743);
xor UO_526 (O_526,N_24617,N_24713);
nand UO_527 (O_527,N_24549,N_24755);
nand UO_528 (O_528,N_24792,N_24824);
nand UO_529 (O_529,N_24376,N_24590);
or UO_530 (O_530,N_24619,N_24968);
and UO_531 (O_531,N_24799,N_24843);
or UO_532 (O_532,N_24622,N_24820);
or UO_533 (O_533,N_24518,N_24645);
nor UO_534 (O_534,N_24578,N_24750);
nand UO_535 (O_535,N_24968,N_24825);
or UO_536 (O_536,N_24938,N_24625);
and UO_537 (O_537,N_24624,N_24952);
nand UO_538 (O_538,N_24861,N_24931);
or UO_539 (O_539,N_24489,N_24562);
nor UO_540 (O_540,N_24945,N_24822);
xnor UO_541 (O_541,N_24760,N_24771);
xor UO_542 (O_542,N_24378,N_24685);
xor UO_543 (O_543,N_24869,N_24756);
and UO_544 (O_544,N_24687,N_24577);
and UO_545 (O_545,N_24900,N_24786);
and UO_546 (O_546,N_24728,N_24396);
nor UO_547 (O_547,N_24812,N_24512);
xnor UO_548 (O_548,N_24734,N_24519);
nand UO_549 (O_549,N_24626,N_24597);
xor UO_550 (O_550,N_24506,N_24443);
nor UO_551 (O_551,N_24472,N_24788);
xor UO_552 (O_552,N_24682,N_24557);
xnor UO_553 (O_553,N_24551,N_24487);
nor UO_554 (O_554,N_24533,N_24526);
xor UO_555 (O_555,N_24957,N_24663);
or UO_556 (O_556,N_24941,N_24825);
or UO_557 (O_557,N_24967,N_24833);
or UO_558 (O_558,N_24634,N_24732);
nor UO_559 (O_559,N_24710,N_24795);
nor UO_560 (O_560,N_24914,N_24577);
and UO_561 (O_561,N_24971,N_24956);
nand UO_562 (O_562,N_24660,N_24565);
nor UO_563 (O_563,N_24485,N_24560);
nand UO_564 (O_564,N_24512,N_24992);
nor UO_565 (O_565,N_24807,N_24516);
and UO_566 (O_566,N_24704,N_24660);
and UO_567 (O_567,N_24836,N_24647);
xnor UO_568 (O_568,N_24729,N_24537);
nand UO_569 (O_569,N_24819,N_24453);
xnor UO_570 (O_570,N_24853,N_24833);
and UO_571 (O_571,N_24672,N_24687);
and UO_572 (O_572,N_24421,N_24784);
or UO_573 (O_573,N_24412,N_24781);
nand UO_574 (O_574,N_24603,N_24777);
or UO_575 (O_575,N_24510,N_24947);
and UO_576 (O_576,N_24711,N_24998);
nor UO_577 (O_577,N_24763,N_24986);
and UO_578 (O_578,N_24883,N_24734);
nand UO_579 (O_579,N_24669,N_24836);
and UO_580 (O_580,N_24871,N_24865);
nand UO_581 (O_581,N_24551,N_24889);
nand UO_582 (O_582,N_24550,N_24603);
nor UO_583 (O_583,N_24840,N_24701);
nand UO_584 (O_584,N_24898,N_24856);
xor UO_585 (O_585,N_24466,N_24743);
or UO_586 (O_586,N_24461,N_24688);
xor UO_587 (O_587,N_24764,N_24860);
nor UO_588 (O_588,N_24913,N_24723);
nor UO_589 (O_589,N_24382,N_24959);
xor UO_590 (O_590,N_24484,N_24966);
nand UO_591 (O_591,N_24655,N_24830);
xnor UO_592 (O_592,N_24541,N_24599);
xnor UO_593 (O_593,N_24707,N_24503);
or UO_594 (O_594,N_24588,N_24640);
nor UO_595 (O_595,N_24673,N_24603);
nand UO_596 (O_596,N_24705,N_24525);
nor UO_597 (O_597,N_24942,N_24728);
nor UO_598 (O_598,N_24379,N_24952);
nand UO_599 (O_599,N_24861,N_24995);
xor UO_600 (O_600,N_24484,N_24701);
xnor UO_601 (O_601,N_24670,N_24795);
nand UO_602 (O_602,N_24644,N_24825);
xor UO_603 (O_603,N_24530,N_24794);
xnor UO_604 (O_604,N_24632,N_24518);
nor UO_605 (O_605,N_24442,N_24875);
or UO_606 (O_606,N_24909,N_24441);
and UO_607 (O_607,N_24812,N_24746);
nand UO_608 (O_608,N_24694,N_24763);
and UO_609 (O_609,N_24836,N_24888);
and UO_610 (O_610,N_24517,N_24705);
nand UO_611 (O_611,N_24992,N_24779);
nand UO_612 (O_612,N_24950,N_24738);
nand UO_613 (O_613,N_24582,N_24756);
nor UO_614 (O_614,N_24830,N_24778);
and UO_615 (O_615,N_24400,N_24893);
nor UO_616 (O_616,N_24610,N_24884);
nor UO_617 (O_617,N_24695,N_24656);
xnor UO_618 (O_618,N_24857,N_24930);
nor UO_619 (O_619,N_24503,N_24897);
xnor UO_620 (O_620,N_24953,N_24738);
or UO_621 (O_621,N_24668,N_24972);
xor UO_622 (O_622,N_24375,N_24504);
or UO_623 (O_623,N_24651,N_24972);
nand UO_624 (O_624,N_24882,N_24931);
or UO_625 (O_625,N_24885,N_24975);
and UO_626 (O_626,N_24938,N_24380);
xnor UO_627 (O_627,N_24701,N_24896);
xnor UO_628 (O_628,N_24636,N_24376);
xor UO_629 (O_629,N_24673,N_24836);
xnor UO_630 (O_630,N_24623,N_24375);
nand UO_631 (O_631,N_24572,N_24980);
xnor UO_632 (O_632,N_24994,N_24903);
or UO_633 (O_633,N_24924,N_24981);
nand UO_634 (O_634,N_24867,N_24421);
xor UO_635 (O_635,N_24411,N_24428);
or UO_636 (O_636,N_24971,N_24910);
or UO_637 (O_637,N_24476,N_24855);
and UO_638 (O_638,N_24643,N_24861);
xor UO_639 (O_639,N_24858,N_24622);
nor UO_640 (O_640,N_24412,N_24515);
and UO_641 (O_641,N_24532,N_24457);
and UO_642 (O_642,N_24955,N_24839);
nand UO_643 (O_643,N_24583,N_24819);
xnor UO_644 (O_644,N_24884,N_24465);
xor UO_645 (O_645,N_24681,N_24672);
nand UO_646 (O_646,N_24904,N_24411);
xor UO_647 (O_647,N_24453,N_24503);
or UO_648 (O_648,N_24701,N_24799);
or UO_649 (O_649,N_24679,N_24402);
nand UO_650 (O_650,N_24805,N_24848);
and UO_651 (O_651,N_24460,N_24945);
nor UO_652 (O_652,N_24963,N_24531);
nor UO_653 (O_653,N_24425,N_24574);
nand UO_654 (O_654,N_24695,N_24706);
xor UO_655 (O_655,N_24640,N_24850);
xor UO_656 (O_656,N_24456,N_24870);
nand UO_657 (O_657,N_24716,N_24499);
and UO_658 (O_658,N_24743,N_24456);
nand UO_659 (O_659,N_24743,N_24586);
xor UO_660 (O_660,N_24438,N_24774);
and UO_661 (O_661,N_24744,N_24641);
or UO_662 (O_662,N_24975,N_24720);
nor UO_663 (O_663,N_24982,N_24853);
and UO_664 (O_664,N_24781,N_24717);
or UO_665 (O_665,N_24605,N_24742);
nor UO_666 (O_666,N_24532,N_24627);
or UO_667 (O_667,N_24750,N_24586);
or UO_668 (O_668,N_24852,N_24428);
and UO_669 (O_669,N_24410,N_24513);
and UO_670 (O_670,N_24913,N_24896);
or UO_671 (O_671,N_24655,N_24606);
nor UO_672 (O_672,N_24420,N_24573);
nand UO_673 (O_673,N_24615,N_24872);
xnor UO_674 (O_674,N_24853,N_24384);
nor UO_675 (O_675,N_24660,N_24976);
and UO_676 (O_676,N_24376,N_24816);
xnor UO_677 (O_677,N_24581,N_24563);
nor UO_678 (O_678,N_24737,N_24907);
and UO_679 (O_679,N_24426,N_24590);
xor UO_680 (O_680,N_24388,N_24423);
nand UO_681 (O_681,N_24921,N_24774);
xor UO_682 (O_682,N_24423,N_24800);
nor UO_683 (O_683,N_24979,N_24409);
or UO_684 (O_684,N_24547,N_24454);
xor UO_685 (O_685,N_24528,N_24552);
nand UO_686 (O_686,N_24446,N_24892);
nor UO_687 (O_687,N_24841,N_24824);
or UO_688 (O_688,N_24494,N_24871);
xnor UO_689 (O_689,N_24728,N_24424);
and UO_690 (O_690,N_24993,N_24939);
nor UO_691 (O_691,N_24967,N_24595);
nor UO_692 (O_692,N_24881,N_24966);
nand UO_693 (O_693,N_24853,N_24761);
xor UO_694 (O_694,N_24426,N_24604);
and UO_695 (O_695,N_24787,N_24877);
xnor UO_696 (O_696,N_24903,N_24976);
nor UO_697 (O_697,N_24805,N_24426);
and UO_698 (O_698,N_24794,N_24590);
nor UO_699 (O_699,N_24863,N_24491);
nor UO_700 (O_700,N_24914,N_24773);
nor UO_701 (O_701,N_24446,N_24625);
nor UO_702 (O_702,N_24893,N_24535);
nor UO_703 (O_703,N_24651,N_24792);
and UO_704 (O_704,N_24774,N_24740);
or UO_705 (O_705,N_24899,N_24816);
xnor UO_706 (O_706,N_24963,N_24596);
xnor UO_707 (O_707,N_24386,N_24720);
or UO_708 (O_708,N_24660,N_24798);
and UO_709 (O_709,N_24483,N_24395);
xnor UO_710 (O_710,N_24825,N_24453);
nor UO_711 (O_711,N_24518,N_24840);
nor UO_712 (O_712,N_24576,N_24599);
or UO_713 (O_713,N_24784,N_24412);
and UO_714 (O_714,N_24684,N_24807);
xnor UO_715 (O_715,N_24926,N_24428);
xnor UO_716 (O_716,N_24552,N_24746);
xnor UO_717 (O_717,N_24619,N_24585);
xnor UO_718 (O_718,N_24737,N_24438);
or UO_719 (O_719,N_24795,N_24617);
xnor UO_720 (O_720,N_24799,N_24482);
nand UO_721 (O_721,N_24949,N_24668);
nor UO_722 (O_722,N_24650,N_24571);
nor UO_723 (O_723,N_24588,N_24755);
nor UO_724 (O_724,N_24413,N_24952);
or UO_725 (O_725,N_24792,N_24571);
nand UO_726 (O_726,N_24441,N_24927);
nor UO_727 (O_727,N_24774,N_24865);
and UO_728 (O_728,N_24913,N_24538);
nor UO_729 (O_729,N_24955,N_24792);
and UO_730 (O_730,N_24778,N_24731);
xnor UO_731 (O_731,N_24695,N_24483);
or UO_732 (O_732,N_24638,N_24811);
and UO_733 (O_733,N_24600,N_24547);
xor UO_734 (O_734,N_24430,N_24606);
nor UO_735 (O_735,N_24930,N_24785);
nor UO_736 (O_736,N_24485,N_24414);
and UO_737 (O_737,N_24530,N_24936);
nand UO_738 (O_738,N_24982,N_24464);
nand UO_739 (O_739,N_24663,N_24502);
or UO_740 (O_740,N_24617,N_24749);
xnor UO_741 (O_741,N_24981,N_24404);
and UO_742 (O_742,N_24975,N_24649);
and UO_743 (O_743,N_24392,N_24556);
nor UO_744 (O_744,N_24622,N_24588);
and UO_745 (O_745,N_24922,N_24382);
nand UO_746 (O_746,N_24507,N_24757);
and UO_747 (O_747,N_24710,N_24805);
nor UO_748 (O_748,N_24630,N_24995);
or UO_749 (O_749,N_24566,N_24452);
or UO_750 (O_750,N_24646,N_24423);
or UO_751 (O_751,N_24996,N_24624);
and UO_752 (O_752,N_24841,N_24802);
nor UO_753 (O_753,N_24934,N_24845);
and UO_754 (O_754,N_24987,N_24909);
nand UO_755 (O_755,N_24471,N_24457);
xor UO_756 (O_756,N_24671,N_24767);
nor UO_757 (O_757,N_24672,N_24834);
or UO_758 (O_758,N_24548,N_24686);
nand UO_759 (O_759,N_24799,N_24905);
nor UO_760 (O_760,N_24697,N_24596);
nand UO_761 (O_761,N_24607,N_24509);
nor UO_762 (O_762,N_24446,N_24804);
nand UO_763 (O_763,N_24423,N_24632);
and UO_764 (O_764,N_24876,N_24770);
and UO_765 (O_765,N_24612,N_24787);
xor UO_766 (O_766,N_24379,N_24778);
or UO_767 (O_767,N_24745,N_24990);
and UO_768 (O_768,N_24707,N_24636);
or UO_769 (O_769,N_24618,N_24403);
or UO_770 (O_770,N_24663,N_24938);
and UO_771 (O_771,N_24976,N_24920);
nand UO_772 (O_772,N_24773,N_24388);
nor UO_773 (O_773,N_24682,N_24849);
and UO_774 (O_774,N_24802,N_24997);
or UO_775 (O_775,N_24761,N_24617);
or UO_776 (O_776,N_24635,N_24617);
or UO_777 (O_777,N_24723,N_24898);
or UO_778 (O_778,N_24438,N_24712);
xnor UO_779 (O_779,N_24610,N_24950);
xor UO_780 (O_780,N_24668,N_24861);
nand UO_781 (O_781,N_24945,N_24562);
nand UO_782 (O_782,N_24970,N_24936);
xnor UO_783 (O_783,N_24715,N_24807);
or UO_784 (O_784,N_24586,N_24680);
nand UO_785 (O_785,N_24765,N_24736);
nand UO_786 (O_786,N_24949,N_24812);
nor UO_787 (O_787,N_24962,N_24540);
nor UO_788 (O_788,N_24739,N_24709);
nor UO_789 (O_789,N_24659,N_24420);
xor UO_790 (O_790,N_24924,N_24930);
xor UO_791 (O_791,N_24497,N_24594);
xnor UO_792 (O_792,N_24593,N_24515);
or UO_793 (O_793,N_24906,N_24490);
nor UO_794 (O_794,N_24436,N_24556);
or UO_795 (O_795,N_24829,N_24704);
or UO_796 (O_796,N_24590,N_24767);
nand UO_797 (O_797,N_24855,N_24735);
xor UO_798 (O_798,N_24581,N_24414);
and UO_799 (O_799,N_24451,N_24596);
or UO_800 (O_800,N_24777,N_24887);
and UO_801 (O_801,N_24920,N_24911);
and UO_802 (O_802,N_24906,N_24467);
nand UO_803 (O_803,N_24974,N_24700);
nand UO_804 (O_804,N_24996,N_24419);
xnor UO_805 (O_805,N_24464,N_24726);
or UO_806 (O_806,N_24428,N_24868);
xor UO_807 (O_807,N_24722,N_24733);
nor UO_808 (O_808,N_24613,N_24805);
nor UO_809 (O_809,N_24603,N_24930);
nand UO_810 (O_810,N_24643,N_24722);
nand UO_811 (O_811,N_24794,N_24475);
and UO_812 (O_812,N_24898,N_24692);
xnor UO_813 (O_813,N_24409,N_24991);
and UO_814 (O_814,N_24463,N_24644);
xnor UO_815 (O_815,N_24915,N_24409);
nand UO_816 (O_816,N_24757,N_24382);
nand UO_817 (O_817,N_24701,N_24536);
xnor UO_818 (O_818,N_24637,N_24735);
and UO_819 (O_819,N_24943,N_24762);
xor UO_820 (O_820,N_24543,N_24912);
nor UO_821 (O_821,N_24969,N_24481);
nand UO_822 (O_822,N_24890,N_24898);
and UO_823 (O_823,N_24584,N_24631);
or UO_824 (O_824,N_24776,N_24640);
nor UO_825 (O_825,N_24652,N_24663);
and UO_826 (O_826,N_24622,N_24634);
nand UO_827 (O_827,N_24377,N_24717);
and UO_828 (O_828,N_24863,N_24624);
or UO_829 (O_829,N_24688,N_24631);
or UO_830 (O_830,N_24562,N_24937);
nand UO_831 (O_831,N_24527,N_24862);
xor UO_832 (O_832,N_24836,N_24543);
nand UO_833 (O_833,N_24487,N_24437);
nor UO_834 (O_834,N_24924,N_24661);
xnor UO_835 (O_835,N_24606,N_24975);
xor UO_836 (O_836,N_24838,N_24563);
xnor UO_837 (O_837,N_24397,N_24673);
nor UO_838 (O_838,N_24674,N_24450);
or UO_839 (O_839,N_24497,N_24503);
nand UO_840 (O_840,N_24645,N_24834);
nor UO_841 (O_841,N_24527,N_24502);
xnor UO_842 (O_842,N_24687,N_24473);
or UO_843 (O_843,N_24800,N_24718);
nand UO_844 (O_844,N_24518,N_24461);
xnor UO_845 (O_845,N_24627,N_24443);
nor UO_846 (O_846,N_24904,N_24881);
or UO_847 (O_847,N_24755,N_24417);
xnor UO_848 (O_848,N_24633,N_24520);
nand UO_849 (O_849,N_24798,N_24609);
nand UO_850 (O_850,N_24408,N_24942);
xnor UO_851 (O_851,N_24557,N_24946);
nand UO_852 (O_852,N_24809,N_24686);
nand UO_853 (O_853,N_24497,N_24392);
and UO_854 (O_854,N_24926,N_24707);
nor UO_855 (O_855,N_24698,N_24869);
or UO_856 (O_856,N_24705,N_24974);
or UO_857 (O_857,N_24766,N_24668);
xnor UO_858 (O_858,N_24725,N_24405);
nand UO_859 (O_859,N_24681,N_24782);
xnor UO_860 (O_860,N_24676,N_24675);
nand UO_861 (O_861,N_24609,N_24578);
or UO_862 (O_862,N_24651,N_24994);
or UO_863 (O_863,N_24883,N_24503);
or UO_864 (O_864,N_24803,N_24982);
nand UO_865 (O_865,N_24862,N_24904);
nand UO_866 (O_866,N_24802,N_24445);
and UO_867 (O_867,N_24829,N_24897);
or UO_868 (O_868,N_24756,N_24712);
nor UO_869 (O_869,N_24579,N_24445);
nor UO_870 (O_870,N_24538,N_24854);
nor UO_871 (O_871,N_24781,N_24996);
nand UO_872 (O_872,N_24884,N_24839);
and UO_873 (O_873,N_24847,N_24785);
and UO_874 (O_874,N_24568,N_24711);
xnor UO_875 (O_875,N_24673,N_24899);
nand UO_876 (O_876,N_24445,N_24757);
xnor UO_877 (O_877,N_24439,N_24905);
xnor UO_878 (O_878,N_24804,N_24897);
xnor UO_879 (O_879,N_24592,N_24441);
or UO_880 (O_880,N_24660,N_24892);
xnor UO_881 (O_881,N_24385,N_24946);
nor UO_882 (O_882,N_24898,N_24878);
or UO_883 (O_883,N_24671,N_24404);
nor UO_884 (O_884,N_24482,N_24958);
or UO_885 (O_885,N_24758,N_24548);
or UO_886 (O_886,N_24494,N_24606);
xor UO_887 (O_887,N_24638,N_24633);
xnor UO_888 (O_888,N_24521,N_24724);
or UO_889 (O_889,N_24405,N_24587);
xor UO_890 (O_890,N_24447,N_24891);
nand UO_891 (O_891,N_24614,N_24617);
and UO_892 (O_892,N_24688,N_24713);
nand UO_893 (O_893,N_24976,N_24921);
nand UO_894 (O_894,N_24904,N_24941);
and UO_895 (O_895,N_24534,N_24898);
and UO_896 (O_896,N_24697,N_24404);
nor UO_897 (O_897,N_24870,N_24768);
nand UO_898 (O_898,N_24833,N_24476);
nand UO_899 (O_899,N_24899,N_24497);
nor UO_900 (O_900,N_24393,N_24865);
nor UO_901 (O_901,N_24770,N_24704);
xor UO_902 (O_902,N_24694,N_24643);
nand UO_903 (O_903,N_24563,N_24659);
and UO_904 (O_904,N_24476,N_24519);
nand UO_905 (O_905,N_24793,N_24471);
nand UO_906 (O_906,N_24446,N_24663);
or UO_907 (O_907,N_24584,N_24697);
or UO_908 (O_908,N_24525,N_24914);
nor UO_909 (O_909,N_24645,N_24866);
xor UO_910 (O_910,N_24805,N_24518);
or UO_911 (O_911,N_24748,N_24502);
and UO_912 (O_912,N_24706,N_24820);
and UO_913 (O_913,N_24815,N_24763);
and UO_914 (O_914,N_24887,N_24641);
nor UO_915 (O_915,N_24572,N_24963);
nand UO_916 (O_916,N_24794,N_24910);
xnor UO_917 (O_917,N_24581,N_24901);
nand UO_918 (O_918,N_24415,N_24617);
or UO_919 (O_919,N_24921,N_24870);
nor UO_920 (O_920,N_24912,N_24785);
xnor UO_921 (O_921,N_24812,N_24808);
nand UO_922 (O_922,N_24394,N_24736);
and UO_923 (O_923,N_24795,N_24872);
nand UO_924 (O_924,N_24460,N_24701);
xor UO_925 (O_925,N_24645,N_24558);
and UO_926 (O_926,N_24717,N_24533);
or UO_927 (O_927,N_24764,N_24910);
nor UO_928 (O_928,N_24613,N_24596);
or UO_929 (O_929,N_24700,N_24828);
xor UO_930 (O_930,N_24450,N_24558);
nand UO_931 (O_931,N_24638,N_24409);
xor UO_932 (O_932,N_24705,N_24774);
or UO_933 (O_933,N_24803,N_24747);
xnor UO_934 (O_934,N_24732,N_24778);
and UO_935 (O_935,N_24880,N_24811);
xor UO_936 (O_936,N_24801,N_24569);
nor UO_937 (O_937,N_24818,N_24458);
or UO_938 (O_938,N_24641,N_24416);
nand UO_939 (O_939,N_24631,N_24831);
nor UO_940 (O_940,N_24401,N_24448);
or UO_941 (O_941,N_24577,N_24862);
nand UO_942 (O_942,N_24629,N_24755);
or UO_943 (O_943,N_24453,N_24828);
xor UO_944 (O_944,N_24709,N_24520);
xnor UO_945 (O_945,N_24654,N_24785);
xor UO_946 (O_946,N_24703,N_24648);
and UO_947 (O_947,N_24925,N_24905);
xor UO_948 (O_948,N_24790,N_24833);
or UO_949 (O_949,N_24723,N_24803);
nand UO_950 (O_950,N_24502,N_24704);
or UO_951 (O_951,N_24630,N_24499);
and UO_952 (O_952,N_24674,N_24765);
nand UO_953 (O_953,N_24473,N_24642);
xnor UO_954 (O_954,N_24948,N_24421);
or UO_955 (O_955,N_24864,N_24388);
and UO_956 (O_956,N_24623,N_24868);
or UO_957 (O_957,N_24991,N_24754);
nand UO_958 (O_958,N_24967,N_24900);
xnor UO_959 (O_959,N_24892,N_24961);
nor UO_960 (O_960,N_24621,N_24746);
or UO_961 (O_961,N_24711,N_24950);
or UO_962 (O_962,N_24847,N_24838);
nor UO_963 (O_963,N_24585,N_24770);
nor UO_964 (O_964,N_24503,N_24695);
xor UO_965 (O_965,N_24584,N_24901);
or UO_966 (O_966,N_24744,N_24830);
or UO_967 (O_967,N_24695,N_24689);
nor UO_968 (O_968,N_24411,N_24776);
xor UO_969 (O_969,N_24758,N_24723);
nand UO_970 (O_970,N_24955,N_24769);
nand UO_971 (O_971,N_24878,N_24409);
nand UO_972 (O_972,N_24653,N_24769);
or UO_973 (O_973,N_24477,N_24873);
and UO_974 (O_974,N_24857,N_24385);
nand UO_975 (O_975,N_24912,N_24743);
or UO_976 (O_976,N_24657,N_24508);
or UO_977 (O_977,N_24918,N_24920);
or UO_978 (O_978,N_24420,N_24386);
xor UO_979 (O_979,N_24853,N_24695);
xnor UO_980 (O_980,N_24740,N_24918);
nand UO_981 (O_981,N_24735,N_24528);
or UO_982 (O_982,N_24935,N_24499);
or UO_983 (O_983,N_24761,N_24634);
xor UO_984 (O_984,N_24982,N_24765);
xor UO_985 (O_985,N_24416,N_24411);
and UO_986 (O_986,N_24427,N_24974);
or UO_987 (O_987,N_24533,N_24569);
nand UO_988 (O_988,N_24548,N_24908);
and UO_989 (O_989,N_24945,N_24931);
xor UO_990 (O_990,N_24768,N_24990);
nand UO_991 (O_991,N_24618,N_24825);
nor UO_992 (O_992,N_24705,N_24647);
or UO_993 (O_993,N_24867,N_24909);
nor UO_994 (O_994,N_24558,N_24910);
nand UO_995 (O_995,N_24906,N_24692);
nor UO_996 (O_996,N_24607,N_24742);
or UO_997 (O_997,N_24448,N_24392);
or UO_998 (O_998,N_24660,N_24380);
nand UO_999 (O_999,N_24518,N_24410);
nand UO_1000 (O_1000,N_24804,N_24816);
or UO_1001 (O_1001,N_24400,N_24706);
nand UO_1002 (O_1002,N_24638,N_24522);
nand UO_1003 (O_1003,N_24470,N_24512);
nor UO_1004 (O_1004,N_24816,N_24487);
xor UO_1005 (O_1005,N_24481,N_24923);
nand UO_1006 (O_1006,N_24902,N_24492);
nand UO_1007 (O_1007,N_24700,N_24917);
xor UO_1008 (O_1008,N_24463,N_24861);
nand UO_1009 (O_1009,N_24969,N_24977);
or UO_1010 (O_1010,N_24570,N_24411);
nor UO_1011 (O_1011,N_24689,N_24829);
or UO_1012 (O_1012,N_24805,N_24519);
nand UO_1013 (O_1013,N_24772,N_24841);
and UO_1014 (O_1014,N_24494,N_24402);
nor UO_1015 (O_1015,N_24582,N_24599);
xor UO_1016 (O_1016,N_24405,N_24421);
xor UO_1017 (O_1017,N_24931,N_24968);
xnor UO_1018 (O_1018,N_24825,N_24454);
and UO_1019 (O_1019,N_24633,N_24593);
or UO_1020 (O_1020,N_24957,N_24946);
nand UO_1021 (O_1021,N_24437,N_24847);
nand UO_1022 (O_1022,N_24670,N_24505);
and UO_1023 (O_1023,N_24849,N_24978);
nor UO_1024 (O_1024,N_24715,N_24995);
and UO_1025 (O_1025,N_24956,N_24802);
or UO_1026 (O_1026,N_24781,N_24864);
nor UO_1027 (O_1027,N_24454,N_24647);
xnor UO_1028 (O_1028,N_24602,N_24984);
xnor UO_1029 (O_1029,N_24535,N_24873);
nor UO_1030 (O_1030,N_24949,N_24982);
xor UO_1031 (O_1031,N_24678,N_24730);
and UO_1032 (O_1032,N_24607,N_24824);
nand UO_1033 (O_1033,N_24889,N_24997);
xnor UO_1034 (O_1034,N_24522,N_24902);
or UO_1035 (O_1035,N_24605,N_24445);
nand UO_1036 (O_1036,N_24579,N_24591);
nand UO_1037 (O_1037,N_24580,N_24516);
nand UO_1038 (O_1038,N_24656,N_24812);
nor UO_1039 (O_1039,N_24510,N_24648);
xnor UO_1040 (O_1040,N_24494,N_24375);
nand UO_1041 (O_1041,N_24499,N_24857);
xnor UO_1042 (O_1042,N_24616,N_24398);
xor UO_1043 (O_1043,N_24869,N_24930);
or UO_1044 (O_1044,N_24518,N_24567);
xor UO_1045 (O_1045,N_24520,N_24638);
xor UO_1046 (O_1046,N_24988,N_24822);
xnor UO_1047 (O_1047,N_24643,N_24930);
nor UO_1048 (O_1048,N_24670,N_24677);
or UO_1049 (O_1049,N_24735,N_24802);
or UO_1050 (O_1050,N_24683,N_24947);
or UO_1051 (O_1051,N_24631,N_24470);
and UO_1052 (O_1052,N_24512,N_24649);
xnor UO_1053 (O_1053,N_24446,N_24812);
nor UO_1054 (O_1054,N_24506,N_24834);
nor UO_1055 (O_1055,N_24782,N_24995);
nor UO_1056 (O_1056,N_24406,N_24982);
or UO_1057 (O_1057,N_24630,N_24770);
and UO_1058 (O_1058,N_24501,N_24483);
or UO_1059 (O_1059,N_24667,N_24808);
xnor UO_1060 (O_1060,N_24482,N_24864);
nor UO_1061 (O_1061,N_24471,N_24715);
and UO_1062 (O_1062,N_24749,N_24666);
and UO_1063 (O_1063,N_24524,N_24509);
nand UO_1064 (O_1064,N_24599,N_24555);
nor UO_1065 (O_1065,N_24941,N_24640);
nand UO_1066 (O_1066,N_24920,N_24872);
and UO_1067 (O_1067,N_24891,N_24621);
or UO_1068 (O_1068,N_24878,N_24866);
or UO_1069 (O_1069,N_24477,N_24604);
and UO_1070 (O_1070,N_24714,N_24832);
or UO_1071 (O_1071,N_24592,N_24932);
xnor UO_1072 (O_1072,N_24625,N_24506);
or UO_1073 (O_1073,N_24853,N_24443);
and UO_1074 (O_1074,N_24980,N_24821);
nor UO_1075 (O_1075,N_24924,N_24591);
or UO_1076 (O_1076,N_24700,N_24447);
nor UO_1077 (O_1077,N_24871,N_24689);
xor UO_1078 (O_1078,N_24693,N_24565);
or UO_1079 (O_1079,N_24765,N_24958);
or UO_1080 (O_1080,N_24969,N_24947);
or UO_1081 (O_1081,N_24470,N_24903);
nor UO_1082 (O_1082,N_24378,N_24742);
xnor UO_1083 (O_1083,N_24569,N_24789);
nor UO_1084 (O_1084,N_24394,N_24619);
nor UO_1085 (O_1085,N_24376,N_24731);
nor UO_1086 (O_1086,N_24862,N_24615);
nor UO_1087 (O_1087,N_24996,N_24682);
xor UO_1088 (O_1088,N_24864,N_24565);
and UO_1089 (O_1089,N_24611,N_24899);
and UO_1090 (O_1090,N_24585,N_24488);
or UO_1091 (O_1091,N_24906,N_24851);
or UO_1092 (O_1092,N_24820,N_24481);
nor UO_1093 (O_1093,N_24832,N_24594);
and UO_1094 (O_1094,N_24557,N_24602);
nor UO_1095 (O_1095,N_24508,N_24558);
and UO_1096 (O_1096,N_24717,N_24813);
xnor UO_1097 (O_1097,N_24454,N_24545);
or UO_1098 (O_1098,N_24710,N_24540);
and UO_1099 (O_1099,N_24505,N_24652);
xor UO_1100 (O_1100,N_24724,N_24538);
nand UO_1101 (O_1101,N_24716,N_24588);
nor UO_1102 (O_1102,N_24873,N_24863);
nor UO_1103 (O_1103,N_24636,N_24703);
and UO_1104 (O_1104,N_24943,N_24917);
xnor UO_1105 (O_1105,N_24848,N_24895);
xor UO_1106 (O_1106,N_24489,N_24859);
xor UO_1107 (O_1107,N_24688,N_24740);
nand UO_1108 (O_1108,N_24785,N_24888);
nand UO_1109 (O_1109,N_24754,N_24718);
nor UO_1110 (O_1110,N_24666,N_24771);
nor UO_1111 (O_1111,N_24929,N_24801);
nand UO_1112 (O_1112,N_24702,N_24383);
nor UO_1113 (O_1113,N_24954,N_24787);
xnor UO_1114 (O_1114,N_24471,N_24492);
and UO_1115 (O_1115,N_24563,N_24539);
and UO_1116 (O_1116,N_24664,N_24597);
or UO_1117 (O_1117,N_24880,N_24667);
and UO_1118 (O_1118,N_24500,N_24934);
or UO_1119 (O_1119,N_24868,N_24767);
or UO_1120 (O_1120,N_24928,N_24979);
and UO_1121 (O_1121,N_24429,N_24878);
xor UO_1122 (O_1122,N_24606,N_24827);
xnor UO_1123 (O_1123,N_24808,N_24394);
xnor UO_1124 (O_1124,N_24929,N_24743);
xor UO_1125 (O_1125,N_24484,N_24565);
or UO_1126 (O_1126,N_24941,N_24774);
xor UO_1127 (O_1127,N_24976,N_24742);
nor UO_1128 (O_1128,N_24958,N_24941);
or UO_1129 (O_1129,N_24502,N_24912);
xnor UO_1130 (O_1130,N_24402,N_24481);
and UO_1131 (O_1131,N_24406,N_24748);
or UO_1132 (O_1132,N_24595,N_24912);
nor UO_1133 (O_1133,N_24759,N_24811);
and UO_1134 (O_1134,N_24740,N_24449);
and UO_1135 (O_1135,N_24819,N_24975);
and UO_1136 (O_1136,N_24669,N_24962);
or UO_1137 (O_1137,N_24902,N_24892);
or UO_1138 (O_1138,N_24380,N_24375);
nor UO_1139 (O_1139,N_24985,N_24424);
xnor UO_1140 (O_1140,N_24391,N_24639);
nor UO_1141 (O_1141,N_24455,N_24445);
xor UO_1142 (O_1142,N_24829,N_24445);
nand UO_1143 (O_1143,N_24740,N_24887);
and UO_1144 (O_1144,N_24931,N_24971);
or UO_1145 (O_1145,N_24419,N_24903);
xor UO_1146 (O_1146,N_24795,N_24716);
xor UO_1147 (O_1147,N_24633,N_24858);
and UO_1148 (O_1148,N_24626,N_24697);
nand UO_1149 (O_1149,N_24828,N_24631);
or UO_1150 (O_1150,N_24834,N_24580);
or UO_1151 (O_1151,N_24599,N_24626);
nor UO_1152 (O_1152,N_24657,N_24618);
and UO_1153 (O_1153,N_24465,N_24668);
and UO_1154 (O_1154,N_24680,N_24543);
nor UO_1155 (O_1155,N_24836,N_24644);
nand UO_1156 (O_1156,N_24852,N_24885);
and UO_1157 (O_1157,N_24932,N_24638);
or UO_1158 (O_1158,N_24863,N_24902);
and UO_1159 (O_1159,N_24770,N_24754);
and UO_1160 (O_1160,N_24407,N_24389);
and UO_1161 (O_1161,N_24658,N_24842);
or UO_1162 (O_1162,N_24491,N_24860);
and UO_1163 (O_1163,N_24435,N_24506);
and UO_1164 (O_1164,N_24466,N_24675);
xor UO_1165 (O_1165,N_24554,N_24727);
and UO_1166 (O_1166,N_24851,N_24831);
and UO_1167 (O_1167,N_24831,N_24916);
and UO_1168 (O_1168,N_24877,N_24694);
xor UO_1169 (O_1169,N_24804,N_24738);
nor UO_1170 (O_1170,N_24977,N_24652);
xor UO_1171 (O_1171,N_24855,N_24562);
or UO_1172 (O_1172,N_24772,N_24509);
nor UO_1173 (O_1173,N_24987,N_24420);
nor UO_1174 (O_1174,N_24735,N_24798);
xnor UO_1175 (O_1175,N_24875,N_24942);
xnor UO_1176 (O_1176,N_24796,N_24612);
nand UO_1177 (O_1177,N_24530,N_24944);
and UO_1178 (O_1178,N_24945,N_24876);
or UO_1179 (O_1179,N_24939,N_24562);
nand UO_1180 (O_1180,N_24608,N_24425);
nor UO_1181 (O_1181,N_24632,N_24637);
or UO_1182 (O_1182,N_24959,N_24907);
or UO_1183 (O_1183,N_24594,N_24745);
nand UO_1184 (O_1184,N_24794,N_24509);
nor UO_1185 (O_1185,N_24538,N_24973);
nand UO_1186 (O_1186,N_24564,N_24908);
and UO_1187 (O_1187,N_24401,N_24375);
and UO_1188 (O_1188,N_24627,N_24610);
or UO_1189 (O_1189,N_24809,N_24636);
xor UO_1190 (O_1190,N_24969,N_24574);
and UO_1191 (O_1191,N_24989,N_24887);
nor UO_1192 (O_1192,N_24935,N_24839);
nand UO_1193 (O_1193,N_24434,N_24420);
or UO_1194 (O_1194,N_24864,N_24926);
xnor UO_1195 (O_1195,N_24418,N_24999);
xnor UO_1196 (O_1196,N_24722,N_24424);
and UO_1197 (O_1197,N_24813,N_24827);
nand UO_1198 (O_1198,N_24796,N_24787);
nand UO_1199 (O_1199,N_24682,N_24773);
nand UO_1200 (O_1200,N_24735,N_24853);
xor UO_1201 (O_1201,N_24714,N_24456);
and UO_1202 (O_1202,N_24723,N_24630);
and UO_1203 (O_1203,N_24528,N_24494);
and UO_1204 (O_1204,N_24856,N_24611);
or UO_1205 (O_1205,N_24511,N_24395);
and UO_1206 (O_1206,N_24721,N_24825);
and UO_1207 (O_1207,N_24820,N_24522);
xor UO_1208 (O_1208,N_24627,N_24777);
nor UO_1209 (O_1209,N_24906,N_24460);
xor UO_1210 (O_1210,N_24568,N_24816);
or UO_1211 (O_1211,N_24555,N_24518);
xnor UO_1212 (O_1212,N_24940,N_24839);
and UO_1213 (O_1213,N_24563,N_24953);
nor UO_1214 (O_1214,N_24547,N_24394);
nor UO_1215 (O_1215,N_24941,N_24852);
and UO_1216 (O_1216,N_24957,N_24876);
nor UO_1217 (O_1217,N_24907,N_24801);
nor UO_1218 (O_1218,N_24462,N_24444);
nand UO_1219 (O_1219,N_24754,N_24916);
or UO_1220 (O_1220,N_24376,N_24923);
and UO_1221 (O_1221,N_24749,N_24639);
nand UO_1222 (O_1222,N_24911,N_24664);
xor UO_1223 (O_1223,N_24833,N_24467);
xor UO_1224 (O_1224,N_24543,N_24638);
xnor UO_1225 (O_1225,N_24401,N_24868);
xor UO_1226 (O_1226,N_24376,N_24484);
or UO_1227 (O_1227,N_24780,N_24941);
or UO_1228 (O_1228,N_24428,N_24957);
or UO_1229 (O_1229,N_24518,N_24897);
nand UO_1230 (O_1230,N_24579,N_24638);
nand UO_1231 (O_1231,N_24890,N_24955);
nand UO_1232 (O_1232,N_24709,N_24444);
xor UO_1233 (O_1233,N_24795,N_24626);
nor UO_1234 (O_1234,N_24849,N_24729);
nor UO_1235 (O_1235,N_24546,N_24676);
nor UO_1236 (O_1236,N_24875,N_24845);
nand UO_1237 (O_1237,N_24569,N_24490);
nor UO_1238 (O_1238,N_24640,N_24901);
nor UO_1239 (O_1239,N_24848,N_24981);
nand UO_1240 (O_1240,N_24844,N_24569);
and UO_1241 (O_1241,N_24382,N_24396);
xnor UO_1242 (O_1242,N_24625,N_24848);
nor UO_1243 (O_1243,N_24587,N_24499);
and UO_1244 (O_1244,N_24919,N_24770);
or UO_1245 (O_1245,N_24607,N_24957);
nor UO_1246 (O_1246,N_24691,N_24563);
or UO_1247 (O_1247,N_24818,N_24990);
nand UO_1248 (O_1248,N_24510,N_24650);
nor UO_1249 (O_1249,N_24837,N_24734);
nand UO_1250 (O_1250,N_24592,N_24992);
and UO_1251 (O_1251,N_24400,N_24666);
nor UO_1252 (O_1252,N_24792,N_24455);
nor UO_1253 (O_1253,N_24787,N_24672);
or UO_1254 (O_1254,N_24669,N_24752);
xnor UO_1255 (O_1255,N_24375,N_24551);
or UO_1256 (O_1256,N_24712,N_24832);
nand UO_1257 (O_1257,N_24533,N_24628);
or UO_1258 (O_1258,N_24529,N_24708);
and UO_1259 (O_1259,N_24524,N_24988);
xor UO_1260 (O_1260,N_24992,N_24499);
nor UO_1261 (O_1261,N_24617,N_24462);
nor UO_1262 (O_1262,N_24592,N_24482);
and UO_1263 (O_1263,N_24625,N_24388);
nor UO_1264 (O_1264,N_24750,N_24459);
nor UO_1265 (O_1265,N_24969,N_24585);
xnor UO_1266 (O_1266,N_24964,N_24945);
nor UO_1267 (O_1267,N_24887,N_24555);
nor UO_1268 (O_1268,N_24480,N_24607);
xor UO_1269 (O_1269,N_24821,N_24528);
or UO_1270 (O_1270,N_24474,N_24678);
and UO_1271 (O_1271,N_24472,N_24944);
nand UO_1272 (O_1272,N_24492,N_24517);
or UO_1273 (O_1273,N_24951,N_24634);
and UO_1274 (O_1274,N_24578,N_24961);
or UO_1275 (O_1275,N_24849,N_24718);
and UO_1276 (O_1276,N_24849,N_24621);
nand UO_1277 (O_1277,N_24617,N_24709);
nor UO_1278 (O_1278,N_24736,N_24800);
and UO_1279 (O_1279,N_24626,N_24800);
xnor UO_1280 (O_1280,N_24827,N_24584);
or UO_1281 (O_1281,N_24415,N_24684);
nor UO_1282 (O_1282,N_24773,N_24399);
xor UO_1283 (O_1283,N_24968,N_24844);
nand UO_1284 (O_1284,N_24566,N_24710);
nand UO_1285 (O_1285,N_24967,N_24435);
and UO_1286 (O_1286,N_24659,N_24575);
or UO_1287 (O_1287,N_24952,N_24640);
nand UO_1288 (O_1288,N_24891,N_24480);
and UO_1289 (O_1289,N_24694,N_24764);
nor UO_1290 (O_1290,N_24951,N_24763);
and UO_1291 (O_1291,N_24532,N_24405);
nand UO_1292 (O_1292,N_24895,N_24809);
or UO_1293 (O_1293,N_24764,N_24408);
or UO_1294 (O_1294,N_24433,N_24678);
or UO_1295 (O_1295,N_24546,N_24673);
nor UO_1296 (O_1296,N_24927,N_24831);
and UO_1297 (O_1297,N_24641,N_24635);
and UO_1298 (O_1298,N_24675,N_24407);
or UO_1299 (O_1299,N_24945,N_24536);
and UO_1300 (O_1300,N_24773,N_24394);
nor UO_1301 (O_1301,N_24608,N_24966);
or UO_1302 (O_1302,N_24928,N_24775);
or UO_1303 (O_1303,N_24541,N_24507);
nand UO_1304 (O_1304,N_24449,N_24662);
nand UO_1305 (O_1305,N_24907,N_24719);
nand UO_1306 (O_1306,N_24884,N_24555);
or UO_1307 (O_1307,N_24563,N_24504);
or UO_1308 (O_1308,N_24948,N_24742);
or UO_1309 (O_1309,N_24417,N_24563);
or UO_1310 (O_1310,N_24508,N_24482);
nor UO_1311 (O_1311,N_24652,N_24863);
and UO_1312 (O_1312,N_24761,N_24455);
nor UO_1313 (O_1313,N_24824,N_24994);
nand UO_1314 (O_1314,N_24653,N_24937);
or UO_1315 (O_1315,N_24451,N_24602);
or UO_1316 (O_1316,N_24459,N_24875);
or UO_1317 (O_1317,N_24758,N_24620);
nand UO_1318 (O_1318,N_24572,N_24823);
or UO_1319 (O_1319,N_24653,N_24409);
nand UO_1320 (O_1320,N_24661,N_24734);
or UO_1321 (O_1321,N_24408,N_24667);
and UO_1322 (O_1322,N_24489,N_24693);
nand UO_1323 (O_1323,N_24791,N_24906);
nand UO_1324 (O_1324,N_24899,N_24388);
nand UO_1325 (O_1325,N_24492,N_24962);
nor UO_1326 (O_1326,N_24507,N_24664);
xor UO_1327 (O_1327,N_24964,N_24543);
nand UO_1328 (O_1328,N_24566,N_24740);
xor UO_1329 (O_1329,N_24979,N_24656);
xnor UO_1330 (O_1330,N_24793,N_24797);
or UO_1331 (O_1331,N_24645,N_24766);
or UO_1332 (O_1332,N_24521,N_24484);
nand UO_1333 (O_1333,N_24448,N_24864);
nor UO_1334 (O_1334,N_24953,N_24577);
xnor UO_1335 (O_1335,N_24855,N_24939);
xor UO_1336 (O_1336,N_24959,N_24455);
xor UO_1337 (O_1337,N_24948,N_24707);
xnor UO_1338 (O_1338,N_24440,N_24404);
nor UO_1339 (O_1339,N_24848,N_24868);
nor UO_1340 (O_1340,N_24562,N_24935);
nand UO_1341 (O_1341,N_24395,N_24866);
nor UO_1342 (O_1342,N_24709,N_24676);
nor UO_1343 (O_1343,N_24694,N_24890);
nor UO_1344 (O_1344,N_24514,N_24565);
xnor UO_1345 (O_1345,N_24811,N_24774);
and UO_1346 (O_1346,N_24438,N_24602);
or UO_1347 (O_1347,N_24600,N_24565);
nor UO_1348 (O_1348,N_24462,N_24896);
nor UO_1349 (O_1349,N_24425,N_24784);
nor UO_1350 (O_1350,N_24741,N_24914);
nand UO_1351 (O_1351,N_24942,N_24756);
nor UO_1352 (O_1352,N_24516,N_24735);
nor UO_1353 (O_1353,N_24512,N_24506);
nor UO_1354 (O_1354,N_24701,N_24416);
nand UO_1355 (O_1355,N_24538,N_24791);
nor UO_1356 (O_1356,N_24699,N_24421);
and UO_1357 (O_1357,N_24531,N_24898);
nor UO_1358 (O_1358,N_24519,N_24697);
nor UO_1359 (O_1359,N_24791,N_24773);
nor UO_1360 (O_1360,N_24644,N_24417);
nand UO_1361 (O_1361,N_24582,N_24851);
and UO_1362 (O_1362,N_24696,N_24595);
nand UO_1363 (O_1363,N_24397,N_24441);
and UO_1364 (O_1364,N_24438,N_24816);
and UO_1365 (O_1365,N_24675,N_24714);
xnor UO_1366 (O_1366,N_24931,N_24397);
and UO_1367 (O_1367,N_24455,N_24719);
nor UO_1368 (O_1368,N_24417,N_24997);
nor UO_1369 (O_1369,N_24453,N_24921);
nor UO_1370 (O_1370,N_24517,N_24430);
xnor UO_1371 (O_1371,N_24843,N_24651);
nand UO_1372 (O_1372,N_24782,N_24719);
and UO_1373 (O_1373,N_24985,N_24707);
and UO_1374 (O_1374,N_24662,N_24515);
or UO_1375 (O_1375,N_24478,N_24570);
xor UO_1376 (O_1376,N_24868,N_24509);
and UO_1377 (O_1377,N_24924,N_24646);
nor UO_1378 (O_1378,N_24676,N_24573);
xor UO_1379 (O_1379,N_24709,N_24620);
xnor UO_1380 (O_1380,N_24892,N_24763);
nand UO_1381 (O_1381,N_24960,N_24439);
nor UO_1382 (O_1382,N_24537,N_24495);
nand UO_1383 (O_1383,N_24839,N_24988);
and UO_1384 (O_1384,N_24636,N_24845);
nand UO_1385 (O_1385,N_24735,N_24382);
or UO_1386 (O_1386,N_24837,N_24649);
or UO_1387 (O_1387,N_24788,N_24874);
xnor UO_1388 (O_1388,N_24592,N_24928);
nand UO_1389 (O_1389,N_24874,N_24534);
xor UO_1390 (O_1390,N_24669,N_24722);
xor UO_1391 (O_1391,N_24901,N_24735);
nor UO_1392 (O_1392,N_24391,N_24710);
xor UO_1393 (O_1393,N_24804,N_24537);
and UO_1394 (O_1394,N_24762,N_24832);
nor UO_1395 (O_1395,N_24660,N_24922);
and UO_1396 (O_1396,N_24557,N_24636);
and UO_1397 (O_1397,N_24495,N_24985);
and UO_1398 (O_1398,N_24739,N_24996);
nand UO_1399 (O_1399,N_24843,N_24709);
or UO_1400 (O_1400,N_24503,N_24432);
and UO_1401 (O_1401,N_24904,N_24793);
nor UO_1402 (O_1402,N_24635,N_24562);
nor UO_1403 (O_1403,N_24740,N_24467);
or UO_1404 (O_1404,N_24547,N_24695);
xor UO_1405 (O_1405,N_24503,N_24408);
xnor UO_1406 (O_1406,N_24960,N_24932);
and UO_1407 (O_1407,N_24689,N_24751);
xor UO_1408 (O_1408,N_24971,N_24853);
nor UO_1409 (O_1409,N_24718,N_24866);
or UO_1410 (O_1410,N_24947,N_24858);
or UO_1411 (O_1411,N_24921,N_24756);
nand UO_1412 (O_1412,N_24622,N_24705);
or UO_1413 (O_1413,N_24874,N_24935);
xnor UO_1414 (O_1414,N_24465,N_24795);
or UO_1415 (O_1415,N_24516,N_24625);
or UO_1416 (O_1416,N_24560,N_24659);
xnor UO_1417 (O_1417,N_24832,N_24554);
nor UO_1418 (O_1418,N_24528,N_24811);
or UO_1419 (O_1419,N_24967,N_24661);
and UO_1420 (O_1420,N_24679,N_24399);
nand UO_1421 (O_1421,N_24774,N_24385);
nand UO_1422 (O_1422,N_24828,N_24472);
nor UO_1423 (O_1423,N_24973,N_24474);
nand UO_1424 (O_1424,N_24807,N_24536);
xor UO_1425 (O_1425,N_24629,N_24715);
xnor UO_1426 (O_1426,N_24785,N_24403);
or UO_1427 (O_1427,N_24450,N_24936);
or UO_1428 (O_1428,N_24532,N_24809);
nand UO_1429 (O_1429,N_24961,N_24941);
or UO_1430 (O_1430,N_24382,N_24662);
nor UO_1431 (O_1431,N_24463,N_24787);
or UO_1432 (O_1432,N_24862,N_24572);
nor UO_1433 (O_1433,N_24613,N_24917);
xnor UO_1434 (O_1434,N_24467,N_24411);
xnor UO_1435 (O_1435,N_24608,N_24578);
nand UO_1436 (O_1436,N_24632,N_24888);
nand UO_1437 (O_1437,N_24631,N_24583);
nand UO_1438 (O_1438,N_24825,N_24915);
xnor UO_1439 (O_1439,N_24986,N_24405);
or UO_1440 (O_1440,N_24522,N_24443);
xnor UO_1441 (O_1441,N_24589,N_24827);
or UO_1442 (O_1442,N_24698,N_24592);
nor UO_1443 (O_1443,N_24805,N_24913);
or UO_1444 (O_1444,N_24568,N_24893);
nand UO_1445 (O_1445,N_24617,N_24816);
or UO_1446 (O_1446,N_24719,N_24918);
and UO_1447 (O_1447,N_24845,N_24941);
nor UO_1448 (O_1448,N_24989,N_24792);
and UO_1449 (O_1449,N_24807,N_24892);
and UO_1450 (O_1450,N_24924,N_24587);
nor UO_1451 (O_1451,N_24995,N_24569);
and UO_1452 (O_1452,N_24695,N_24683);
nor UO_1453 (O_1453,N_24859,N_24502);
nand UO_1454 (O_1454,N_24381,N_24732);
xor UO_1455 (O_1455,N_24488,N_24550);
or UO_1456 (O_1456,N_24508,N_24519);
nand UO_1457 (O_1457,N_24475,N_24701);
xnor UO_1458 (O_1458,N_24912,N_24493);
or UO_1459 (O_1459,N_24910,N_24923);
nor UO_1460 (O_1460,N_24950,N_24383);
and UO_1461 (O_1461,N_24625,N_24710);
or UO_1462 (O_1462,N_24766,N_24812);
nor UO_1463 (O_1463,N_24905,N_24415);
and UO_1464 (O_1464,N_24819,N_24976);
and UO_1465 (O_1465,N_24685,N_24965);
or UO_1466 (O_1466,N_24502,N_24455);
xnor UO_1467 (O_1467,N_24904,N_24858);
xor UO_1468 (O_1468,N_24888,N_24782);
xor UO_1469 (O_1469,N_24401,N_24404);
xor UO_1470 (O_1470,N_24524,N_24767);
or UO_1471 (O_1471,N_24654,N_24819);
or UO_1472 (O_1472,N_24805,N_24524);
nor UO_1473 (O_1473,N_24973,N_24588);
nor UO_1474 (O_1474,N_24632,N_24960);
nand UO_1475 (O_1475,N_24762,N_24852);
nand UO_1476 (O_1476,N_24969,N_24763);
or UO_1477 (O_1477,N_24560,N_24825);
xor UO_1478 (O_1478,N_24884,N_24493);
xnor UO_1479 (O_1479,N_24861,N_24512);
xnor UO_1480 (O_1480,N_24991,N_24796);
or UO_1481 (O_1481,N_24424,N_24504);
or UO_1482 (O_1482,N_24617,N_24814);
and UO_1483 (O_1483,N_24718,N_24801);
or UO_1484 (O_1484,N_24928,N_24401);
xnor UO_1485 (O_1485,N_24617,N_24688);
xor UO_1486 (O_1486,N_24429,N_24458);
xnor UO_1487 (O_1487,N_24993,N_24882);
or UO_1488 (O_1488,N_24888,N_24507);
nor UO_1489 (O_1489,N_24640,N_24804);
or UO_1490 (O_1490,N_24934,N_24548);
nor UO_1491 (O_1491,N_24937,N_24802);
nor UO_1492 (O_1492,N_24939,N_24506);
nor UO_1493 (O_1493,N_24697,N_24786);
or UO_1494 (O_1494,N_24949,N_24810);
nand UO_1495 (O_1495,N_24623,N_24767);
xnor UO_1496 (O_1496,N_24855,N_24974);
and UO_1497 (O_1497,N_24922,N_24668);
nand UO_1498 (O_1498,N_24576,N_24981);
and UO_1499 (O_1499,N_24534,N_24593);
xor UO_1500 (O_1500,N_24605,N_24496);
or UO_1501 (O_1501,N_24689,N_24653);
or UO_1502 (O_1502,N_24749,N_24423);
nor UO_1503 (O_1503,N_24472,N_24595);
xnor UO_1504 (O_1504,N_24551,N_24761);
and UO_1505 (O_1505,N_24613,N_24581);
xor UO_1506 (O_1506,N_24998,N_24708);
nor UO_1507 (O_1507,N_24607,N_24553);
xor UO_1508 (O_1508,N_24903,N_24403);
or UO_1509 (O_1509,N_24796,N_24600);
nand UO_1510 (O_1510,N_24892,N_24395);
nor UO_1511 (O_1511,N_24537,N_24597);
nand UO_1512 (O_1512,N_24473,N_24919);
and UO_1513 (O_1513,N_24845,N_24766);
xnor UO_1514 (O_1514,N_24381,N_24603);
and UO_1515 (O_1515,N_24861,N_24875);
or UO_1516 (O_1516,N_24829,N_24910);
xnor UO_1517 (O_1517,N_24591,N_24722);
or UO_1518 (O_1518,N_24954,N_24808);
and UO_1519 (O_1519,N_24748,N_24462);
or UO_1520 (O_1520,N_24985,N_24979);
nor UO_1521 (O_1521,N_24905,N_24491);
nand UO_1522 (O_1522,N_24910,N_24715);
xor UO_1523 (O_1523,N_24655,N_24978);
or UO_1524 (O_1524,N_24934,N_24999);
xor UO_1525 (O_1525,N_24562,N_24986);
and UO_1526 (O_1526,N_24679,N_24695);
xnor UO_1527 (O_1527,N_24520,N_24675);
xor UO_1528 (O_1528,N_24840,N_24492);
xor UO_1529 (O_1529,N_24417,N_24633);
xnor UO_1530 (O_1530,N_24671,N_24964);
xor UO_1531 (O_1531,N_24378,N_24915);
nand UO_1532 (O_1532,N_24409,N_24752);
nor UO_1533 (O_1533,N_24865,N_24890);
nand UO_1534 (O_1534,N_24818,N_24706);
or UO_1535 (O_1535,N_24771,N_24745);
xnor UO_1536 (O_1536,N_24659,N_24858);
nand UO_1537 (O_1537,N_24989,N_24478);
nor UO_1538 (O_1538,N_24433,N_24913);
nand UO_1539 (O_1539,N_24913,N_24867);
nor UO_1540 (O_1540,N_24664,N_24482);
or UO_1541 (O_1541,N_24555,N_24701);
nand UO_1542 (O_1542,N_24832,N_24895);
xor UO_1543 (O_1543,N_24668,N_24937);
or UO_1544 (O_1544,N_24687,N_24589);
nor UO_1545 (O_1545,N_24796,N_24552);
nor UO_1546 (O_1546,N_24781,N_24641);
nand UO_1547 (O_1547,N_24764,N_24788);
nor UO_1548 (O_1548,N_24644,N_24693);
xnor UO_1549 (O_1549,N_24441,N_24625);
nor UO_1550 (O_1550,N_24425,N_24899);
and UO_1551 (O_1551,N_24427,N_24486);
nor UO_1552 (O_1552,N_24714,N_24510);
and UO_1553 (O_1553,N_24704,N_24961);
xnor UO_1554 (O_1554,N_24839,N_24566);
nand UO_1555 (O_1555,N_24883,N_24824);
nand UO_1556 (O_1556,N_24546,N_24408);
nor UO_1557 (O_1557,N_24495,N_24525);
xnor UO_1558 (O_1558,N_24614,N_24534);
nand UO_1559 (O_1559,N_24944,N_24985);
or UO_1560 (O_1560,N_24575,N_24637);
xor UO_1561 (O_1561,N_24723,N_24767);
nand UO_1562 (O_1562,N_24804,N_24705);
nand UO_1563 (O_1563,N_24570,N_24621);
and UO_1564 (O_1564,N_24488,N_24812);
and UO_1565 (O_1565,N_24575,N_24940);
xnor UO_1566 (O_1566,N_24776,N_24512);
nand UO_1567 (O_1567,N_24979,N_24410);
xor UO_1568 (O_1568,N_24535,N_24500);
or UO_1569 (O_1569,N_24463,N_24772);
or UO_1570 (O_1570,N_24924,N_24487);
xnor UO_1571 (O_1571,N_24916,N_24608);
or UO_1572 (O_1572,N_24856,N_24829);
xor UO_1573 (O_1573,N_24724,N_24861);
nand UO_1574 (O_1574,N_24556,N_24797);
nand UO_1575 (O_1575,N_24831,N_24799);
nand UO_1576 (O_1576,N_24577,N_24729);
nand UO_1577 (O_1577,N_24880,N_24453);
or UO_1578 (O_1578,N_24556,N_24653);
nand UO_1579 (O_1579,N_24407,N_24783);
or UO_1580 (O_1580,N_24730,N_24954);
nor UO_1581 (O_1581,N_24778,N_24748);
or UO_1582 (O_1582,N_24629,N_24444);
xor UO_1583 (O_1583,N_24384,N_24580);
nand UO_1584 (O_1584,N_24400,N_24756);
xor UO_1585 (O_1585,N_24382,N_24441);
xor UO_1586 (O_1586,N_24517,N_24885);
and UO_1587 (O_1587,N_24722,N_24922);
xor UO_1588 (O_1588,N_24885,N_24976);
nor UO_1589 (O_1589,N_24508,N_24925);
nor UO_1590 (O_1590,N_24500,N_24414);
nor UO_1591 (O_1591,N_24967,N_24859);
nor UO_1592 (O_1592,N_24973,N_24631);
nand UO_1593 (O_1593,N_24933,N_24658);
nor UO_1594 (O_1594,N_24807,N_24596);
or UO_1595 (O_1595,N_24889,N_24942);
xor UO_1596 (O_1596,N_24853,N_24835);
or UO_1597 (O_1597,N_24572,N_24420);
nand UO_1598 (O_1598,N_24847,N_24476);
nor UO_1599 (O_1599,N_24580,N_24653);
or UO_1600 (O_1600,N_24690,N_24482);
xor UO_1601 (O_1601,N_24874,N_24937);
and UO_1602 (O_1602,N_24540,N_24783);
nor UO_1603 (O_1603,N_24460,N_24976);
and UO_1604 (O_1604,N_24376,N_24931);
nand UO_1605 (O_1605,N_24962,N_24399);
or UO_1606 (O_1606,N_24596,N_24921);
nand UO_1607 (O_1607,N_24985,N_24745);
and UO_1608 (O_1608,N_24862,N_24832);
nor UO_1609 (O_1609,N_24696,N_24581);
nand UO_1610 (O_1610,N_24642,N_24511);
nor UO_1611 (O_1611,N_24616,N_24765);
and UO_1612 (O_1612,N_24812,N_24422);
or UO_1613 (O_1613,N_24843,N_24859);
and UO_1614 (O_1614,N_24380,N_24722);
xor UO_1615 (O_1615,N_24536,N_24825);
xnor UO_1616 (O_1616,N_24510,N_24527);
xnor UO_1617 (O_1617,N_24590,N_24823);
nor UO_1618 (O_1618,N_24461,N_24539);
xnor UO_1619 (O_1619,N_24993,N_24566);
nor UO_1620 (O_1620,N_24900,N_24949);
or UO_1621 (O_1621,N_24871,N_24856);
nand UO_1622 (O_1622,N_24491,N_24622);
nor UO_1623 (O_1623,N_24497,N_24929);
or UO_1624 (O_1624,N_24560,N_24513);
or UO_1625 (O_1625,N_24642,N_24493);
nor UO_1626 (O_1626,N_24895,N_24875);
nor UO_1627 (O_1627,N_24794,N_24752);
nor UO_1628 (O_1628,N_24865,N_24711);
nor UO_1629 (O_1629,N_24796,N_24825);
or UO_1630 (O_1630,N_24962,N_24592);
xnor UO_1631 (O_1631,N_24886,N_24778);
and UO_1632 (O_1632,N_24541,N_24795);
nand UO_1633 (O_1633,N_24816,N_24724);
xnor UO_1634 (O_1634,N_24624,N_24886);
and UO_1635 (O_1635,N_24833,N_24826);
nor UO_1636 (O_1636,N_24656,N_24853);
xor UO_1637 (O_1637,N_24724,N_24614);
and UO_1638 (O_1638,N_24855,N_24823);
and UO_1639 (O_1639,N_24987,N_24849);
or UO_1640 (O_1640,N_24833,N_24452);
xor UO_1641 (O_1641,N_24950,N_24712);
xor UO_1642 (O_1642,N_24623,N_24797);
and UO_1643 (O_1643,N_24573,N_24907);
nand UO_1644 (O_1644,N_24582,N_24498);
or UO_1645 (O_1645,N_24479,N_24436);
and UO_1646 (O_1646,N_24712,N_24569);
or UO_1647 (O_1647,N_24752,N_24509);
nand UO_1648 (O_1648,N_24953,N_24442);
xor UO_1649 (O_1649,N_24484,N_24921);
xor UO_1650 (O_1650,N_24901,N_24423);
nor UO_1651 (O_1651,N_24828,N_24737);
nor UO_1652 (O_1652,N_24612,N_24804);
and UO_1653 (O_1653,N_24589,N_24897);
xor UO_1654 (O_1654,N_24873,N_24926);
or UO_1655 (O_1655,N_24695,N_24646);
and UO_1656 (O_1656,N_24961,N_24474);
or UO_1657 (O_1657,N_24975,N_24741);
and UO_1658 (O_1658,N_24498,N_24507);
and UO_1659 (O_1659,N_24873,N_24375);
xor UO_1660 (O_1660,N_24876,N_24602);
nand UO_1661 (O_1661,N_24556,N_24680);
xor UO_1662 (O_1662,N_24403,N_24550);
xnor UO_1663 (O_1663,N_24539,N_24631);
nor UO_1664 (O_1664,N_24491,N_24418);
nand UO_1665 (O_1665,N_24997,N_24485);
nor UO_1666 (O_1666,N_24663,N_24638);
or UO_1667 (O_1667,N_24710,N_24973);
xor UO_1668 (O_1668,N_24657,N_24546);
or UO_1669 (O_1669,N_24503,N_24899);
xnor UO_1670 (O_1670,N_24944,N_24788);
and UO_1671 (O_1671,N_24605,N_24682);
or UO_1672 (O_1672,N_24415,N_24437);
xor UO_1673 (O_1673,N_24837,N_24401);
nor UO_1674 (O_1674,N_24985,N_24751);
nand UO_1675 (O_1675,N_24713,N_24814);
xor UO_1676 (O_1676,N_24748,N_24623);
nor UO_1677 (O_1677,N_24414,N_24626);
nor UO_1678 (O_1678,N_24937,N_24865);
or UO_1679 (O_1679,N_24835,N_24860);
xnor UO_1680 (O_1680,N_24992,N_24963);
nor UO_1681 (O_1681,N_24406,N_24578);
nor UO_1682 (O_1682,N_24559,N_24841);
or UO_1683 (O_1683,N_24578,N_24679);
and UO_1684 (O_1684,N_24677,N_24879);
and UO_1685 (O_1685,N_24856,N_24641);
xnor UO_1686 (O_1686,N_24745,N_24993);
or UO_1687 (O_1687,N_24673,N_24767);
or UO_1688 (O_1688,N_24590,N_24867);
nand UO_1689 (O_1689,N_24428,N_24879);
xnor UO_1690 (O_1690,N_24842,N_24858);
nand UO_1691 (O_1691,N_24801,N_24620);
nand UO_1692 (O_1692,N_24540,N_24733);
nand UO_1693 (O_1693,N_24863,N_24597);
nand UO_1694 (O_1694,N_24586,N_24419);
or UO_1695 (O_1695,N_24986,N_24645);
or UO_1696 (O_1696,N_24952,N_24468);
or UO_1697 (O_1697,N_24757,N_24858);
or UO_1698 (O_1698,N_24473,N_24689);
nor UO_1699 (O_1699,N_24889,N_24590);
xor UO_1700 (O_1700,N_24677,N_24986);
or UO_1701 (O_1701,N_24763,N_24888);
xnor UO_1702 (O_1702,N_24824,N_24506);
nor UO_1703 (O_1703,N_24692,N_24946);
or UO_1704 (O_1704,N_24476,N_24938);
or UO_1705 (O_1705,N_24606,N_24669);
xor UO_1706 (O_1706,N_24479,N_24785);
or UO_1707 (O_1707,N_24508,N_24946);
xnor UO_1708 (O_1708,N_24529,N_24449);
nor UO_1709 (O_1709,N_24468,N_24835);
or UO_1710 (O_1710,N_24690,N_24524);
xor UO_1711 (O_1711,N_24592,N_24853);
or UO_1712 (O_1712,N_24567,N_24878);
xnor UO_1713 (O_1713,N_24659,N_24705);
nor UO_1714 (O_1714,N_24775,N_24404);
or UO_1715 (O_1715,N_24951,N_24724);
and UO_1716 (O_1716,N_24647,N_24481);
or UO_1717 (O_1717,N_24573,N_24523);
and UO_1718 (O_1718,N_24848,N_24722);
nand UO_1719 (O_1719,N_24385,N_24551);
nand UO_1720 (O_1720,N_24517,N_24499);
or UO_1721 (O_1721,N_24601,N_24894);
nor UO_1722 (O_1722,N_24767,N_24496);
nand UO_1723 (O_1723,N_24773,N_24459);
nand UO_1724 (O_1724,N_24746,N_24826);
or UO_1725 (O_1725,N_24530,N_24688);
nand UO_1726 (O_1726,N_24821,N_24832);
nor UO_1727 (O_1727,N_24459,N_24849);
and UO_1728 (O_1728,N_24711,N_24910);
or UO_1729 (O_1729,N_24756,N_24727);
or UO_1730 (O_1730,N_24740,N_24679);
nor UO_1731 (O_1731,N_24453,N_24783);
or UO_1732 (O_1732,N_24408,N_24700);
and UO_1733 (O_1733,N_24974,N_24646);
and UO_1734 (O_1734,N_24408,N_24540);
nor UO_1735 (O_1735,N_24973,N_24404);
nor UO_1736 (O_1736,N_24727,N_24861);
nand UO_1737 (O_1737,N_24735,N_24383);
xnor UO_1738 (O_1738,N_24744,N_24533);
xnor UO_1739 (O_1739,N_24875,N_24617);
or UO_1740 (O_1740,N_24798,N_24903);
nand UO_1741 (O_1741,N_24928,N_24584);
or UO_1742 (O_1742,N_24993,N_24897);
or UO_1743 (O_1743,N_24990,N_24443);
or UO_1744 (O_1744,N_24681,N_24439);
or UO_1745 (O_1745,N_24595,N_24970);
and UO_1746 (O_1746,N_24554,N_24697);
and UO_1747 (O_1747,N_24726,N_24408);
nand UO_1748 (O_1748,N_24879,N_24776);
nor UO_1749 (O_1749,N_24654,N_24646);
xnor UO_1750 (O_1750,N_24663,N_24621);
xnor UO_1751 (O_1751,N_24886,N_24432);
nor UO_1752 (O_1752,N_24991,N_24779);
or UO_1753 (O_1753,N_24535,N_24851);
or UO_1754 (O_1754,N_24659,N_24786);
xor UO_1755 (O_1755,N_24410,N_24916);
nor UO_1756 (O_1756,N_24386,N_24959);
and UO_1757 (O_1757,N_24786,N_24876);
nand UO_1758 (O_1758,N_24654,N_24649);
nor UO_1759 (O_1759,N_24547,N_24965);
nor UO_1760 (O_1760,N_24518,N_24466);
and UO_1761 (O_1761,N_24596,N_24562);
xnor UO_1762 (O_1762,N_24638,N_24584);
xor UO_1763 (O_1763,N_24805,N_24627);
and UO_1764 (O_1764,N_24735,N_24645);
or UO_1765 (O_1765,N_24559,N_24697);
and UO_1766 (O_1766,N_24890,N_24567);
nand UO_1767 (O_1767,N_24548,N_24904);
or UO_1768 (O_1768,N_24865,N_24908);
or UO_1769 (O_1769,N_24571,N_24780);
nor UO_1770 (O_1770,N_24873,N_24709);
nand UO_1771 (O_1771,N_24867,N_24885);
xor UO_1772 (O_1772,N_24793,N_24931);
and UO_1773 (O_1773,N_24533,N_24793);
xnor UO_1774 (O_1774,N_24482,N_24543);
or UO_1775 (O_1775,N_24503,N_24520);
xor UO_1776 (O_1776,N_24628,N_24457);
nor UO_1777 (O_1777,N_24618,N_24506);
and UO_1778 (O_1778,N_24929,N_24816);
and UO_1779 (O_1779,N_24390,N_24676);
and UO_1780 (O_1780,N_24551,N_24852);
or UO_1781 (O_1781,N_24945,N_24726);
nor UO_1782 (O_1782,N_24874,N_24852);
or UO_1783 (O_1783,N_24807,N_24473);
nand UO_1784 (O_1784,N_24756,N_24541);
and UO_1785 (O_1785,N_24566,N_24992);
nor UO_1786 (O_1786,N_24523,N_24997);
nor UO_1787 (O_1787,N_24591,N_24863);
nor UO_1788 (O_1788,N_24485,N_24668);
nor UO_1789 (O_1789,N_24602,N_24525);
and UO_1790 (O_1790,N_24413,N_24790);
xor UO_1791 (O_1791,N_24377,N_24731);
nand UO_1792 (O_1792,N_24869,N_24964);
or UO_1793 (O_1793,N_24908,N_24526);
nor UO_1794 (O_1794,N_24987,N_24380);
and UO_1795 (O_1795,N_24887,N_24880);
xnor UO_1796 (O_1796,N_24890,N_24502);
or UO_1797 (O_1797,N_24696,N_24613);
or UO_1798 (O_1798,N_24833,N_24793);
xor UO_1799 (O_1799,N_24648,N_24742);
nor UO_1800 (O_1800,N_24833,N_24617);
xor UO_1801 (O_1801,N_24827,N_24963);
xnor UO_1802 (O_1802,N_24629,N_24805);
or UO_1803 (O_1803,N_24664,N_24525);
or UO_1804 (O_1804,N_24610,N_24631);
nor UO_1805 (O_1805,N_24681,N_24678);
nor UO_1806 (O_1806,N_24979,N_24552);
or UO_1807 (O_1807,N_24771,N_24907);
nor UO_1808 (O_1808,N_24459,N_24918);
xnor UO_1809 (O_1809,N_24511,N_24825);
and UO_1810 (O_1810,N_24581,N_24725);
nor UO_1811 (O_1811,N_24760,N_24380);
nand UO_1812 (O_1812,N_24605,N_24539);
nand UO_1813 (O_1813,N_24640,N_24575);
nor UO_1814 (O_1814,N_24722,N_24727);
nand UO_1815 (O_1815,N_24754,N_24554);
nor UO_1816 (O_1816,N_24886,N_24946);
and UO_1817 (O_1817,N_24376,N_24930);
or UO_1818 (O_1818,N_24390,N_24920);
xnor UO_1819 (O_1819,N_24696,N_24784);
or UO_1820 (O_1820,N_24577,N_24651);
xnor UO_1821 (O_1821,N_24652,N_24848);
nand UO_1822 (O_1822,N_24894,N_24808);
nor UO_1823 (O_1823,N_24823,N_24761);
xnor UO_1824 (O_1824,N_24531,N_24734);
nor UO_1825 (O_1825,N_24485,N_24677);
and UO_1826 (O_1826,N_24991,N_24933);
xor UO_1827 (O_1827,N_24481,N_24728);
xor UO_1828 (O_1828,N_24691,N_24528);
nor UO_1829 (O_1829,N_24711,N_24573);
or UO_1830 (O_1830,N_24792,N_24820);
nand UO_1831 (O_1831,N_24659,N_24719);
and UO_1832 (O_1832,N_24541,N_24515);
xor UO_1833 (O_1833,N_24439,N_24988);
nor UO_1834 (O_1834,N_24582,N_24416);
nor UO_1835 (O_1835,N_24383,N_24960);
nor UO_1836 (O_1836,N_24485,N_24533);
nor UO_1837 (O_1837,N_24660,N_24905);
nor UO_1838 (O_1838,N_24476,N_24751);
nor UO_1839 (O_1839,N_24377,N_24846);
nor UO_1840 (O_1840,N_24772,N_24434);
xnor UO_1841 (O_1841,N_24874,N_24569);
xnor UO_1842 (O_1842,N_24815,N_24765);
nor UO_1843 (O_1843,N_24564,N_24620);
or UO_1844 (O_1844,N_24518,N_24451);
xor UO_1845 (O_1845,N_24668,N_24493);
nor UO_1846 (O_1846,N_24910,N_24996);
and UO_1847 (O_1847,N_24844,N_24436);
xnor UO_1848 (O_1848,N_24437,N_24482);
xnor UO_1849 (O_1849,N_24973,N_24598);
nand UO_1850 (O_1850,N_24778,N_24473);
nand UO_1851 (O_1851,N_24770,N_24817);
xor UO_1852 (O_1852,N_24861,N_24834);
nand UO_1853 (O_1853,N_24558,N_24632);
and UO_1854 (O_1854,N_24941,N_24829);
or UO_1855 (O_1855,N_24602,N_24450);
nand UO_1856 (O_1856,N_24881,N_24687);
nor UO_1857 (O_1857,N_24642,N_24955);
and UO_1858 (O_1858,N_24690,N_24921);
and UO_1859 (O_1859,N_24958,N_24504);
nand UO_1860 (O_1860,N_24844,N_24697);
nor UO_1861 (O_1861,N_24939,N_24800);
nor UO_1862 (O_1862,N_24440,N_24561);
or UO_1863 (O_1863,N_24878,N_24618);
and UO_1864 (O_1864,N_24560,N_24525);
nor UO_1865 (O_1865,N_24977,N_24478);
nor UO_1866 (O_1866,N_24915,N_24400);
nand UO_1867 (O_1867,N_24663,N_24477);
nor UO_1868 (O_1868,N_24698,N_24582);
and UO_1869 (O_1869,N_24690,N_24502);
and UO_1870 (O_1870,N_24659,N_24818);
xor UO_1871 (O_1871,N_24466,N_24573);
and UO_1872 (O_1872,N_24521,N_24443);
and UO_1873 (O_1873,N_24519,N_24954);
nand UO_1874 (O_1874,N_24996,N_24585);
and UO_1875 (O_1875,N_24719,N_24996);
nand UO_1876 (O_1876,N_24459,N_24825);
or UO_1877 (O_1877,N_24890,N_24393);
xor UO_1878 (O_1878,N_24390,N_24706);
nand UO_1879 (O_1879,N_24930,N_24737);
and UO_1880 (O_1880,N_24444,N_24759);
xor UO_1881 (O_1881,N_24505,N_24447);
nand UO_1882 (O_1882,N_24773,N_24464);
nand UO_1883 (O_1883,N_24746,N_24981);
and UO_1884 (O_1884,N_24563,N_24764);
or UO_1885 (O_1885,N_24858,N_24537);
nand UO_1886 (O_1886,N_24495,N_24610);
xor UO_1887 (O_1887,N_24778,N_24895);
and UO_1888 (O_1888,N_24660,N_24794);
nand UO_1889 (O_1889,N_24701,N_24859);
nor UO_1890 (O_1890,N_24878,N_24687);
nor UO_1891 (O_1891,N_24397,N_24968);
and UO_1892 (O_1892,N_24416,N_24735);
xor UO_1893 (O_1893,N_24988,N_24729);
nand UO_1894 (O_1894,N_24508,N_24808);
or UO_1895 (O_1895,N_24780,N_24569);
nand UO_1896 (O_1896,N_24410,N_24971);
nor UO_1897 (O_1897,N_24421,N_24525);
nor UO_1898 (O_1898,N_24687,N_24507);
or UO_1899 (O_1899,N_24675,N_24773);
or UO_1900 (O_1900,N_24677,N_24903);
xnor UO_1901 (O_1901,N_24925,N_24856);
nor UO_1902 (O_1902,N_24961,N_24684);
nor UO_1903 (O_1903,N_24544,N_24807);
and UO_1904 (O_1904,N_24801,N_24594);
or UO_1905 (O_1905,N_24909,N_24552);
xnor UO_1906 (O_1906,N_24879,N_24400);
xnor UO_1907 (O_1907,N_24530,N_24985);
nor UO_1908 (O_1908,N_24646,N_24722);
or UO_1909 (O_1909,N_24514,N_24937);
or UO_1910 (O_1910,N_24670,N_24441);
xor UO_1911 (O_1911,N_24568,N_24719);
and UO_1912 (O_1912,N_24587,N_24603);
nand UO_1913 (O_1913,N_24408,N_24709);
xnor UO_1914 (O_1914,N_24764,N_24735);
and UO_1915 (O_1915,N_24898,N_24495);
nand UO_1916 (O_1916,N_24834,N_24924);
or UO_1917 (O_1917,N_24972,N_24459);
nor UO_1918 (O_1918,N_24998,N_24420);
nand UO_1919 (O_1919,N_24509,N_24578);
and UO_1920 (O_1920,N_24444,N_24708);
or UO_1921 (O_1921,N_24713,N_24930);
or UO_1922 (O_1922,N_24856,N_24435);
nor UO_1923 (O_1923,N_24447,N_24964);
nor UO_1924 (O_1924,N_24395,N_24938);
xnor UO_1925 (O_1925,N_24391,N_24704);
xor UO_1926 (O_1926,N_24925,N_24723);
or UO_1927 (O_1927,N_24392,N_24828);
nand UO_1928 (O_1928,N_24847,N_24793);
nand UO_1929 (O_1929,N_24947,N_24423);
nor UO_1930 (O_1930,N_24680,N_24620);
and UO_1931 (O_1931,N_24812,N_24829);
xor UO_1932 (O_1932,N_24664,N_24583);
or UO_1933 (O_1933,N_24855,N_24947);
xor UO_1934 (O_1934,N_24486,N_24860);
and UO_1935 (O_1935,N_24909,N_24583);
and UO_1936 (O_1936,N_24636,N_24967);
nor UO_1937 (O_1937,N_24491,N_24797);
nand UO_1938 (O_1938,N_24628,N_24668);
and UO_1939 (O_1939,N_24620,N_24440);
or UO_1940 (O_1940,N_24635,N_24544);
and UO_1941 (O_1941,N_24918,N_24565);
or UO_1942 (O_1942,N_24992,N_24826);
and UO_1943 (O_1943,N_24942,N_24530);
nand UO_1944 (O_1944,N_24413,N_24724);
xnor UO_1945 (O_1945,N_24459,N_24760);
nand UO_1946 (O_1946,N_24581,N_24738);
or UO_1947 (O_1947,N_24697,N_24601);
or UO_1948 (O_1948,N_24625,N_24948);
nand UO_1949 (O_1949,N_24723,N_24980);
or UO_1950 (O_1950,N_24743,N_24765);
or UO_1951 (O_1951,N_24456,N_24406);
nor UO_1952 (O_1952,N_24504,N_24719);
or UO_1953 (O_1953,N_24568,N_24543);
xor UO_1954 (O_1954,N_24377,N_24831);
or UO_1955 (O_1955,N_24393,N_24390);
nand UO_1956 (O_1956,N_24701,N_24889);
or UO_1957 (O_1957,N_24404,N_24927);
nor UO_1958 (O_1958,N_24725,N_24701);
and UO_1959 (O_1959,N_24663,N_24844);
or UO_1960 (O_1960,N_24738,N_24396);
xnor UO_1961 (O_1961,N_24663,N_24667);
nor UO_1962 (O_1962,N_24888,N_24951);
nor UO_1963 (O_1963,N_24926,N_24701);
or UO_1964 (O_1964,N_24704,N_24457);
nor UO_1965 (O_1965,N_24785,N_24506);
and UO_1966 (O_1966,N_24575,N_24481);
nand UO_1967 (O_1967,N_24465,N_24979);
and UO_1968 (O_1968,N_24787,N_24519);
or UO_1969 (O_1969,N_24983,N_24843);
or UO_1970 (O_1970,N_24447,N_24727);
or UO_1971 (O_1971,N_24507,N_24908);
nor UO_1972 (O_1972,N_24754,N_24764);
xor UO_1973 (O_1973,N_24965,N_24682);
and UO_1974 (O_1974,N_24407,N_24686);
nor UO_1975 (O_1975,N_24595,N_24674);
xnor UO_1976 (O_1976,N_24679,N_24527);
and UO_1977 (O_1977,N_24877,N_24703);
or UO_1978 (O_1978,N_24926,N_24717);
or UO_1979 (O_1979,N_24762,N_24521);
nand UO_1980 (O_1980,N_24486,N_24830);
or UO_1981 (O_1981,N_24834,N_24380);
nor UO_1982 (O_1982,N_24578,N_24395);
xor UO_1983 (O_1983,N_24425,N_24838);
nor UO_1984 (O_1984,N_24770,N_24480);
or UO_1985 (O_1985,N_24548,N_24889);
and UO_1986 (O_1986,N_24458,N_24426);
nand UO_1987 (O_1987,N_24819,N_24909);
or UO_1988 (O_1988,N_24744,N_24918);
and UO_1989 (O_1989,N_24703,N_24823);
and UO_1990 (O_1990,N_24580,N_24865);
nor UO_1991 (O_1991,N_24933,N_24987);
nand UO_1992 (O_1992,N_24945,N_24745);
nor UO_1993 (O_1993,N_24396,N_24616);
and UO_1994 (O_1994,N_24513,N_24389);
nor UO_1995 (O_1995,N_24661,N_24928);
nor UO_1996 (O_1996,N_24561,N_24451);
or UO_1997 (O_1997,N_24836,N_24551);
xnor UO_1998 (O_1998,N_24510,N_24519);
or UO_1999 (O_1999,N_24836,N_24840);
xor UO_2000 (O_2000,N_24465,N_24701);
xor UO_2001 (O_2001,N_24501,N_24943);
xnor UO_2002 (O_2002,N_24847,N_24986);
nor UO_2003 (O_2003,N_24790,N_24679);
nand UO_2004 (O_2004,N_24971,N_24950);
and UO_2005 (O_2005,N_24436,N_24829);
nor UO_2006 (O_2006,N_24612,N_24948);
nand UO_2007 (O_2007,N_24564,N_24772);
nor UO_2008 (O_2008,N_24721,N_24961);
xnor UO_2009 (O_2009,N_24926,N_24975);
or UO_2010 (O_2010,N_24620,N_24971);
or UO_2011 (O_2011,N_24910,N_24819);
and UO_2012 (O_2012,N_24712,N_24398);
nor UO_2013 (O_2013,N_24709,N_24936);
xor UO_2014 (O_2014,N_24707,N_24977);
nor UO_2015 (O_2015,N_24806,N_24952);
nand UO_2016 (O_2016,N_24588,N_24745);
nand UO_2017 (O_2017,N_24427,N_24610);
nand UO_2018 (O_2018,N_24573,N_24490);
and UO_2019 (O_2019,N_24766,N_24983);
nand UO_2020 (O_2020,N_24868,N_24462);
nand UO_2021 (O_2021,N_24654,N_24632);
or UO_2022 (O_2022,N_24538,N_24420);
nand UO_2023 (O_2023,N_24552,N_24499);
nand UO_2024 (O_2024,N_24633,N_24882);
nand UO_2025 (O_2025,N_24415,N_24962);
nor UO_2026 (O_2026,N_24675,N_24685);
xor UO_2027 (O_2027,N_24611,N_24974);
nand UO_2028 (O_2028,N_24476,N_24443);
or UO_2029 (O_2029,N_24670,N_24579);
nand UO_2030 (O_2030,N_24750,N_24564);
and UO_2031 (O_2031,N_24900,N_24898);
or UO_2032 (O_2032,N_24665,N_24741);
nand UO_2033 (O_2033,N_24897,N_24771);
and UO_2034 (O_2034,N_24486,N_24667);
xor UO_2035 (O_2035,N_24536,N_24757);
xor UO_2036 (O_2036,N_24875,N_24519);
nor UO_2037 (O_2037,N_24827,N_24590);
xnor UO_2038 (O_2038,N_24938,N_24939);
nor UO_2039 (O_2039,N_24754,N_24422);
xor UO_2040 (O_2040,N_24688,N_24471);
nand UO_2041 (O_2041,N_24509,N_24866);
xor UO_2042 (O_2042,N_24419,N_24797);
or UO_2043 (O_2043,N_24784,N_24778);
nor UO_2044 (O_2044,N_24382,N_24645);
xnor UO_2045 (O_2045,N_24491,N_24438);
nand UO_2046 (O_2046,N_24421,N_24583);
nand UO_2047 (O_2047,N_24697,N_24587);
or UO_2048 (O_2048,N_24927,N_24767);
and UO_2049 (O_2049,N_24657,N_24840);
nand UO_2050 (O_2050,N_24538,N_24656);
nand UO_2051 (O_2051,N_24860,N_24984);
nand UO_2052 (O_2052,N_24770,N_24872);
nor UO_2053 (O_2053,N_24715,N_24736);
xor UO_2054 (O_2054,N_24715,N_24682);
nand UO_2055 (O_2055,N_24434,N_24411);
nand UO_2056 (O_2056,N_24700,N_24719);
xor UO_2057 (O_2057,N_24786,N_24636);
nand UO_2058 (O_2058,N_24642,N_24864);
xnor UO_2059 (O_2059,N_24767,N_24884);
nor UO_2060 (O_2060,N_24914,N_24945);
xor UO_2061 (O_2061,N_24895,N_24500);
xnor UO_2062 (O_2062,N_24750,N_24812);
nor UO_2063 (O_2063,N_24575,N_24502);
and UO_2064 (O_2064,N_24463,N_24895);
nor UO_2065 (O_2065,N_24378,N_24898);
or UO_2066 (O_2066,N_24748,N_24741);
or UO_2067 (O_2067,N_24830,N_24651);
xor UO_2068 (O_2068,N_24746,N_24830);
nor UO_2069 (O_2069,N_24674,N_24892);
nor UO_2070 (O_2070,N_24410,N_24704);
xnor UO_2071 (O_2071,N_24595,N_24989);
nor UO_2072 (O_2072,N_24955,N_24880);
or UO_2073 (O_2073,N_24623,N_24695);
xnor UO_2074 (O_2074,N_24697,N_24807);
or UO_2075 (O_2075,N_24826,N_24815);
and UO_2076 (O_2076,N_24774,N_24570);
xnor UO_2077 (O_2077,N_24776,N_24574);
and UO_2078 (O_2078,N_24800,N_24693);
nand UO_2079 (O_2079,N_24967,N_24565);
nor UO_2080 (O_2080,N_24737,N_24451);
nor UO_2081 (O_2081,N_24958,N_24980);
nand UO_2082 (O_2082,N_24659,N_24871);
and UO_2083 (O_2083,N_24380,N_24670);
xnor UO_2084 (O_2084,N_24646,N_24386);
nor UO_2085 (O_2085,N_24393,N_24816);
nor UO_2086 (O_2086,N_24433,N_24422);
and UO_2087 (O_2087,N_24421,N_24808);
nand UO_2088 (O_2088,N_24626,N_24861);
or UO_2089 (O_2089,N_24742,N_24693);
nand UO_2090 (O_2090,N_24968,N_24410);
and UO_2091 (O_2091,N_24850,N_24911);
nor UO_2092 (O_2092,N_24693,N_24916);
or UO_2093 (O_2093,N_24943,N_24850);
nor UO_2094 (O_2094,N_24949,N_24447);
nor UO_2095 (O_2095,N_24526,N_24941);
and UO_2096 (O_2096,N_24413,N_24574);
nand UO_2097 (O_2097,N_24990,N_24464);
and UO_2098 (O_2098,N_24825,N_24603);
nand UO_2099 (O_2099,N_24850,N_24807);
nand UO_2100 (O_2100,N_24890,N_24895);
and UO_2101 (O_2101,N_24766,N_24997);
and UO_2102 (O_2102,N_24404,N_24625);
or UO_2103 (O_2103,N_24783,N_24751);
nand UO_2104 (O_2104,N_24456,N_24534);
nor UO_2105 (O_2105,N_24437,N_24909);
or UO_2106 (O_2106,N_24606,N_24598);
and UO_2107 (O_2107,N_24983,N_24710);
and UO_2108 (O_2108,N_24901,N_24884);
nor UO_2109 (O_2109,N_24517,N_24962);
nand UO_2110 (O_2110,N_24602,N_24385);
xnor UO_2111 (O_2111,N_24783,N_24460);
and UO_2112 (O_2112,N_24697,N_24749);
or UO_2113 (O_2113,N_24529,N_24581);
and UO_2114 (O_2114,N_24502,N_24388);
xnor UO_2115 (O_2115,N_24805,N_24824);
and UO_2116 (O_2116,N_24892,N_24932);
or UO_2117 (O_2117,N_24779,N_24649);
nor UO_2118 (O_2118,N_24713,N_24682);
xnor UO_2119 (O_2119,N_24852,N_24553);
xor UO_2120 (O_2120,N_24647,N_24916);
or UO_2121 (O_2121,N_24923,N_24780);
and UO_2122 (O_2122,N_24845,N_24886);
xor UO_2123 (O_2123,N_24725,N_24595);
nand UO_2124 (O_2124,N_24655,N_24701);
and UO_2125 (O_2125,N_24682,N_24462);
nand UO_2126 (O_2126,N_24709,N_24830);
and UO_2127 (O_2127,N_24490,N_24659);
or UO_2128 (O_2128,N_24665,N_24430);
or UO_2129 (O_2129,N_24769,N_24912);
or UO_2130 (O_2130,N_24505,N_24918);
xnor UO_2131 (O_2131,N_24802,N_24556);
xor UO_2132 (O_2132,N_24829,N_24914);
nor UO_2133 (O_2133,N_24526,N_24716);
and UO_2134 (O_2134,N_24724,N_24991);
and UO_2135 (O_2135,N_24543,N_24986);
nand UO_2136 (O_2136,N_24705,N_24865);
nand UO_2137 (O_2137,N_24402,N_24592);
nand UO_2138 (O_2138,N_24661,N_24558);
or UO_2139 (O_2139,N_24476,N_24623);
or UO_2140 (O_2140,N_24744,N_24601);
nand UO_2141 (O_2141,N_24977,N_24728);
or UO_2142 (O_2142,N_24419,N_24482);
nor UO_2143 (O_2143,N_24475,N_24927);
xor UO_2144 (O_2144,N_24714,N_24666);
and UO_2145 (O_2145,N_24725,N_24909);
xnor UO_2146 (O_2146,N_24380,N_24552);
xnor UO_2147 (O_2147,N_24378,N_24710);
and UO_2148 (O_2148,N_24708,N_24390);
or UO_2149 (O_2149,N_24791,N_24683);
nor UO_2150 (O_2150,N_24540,N_24593);
nor UO_2151 (O_2151,N_24749,N_24417);
xor UO_2152 (O_2152,N_24416,N_24679);
nand UO_2153 (O_2153,N_24544,N_24888);
nand UO_2154 (O_2154,N_24606,N_24809);
and UO_2155 (O_2155,N_24591,N_24566);
xnor UO_2156 (O_2156,N_24752,N_24778);
nand UO_2157 (O_2157,N_24943,N_24385);
nand UO_2158 (O_2158,N_24601,N_24835);
xor UO_2159 (O_2159,N_24588,N_24380);
nand UO_2160 (O_2160,N_24884,N_24625);
nand UO_2161 (O_2161,N_24889,N_24650);
nor UO_2162 (O_2162,N_24707,N_24776);
nand UO_2163 (O_2163,N_24525,N_24908);
nor UO_2164 (O_2164,N_24951,N_24943);
and UO_2165 (O_2165,N_24535,N_24762);
and UO_2166 (O_2166,N_24733,N_24885);
nand UO_2167 (O_2167,N_24550,N_24534);
xnor UO_2168 (O_2168,N_24513,N_24864);
xor UO_2169 (O_2169,N_24874,N_24640);
nand UO_2170 (O_2170,N_24719,N_24757);
or UO_2171 (O_2171,N_24703,N_24549);
nor UO_2172 (O_2172,N_24683,N_24808);
xnor UO_2173 (O_2173,N_24381,N_24869);
and UO_2174 (O_2174,N_24421,N_24788);
or UO_2175 (O_2175,N_24445,N_24720);
nor UO_2176 (O_2176,N_24847,N_24736);
xor UO_2177 (O_2177,N_24514,N_24754);
nand UO_2178 (O_2178,N_24574,N_24754);
nand UO_2179 (O_2179,N_24853,N_24961);
nand UO_2180 (O_2180,N_24436,N_24784);
nand UO_2181 (O_2181,N_24656,N_24736);
nand UO_2182 (O_2182,N_24755,N_24497);
nor UO_2183 (O_2183,N_24796,N_24682);
and UO_2184 (O_2184,N_24733,N_24840);
xnor UO_2185 (O_2185,N_24387,N_24402);
or UO_2186 (O_2186,N_24881,N_24463);
and UO_2187 (O_2187,N_24885,N_24437);
nor UO_2188 (O_2188,N_24634,N_24972);
nor UO_2189 (O_2189,N_24488,N_24950);
xnor UO_2190 (O_2190,N_24476,N_24863);
or UO_2191 (O_2191,N_24552,N_24404);
xor UO_2192 (O_2192,N_24544,N_24703);
and UO_2193 (O_2193,N_24640,N_24593);
xnor UO_2194 (O_2194,N_24947,N_24495);
xnor UO_2195 (O_2195,N_24504,N_24697);
xnor UO_2196 (O_2196,N_24714,N_24807);
nor UO_2197 (O_2197,N_24945,N_24603);
xor UO_2198 (O_2198,N_24522,N_24503);
nor UO_2199 (O_2199,N_24935,N_24895);
and UO_2200 (O_2200,N_24897,N_24592);
and UO_2201 (O_2201,N_24415,N_24816);
nand UO_2202 (O_2202,N_24666,N_24845);
nand UO_2203 (O_2203,N_24791,N_24491);
nand UO_2204 (O_2204,N_24693,N_24782);
and UO_2205 (O_2205,N_24498,N_24617);
nand UO_2206 (O_2206,N_24710,N_24986);
xor UO_2207 (O_2207,N_24696,N_24934);
nand UO_2208 (O_2208,N_24564,N_24677);
and UO_2209 (O_2209,N_24684,N_24581);
and UO_2210 (O_2210,N_24808,N_24554);
xnor UO_2211 (O_2211,N_24939,N_24628);
nor UO_2212 (O_2212,N_24742,N_24475);
or UO_2213 (O_2213,N_24961,N_24848);
or UO_2214 (O_2214,N_24835,N_24440);
or UO_2215 (O_2215,N_24965,N_24998);
or UO_2216 (O_2216,N_24858,N_24915);
xnor UO_2217 (O_2217,N_24570,N_24880);
xor UO_2218 (O_2218,N_24742,N_24896);
nand UO_2219 (O_2219,N_24796,N_24391);
or UO_2220 (O_2220,N_24405,N_24960);
and UO_2221 (O_2221,N_24494,N_24557);
nor UO_2222 (O_2222,N_24547,N_24467);
and UO_2223 (O_2223,N_24538,N_24698);
nor UO_2224 (O_2224,N_24529,N_24849);
xor UO_2225 (O_2225,N_24872,N_24449);
xnor UO_2226 (O_2226,N_24568,N_24714);
and UO_2227 (O_2227,N_24997,N_24794);
nor UO_2228 (O_2228,N_24823,N_24647);
and UO_2229 (O_2229,N_24413,N_24978);
or UO_2230 (O_2230,N_24611,N_24928);
or UO_2231 (O_2231,N_24422,N_24843);
or UO_2232 (O_2232,N_24430,N_24673);
or UO_2233 (O_2233,N_24461,N_24501);
nand UO_2234 (O_2234,N_24525,N_24433);
nand UO_2235 (O_2235,N_24639,N_24714);
or UO_2236 (O_2236,N_24911,N_24829);
nor UO_2237 (O_2237,N_24749,N_24624);
nor UO_2238 (O_2238,N_24870,N_24595);
xor UO_2239 (O_2239,N_24569,N_24694);
or UO_2240 (O_2240,N_24434,N_24582);
xnor UO_2241 (O_2241,N_24614,N_24378);
or UO_2242 (O_2242,N_24473,N_24654);
nand UO_2243 (O_2243,N_24567,N_24544);
and UO_2244 (O_2244,N_24836,N_24388);
and UO_2245 (O_2245,N_24852,N_24871);
xor UO_2246 (O_2246,N_24473,N_24860);
or UO_2247 (O_2247,N_24610,N_24715);
nand UO_2248 (O_2248,N_24734,N_24565);
or UO_2249 (O_2249,N_24480,N_24893);
nor UO_2250 (O_2250,N_24398,N_24842);
nand UO_2251 (O_2251,N_24888,N_24612);
or UO_2252 (O_2252,N_24385,N_24951);
nor UO_2253 (O_2253,N_24487,N_24826);
xor UO_2254 (O_2254,N_24451,N_24666);
nor UO_2255 (O_2255,N_24518,N_24928);
nor UO_2256 (O_2256,N_24707,N_24402);
or UO_2257 (O_2257,N_24862,N_24474);
or UO_2258 (O_2258,N_24483,N_24508);
nor UO_2259 (O_2259,N_24505,N_24719);
or UO_2260 (O_2260,N_24697,N_24522);
or UO_2261 (O_2261,N_24678,N_24958);
xnor UO_2262 (O_2262,N_24745,N_24524);
and UO_2263 (O_2263,N_24804,N_24578);
or UO_2264 (O_2264,N_24807,N_24566);
nor UO_2265 (O_2265,N_24531,N_24498);
or UO_2266 (O_2266,N_24533,N_24500);
nand UO_2267 (O_2267,N_24522,N_24423);
and UO_2268 (O_2268,N_24390,N_24852);
or UO_2269 (O_2269,N_24719,N_24765);
nand UO_2270 (O_2270,N_24651,N_24826);
and UO_2271 (O_2271,N_24418,N_24564);
or UO_2272 (O_2272,N_24815,N_24977);
nor UO_2273 (O_2273,N_24524,N_24846);
nand UO_2274 (O_2274,N_24621,N_24450);
or UO_2275 (O_2275,N_24389,N_24460);
and UO_2276 (O_2276,N_24585,N_24869);
xor UO_2277 (O_2277,N_24598,N_24841);
nor UO_2278 (O_2278,N_24989,N_24947);
xnor UO_2279 (O_2279,N_24426,N_24812);
nor UO_2280 (O_2280,N_24941,N_24608);
xor UO_2281 (O_2281,N_24853,N_24861);
xor UO_2282 (O_2282,N_24574,N_24934);
xnor UO_2283 (O_2283,N_24769,N_24783);
nor UO_2284 (O_2284,N_24646,N_24393);
xor UO_2285 (O_2285,N_24423,N_24877);
xnor UO_2286 (O_2286,N_24577,N_24894);
nor UO_2287 (O_2287,N_24637,N_24817);
or UO_2288 (O_2288,N_24471,N_24772);
or UO_2289 (O_2289,N_24633,N_24473);
xor UO_2290 (O_2290,N_24862,N_24769);
nor UO_2291 (O_2291,N_24433,N_24669);
xnor UO_2292 (O_2292,N_24647,N_24828);
nand UO_2293 (O_2293,N_24576,N_24706);
nor UO_2294 (O_2294,N_24594,N_24925);
xor UO_2295 (O_2295,N_24792,N_24816);
nor UO_2296 (O_2296,N_24909,N_24447);
or UO_2297 (O_2297,N_24698,N_24969);
nor UO_2298 (O_2298,N_24736,N_24486);
xor UO_2299 (O_2299,N_24812,N_24866);
xnor UO_2300 (O_2300,N_24639,N_24854);
or UO_2301 (O_2301,N_24919,N_24490);
or UO_2302 (O_2302,N_24633,N_24440);
nand UO_2303 (O_2303,N_24824,N_24629);
and UO_2304 (O_2304,N_24699,N_24765);
nand UO_2305 (O_2305,N_24633,N_24412);
and UO_2306 (O_2306,N_24825,N_24436);
or UO_2307 (O_2307,N_24583,N_24976);
or UO_2308 (O_2308,N_24847,N_24584);
and UO_2309 (O_2309,N_24964,N_24939);
nor UO_2310 (O_2310,N_24538,N_24527);
and UO_2311 (O_2311,N_24717,N_24994);
nor UO_2312 (O_2312,N_24871,N_24975);
nand UO_2313 (O_2313,N_24697,N_24598);
nand UO_2314 (O_2314,N_24990,N_24391);
and UO_2315 (O_2315,N_24803,N_24862);
nor UO_2316 (O_2316,N_24448,N_24533);
xnor UO_2317 (O_2317,N_24455,N_24472);
or UO_2318 (O_2318,N_24742,N_24601);
or UO_2319 (O_2319,N_24785,N_24806);
or UO_2320 (O_2320,N_24580,N_24774);
nand UO_2321 (O_2321,N_24681,N_24968);
or UO_2322 (O_2322,N_24729,N_24712);
nand UO_2323 (O_2323,N_24453,N_24413);
nand UO_2324 (O_2324,N_24378,N_24544);
nor UO_2325 (O_2325,N_24807,N_24878);
or UO_2326 (O_2326,N_24557,N_24413);
xor UO_2327 (O_2327,N_24973,N_24523);
xor UO_2328 (O_2328,N_24393,N_24447);
or UO_2329 (O_2329,N_24979,N_24865);
nor UO_2330 (O_2330,N_24957,N_24800);
xor UO_2331 (O_2331,N_24709,N_24664);
or UO_2332 (O_2332,N_24890,N_24519);
and UO_2333 (O_2333,N_24654,N_24879);
nor UO_2334 (O_2334,N_24561,N_24883);
and UO_2335 (O_2335,N_24546,N_24945);
nor UO_2336 (O_2336,N_24407,N_24734);
xor UO_2337 (O_2337,N_24936,N_24606);
and UO_2338 (O_2338,N_24629,N_24883);
or UO_2339 (O_2339,N_24901,N_24715);
nor UO_2340 (O_2340,N_24997,N_24506);
xnor UO_2341 (O_2341,N_24551,N_24465);
nor UO_2342 (O_2342,N_24615,N_24445);
nor UO_2343 (O_2343,N_24487,N_24776);
nand UO_2344 (O_2344,N_24511,N_24657);
xnor UO_2345 (O_2345,N_24906,N_24990);
nor UO_2346 (O_2346,N_24984,N_24378);
xor UO_2347 (O_2347,N_24969,N_24960);
or UO_2348 (O_2348,N_24593,N_24927);
nor UO_2349 (O_2349,N_24744,N_24713);
xnor UO_2350 (O_2350,N_24473,N_24536);
or UO_2351 (O_2351,N_24712,N_24782);
nor UO_2352 (O_2352,N_24876,N_24685);
nor UO_2353 (O_2353,N_24610,N_24531);
and UO_2354 (O_2354,N_24950,N_24746);
nand UO_2355 (O_2355,N_24908,N_24784);
and UO_2356 (O_2356,N_24545,N_24699);
nor UO_2357 (O_2357,N_24557,N_24991);
and UO_2358 (O_2358,N_24981,N_24379);
or UO_2359 (O_2359,N_24964,N_24523);
xor UO_2360 (O_2360,N_24787,N_24848);
xor UO_2361 (O_2361,N_24605,N_24598);
and UO_2362 (O_2362,N_24551,N_24455);
or UO_2363 (O_2363,N_24650,N_24440);
and UO_2364 (O_2364,N_24926,N_24462);
nor UO_2365 (O_2365,N_24573,N_24810);
or UO_2366 (O_2366,N_24645,N_24451);
or UO_2367 (O_2367,N_24886,N_24452);
nor UO_2368 (O_2368,N_24418,N_24760);
or UO_2369 (O_2369,N_24718,N_24812);
and UO_2370 (O_2370,N_24574,N_24756);
nor UO_2371 (O_2371,N_24694,N_24878);
nor UO_2372 (O_2372,N_24692,N_24563);
xnor UO_2373 (O_2373,N_24439,N_24426);
xnor UO_2374 (O_2374,N_24828,N_24683);
and UO_2375 (O_2375,N_24449,N_24793);
or UO_2376 (O_2376,N_24713,N_24706);
xor UO_2377 (O_2377,N_24869,N_24752);
nand UO_2378 (O_2378,N_24758,N_24498);
or UO_2379 (O_2379,N_24620,N_24685);
nor UO_2380 (O_2380,N_24989,N_24394);
nor UO_2381 (O_2381,N_24885,N_24758);
nand UO_2382 (O_2382,N_24514,N_24931);
and UO_2383 (O_2383,N_24603,N_24796);
and UO_2384 (O_2384,N_24872,N_24541);
nor UO_2385 (O_2385,N_24987,N_24554);
or UO_2386 (O_2386,N_24431,N_24579);
or UO_2387 (O_2387,N_24487,N_24845);
and UO_2388 (O_2388,N_24631,N_24742);
and UO_2389 (O_2389,N_24959,N_24463);
nand UO_2390 (O_2390,N_24693,N_24422);
nand UO_2391 (O_2391,N_24384,N_24705);
and UO_2392 (O_2392,N_24973,N_24639);
xnor UO_2393 (O_2393,N_24709,N_24385);
xnor UO_2394 (O_2394,N_24611,N_24706);
nand UO_2395 (O_2395,N_24453,N_24742);
nand UO_2396 (O_2396,N_24424,N_24846);
and UO_2397 (O_2397,N_24610,N_24579);
and UO_2398 (O_2398,N_24823,N_24683);
or UO_2399 (O_2399,N_24958,N_24634);
nor UO_2400 (O_2400,N_24438,N_24833);
or UO_2401 (O_2401,N_24523,N_24489);
xnor UO_2402 (O_2402,N_24743,N_24652);
and UO_2403 (O_2403,N_24926,N_24441);
nand UO_2404 (O_2404,N_24690,N_24472);
nor UO_2405 (O_2405,N_24949,N_24805);
or UO_2406 (O_2406,N_24880,N_24733);
nor UO_2407 (O_2407,N_24466,N_24881);
and UO_2408 (O_2408,N_24411,N_24591);
and UO_2409 (O_2409,N_24811,N_24504);
or UO_2410 (O_2410,N_24959,N_24890);
nand UO_2411 (O_2411,N_24703,N_24963);
xnor UO_2412 (O_2412,N_24816,N_24453);
nand UO_2413 (O_2413,N_24390,N_24576);
nor UO_2414 (O_2414,N_24442,N_24424);
xnor UO_2415 (O_2415,N_24883,N_24449);
nand UO_2416 (O_2416,N_24388,N_24389);
or UO_2417 (O_2417,N_24431,N_24742);
or UO_2418 (O_2418,N_24940,N_24545);
and UO_2419 (O_2419,N_24559,N_24402);
xnor UO_2420 (O_2420,N_24893,N_24656);
or UO_2421 (O_2421,N_24412,N_24411);
or UO_2422 (O_2422,N_24755,N_24606);
or UO_2423 (O_2423,N_24452,N_24380);
or UO_2424 (O_2424,N_24532,N_24908);
nor UO_2425 (O_2425,N_24967,N_24614);
and UO_2426 (O_2426,N_24875,N_24592);
xnor UO_2427 (O_2427,N_24859,N_24733);
or UO_2428 (O_2428,N_24500,N_24571);
xnor UO_2429 (O_2429,N_24413,N_24827);
xnor UO_2430 (O_2430,N_24435,N_24993);
nor UO_2431 (O_2431,N_24979,N_24674);
xor UO_2432 (O_2432,N_24858,N_24407);
or UO_2433 (O_2433,N_24397,N_24612);
xor UO_2434 (O_2434,N_24698,N_24765);
or UO_2435 (O_2435,N_24570,N_24779);
xnor UO_2436 (O_2436,N_24930,N_24579);
nor UO_2437 (O_2437,N_24391,N_24844);
nor UO_2438 (O_2438,N_24789,N_24891);
xor UO_2439 (O_2439,N_24597,N_24745);
and UO_2440 (O_2440,N_24839,N_24915);
and UO_2441 (O_2441,N_24929,N_24506);
xnor UO_2442 (O_2442,N_24443,N_24667);
and UO_2443 (O_2443,N_24672,N_24986);
xor UO_2444 (O_2444,N_24845,N_24732);
or UO_2445 (O_2445,N_24579,N_24641);
or UO_2446 (O_2446,N_24465,N_24845);
nand UO_2447 (O_2447,N_24722,N_24901);
nand UO_2448 (O_2448,N_24893,N_24629);
nor UO_2449 (O_2449,N_24472,N_24381);
nand UO_2450 (O_2450,N_24570,N_24983);
and UO_2451 (O_2451,N_24781,N_24896);
and UO_2452 (O_2452,N_24816,N_24948);
nor UO_2453 (O_2453,N_24601,N_24417);
or UO_2454 (O_2454,N_24997,N_24565);
xnor UO_2455 (O_2455,N_24448,N_24975);
and UO_2456 (O_2456,N_24733,N_24427);
xnor UO_2457 (O_2457,N_24888,N_24391);
nand UO_2458 (O_2458,N_24808,N_24709);
and UO_2459 (O_2459,N_24633,N_24529);
nand UO_2460 (O_2460,N_24926,N_24471);
and UO_2461 (O_2461,N_24856,N_24872);
xnor UO_2462 (O_2462,N_24975,N_24632);
nor UO_2463 (O_2463,N_24650,N_24929);
nand UO_2464 (O_2464,N_24663,N_24715);
xor UO_2465 (O_2465,N_24950,N_24407);
nor UO_2466 (O_2466,N_24425,N_24764);
nand UO_2467 (O_2467,N_24839,N_24942);
nor UO_2468 (O_2468,N_24583,N_24603);
or UO_2469 (O_2469,N_24658,N_24489);
and UO_2470 (O_2470,N_24504,N_24632);
nand UO_2471 (O_2471,N_24548,N_24666);
nor UO_2472 (O_2472,N_24432,N_24945);
xnor UO_2473 (O_2473,N_24886,N_24929);
nor UO_2474 (O_2474,N_24937,N_24777);
xor UO_2475 (O_2475,N_24983,N_24399);
nand UO_2476 (O_2476,N_24415,N_24555);
xor UO_2477 (O_2477,N_24636,N_24379);
or UO_2478 (O_2478,N_24712,N_24942);
nand UO_2479 (O_2479,N_24635,N_24733);
nand UO_2480 (O_2480,N_24381,N_24793);
and UO_2481 (O_2481,N_24652,N_24691);
and UO_2482 (O_2482,N_24787,N_24493);
nor UO_2483 (O_2483,N_24635,N_24435);
nor UO_2484 (O_2484,N_24928,N_24375);
or UO_2485 (O_2485,N_24705,N_24786);
and UO_2486 (O_2486,N_24776,N_24889);
and UO_2487 (O_2487,N_24704,N_24945);
xnor UO_2488 (O_2488,N_24867,N_24811);
xor UO_2489 (O_2489,N_24700,N_24672);
nand UO_2490 (O_2490,N_24427,N_24601);
xor UO_2491 (O_2491,N_24473,N_24507);
or UO_2492 (O_2492,N_24786,N_24906);
and UO_2493 (O_2493,N_24637,N_24776);
nand UO_2494 (O_2494,N_24500,N_24911);
nand UO_2495 (O_2495,N_24416,N_24664);
or UO_2496 (O_2496,N_24425,N_24622);
and UO_2497 (O_2497,N_24859,N_24854);
and UO_2498 (O_2498,N_24573,N_24630);
nand UO_2499 (O_2499,N_24890,N_24941);
and UO_2500 (O_2500,N_24638,N_24533);
or UO_2501 (O_2501,N_24708,N_24459);
nor UO_2502 (O_2502,N_24409,N_24515);
nor UO_2503 (O_2503,N_24847,N_24571);
xor UO_2504 (O_2504,N_24775,N_24380);
and UO_2505 (O_2505,N_24674,N_24437);
nand UO_2506 (O_2506,N_24376,N_24990);
or UO_2507 (O_2507,N_24538,N_24963);
and UO_2508 (O_2508,N_24736,N_24918);
nor UO_2509 (O_2509,N_24747,N_24574);
and UO_2510 (O_2510,N_24381,N_24467);
nand UO_2511 (O_2511,N_24807,N_24439);
or UO_2512 (O_2512,N_24628,N_24617);
nor UO_2513 (O_2513,N_24385,N_24612);
or UO_2514 (O_2514,N_24555,N_24937);
xnor UO_2515 (O_2515,N_24538,N_24543);
nor UO_2516 (O_2516,N_24472,N_24999);
xor UO_2517 (O_2517,N_24831,N_24811);
xnor UO_2518 (O_2518,N_24899,N_24920);
nand UO_2519 (O_2519,N_24721,N_24549);
or UO_2520 (O_2520,N_24559,N_24967);
and UO_2521 (O_2521,N_24505,N_24909);
xor UO_2522 (O_2522,N_24938,N_24838);
and UO_2523 (O_2523,N_24720,N_24721);
or UO_2524 (O_2524,N_24464,N_24435);
nand UO_2525 (O_2525,N_24587,N_24627);
nor UO_2526 (O_2526,N_24858,N_24691);
xor UO_2527 (O_2527,N_24413,N_24583);
nand UO_2528 (O_2528,N_24723,N_24665);
or UO_2529 (O_2529,N_24699,N_24820);
nand UO_2530 (O_2530,N_24464,N_24405);
nor UO_2531 (O_2531,N_24398,N_24519);
nor UO_2532 (O_2532,N_24659,N_24483);
nand UO_2533 (O_2533,N_24410,N_24713);
nand UO_2534 (O_2534,N_24574,N_24486);
xor UO_2535 (O_2535,N_24426,N_24774);
and UO_2536 (O_2536,N_24726,N_24732);
or UO_2537 (O_2537,N_24690,N_24834);
and UO_2538 (O_2538,N_24584,N_24396);
or UO_2539 (O_2539,N_24985,N_24860);
and UO_2540 (O_2540,N_24962,N_24833);
nand UO_2541 (O_2541,N_24824,N_24905);
and UO_2542 (O_2542,N_24480,N_24489);
and UO_2543 (O_2543,N_24624,N_24739);
xor UO_2544 (O_2544,N_24592,N_24523);
or UO_2545 (O_2545,N_24794,N_24974);
xnor UO_2546 (O_2546,N_24821,N_24805);
nor UO_2547 (O_2547,N_24580,N_24586);
and UO_2548 (O_2548,N_24914,N_24640);
and UO_2549 (O_2549,N_24388,N_24806);
and UO_2550 (O_2550,N_24586,N_24381);
xnor UO_2551 (O_2551,N_24580,N_24991);
xnor UO_2552 (O_2552,N_24642,N_24763);
or UO_2553 (O_2553,N_24925,N_24870);
nand UO_2554 (O_2554,N_24784,N_24531);
or UO_2555 (O_2555,N_24919,N_24765);
or UO_2556 (O_2556,N_24560,N_24739);
nor UO_2557 (O_2557,N_24835,N_24478);
or UO_2558 (O_2558,N_24398,N_24594);
xor UO_2559 (O_2559,N_24781,N_24909);
nor UO_2560 (O_2560,N_24799,N_24518);
nor UO_2561 (O_2561,N_24440,N_24961);
xor UO_2562 (O_2562,N_24977,N_24382);
xor UO_2563 (O_2563,N_24588,N_24576);
nand UO_2564 (O_2564,N_24422,N_24746);
xnor UO_2565 (O_2565,N_24440,N_24873);
and UO_2566 (O_2566,N_24745,N_24989);
or UO_2567 (O_2567,N_24865,N_24627);
or UO_2568 (O_2568,N_24716,N_24625);
nor UO_2569 (O_2569,N_24820,N_24619);
or UO_2570 (O_2570,N_24442,N_24769);
or UO_2571 (O_2571,N_24839,N_24986);
nand UO_2572 (O_2572,N_24839,N_24618);
nand UO_2573 (O_2573,N_24623,N_24745);
and UO_2574 (O_2574,N_24952,N_24602);
or UO_2575 (O_2575,N_24588,N_24636);
nor UO_2576 (O_2576,N_24431,N_24918);
or UO_2577 (O_2577,N_24817,N_24930);
nand UO_2578 (O_2578,N_24539,N_24524);
and UO_2579 (O_2579,N_24771,N_24847);
nand UO_2580 (O_2580,N_24470,N_24753);
nor UO_2581 (O_2581,N_24843,N_24557);
and UO_2582 (O_2582,N_24742,N_24864);
or UO_2583 (O_2583,N_24724,N_24906);
and UO_2584 (O_2584,N_24727,N_24599);
nand UO_2585 (O_2585,N_24945,N_24859);
xor UO_2586 (O_2586,N_24962,N_24944);
nand UO_2587 (O_2587,N_24389,N_24864);
or UO_2588 (O_2588,N_24628,N_24777);
and UO_2589 (O_2589,N_24594,N_24999);
xor UO_2590 (O_2590,N_24661,N_24538);
nor UO_2591 (O_2591,N_24433,N_24634);
or UO_2592 (O_2592,N_24755,N_24963);
or UO_2593 (O_2593,N_24645,N_24659);
xnor UO_2594 (O_2594,N_24692,N_24999);
nand UO_2595 (O_2595,N_24620,N_24512);
xor UO_2596 (O_2596,N_24658,N_24823);
or UO_2597 (O_2597,N_24644,N_24963);
nor UO_2598 (O_2598,N_24415,N_24731);
and UO_2599 (O_2599,N_24773,N_24856);
xnor UO_2600 (O_2600,N_24709,N_24736);
and UO_2601 (O_2601,N_24866,N_24959);
nor UO_2602 (O_2602,N_24447,N_24509);
nand UO_2603 (O_2603,N_24762,N_24502);
or UO_2604 (O_2604,N_24416,N_24602);
nor UO_2605 (O_2605,N_24525,N_24745);
nand UO_2606 (O_2606,N_24577,N_24837);
xnor UO_2607 (O_2607,N_24531,N_24493);
nand UO_2608 (O_2608,N_24399,N_24701);
nor UO_2609 (O_2609,N_24997,N_24627);
nor UO_2610 (O_2610,N_24445,N_24433);
nand UO_2611 (O_2611,N_24626,N_24988);
or UO_2612 (O_2612,N_24434,N_24385);
nor UO_2613 (O_2613,N_24643,N_24912);
or UO_2614 (O_2614,N_24669,N_24901);
nor UO_2615 (O_2615,N_24754,N_24430);
nor UO_2616 (O_2616,N_24793,N_24643);
or UO_2617 (O_2617,N_24782,N_24529);
or UO_2618 (O_2618,N_24739,N_24537);
and UO_2619 (O_2619,N_24847,N_24705);
or UO_2620 (O_2620,N_24458,N_24777);
xor UO_2621 (O_2621,N_24830,N_24525);
or UO_2622 (O_2622,N_24917,N_24441);
and UO_2623 (O_2623,N_24526,N_24880);
or UO_2624 (O_2624,N_24933,N_24997);
nand UO_2625 (O_2625,N_24905,N_24513);
nor UO_2626 (O_2626,N_24733,N_24620);
nand UO_2627 (O_2627,N_24869,N_24837);
nand UO_2628 (O_2628,N_24977,N_24673);
and UO_2629 (O_2629,N_24838,N_24375);
nor UO_2630 (O_2630,N_24412,N_24846);
and UO_2631 (O_2631,N_24715,N_24760);
and UO_2632 (O_2632,N_24806,N_24693);
xnor UO_2633 (O_2633,N_24758,N_24927);
or UO_2634 (O_2634,N_24530,N_24945);
nor UO_2635 (O_2635,N_24733,N_24500);
and UO_2636 (O_2636,N_24482,N_24497);
nor UO_2637 (O_2637,N_24699,N_24378);
and UO_2638 (O_2638,N_24440,N_24738);
and UO_2639 (O_2639,N_24542,N_24894);
xnor UO_2640 (O_2640,N_24785,N_24396);
or UO_2641 (O_2641,N_24917,N_24443);
xnor UO_2642 (O_2642,N_24542,N_24578);
xnor UO_2643 (O_2643,N_24504,N_24615);
xor UO_2644 (O_2644,N_24401,N_24793);
or UO_2645 (O_2645,N_24494,N_24555);
nor UO_2646 (O_2646,N_24716,N_24421);
nor UO_2647 (O_2647,N_24443,N_24469);
nand UO_2648 (O_2648,N_24993,N_24783);
xor UO_2649 (O_2649,N_24519,N_24642);
or UO_2650 (O_2650,N_24808,N_24673);
and UO_2651 (O_2651,N_24452,N_24555);
nand UO_2652 (O_2652,N_24390,N_24724);
and UO_2653 (O_2653,N_24589,N_24546);
or UO_2654 (O_2654,N_24997,N_24765);
or UO_2655 (O_2655,N_24876,N_24680);
or UO_2656 (O_2656,N_24855,N_24960);
or UO_2657 (O_2657,N_24441,N_24688);
and UO_2658 (O_2658,N_24692,N_24680);
nand UO_2659 (O_2659,N_24693,N_24804);
and UO_2660 (O_2660,N_24819,N_24633);
xnor UO_2661 (O_2661,N_24440,N_24750);
nor UO_2662 (O_2662,N_24541,N_24724);
nand UO_2663 (O_2663,N_24951,N_24960);
xnor UO_2664 (O_2664,N_24965,N_24532);
xnor UO_2665 (O_2665,N_24399,N_24783);
nand UO_2666 (O_2666,N_24917,N_24777);
xor UO_2667 (O_2667,N_24439,N_24682);
nand UO_2668 (O_2668,N_24857,N_24517);
and UO_2669 (O_2669,N_24446,N_24621);
nand UO_2670 (O_2670,N_24997,N_24914);
and UO_2671 (O_2671,N_24799,N_24744);
nor UO_2672 (O_2672,N_24600,N_24940);
and UO_2673 (O_2673,N_24885,N_24982);
or UO_2674 (O_2674,N_24422,N_24993);
or UO_2675 (O_2675,N_24468,N_24430);
and UO_2676 (O_2676,N_24930,N_24838);
or UO_2677 (O_2677,N_24712,N_24810);
and UO_2678 (O_2678,N_24633,N_24378);
and UO_2679 (O_2679,N_24671,N_24599);
and UO_2680 (O_2680,N_24492,N_24775);
nor UO_2681 (O_2681,N_24704,N_24543);
nor UO_2682 (O_2682,N_24737,N_24840);
xnor UO_2683 (O_2683,N_24930,N_24576);
and UO_2684 (O_2684,N_24981,N_24474);
nand UO_2685 (O_2685,N_24639,N_24466);
xor UO_2686 (O_2686,N_24776,N_24713);
nor UO_2687 (O_2687,N_24462,N_24412);
nor UO_2688 (O_2688,N_24836,N_24567);
or UO_2689 (O_2689,N_24447,N_24479);
nand UO_2690 (O_2690,N_24930,N_24436);
or UO_2691 (O_2691,N_24657,N_24750);
nand UO_2692 (O_2692,N_24443,N_24790);
xor UO_2693 (O_2693,N_24943,N_24993);
xor UO_2694 (O_2694,N_24977,N_24523);
nor UO_2695 (O_2695,N_24556,N_24669);
or UO_2696 (O_2696,N_24735,N_24707);
and UO_2697 (O_2697,N_24981,N_24500);
xor UO_2698 (O_2698,N_24820,N_24472);
and UO_2699 (O_2699,N_24750,N_24419);
and UO_2700 (O_2700,N_24385,N_24578);
xor UO_2701 (O_2701,N_24852,N_24454);
or UO_2702 (O_2702,N_24591,N_24568);
or UO_2703 (O_2703,N_24489,N_24414);
xor UO_2704 (O_2704,N_24528,N_24955);
nor UO_2705 (O_2705,N_24916,N_24531);
nor UO_2706 (O_2706,N_24520,N_24409);
nand UO_2707 (O_2707,N_24594,N_24906);
or UO_2708 (O_2708,N_24480,N_24824);
or UO_2709 (O_2709,N_24915,N_24448);
xor UO_2710 (O_2710,N_24951,N_24846);
nor UO_2711 (O_2711,N_24996,N_24633);
or UO_2712 (O_2712,N_24804,N_24758);
or UO_2713 (O_2713,N_24836,N_24586);
nor UO_2714 (O_2714,N_24653,N_24940);
nor UO_2715 (O_2715,N_24435,N_24894);
or UO_2716 (O_2716,N_24757,N_24408);
nor UO_2717 (O_2717,N_24700,N_24585);
nand UO_2718 (O_2718,N_24822,N_24894);
nor UO_2719 (O_2719,N_24683,N_24916);
xor UO_2720 (O_2720,N_24943,N_24505);
nor UO_2721 (O_2721,N_24827,N_24886);
xnor UO_2722 (O_2722,N_24898,N_24467);
nor UO_2723 (O_2723,N_24578,N_24407);
xnor UO_2724 (O_2724,N_24418,N_24646);
xor UO_2725 (O_2725,N_24530,N_24830);
or UO_2726 (O_2726,N_24705,N_24471);
or UO_2727 (O_2727,N_24841,N_24393);
nor UO_2728 (O_2728,N_24510,N_24533);
xnor UO_2729 (O_2729,N_24780,N_24766);
and UO_2730 (O_2730,N_24675,N_24535);
nand UO_2731 (O_2731,N_24573,N_24441);
nor UO_2732 (O_2732,N_24523,N_24452);
nand UO_2733 (O_2733,N_24977,N_24794);
xnor UO_2734 (O_2734,N_24911,N_24626);
or UO_2735 (O_2735,N_24744,N_24715);
or UO_2736 (O_2736,N_24821,N_24502);
and UO_2737 (O_2737,N_24720,N_24626);
nand UO_2738 (O_2738,N_24434,N_24939);
nand UO_2739 (O_2739,N_24586,N_24849);
and UO_2740 (O_2740,N_24481,N_24979);
and UO_2741 (O_2741,N_24663,N_24928);
nand UO_2742 (O_2742,N_24949,N_24511);
nand UO_2743 (O_2743,N_24855,N_24493);
nand UO_2744 (O_2744,N_24445,N_24495);
or UO_2745 (O_2745,N_24882,N_24712);
nand UO_2746 (O_2746,N_24849,N_24710);
and UO_2747 (O_2747,N_24640,N_24909);
nand UO_2748 (O_2748,N_24963,N_24979);
or UO_2749 (O_2749,N_24530,N_24724);
and UO_2750 (O_2750,N_24669,N_24973);
and UO_2751 (O_2751,N_24779,N_24499);
and UO_2752 (O_2752,N_24456,N_24792);
xor UO_2753 (O_2753,N_24720,N_24610);
nand UO_2754 (O_2754,N_24411,N_24712);
nand UO_2755 (O_2755,N_24422,N_24804);
and UO_2756 (O_2756,N_24559,N_24797);
xnor UO_2757 (O_2757,N_24658,N_24440);
xnor UO_2758 (O_2758,N_24596,N_24493);
or UO_2759 (O_2759,N_24749,N_24710);
nor UO_2760 (O_2760,N_24474,N_24708);
nand UO_2761 (O_2761,N_24416,N_24693);
and UO_2762 (O_2762,N_24736,N_24600);
xor UO_2763 (O_2763,N_24924,N_24805);
or UO_2764 (O_2764,N_24412,N_24642);
and UO_2765 (O_2765,N_24512,N_24467);
and UO_2766 (O_2766,N_24653,N_24692);
xnor UO_2767 (O_2767,N_24463,N_24675);
nand UO_2768 (O_2768,N_24556,N_24431);
xor UO_2769 (O_2769,N_24461,N_24580);
or UO_2770 (O_2770,N_24429,N_24485);
nand UO_2771 (O_2771,N_24387,N_24420);
xnor UO_2772 (O_2772,N_24447,N_24439);
xor UO_2773 (O_2773,N_24453,N_24841);
nor UO_2774 (O_2774,N_24642,N_24456);
or UO_2775 (O_2775,N_24496,N_24452);
nand UO_2776 (O_2776,N_24798,N_24447);
nand UO_2777 (O_2777,N_24577,N_24416);
nor UO_2778 (O_2778,N_24380,N_24574);
nor UO_2779 (O_2779,N_24434,N_24475);
and UO_2780 (O_2780,N_24863,N_24952);
and UO_2781 (O_2781,N_24738,N_24818);
nand UO_2782 (O_2782,N_24638,N_24547);
nor UO_2783 (O_2783,N_24997,N_24464);
nor UO_2784 (O_2784,N_24562,N_24574);
or UO_2785 (O_2785,N_24469,N_24749);
nor UO_2786 (O_2786,N_24925,N_24475);
nand UO_2787 (O_2787,N_24662,N_24551);
xor UO_2788 (O_2788,N_24568,N_24570);
nand UO_2789 (O_2789,N_24858,N_24448);
or UO_2790 (O_2790,N_24995,N_24873);
or UO_2791 (O_2791,N_24678,N_24464);
nand UO_2792 (O_2792,N_24849,N_24872);
nand UO_2793 (O_2793,N_24910,N_24710);
xor UO_2794 (O_2794,N_24646,N_24996);
xor UO_2795 (O_2795,N_24496,N_24618);
nor UO_2796 (O_2796,N_24398,N_24986);
or UO_2797 (O_2797,N_24609,N_24452);
and UO_2798 (O_2798,N_24458,N_24445);
nand UO_2799 (O_2799,N_24868,N_24880);
and UO_2800 (O_2800,N_24532,N_24453);
nand UO_2801 (O_2801,N_24706,N_24433);
nand UO_2802 (O_2802,N_24509,N_24547);
or UO_2803 (O_2803,N_24561,N_24751);
nand UO_2804 (O_2804,N_24851,N_24383);
nor UO_2805 (O_2805,N_24494,N_24450);
xnor UO_2806 (O_2806,N_24711,N_24509);
xor UO_2807 (O_2807,N_24539,N_24700);
nor UO_2808 (O_2808,N_24770,N_24985);
nand UO_2809 (O_2809,N_24969,N_24820);
nand UO_2810 (O_2810,N_24467,N_24856);
nor UO_2811 (O_2811,N_24791,N_24978);
nand UO_2812 (O_2812,N_24727,N_24763);
or UO_2813 (O_2813,N_24759,N_24531);
or UO_2814 (O_2814,N_24828,N_24579);
nand UO_2815 (O_2815,N_24431,N_24883);
xnor UO_2816 (O_2816,N_24842,N_24782);
xor UO_2817 (O_2817,N_24676,N_24840);
xor UO_2818 (O_2818,N_24621,N_24592);
nand UO_2819 (O_2819,N_24903,N_24932);
nor UO_2820 (O_2820,N_24809,N_24751);
nand UO_2821 (O_2821,N_24951,N_24994);
nand UO_2822 (O_2822,N_24610,N_24817);
xor UO_2823 (O_2823,N_24733,N_24668);
or UO_2824 (O_2824,N_24871,N_24851);
nand UO_2825 (O_2825,N_24439,N_24627);
or UO_2826 (O_2826,N_24477,N_24536);
and UO_2827 (O_2827,N_24706,N_24770);
or UO_2828 (O_2828,N_24689,N_24574);
nor UO_2829 (O_2829,N_24784,N_24499);
or UO_2830 (O_2830,N_24717,N_24376);
xnor UO_2831 (O_2831,N_24505,N_24672);
xor UO_2832 (O_2832,N_24392,N_24728);
nor UO_2833 (O_2833,N_24508,N_24973);
nor UO_2834 (O_2834,N_24956,N_24551);
nor UO_2835 (O_2835,N_24658,N_24637);
nand UO_2836 (O_2836,N_24455,N_24904);
xor UO_2837 (O_2837,N_24386,N_24648);
nand UO_2838 (O_2838,N_24730,N_24390);
or UO_2839 (O_2839,N_24978,N_24969);
nor UO_2840 (O_2840,N_24641,N_24552);
nor UO_2841 (O_2841,N_24402,N_24737);
nand UO_2842 (O_2842,N_24471,N_24696);
and UO_2843 (O_2843,N_24999,N_24822);
or UO_2844 (O_2844,N_24395,N_24831);
xor UO_2845 (O_2845,N_24861,N_24381);
nand UO_2846 (O_2846,N_24487,N_24789);
nand UO_2847 (O_2847,N_24715,N_24842);
and UO_2848 (O_2848,N_24499,N_24875);
nand UO_2849 (O_2849,N_24622,N_24418);
or UO_2850 (O_2850,N_24508,N_24974);
nor UO_2851 (O_2851,N_24868,N_24826);
or UO_2852 (O_2852,N_24477,N_24457);
or UO_2853 (O_2853,N_24891,N_24734);
nor UO_2854 (O_2854,N_24796,N_24823);
and UO_2855 (O_2855,N_24883,N_24960);
nand UO_2856 (O_2856,N_24427,N_24433);
and UO_2857 (O_2857,N_24894,N_24583);
nor UO_2858 (O_2858,N_24849,N_24846);
and UO_2859 (O_2859,N_24626,N_24417);
nand UO_2860 (O_2860,N_24851,N_24874);
nand UO_2861 (O_2861,N_24510,N_24507);
or UO_2862 (O_2862,N_24624,N_24574);
or UO_2863 (O_2863,N_24817,N_24475);
and UO_2864 (O_2864,N_24776,N_24490);
nor UO_2865 (O_2865,N_24631,N_24481);
xnor UO_2866 (O_2866,N_24774,N_24594);
or UO_2867 (O_2867,N_24479,N_24678);
nor UO_2868 (O_2868,N_24695,N_24432);
or UO_2869 (O_2869,N_24948,N_24686);
or UO_2870 (O_2870,N_24452,N_24739);
xnor UO_2871 (O_2871,N_24783,N_24420);
nor UO_2872 (O_2872,N_24542,N_24701);
nand UO_2873 (O_2873,N_24720,N_24400);
or UO_2874 (O_2874,N_24597,N_24754);
or UO_2875 (O_2875,N_24914,N_24894);
or UO_2876 (O_2876,N_24865,N_24403);
nand UO_2877 (O_2877,N_24906,N_24394);
and UO_2878 (O_2878,N_24581,N_24886);
or UO_2879 (O_2879,N_24675,N_24622);
nand UO_2880 (O_2880,N_24670,N_24524);
nand UO_2881 (O_2881,N_24400,N_24760);
and UO_2882 (O_2882,N_24922,N_24729);
nor UO_2883 (O_2883,N_24722,N_24438);
nand UO_2884 (O_2884,N_24926,N_24770);
xnor UO_2885 (O_2885,N_24491,N_24947);
nor UO_2886 (O_2886,N_24579,N_24978);
xnor UO_2887 (O_2887,N_24515,N_24913);
or UO_2888 (O_2888,N_24689,N_24670);
or UO_2889 (O_2889,N_24969,N_24778);
nand UO_2890 (O_2890,N_24823,N_24962);
nand UO_2891 (O_2891,N_24529,N_24448);
xor UO_2892 (O_2892,N_24868,N_24524);
nand UO_2893 (O_2893,N_24597,N_24908);
or UO_2894 (O_2894,N_24553,N_24967);
xor UO_2895 (O_2895,N_24882,N_24473);
nor UO_2896 (O_2896,N_24686,N_24382);
nor UO_2897 (O_2897,N_24442,N_24834);
nand UO_2898 (O_2898,N_24800,N_24408);
or UO_2899 (O_2899,N_24575,N_24817);
xor UO_2900 (O_2900,N_24613,N_24656);
xor UO_2901 (O_2901,N_24423,N_24709);
xnor UO_2902 (O_2902,N_24734,N_24852);
and UO_2903 (O_2903,N_24964,N_24997);
xor UO_2904 (O_2904,N_24764,N_24911);
and UO_2905 (O_2905,N_24688,N_24612);
and UO_2906 (O_2906,N_24998,N_24566);
nor UO_2907 (O_2907,N_24679,N_24545);
and UO_2908 (O_2908,N_24915,N_24576);
xor UO_2909 (O_2909,N_24663,N_24436);
nand UO_2910 (O_2910,N_24988,N_24535);
xnor UO_2911 (O_2911,N_24690,N_24580);
nand UO_2912 (O_2912,N_24986,N_24853);
and UO_2913 (O_2913,N_24896,N_24966);
nand UO_2914 (O_2914,N_24934,N_24644);
xnor UO_2915 (O_2915,N_24960,N_24688);
or UO_2916 (O_2916,N_24727,N_24859);
nand UO_2917 (O_2917,N_24409,N_24746);
xnor UO_2918 (O_2918,N_24934,N_24590);
or UO_2919 (O_2919,N_24486,N_24677);
and UO_2920 (O_2920,N_24761,N_24539);
xor UO_2921 (O_2921,N_24495,N_24783);
nor UO_2922 (O_2922,N_24977,N_24951);
nand UO_2923 (O_2923,N_24777,N_24705);
and UO_2924 (O_2924,N_24712,N_24860);
nor UO_2925 (O_2925,N_24760,N_24962);
nand UO_2926 (O_2926,N_24609,N_24623);
nor UO_2927 (O_2927,N_24382,N_24647);
xnor UO_2928 (O_2928,N_24989,N_24449);
and UO_2929 (O_2929,N_24714,N_24834);
or UO_2930 (O_2930,N_24594,N_24511);
and UO_2931 (O_2931,N_24800,N_24738);
nor UO_2932 (O_2932,N_24882,N_24514);
and UO_2933 (O_2933,N_24444,N_24967);
nor UO_2934 (O_2934,N_24672,N_24917);
xor UO_2935 (O_2935,N_24588,N_24877);
and UO_2936 (O_2936,N_24905,N_24896);
nand UO_2937 (O_2937,N_24692,N_24723);
and UO_2938 (O_2938,N_24438,N_24642);
or UO_2939 (O_2939,N_24913,N_24567);
xnor UO_2940 (O_2940,N_24781,N_24778);
xor UO_2941 (O_2941,N_24921,N_24925);
nor UO_2942 (O_2942,N_24520,N_24608);
xor UO_2943 (O_2943,N_24385,N_24739);
nor UO_2944 (O_2944,N_24625,N_24456);
or UO_2945 (O_2945,N_24937,N_24434);
and UO_2946 (O_2946,N_24669,N_24428);
or UO_2947 (O_2947,N_24451,N_24490);
nor UO_2948 (O_2948,N_24970,N_24573);
xnor UO_2949 (O_2949,N_24646,N_24887);
xor UO_2950 (O_2950,N_24472,N_24989);
and UO_2951 (O_2951,N_24700,N_24893);
nor UO_2952 (O_2952,N_24732,N_24997);
or UO_2953 (O_2953,N_24630,N_24775);
or UO_2954 (O_2954,N_24793,N_24721);
nor UO_2955 (O_2955,N_24443,N_24560);
nand UO_2956 (O_2956,N_24729,N_24946);
nand UO_2957 (O_2957,N_24874,N_24667);
nand UO_2958 (O_2958,N_24438,N_24522);
nand UO_2959 (O_2959,N_24440,N_24604);
xor UO_2960 (O_2960,N_24621,N_24854);
nor UO_2961 (O_2961,N_24888,N_24697);
or UO_2962 (O_2962,N_24869,N_24710);
nor UO_2963 (O_2963,N_24731,N_24789);
nor UO_2964 (O_2964,N_24736,N_24487);
or UO_2965 (O_2965,N_24835,N_24961);
and UO_2966 (O_2966,N_24831,N_24509);
and UO_2967 (O_2967,N_24884,N_24995);
and UO_2968 (O_2968,N_24646,N_24621);
nor UO_2969 (O_2969,N_24969,N_24617);
nand UO_2970 (O_2970,N_24409,N_24488);
nand UO_2971 (O_2971,N_24538,N_24906);
and UO_2972 (O_2972,N_24701,N_24514);
nand UO_2973 (O_2973,N_24706,N_24468);
xor UO_2974 (O_2974,N_24844,N_24599);
xor UO_2975 (O_2975,N_24425,N_24953);
nand UO_2976 (O_2976,N_24831,N_24677);
or UO_2977 (O_2977,N_24693,N_24536);
and UO_2978 (O_2978,N_24663,N_24880);
nor UO_2979 (O_2979,N_24963,N_24639);
nor UO_2980 (O_2980,N_24846,N_24406);
nand UO_2981 (O_2981,N_24539,N_24685);
or UO_2982 (O_2982,N_24581,N_24922);
nand UO_2983 (O_2983,N_24841,N_24837);
or UO_2984 (O_2984,N_24638,N_24471);
nor UO_2985 (O_2985,N_24633,N_24489);
nand UO_2986 (O_2986,N_24657,N_24908);
and UO_2987 (O_2987,N_24692,N_24981);
or UO_2988 (O_2988,N_24618,N_24976);
xnor UO_2989 (O_2989,N_24856,N_24946);
and UO_2990 (O_2990,N_24486,N_24926);
or UO_2991 (O_2991,N_24473,N_24640);
nor UO_2992 (O_2992,N_24474,N_24747);
and UO_2993 (O_2993,N_24972,N_24611);
nand UO_2994 (O_2994,N_24550,N_24618);
nand UO_2995 (O_2995,N_24636,N_24434);
and UO_2996 (O_2996,N_24459,N_24735);
nor UO_2997 (O_2997,N_24797,N_24913);
or UO_2998 (O_2998,N_24811,N_24901);
nand UO_2999 (O_2999,N_24469,N_24851);
endmodule