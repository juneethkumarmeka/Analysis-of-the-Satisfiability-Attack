module basic_750_5000_1000_5_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_380,In_432);
nand U1 (N_1,In_636,In_334);
and U2 (N_2,In_137,In_514);
nand U3 (N_3,In_725,In_675);
nor U4 (N_4,In_720,In_18);
nor U5 (N_5,In_742,In_148);
or U6 (N_6,In_438,In_38);
and U7 (N_7,In_339,In_537);
nor U8 (N_8,In_167,In_723);
or U9 (N_9,In_409,In_541);
xnor U10 (N_10,In_652,In_462);
nor U11 (N_11,In_558,In_143);
nand U12 (N_12,In_121,In_208);
or U13 (N_13,In_543,In_215);
nand U14 (N_14,In_431,In_65);
xor U15 (N_15,In_98,In_175);
nand U16 (N_16,In_707,In_637);
nor U17 (N_17,In_299,In_82);
and U18 (N_18,In_113,In_613);
or U19 (N_19,In_147,In_461);
nand U20 (N_20,In_110,In_269);
nand U21 (N_21,In_151,In_684);
nand U22 (N_22,In_224,In_1);
or U23 (N_23,In_197,In_746);
nor U24 (N_24,In_406,In_150);
nor U25 (N_25,In_72,In_195);
nor U26 (N_26,In_223,In_658);
or U27 (N_27,In_357,In_252);
nand U28 (N_28,In_233,In_459);
nor U29 (N_29,In_39,In_211);
and U30 (N_30,In_539,In_592);
or U31 (N_31,In_122,In_21);
and U32 (N_32,In_32,In_434);
nor U33 (N_33,In_338,In_129);
and U34 (N_34,In_555,In_285);
or U35 (N_35,In_375,In_293);
nor U36 (N_36,In_10,In_739);
nand U37 (N_37,In_286,In_427);
nor U38 (N_38,In_521,In_458);
nor U39 (N_39,In_216,In_593);
nor U40 (N_40,In_672,In_29);
nor U41 (N_41,In_45,In_489);
or U42 (N_42,In_342,In_388);
or U43 (N_43,In_303,In_628);
nand U44 (N_44,In_41,In_439);
nor U45 (N_45,In_727,In_691);
or U46 (N_46,In_378,In_369);
nor U47 (N_47,In_625,In_306);
or U48 (N_48,In_315,In_212);
nor U49 (N_49,In_231,In_565);
nand U50 (N_50,In_271,In_559);
or U51 (N_51,In_57,In_476);
nor U52 (N_52,In_444,In_264);
nand U53 (N_53,In_296,In_107);
nor U54 (N_54,In_411,In_356);
and U55 (N_55,In_160,In_717);
and U56 (N_56,In_103,In_141);
and U57 (N_57,In_446,In_59);
and U58 (N_58,In_397,In_572);
or U59 (N_59,In_133,In_683);
nand U60 (N_60,In_573,In_712);
nand U61 (N_61,In_687,In_347);
nor U62 (N_62,In_101,In_258);
nand U63 (N_63,In_609,In_326);
or U64 (N_64,In_420,In_520);
and U65 (N_65,In_574,In_656);
and U66 (N_66,In_88,In_726);
and U67 (N_67,In_620,In_100);
and U68 (N_68,In_482,In_700);
nand U69 (N_69,In_740,In_49);
nand U70 (N_70,In_177,In_733);
and U71 (N_71,In_582,In_692);
nand U72 (N_72,In_185,In_260);
nor U73 (N_73,In_2,In_423);
nor U74 (N_74,In_545,In_635);
xnor U75 (N_75,In_118,In_19);
nand U76 (N_76,In_703,In_352);
and U77 (N_77,In_256,In_578);
or U78 (N_78,In_71,In_506);
or U79 (N_79,In_11,In_350);
nor U80 (N_80,In_627,In_580);
or U81 (N_81,In_517,In_679);
nor U82 (N_82,In_94,In_77);
nand U83 (N_83,In_157,In_152);
nand U84 (N_84,In_75,In_161);
and U85 (N_85,In_144,In_297);
and U86 (N_86,In_666,In_166);
and U87 (N_87,In_332,In_648);
nand U88 (N_88,In_589,In_393);
nor U89 (N_89,In_435,In_305);
nand U90 (N_90,In_415,In_78);
nor U91 (N_91,In_651,In_382);
nor U92 (N_92,In_486,In_288);
nor U93 (N_93,In_721,In_287);
or U94 (N_94,In_660,In_280);
nand U95 (N_95,In_608,In_669);
nor U96 (N_96,In_0,In_206);
or U97 (N_97,In_340,In_569);
nand U98 (N_98,In_52,In_405);
nand U99 (N_99,In_320,In_642);
xnor U100 (N_100,In_394,In_523);
nor U101 (N_101,In_452,In_467);
or U102 (N_102,In_502,In_630);
nor U103 (N_103,In_54,In_87);
nand U104 (N_104,In_464,In_43);
nor U105 (N_105,In_599,In_64);
nor U106 (N_106,In_79,In_222);
nor U107 (N_107,In_67,In_6);
and U108 (N_108,In_645,In_668);
nor U109 (N_109,In_86,In_90);
nand U110 (N_110,In_585,In_581);
and U111 (N_111,In_304,In_492);
nand U112 (N_112,In_528,In_294);
nor U113 (N_113,In_263,In_734);
and U114 (N_114,In_566,In_243);
nand U115 (N_115,In_300,In_198);
or U116 (N_116,In_190,In_188);
xor U117 (N_117,In_196,In_661);
nor U118 (N_118,In_116,In_327);
nor U119 (N_119,In_261,In_310);
xor U120 (N_120,In_653,In_532);
and U121 (N_121,In_191,In_426);
or U122 (N_122,In_629,In_549);
nor U123 (N_123,In_248,In_500);
nand U124 (N_124,In_50,In_99);
nor U125 (N_125,In_632,In_236);
nor U126 (N_126,In_265,In_722);
nor U127 (N_127,In_448,In_207);
nand U128 (N_128,In_404,In_105);
or U129 (N_129,In_371,In_253);
or U130 (N_130,In_719,In_618);
or U131 (N_131,In_445,In_709);
and U132 (N_132,In_579,In_571);
nor U133 (N_133,In_324,In_372);
nor U134 (N_134,In_173,In_227);
or U135 (N_135,In_384,In_670);
and U136 (N_136,In_267,In_182);
or U137 (N_137,In_655,In_37);
or U138 (N_138,In_540,In_594);
nor U139 (N_139,In_422,In_176);
nor U140 (N_140,In_268,In_363);
nor U141 (N_141,In_346,In_586);
or U142 (N_142,In_205,In_355);
and U143 (N_143,In_368,In_46);
nor U144 (N_144,In_515,In_55);
nand U145 (N_145,In_364,In_5);
nor U146 (N_146,In_536,In_178);
and U147 (N_147,In_659,In_131);
or U148 (N_148,In_12,In_605);
nor U149 (N_149,In_309,In_91);
or U150 (N_150,In_485,In_527);
nor U151 (N_151,In_146,In_60);
or U152 (N_152,In_504,In_123);
and U153 (N_153,In_158,In_447);
xor U154 (N_154,In_272,In_449);
nor U155 (N_155,In_465,In_187);
nor U156 (N_156,In_563,In_76);
nor U157 (N_157,In_495,In_257);
nor U158 (N_158,In_179,In_391);
or U159 (N_159,In_440,In_729);
nand U160 (N_160,In_621,In_240);
or U161 (N_161,In_16,In_525);
and U162 (N_162,In_27,In_155);
and U163 (N_163,In_376,In_387);
or U164 (N_164,In_4,In_136);
or U165 (N_165,In_451,In_557);
nand U166 (N_166,In_612,In_181);
and U167 (N_167,In_481,In_92);
nor U168 (N_168,In_362,In_199);
or U169 (N_169,In_153,In_53);
or U170 (N_170,In_398,In_744);
nand U171 (N_171,In_183,In_622);
nor U172 (N_172,In_576,In_508);
nand U173 (N_173,In_169,In_171);
and U174 (N_174,In_381,In_314);
or U175 (N_175,In_48,In_724);
and U176 (N_176,In_441,In_473);
nor U177 (N_177,In_311,In_681);
nand U178 (N_178,In_9,In_493);
or U179 (N_179,In_511,In_403);
or U180 (N_180,In_61,In_322);
nand U181 (N_181,In_93,In_682);
and U182 (N_182,In_202,In_619);
or U183 (N_183,In_194,In_238);
and U184 (N_184,In_662,In_125);
nor U185 (N_185,In_400,In_436);
and U186 (N_186,In_551,In_336);
nor U187 (N_187,In_385,In_698);
nor U188 (N_188,In_126,In_716);
and U189 (N_189,In_164,In_189);
or U190 (N_190,In_307,In_213);
or U191 (N_191,In_643,In_230);
or U192 (N_192,In_412,In_225);
or U193 (N_193,In_31,In_442);
nor U194 (N_194,In_603,In_533);
xnor U195 (N_195,In_650,In_278);
and U196 (N_196,In_598,In_30);
nand U197 (N_197,In_354,In_289);
nor U198 (N_198,In_453,In_325);
or U199 (N_199,In_301,In_399);
or U200 (N_200,In_313,In_170);
or U201 (N_201,In_298,In_583);
or U202 (N_202,In_702,In_455);
and U203 (N_203,In_497,In_254);
and U204 (N_204,In_713,In_249);
or U205 (N_205,In_550,In_114);
nand U206 (N_206,In_134,In_180);
nor U207 (N_207,In_730,In_737);
or U208 (N_208,In_499,In_657);
and U209 (N_209,In_624,In_244);
nor U210 (N_210,In_51,In_163);
and U211 (N_211,In_84,In_36);
or U212 (N_212,In_358,In_44);
nand U213 (N_213,In_117,In_33);
or U214 (N_214,In_245,In_510);
nand U215 (N_215,In_654,In_247);
and U216 (N_216,In_119,In_17);
or U217 (N_217,In_677,In_7);
or U218 (N_218,In_475,In_359);
nor U219 (N_219,In_132,In_209);
or U220 (N_220,In_561,In_291);
and U221 (N_221,In_673,In_204);
nand U222 (N_222,In_748,In_590);
nor U223 (N_223,In_496,In_688);
or U224 (N_224,In_745,In_604);
nor U225 (N_225,In_425,In_693);
nor U226 (N_226,In_273,In_58);
nor U227 (N_227,In_328,In_477);
and U228 (N_228,In_106,In_646);
nor U229 (N_229,In_102,In_124);
xnor U230 (N_230,In_747,In_705);
nand U231 (N_231,In_414,In_680);
or U232 (N_232,In_331,In_584);
nor U233 (N_233,In_250,In_221);
nor U234 (N_234,In_210,In_468);
nor U235 (N_235,In_239,In_417);
nand U236 (N_236,In_410,In_649);
nand U237 (N_237,In_95,In_139);
or U238 (N_238,In_374,In_483);
or U239 (N_239,In_749,In_591);
or U240 (N_240,In_295,In_567);
nor U241 (N_241,In_353,In_140);
nand U242 (N_242,In_575,In_15);
nand U243 (N_243,In_47,In_149);
or U244 (N_244,In_443,In_373);
nand U245 (N_245,In_63,In_81);
and U246 (N_246,In_469,In_266);
or U247 (N_247,In_111,In_274);
or U248 (N_248,In_42,In_130);
nand U249 (N_249,In_323,In_466);
nand U250 (N_250,In_547,In_68);
nor U251 (N_251,In_664,In_83);
or U252 (N_252,In_456,In_507);
nor U253 (N_253,In_217,In_487);
nand U254 (N_254,In_290,In_647);
and U255 (N_255,In_321,In_142);
nor U256 (N_256,In_743,In_135);
nand U257 (N_257,In_23,In_470);
nor U258 (N_258,In_120,In_715);
nor U259 (N_259,In_214,In_626);
and U260 (N_260,In_513,In_351);
or U261 (N_261,In_524,In_615);
nand U262 (N_262,In_108,In_600);
or U263 (N_263,In_710,In_552);
nand U264 (N_264,In_478,In_348);
nand U265 (N_265,In_366,In_494);
xnor U266 (N_266,In_542,In_562);
and U267 (N_267,In_588,In_73);
nand U268 (N_268,In_704,In_229);
nor U269 (N_269,In_546,In_519);
xnor U270 (N_270,In_556,In_40);
nor U271 (N_271,In_262,In_345);
and U272 (N_272,In_408,In_738);
or U273 (N_273,In_127,In_663);
or U274 (N_274,In_276,In_246);
and U275 (N_275,In_112,In_741);
and U276 (N_276,In_623,In_219);
nor U277 (N_277,In_731,In_365);
nor U278 (N_278,In_292,In_275);
nor U279 (N_279,In_28,In_318);
nand U280 (N_280,In_474,In_450);
nand U281 (N_281,In_644,In_498);
or U282 (N_282,In_428,In_154);
nor U283 (N_283,In_530,In_501);
nand U284 (N_284,In_281,In_595);
and U285 (N_285,In_317,In_472);
nor U286 (N_286,In_568,In_735);
or U287 (N_287,In_14,In_529);
nor U288 (N_288,In_695,In_512);
nor U289 (N_289,In_335,In_341);
nor U290 (N_290,In_544,In_479);
nor U291 (N_291,In_505,In_282);
and U292 (N_292,In_193,In_25);
nor U293 (N_293,In_602,In_418);
nor U294 (N_294,In_437,In_34);
and U295 (N_295,In_711,In_690);
or U296 (N_296,In_138,In_607);
nor U297 (N_297,In_242,In_66);
or U298 (N_298,In_696,In_548);
or U299 (N_299,In_333,In_8);
nand U300 (N_300,In_401,In_611);
nand U301 (N_301,In_172,In_97);
nand U302 (N_302,In_69,In_516);
and U303 (N_303,In_367,In_184);
xnor U304 (N_304,In_699,In_316);
or U305 (N_305,In_728,In_85);
nand U306 (N_306,In_503,In_606);
and U307 (N_307,In_518,In_685);
and U308 (N_308,In_200,In_732);
and U309 (N_309,In_641,In_251);
and U310 (N_310,In_631,In_330);
nor U311 (N_311,In_706,In_471);
nand U312 (N_312,In_255,In_74);
or U313 (N_313,In_667,In_237);
and U314 (N_314,In_676,In_156);
or U315 (N_315,In_203,In_168);
nor U316 (N_316,In_454,In_714);
and U317 (N_317,In_201,In_560);
and U318 (N_318,In_457,In_421);
and U319 (N_319,In_694,In_531);
nor U320 (N_320,In_689,In_174);
nand U321 (N_321,In_597,In_538);
nand U322 (N_322,In_270,In_671);
nand U323 (N_323,In_416,In_226);
or U324 (N_324,In_115,In_159);
nand U325 (N_325,In_617,In_402);
or U326 (N_326,In_277,In_284);
nand U327 (N_327,In_616,In_488);
and U328 (N_328,In_232,In_553);
and U329 (N_329,In_665,In_708);
and U330 (N_330,In_370,In_241);
or U331 (N_331,In_89,In_302);
or U332 (N_332,In_162,In_109);
nor U333 (N_333,In_392,In_22);
and U334 (N_334,In_718,In_308);
and U335 (N_335,In_80,In_70);
nor U336 (N_336,In_377,In_283);
and U337 (N_337,In_395,In_463);
and U338 (N_338,In_736,In_491);
nand U339 (N_339,In_633,In_697);
nand U340 (N_340,In_165,In_526);
or U341 (N_341,In_234,In_56);
or U342 (N_342,In_319,In_379);
nand U343 (N_343,In_62,In_610);
nor U344 (N_344,In_349,In_24);
nor U345 (N_345,In_128,In_35);
nor U346 (N_346,In_433,In_104);
or U347 (N_347,In_343,In_390);
and U348 (N_348,In_361,In_26);
nor U349 (N_349,In_678,In_587);
or U350 (N_350,In_279,In_192);
or U351 (N_351,In_344,In_614);
nor U352 (N_352,In_429,In_490);
and U353 (N_353,In_596,In_430);
or U354 (N_354,In_601,In_235);
nand U355 (N_355,In_228,In_360);
xor U356 (N_356,In_329,In_640);
or U357 (N_357,In_570,In_577);
nand U358 (N_358,In_312,In_383);
and U359 (N_359,In_407,In_674);
nor U360 (N_360,In_535,In_484);
nor U361 (N_361,In_639,In_419);
nor U362 (N_362,In_186,In_460);
nand U363 (N_363,In_424,In_701);
or U364 (N_364,In_509,In_145);
nand U365 (N_365,In_218,In_534);
nor U366 (N_366,In_389,In_638);
nand U367 (N_367,In_96,In_3);
and U368 (N_368,In_13,In_386);
nand U369 (N_369,In_634,In_522);
and U370 (N_370,In_259,In_564);
or U371 (N_371,In_480,In_686);
nand U372 (N_372,In_20,In_337);
or U373 (N_373,In_413,In_396);
and U374 (N_374,In_220,In_554);
or U375 (N_375,In_338,In_248);
or U376 (N_376,In_5,In_356);
and U377 (N_377,In_496,In_621);
nand U378 (N_378,In_331,In_634);
nand U379 (N_379,In_154,In_613);
nand U380 (N_380,In_431,In_378);
or U381 (N_381,In_671,In_626);
or U382 (N_382,In_180,In_521);
nor U383 (N_383,In_354,In_524);
nand U384 (N_384,In_732,In_388);
nand U385 (N_385,In_524,In_461);
nor U386 (N_386,In_74,In_700);
nor U387 (N_387,In_536,In_406);
or U388 (N_388,In_140,In_667);
xor U389 (N_389,In_169,In_257);
nand U390 (N_390,In_68,In_330);
or U391 (N_391,In_219,In_290);
nor U392 (N_392,In_317,In_177);
or U393 (N_393,In_685,In_266);
nor U394 (N_394,In_110,In_300);
nor U395 (N_395,In_506,In_422);
nor U396 (N_396,In_348,In_38);
nor U397 (N_397,In_662,In_413);
and U398 (N_398,In_435,In_216);
or U399 (N_399,In_276,In_144);
or U400 (N_400,In_93,In_16);
or U401 (N_401,In_709,In_594);
nor U402 (N_402,In_407,In_747);
nand U403 (N_403,In_65,In_407);
and U404 (N_404,In_79,In_234);
or U405 (N_405,In_666,In_78);
nor U406 (N_406,In_536,In_653);
nor U407 (N_407,In_705,In_156);
or U408 (N_408,In_332,In_50);
nor U409 (N_409,In_704,In_455);
nor U410 (N_410,In_188,In_218);
or U411 (N_411,In_311,In_260);
nor U412 (N_412,In_180,In_495);
nor U413 (N_413,In_127,In_510);
nor U414 (N_414,In_556,In_610);
nand U415 (N_415,In_208,In_400);
nand U416 (N_416,In_439,In_427);
and U417 (N_417,In_705,In_633);
nand U418 (N_418,In_627,In_576);
or U419 (N_419,In_158,In_457);
nor U420 (N_420,In_546,In_746);
and U421 (N_421,In_599,In_673);
or U422 (N_422,In_11,In_232);
nand U423 (N_423,In_481,In_79);
nand U424 (N_424,In_193,In_252);
and U425 (N_425,In_199,In_673);
or U426 (N_426,In_401,In_711);
nor U427 (N_427,In_742,In_679);
and U428 (N_428,In_215,In_332);
or U429 (N_429,In_677,In_548);
nand U430 (N_430,In_657,In_503);
and U431 (N_431,In_144,In_358);
or U432 (N_432,In_272,In_296);
and U433 (N_433,In_398,In_225);
nor U434 (N_434,In_679,In_51);
nand U435 (N_435,In_726,In_176);
and U436 (N_436,In_444,In_81);
nor U437 (N_437,In_613,In_254);
or U438 (N_438,In_181,In_367);
or U439 (N_439,In_495,In_45);
nand U440 (N_440,In_395,In_131);
and U441 (N_441,In_591,In_511);
or U442 (N_442,In_125,In_391);
and U443 (N_443,In_0,In_42);
and U444 (N_444,In_195,In_344);
nand U445 (N_445,In_194,In_728);
or U446 (N_446,In_343,In_42);
and U447 (N_447,In_126,In_638);
and U448 (N_448,In_186,In_149);
or U449 (N_449,In_221,In_503);
nand U450 (N_450,In_287,In_78);
nor U451 (N_451,In_43,In_364);
and U452 (N_452,In_76,In_629);
or U453 (N_453,In_332,In_79);
or U454 (N_454,In_25,In_598);
or U455 (N_455,In_190,In_299);
nand U456 (N_456,In_73,In_604);
nor U457 (N_457,In_106,In_25);
and U458 (N_458,In_128,In_380);
nor U459 (N_459,In_551,In_480);
nand U460 (N_460,In_401,In_333);
or U461 (N_461,In_686,In_243);
nand U462 (N_462,In_287,In_294);
and U463 (N_463,In_724,In_731);
nand U464 (N_464,In_445,In_379);
nand U465 (N_465,In_462,In_485);
nor U466 (N_466,In_574,In_134);
nand U467 (N_467,In_441,In_95);
nor U468 (N_468,In_34,In_165);
nand U469 (N_469,In_250,In_451);
and U470 (N_470,In_476,In_140);
nor U471 (N_471,In_179,In_61);
nor U472 (N_472,In_273,In_569);
nand U473 (N_473,In_276,In_103);
nor U474 (N_474,In_538,In_383);
nand U475 (N_475,In_98,In_299);
nand U476 (N_476,In_91,In_547);
and U477 (N_477,In_470,In_153);
nand U478 (N_478,In_375,In_585);
and U479 (N_479,In_314,In_547);
nand U480 (N_480,In_25,In_559);
nand U481 (N_481,In_281,In_324);
or U482 (N_482,In_492,In_180);
and U483 (N_483,In_23,In_350);
nand U484 (N_484,In_182,In_30);
nor U485 (N_485,In_551,In_296);
or U486 (N_486,In_224,In_352);
xor U487 (N_487,In_95,In_276);
and U488 (N_488,In_285,In_220);
nor U489 (N_489,In_390,In_649);
and U490 (N_490,In_360,In_192);
and U491 (N_491,In_65,In_728);
or U492 (N_492,In_218,In_315);
and U493 (N_493,In_240,In_511);
and U494 (N_494,In_463,In_94);
and U495 (N_495,In_279,In_289);
nand U496 (N_496,In_664,In_612);
or U497 (N_497,In_66,In_215);
nand U498 (N_498,In_549,In_618);
and U499 (N_499,In_358,In_433);
and U500 (N_500,In_523,In_35);
and U501 (N_501,In_96,In_32);
and U502 (N_502,In_186,In_531);
nor U503 (N_503,In_695,In_261);
nand U504 (N_504,In_738,In_696);
or U505 (N_505,In_641,In_406);
nor U506 (N_506,In_622,In_549);
nand U507 (N_507,In_413,In_357);
or U508 (N_508,In_12,In_622);
nor U509 (N_509,In_600,In_58);
or U510 (N_510,In_708,In_487);
nand U511 (N_511,In_702,In_135);
nor U512 (N_512,In_671,In_262);
nand U513 (N_513,In_493,In_598);
or U514 (N_514,In_156,In_277);
and U515 (N_515,In_36,In_277);
nor U516 (N_516,In_476,In_257);
nand U517 (N_517,In_703,In_346);
nor U518 (N_518,In_313,In_336);
or U519 (N_519,In_150,In_270);
or U520 (N_520,In_292,In_82);
nor U521 (N_521,In_370,In_681);
nor U522 (N_522,In_747,In_156);
or U523 (N_523,In_129,In_287);
nand U524 (N_524,In_286,In_505);
nand U525 (N_525,In_450,In_82);
or U526 (N_526,In_12,In_111);
nand U527 (N_527,In_3,In_305);
nor U528 (N_528,In_213,In_517);
nand U529 (N_529,In_92,In_699);
or U530 (N_530,In_444,In_419);
nor U531 (N_531,In_55,In_34);
and U532 (N_532,In_143,In_505);
or U533 (N_533,In_30,In_84);
or U534 (N_534,In_480,In_568);
nand U535 (N_535,In_310,In_452);
nor U536 (N_536,In_109,In_158);
or U537 (N_537,In_428,In_114);
or U538 (N_538,In_363,In_630);
and U539 (N_539,In_384,In_39);
or U540 (N_540,In_591,In_518);
and U541 (N_541,In_151,In_254);
nor U542 (N_542,In_445,In_516);
xnor U543 (N_543,In_402,In_533);
or U544 (N_544,In_423,In_688);
nor U545 (N_545,In_359,In_599);
and U546 (N_546,In_392,In_401);
nand U547 (N_547,In_105,In_727);
and U548 (N_548,In_124,In_161);
or U549 (N_549,In_534,In_671);
nand U550 (N_550,In_273,In_703);
nand U551 (N_551,In_709,In_11);
nand U552 (N_552,In_274,In_660);
and U553 (N_553,In_67,In_635);
nand U554 (N_554,In_240,In_196);
nand U555 (N_555,In_138,In_617);
or U556 (N_556,In_223,In_165);
nand U557 (N_557,In_389,In_10);
nor U558 (N_558,In_564,In_406);
or U559 (N_559,In_466,In_336);
nand U560 (N_560,In_204,In_697);
nand U561 (N_561,In_567,In_504);
nor U562 (N_562,In_186,In_570);
and U563 (N_563,In_113,In_594);
nand U564 (N_564,In_569,In_98);
and U565 (N_565,In_265,In_157);
or U566 (N_566,In_239,In_126);
or U567 (N_567,In_3,In_399);
and U568 (N_568,In_438,In_277);
and U569 (N_569,In_430,In_137);
nand U570 (N_570,In_743,In_29);
or U571 (N_571,In_492,In_43);
nor U572 (N_572,In_44,In_262);
and U573 (N_573,In_356,In_145);
nor U574 (N_574,In_691,In_266);
and U575 (N_575,In_728,In_102);
or U576 (N_576,In_444,In_87);
nand U577 (N_577,In_338,In_451);
and U578 (N_578,In_555,In_109);
nand U579 (N_579,In_106,In_183);
and U580 (N_580,In_428,In_424);
nor U581 (N_581,In_190,In_167);
and U582 (N_582,In_439,In_616);
and U583 (N_583,In_560,In_433);
nand U584 (N_584,In_689,In_459);
nand U585 (N_585,In_547,In_495);
and U586 (N_586,In_423,In_84);
nand U587 (N_587,In_744,In_320);
and U588 (N_588,In_176,In_623);
nand U589 (N_589,In_209,In_319);
nor U590 (N_590,In_318,In_592);
nor U591 (N_591,In_87,In_279);
nand U592 (N_592,In_253,In_394);
and U593 (N_593,In_310,In_531);
and U594 (N_594,In_565,In_497);
nor U595 (N_595,In_346,In_24);
and U596 (N_596,In_193,In_605);
nand U597 (N_597,In_737,In_100);
nand U598 (N_598,In_62,In_411);
or U599 (N_599,In_283,In_311);
or U600 (N_600,In_163,In_423);
nand U601 (N_601,In_445,In_573);
and U602 (N_602,In_173,In_613);
or U603 (N_603,In_271,In_36);
nor U604 (N_604,In_609,In_563);
nor U605 (N_605,In_634,In_231);
or U606 (N_606,In_661,In_107);
nand U607 (N_607,In_530,In_678);
or U608 (N_608,In_586,In_373);
or U609 (N_609,In_492,In_132);
nor U610 (N_610,In_396,In_549);
and U611 (N_611,In_158,In_21);
or U612 (N_612,In_423,In_578);
nand U613 (N_613,In_258,In_712);
and U614 (N_614,In_737,In_649);
or U615 (N_615,In_183,In_40);
and U616 (N_616,In_270,In_507);
nor U617 (N_617,In_94,In_536);
nand U618 (N_618,In_233,In_208);
nor U619 (N_619,In_529,In_298);
and U620 (N_620,In_730,In_123);
nor U621 (N_621,In_714,In_116);
nand U622 (N_622,In_410,In_173);
and U623 (N_623,In_28,In_648);
or U624 (N_624,In_50,In_104);
or U625 (N_625,In_482,In_241);
and U626 (N_626,In_549,In_742);
nor U627 (N_627,In_486,In_680);
nand U628 (N_628,In_284,In_202);
nand U629 (N_629,In_170,In_402);
and U630 (N_630,In_416,In_602);
or U631 (N_631,In_633,In_193);
nand U632 (N_632,In_540,In_574);
nand U633 (N_633,In_411,In_338);
and U634 (N_634,In_667,In_619);
nand U635 (N_635,In_466,In_607);
or U636 (N_636,In_336,In_556);
nand U637 (N_637,In_231,In_141);
and U638 (N_638,In_544,In_579);
or U639 (N_639,In_509,In_364);
nor U640 (N_640,In_622,In_366);
and U641 (N_641,In_501,In_546);
nor U642 (N_642,In_45,In_233);
or U643 (N_643,In_718,In_464);
or U644 (N_644,In_714,In_14);
nand U645 (N_645,In_47,In_414);
nor U646 (N_646,In_615,In_45);
or U647 (N_647,In_1,In_674);
and U648 (N_648,In_665,In_247);
and U649 (N_649,In_418,In_166);
and U650 (N_650,In_378,In_552);
or U651 (N_651,In_178,In_287);
nand U652 (N_652,In_732,In_374);
and U653 (N_653,In_231,In_137);
nand U654 (N_654,In_568,In_313);
or U655 (N_655,In_125,In_367);
or U656 (N_656,In_525,In_286);
and U657 (N_657,In_254,In_198);
nor U658 (N_658,In_89,In_361);
nor U659 (N_659,In_370,In_492);
and U660 (N_660,In_391,In_138);
nand U661 (N_661,In_339,In_596);
nor U662 (N_662,In_145,In_667);
nor U663 (N_663,In_631,In_336);
or U664 (N_664,In_34,In_483);
nand U665 (N_665,In_607,In_659);
nand U666 (N_666,In_234,In_80);
or U667 (N_667,In_655,In_555);
nand U668 (N_668,In_563,In_657);
or U669 (N_669,In_153,In_565);
or U670 (N_670,In_1,In_237);
nor U671 (N_671,In_214,In_228);
nor U672 (N_672,In_522,In_83);
or U673 (N_673,In_287,In_273);
or U674 (N_674,In_600,In_597);
nor U675 (N_675,In_506,In_135);
nor U676 (N_676,In_100,In_691);
and U677 (N_677,In_277,In_419);
nor U678 (N_678,In_126,In_700);
and U679 (N_679,In_468,In_29);
nand U680 (N_680,In_390,In_661);
and U681 (N_681,In_646,In_266);
or U682 (N_682,In_164,In_294);
nand U683 (N_683,In_569,In_87);
or U684 (N_684,In_56,In_295);
nor U685 (N_685,In_623,In_327);
nand U686 (N_686,In_380,In_663);
nand U687 (N_687,In_222,In_443);
nor U688 (N_688,In_189,In_96);
nor U689 (N_689,In_477,In_72);
or U690 (N_690,In_208,In_56);
nor U691 (N_691,In_212,In_382);
nand U692 (N_692,In_637,In_212);
nor U693 (N_693,In_243,In_188);
nor U694 (N_694,In_605,In_273);
nand U695 (N_695,In_317,In_257);
and U696 (N_696,In_645,In_64);
and U697 (N_697,In_413,In_120);
or U698 (N_698,In_227,In_564);
or U699 (N_699,In_561,In_20);
or U700 (N_700,In_590,In_458);
nand U701 (N_701,In_279,In_202);
or U702 (N_702,In_711,In_388);
nand U703 (N_703,In_708,In_53);
nand U704 (N_704,In_519,In_115);
and U705 (N_705,In_600,In_2);
and U706 (N_706,In_368,In_335);
or U707 (N_707,In_35,In_14);
or U708 (N_708,In_627,In_391);
or U709 (N_709,In_185,In_557);
and U710 (N_710,In_406,In_439);
and U711 (N_711,In_719,In_668);
xnor U712 (N_712,In_8,In_682);
nor U713 (N_713,In_297,In_585);
and U714 (N_714,In_464,In_580);
or U715 (N_715,In_429,In_307);
and U716 (N_716,In_502,In_280);
nand U717 (N_717,In_376,In_346);
or U718 (N_718,In_589,In_555);
nand U719 (N_719,In_271,In_45);
nor U720 (N_720,In_235,In_553);
or U721 (N_721,In_658,In_717);
or U722 (N_722,In_526,In_204);
nor U723 (N_723,In_306,In_14);
or U724 (N_724,In_640,In_176);
nor U725 (N_725,In_715,In_722);
and U726 (N_726,In_256,In_432);
and U727 (N_727,In_673,In_565);
nand U728 (N_728,In_167,In_142);
and U729 (N_729,In_250,In_91);
and U730 (N_730,In_259,In_602);
nand U731 (N_731,In_50,In_87);
or U732 (N_732,In_418,In_191);
nand U733 (N_733,In_499,In_737);
or U734 (N_734,In_31,In_402);
and U735 (N_735,In_424,In_442);
nand U736 (N_736,In_174,In_337);
nor U737 (N_737,In_672,In_1);
and U738 (N_738,In_380,In_463);
nand U739 (N_739,In_612,In_538);
nand U740 (N_740,In_451,In_324);
or U741 (N_741,In_80,In_713);
or U742 (N_742,In_116,In_646);
nor U743 (N_743,In_443,In_461);
or U744 (N_744,In_67,In_91);
nor U745 (N_745,In_48,In_470);
or U746 (N_746,In_211,In_99);
or U747 (N_747,In_599,In_608);
nor U748 (N_748,In_332,In_375);
or U749 (N_749,In_69,In_329);
nor U750 (N_750,In_29,In_243);
and U751 (N_751,In_298,In_271);
and U752 (N_752,In_723,In_479);
nor U753 (N_753,In_114,In_398);
or U754 (N_754,In_226,In_615);
nand U755 (N_755,In_744,In_90);
nor U756 (N_756,In_712,In_429);
or U757 (N_757,In_356,In_570);
nand U758 (N_758,In_85,In_601);
or U759 (N_759,In_656,In_702);
and U760 (N_760,In_730,In_183);
nor U761 (N_761,In_577,In_544);
nor U762 (N_762,In_254,In_73);
and U763 (N_763,In_635,In_219);
or U764 (N_764,In_419,In_332);
or U765 (N_765,In_273,In_533);
and U766 (N_766,In_660,In_461);
or U767 (N_767,In_310,In_184);
nor U768 (N_768,In_50,In_19);
and U769 (N_769,In_185,In_165);
nand U770 (N_770,In_150,In_658);
or U771 (N_771,In_469,In_620);
nand U772 (N_772,In_525,In_373);
and U773 (N_773,In_743,In_170);
nand U774 (N_774,In_446,In_517);
nand U775 (N_775,In_120,In_231);
or U776 (N_776,In_366,In_54);
or U777 (N_777,In_571,In_544);
nor U778 (N_778,In_537,In_649);
and U779 (N_779,In_361,In_701);
and U780 (N_780,In_690,In_304);
nand U781 (N_781,In_383,In_451);
nand U782 (N_782,In_606,In_406);
nand U783 (N_783,In_251,In_212);
or U784 (N_784,In_20,In_681);
or U785 (N_785,In_725,In_683);
and U786 (N_786,In_59,In_395);
nand U787 (N_787,In_111,In_333);
and U788 (N_788,In_172,In_664);
nand U789 (N_789,In_387,In_415);
or U790 (N_790,In_622,In_406);
nand U791 (N_791,In_565,In_42);
or U792 (N_792,In_405,In_552);
nand U793 (N_793,In_352,In_493);
and U794 (N_794,In_148,In_224);
nor U795 (N_795,In_479,In_224);
or U796 (N_796,In_314,In_354);
nand U797 (N_797,In_216,In_699);
nor U798 (N_798,In_680,In_547);
nand U799 (N_799,In_178,In_334);
or U800 (N_800,In_708,In_125);
nand U801 (N_801,In_451,In_727);
or U802 (N_802,In_204,In_212);
nor U803 (N_803,In_289,In_262);
or U804 (N_804,In_337,In_282);
nor U805 (N_805,In_160,In_657);
and U806 (N_806,In_566,In_739);
and U807 (N_807,In_274,In_732);
nor U808 (N_808,In_513,In_704);
or U809 (N_809,In_569,In_109);
or U810 (N_810,In_380,In_14);
and U811 (N_811,In_176,In_530);
nor U812 (N_812,In_391,In_131);
or U813 (N_813,In_486,In_655);
and U814 (N_814,In_476,In_567);
nand U815 (N_815,In_255,In_685);
xnor U816 (N_816,In_550,In_207);
nor U817 (N_817,In_435,In_264);
or U818 (N_818,In_550,In_450);
xor U819 (N_819,In_30,In_340);
nor U820 (N_820,In_122,In_69);
and U821 (N_821,In_339,In_19);
or U822 (N_822,In_173,In_71);
nor U823 (N_823,In_638,In_627);
and U824 (N_824,In_506,In_538);
or U825 (N_825,In_127,In_71);
or U826 (N_826,In_273,In_409);
and U827 (N_827,In_429,In_513);
nor U828 (N_828,In_428,In_483);
or U829 (N_829,In_702,In_741);
and U830 (N_830,In_558,In_429);
or U831 (N_831,In_108,In_123);
and U832 (N_832,In_415,In_182);
or U833 (N_833,In_408,In_348);
and U834 (N_834,In_200,In_94);
or U835 (N_835,In_602,In_244);
nand U836 (N_836,In_258,In_575);
or U837 (N_837,In_169,In_456);
nor U838 (N_838,In_344,In_442);
or U839 (N_839,In_452,In_463);
or U840 (N_840,In_709,In_649);
nor U841 (N_841,In_337,In_611);
and U842 (N_842,In_30,In_603);
and U843 (N_843,In_682,In_301);
and U844 (N_844,In_584,In_439);
nor U845 (N_845,In_167,In_246);
and U846 (N_846,In_440,In_132);
nand U847 (N_847,In_137,In_571);
nor U848 (N_848,In_592,In_551);
or U849 (N_849,In_339,In_676);
or U850 (N_850,In_158,In_557);
nor U851 (N_851,In_379,In_638);
or U852 (N_852,In_736,In_671);
and U853 (N_853,In_385,In_428);
and U854 (N_854,In_672,In_653);
nand U855 (N_855,In_740,In_444);
nor U856 (N_856,In_141,In_41);
nor U857 (N_857,In_499,In_183);
or U858 (N_858,In_37,In_248);
and U859 (N_859,In_683,In_169);
or U860 (N_860,In_615,In_527);
nor U861 (N_861,In_275,In_204);
or U862 (N_862,In_168,In_273);
nand U863 (N_863,In_290,In_257);
nor U864 (N_864,In_474,In_257);
nand U865 (N_865,In_435,In_669);
or U866 (N_866,In_739,In_465);
nor U867 (N_867,In_113,In_405);
or U868 (N_868,In_138,In_433);
nor U869 (N_869,In_466,In_290);
or U870 (N_870,In_148,In_59);
or U871 (N_871,In_660,In_166);
or U872 (N_872,In_609,In_505);
nand U873 (N_873,In_527,In_67);
and U874 (N_874,In_668,In_599);
or U875 (N_875,In_583,In_669);
nor U876 (N_876,In_695,In_223);
nor U877 (N_877,In_660,In_581);
nor U878 (N_878,In_610,In_525);
nor U879 (N_879,In_122,In_96);
and U880 (N_880,In_83,In_706);
nand U881 (N_881,In_734,In_405);
nor U882 (N_882,In_273,In_125);
and U883 (N_883,In_315,In_717);
or U884 (N_884,In_473,In_175);
nand U885 (N_885,In_155,In_522);
and U886 (N_886,In_176,In_418);
xor U887 (N_887,In_539,In_226);
nand U888 (N_888,In_190,In_746);
and U889 (N_889,In_726,In_560);
nand U890 (N_890,In_536,In_531);
nor U891 (N_891,In_661,In_697);
or U892 (N_892,In_79,In_544);
and U893 (N_893,In_491,In_1);
or U894 (N_894,In_160,In_378);
nor U895 (N_895,In_724,In_271);
nor U896 (N_896,In_40,In_58);
and U897 (N_897,In_271,In_281);
nor U898 (N_898,In_374,In_209);
nand U899 (N_899,In_239,In_482);
and U900 (N_900,In_403,In_349);
xor U901 (N_901,In_17,In_584);
and U902 (N_902,In_495,In_76);
nor U903 (N_903,In_421,In_141);
nor U904 (N_904,In_141,In_187);
nand U905 (N_905,In_333,In_423);
or U906 (N_906,In_72,In_724);
and U907 (N_907,In_109,In_718);
nand U908 (N_908,In_11,In_100);
nor U909 (N_909,In_240,In_670);
or U910 (N_910,In_303,In_275);
and U911 (N_911,In_54,In_276);
or U912 (N_912,In_706,In_288);
nor U913 (N_913,In_174,In_519);
nor U914 (N_914,In_350,In_453);
or U915 (N_915,In_401,In_146);
nand U916 (N_916,In_632,In_687);
or U917 (N_917,In_290,In_33);
or U918 (N_918,In_506,In_730);
or U919 (N_919,In_350,In_94);
and U920 (N_920,In_681,In_472);
and U921 (N_921,In_711,In_623);
nand U922 (N_922,In_370,In_334);
nor U923 (N_923,In_662,In_17);
nor U924 (N_924,In_588,In_84);
nand U925 (N_925,In_313,In_594);
and U926 (N_926,In_638,In_667);
nor U927 (N_927,In_203,In_378);
and U928 (N_928,In_557,In_462);
nor U929 (N_929,In_419,In_126);
xnor U930 (N_930,In_269,In_589);
and U931 (N_931,In_192,In_257);
or U932 (N_932,In_469,In_734);
nor U933 (N_933,In_213,In_296);
nor U934 (N_934,In_470,In_715);
and U935 (N_935,In_109,In_52);
nand U936 (N_936,In_243,In_540);
and U937 (N_937,In_293,In_9);
nor U938 (N_938,In_353,In_522);
and U939 (N_939,In_559,In_631);
nor U940 (N_940,In_121,In_53);
and U941 (N_941,In_249,In_412);
or U942 (N_942,In_414,In_251);
or U943 (N_943,In_533,In_124);
or U944 (N_944,In_66,In_410);
nor U945 (N_945,In_692,In_98);
and U946 (N_946,In_304,In_524);
and U947 (N_947,In_179,In_347);
and U948 (N_948,In_469,In_387);
nor U949 (N_949,In_642,In_567);
or U950 (N_950,In_168,In_15);
and U951 (N_951,In_670,In_125);
or U952 (N_952,In_377,In_430);
or U953 (N_953,In_54,In_323);
or U954 (N_954,In_499,In_605);
nor U955 (N_955,In_173,In_680);
and U956 (N_956,In_540,In_646);
nand U957 (N_957,In_195,In_523);
nor U958 (N_958,In_1,In_675);
and U959 (N_959,In_128,In_738);
or U960 (N_960,In_139,In_617);
nand U961 (N_961,In_258,In_639);
and U962 (N_962,In_669,In_568);
and U963 (N_963,In_89,In_648);
nor U964 (N_964,In_465,In_204);
and U965 (N_965,In_391,In_499);
and U966 (N_966,In_121,In_542);
nand U967 (N_967,In_430,In_586);
nand U968 (N_968,In_629,In_153);
nor U969 (N_969,In_136,In_206);
nand U970 (N_970,In_670,In_177);
nand U971 (N_971,In_74,In_602);
nand U972 (N_972,In_638,In_660);
or U973 (N_973,In_552,In_588);
and U974 (N_974,In_51,In_370);
nor U975 (N_975,In_590,In_495);
nor U976 (N_976,In_444,In_154);
nand U977 (N_977,In_584,In_236);
nand U978 (N_978,In_565,In_184);
and U979 (N_979,In_190,In_367);
nor U980 (N_980,In_51,In_560);
and U981 (N_981,In_128,In_463);
nor U982 (N_982,In_385,In_616);
or U983 (N_983,In_408,In_557);
or U984 (N_984,In_656,In_705);
and U985 (N_985,In_65,In_107);
or U986 (N_986,In_176,In_735);
nand U987 (N_987,In_105,In_154);
or U988 (N_988,In_484,In_214);
and U989 (N_989,In_293,In_312);
nand U990 (N_990,In_367,In_692);
nand U991 (N_991,In_315,In_428);
nor U992 (N_992,In_511,In_157);
or U993 (N_993,In_523,In_412);
nand U994 (N_994,In_92,In_30);
nor U995 (N_995,In_86,In_121);
and U996 (N_996,In_557,In_149);
or U997 (N_997,In_641,In_644);
or U998 (N_998,In_94,In_367);
nor U999 (N_999,In_575,In_712);
nand U1000 (N_1000,N_921,N_205);
nor U1001 (N_1001,N_407,N_124);
nor U1002 (N_1002,N_94,N_633);
and U1003 (N_1003,N_43,N_965);
and U1004 (N_1004,N_811,N_917);
nor U1005 (N_1005,N_226,N_121);
and U1006 (N_1006,N_31,N_68);
and U1007 (N_1007,N_989,N_148);
nor U1008 (N_1008,N_256,N_618);
nor U1009 (N_1009,N_319,N_351);
nand U1010 (N_1010,N_600,N_398);
and U1011 (N_1011,N_262,N_301);
nand U1012 (N_1012,N_732,N_76);
nor U1013 (N_1013,N_418,N_563);
nand U1014 (N_1014,N_964,N_945);
nor U1015 (N_1015,N_234,N_362);
nor U1016 (N_1016,N_267,N_943);
nor U1017 (N_1017,N_796,N_413);
nand U1018 (N_1018,N_966,N_665);
or U1019 (N_1019,N_602,N_61);
xor U1020 (N_1020,N_603,N_706);
or U1021 (N_1021,N_955,N_38);
nand U1022 (N_1022,N_176,N_909);
or U1023 (N_1023,N_74,N_0);
nand U1024 (N_1024,N_568,N_961);
and U1025 (N_1025,N_192,N_860);
nor U1026 (N_1026,N_388,N_824);
nor U1027 (N_1027,N_528,N_952);
nand U1028 (N_1028,N_367,N_577);
and U1029 (N_1029,N_631,N_999);
and U1030 (N_1030,N_66,N_988);
nand U1031 (N_1031,N_346,N_873);
and U1032 (N_1032,N_116,N_165);
nor U1033 (N_1033,N_73,N_459);
or U1034 (N_1034,N_555,N_562);
nor U1035 (N_1035,N_167,N_553);
nand U1036 (N_1036,N_39,N_72);
nand U1037 (N_1037,N_708,N_455);
or U1038 (N_1038,N_545,N_894);
nand U1039 (N_1039,N_549,N_380);
nor U1040 (N_1040,N_419,N_431);
or U1041 (N_1041,N_463,N_172);
or U1042 (N_1042,N_721,N_100);
nor U1043 (N_1043,N_173,N_643);
or U1044 (N_1044,N_120,N_79);
nor U1045 (N_1045,N_668,N_793);
and U1046 (N_1046,N_350,N_349);
or U1047 (N_1047,N_402,N_26);
nand U1048 (N_1048,N_792,N_742);
nand U1049 (N_1049,N_330,N_804);
nor U1050 (N_1050,N_953,N_834);
nand U1051 (N_1051,N_64,N_881);
nand U1052 (N_1052,N_758,N_470);
nand U1053 (N_1053,N_456,N_644);
nand U1054 (N_1054,N_838,N_490);
nand U1055 (N_1055,N_161,N_839);
or U1056 (N_1056,N_198,N_133);
nor U1057 (N_1057,N_483,N_233);
and U1058 (N_1058,N_168,N_283);
or U1059 (N_1059,N_272,N_412);
and U1060 (N_1060,N_71,N_523);
nand U1061 (N_1061,N_381,N_669);
or U1062 (N_1062,N_69,N_693);
nand U1063 (N_1063,N_18,N_847);
nand U1064 (N_1064,N_199,N_481);
nor U1065 (N_1065,N_104,N_806);
nand U1066 (N_1066,N_931,N_960);
or U1067 (N_1067,N_296,N_281);
nand U1068 (N_1068,N_58,N_162);
and U1069 (N_1069,N_813,N_322);
or U1070 (N_1070,N_801,N_780);
nand U1071 (N_1071,N_674,N_489);
nor U1072 (N_1072,N_971,N_348);
or U1073 (N_1073,N_342,N_580);
nor U1074 (N_1074,N_652,N_241);
or U1075 (N_1075,N_33,N_190);
nand U1076 (N_1076,N_962,N_185);
nand U1077 (N_1077,N_186,N_50);
and U1078 (N_1078,N_289,N_940);
or U1079 (N_1079,N_635,N_27);
nor U1080 (N_1080,N_710,N_898);
nor U1081 (N_1081,N_376,N_313);
and U1082 (N_1082,N_62,N_550);
nand U1083 (N_1083,N_731,N_95);
nand U1084 (N_1084,N_129,N_439);
and U1085 (N_1085,N_959,N_88);
nor U1086 (N_1086,N_585,N_466);
nand U1087 (N_1087,N_410,N_458);
nand U1088 (N_1088,N_273,N_210);
nor U1089 (N_1089,N_612,N_164);
nand U1090 (N_1090,N_111,N_401);
nor U1091 (N_1091,N_519,N_253);
and U1092 (N_1092,N_609,N_878);
nor U1093 (N_1093,N_559,N_451);
nor U1094 (N_1094,N_540,N_408);
or U1095 (N_1095,N_872,N_913);
and U1096 (N_1096,N_981,N_740);
nor U1097 (N_1097,N_464,N_448);
and U1098 (N_1098,N_462,N_25);
or U1099 (N_1099,N_151,N_125);
or U1100 (N_1100,N_781,N_227);
nor U1101 (N_1101,N_251,N_903);
or U1102 (N_1102,N_696,N_181);
or U1103 (N_1103,N_394,N_369);
nand U1104 (N_1104,N_911,N_799);
and U1105 (N_1105,N_853,N_440);
xor U1106 (N_1106,N_591,N_189);
and U1107 (N_1107,N_773,N_35);
nand U1108 (N_1108,N_86,N_195);
and U1109 (N_1109,N_787,N_307);
and U1110 (N_1110,N_744,N_219);
or U1111 (N_1111,N_373,N_904);
nand U1112 (N_1112,N_311,N_75);
nor U1113 (N_1113,N_356,N_521);
nor U1114 (N_1114,N_237,N_637);
nor U1115 (N_1115,N_496,N_321);
nand U1116 (N_1116,N_686,N_768);
nand U1117 (N_1117,N_541,N_77);
and U1118 (N_1118,N_323,N_374);
and U1119 (N_1119,N_471,N_247);
nand U1120 (N_1120,N_386,N_264);
nand U1121 (N_1121,N_250,N_750);
nor U1122 (N_1122,N_209,N_814);
or U1123 (N_1123,N_715,N_359);
or U1124 (N_1124,N_868,N_856);
or U1125 (N_1125,N_187,N_12);
and U1126 (N_1126,N_888,N_132);
and U1127 (N_1127,N_8,N_701);
nor U1128 (N_1128,N_970,N_239);
nand U1129 (N_1129,N_926,N_942);
nor U1130 (N_1130,N_968,N_302);
or U1131 (N_1131,N_820,N_547);
nand U1132 (N_1132,N_685,N_554);
or U1133 (N_1133,N_285,N_223);
and U1134 (N_1134,N_835,N_918);
and U1135 (N_1135,N_501,N_784);
and U1136 (N_1136,N_821,N_557);
nand U1137 (N_1137,N_759,N_163);
nand U1138 (N_1138,N_919,N_973);
or U1139 (N_1139,N_716,N_535);
nor U1140 (N_1140,N_42,N_67);
and U1141 (N_1141,N_733,N_22);
nand U1142 (N_1142,N_436,N_276);
nor U1143 (N_1143,N_864,N_235);
nor U1144 (N_1144,N_150,N_421);
or U1145 (N_1145,N_294,N_836);
nor U1146 (N_1146,N_308,N_145);
or U1147 (N_1147,N_995,N_135);
nand U1148 (N_1148,N_101,N_450);
or U1149 (N_1149,N_475,N_513);
nor U1150 (N_1150,N_983,N_975);
or U1151 (N_1151,N_128,N_984);
xor U1152 (N_1152,N_2,N_404);
nand U1153 (N_1153,N_850,N_4);
nor U1154 (N_1154,N_682,N_880);
nand U1155 (N_1155,N_867,N_400);
nor U1156 (N_1156,N_762,N_772);
nand U1157 (N_1157,N_560,N_632);
nor U1158 (N_1158,N_152,N_149);
nor U1159 (N_1159,N_170,N_790);
nand U1160 (N_1160,N_977,N_106);
nand U1161 (N_1161,N_608,N_240);
and U1162 (N_1162,N_108,N_17);
nand U1163 (N_1163,N_117,N_309);
nor U1164 (N_1164,N_6,N_429);
nand U1165 (N_1165,N_218,N_217);
and U1166 (N_1166,N_833,N_862);
and U1167 (N_1167,N_390,N_510);
nor U1168 (N_1168,N_681,N_211);
nand U1169 (N_1169,N_684,N_908);
xnor U1170 (N_1170,N_957,N_927);
nor U1171 (N_1171,N_582,N_902);
nand U1172 (N_1172,N_675,N_905);
nand U1173 (N_1173,N_461,N_761);
and U1174 (N_1174,N_654,N_409);
nor U1175 (N_1175,N_244,N_507);
nand U1176 (N_1176,N_288,N_907);
and U1177 (N_1177,N_385,N_756);
nand U1178 (N_1178,N_131,N_280);
or U1179 (N_1179,N_20,N_432);
nor U1180 (N_1180,N_819,N_874);
nor U1181 (N_1181,N_855,N_454);
nor U1182 (N_1182,N_59,N_147);
or U1183 (N_1183,N_651,N_538);
or U1184 (N_1184,N_822,N_341);
nor U1185 (N_1185,N_208,N_816);
xnor U1186 (N_1186,N_594,N_869);
and U1187 (N_1187,N_883,N_937);
or U1188 (N_1188,N_785,N_689);
nor U1189 (N_1189,N_987,N_96);
and U1190 (N_1190,N_84,N_664);
nor U1191 (N_1191,N_656,N_809);
or U1192 (N_1192,N_316,N_137);
or U1193 (N_1193,N_976,N_265);
nand U1194 (N_1194,N_468,N_641);
nand U1195 (N_1195,N_727,N_37);
and U1196 (N_1196,N_194,N_314);
nand U1197 (N_1197,N_561,N_719);
or U1198 (N_1198,N_741,N_534);
nand U1199 (N_1199,N_224,N_658);
or U1200 (N_1200,N_391,N_425);
or U1201 (N_1201,N_415,N_551);
or U1202 (N_1202,N_938,N_246);
and U1203 (N_1203,N_5,N_889);
or U1204 (N_1204,N_846,N_766);
nand U1205 (N_1205,N_406,N_574);
and U1206 (N_1206,N_599,N_21);
or U1207 (N_1207,N_478,N_845);
and U1208 (N_1208,N_191,N_969);
or U1209 (N_1209,N_579,N_118);
and U1210 (N_1210,N_228,N_980);
nor U1211 (N_1211,N_718,N_422);
nor U1212 (N_1212,N_520,N_500);
and U1213 (N_1213,N_530,N_688);
or U1214 (N_1214,N_449,N_692);
or U1215 (N_1215,N_653,N_986);
and U1216 (N_1216,N_922,N_666);
nand U1217 (N_1217,N_63,N_403);
or U1218 (N_1218,N_760,N_213);
and U1219 (N_1219,N_769,N_357);
and U1220 (N_1220,N_60,N_434);
nor U1221 (N_1221,N_82,N_569);
nor U1222 (N_1222,N_858,N_645);
nand U1223 (N_1223,N_748,N_606);
and U1224 (N_1224,N_315,N_243);
nor U1225 (N_1225,N_140,N_212);
or U1226 (N_1226,N_155,N_502);
nand U1227 (N_1227,N_144,N_472);
or U1228 (N_1228,N_998,N_427);
and U1229 (N_1229,N_730,N_438);
nand U1230 (N_1230,N_370,N_640);
nor U1231 (N_1231,N_638,N_372);
nor U1232 (N_1232,N_932,N_915);
or U1233 (N_1233,N_395,N_642);
and U1234 (N_1234,N_363,N_737);
xor U1235 (N_1235,N_136,N_593);
nand U1236 (N_1236,N_126,N_32);
nor U1237 (N_1237,N_586,N_329);
or U1238 (N_1238,N_486,N_798);
and U1239 (N_1239,N_476,N_179);
nor U1240 (N_1240,N_484,N_544);
and U1241 (N_1241,N_615,N_829);
nor U1242 (N_1242,N_728,N_863);
and U1243 (N_1243,N_335,N_879);
nand U1244 (N_1244,N_935,N_452);
xnor U1245 (N_1245,N_215,N_947);
nand U1246 (N_1246,N_512,N_85);
nand U1247 (N_1247,N_556,N_153);
and U1248 (N_1248,N_503,N_789);
and U1249 (N_1249,N_830,N_746);
or U1250 (N_1250,N_34,N_663);
and U1251 (N_1251,N_340,N_724);
nand U1252 (N_1252,N_703,N_389);
or U1253 (N_1253,N_54,N_885);
or U1254 (N_1254,N_269,N_352);
nand U1255 (N_1255,N_617,N_920);
or U1256 (N_1256,N_776,N_447);
nand U1257 (N_1257,N_711,N_382);
nor U1258 (N_1258,N_277,N_259);
or U1259 (N_1259,N_229,N_777);
or U1260 (N_1260,N_10,N_791);
or U1261 (N_1261,N_442,N_779);
or U1262 (N_1262,N_159,N_517);
or U1263 (N_1263,N_647,N_182);
and U1264 (N_1264,N_474,N_428);
or U1265 (N_1265,N_130,N_592);
and U1266 (N_1266,N_683,N_102);
and U1267 (N_1267,N_713,N_709);
nor U1268 (N_1268,N_119,N_575);
nor U1269 (N_1269,N_331,N_297);
nand U1270 (N_1270,N_705,N_53);
nor U1271 (N_1271,N_725,N_207);
nor U1272 (N_1272,N_677,N_399);
and U1273 (N_1273,N_837,N_893);
or U1274 (N_1274,N_671,N_912);
nand U1275 (N_1275,N_840,N_249);
or U1276 (N_1276,N_354,N_200);
nor U1277 (N_1277,N_169,N_877);
nor U1278 (N_1278,N_795,N_807);
or U1279 (N_1279,N_304,N_36);
nand U1280 (N_1280,N_948,N_702);
or U1281 (N_1281,N_584,N_979);
nand U1282 (N_1282,N_158,N_852);
and U1283 (N_1283,N_467,N_92);
nand U1284 (N_1284,N_291,N_254);
nand U1285 (N_1285,N_723,N_950);
or U1286 (N_1286,N_891,N_951);
nor U1287 (N_1287,N_825,N_581);
or U1288 (N_1288,N_598,N_112);
and U1289 (N_1289,N_659,N_890);
and U1290 (N_1290,N_783,N_997);
nor U1291 (N_1291,N_270,N_616);
nand U1292 (N_1292,N_994,N_527);
nand U1293 (N_1293,N_596,N_343);
nor U1294 (N_1294,N_368,N_146);
nor U1295 (N_1295,N_589,N_24);
or U1296 (N_1296,N_28,N_714);
and U1297 (N_1297,N_377,N_231);
nand U1298 (N_1298,N_849,N_156);
nor U1299 (N_1299,N_230,N_91);
or U1300 (N_1300,N_661,N_626);
and U1301 (N_1301,N_771,N_261);
nor U1302 (N_1302,N_974,N_765);
nand U1303 (N_1303,N_55,N_396);
nor U1304 (N_1304,N_423,N_558);
nand U1305 (N_1305,N_360,N_622);
or U1306 (N_1306,N_49,N_972);
nor U1307 (N_1307,N_720,N_634);
nor U1308 (N_1308,N_899,N_263);
nand U1309 (N_1309,N_958,N_48);
or U1310 (N_1310,N_320,N_258);
and U1311 (N_1311,N_287,N_242);
or U1312 (N_1312,N_9,N_498);
or U1313 (N_1313,N_949,N_41);
nor U1314 (N_1314,N_326,N_344);
and U1315 (N_1315,N_722,N_993);
and U1316 (N_1316,N_623,N_14);
nand U1317 (N_1317,N_667,N_266);
or U1318 (N_1318,N_735,N_56);
nand U1319 (N_1319,N_51,N_946);
or U1320 (N_1320,N_924,N_110);
nor U1321 (N_1321,N_87,N_646);
nand U1322 (N_1322,N_479,N_817);
nand U1323 (N_1323,N_138,N_196);
nand U1324 (N_1324,N_886,N_605);
and U1325 (N_1325,N_704,N_810);
nor U1326 (N_1326,N_52,N_859);
nand U1327 (N_1327,N_292,N_23);
nor U1328 (N_1328,N_698,N_587);
nor U1329 (N_1329,N_397,N_441);
and U1330 (N_1330,N_788,N_597);
and U1331 (N_1331,N_392,N_487);
nor U1332 (N_1332,N_364,N_183);
nand U1333 (N_1333,N_40,N_778);
nor U1334 (N_1334,N_566,N_16);
nor U1335 (N_1335,N_539,N_497);
and U1336 (N_1336,N_445,N_3);
nor U1337 (N_1337,N_333,N_160);
or U1338 (N_1338,N_786,N_271);
or U1339 (N_1339,N_516,N_284);
nand U1340 (N_1340,N_184,N_255);
or U1341 (N_1341,N_290,N_805);
or U1342 (N_1342,N_601,N_405);
nor U1343 (N_1343,N_332,N_318);
nor U1344 (N_1344,N_424,N_166);
nand U1345 (N_1345,N_738,N_749);
nor U1346 (N_1346,N_514,N_298);
or U1347 (N_1347,N_383,N_743);
and U1348 (N_1348,N_203,N_828);
and U1349 (N_1349,N_515,N_956);
nor U1350 (N_1350,N_393,N_78);
and U1351 (N_1351,N_473,N_990);
and U1352 (N_1352,N_595,N_303);
nand U1353 (N_1353,N_300,N_763);
and U1354 (N_1354,N_655,N_252);
and U1355 (N_1355,N_992,N_375);
and U1356 (N_1356,N_232,N_57);
or U1357 (N_1357,N_607,N_443);
and U1358 (N_1358,N_293,N_134);
or U1359 (N_1359,N_371,N_752);
nand U1360 (N_1360,N_925,N_529);
nand U1361 (N_1361,N_624,N_214);
and U1362 (N_1362,N_411,N_446);
and U1363 (N_1363,N_628,N_127);
or U1364 (N_1364,N_305,N_143);
and U1365 (N_1365,N_871,N_142);
nand U1366 (N_1366,N_80,N_896);
nand U1367 (N_1367,N_794,N_220);
nand U1368 (N_1368,N_842,N_295);
nand U1369 (N_1369,N_754,N_494);
and U1370 (N_1370,N_511,N_670);
nor U1371 (N_1371,N_103,N_536);
or U1372 (N_1372,N_509,N_866);
nor U1373 (N_1373,N_895,N_542);
and U1374 (N_1374,N_699,N_831);
and U1375 (N_1375,N_650,N_414);
or U1376 (N_1376,N_870,N_353);
nor U1377 (N_1377,N_115,N_691);
and U1378 (N_1378,N_954,N_844);
nor U1379 (N_1379,N_44,N_107);
and U1380 (N_1380,N_236,N_437);
nor U1381 (N_1381,N_611,N_430);
and U1382 (N_1382,N_673,N_327);
or U1383 (N_1383,N_770,N_571);
nand U1384 (N_1384,N_47,N_206);
nor U1385 (N_1385,N_522,N_306);
or U1386 (N_1386,N_901,N_312);
nand U1387 (N_1387,N_832,N_90);
nor U1388 (N_1388,N_157,N_93);
nand U1389 (N_1389,N_757,N_433);
or U1390 (N_1390,N_324,N_345);
xnor U1391 (N_1391,N_109,N_482);
nand U1392 (N_1392,N_275,N_590);
or U1393 (N_1393,N_387,N_420);
nor U1394 (N_1394,N_45,N_13);
and U1395 (N_1395,N_660,N_736);
nand U1396 (N_1396,N_417,N_639);
nand U1397 (N_1397,N_531,N_588);
nor U1398 (N_1398,N_808,N_914);
or U1399 (N_1399,N_576,N_726);
nor U1400 (N_1400,N_416,N_268);
nor U1401 (N_1401,N_578,N_564);
nor U1402 (N_1402,N_491,N_755);
and U1403 (N_1403,N_493,N_83);
nand U1404 (N_1404,N_279,N_89);
nand U1405 (N_1405,N_882,N_141);
or U1406 (N_1406,N_30,N_774);
nor U1407 (N_1407,N_245,N_906);
nand U1408 (N_1408,N_216,N_532);
or U1409 (N_1409,N_697,N_614);
nand U1410 (N_1410,N_175,N_629);
nand U1411 (N_1411,N_797,N_767);
nor U1412 (N_1412,N_843,N_325);
nor U1413 (N_1413,N_286,N_488);
or U1414 (N_1414,N_676,N_941);
nand U1415 (N_1415,N_851,N_379);
nor U1416 (N_1416,N_672,N_818);
nand U1417 (N_1417,N_546,N_619);
and U1418 (N_1418,N_729,N_465);
or U1419 (N_1419,N_1,N_355);
nand U1420 (N_1420,N_29,N_700);
nor U1421 (N_1421,N_384,N_841);
or U1422 (N_1422,N_620,N_453);
and U1423 (N_1423,N_854,N_366);
nand U1424 (N_1424,N_690,N_19);
nor U1425 (N_1425,N_996,N_567);
nor U1426 (N_1426,N_892,N_225);
nand U1427 (N_1427,N_707,N_900);
nor U1428 (N_1428,N_800,N_751);
nor U1429 (N_1429,N_627,N_694);
or U1430 (N_1430,N_506,N_11);
or U1431 (N_1431,N_505,N_222);
nor U1432 (N_1432,N_260,N_848);
nand U1433 (N_1433,N_188,N_687);
or U1434 (N_1434,N_282,N_444);
nor U1435 (N_1435,N_278,N_193);
and U1436 (N_1436,N_717,N_7);
and U1437 (N_1437,N_221,N_827);
nand U1438 (N_1438,N_201,N_991);
nor U1439 (N_1439,N_204,N_123);
nor U1440 (N_1440,N_378,N_939);
nand U1441 (N_1441,N_525,N_963);
nor U1442 (N_1442,N_630,N_610);
nand U1443 (N_1443,N_499,N_712);
nand U1444 (N_1444,N_910,N_815);
and U1445 (N_1445,N_526,N_621);
and U1446 (N_1446,N_923,N_695);
nor U1447 (N_1447,N_929,N_202);
xnor U1448 (N_1448,N_337,N_435);
nand U1449 (N_1449,N_570,N_197);
nor U1450 (N_1450,N_347,N_105);
and U1451 (N_1451,N_930,N_861);
and U1452 (N_1452,N_985,N_492);
and U1453 (N_1453,N_933,N_775);
and U1454 (N_1454,N_524,N_70);
and U1455 (N_1455,N_823,N_154);
or U1456 (N_1456,N_177,N_65);
or U1457 (N_1457,N_887,N_543);
nand U1458 (N_1458,N_457,N_548);
nor U1459 (N_1459,N_604,N_648);
nand U1460 (N_1460,N_15,N_114);
nor U1461 (N_1461,N_928,N_334);
nor U1462 (N_1462,N_739,N_764);
nand U1463 (N_1463,N_180,N_875);
and U1464 (N_1464,N_46,N_122);
or U1465 (N_1465,N_338,N_495);
or U1466 (N_1466,N_533,N_745);
or U1467 (N_1467,N_636,N_678);
nor U1468 (N_1468,N_884,N_98);
nor U1469 (N_1469,N_944,N_934);
nand U1470 (N_1470,N_583,N_460);
and U1471 (N_1471,N_81,N_365);
and U1472 (N_1472,N_897,N_613);
nand U1473 (N_1473,N_753,N_174);
nand U1474 (N_1474,N_679,N_518);
or U1475 (N_1475,N_537,N_782);
or U1476 (N_1476,N_916,N_865);
and U1477 (N_1477,N_361,N_680);
or U1478 (N_1478,N_936,N_734);
nor U1479 (N_1479,N_328,N_978);
or U1480 (N_1480,N_257,N_480);
and U1481 (N_1481,N_649,N_299);
and U1482 (N_1482,N_485,N_802);
or U1483 (N_1483,N_572,N_504);
nor U1484 (N_1484,N_178,N_508);
nand U1485 (N_1485,N_274,N_552);
nor U1486 (N_1486,N_803,N_171);
nor U1487 (N_1487,N_248,N_747);
or U1488 (N_1488,N_982,N_812);
and U1489 (N_1489,N_967,N_857);
nor U1490 (N_1490,N_662,N_97);
nor U1491 (N_1491,N_339,N_317);
nor U1492 (N_1492,N_99,N_469);
nor U1493 (N_1493,N_113,N_876);
and U1494 (N_1494,N_139,N_477);
nand U1495 (N_1495,N_565,N_625);
or U1496 (N_1496,N_336,N_826);
and U1497 (N_1497,N_238,N_657);
nor U1498 (N_1498,N_358,N_426);
nor U1499 (N_1499,N_310,N_573);
nand U1500 (N_1500,N_699,N_751);
or U1501 (N_1501,N_182,N_148);
or U1502 (N_1502,N_967,N_680);
and U1503 (N_1503,N_394,N_499);
or U1504 (N_1504,N_387,N_676);
nand U1505 (N_1505,N_733,N_169);
or U1506 (N_1506,N_381,N_865);
or U1507 (N_1507,N_273,N_432);
nand U1508 (N_1508,N_687,N_479);
nor U1509 (N_1509,N_756,N_413);
or U1510 (N_1510,N_964,N_259);
and U1511 (N_1511,N_67,N_308);
and U1512 (N_1512,N_677,N_128);
or U1513 (N_1513,N_707,N_291);
nand U1514 (N_1514,N_188,N_922);
nand U1515 (N_1515,N_889,N_57);
nand U1516 (N_1516,N_636,N_217);
nand U1517 (N_1517,N_227,N_533);
nand U1518 (N_1518,N_421,N_831);
nand U1519 (N_1519,N_175,N_14);
nand U1520 (N_1520,N_53,N_220);
or U1521 (N_1521,N_860,N_104);
nor U1522 (N_1522,N_661,N_474);
nand U1523 (N_1523,N_595,N_443);
nand U1524 (N_1524,N_500,N_928);
nand U1525 (N_1525,N_593,N_351);
and U1526 (N_1526,N_642,N_966);
nand U1527 (N_1527,N_415,N_912);
or U1528 (N_1528,N_972,N_486);
and U1529 (N_1529,N_142,N_445);
and U1530 (N_1530,N_223,N_518);
nand U1531 (N_1531,N_698,N_704);
nor U1532 (N_1532,N_173,N_497);
nand U1533 (N_1533,N_967,N_217);
or U1534 (N_1534,N_309,N_441);
and U1535 (N_1535,N_458,N_230);
or U1536 (N_1536,N_746,N_821);
nor U1537 (N_1537,N_946,N_622);
nor U1538 (N_1538,N_401,N_978);
or U1539 (N_1539,N_747,N_977);
nor U1540 (N_1540,N_825,N_846);
nand U1541 (N_1541,N_721,N_648);
nor U1542 (N_1542,N_51,N_784);
and U1543 (N_1543,N_296,N_331);
nor U1544 (N_1544,N_65,N_465);
and U1545 (N_1545,N_977,N_593);
nand U1546 (N_1546,N_262,N_81);
and U1547 (N_1547,N_252,N_99);
nand U1548 (N_1548,N_457,N_18);
nand U1549 (N_1549,N_789,N_110);
nor U1550 (N_1550,N_788,N_185);
and U1551 (N_1551,N_726,N_611);
or U1552 (N_1552,N_296,N_368);
nand U1553 (N_1553,N_750,N_354);
and U1554 (N_1554,N_724,N_746);
and U1555 (N_1555,N_433,N_519);
nor U1556 (N_1556,N_8,N_279);
nor U1557 (N_1557,N_309,N_423);
nand U1558 (N_1558,N_547,N_653);
nor U1559 (N_1559,N_105,N_313);
or U1560 (N_1560,N_368,N_110);
nor U1561 (N_1561,N_711,N_587);
or U1562 (N_1562,N_222,N_92);
nand U1563 (N_1563,N_314,N_608);
or U1564 (N_1564,N_102,N_672);
nor U1565 (N_1565,N_300,N_660);
nand U1566 (N_1566,N_306,N_815);
nand U1567 (N_1567,N_139,N_869);
and U1568 (N_1568,N_933,N_82);
and U1569 (N_1569,N_105,N_332);
nand U1570 (N_1570,N_464,N_139);
and U1571 (N_1571,N_410,N_513);
or U1572 (N_1572,N_892,N_58);
nand U1573 (N_1573,N_225,N_317);
or U1574 (N_1574,N_234,N_937);
and U1575 (N_1575,N_903,N_506);
nand U1576 (N_1576,N_80,N_773);
and U1577 (N_1577,N_342,N_361);
nand U1578 (N_1578,N_484,N_367);
nand U1579 (N_1579,N_419,N_555);
or U1580 (N_1580,N_744,N_673);
or U1581 (N_1581,N_504,N_173);
or U1582 (N_1582,N_868,N_851);
and U1583 (N_1583,N_239,N_733);
or U1584 (N_1584,N_726,N_830);
or U1585 (N_1585,N_153,N_945);
nor U1586 (N_1586,N_538,N_646);
nand U1587 (N_1587,N_781,N_569);
nor U1588 (N_1588,N_990,N_299);
nor U1589 (N_1589,N_854,N_231);
or U1590 (N_1590,N_416,N_340);
or U1591 (N_1591,N_150,N_768);
and U1592 (N_1592,N_970,N_149);
or U1593 (N_1593,N_447,N_304);
nand U1594 (N_1594,N_476,N_320);
nand U1595 (N_1595,N_351,N_691);
nor U1596 (N_1596,N_202,N_830);
and U1597 (N_1597,N_424,N_108);
and U1598 (N_1598,N_682,N_170);
and U1599 (N_1599,N_662,N_913);
and U1600 (N_1600,N_826,N_40);
and U1601 (N_1601,N_916,N_370);
nand U1602 (N_1602,N_159,N_539);
or U1603 (N_1603,N_718,N_680);
nor U1604 (N_1604,N_208,N_863);
nand U1605 (N_1605,N_977,N_482);
nand U1606 (N_1606,N_829,N_15);
and U1607 (N_1607,N_331,N_734);
or U1608 (N_1608,N_90,N_259);
nand U1609 (N_1609,N_859,N_911);
and U1610 (N_1610,N_136,N_0);
nor U1611 (N_1611,N_222,N_978);
nor U1612 (N_1612,N_394,N_836);
nand U1613 (N_1613,N_798,N_596);
and U1614 (N_1614,N_748,N_275);
nor U1615 (N_1615,N_890,N_521);
and U1616 (N_1616,N_667,N_755);
or U1617 (N_1617,N_243,N_801);
or U1618 (N_1618,N_332,N_776);
and U1619 (N_1619,N_524,N_145);
nor U1620 (N_1620,N_498,N_452);
nor U1621 (N_1621,N_601,N_901);
or U1622 (N_1622,N_318,N_515);
or U1623 (N_1623,N_102,N_700);
and U1624 (N_1624,N_469,N_664);
or U1625 (N_1625,N_653,N_651);
nand U1626 (N_1626,N_97,N_487);
and U1627 (N_1627,N_197,N_503);
and U1628 (N_1628,N_888,N_749);
nand U1629 (N_1629,N_871,N_164);
and U1630 (N_1630,N_563,N_314);
and U1631 (N_1631,N_786,N_559);
nand U1632 (N_1632,N_223,N_645);
and U1633 (N_1633,N_301,N_105);
nor U1634 (N_1634,N_504,N_977);
and U1635 (N_1635,N_700,N_874);
nor U1636 (N_1636,N_117,N_855);
nor U1637 (N_1637,N_573,N_259);
nand U1638 (N_1638,N_912,N_475);
or U1639 (N_1639,N_883,N_21);
and U1640 (N_1640,N_967,N_481);
and U1641 (N_1641,N_287,N_687);
nor U1642 (N_1642,N_307,N_572);
nand U1643 (N_1643,N_577,N_391);
and U1644 (N_1644,N_154,N_880);
or U1645 (N_1645,N_920,N_396);
or U1646 (N_1646,N_573,N_260);
nand U1647 (N_1647,N_492,N_157);
and U1648 (N_1648,N_706,N_784);
and U1649 (N_1649,N_469,N_153);
or U1650 (N_1650,N_542,N_642);
and U1651 (N_1651,N_462,N_484);
and U1652 (N_1652,N_931,N_523);
nand U1653 (N_1653,N_612,N_940);
nand U1654 (N_1654,N_740,N_230);
nand U1655 (N_1655,N_397,N_936);
and U1656 (N_1656,N_132,N_851);
nand U1657 (N_1657,N_964,N_572);
nor U1658 (N_1658,N_689,N_186);
and U1659 (N_1659,N_904,N_886);
nor U1660 (N_1660,N_296,N_941);
and U1661 (N_1661,N_374,N_828);
nor U1662 (N_1662,N_437,N_797);
and U1663 (N_1663,N_203,N_35);
nor U1664 (N_1664,N_525,N_513);
nand U1665 (N_1665,N_967,N_779);
nor U1666 (N_1666,N_102,N_745);
or U1667 (N_1667,N_342,N_373);
nor U1668 (N_1668,N_39,N_241);
and U1669 (N_1669,N_719,N_4);
or U1670 (N_1670,N_641,N_924);
nand U1671 (N_1671,N_637,N_607);
nor U1672 (N_1672,N_896,N_310);
or U1673 (N_1673,N_350,N_71);
and U1674 (N_1674,N_797,N_760);
nor U1675 (N_1675,N_358,N_684);
nor U1676 (N_1676,N_427,N_821);
nand U1677 (N_1677,N_114,N_106);
nand U1678 (N_1678,N_711,N_50);
and U1679 (N_1679,N_874,N_188);
or U1680 (N_1680,N_337,N_9);
or U1681 (N_1681,N_229,N_959);
nor U1682 (N_1682,N_259,N_581);
nand U1683 (N_1683,N_551,N_507);
nand U1684 (N_1684,N_720,N_878);
nor U1685 (N_1685,N_496,N_36);
and U1686 (N_1686,N_156,N_237);
or U1687 (N_1687,N_497,N_917);
or U1688 (N_1688,N_57,N_650);
or U1689 (N_1689,N_124,N_422);
nor U1690 (N_1690,N_887,N_690);
and U1691 (N_1691,N_712,N_55);
nor U1692 (N_1692,N_834,N_917);
nor U1693 (N_1693,N_32,N_368);
and U1694 (N_1694,N_476,N_616);
and U1695 (N_1695,N_524,N_59);
nand U1696 (N_1696,N_309,N_793);
nand U1697 (N_1697,N_680,N_130);
and U1698 (N_1698,N_516,N_638);
or U1699 (N_1699,N_307,N_769);
or U1700 (N_1700,N_478,N_454);
nand U1701 (N_1701,N_743,N_746);
nand U1702 (N_1702,N_655,N_707);
or U1703 (N_1703,N_348,N_926);
or U1704 (N_1704,N_119,N_464);
or U1705 (N_1705,N_243,N_728);
nor U1706 (N_1706,N_295,N_915);
and U1707 (N_1707,N_78,N_638);
and U1708 (N_1708,N_175,N_781);
nor U1709 (N_1709,N_852,N_449);
or U1710 (N_1710,N_828,N_779);
and U1711 (N_1711,N_914,N_880);
or U1712 (N_1712,N_518,N_33);
nand U1713 (N_1713,N_517,N_25);
and U1714 (N_1714,N_800,N_298);
nand U1715 (N_1715,N_812,N_117);
and U1716 (N_1716,N_946,N_742);
or U1717 (N_1717,N_215,N_570);
or U1718 (N_1718,N_405,N_303);
and U1719 (N_1719,N_256,N_343);
or U1720 (N_1720,N_86,N_808);
nand U1721 (N_1721,N_17,N_899);
nor U1722 (N_1722,N_906,N_775);
nand U1723 (N_1723,N_343,N_787);
nor U1724 (N_1724,N_63,N_179);
and U1725 (N_1725,N_162,N_328);
and U1726 (N_1726,N_867,N_990);
nand U1727 (N_1727,N_869,N_243);
or U1728 (N_1728,N_795,N_435);
and U1729 (N_1729,N_943,N_35);
and U1730 (N_1730,N_243,N_251);
nand U1731 (N_1731,N_225,N_263);
nand U1732 (N_1732,N_758,N_766);
nand U1733 (N_1733,N_219,N_849);
or U1734 (N_1734,N_803,N_60);
or U1735 (N_1735,N_604,N_859);
nor U1736 (N_1736,N_172,N_929);
nand U1737 (N_1737,N_946,N_746);
or U1738 (N_1738,N_238,N_214);
nand U1739 (N_1739,N_101,N_559);
nand U1740 (N_1740,N_686,N_51);
nor U1741 (N_1741,N_819,N_810);
nor U1742 (N_1742,N_184,N_985);
nor U1743 (N_1743,N_580,N_343);
and U1744 (N_1744,N_207,N_827);
nor U1745 (N_1745,N_18,N_542);
or U1746 (N_1746,N_558,N_352);
or U1747 (N_1747,N_397,N_925);
and U1748 (N_1748,N_722,N_377);
or U1749 (N_1749,N_931,N_865);
or U1750 (N_1750,N_367,N_747);
nor U1751 (N_1751,N_303,N_490);
nor U1752 (N_1752,N_604,N_878);
nand U1753 (N_1753,N_726,N_505);
and U1754 (N_1754,N_807,N_73);
nor U1755 (N_1755,N_354,N_167);
nand U1756 (N_1756,N_530,N_718);
and U1757 (N_1757,N_907,N_116);
or U1758 (N_1758,N_307,N_282);
nand U1759 (N_1759,N_480,N_216);
and U1760 (N_1760,N_869,N_753);
nand U1761 (N_1761,N_570,N_990);
or U1762 (N_1762,N_103,N_670);
or U1763 (N_1763,N_864,N_820);
and U1764 (N_1764,N_658,N_461);
and U1765 (N_1765,N_20,N_15);
nor U1766 (N_1766,N_855,N_875);
xor U1767 (N_1767,N_614,N_241);
or U1768 (N_1768,N_588,N_872);
nor U1769 (N_1769,N_789,N_401);
nand U1770 (N_1770,N_223,N_913);
nor U1771 (N_1771,N_382,N_44);
nand U1772 (N_1772,N_969,N_452);
or U1773 (N_1773,N_870,N_815);
or U1774 (N_1774,N_474,N_116);
or U1775 (N_1775,N_230,N_576);
and U1776 (N_1776,N_564,N_519);
and U1777 (N_1777,N_532,N_823);
nor U1778 (N_1778,N_849,N_726);
or U1779 (N_1779,N_328,N_304);
nand U1780 (N_1780,N_935,N_873);
and U1781 (N_1781,N_848,N_632);
and U1782 (N_1782,N_347,N_672);
nor U1783 (N_1783,N_522,N_332);
nor U1784 (N_1784,N_586,N_282);
and U1785 (N_1785,N_868,N_900);
xnor U1786 (N_1786,N_850,N_880);
nand U1787 (N_1787,N_803,N_223);
nor U1788 (N_1788,N_527,N_668);
nand U1789 (N_1789,N_722,N_241);
nand U1790 (N_1790,N_316,N_786);
nor U1791 (N_1791,N_101,N_284);
nor U1792 (N_1792,N_77,N_449);
nor U1793 (N_1793,N_865,N_467);
nor U1794 (N_1794,N_55,N_616);
and U1795 (N_1795,N_576,N_557);
and U1796 (N_1796,N_769,N_601);
nand U1797 (N_1797,N_689,N_246);
nand U1798 (N_1798,N_236,N_514);
and U1799 (N_1799,N_122,N_154);
or U1800 (N_1800,N_696,N_805);
and U1801 (N_1801,N_494,N_127);
and U1802 (N_1802,N_327,N_669);
or U1803 (N_1803,N_269,N_764);
or U1804 (N_1804,N_266,N_292);
and U1805 (N_1805,N_116,N_38);
nor U1806 (N_1806,N_289,N_65);
nor U1807 (N_1807,N_626,N_880);
nand U1808 (N_1808,N_789,N_548);
nor U1809 (N_1809,N_76,N_988);
and U1810 (N_1810,N_763,N_338);
or U1811 (N_1811,N_964,N_470);
nand U1812 (N_1812,N_89,N_496);
nand U1813 (N_1813,N_837,N_88);
and U1814 (N_1814,N_685,N_546);
nand U1815 (N_1815,N_519,N_321);
nand U1816 (N_1816,N_62,N_528);
and U1817 (N_1817,N_627,N_255);
nand U1818 (N_1818,N_233,N_535);
nor U1819 (N_1819,N_68,N_210);
nand U1820 (N_1820,N_870,N_761);
and U1821 (N_1821,N_406,N_39);
xor U1822 (N_1822,N_381,N_606);
and U1823 (N_1823,N_482,N_557);
or U1824 (N_1824,N_101,N_976);
nor U1825 (N_1825,N_922,N_219);
and U1826 (N_1826,N_794,N_554);
and U1827 (N_1827,N_436,N_661);
and U1828 (N_1828,N_904,N_735);
or U1829 (N_1829,N_832,N_731);
nor U1830 (N_1830,N_752,N_121);
nand U1831 (N_1831,N_36,N_734);
nor U1832 (N_1832,N_103,N_443);
nand U1833 (N_1833,N_433,N_74);
and U1834 (N_1834,N_28,N_456);
and U1835 (N_1835,N_936,N_371);
nand U1836 (N_1836,N_410,N_567);
nand U1837 (N_1837,N_110,N_968);
and U1838 (N_1838,N_176,N_788);
and U1839 (N_1839,N_732,N_157);
nand U1840 (N_1840,N_156,N_730);
nand U1841 (N_1841,N_829,N_604);
nor U1842 (N_1842,N_255,N_313);
nand U1843 (N_1843,N_133,N_565);
nand U1844 (N_1844,N_424,N_653);
or U1845 (N_1845,N_676,N_449);
nor U1846 (N_1846,N_806,N_376);
nor U1847 (N_1847,N_941,N_276);
nor U1848 (N_1848,N_46,N_210);
or U1849 (N_1849,N_852,N_733);
and U1850 (N_1850,N_156,N_332);
xnor U1851 (N_1851,N_895,N_853);
xnor U1852 (N_1852,N_35,N_711);
nor U1853 (N_1853,N_819,N_29);
nor U1854 (N_1854,N_193,N_798);
and U1855 (N_1855,N_525,N_536);
and U1856 (N_1856,N_801,N_714);
nor U1857 (N_1857,N_89,N_908);
or U1858 (N_1858,N_304,N_392);
nor U1859 (N_1859,N_817,N_483);
nand U1860 (N_1860,N_811,N_184);
nand U1861 (N_1861,N_229,N_196);
and U1862 (N_1862,N_227,N_387);
or U1863 (N_1863,N_796,N_931);
nor U1864 (N_1864,N_578,N_160);
and U1865 (N_1865,N_936,N_671);
nor U1866 (N_1866,N_880,N_716);
nand U1867 (N_1867,N_384,N_178);
and U1868 (N_1868,N_482,N_963);
nor U1869 (N_1869,N_706,N_696);
or U1870 (N_1870,N_203,N_935);
or U1871 (N_1871,N_931,N_847);
or U1872 (N_1872,N_531,N_755);
and U1873 (N_1873,N_667,N_540);
nand U1874 (N_1874,N_547,N_665);
or U1875 (N_1875,N_86,N_501);
nor U1876 (N_1876,N_649,N_29);
or U1877 (N_1877,N_101,N_517);
nor U1878 (N_1878,N_95,N_967);
nor U1879 (N_1879,N_248,N_850);
and U1880 (N_1880,N_917,N_977);
and U1881 (N_1881,N_154,N_13);
nor U1882 (N_1882,N_954,N_769);
and U1883 (N_1883,N_452,N_794);
nor U1884 (N_1884,N_255,N_50);
nand U1885 (N_1885,N_329,N_925);
or U1886 (N_1886,N_967,N_922);
and U1887 (N_1887,N_529,N_947);
and U1888 (N_1888,N_158,N_219);
nand U1889 (N_1889,N_408,N_874);
nor U1890 (N_1890,N_376,N_563);
or U1891 (N_1891,N_751,N_474);
and U1892 (N_1892,N_48,N_825);
and U1893 (N_1893,N_665,N_831);
nand U1894 (N_1894,N_224,N_538);
or U1895 (N_1895,N_53,N_311);
nand U1896 (N_1896,N_364,N_636);
nand U1897 (N_1897,N_356,N_919);
and U1898 (N_1898,N_633,N_771);
nand U1899 (N_1899,N_274,N_413);
or U1900 (N_1900,N_482,N_280);
and U1901 (N_1901,N_658,N_896);
nor U1902 (N_1902,N_523,N_143);
and U1903 (N_1903,N_764,N_870);
nor U1904 (N_1904,N_811,N_903);
nand U1905 (N_1905,N_184,N_990);
or U1906 (N_1906,N_963,N_186);
nor U1907 (N_1907,N_540,N_945);
or U1908 (N_1908,N_183,N_325);
or U1909 (N_1909,N_402,N_993);
nand U1910 (N_1910,N_223,N_529);
nor U1911 (N_1911,N_694,N_304);
nor U1912 (N_1912,N_496,N_783);
nor U1913 (N_1913,N_415,N_419);
nor U1914 (N_1914,N_427,N_51);
nor U1915 (N_1915,N_249,N_734);
or U1916 (N_1916,N_135,N_37);
nor U1917 (N_1917,N_479,N_206);
or U1918 (N_1918,N_657,N_354);
nor U1919 (N_1919,N_843,N_992);
and U1920 (N_1920,N_308,N_453);
and U1921 (N_1921,N_929,N_279);
and U1922 (N_1922,N_61,N_993);
nor U1923 (N_1923,N_721,N_713);
and U1924 (N_1924,N_568,N_710);
nand U1925 (N_1925,N_738,N_405);
xnor U1926 (N_1926,N_273,N_864);
nor U1927 (N_1927,N_248,N_899);
or U1928 (N_1928,N_588,N_194);
nor U1929 (N_1929,N_401,N_403);
nor U1930 (N_1930,N_444,N_518);
or U1931 (N_1931,N_79,N_391);
and U1932 (N_1932,N_414,N_406);
or U1933 (N_1933,N_453,N_304);
or U1934 (N_1934,N_658,N_730);
nor U1935 (N_1935,N_328,N_758);
xnor U1936 (N_1936,N_398,N_654);
and U1937 (N_1937,N_486,N_872);
or U1938 (N_1938,N_853,N_288);
nor U1939 (N_1939,N_578,N_831);
nand U1940 (N_1940,N_332,N_822);
or U1941 (N_1941,N_521,N_256);
and U1942 (N_1942,N_954,N_659);
or U1943 (N_1943,N_791,N_15);
and U1944 (N_1944,N_178,N_549);
and U1945 (N_1945,N_993,N_758);
nand U1946 (N_1946,N_569,N_697);
nand U1947 (N_1947,N_108,N_200);
nand U1948 (N_1948,N_847,N_597);
nand U1949 (N_1949,N_797,N_249);
nor U1950 (N_1950,N_579,N_41);
and U1951 (N_1951,N_181,N_199);
or U1952 (N_1952,N_220,N_90);
and U1953 (N_1953,N_459,N_629);
or U1954 (N_1954,N_517,N_255);
or U1955 (N_1955,N_837,N_699);
nor U1956 (N_1956,N_963,N_106);
or U1957 (N_1957,N_790,N_86);
nor U1958 (N_1958,N_949,N_257);
or U1959 (N_1959,N_881,N_966);
or U1960 (N_1960,N_206,N_508);
or U1961 (N_1961,N_623,N_62);
and U1962 (N_1962,N_144,N_524);
nand U1963 (N_1963,N_67,N_673);
nor U1964 (N_1964,N_386,N_688);
or U1965 (N_1965,N_681,N_67);
nand U1966 (N_1966,N_391,N_801);
and U1967 (N_1967,N_1,N_516);
and U1968 (N_1968,N_106,N_107);
and U1969 (N_1969,N_499,N_925);
or U1970 (N_1970,N_713,N_531);
xnor U1971 (N_1971,N_313,N_548);
nand U1972 (N_1972,N_542,N_231);
nor U1973 (N_1973,N_342,N_743);
and U1974 (N_1974,N_460,N_923);
or U1975 (N_1975,N_792,N_235);
nor U1976 (N_1976,N_916,N_329);
or U1977 (N_1977,N_343,N_321);
nor U1978 (N_1978,N_37,N_450);
or U1979 (N_1979,N_210,N_347);
or U1980 (N_1980,N_232,N_357);
nand U1981 (N_1981,N_91,N_990);
nand U1982 (N_1982,N_696,N_694);
or U1983 (N_1983,N_303,N_855);
and U1984 (N_1984,N_142,N_210);
nor U1985 (N_1985,N_388,N_951);
nor U1986 (N_1986,N_707,N_202);
nand U1987 (N_1987,N_344,N_27);
nand U1988 (N_1988,N_557,N_564);
or U1989 (N_1989,N_726,N_869);
or U1990 (N_1990,N_216,N_296);
nor U1991 (N_1991,N_632,N_182);
nand U1992 (N_1992,N_306,N_593);
or U1993 (N_1993,N_60,N_970);
and U1994 (N_1994,N_587,N_77);
or U1995 (N_1995,N_172,N_97);
and U1996 (N_1996,N_268,N_157);
and U1997 (N_1997,N_721,N_373);
nor U1998 (N_1998,N_984,N_832);
or U1999 (N_1999,N_51,N_74);
nand U2000 (N_2000,N_1816,N_1351);
or U2001 (N_2001,N_1422,N_1118);
and U2002 (N_2002,N_1829,N_1628);
nand U2003 (N_2003,N_1898,N_1493);
or U2004 (N_2004,N_1059,N_1964);
nor U2005 (N_2005,N_1764,N_1657);
nand U2006 (N_2006,N_1874,N_1935);
and U2007 (N_2007,N_1592,N_1536);
or U2008 (N_2008,N_1086,N_1809);
or U2009 (N_2009,N_1116,N_1355);
nand U2010 (N_2010,N_1113,N_1019);
and U2011 (N_2011,N_1565,N_1103);
nor U2012 (N_2012,N_1184,N_1044);
xor U2013 (N_2013,N_1121,N_1675);
and U2014 (N_2014,N_1597,N_1230);
and U2015 (N_2015,N_1210,N_1265);
xor U2016 (N_2016,N_1552,N_1715);
nor U2017 (N_2017,N_1153,N_1143);
nor U2018 (N_2018,N_1582,N_1489);
nand U2019 (N_2019,N_1701,N_1421);
and U2020 (N_2020,N_1713,N_1138);
or U2021 (N_2021,N_1226,N_1278);
nand U2022 (N_2022,N_1036,N_1728);
nand U2023 (N_2023,N_1252,N_1947);
or U2024 (N_2024,N_1216,N_1432);
nand U2025 (N_2025,N_1100,N_1128);
and U2026 (N_2026,N_1000,N_1900);
and U2027 (N_2027,N_1570,N_1065);
nor U2028 (N_2028,N_1533,N_1320);
nand U2029 (N_2029,N_1682,N_1600);
or U2030 (N_2030,N_1419,N_1613);
and U2031 (N_2031,N_1304,N_1798);
nor U2032 (N_2032,N_1013,N_1211);
nor U2033 (N_2033,N_1806,N_1703);
nor U2034 (N_2034,N_1585,N_1665);
or U2035 (N_2035,N_1788,N_1733);
or U2036 (N_2036,N_1574,N_1295);
nand U2037 (N_2037,N_1050,N_1659);
and U2038 (N_2038,N_1073,N_1054);
and U2039 (N_2039,N_1306,N_1417);
and U2040 (N_2040,N_1404,N_1207);
or U2041 (N_2041,N_1077,N_1316);
or U2042 (N_2042,N_1313,N_1603);
or U2043 (N_2043,N_1923,N_1812);
and U2044 (N_2044,N_1152,N_1414);
and U2045 (N_2045,N_1609,N_1003);
and U2046 (N_2046,N_1009,N_1068);
nor U2047 (N_2047,N_1174,N_1511);
and U2048 (N_2048,N_1443,N_1890);
and U2049 (N_2049,N_1260,N_1310);
or U2050 (N_2050,N_1276,N_1527);
nand U2051 (N_2051,N_1460,N_1187);
or U2052 (N_2052,N_1450,N_1672);
nand U2053 (N_2053,N_1225,N_1602);
nor U2054 (N_2054,N_1670,N_1357);
and U2055 (N_2055,N_1749,N_1752);
and U2056 (N_2056,N_1637,N_1215);
nand U2057 (N_2057,N_1409,N_1641);
nor U2058 (N_2058,N_1429,N_1286);
nor U2059 (N_2059,N_1283,N_1828);
and U2060 (N_2060,N_1905,N_1497);
or U2061 (N_2061,N_1040,N_1677);
nor U2062 (N_2062,N_1022,N_1244);
and U2063 (N_2063,N_1158,N_1366);
nor U2064 (N_2064,N_1302,N_1478);
and U2065 (N_2065,N_1714,N_1712);
nor U2066 (N_2066,N_1522,N_1643);
or U2067 (N_2067,N_1024,N_1888);
and U2068 (N_2068,N_1399,N_1902);
nand U2069 (N_2069,N_1862,N_1614);
or U2070 (N_2070,N_1605,N_1767);
nand U2071 (N_2071,N_1688,N_1931);
and U2072 (N_2072,N_1893,N_1243);
or U2073 (N_2073,N_1826,N_1157);
and U2074 (N_2074,N_1288,N_1342);
or U2075 (N_2075,N_1078,N_1966);
nand U2076 (N_2076,N_1198,N_1285);
and U2077 (N_2077,N_1651,N_1769);
and U2078 (N_2078,N_1615,N_1946);
and U2079 (N_2079,N_1411,N_1365);
nand U2080 (N_2080,N_1638,N_1123);
nor U2081 (N_2081,N_1831,N_1940);
and U2082 (N_2082,N_1624,N_1621);
nor U2083 (N_2083,N_1861,N_1937);
or U2084 (N_2084,N_1748,N_1977);
nand U2085 (N_2085,N_1192,N_1755);
and U2086 (N_2086,N_1704,N_1162);
or U2087 (N_2087,N_1047,N_1181);
or U2088 (N_2088,N_1319,N_1642);
nand U2089 (N_2089,N_1878,N_1096);
or U2090 (N_2090,N_1502,N_1515);
and U2091 (N_2091,N_1245,N_1989);
nand U2092 (N_2092,N_1870,N_1032);
or U2093 (N_2093,N_1514,N_1783);
nand U2094 (N_2094,N_1027,N_1154);
or U2095 (N_2095,N_1418,N_1132);
nor U2096 (N_2096,N_1996,N_1348);
and U2097 (N_2097,N_1089,N_1879);
nand U2098 (N_2098,N_1736,N_1988);
nor U2099 (N_2099,N_1063,N_1526);
nand U2100 (N_2100,N_1897,N_1978);
nand U2101 (N_2101,N_1340,N_1884);
nor U2102 (N_2102,N_1082,N_1377);
nor U2103 (N_2103,N_1137,N_1636);
or U2104 (N_2104,N_1135,N_1745);
and U2105 (N_2105,N_1317,N_1454);
and U2106 (N_2106,N_1049,N_1477);
nand U2107 (N_2107,N_1370,N_1982);
or U2108 (N_2108,N_1492,N_1667);
nand U2109 (N_2109,N_1516,N_1479);
and U2110 (N_2110,N_1075,N_1531);
and U2111 (N_2111,N_1336,N_1991);
nor U2112 (N_2112,N_1470,N_1620);
or U2113 (N_2113,N_1719,N_1384);
nand U2114 (N_2114,N_1622,N_1953);
and U2115 (N_2115,N_1508,N_1997);
and U2116 (N_2116,N_1220,N_1176);
nand U2117 (N_2117,N_1484,N_1420);
nor U2118 (N_2118,N_1505,N_1741);
nand U2119 (N_2119,N_1679,N_1165);
nand U2120 (N_2120,N_1026,N_1580);
nand U2121 (N_2121,N_1410,N_1892);
nor U2122 (N_2122,N_1030,N_1309);
nor U2123 (N_2123,N_1164,N_1841);
nor U2124 (N_2124,N_1494,N_1237);
nor U2125 (N_2125,N_1818,N_1510);
and U2126 (N_2126,N_1209,N_1335);
nor U2127 (N_2127,N_1392,N_1463);
nand U2128 (N_2128,N_1750,N_1326);
and U2129 (N_2129,N_1579,N_1687);
nor U2130 (N_2130,N_1822,N_1524);
and U2131 (N_2131,N_1765,N_1794);
or U2132 (N_2132,N_1932,N_1178);
nor U2133 (N_2133,N_1771,N_1218);
and U2134 (N_2134,N_1746,N_1438);
and U2135 (N_2135,N_1466,N_1800);
nand U2136 (N_2136,N_1199,N_1567);
or U2137 (N_2137,N_1721,N_1588);
nand U2138 (N_2138,N_1858,N_1876);
nor U2139 (N_2139,N_1254,N_1683);
nand U2140 (N_2140,N_1016,N_1911);
nand U2141 (N_2141,N_1980,N_1819);
nor U2142 (N_2142,N_1431,N_1127);
or U2143 (N_2143,N_1805,N_1412);
and U2144 (N_2144,N_1074,N_1247);
or U2145 (N_2145,N_1648,N_1272);
nand U2146 (N_2146,N_1266,N_1029);
or U2147 (N_2147,N_1994,N_1233);
or U2148 (N_2148,N_1166,N_1070);
nand U2149 (N_2149,N_1048,N_1590);
nand U2150 (N_2150,N_1148,N_1744);
nor U2151 (N_2151,N_1668,N_1426);
and U2152 (N_2152,N_1179,N_1232);
nor U2153 (N_2153,N_1601,N_1248);
nor U2154 (N_2154,N_1984,N_1042);
or U2155 (N_2155,N_1852,N_1180);
and U2156 (N_2156,N_1617,N_1720);
nor U2157 (N_2157,N_1844,N_1859);
nand U2158 (N_2158,N_1102,N_1802);
nand U2159 (N_2159,N_1041,N_1408);
nand U2160 (N_2160,N_1094,N_1627);
nor U2161 (N_2161,N_1223,N_1832);
nor U2162 (N_2162,N_1847,N_1710);
nand U2163 (N_2163,N_1145,N_1358);
and U2164 (N_2164,N_1033,N_1200);
and U2165 (N_2165,N_1448,N_1398);
nor U2166 (N_2166,N_1445,N_1891);
nor U2167 (N_2167,N_1772,N_1396);
and U2168 (N_2168,N_1471,N_1894);
nand U2169 (N_2169,N_1632,N_1866);
nand U2170 (N_2170,N_1294,N_1985);
and U2171 (N_2171,N_1051,N_1534);
nor U2172 (N_2172,N_1343,N_1589);
nand U2173 (N_2173,N_1287,N_1954);
nor U2174 (N_2174,N_1518,N_1095);
or U2175 (N_2175,N_1444,N_1101);
nand U2176 (N_2176,N_1452,N_1722);
or U2177 (N_2177,N_1385,N_1191);
and U2178 (N_2178,N_1405,N_1691);
and U2179 (N_2179,N_1246,N_1539);
nand U2180 (N_2180,N_1056,N_1299);
nor U2181 (N_2181,N_1387,N_1811);
xnor U2182 (N_2182,N_1882,N_1895);
and U2183 (N_2183,N_1833,N_1099);
or U2184 (N_2184,N_1924,N_1119);
nor U2185 (N_2185,N_1388,N_1616);
and U2186 (N_2186,N_1513,N_1052);
nand U2187 (N_2187,N_1079,N_1175);
nor U2188 (N_2188,N_1021,N_1725);
and U2189 (N_2189,N_1727,N_1034);
or U2190 (N_2190,N_1877,N_1427);
and U2191 (N_2191,N_1799,N_1548);
nand U2192 (N_2192,N_1674,N_1920);
nor U2193 (N_2193,N_1425,N_1259);
nand U2194 (N_2194,N_1381,N_1383);
nand U2195 (N_2195,N_1606,N_1347);
nand U2196 (N_2196,N_1066,N_1360);
or U2197 (N_2197,N_1705,N_1647);
or U2198 (N_2198,N_1723,N_1129);
or U2199 (N_2199,N_1650,N_1130);
or U2200 (N_2200,N_1992,N_1221);
nor U2201 (N_2201,N_1731,N_1664);
and U2202 (N_2202,N_1407,N_1639);
nand U2203 (N_2203,N_1329,N_1685);
or U2204 (N_2204,N_1436,N_1375);
or U2205 (N_2205,N_1491,N_1053);
xor U2206 (N_2206,N_1367,N_1442);
nand U2207 (N_2207,N_1969,N_1007);
or U2208 (N_2208,N_1564,N_1971);
nand U2209 (N_2209,N_1228,N_1255);
nor U2210 (N_2210,N_1631,N_1023);
or U2211 (N_2211,N_1171,N_1694);
and U2212 (N_2212,N_1577,N_1453);
and U2213 (N_2213,N_1440,N_1371);
and U2214 (N_2214,N_1553,N_1857);
or U2215 (N_2215,N_1069,N_1963);
nand U2216 (N_2216,N_1031,N_1568);
nand U2217 (N_2217,N_1406,N_1393);
nand U2218 (N_2218,N_1774,N_1311);
nand U2219 (N_2219,N_1110,N_1057);
or U2220 (N_2220,N_1693,N_1532);
nor U2221 (N_2221,N_1386,N_1901);
nand U2222 (N_2222,N_1836,N_1768);
or U2223 (N_2223,N_1521,N_1333);
xnor U2224 (N_2224,N_1608,N_1644);
nand U2225 (N_2225,N_1656,N_1562);
or U2226 (N_2226,N_1766,N_1530);
nor U2227 (N_2227,N_1775,N_1757);
nand U2228 (N_2228,N_1067,N_1280);
or U2229 (N_2229,N_1754,N_1362);
nor U2230 (N_2230,N_1908,N_1274);
nor U2231 (N_2231,N_1883,N_1625);
nand U2232 (N_2232,N_1555,N_1229);
nor U2233 (N_2233,N_1927,N_1331);
nand U2234 (N_2234,N_1382,N_1778);
and U2235 (N_2235,N_1610,N_1760);
and U2236 (N_2236,N_1341,N_1212);
nor U2237 (N_2237,N_1010,N_1784);
nor U2238 (N_2238,N_1441,N_1297);
nor U2239 (N_2239,N_1842,N_1979);
nand U2240 (N_2240,N_1576,N_1885);
or U2241 (N_2241,N_1481,N_1661);
and U2242 (N_2242,N_1186,N_1517);
or U2243 (N_2243,N_1433,N_1446);
and U2244 (N_2244,N_1213,N_1655);
and U2245 (N_2245,N_1827,N_1763);
nor U2246 (N_2246,N_1324,N_1835);
nand U2247 (N_2247,N_1361,N_1965);
and U2248 (N_2248,N_1626,N_1640);
or U2249 (N_2249,N_1104,N_1843);
and U2250 (N_2250,N_1364,N_1630);
or U2251 (N_2251,N_1261,N_1017);
nor U2252 (N_2252,N_1476,N_1787);
and U2253 (N_2253,N_1087,N_1743);
or U2254 (N_2254,N_1379,N_1612);
and U2255 (N_2255,N_1993,N_1144);
and U2256 (N_2256,N_1934,N_1190);
nand U2257 (N_2257,N_1867,N_1338);
nor U2258 (N_2258,N_1240,N_1962);
and U2259 (N_2259,N_1863,N_1005);
and U2260 (N_2260,N_1195,N_1975);
and U2261 (N_2261,N_1762,N_1973);
or U2262 (N_2262,N_1345,N_1334);
nand U2263 (N_2263,N_1015,N_1234);
or U2264 (N_2264,N_1595,N_1566);
and U2265 (N_2265,N_1008,N_1439);
nand U2266 (N_2266,N_1730,N_1793);
nor U2267 (N_2267,N_1424,N_1035);
or U2268 (N_2268,N_1235,N_1456);
nand U2269 (N_2269,N_1193,N_1461);
nor U2270 (N_2270,N_1270,N_1584);
or U2271 (N_2271,N_1596,N_1196);
and U2272 (N_2272,N_1170,N_1671);
nand U2273 (N_2273,N_1084,N_1950);
nor U2274 (N_2274,N_1785,N_1282);
or U2275 (N_2275,N_1167,N_1141);
nand U2276 (N_2276,N_1374,N_1117);
nand U2277 (N_2277,N_1974,N_1458);
nor U2278 (N_2278,N_1607,N_1604);
nor U2279 (N_2279,N_1970,N_1168);
and U2280 (N_2280,N_1483,N_1653);
nand U2281 (N_2281,N_1149,N_1995);
nand U2282 (N_2282,N_1114,N_1330);
nand U2283 (N_2283,N_1817,N_1290);
nor U2284 (N_2284,N_1435,N_1353);
nand U2285 (N_2285,N_1729,N_1155);
or U2286 (N_2286,N_1293,N_1557);
nand U2287 (N_2287,N_1006,N_1043);
or U2288 (N_2288,N_1758,N_1359);
or U2289 (N_2289,N_1133,N_1416);
or U2290 (N_2290,N_1938,N_1352);
nor U2291 (N_2291,N_1915,N_1998);
and U2292 (N_2292,N_1538,N_1945);
and U2293 (N_2293,N_1550,N_1904);
nand U2294 (N_2294,N_1002,N_1792);
nand U2295 (N_2295,N_1961,N_1372);
nand U2296 (N_2296,N_1735,N_1761);
nand U2297 (N_2297,N_1807,N_1140);
nand U2298 (N_2298,N_1929,N_1300);
and U2299 (N_2299,N_1125,N_1437);
nor U2300 (N_2300,N_1160,N_1919);
and U2301 (N_2301,N_1673,N_1854);
and U2302 (N_2302,N_1853,N_1107);
and U2303 (N_2303,N_1189,N_1810);
nor U2304 (N_2304,N_1848,N_1081);
nor U2305 (N_2305,N_1868,N_1916);
nand U2306 (N_2306,N_1473,N_1262);
nand U2307 (N_2307,N_1380,N_1368);
and U2308 (N_2308,N_1093,N_1958);
nand U2309 (N_2309,N_1298,N_1004);
xnor U2310 (N_2310,N_1231,N_1561);
nand U2311 (N_2311,N_1753,N_1296);
nand U2312 (N_2312,N_1824,N_1291);
or U2313 (N_2313,N_1777,N_1599);
and U2314 (N_2314,N_1142,N_1447);
nor U2315 (N_2315,N_1263,N_1899);
or U2316 (N_2316,N_1486,N_1666);
or U2317 (N_2317,N_1558,N_1038);
nor U2318 (N_2318,N_1840,N_1279);
nor U2319 (N_2319,N_1987,N_1455);
nand U2320 (N_2320,N_1378,N_1236);
and U2321 (N_2321,N_1808,N_1151);
or U2322 (N_2322,N_1500,N_1020);
nand U2323 (N_2323,N_1303,N_1990);
xnor U2324 (N_2324,N_1849,N_1415);
nand U2325 (N_2325,N_1238,N_1001);
and U2326 (N_2326,N_1339,N_1205);
nor U2327 (N_2327,N_1413,N_1242);
nor U2328 (N_2328,N_1188,N_1485);
and U2329 (N_2329,N_1623,N_1726);
or U2330 (N_2330,N_1045,N_1575);
and U2331 (N_2331,N_1434,N_1480);
nand U2332 (N_2332,N_1781,N_1948);
or U2333 (N_2333,N_1569,N_1537);
nor U2334 (N_2334,N_1921,N_1776);
and U2335 (N_2335,N_1062,N_1855);
and U2336 (N_2336,N_1837,N_1202);
nand U2337 (N_2337,N_1354,N_1519);
or U2338 (N_2338,N_1939,N_1563);
or U2339 (N_2339,N_1462,N_1556);
or U2340 (N_2340,N_1523,N_1711);
nor U2341 (N_2341,N_1284,N_1815);
or U2342 (N_2342,N_1203,N_1737);
nor U2343 (N_2343,N_1797,N_1039);
or U2344 (N_2344,N_1449,N_1591);
nand U2345 (N_2345,N_1163,N_1076);
nand U2346 (N_2346,N_1740,N_1327);
nand U2347 (N_2347,N_1560,N_1503);
nor U2348 (N_2348,N_1789,N_1838);
or U2349 (N_2349,N_1182,N_1790);
nor U2350 (N_2350,N_1150,N_1402);
or U2351 (N_2351,N_1633,N_1999);
or U2352 (N_2352,N_1684,N_1654);
nand U2353 (N_2353,N_1097,N_1696);
nor U2354 (N_2354,N_1080,N_1267);
and U2355 (N_2355,N_1391,N_1554);
nand U2356 (N_2356,N_1942,N_1541);
and U2357 (N_2357,N_1172,N_1308);
nor U2358 (N_2358,N_1706,N_1943);
nand U2359 (N_2359,N_1658,N_1060);
and U2360 (N_2360,N_1864,N_1635);
and U2361 (N_2361,N_1545,N_1472);
and U2362 (N_2362,N_1430,N_1273);
nand U2363 (N_2363,N_1618,N_1350);
and U2364 (N_2364,N_1928,N_1147);
and U2365 (N_2365,N_1106,N_1305);
and U2366 (N_2366,N_1528,N_1860);
or U2367 (N_2367,N_1126,N_1346);
nor U2368 (N_2368,N_1583,N_1944);
or U2369 (N_2369,N_1791,N_1459);
nand U2370 (N_2370,N_1681,N_1571);
or U2371 (N_2371,N_1504,N_1495);
nor U2372 (N_2372,N_1194,N_1593);
and U2373 (N_2373,N_1540,N_1930);
nand U2374 (N_2374,N_1482,N_1886);
xor U2375 (N_2375,N_1669,N_1686);
or U2376 (N_2376,N_1124,N_1851);
and U2377 (N_2377,N_1258,N_1551);
or U2378 (N_2378,N_1108,N_1896);
and U2379 (N_2379,N_1159,N_1543);
nor U2380 (N_2380,N_1269,N_1779);
and U2381 (N_2381,N_1256,N_1717);
and U2382 (N_2382,N_1702,N_1825);
nor U2383 (N_2383,N_1887,N_1156);
nand U2384 (N_2384,N_1689,N_1547);
nand U2385 (N_2385,N_1880,N_1423);
nand U2386 (N_2386,N_1249,N_1529);
and U2387 (N_2387,N_1549,N_1846);
and U2388 (N_2388,N_1217,N_1268);
or U2389 (N_2389,N_1376,N_1692);
nor U2390 (N_2390,N_1718,N_1349);
and U2391 (N_2391,N_1594,N_1312);
and U2392 (N_2392,N_1253,N_1738);
or U2393 (N_2393,N_1676,N_1390);
and U2394 (N_2394,N_1660,N_1956);
or U2395 (N_2395,N_1951,N_1801);
nand U2396 (N_2396,N_1307,N_1917);
nand U2397 (N_2397,N_1821,N_1014);
nand U2398 (N_2398,N_1085,N_1373);
nor U2399 (N_2399,N_1131,N_1321);
or U2400 (N_2400,N_1509,N_1487);
or U2401 (N_2401,N_1325,N_1872);
or U2402 (N_2402,N_1090,N_1092);
nor U2403 (N_2403,N_1814,N_1091);
and U2404 (N_2404,N_1115,N_1264);
nand U2405 (N_2405,N_1201,N_1088);
and U2406 (N_2406,N_1139,N_1292);
and U2407 (N_2407,N_1257,N_1525);
or U2408 (N_2408,N_1469,N_1337);
nand U2409 (N_2409,N_1910,N_1922);
nand U2410 (N_2410,N_1598,N_1018);
or U2411 (N_2411,N_1451,N_1955);
or U2412 (N_2412,N_1315,N_1611);
or U2413 (N_2413,N_1739,N_1251);
and U2414 (N_2414,N_1869,N_1873);
and U2415 (N_2415,N_1136,N_1122);
or U2416 (N_2416,N_1394,N_1936);
nand U2417 (N_2417,N_1795,N_1823);
nor U2418 (N_2418,N_1281,N_1850);
nor U2419 (N_2419,N_1732,N_1957);
and U2420 (N_2420,N_1208,N_1586);
nand U2421 (N_2421,N_1356,N_1986);
nand U2422 (N_2422,N_1177,N_1903);
nand U2423 (N_2423,N_1634,N_1949);
or U2424 (N_2424,N_1064,N_1072);
nor U2425 (N_2425,N_1542,N_1173);
and U2426 (N_2426,N_1770,N_1759);
or U2427 (N_2427,N_1395,N_1112);
nor U2428 (N_2428,N_1981,N_1120);
nor U2429 (N_2429,N_1322,N_1046);
nor U2430 (N_2430,N_1206,N_1941);
nor U2431 (N_2431,N_1465,N_1960);
nand U2432 (N_2432,N_1959,N_1581);
nand U2433 (N_2433,N_1933,N_1464);
or U2434 (N_2434,N_1709,N_1028);
nor U2435 (N_2435,N_1314,N_1906);
and U2436 (N_2436,N_1619,N_1839);
or U2437 (N_2437,N_1926,N_1227);
nand U2438 (N_2438,N_1474,N_1250);
nand U2439 (N_2439,N_1803,N_1983);
and U2440 (N_2440,N_1224,N_1724);
nor U2441 (N_2441,N_1403,N_1134);
nor U2442 (N_2442,N_1457,N_1275);
nand U2443 (N_2443,N_1183,N_1222);
nor U2444 (N_2444,N_1796,N_1490);
nor U2445 (N_2445,N_1968,N_1914);
nand U2446 (N_2446,N_1925,N_1559);
and U2447 (N_2447,N_1780,N_1813);
or U2448 (N_2448,N_1952,N_1012);
or U2449 (N_2449,N_1083,N_1499);
or U2450 (N_2450,N_1058,N_1652);
or U2451 (N_2451,N_1856,N_1197);
or U2452 (N_2452,N_1098,N_1544);
or U2453 (N_2453,N_1716,N_1865);
or U2454 (N_2454,N_1834,N_1498);
or U2455 (N_2455,N_1467,N_1520);
nand U2456 (N_2456,N_1972,N_1804);
nand U2457 (N_2457,N_1507,N_1967);
nand U2458 (N_2458,N_1025,N_1976);
or U2459 (N_2459,N_1037,N_1680);
and U2460 (N_2460,N_1071,N_1782);
nor U2461 (N_2461,N_1332,N_1572);
xnor U2462 (N_2462,N_1699,N_1662);
or U2463 (N_2463,N_1773,N_1707);
nand U2464 (N_2464,N_1105,N_1663);
or U2465 (N_2465,N_1909,N_1756);
nand U2466 (N_2466,N_1428,N_1845);
nor U2467 (N_2467,N_1646,N_1328);
or U2468 (N_2468,N_1055,N_1678);
or U2469 (N_2469,N_1475,N_1239);
and U2470 (N_2470,N_1397,N_1496);
nand U2471 (N_2471,N_1573,N_1161);
and U2472 (N_2472,N_1742,N_1146);
or U2473 (N_2473,N_1830,N_1468);
nor U2474 (N_2474,N_1369,N_1301);
or U2475 (N_2475,N_1363,N_1488);
and U2476 (N_2476,N_1401,N_1645);
or U2477 (N_2477,N_1389,N_1241);
nor U2478 (N_2478,N_1578,N_1698);
xor U2479 (N_2479,N_1734,N_1907);
nor U2480 (N_2480,N_1820,N_1690);
nor U2481 (N_2481,N_1185,N_1913);
nor U2482 (N_2482,N_1875,N_1109);
nand U2483 (N_2483,N_1649,N_1695);
nand U2484 (N_2484,N_1169,N_1697);
nand U2485 (N_2485,N_1344,N_1011);
and U2486 (N_2486,N_1708,N_1881);
nand U2487 (N_2487,N_1747,N_1535);
or U2488 (N_2488,N_1912,N_1061);
nand U2489 (N_2489,N_1751,N_1700);
and U2490 (N_2490,N_1214,N_1400);
nand U2491 (N_2491,N_1629,N_1318);
nor U2492 (N_2492,N_1111,N_1271);
or U2493 (N_2493,N_1587,N_1918);
nand U2494 (N_2494,N_1871,N_1219);
nor U2495 (N_2495,N_1289,N_1889);
and U2496 (N_2496,N_1546,N_1204);
and U2497 (N_2497,N_1501,N_1323);
and U2498 (N_2498,N_1512,N_1277);
or U2499 (N_2499,N_1506,N_1786);
or U2500 (N_2500,N_1628,N_1426);
or U2501 (N_2501,N_1688,N_1990);
nor U2502 (N_2502,N_1376,N_1506);
nand U2503 (N_2503,N_1434,N_1417);
and U2504 (N_2504,N_1691,N_1434);
nand U2505 (N_2505,N_1406,N_1340);
nand U2506 (N_2506,N_1152,N_1135);
or U2507 (N_2507,N_1239,N_1981);
or U2508 (N_2508,N_1377,N_1960);
and U2509 (N_2509,N_1076,N_1368);
nor U2510 (N_2510,N_1857,N_1660);
nand U2511 (N_2511,N_1642,N_1203);
nor U2512 (N_2512,N_1359,N_1801);
xor U2513 (N_2513,N_1699,N_1526);
nand U2514 (N_2514,N_1770,N_1344);
and U2515 (N_2515,N_1723,N_1904);
nor U2516 (N_2516,N_1498,N_1018);
or U2517 (N_2517,N_1732,N_1390);
nand U2518 (N_2518,N_1302,N_1155);
nand U2519 (N_2519,N_1373,N_1205);
nor U2520 (N_2520,N_1740,N_1697);
nand U2521 (N_2521,N_1083,N_1931);
or U2522 (N_2522,N_1784,N_1939);
nor U2523 (N_2523,N_1925,N_1742);
and U2524 (N_2524,N_1958,N_1504);
and U2525 (N_2525,N_1591,N_1066);
or U2526 (N_2526,N_1209,N_1955);
or U2527 (N_2527,N_1175,N_1831);
and U2528 (N_2528,N_1201,N_1921);
nor U2529 (N_2529,N_1300,N_1731);
nor U2530 (N_2530,N_1748,N_1292);
or U2531 (N_2531,N_1357,N_1016);
or U2532 (N_2532,N_1325,N_1654);
nand U2533 (N_2533,N_1823,N_1852);
xnor U2534 (N_2534,N_1827,N_1617);
or U2535 (N_2535,N_1378,N_1465);
and U2536 (N_2536,N_1161,N_1453);
or U2537 (N_2537,N_1908,N_1732);
and U2538 (N_2538,N_1814,N_1754);
or U2539 (N_2539,N_1959,N_1733);
nor U2540 (N_2540,N_1236,N_1031);
nand U2541 (N_2541,N_1210,N_1541);
nand U2542 (N_2542,N_1379,N_1268);
or U2543 (N_2543,N_1787,N_1961);
or U2544 (N_2544,N_1194,N_1009);
nor U2545 (N_2545,N_1553,N_1412);
nand U2546 (N_2546,N_1680,N_1573);
and U2547 (N_2547,N_1856,N_1731);
nor U2548 (N_2548,N_1763,N_1692);
nor U2549 (N_2549,N_1594,N_1844);
nand U2550 (N_2550,N_1696,N_1559);
xor U2551 (N_2551,N_1061,N_1826);
or U2552 (N_2552,N_1161,N_1731);
or U2553 (N_2553,N_1055,N_1506);
nand U2554 (N_2554,N_1504,N_1518);
nand U2555 (N_2555,N_1517,N_1057);
and U2556 (N_2556,N_1446,N_1927);
nor U2557 (N_2557,N_1837,N_1188);
nor U2558 (N_2558,N_1300,N_1943);
nor U2559 (N_2559,N_1080,N_1140);
or U2560 (N_2560,N_1827,N_1325);
and U2561 (N_2561,N_1089,N_1504);
and U2562 (N_2562,N_1947,N_1198);
nand U2563 (N_2563,N_1974,N_1852);
and U2564 (N_2564,N_1687,N_1846);
nand U2565 (N_2565,N_1370,N_1537);
nor U2566 (N_2566,N_1835,N_1708);
nor U2567 (N_2567,N_1646,N_1001);
xnor U2568 (N_2568,N_1852,N_1563);
and U2569 (N_2569,N_1978,N_1972);
and U2570 (N_2570,N_1874,N_1465);
and U2571 (N_2571,N_1053,N_1584);
or U2572 (N_2572,N_1049,N_1108);
or U2573 (N_2573,N_1472,N_1785);
or U2574 (N_2574,N_1640,N_1062);
or U2575 (N_2575,N_1869,N_1426);
nor U2576 (N_2576,N_1389,N_1937);
or U2577 (N_2577,N_1520,N_1603);
and U2578 (N_2578,N_1261,N_1927);
or U2579 (N_2579,N_1865,N_1588);
nand U2580 (N_2580,N_1987,N_1593);
xnor U2581 (N_2581,N_1515,N_1689);
and U2582 (N_2582,N_1651,N_1793);
nor U2583 (N_2583,N_1099,N_1112);
nor U2584 (N_2584,N_1258,N_1775);
nor U2585 (N_2585,N_1431,N_1463);
nand U2586 (N_2586,N_1355,N_1747);
and U2587 (N_2587,N_1222,N_1147);
nor U2588 (N_2588,N_1815,N_1758);
and U2589 (N_2589,N_1888,N_1906);
nor U2590 (N_2590,N_1317,N_1519);
or U2591 (N_2591,N_1103,N_1111);
and U2592 (N_2592,N_1252,N_1651);
or U2593 (N_2593,N_1723,N_1550);
and U2594 (N_2594,N_1631,N_1275);
nand U2595 (N_2595,N_1860,N_1559);
nand U2596 (N_2596,N_1405,N_1529);
and U2597 (N_2597,N_1792,N_1256);
nand U2598 (N_2598,N_1053,N_1169);
and U2599 (N_2599,N_1967,N_1295);
or U2600 (N_2600,N_1590,N_1354);
nor U2601 (N_2601,N_1598,N_1030);
xnor U2602 (N_2602,N_1010,N_1967);
and U2603 (N_2603,N_1536,N_1152);
nor U2604 (N_2604,N_1104,N_1191);
nand U2605 (N_2605,N_1455,N_1983);
or U2606 (N_2606,N_1370,N_1102);
nand U2607 (N_2607,N_1935,N_1997);
nand U2608 (N_2608,N_1922,N_1875);
and U2609 (N_2609,N_1989,N_1070);
nor U2610 (N_2610,N_1494,N_1566);
nand U2611 (N_2611,N_1459,N_1061);
nor U2612 (N_2612,N_1200,N_1176);
nand U2613 (N_2613,N_1331,N_1018);
or U2614 (N_2614,N_1258,N_1440);
or U2615 (N_2615,N_1928,N_1615);
or U2616 (N_2616,N_1880,N_1722);
nand U2617 (N_2617,N_1047,N_1738);
and U2618 (N_2618,N_1386,N_1320);
and U2619 (N_2619,N_1066,N_1156);
or U2620 (N_2620,N_1836,N_1056);
or U2621 (N_2621,N_1706,N_1445);
and U2622 (N_2622,N_1452,N_1391);
and U2623 (N_2623,N_1884,N_1790);
or U2624 (N_2624,N_1779,N_1541);
nand U2625 (N_2625,N_1352,N_1172);
or U2626 (N_2626,N_1429,N_1599);
nor U2627 (N_2627,N_1846,N_1745);
and U2628 (N_2628,N_1649,N_1444);
nand U2629 (N_2629,N_1853,N_1349);
or U2630 (N_2630,N_1909,N_1461);
and U2631 (N_2631,N_1531,N_1258);
nor U2632 (N_2632,N_1704,N_1055);
nand U2633 (N_2633,N_1519,N_1198);
nand U2634 (N_2634,N_1401,N_1131);
nor U2635 (N_2635,N_1770,N_1351);
and U2636 (N_2636,N_1865,N_1876);
or U2637 (N_2637,N_1069,N_1427);
and U2638 (N_2638,N_1156,N_1890);
or U2639 (N_2639,N_1324,N_1099);
and U2640 (N_2640,N_1167,N_1964);
nor U2641 (N_2641,N_1659,N_1559);
nand U2642 (N_2642,N_1566,N_1035);
or U2643 (N_2643,N_1657,N_1137);
nand U2644 (N_2644,N_1989,N_1563);
xor U2645 (N_2645,N_1790,N_1089);
nand U2646 (N_2646,N_1387,N_1376);
nor U2647 (N_2647,N_1564,N_1734);
or U2648 (N_2648,N_1268,N_1476);
and U2649 (N_2649,N_1886,N_1869);
nand U2650 (N_2650,N_1801,N_1777);
and U2651 (N_2651,N_1247,N_1062);
and U2652 (N_2652,N_1304,N_1414);
nand U2653 (N_2653,N_1254,N_1857);
and U2654 (N_2654,N_1010,N_1239);
nor U2655 (N_2655,N_1439,N_1824);
and U2656 (N_2656,N_1112,N_1399);
nand U2657 (N_2657,N_1968,N_1655);
and U2658 (N_2658,N_1332,N_1752);
and U2659 (N_2659,N_1259,N_1702);
or U2660 (N_2660,N_1794,N_1180);
nand U2661 (N_2661,N_1607,N_1949);
or U2662 (N_2662,N_1792,N_1104);
nor U2663 (N_2663,N_1568,N_1932);
nor U2664 (N_2664,N_1045,N_1734);
and U2665 (N_2665,N_1037,N_1873);
or U2666 (N_2666,N_1880,N_1287);
and U2667 (N_2667,N_1407,N_1273);
or U2668 (N_2668,N_1971,N_1574);
or U2669 (N_2669,N_1372,N_1252);
or U2670 (N_2670,N_1644,N_1859);
and U2671 (N_2671,N_1871,N_1417);
or U2672 (N_2672,N_1294,N_1533);
and U2673 (N_2673,N_1641,N_1555);
or U2674 (N_2674,N_1237,N_1696);
nand U2675 (N_2675,N_1257,N_1589);
or U2676 (N_2676,N_1455,N_1973);
or U2677 (N_2677,N_1757,N_1834);
nand U2678 (N_2678,N_1683,N_1276);
and U2679 (N_2679,N_1618,N_1796);
nor U2680 (N_2680,N_1990,N_1205);
and U2681 (N_2681,N_1243,N_1026);
and U2682 (N_2682,N_1272,N_1183);
nand U2683 (N_2683,N_1556,N_1365);
nand U2684 (N_2684,N_1900,N_1493);
nand U2685 (N_2685,N_1997,N_1168);
and U2686 (N_2686,N_1712,N_1785);
nor U2687 (N_2687,N_1213,N_1311);
nor U2688 (N_2688,N_1567,N_1248);
nand U2689 (N_2689,N_1673,N_1408);
or U2690 (N_2690,N_1272,N_1545);
nor U2691 (N_2691,N_1206,N_1030);
or U2692 (N_2692,N_1231,N_1715);
and U2693 (N_2693,N_1158,N_1810);
nand U2694 (N_2694,N_1598,N_1468);
nand U2695 (N_2695,N_1460,N_1715);
nor U2696 (N_2696,N_1065,N_1807);
or U2697 (N_2697,N_1156,N_1603);
nor U2698 (N_2698,N_1801,N_1572);
or U2699 (N_2699,N_1604,N_1027);
nor U2700 (N_2700,N_1443,N_1197);
nor U2701 (N_2701,N_1237,N_1386);
nand U2702 (N_2702,N_1825,N_1601);
or U2703 (N_2703,N_1039,N_1859);
nand U2704 (N_2704,N_1481,N_1083);
xor U2705 (N_2705,N_1334,N_1897);
nor U2706 (N_2706,N_1165,N_1189);
nand U2707 (N_2707,N_1416,N_1460);
nor U2708 (N_2708,N_1670,N_1320);
nand U2709 (N_2709,N_1945,N_1347);
or U2710 (N_2710,N_1142,N_1847);
nand U2711 (N_2711,N_1871,N_1155);
and U2712 (N_2712,N_1177,N_1880);
nor U2713 (N_2713,N_1668,N_1474);
or U2714 (N_2714,N_1724,N_1843);
nor U2715 (N_2715,N_1431,N_1347);
nand U2716 (N_2716,N_1934,N_1694);
nand U2717 (N_2717,N_1870,N_1889);
and U2718 (N_2718,N_1622,N_1960);
nand U2719 (N_2719,N_1493,N_1592);
nand U2720 (N_2720,N_1554,N_1433);
and U2721 (N_2721,N_1360,N_1346);
or U2722 (N_2722,N_1811,N_1400);
and U2723 (N_2723,N_1631,N_1782);
nor U2724 (N_2724,N_1591,N_1434);
nand U2725 (N_2725,N_1421,N_1328);
nand U2726 (N_2726,N_1335,N_1968);
nand U2727 (N_2727,N_1724,N_1529);
nor U2728 (N_2728,N_1783,N_1040);
and U2729 (N_2729,N_1878,N_1946);
and U2730 (N_2730,N_1770,N_1962);
and U2731 (N_2731,N_1737,N_1657);
and U2732 (N_2732,N_1110,N_1728);
nand U2733 (N_2733,N_1595,N_1966);
nor U2734 (N_2734,N_1035,N_1267);
and U2735 (N_2735,N_1793,N_1596);
nand U2736 (N_2736,N_1320,N_1736);
and U2737 (N_2737,N_1539,N_1392);
nor U2738 (N_2738,N_1077,N_1079);
and U2739 (N_2739,N_1249,N_1038);
nor U2740 (N_2740,N_1700,N_1474);
xnor U2741 (N_2741,N_1276,N_1514);
nand U2742 (N_2742,N_1907,N_1973);
nor U2743 (N_2743,N_1123,N_1158);
or U2744 (N_2744,N_1178,N_1954);
nor U2745 (N_2745,N_1958,N_1967);
or U2746 (N_2746,N_1090,N_1618);
and U2747 (N_2747,N_1402,N_1787);
or U2748 (N_2748,N_1572,N_1046);
nor U2749 (N_2749,N_1354,N_1643);
or U2750 (N_2750,N_1577,N_1671);
nand U2751 (N_2751,N_1406,N_1207);
nand U2752 (N_2752,N_1532,N_1585);
or U2753 (N_2753,N_1525,N_1799);
and U2754 (N_2754,N_1963,N_1429);
or U2755 (N_2755,N_1607,N_1163);
nand U2756 (N_2756,N_1141,N_1697);
nand U2757 (N_2757,N_1290,N_1889);
nand U2758 (N_2758,N_1636,N_1610);
and U2759 (N_2759,N_1750,N_1737);
and U2760 (N_2760,N_1958,N_1111);
and U2761 (N_2761,N_1774,N_1737);
nand U2762 (N_2762,N_1635,N_1163);
nand U2763 (N_2763,N_1087,N_1735);
nor U2764 (N_2764,N_1715,N_1849);
nor U2765 (N_2765,N_1973,N_1394);
nor U2766 (N_2766,N_1266,N_1357);
or U2767 (N_2767,N_1675,N_1332);
and U2768 (N_2768,N_1537,N_1850);
and U2769 (N_2769,N_1776,N_1346);
nor U2770 (N_2770,N_1985,N_1577);
or U2771 (N_2771,N_1196,N_1929);
xor U2772 (N_2772,N_1360,N_1659);
or U2773 (N_2773,N_1214,N_1365);
and U2774 (N_2774,N_1153,N_1888);
nor U2775 (N_2775,N_1129,N_1392);
nand U2776 (N_2776,N_1688,N_1158);
nor U2777 (N_2777,N_1428,N_1741);
nand U2778 (N_2778,N_1966,N_1785);
or U2779 (N_2779,N_1276,N_1910);
nand U2780 (N_2780,N_1182,N_1350);
nor U2781 (N_2781,N_1569,N_1053);
and U2782 (N_2782,N_1686,N_1298);
nor U2783 (N_2783,N_1992,N_1128);
nor U2784 (N_2784,N_1831,N_1510);
or U2785 (N_2785,N_1049,N_1298);
and U2786 (N_2786,N_1181,N_1088);
nor U2787 (N_2787,N_1396,N_1643);
and U2788 (N_2788,N_1160,N_1645);
nand U2789 (N_2789,N_1092,N_1591);
nand U2790 (N_2790,N_1226,N_1031);
nor U2791 (N_2791,N_1595,N_1806);
nand U2792 (N_2792,N_1180,N_1319);
or U2793 (N_2793,N_1157,N_1632);
or U2794 (N_2794,N_1110,N_1131);
nor U2795 (N_2795,N_1400,N_1761);
and U2796 (N_2796,N_1471,N_1103);
nand U2797 (N_2797,N_1298,N_1077);
nand U2798 (N_2798,N_1896,N_1294);
or U2799 (N_2799,N_1684,N_1843);
nand U2800 (N_2800,N_1704,N_1036);
nor U2801 (N_2801,N_1162,N_1133);
and U2802 (N_2802,N_1962,N_1539);
nor U2803 (N_2803,N_1736,N_1960);
nor U2804 (N_2804,N_1372,N_1972);
xor U2805 (N_2805,N_1085,N_1615);
nor U2806 (N_2806,N_1220,N_1060);
nor U2807 (N_2807,N_1582,N_1312);
nor U2808 (N_2808,N_1756,N_1860);
or U2809 (N_2809,N_1707,N_1245);
and U2810 (N_2810,N_1157,N_1934);
nor U2811 (N_2811,N_1933,N_1638);
nand U2812 (N_2812,N_1332,N_1184);
and U2813 (N_2813,N_1421,N_1316);
nand U2814 (N_2814,N_1210,N_1468);
or U2815 (N_2815,N_1072,N_1419);
or U2816 (N_2816,N_1899,N_1154);
nor U2817 (N_2817,N_1176,N_1293);
nor U2818 (N_2818,N_1012,N_1771);
xor U2819 (N_2819,N_1710,N_1210);
and U2820 (N_2820,N_1540,N_1493);
or U2821 (N_2821,N_1919,N_1287);
nor U2822 (N_2822,N_1393,N_1132);
nor U2823 (N_2823,N_1537,N_1651);
nand U2824 (N_2824,N_1039,N_1345);
and U2825 (N_2825,N_1426,N_1661);
or U2826 (N_2826,N_1687,N_1380);
xor U2827 (N_2827,N_1715,N_1305);
and U2828 (N_2828,N_1363,N_1278);
and U2829 (N_2829,N_1274,N_1539);
nand U2830 (N_2830,N_1942,N_1069);
or U2831 (N_2831,N_1391,N_1209);
nor U2832 (N_2832,N_1972,N_1878);
and U2833 (N_2833,N_1478,N_1161);
and U2834 (N_2834,N_1431,N_1686);
and U2835 (N_2835,N_1689,N_1920);
nor U2836 (N_2836,N_1221,N_1770);
nor U2837 (N_2837,N_1928,N_1112);
nor U2838 (N_2838,N_1242,N_1014);
and U2839 (N_2839,N_1773,N_1085);
or U2840 (N_2840,N_1982,N_1730);
nor U2841 (N_2841,N_1262,N_1110);
and U2842 (N_2842,N_1412,N_1715);
xnor U2843 (N_2843,N_1982,N_1058);
or U2844 (N_2844,N_1771,N_1209);
or U2845 (N_2845,N_1706,N_1039);
nor U2846 (N_2846,N_1945,N_1851);
xnor U2847 (N_2847,N_1037,N_1581);
nand U2848 (N_2848,N_1424,N_1832);
nand U2849 (N_2849,N_1918,N_1410);
nor U2850 (N_2850,N_1523,N_1421);
nand U2851 (N_2851,N_1907,N_1622);
nor U2852 (N_2852,N_1552,N_1289);
and U2853 (N_2853,N_1081,N_1047);
nand U2854 (N_2854,N_1204,N_1375);
or U2855 (N_2855,N_1184,N_1786);
nor U2856 (N_2856,N_1369,N_1626);
and U2857 (N_2857,N_1627,N_1651);
nand U2858 (N_2858,N_1054,N_1570);
nand U2859 (N_2859,N_1204,N_1978);
or U2860 (N_2860,N_1600,N_1935);
nand U2861 (N_2861,N_1509,N_1031);
nand U2862 (N_2862,N_1770,N_1543);
nor U2863 (N_2863,N_1683,N_1661);
xnor U2864 (N_2864,N_1400,N_1697);
or U2865 (N_2865,N_1432,N_1664);
nor U2866 (N_2866,N_1285,N_1520);
and U2867 (N_2867,N_1208,N_1955);
or U2868 (N_2868,N_1047,N_1370);
or U2869 (N_2869,N_1625,N_1295);
or U2870 (N_2870,N_1298,N_1844);
or U2871 (N_2871,N_1595,N_1080);
nor U2872 (N_2872,N_1635,N_1189);
nand U2873 (N_2873,N_1090,N_1959);
and U2874 (N_2874,N_1174,N_1718);
nor U2875 (N_2875,N_1174,N_1505);
and U2876 (N_2876,N_1551,N_1869);
and U2877 (N_2877,N_1454,N_1787);
nor U2878 (N_2878,N_1594,N_1623);
nor U2879 (N_2879,N_1452,N_1064);
nand U2880 (N_2880,N_1007,N_1457);
and U2881 (N_2881,N_1983,N_1574);
nor U2882 (N_2882,N_1280,N_1876);
nor U2883 (N_2883,N_1968,N_1547);
nor U2884 (N_2884,N_1681,N_1278);
nand U2885 (N_2885,N_1464,N_1144);
nand U2886 (N_2886,N_1945,N_1978);
or U2887 (N_2887,N_1152,N_1608);
nand U2888 (N_2888,N_1031,N_1793);
or U2889 (N_2889,N_1391,N_1586);
or U2890 (N_2890,N_1087,N_1550);
and U2891 (N_2891,N_1283,N_1000);
or U2892 (N_2892,N_1113,N_1050);
and U2893 (N_2893,N_1128,N_1519);
or U2894 (N_2894,N_1632,N_1623);
nor U2895 (N_2895,N_1176,N_1235);
nand U2896 (N_2896,N_1144,N_1649);
or U2897 (N_2897,N_1863,N_1030);
nand U2898 (N_2898,N_1231,N_1115);
or U2899 (N_2899,N_1476,N_1358);
or U2900 (N_2900,N_1148,N_1189);
and U2901 (N_2901,N_1511,N_1683);
or U2902 (N_2902,N_1200,N_1905);
and U2903 (N_2903,N_1638,N_1401);
nor U2904 (N_2904,N_1954,N_1556);
nor U2905 (N_2905,N_1346,N_1580);
nand U2906 (N_2906,N_1110,N_1433);
nor U2907 (N_2907,N_1928,N_1494);
nor U2908 (N_2908,N_1150,N_1741);
nor U2909 (N_2909,N_1353,N_1510);
nand U2910 (N_2910,N_1292,N_1321);
nor U2911 (N_2911,N_1097,N_1297);
and U2912 (N_2912,N_1498,N_1752);
and U2913 (N_2913,N_1377,N_1844);
nor U2914 (N_2914,N_1068,N_1097);
nand U2915 (N_2915,N_1076,N_1296);
nand U2916 (N_2916,N_1800,N_1879);
and U2917 (N_2917,N_1233,N_1225);
or U2918 (N_2918,N_1279,N_1413);
and U2919 (N_2919,N_1520,N_1054);
or U2920 (N_2920,N_1247,N_1376);
and U2921 (N_2921,N_1942,N_1999);
nand U2922 (N_2922,N_1888,N_1430);
and U2923 (N_2923,N_1344,N_1400);
and U2924 (N_2924,N_1888,N_1351);
and U2925 (N_2925,N_1906,N_1024);
and U2926 (N_2926,N_1652,N_1483);
nand U2927 (N_2927,N_1680,N_1018);
or U2928 (N_2928,N_1512,N_1688);
or U2929 (N_2929,N_1289,N_1219);
nor U2930 (N_2930,N_1587,N_1872);
or U2931 (N_2931,N_1760,N_1109);
and U2932 (N_2932,N_1812,N_1612);
nor U2933 (N_2933,N_1605,N_1962);
and U2934 (N_2934,N_1377,N_1673);
nand U2935 (N_2935,N_1571,N_1797);
nand U2936 (N_2936,N_1977,N_1624);
nand U2937 (N_2937,N_1263,N_1563);
or U2938 (N_2938,N_1464,N_1033);
and U2939 (N_2939,N_1851,N_1183);
and U2940 (N_2940,N_1916,N_1901);
and U2941 (N_2941,N_1746,N_1122);
or U2942 (N_2942,N_1633,N_1362);
nand U2943 (N_2943,N_1583,N_1911);
nor U2944 (N_2944,N_1058,N_1372);
or U2945 (N_2945,N_1561,N_1668);
nor U2946 (N_2946,N_1717,N_1787);
or U2947 (N_2947,N_1584,N_1614);
and U2948 (N_2948,N_1544,N_1762);
nand U2949 (N_2949,N_1131,N_1922);
or U2950 (N_2950,N_1710,N_1725);
nor U2951 (N_2951,N_1583,N_1376);
and U2952 (N_2952,N_1396,N_1191);
nand U2953 (N_2953,N_1828,N_1034);
or U2954 (N_2954,N_1517,N_1525);
or U2955 (N_2955,N_1539,N_1025);
and U2956 (N_2956,N_1023,N_1788);
and U2957 (N_2957,N_1194,N_1074);
nor U2958 (N_2958,N_1016,N_1505);
or U2959 (N_2959,N_1524,N_1241);
and U2960 (N_2960,N_1582,N_1169);
nand U2961 (N_2961,N_1036,N_1143);
and U2962 (N_2962,N_1406,N_1162);
and U2963 (N_2963,N_1516,N_1541);
and U2964 (N_2964,N_1348,N_1808);
or U2965 (N_2965,N_1878,N_1897);
and U2966 (N_2966,N_1077,N_1145);
or U2967 (N_2967,N_1679,N_1273);
and U2968 (N_2968,N_1884,N_1115);
and U2969 (N_2969,N_1728,N_1493);
nor U2970 (N_2970,N_1417,N_1187);
or U2971 (N_2971,N_1357,N_1103);
nor U2972 (N_2972,N_1848,N_1822);
nand U2973 (N_2973,N_1542,N_1480);
or U2974 (N_2974,N_1181,N_1005);
or U2975 (N_2975,N_1435,N_1841);
nand U2976 (N_2976,N_1509,N_1984);
and U2977 (N_2977,N_1338,N_1948);
or U2978 (N_2978,N_1949,N_1809);
and U2979 (N_2979,N_1133,N_1794);
nand U2980 (N_2980,N_1775,N_1435);
and U2981 (N_2981,N_1007,N_1629);
and U2982 (N_2982,N_1639,N_1975);
or U2983 (N_2983,N_1241,N_1438);
nor U2984 (N_2984,N_1097,N_1490);
and U2985 (N_2985,N_1275,N_1921);
nand U2986 (N_2986,N_1390,N_1865);
nand U2987 (N_2987,N_1610,N_1347);
or U2988 (N_2988,N_1266,N_1709);
nand U2989 (N_2989,N_1149,N_1301);
nor U2990 (N_2990,N_1100,N_1039);
and U2991 (N_2991,N_1445,N_1111);
nor U2992 (N_2992,N_1679,N_1784);
or U2993 (N_2993,N_1852,N_1878);
or U2994 (N_2994,N_1517,N_1905);
nand U2995 (N_2995,N_1564,N_1556);
and U2996 (N_2996,N_1326,N_1960);
or U2997 (N_2997,N_1843,N_1719);
or U2998 (N_2998,N_1686,N_1519);
and U2999 (N_2999,N_1235,N_1505);
nand U3000 (N_3000,N_2139,N_2870);
and U3001 (N_3001,N_2938,N_2727);
nor U3002 (N_3002,N_2595,N_2609);
nand U3003 (N_3003,N_2535,N_2022);
and U3004 (N_3004,N_2885,N_2882);
and U3005 (N_3005,N_2538,N_2778);
nor U3006 (N_3006,N_2430,N_2631);
and U3007 (N_3007,N_2165,N_2889);
and U3008 (N_3008,N_2436,N_2724);
nor U3009 (N_3009,N_2438,N_2886);
nor U3010 (N_3010,N_2704,N_2963);
nor U3011 (N_3011,N_2991,N_2834);
nor U3012 (N_3012,N_2844,N_2170);
and U3013 (N_3013,N_2649,N_2426);
or U3014 (N_3014,N_2010,N_2659);
or U3015 (N_3015,N_2157,N_2337);
nand U3016 (N_3016,N_2239,N_2113);
or U3017 (N_3017,N_2909,N_2439);
and U3018 (N_3018,N_2247,N_2057);
and U3019 (N_3019,N_2795,N_2248);
nor U3020 (N_3020,N_2068,N_2894);
or U3021 (N_3021,N_2148,N_2106);
or U3022 (N_3022,N_2543,N_2103);
and U3023 (N_3023,N_2092,N_2335);
nor U3024 (N_3024,N_2959,N_2643);
and U3025 (N_3025,N_2933,N_2446);
nand U3026 (N_3026,N_2822,N_2536);
nand U3027 (N_3027,N_2379,N_2561);
and U3028 (N_3028,N_2389,N_2458);
nor U3029 (N_3029,N_2851,N_2799);
or U3030 (N_3030,N_2982,N_2222);
nor U3031 (N_3031,N_2792,N_2617);
nor U3032 (N_3032,N_2987,N_2890);
nand U3033 (N_3033,N_2108,N_2235);
or U3034 (N_3034,N_2062,N_2739);
nor U3035 (N_3035,N_2860,N_2603);
and U3036 (N_3036,N_2231,N_2677);
nor U3037 (N_3037,N_2114,N_2221);
nand U3038 (N_3038,N_2619,N_2519);
or U3039 (N_3039,N_2474,N_2788);
nor U3040 (N_3040,N_2350,N_2315);
xor U3041 (N_3041,N_2263,N_2797);
or U3042 (N_3042,N_2416,N_2624);
and U3043 (N_3043,N_2391,N_2722);
nor U3044 (N_3044,N_2840,N_2411);
or U3045 (N_3045,N_2490,N_2692);
or U3046 (N_3046,N_2548,N_2947);
nand U3047 (N_3047,N_2550,N_2997);
and U3048 (N_3048,N_2915,N_2555);
and U3049 (N_3049,N_2050,N_2695);
nor U3050 (N_3050,N_2293,N_2489);
nand U3051 (N_3051,N_2485,N_2121);
nor U3052 (N_3052,N_2162,N_2807);
or U3053 (N_3053,N_2751,N_2852);
or U3054 (N_3054,N_2960,N_2793);
nor U3055 (N_3055,N_2151,N_2861);
and U3056 (N_3056,N_2937,N_2819);
nand U3057 (N_3057,N_2185,N_2154);
and U3058 (N_3058,N_2575,N_2848);
nand U3059 (N_3059,N_2591,N_2412);
nor U3060 (N_3060,N_2444,N_2559);
or U3061 (N_3061,N_2770,N_2160);
nand U3062 (N_3062,N_2351,N_2689);
and U3063 (N_3063,N_2499,N_2357);
nand U3064 (N_3064,N_2204,N_2186);
nand U3065 (N_3065,N_2005,N_2829);
nand U3066 (N_3066,N_2912,N_2396);
nor U3067 (N_3067,N_2502,N_2847);
or U3068 (N_3068,N_2081,N_2230);
or U3069 (N_3069,N_2224,N_2195);
nand U3070 (N_3070,N_2283,N_2237);
nand U3071 (N_3071,N_2496,N_2245);
nand U3072 (N_3072,N_2957,N_2642);
and U3073 (N_3073,N_2873,N_2266);
nor U3074 (N_3074,N_2945,N_2850);
nor U3075 (N_3075,N_2598,N_2082);
nor U3076 (N_3076,N_2332,N_2632);
or U3077 (N_3077,N_2791,N_2383);
nand U3078 (N_3078,N_2863,N_2084);
and U3079 (N_3079,N_2137,N_2336);
nor U3080 (N_3080,N_2422,N_2299);
nor U3081 (N_3081,N_2107,N_2680);
nand U3082 (N_3082,N_2817,N_2949);
and U3083 (N_3083,N_2152,N_2064);
nor U3084 (N_3084,N_2765,N_2029);
and U3085 (N_3085,N_2918,N_2355);
and U3086 (N_3086,N_2046,N_2188);
or U3087 (N_3087,N_2942,N_2897);
nand U3088 (N_3088,N_2356,N_2887);
and U3089 (N_3089,N_2639,N_2806);
or U3090 (N_3090,N_2725,N_2986);
nor U3091 (N_3091,N_2405,N_2988);
nand U3092 (N_3092,N_2976,N_2451);
xnor U3093 (N_3093,N_2243,N_2774);
nor U3094 (N_3094,N_2993,N_2922);
nor U3095 (N_3095,N_2600,N_2483);
and U3096 (N_3096,N_2189,N_2066);
or U3097 (N_3097,N_2212,N_2261);
or U3098 (N_3098,N_2480,N_2701);
and U3099 (N_3099,N_2572,N_2839);
and U3100 (N_3100,N_2827,N_2622);
or U3101 (N_3101,N_2524,N_2043);
nand U3102 (N_3102,N_2143,N_2415);
nand U3103 (N_3103,N_2463,N_2265);
or U3104 (N_3104,N_2719,N_2259);
nor U3105 (N_3105,N_2734,N_2091);
nand U3106 (N_3106,N_2373,N_2159);
and U3107 (N_3107,N_2698,N_2130);
nand U3108 (N_3108,N_2638,N_2876);
or U3109 (N_3109,N_2599,N_2175);
and U3110 (N_3110,N_2920,N_2849);
nand U3111 (N_3111,N_2821,N_2891);
xor U3112 (N_3112,N_2833,N_2408);
nor U3113 (N_3113,N_2054,N_2551);
or U3114 (N_3114,N_2295,N_2634);
and U3115 (N_3115,N_2055,N_2205);
nor U3116 (N_3116,N_2290,N_2627);
nor U3117 (N_3117,N_2709,N_2494);
and U3118 (N_3118,N_2517,N_2545);
and U3119 (N_3119,N_2500,N_2941);
nor U3120 (N_3120,N_2635,N_2060);
nand U3121 (N_3121,N_2378,N_2122);
nor U3122 (N_3122,N_2990,N_2690);
and U3123 (N_3123,N_2419,N_2363);
nor U3124 (N_3124,N_2906,N_2999);
nor U3125 (N_3125,N_2961,N_2712);
nand U3126 (N_3126,N_2656,N_2333);
nand U3127 (N_3127,N_2343,N_2823);
or U3128 (N_3128,N_2604,N_2155);
nor U3129 (N_3129,N_2981,N_2174);
nand U3130 (N_3130,N_2164,N_2972);
nor U3131 (N_3131,N_2297,N_2589);
and U3132 (N_3132,N_2470,N_2327);
nand U3133 (N_3133,N_2063,N_2460);
or U3134 (N_3134,N_2488,N_2233);
nor U3135 (N_3135,N_2039,N_2781);
nor U3136 (N_3136,N_2684,N_2220);
and U3137 (N_3137,N_2581,N_2525);
or U3138 (N_3138,N_2662,N_2950);
nand U3139 (N_3139,N_2686,N_2877);
nor U3140 (N_3140,N_2843,N_2073);
or U3141 (N_3141,N_2296,N_2720);
and U3142 (N_3142,N_2520,N_2354);
nand U3143 (N_3143,N_2741,N_2896);
nor U3144 (N_3144,N_2144,N_2199);
or U3145 (N_3145,N_2207,N_2284);
nor U3146 (N_3146,N_2934,N_2418);
nor U3147 (N_3147,N_2880,N_2650);
nand U3148 (N_3148,N_2370,N_2455);
nor U3149 (N_3149,N_2755,N_2994);
and U3150 (N_3150,N_2209,N_2171);
and U3151 (N_3151,N_2557,N_2747);
and U3152 (N_3152,N_2710,N_2161);
or U3153 (N_3153,N_2508,N_2789);
or U3154 (N_3154,N_2443,N_2365);
and U3155 (N_3155,N_2842,N_2256);
nand U3156 (N_3156,N_2948,N_2711);
and U3157 (N_3157,N_2276,N_2726);
or U3158 (N_3158,N_2099,N_2392);
nand U3159 (N_3159,N_2067,N_2413);
nand U3160 (N_3160,N_2738,N_2172);
nand U3161 (N_3161,N_2601,N_2878);
nand U3162 (N_3162,N_2919,N_2069);
and U3163 (N_3163,N_2825,N_2824);
or U3164 (N_3164,N_2750,N_2679);
or U3165 (N_3165,N_2281,N_2448);
and U3166 (N_3166,N_2181,N_2133);
or U3167 (N_3167,N_2729,N_2682);
or U3168 (N_3168,N_2664,N_2895);
or U3169 (N_3169,N_2119,N_2539);
nand U3170 (N_3170,N_2404,N_2226);
nand U3171 (N_3171,N_2621,N_2102);
and U3172 (N_3172,N_2615,N_2045);
and U3173 (N_3173,N_2362,N_2706);
or U3174 (N_3174,N_2298,N_2393);
or U3175 (N_3175,N_2998,N_2964);
or U3176 (N_3176,N_2969,N_2110);
or U3177 (N_3177,N_2104,N_2678);
or U3178 (N_3178,N_2385,N_2759);
and U3179 (N_3179,N_2308,N_2112);
nor U3180 (N_3180,N_2970,N_2124);
nor U3181 (N_3181,N_2374,N_2246);
nor U3182 (N_3182,N_2128,N_2253);
nand U3183 (N_3183,N_2903,N_2504);
or U3184 (N_3184,N_2252,N_2434);
and U3185 (N_3185,N_2407,N_2578);
nand U3186 (N_3186,N_2673,N_2697);
nor U3187 (N_3187,N_2796,N_2316);
nand U3188 (N_3188,N_2040,N_2808);
nor U3189 (N_3189,N_2531,N_2021);
and U3190 (N_3190,N_2648,N_2995);
and U3191 (N_3191,N_2240,N_2614);
nand U3192 (N_3192,N_2790,N_2804);
nor U3193 (N_3193,N_2086,N_2372);
or U3194 (N_3194,N_2482,N_2241);
and U3195 (N_3195,N_2592,N_2280);
and U3196 (N_3196,N_2925,N_2210);
nand U3197 (N_3197,N_2360,N_2244);
nor U3198 (N_3198,N_2930,N_2640);
nor U3199 (N_3199,N_2854,N_2973);
and U3200 (N_3200,N_2492,N_2013);
and U3201 (N_3201,N_2767,N_2567);
and U3202 (N_3202,N_2588,N_2163);
and U3203 (N_3203,N_2657,N_2105);
or U3204 (N_3204,N_2194,N_2071);
nor U3205 (N_3205,N_2566,N_2613);
nor U3206 (N_3206,N_2319,N_2743);
nor U3207 (N_3207,N_2272,N_2579);
nand U3208 (N_3208,N_2397,N_2794);
nor U3209 (N_3209,N_2359,N_2429);
nor U3210 (N_3210,N_2801,N_2707);
nor U3211 (N_3211,N_2893,N_2223);
nor U3212 (N_3212,N_2775,N_2902);
and U3213 (N_3213,N_2138,N_2671);
and U3214 (N_3214,N_2527,N_2249);
nand U3215 (N_3215,N_2503,N_2753);
or U3216 (N_3216,N_2401,N_2708);
nor U3217 (N_3217,N_2730,N_2735);
or U3218 (N_3218,N_2116,N_2117);
nor U3219 (N_3219,N_2493,N_2779);
nand U3220 (N_3220,N_2011,N_2344);
or U3221 (N_3221,N_2236,N_2001);
nor U3222 (N_3222,N_2655,N_2618);
nor U3223 (N_3223,N_2330,N_2254);
nor U3224 (N_3224,N_2688,N_2810);
nand U3225 (N_3225,N_2962,N_2345);
nand U3226 (N_3226,N_2270,N_2556);
nand U3227 (N_3227,N_2544,N_2610);
or U3228 (N_3228,N_2835,N_2452);
nor U3229 (N_3229,N_2685,N_2633);
or U3230 (N_3230,N_2424,N_2399);
nand U3231 (N_3231,N_2660,N_2645);
nor U3232 (N_3232,N_2783,N_2025);
and U3233 (N_3233,N_2658,N_2506);
or U3234 (N_3234,N_2009,N_2065);
and U3235 (N_3235,N_2179,N_2560);
nand U3236 (N_3236,N_2554,N_2958);
nand U3237 (N_3237,N_2654,N_2714);
or U3238 (N_3238,N_2441,N_2070);
nand U3239 (N_3239,N_2892,N_2042);
or U3240 (N_3240,N_2202,N_2331);
or U3241 (N_3241,N_2552,N_2951);
nand U3242 (N_3242,N_2992,N_2868);
and U3243 (N_3243,N_2713,N_2264);
or U3244 (N_3244,N_2167,N_2924);
and U3245 (N_3245,N_2549,N_2715);
nand U3246 (N_3246,N_2038,N_2289);
or U3247 (N_3247,N_2232,N_2927);
nor U3248 (N_3248,N_2929,N_2611);
or U3249 (N_3249,N_2910,N_2647);
or U3250 (N_3250,N_2101,N_2921);
xor U3251 (N_3251,N_2288,N_2899);
nor U3252 (N_3252,N_2364,N_2203);
and U3253 (N_3253,N_2487,N_2014);
or U3254 (N_3254,N_2898,N_2862);
nor U3255 (N_3255,N_2563,N_2190);
nand U3256 (N_3256,N_2523,N_2597);
nand U3257 (N_3257,N_2769,N_2007);
or U3258 (N_3258,N_2433,N_2800);
or U3259 (N_3259,N_2883,N_2558);
and U3260 (N_3260,N_2352,N_2809);
and U3261 (N_3261,N_2637,N_2608);
and U3262 (N_3262,N_2510,N_2653);
nand U3263 (N_3263,N_2278,N_2349);
or U3264 (N_3264,N_2177,N_2300);
or U3265 (N_3265,N_2037,N_2568);
nor U3266 (N_3266,N_2375,N_2376);
and U3267 (N_3267,N_2855,N_2085);
nor U3268 (N_3268,N_2498,N_2571);
nand U3269 (N_3269,N_2590,N_2464);
nand U3270 (N_3270,N_2271,N_2242);
nand U3271 (N_3271,N_2497,N_2462);
nand U3272 (N_3272,N_2745,N_2030);
nand U3273 (N_3273,N_2904,N_2478);
nand U3274 (N_3274,N_2317,N_2716);
and U3275 (N_3275,N_2388,N_2667);
and U3276 (N_3276,N_2017,N_2913);
and U3277 (N_3277,N_2282,N_2307);
nor U3278 (N_3278,N_2465,N_2340);
nand U3279 (N_3279,N_2780,N_2428);
and U3280 (N_3280,N_2310,N_2785);
and U3281 (N_3281,N_2454,N_2140);
and U3282 (N_3282,N_2024,N_2534);
and U3283 (N_3283,N_2100,N_2513);
nor U3284 (N_3284,N_2768,N_2732);
or U3285 (N_3285,N_2573,N_2594);
nor U3286 (N_3286,N_2326,N_2845);
nand U3287 (N_3287,N_2512,N_2234);
or U3288 (N_3288,N_2277,N_2507);
or U3289 (N_3289,N_2200,N_2096);
nor U3290 (N_3290,N_2926,N_2731);
or U3291 (N_3291,N_2314,N_2472);
nand U3292 (N_3292,N_2437,N_2760);
nor U3293 (N_3293,N_2328,N_2742);
or U3294 (N_3294,N_2187,N_2156);
or U3295 (N_3295,N_2865,N_2312);
nand U3296 (N_3296,N_2000,N_2495);
nor U3297 (N_3297,N_2180,N_2127);
nor U3298 (N_3298,N_2219,N_2593);
or U3299 (N_3299,N_2955,N_2358);
or U3300 (N_3300,N_2291,N_2198);
nand U3301 (N_3301,N_2053,N_2320);
nand U3302 (N_3302,N_2888,N_2917);
or U3303 (N_3303,N_2736,N_2700);
nor U3304 (N_3304,N_2079,N_2923);
or U3305 (N_3305,N_2268,N_2518);
nand U3306 (N_3306,N_2620,N_2078);
and U3307 (N_3307,N_2329,N_2943);
and U3308 (N_3308,N_2032,N_2425);
and U3309 (N_3309,N_2953,N_2292);
and U3310 (N_3310,N_2874,N_2574);
nor U3311 (N_3311,N_2041,N_2125);
or U3312 (N_3312,N_2120,N_2651);
nor U3313 (N_3313,N_2182,N_2208);
nor U3314 (N_3314,N_2178,N_2158);
nand U3315 (N_3315,N_2733,N_2002);
nor U3316 (N_3316,N_2744,N_2306);
and U3317 (N_3317,N_2665,N_2059);
nor U3318 (N_3318,N_2456,N_2675);
nand U3319 (N_3319,N_2628,N_2818);
nor U3320 (N_3320,N_2939,N_2145);
nor U3321 (N_3321,N_2353,N_2931);
or U3322 (N_3322,N_2699,N_2968);
or U3323 (N_3323,N_2871,N_2625);
nor U3324 (N_3324,N_2406,N_2696);
nor U3325 (N_3325,N_2322,N_2811);
or U3326 (N_3326,N_2126,N_2872);
and U3327 (N_3327,N_2131,N_2473);
nand U3328 (N_3328,N_2944,N_2914);
nor U3329 (N_3329,N_2864,N_2090);
nand U3330 (N_3330,N_2303,N_2251);
nand U3331 (N_3331,N_2227,N_2900);
nor U3332 (N_3332,N_2176,N_2836);
nand U3333 (N_3333,N_2479,N_2257);
nor U3334 (N_3334,N_2481,N_2989);
and U3335 (N_3335,N_2616,N_2153);
and U3336 (N_3336,N_2582,N_2979);
nand U3337 (N_3337,N_2773,N_2975);
or U3338 (N_3338,N_2260,N_2192);
nand U3339 (N_3339,N_2390,N_2723);
or U3340 (N_3340,N_2048,N_2398);
and U3341 (N_3341,N_2382,N_2533);
or U3342 (N_3342,N_2812,N_2977);
and U3343 (N_3343,N_2605,N_2394);
nand U3344 (N_3344,N_2717,N_2471);
or U3345 (N_3345,N_2229,N_2875);
and U3346 (N_3346,N_2629,N_2787);
nor U3347 (N_3347,N_2761,N_2440);
nor U3348 (N_3348,N_2928,N_2838);
and U3349 (N_3349,N_2771,N_2905);
or U3350 (N_3350,N_2830,N_2748);
and U3351 (N_3351,N_2269,N_2776);
or U3352 (N_3352,N_2476,N_2516);
nor U3353 (N_3353,N_2828,N_2757);
and U3354 (N_3354,N_2400,N_2466);
or U3355 (N_3355,N_2089,N_2772);
nand U3356 (N_3356,N_2028,N_2369);
nor U3357 (N_3357,N_2285,N_2996);
or U3358 (N_3358,N_2974,N_2586);
nand U3359 (N_3359,N_2668,N_2088);
xor U3360 (N_3360,N_2324,N_2623);
and U3361 (N_3361,N_2012,N_2129);
nor U3362 (N_3362,N_2403,N_2841);
nand U3363 (N_3363,N_2342,N_2541);
nor U3364 (N_3364,N_2169,N_2077);
nor U3365 (N_3365,N_2607,N_2134);
nor U3366 (N_3366,N_2644,N_2371);
nor U3367 (N_3367,N_2672,N_2166);
or U3368 (N_3368,N_2967,N_2453);
or U3369 (N_3369,N_2457,N_2368);
and U3370 (N_3370,N_2173,N_2484);
nor U3371 (N_3371,N_2132,N_2703);
and U3372 (N_3372,N_2003,N_2971);
or U3373 (N_3373,N_2076,N_2141);
or U3374 (N_3374,N_2866,N_2047);
or U3375 (N_3375,N_2211,N_2080);
or U3376 (N_3376,N_2530,N_2417);
nor U3377 (N_3377,N_2031,N_2094);
or U3378 (N_3378,N_2565,N_2641);
and U3379 (N_3379,N_2820,N_2669);
nor U3380 (N_3380,N_2409,N_2147);
nor U3381 (N_3381,N_2196,N_2146);
or U3382 (N_3382,N_2072,N_2758);
and U3383 (N_3383,N_2008,N_2526);
nand U3384 (N_3384,N_2238,N_2802);
nor U3385 (N_3385,N_2338,N_2764);
nand U3386 (N_3386,N_2718,N_2683);
nand U3387 (N_3387,N_2983,N_2932);
nor U3388 (N_3388,N_2681,N_2255);
and U3389 (N_3389,N_2274,N_2859);
nor U3390 (N_3390,N_2956,N_2762);
nand U3391 (N_3391,N_2467,N_2505);
nand U3392 (N_3392,N_2846,N_2652);
and U3393 (N_3393,N_2118,N_2213);
and U3394 (N_3394,N_2058,N_2377);
nor U3395 (N_3395,N_2447,N_2461);
and U3396 (N_3396,N_2302,N_2754);
nand U3397 (N_3397,N_2856,N_2435);
nor U3398 (N_3398,N_2115,N_2869);
and U3399 (N_3399,N_2564,N_2075);
xnor U3400 (N_3400,N_2135,N_2035);
or U3401 (N_3401,N_2027,N_2061);
nand U3402 (N_3402,N_2191,N_2149);
or U3403 (N_3403,N_2702,N_2321);
and U3404 (N_3404,N_2168,N_2015);
or U3405 (N_3405,N_2521,N_2334);
nor U3406 (N_3406,N_2432,N_2663);
nand U3407 (N_3407,N_2346,N_2514);
and U3408 (N_3408,N_2410,N_2630);
or U3409 (N_3409,N_2287,N_2313);
nand U3410 (N_3410,N_2311,N_2587);
and U3411 (N_3411,N_2674,N_2570);
and U3412 (N_3412,N_2705,N_2752);
and U3413 (N_3413,N_2074,N_2279);
nor U3414 (N_3414,N_2853,N_2837);
or U3415 (N_3415,N_2273,N_2087);
and U3416 (N_3416,N_2442,N_2056);
and U3417 (N_3417,N_2511,N_2965);
or U3418 (N_3418,N_2217,N_2532);
and U3419 (N_3419,N_2676,N_2946);
nand U3420 (N_3420,N_2911,N_2123);
or U3421 (N_3421,N_2051,N_2509);
nor U3422 (N_3422,N_2380,N_2193);
or U3423 (N_3423,N_2427,N_2916);
nor U3424 (N_3424,N_2262,N_2542);
or U3425 (N_3425,N_2445,N_2515);
nor U3426 (N_3426,N_2309,N_2954);
nand U3427 (N_3427,N_2348,N_2468);
nand U3428 (N_3428,N_2978,N_2936);
nor U3429 (N_3429,N_2867,N_2612);
xor U3430 (N_3430,N_2553,N_2813);
or U3431 (N_3431,N_2402,N_2305);
nand U3432 (N_3432,N_2687,N_2150);
nand U3433 (N_3433,N_2228,N_2966);
nor U3434 (N_3434,N_2201,N_2547);
or U3435 (N_3435,N_2777,N_2583);
and U3436 (N_3436,N_2537,N_2095);
or U3437 (N_3437,N_2183,N_2984);
nor U3438 (N_3438,N_2395,N_2585);
or U3439 (N_3439,N_2339,N_2049);
nor U3440 (N_3440,N_2036,N_2857);
or U3441 (N_3441,N_2626,N_2577);
nor U3442 (N_3442,N_2884,N_2093);
nand U3443 (N_3443,N_2606,N_2477);
nor U3444 (N_3444,N_2475,N_2004);
or U3445 (N_3445,N_2881,N_2033);
nand U3446 (N_3446,N_2044,N_2985);
nor U3447 (N_3447,N_2459,N_2749);
xnor U3448 (N_3448,N_2323,N_2109);
nand U3449 (N_3449,N_2740,N_2216);
and U3450 (N_3450,N_2414,N_2423);
nand U3451 (N_3451,N_2486,N_2798);
and U3452 (N_3452,N_2952,N_2816);
and U3453 (N_3453,N_2301,N_2562);
nor U3454 (N_3454,N_2661,N_2784);
or U3455 (N_3455,N_2501,N_2596);
or U3456 (N_3456,N_2569,N_2026);
or U3457 (N_3457,N_2386,N_2522);
nor U3458 (N_3458,N_2018,N_2214);
nor U3459 (N_3459,N_2670,N_2805);
nand U3460 (N_3460,N_2907,N_2347);
nand U3461 (N_3461,N_2097,N_2052);
nand U3462 (N_3462,N_2020,N_2098);
nor U3463 (N_3463,N_2693,N_2858);
nand U3464 (N_3464,N_2275,N_2826);
or U3465 (N_3465,N_2341,N_2746);
and U3466 (N_3466,N_2366,N_2737);
nor U3467 (N_3467,N_2901,N_2381);
nand U3468 (N_3468,N_2766,N_2361);
nor U3469 (N_3469,N_2294,N_2832);
nand U3470 (N_3470,N_2491,N_2136);
nand U3471 (N_3471,N_2016,N_2763);
and U3472 (N_3472,N_2908,N_2258);
and U3473 (N_3473,N_2387,N_2576);
or U3474 (N_3474,N_2197,N_2646);
nand U3475 (N_3475,N_2529,N_2546);
or U3476 (N_3476,N_2019,N_2286);
nand U3477 (N_3477,N_2721,N_2215);
nand U3478 (N_3478,N_2206,N_2225);
nor U3479 (N_3479,N_2584,N_2602);
and U3480 (N_3480,N_2540,N_2728);
and U3481 (N_3481,N_2666,N_2420);
nor U3482 (N_3482,N_2815,N_2142);
or U3483 (N_3483,N_2782,N_2367);
nand U3484 (N_3484,N_2384,N_2691);
or U3485 (N_3485,N_2184,N_2006);
nand U3486 (N_3486,N_2469,N_2756);
nor U3487 (N_3487,N_2814,N_2935);
nand U3488 (N_3488,N_2218,N_2879);
or U3489 (N_3489,N_2318,N_2449);
or U3490 (N_3490,N_2250,N_2023);
nand U3491 (N_3491,N_2034,N_2267);
nor U3492 (N_3492,N_2528,N_2325);
xor U3493 (N_3493,N_2940,N_2831);
and U3494 (N_3494,N_2304,N_2636);
nor U3495 (N_3495,N_2694,N_2803);
nand U3496 (N_3496,N_2786,N_2421);
and U3497 (N_3497,N_2431,N_2450);
or U3498 (N_3498,N_2083,N_2111);
nor U3499 (N_3499,N_2980,N_2580);
nand U3500 (N_3500,N_2604,N_2313);
nor U3501 (N_3501,N_2636,N_2198);
and U3502 (N_3502,N_2359,N_2948);
and U3503 (N_3503,N_2849,N_2412);
or U3504 (N_3504,N_2084,N_2128);
or U3505 (N_3505,N_2641,N_2290);
or U3506 (N_3506,N_2097,N_2884);
nand U3507 (N_3507,N_2627,N_2034);
or U3508 (N_3508,N_2629,N_2597);
nor U3509 (N_3509,N_2869,N_2579);
and U3510 (N_3510,N_2908,N_2604);
and U3511 (N_3511,N_2218,N_2731);
nor U3512 (N_3512,N_2017,N_2898);
nand U3513 (N_3513,N_2809,N_2059);
and U3514 (N_3514,N_2512,N_2094);
nand U3515 (N_3515,N_2283,N_2558);
nor U3516 (N_3516,N_2768,N_2051);
nand U3517 (N_3517,N_2457,N_2524);
or U3518 (N_3518,N_2154,N_2327);
or U3519 (N_3519,N_2657,N_2065);
nand U3520 (N_3520,N_2231,N_2325);
nand U3521 (N_3521,N_2758,N_2861);
nand U3522 (N_3522,N_2246,N_2154);
nor U3523 (N_3523,N_2214,N_2807);
nand U3524 (N_3524,N_2396,N_2354);
nand U3525 (N_3525,N_2552,N_2888);
nand U3526 (N_3526,N_2063,N_2589);
and U3527 (N_3527,N_2325,N_2611);
or U3528 (N_3528,N_2006,N_2318);
and U3529 (N_3529,N_2968,N_2487);
nand U3530 (N_3530,N_2296,N_2938);
and U3531 (N_3531,N_2570,N_2400);
nand U3532 (N_3532,N_2545,N_2182);
nand U3533 (N_3533,N_2532,N_2318);
and U3534 (N_3534,N_2410,N_2731);
nor U3535 (N_3535,N_2915,N_2252);
or U3536 (N_3536,N_2630,N_2657);
nand U3537 (N_3537,N_2540,N_2455);
nor U3538 (N_3538,N_2724,N_2299);
or U3539 (N_3539,N_2032,N_2766);
or U3540 (N_3540,N_2343,N_2387);
or U3541 (N_3541,N_2588,N_2020);
or U3542 (N_3542,N_2137,N_2238);
nor U3543 (N_3543,N_2725,N_2616);
nor U3544 (N_3544,N_2287,N_2345);
or U3545 (N_3545,N_2574,N_2248);
nor U3546 (N_3546,N_2977,N_2355);
and U3547 (N_3547,N_2023,N_2625);
and U3548 (N_3548,N_2538,N_2676);
and U3549 (N_3549,N_2198,N_2025);
or U3550 (N_3550,N_2279,N_2674);
nand U3551 (N_3551,N_2370,N_2744);
and U3552 (N_3552,N_2244,N_2153);
and U3553 (N_3553,N_2014,N_2040);
nand U3554 (N_3554,N_2154,N_2746);
nor U3555 (N_3555,N_2490,N_2813);
or U3556 (N_3556,N_2401,N_2309);
nand U3557 (N_3557,N_2655,N_2333);
nor U3558 (N_3558,N_2613,N_2746);
and U3559 (N_3559,N_2218,N_2913);
and U3560 (N_3560,N_2100,N_2373);
nand U3561 (N_3561,N_2975,N_2794);
or U3562 (N_3562,N_2221,N_2406);
nand U3563 (N_3563,N_2160,N_2408);
nor U3564 (N_3564,N_2539,N_2343);
or U3565 (N_3565,N_2393,N_2736);
nor U3566 (N_3566,N_2128,N_2052);
or U3567 (N_3567,N_2230,N_2128);
nor U3568 (N_3568,N_2581,N_2357);
nand U3569 (N_3569,N_2110,N_2316);
and U3570 (N_3570,N_2471,N_2288);
or U3571 (N_3571,N_2296,N_2982);
nor U3572 (N_3572,N_2133,N_2533);
or U3573 (N_3573,N_2005,N_2860);
and U3574 (N_3574,N_2713,N_2864);
and U3575 (N_3575,N_2042,N_2543);
nor U3576 (N_3576,N_2016,N_2594);
nand U3577 (N_3577,N_2558,N_2504);
nand U3578 (N_3578,N_2184,N_2777);
nand U3579 (N_3579,N_2214,N_2321);
nor U3580 (N_3580,N_2006,N_2083);
and U3581 (N_3581,N_2841,N_2008);
nor U3582 (N_3582,N_2058,N_2226);
nand U3583 (N_3583,N_2470,N_2607);
nand U3584 (N_3584,N_2169,N_2913);
and U3585 (N_3585,N_2678,N_2153);
or U3586 (N_3586,N_2696,N_2694);
and U3587 (N_3587,N_2723,N_2658);
nor U3588 (N_3588,N_2951,N_2180);
and U3589 (N_3589,N_2028,N_2871);
or U3590 (N_3590,N_2367,N_2604);
or U3591 (N_3591,N_2342,N_2294);
and U3592 (N_3592,N_2216,N_2401);
nor U3593 (N_3593,N_2201,N_2482);
nand U3594 (N_3594,N_2055,N_2922);
nand U3595 (N_3595,N_2984,N_2101);
nor U3596 (N_3596,N_2586,N_2626);
and U3597 (N_3597,N_2808,N_2381);
nor U3598 (N_3598,N_2900,N_2843);
or U3599 (N_3599,N_2202,N_2195);
nor U3600 (N_3600,N_2146,N_2724);
nor U3601 (N_3601,N_2865,N_2622);
nor U3602 (N_3602,N_2009,N_2673);
xnor U3603 (N_3603,N_2769,N_2625);
nand U3604 (N_3604,N_2272,N_2899);
xor U3605 (N_3605,N_2115,N_2062);
nand U3606 (N_3606,N_2897,N_2708);
and U3607 (N_3607,N_2407,N_2327);
or U3608 (N_3608,N_2446,N_2492);
nor U3609 (N_3609,N_2777,N_2046);
and U3610 (N_3610,N_2572,N_2570);
or U3611 (N_3611,N_2849,N_2903);
or U3612 (N_3612,N_2904,N_2235);
or U3613 (N_3613,N_2470,N_2572);
nor U3614 (N_3614,N_2924,N_2078);
and U3615 (N_3615,N_2779,N_2280);
and U3616 (N_3616,N_2542,N_2446);
or U3617 (N_3617,N_2430,N_2743);
nor U3618 (N_3618,N_2077,N_2722);
or U3619 (N_3619,N_2453,N_2355);
and U3620 (N_3620,N_2216,N_2523);
nor U3621 (N_3621,N_2583,N_2134);
and U3622 (N_3622,N_2553,N_2981);
or U3623 (N_3623,N_2968,N_2607);
or U3624 (N_3624,N_2928,N_2619);
nand U3625 (N_3625,N_2144,N_2320);
or U3626 (N_3626,N_2385,N_2313);
nand U3627 (N_3627,N_2515,N_2633);
nand U3628 (N_3628,N_2963,N_2113);
nand U3629 (N_3629,N_2167,N_2259);
nor U3630 (N_3630,N_2455,N_2575);
nor U3631 (N_3631,N_2031,N_2389);
nor U3632 (N_3632,N_2558,N_2866);
nor U3633 (N_3633,N_2366,N_2139);
nor U3634 (N_3634,N_2740,N_2633);
nor U3635 (N_3635,N_2990,N_2353);
nor U3636 (N_3636,N_2767,N_2116);
nand U3637 (N_3637,N_2031,N_2636);
or U3638 (N_3638,N_2527,N_2718);
nor U3639 (N_3639,N_2907,N_2863);
nand U3640 (N_3640,N_2019,N_2457);
nor U3641 (N_3641,N_2251,N_2078);
nor U3642 (N_3642,N_2900,N_2333);
nor U3643 (N_3643,N_2259,N_2964);
nand U3644 (N_3644,N_2434,N_2179);
or U3645 (N_3645,N_2320,N_2899);
or U3646 (N_3646,N_2226,N_2447);
or U3647 (N_3647,N_2731,N_2395);
nor U3648 (N_3648,N_2756,N_2649);
or U3649 (N_3649,N_2329,N_2848);
nand U3650 (N_3650,N_2564,N_2862);
or U3651 (N_3651,N_2139,N_2164);
nor U3652 (N_3652,N_2802,N_2944);
or U3653 (N_3653,N_2413,N_2049);
nor U3654 (N_3654,N_2172,N_2300);
and U3655 (N_3655,N_2570,N_2026);
or U3656 (N_3656,N_2726,N_2141);
nand U3657 (N_3657,N_2718,N_2041);
or U3658 (N_3658,N_2540,N_2535);
or U3659 (N_3659,N_2655,N_2041);
nor U3660 (N_3660,N_2029,N_2012);
and U3661 (N_3661,N_2279,N_2839);
nand U3662 (N_3662,N_2922,N_2348);
and U3663 (N_3663,N_2447,N_2652);
and U3664 (N_3664,N_2413,N_2133);
and U3665 (N_3665,N_2057,N_2185);
nor U3666 (N_3666,N_2102,N_2508);
nand U3667 (N_3667,N_2706,N_2093);
and U3668 (N_3668,N_2984,N_2149);
and U3669 (N_3669,N_2845,N_2969);
or U3670 (N_3670,N_2726,N_2264);
or U3671 (N_3671,N_2200,N_2774);
nor U3672 (N_3672,N_2232,N_2570);
nor U3673 (N_3673,N_2470,N_2263);
and U3674 (N_3674,N_2035,N_2010);
nor U3675 (N_3675,N_2016,N_2819);
nand U3676 (N_3676,N_2307,N_2391);
or U3677 (N_3677,N_2111,N_2997);
nand U3678 (N_3678,N_2900,N_2497);
or U3679 (N_3679,N_2989,N_2242);
and U3680 (N_3680,N_2051,N_2510);
nor U3681 (N_3681,N_2091,N_2819);
or U3682 (N_3682,N_2214,N_2070);
nor U3683 (N_3683,N_2798,N_2445);
or U3684 (N_3684,N_2157,N_2613);
xor U3685 (N_3685,N_2427,N_2261);
or U3686 (N_3686,N_2253,N_2306);
and U3687 (N_3687,N_2104,N_2294);
or U3688 (N_3688,N_2202,N_2396);
nand U3689 (N_3689,N_2997,N_2596);
xnor U3690 (N_3690,N_2884,N_2650);
or U3691 (N_3691,N_2252,N_2678);
nand U3692 (N_3692,N_2877,N_2331);
nor U3693 (N_3693,N_2542,N_2933);
or U3694 (N_3694,N_2538,N_2833);
or U3695 (N_3695,N_2401,N_2964);
nor U3696 (N_3696,N_2647,N_2449);
and U3697 (N_3697,N_2916,N_2110);
or U3698 (N_3698,N_2932,N_2166);
nor U3699 (N_3699,N_2308,N_2685);
and U3700 (N_3700,N_2659,N_2555);
nand U3701 (N_3701,N_2578,N_2719);
nor U3702 (N_3702,N_2683,N_2090);
and U3703 (N_3703,N_2887,N_2365);
nand U3704 (N_3704,N_2339,N_2942);
and U3705 (N_3705,N_2952,N_2418);
or U3706 (N_3706,N_2563,N_2460);
and U3707 (N_3707,N_2915,N_2190);
or U3708 (N_3708,N_2385,N_2510);
or U3709 (N_3709,N_2168,N_2734);
nor U3710 (N_3710,N_2146,N_2432);
xor U3711 (N_3711,N_2855,N_2062);
and U3712 (N_3712,N_2496,N_2910);
or U3713 (N_3713,N_2348,N_2274);
nand U3714 (N_3714,N_2050,N_2250);
or U3715 (N_3715,N_2334,N_2406);
nor U3716 (N_3716,N_2150,N_2546);
nor U3717 (N_3717,N_2140,N_2887);
or U3718 (N_3718,N_2793,N_2890);
nor U3719 (N_3719,N_2300,N_2546);
xor U3720 (N_3720,N_2773,N_2442);
and U3721 (N_3721,N_2470,N_2768);
or U3722 (N_3722,N_2950,N_2806);
xnor U3723 (N_3723,N_2033,N_2549);
nand U3724 (N_3724,N_2753,N_2061);
and U3725 (N_3725,N_2829,N_2813);
or U3726 (N_3726,N_2887,N_2281);
nor U3727 (N_3727,N_2055,N_2451);
nor U3728 (N_3728,N_2023,N_2465);
nand U3729 (N_3729,N_2913,N_2288);
and U3730 (N_3730,N_2706,N_2967);
and U3731 (N_3731,N_2441,N_2253);
or U3732 (N_3732,N_2935,N_2377);
nand U3733 (N_3733,N_2421,N_2510);
nand U3734 (N_3734,N_2029,N_2661);
or U3735 (N_3735,N_2546,N_2871);
nand U3736 (N_3736,N_2659,N_2215);
nor U3737 (N_3737,N_2073,N_2913);
or U3738 (N_3738,N_2492,N_2218);
and U3739 (N_3739,N_2804,N_2448);
nor U3740 (N_3740,N_2717,N_2743);
nand U3741 (N_3741,N_2412,N_2831);
and U3742 (N_3742,N_2445,N_2088);
and U3743 (N_3743,N_2529,N_2028);
nand U3744 (N_3744,N_2626,N_2656);
nand U3745 (N_3745,N_2608,N_2880);
nor U3746 (N_3746,N_2509,N_2527);
and U3747 (N_3747,N_2818,N_2715);
and U3748 (N_3748,N_2775,N_2009);
nor U3749 (N_3749,N_2228,N_2498);
and U3750 (N_3750,N_2252,N_2761);
nor U3751 (N_3751,N_2602,N_2299);
or U3752 (N_3752,N_2186,N_2688);
and U3753 (N_3753,N_2507,N_2743);
and U3754 (N_3754,N_2221,N_2215);
nand U3755 (N_3755,N_2973,N_2032);
nand U3756 (N_3756,N_2065,N_2826);
or U3757 (N_3757,N_2887,N_2820);
nand U3758 (N_3758,N_2382,N_2784);
nor U3759 (N_3759,N_2328,N_2113);
nor U3760 (N_3760,N_2833,N_2051);
or U3761 (N_3761,N_2400,N_2645);
or U3762 (N_3762,N_2591,N_2217);
nor U3763 (N_3763,N_2141,N_2234);
nand U3764 (N_3764,N_2061,N_2157);
or U3765 (N_3765,N_2597,N_2091);
or U3766 (N_3766,N_2054,N_2059);
or U3767 (N_3767,N_2600,N_2614);
and U3768 (N_3768,N_2982,N_2577);
nor U3769 (N_3769,N_2154,N_2040);
nand U3770 (N_3770,N_2650,N_2865);
nor U3771 (N_3771,N_2941,N_2459);
and U3772 (N_3772,N_2836,N_2185);
nand U3773 (N_3773,N_2775,N_2629);
nand U3774 (N_3774,N_2667,N_2617);
and U3775 (N_3775,N_2725,N_2137);
nor U3776 (N_3776,N_2620,N_2233);
and U3777 (N_3777,N_2099,N_2108);
nor U3778 (N_3778,N_2490,N_2633);
or U3779 (N_3779,N_2675,N_2165);
or U3780 (N_3780,N_2153,N_2385);
nand U3781 (N_3781,N_2003,N_2551);
and U3782 (N_3782,N_2182,N_2286);
and U3783 (N_3783,N_2991,N_2343);
and U3784 (N_3784,N_2565,N_2219);
nor U3785 (N_3785,N_2380,N_2173);
or U3786 (N_3786,N_2678,N_2218);
nor U3787 (N_3787,N_2990,N_2006);
and U3788 (N_3788,N_2405,N_2901);
nor U3789 (N_3789,N_2091,N_2068);
nor U3790 (N_3790,N_2536,N_2372);
nand U3791 (N_3791,N_2776,N_2311);
nand U3792 (N_3792,N_2348,N_2856);
nand U3793 (N_3793,N_2016,N_2167);
or U3794 (N_3794,N_2265,N_2501);
or U3795 (N_3795,N_2422,N_2508);
nor U3796 (N_3796,N_2716,N_2565);
nand U3797 (N_3797,N_2423,N_2108);
and U3798 (N_3798,N_2368,N_2751);
nand U3799 (N_3799,N_2181,N_2270);
nand U3800 (N_3800,N_2622,N_2952);
nor U3801 (N_3801,N_2297,N_2346);
nor U3802 (N_3802,N_2594,N_2119);
and U3803 (N_3803,N_2263,N_2705);
xnor U3804 (N_3804,N_2222,N_2206);
and U3805 (N_3805,N_2706,N_2063);
and U3806 (N_3806,N_2475,N_2387);
nand U3807 (N_3807,N_2553,N_2025);
nor U3808 (N_3808,N_2398,N_2404);
nand U3809 (N_3809,N_2935,N_2131);
or U3810 (N_3810,N_2470,N_2296);
nand U3811 (N_3811,N_2942,N_2186);
nand U3812 (N_3812,N_2316,N_2285);
or U3813 (N_3813,N_2739,N_2160);
nor U3814 (N_3814,N_2845,N_2404);
nor U3815 (N_3815,N_2724,N_2660);
nand U3816 (N_3816,N_2858,N_2008);
nor U3817 (N_3817,N_2977,N_2819);
and U3818 (N_3818,N_2760,N_2619);
nor U3819 (N_3819,N_2499,N_2149);
and U3820 (N_3820,N_2807,N_2503);
and U3821 (N_3821,N_2040,N_2531);
or U3822 (N_3822,N_2749,N_2414);
nand U3823 (N_3823,N_2828,N_2482);
and U3824 (N_3824,N_2595,N_2153);
nand U3825 (N_3825,N_2173,N_2654);
nor U3826 (N_3826,N_2282,N_2220);
or U3827 (N_3827,N_2705,N_2250);
or U3828 (N_3828,N_2954,N_2079);
and U3829 (N_3829,N_2028,N_2361);
and U3830 (N_3830,N_2954,N_2927);
nand U3831 (N_3831,N_2061,N_2861);
nor U3832 (N_3832,N_2401,N_2493);
nand U3833 (N_3833,N_2591,N_2576);
nand U3834 (N_3834,N_2799,N_2219);
and U3835 (N_3835,N_2784,N_2609);
and U3836 (N_3836,N_2559,N_2525);
and U3837 (N_3837,N_2181,N_2722);
or U3838 (N_3838,N_2034,N_2961);
and U3839 (N_3839,N_2792,N_2529);
xnor U3840 (N_3840,N_2579,N_2762);
and U3841 (N_3841,N_2430,N_2466);
nand U3842 (N_3842,N_2234,N_2537);
nand U3843 (N_3843,N_2045,N_2208);
nand U3844 (N_3844,N_2955,N_2192);
nand U3845 (N_3845,N_2135,N_2847);
nand U3846 (N_3846,N_2550,N_2965);
or U3847 (N_3847,N_2805,N_2080);
and U3848 (N_3848,N_2736,N_2183);
nor U3849 (N_3849,N_2041,N_2145);
and U3850 (N_3850,N_2716,N_2365);
and U3851 (N_3851,N_2028,N_2225);
and U3852 (N_3852,N_2992,N_2027);
and U3853 (N_3853,N_2519,N_2654);
nand U3854 (N_3854,N_2814,N_2932);
nor U3855 (N_3855,N_2726,N_2088);
and U3856 (N_3856,N_2395,N_2736);
nand U3857 (N_3857,N_2953,N_2241);
or U3858 (N_3858,N_2497,N_2251);
nand U3859 (N_3859,N_2280,N_2117);
nor U3860 (N_3860,N_2970,N_2631);
nor U3861 (N_3861,N_2025,N_2710);
and U3862 (N_3862,N_2521,N_2389);
nand U3863 (N_3863,N_2234,N_2661);
and U3864 (N_3864,N_2310,N_2673);
or U3865 (N_3865,N_2051,N_2754);
and U3866 (N_3866,N_2851,N_2024);
and U3867 (N_3867,N_2224,N_2927);
nand U3868 (N_3868,N_2615,N_2249);
nor U3869 (N_3869,N_2600,N_2085);
nor U3870 (N_3870,N_2489,N_2153);
or U3871 (N_3871,N_2588,N_2659);
nand U3872 (N_3872,N_2886,N_2336);
and U3873 (N_3873,N_2620,N_2467);
nor U3874 (N_3874,N_2953,N_2052);
nor U3875 (N_3875,N_2744,N_2934);
nor U3876 (N_3876,N_2004,N_2045);
and U3877 (N_3877,N_2726,N_2240);
nor U3878 (N_3878,N_2267,N_2640);
nand U3879 (N_3879,N_2037,N_2078);
or U3880 (N_3880,N_2525,N_2777);
and U3881 (N_3881,N_2215,N_2013);
nand U3882 (N_3882,N_2563,N_2462);
and U3883 (N_3883,N_2605,N_2363);
nand U3884 (N_3884,N_2372,N_2017);
and U3885 (N_3885,N_2119,N_2761);
and U3886 (N_3886,N_2545,N_2060);
and U3887 (N_3887,N_2703,N_2896);
nand U3888 (N_3888,N_2564,N_2540);
or U3889 (N_3889,N_2664,N_2066);
and U3890 (N_3890,N_2515,N_2440);
and U3891 (N_3891,N_2072,N_2032);
nand U3892 (N_3892,N_2114,N_2335);
nor U3893 (N_3893,N_2610,N_2079);
and U3894 (N_3894,N_2109,N_2098);
or U3895 (N_3895,N_2094,N_2342);
and U3896 (N_3896,N_2924,N_2397);
nand U3897 (N_3897,N_2701,N_2317);
or U3898 (N_3898,N_2055,N_2525);
or U3899 (N_3899,N_2770,N_2630);
or U3900 (N_3900,N_2429,N_2448);
nor U3901 (N_3901,N_2506,N_2272);
nand U3902 (N_3902,N_2548,N_2260);
and U3903 (N_3903,N_2701,N_2224);
or U3904 (N_3904,N_2014,N_2412);
nand U3905 (N_3905,N_2161,N_2427);
and U3906 (N_3906,N_2240,N_2472);
and U3907 (N_3907,N_2943,N_2227);
nor U3908 (N_3908,N_2137,N_2431);
nand U3909 (N_3909,N_2102,N_2379);
and U3910 (N_3910,N_2085,N_2787);
or U3911 (N_3911,N_2918,N_2406);
and U3912 (N_3912,N_2668,N_2898);
nor U3913 (N_3913,N_2529,N_2471);
nand U3914 (N_3914,N_2142,N_2610);
nor U3915 (N_3915,N_2944,N_2259);
and U3916 (N_3916,N_2339,N_2801);
and U3917 (N_3917,N_2093,N_2878);
nand U3918 (N_3918,N_2131,N_2642);
nand U3919 (N_3919,N_2501,N_2328);
nor U3920 (N_3920,N_2497,N_2846);
nor U3921 (N_3921,N_2822,N_2873);
nand U3922 (N_3922,N_2444,N_2780);
and U3923 (N_3923,N_2094,N_2471);
nand U3924 (N_3924,N_2005,N_2898);
nor U3925 (N_3925,N_2400,N_2381);
or U3926 (N_3926,N_2757,N_2228);
nand U3927 (N_3927,N_2406,N_2408);
and U3928 (N_3928,N_2447,N_2102);
nand U3929 (N_3929,N_2568,N_2462);
nand U3930 (N_3930,N_2539,N_2929);
nor U3931 (N_3931,N_2191,N_2488);
or U3932 (N_3932,N_2008,N_2360);
or U3933 (N_3933,N_2512,N_2206);
and U3934 (N_3934,N_2700,N_2272);
nand U3935 (N_3935,N_2889,N_2073);
nor U3936 (N_3936,N_2970,N_2371);
or U3937 (N_3937,N_2623,N_2812);
and U3938 (N_3938,N_2388,N_2473);
nor U3939 (N_3939,N_2012,N_2485);
nor U3940 (N_3940,N_2158,N_2500);
nor U3941 (N_3941,N_2901,N_2536);
and U3942 (N_3942,N_2653,N_2062);
nand U3943 (N_3943,N_2921,N_2440);
nor U3944 (N_3944,N_2754,N_2047);
nand U3945 (N_3945,N_2143,N_2727);
and U3946 (N_3946,N_2868,N_2016);
or U3947 (N_3947,N_2758,N_2406);
nor U3948 (N_3948,N_2243,N_2841);
nor U3949 (N_3949,N_2268,N_2413);
nor U3950 (N_3950,N_2432,N_2518);
or U3951 (N_3951,N_2851,N_2051);
and U3952 (N_3952,N_2105,N_2110);
nand U3953 (N_3953,N_2430,N_2491);
nor U3954 (N_3954,N_2991,N_2046);
or U3955 (N_3955,N_2962,N_2991);
or U3956 (N_3956,N_2887,N_2512);
or U3957 (N_3957,N_2119,N_2181);
and U3958 (N_3958,N_2350,N_2450);
and U3959 (N_3959,N_2687,N_2651);
nand U3960 (N_3960,N_2779,N_2976);
or U3961 (N_3961,N_2775,N_2207);
and U3962 (N_3962,N_2000,N_2848);
nor U3963 (N_3963,N_2559,N_2887);
nor U3964 (N_3964,N_2348,N_2820);
and U3965 (N_3965,N_2696,N_2935);
or U3966 (N_3966,N_2554,N_2586);
nor U3967 (N_3967,N_2945,N_2691);
nand U3968 (N_3968,N_2456,N_2506);
nand U3969 (N_3969,N_2043,N_2401);
or U3970 (N_3970,N_2185,N_2875);
nand U3971 (N_3971,N_2702,N_2616);
nand U3972 (N_3972,N_2393,N_2825);
and U3973 (N_3973,N_2025,N_2614);
and U3974 (N_3974,N_2606,N_2921);
nand U3975 (N_3975,N_2936,N_2850);
or U3976 (N_3976,N_2030,N_2261);
nor U3977 (N_3977,N_2576,N_2302);
nand U3978 (N_3978,N_2972,N_2819);
or U3979 (N_3979,N_2610,N_2914);
nor U3980 (N_3980,N_2035,N_2419);
xor U3981 (N_3981,N_2601,N_2709);
and U3982 (N_3982,N_2434,N_2663);
and U3983 (N_3983,N_2507,N_2746);
or U3984 (N_3984,N_2259,N_2771);
and U3985 (N_3985,N_2350,N_2352);
nand U3986 (N_3986,N_2910,N_2315);
or U3987 (N_3987,N_2823,N_2945);
or U3988 (N_3988,N_2961,N_2303);
and U3989 (N_3989,N_2550,N_2542);
nand U3990 (N_3990,N_2877,N_2133);
nor U3991 (N_3991,N_2644,N_2655);
nor U3992 (N_3992,N_2221,N_2082);
or U3993 (N_3993,N_2554,N_2160);
nand U3994 (N_3994,N_2566,N_2819);
or U3995 (N_3995,N_2946,N_2644);
nor U3996 (N_3996,N_2153,N_2448);
or U3997 (N_3997,N_2305,N_2462);
or U3998 (N_3998,N_2513,N_2775);
or U3999 (N_3999,N_2765,N_2966);
or U4000 (N_4000,N_3925,N_3160);
nand U4001 (N_4001,N_3518,N_3022);
nor U4002 (N_4002,N_3342,N_3037);
nand U4003 (N_4003,N_3118,N_3275);
nor U4004 (N_4004,N_3384,N_3927);
nor U4005 (N_4005,N_3884,N_3104);
nor U4006 (N_4006,N_3206,N_3476);
or U4007 (N_4007,N_3365,N_3871);
and U4008 (N_4008,N_3759,N_3333);
or U4009 (N_4009,N_3303,N_3242);
nor U4010 (N_4010,N_3486,N_3307);
nor U4011 (N_4011,N_3585,N_3708);
nor U4012 (N_4012,N_3077,N_3785);
nand U4013 (N_4013,N_3842,N_3256);
nand U4014 (N_4014,N_3943,N_3316);
and U4015 (N_4015,N_3914,N_3979);
or U4016 (N_4016,N_3687,N_3562);
or U4017 (N_4017,N_3689,N_3598);
nor U4018 (N_4018,N_3050,N_3377);
and U4019 (N_4019,N_3777,N_3720);
or U4020 (N_4020,N_3341,N_3716);
nor U4021 (N_4021,N_3532,N_3738);
and U4022 (N_4022,N_3591,N_3824);
nand U4023 (N_4023,N_3772,N_3346);
and U4024 (N_4024,N_3641,N_3540);
and U4025 (N_4025,N_3144,N_3690);
and U4026 (N_4026,N_3726,N_3220);
or U4027 (N_4027,N_3051,N_3583);
or U4028 (N_4028,N_3041,N_3143);
and U4029 (N_4029,N_3288,N_3944);
nor U4030 (N_4030,N_3425,N_3002);
nand U4031 (N_4031,N_3178,N_3563);
or U4032 (N_4032,N_3323,N_3547);
nor U4033 (N_4033,N_3645,N_3549);
or U4034 (N_4034,N_3017,N_3685);
nor U4035 (N_4035,N_3565,N_3447);
or U4036 (N_4036,N_3497,N_3360);
nand U4037 (N_4037,N_3858,N_3230);
nor U4038 (N_4038,N_3191,N_3816);
or U4039 (N_4039,N_3968,N_3176);
and U4040 (N_4040,N_3947,N_3446);
and U4041 (N_4041,N_3614,N_3308);
nand U4042 (N_4042,N_3366,N_3055);
and U4043 (N_4043,N_3805,N_3950);
and U4044 (N_4044,N_3203,N_3020);
or U4045 (N_4045,N_3092,N_3564);
nand U4046 (N_4046,N_3804,N_3522);
or U4047 (N_4047,N_3321,N_3949);
and U4048 (N_4048,N_3659,N_3875);
or U4049 (N_4049,N_3599,N_3814);
nand U4050 (N_4050,N_3813,N_3309);
or U4051 (N_4051,N_3237,N_3452);
nand U4052 (N_4052,N_3615,N_3215);
nor U4053 (N_4053,N_3015,N_3821);
nand U4054 (N_4054,N_3427,N_3966);
nand U4055 (N_4055,N_3932,N_3196);
or U4056 (N_4056,N_3795,N_3844);
or U4057 (N_4057,N_3586,N_3000);
nor U4058 (N_4058,N_3571,N_3646);
or U4059 (N_4059,N_3657,N_3195);
or U4060 (N_4060,N_3848,N_3575);
and U4061 (N_4061,N_3045,N_3800);
and U4062 (N_4062,N_3998,N_3003);
nand U4063 (N_4063,N_3329,N_3713);
and U4064 (N_4064,N_3379,N_3808);
and U4065 (N_4065,N_3100,N_3721);
nor U4066 (N_4066,N_3747,N_3453);
and U4067 (N_4067,N_3246,N_3724);
or U4068 (N_4068,N_3854,N_3349);
nor U4069 (N_4069,N_3538,N_3515);
nor U4070 (N_4070,N_3737,N_3182);
and U4071 (N_4071,N_3851,N_3873);
nand U4072 (N_4072,N_3027,N_3535);
or U4073 (N_4073,N_3809,N_3415);
nor U4074 (N_4074,N_3146,N_3347);
or U4075 (N_4075,N_3697,N_3324);
or U4076 (N_4076,N_3782,N_3783);
nor U4077 (N_4077,N_3424,N_3976);
nand U4078 (N_4078,N_3674,N_3617);
xnor U4079 (N_4079,N_3572,N_3487);
nor U4080 (N_4080,N_3779,N_3484);
and U4081 (N_4081,N_3358,N_3650);
or U4082 (N_4082,N_3883,N_3870);
nand U4083 (N_4083,N_3581,N_3728);
nor U4084 (N_4084,N_3098,N_3139);
and U4085 (N_4085,N_3802,N_3197);
or U4086 (N_4086,N_3960,N_3744);
nor U4087 (N_4087,N_3555,N_3397);
or U4088 (N_4088,N_3008,N_3985);
nor U4089 (N_4089,N_3315,N_3493);
and U4090 (N_4090,N_3062,N_3418);
nand U4091 (N_4091,N_3394,N_3988);
nand U4092 (N_4092,N_3202,N_3908);
and U4093 (N_4093,N_3428,N_3837);
nand U4094 (N_4094,N_3268,N_3573);
nor U4095 (N_4095,N_3414,N_3924);
nand U4096 (N_4096,N_3669,N_3499);
or U4097 (N_4097,N_3910,N_3495);
nor U4098 (N_4098,N_3221,N_3590);
or U4099 (N_4099,N_3149,N_3094);
nor U4100 (N_4100,N_3161,N_3730);
or U4101 (N_4101,N_3198,N_3337);
nand U4102 (N_4102,N_3336,N_3917);
nor U4103 (N_4103,N_3167,N_3007);
nor U4104 (N_4104,N_3776,N_3594);
nor U4105 (N_4105,N_3370,N_3683);
nand U4106 (N_4106,N_3663,N_3205);
or U4107 (N_4107,N_3480,N_3073);
and U4108 (N_4108,N_3760,N_3520);
nor U4109 (N_4109,N_3799,N_3047);
and U4110 (N_4110,N_3439,N_3469);
or U4111 (N_4111,N_3845,N_3638);
nand U4112 (N_4112,N_3505,N_3667);
and U4113 (N_4113,N_3087,N_3292);
or U4114 (N_4114,N_3529,N_3939);
and U4115 (N_4115,N_3566,N_3934);
nor U4116 (N_4116,N_3417,N_3725);
nand U4117 (N_4117,N_3403,N_3074);
or U4118 (N_4118,N_3817,N_3318);
and U4119 (N_4119,N_3951,N_3931);
and U4120 (N_4120,N_3192,N_3916);
and U4121 (N_4121,N_3209,N_3356);
or U4122 (N_4122,N_3879,N_3955);
nand U4123 (N_4123,N_3963,N_3853);
and U4124 (N_4124,N_3570,N_3135);
or U4125 (N_4125,N_3554,N_3559);
nand U4126 (N_4126,N_3832,N_3282);
nand U4127 (N_4127,N_3742,N_3579);
or U4128 (N_4128,N_3746,N_3300);
and U4129 (N_4129,N_3671,N_3684);
nand U4130 (N_4130,N_3761,N_3830);
or U4131 (N_4131,N_3970,N_3605);
nor U4132 (N_4132,N_3444,N_3408);
or U4133 (N_4133,N_3420,N_3694);
and U4134 (N_4134,N_3576,N_3913);
nand U4135 (N_4135,N_3796,N_3023);
nor U4136 (N_4136,N_3361,N_3232);
nand U4137 (N_4137,N_3276,N_3390);
or U4138 (N_4138,N_3431,N_3102);
nor U4139 (N_4139,N_3185,N_3629);
and U4140 (N_4140,N_3676,N_3700);
nand U4141 (N_4141,N_3903,N_3981);
nor U4142 (N_4142,N_3065,N_3362);
xor U4143 (N_4143,N_3281,N_3291);
and U4144 (N_4144,N_3691,N_3699);
or U4145 (N_4145,N_3501,N_3926);
or U4146 (N_4146,N_3409,N_3274);
nand U4147 (N_4147,N_3537,N_3636);
nor U4148 (N_4148,N_3407,N_3882);
or U4149 (N_4149,N_3187,N_3236);
nor U4150 (N_4150,N_3293,N_3727);
or U4151 (N_4151,N_3899,N_3836);
nand U4152 (N_4152,N_3901,N_3014);
nor U4153 (N_4153,N_3075,N_3709);
nor U4154 (N_4154,N_3359,N_3267);
nor U4155 (N_4155,N_3284,N_3923);
and U4156 (N_4156,N_3625,N_3227);
and U4157 (N_4157,N_3214,N_3113);
and U4158 (N_4158,N_3364,N_3895);
nand U4159 (N_4159,N_3582,N_3516);
nand U4160 (N_4160,N_3855,N_3749);
or U4161 (N_4161,N_3496,N_3768);
nor U4162 (N_4162,N_3775,N_3885);
nand U4163 (N_4163,N_3297,N_3498);
and U4164 (N_4164,N_3387,N_3603);
or U4165 (N_4165,N_3272,N_3611);
or U4166 (N_4166,N_3353,N_3306);
nor U4167 (N_4167,N_3886,N_3770);
nand U4168 (N_4168,N_3399,N_3867);
and U4169 (N_4169,N_3440,N_3794);
nand U4170 (N_4170,N_3219,N_3517);
nor U4171 (N_4171,N_3054,N_3299);
xnor U4172 (N_4172,N_3894,N_3595);
nor U4173 (N_4173,N_3208,N_3376);
nor U4174 (N_4174,N_3791,N_3652);
nand U4175 (N_4175,N_3437,N_3451);
nand U4176 (N_4176,N_3183,N_3642);
nand U4177 (N_4177,N_3071,N_3896);
nand U4178 (N_4178,N_3878,N_3287);
nand U4179 (N_4179,N_3758,N_3490);
nor U4180 (N_4180,N_3577,N_3980);
nor U4181 (N_4181,N_3890,N_3477);
nand U4182 (N_4182,N_3504,N_3545);
nand U4183 (N_4183,N_3097,N_3637);
and U4184 (N_4184,N_3632,N_3864);
and U4185 (N_4185,N_3238,N_3217);
and U4186 (N_4186,N_3673,N_3345);
nor U4187 (N_4187,N_3166,N_3722);
and U4188 (N_4188,N_3240,N_3393);
and U4189 (N_4189,N_3874,N_3371);
nand U4190 (N_4190,N_3588,N_3600);
nor U4191 (N_4191,N_3235,N_3168);
nand U4192 (N_4192,N_3525,N_3987);
nor U4193 (N_4193,N_3500,N_3259);
or U4194 (N_4194,N_3004,N_3462);
or U4195 (N_4195,N_3269,N_3952);
or U4196 (N_4196,N_3546,N_3946);
nand U4197 (N_4197,N_3429,N_3921);
and U4198 (N_4198,N_3177,N_3126);
and U4199 (N_4199,N_3343,N_3954);
and U4200 (N_4200,N_3790,N_3682);
and U4201 (N_4201,N_3430,N_3865);
or U4202 (N_4202,N_3466,N_3843);
nor U4203 (N_4203,N_3624,N_3450);
nand U4204 (N_4204,N_3148,N_3762);
and U4205 (N_4205,N_3378,N_3159);
nand U4206 (N_4206,N_3911,N_3031);
and U4207 (N_4207,N_3029,N_3681);
nor U4208 (N_4208,N_3155,N_3717);
nand U4209 (N_4209,N_3491,N_3807);
nor U4210 (N_4210,N_3043,N_3862);
and U4211 (N_4211,N_3613,N_3186);
and U4212 (N_4212,N_3257,N_3654);
nand U4213 (N_4213,N_3088,N_3038);
or U4214 (N_4214,N_3357,N_3511);
nor U4215 (N_4215,N_3769,N_3763);
and U4216 (N_4216,N_3578,N_3422);
nand U4217 (N_4217,N_3834,N_3188);
nor U4218 (N_4218,N_3906,N_3295);
and U4219 (N_4219,N_3369,N_3125);
and U4220 (N_4220,N_3999,N_3052);
or U4221 (N_4221,N_3124,N_3648);
nand U4222 (N_4222,N_3852,N_3695);
nor U4223 (N_4223,N_3290,N_3766);
or U4224 (N_4224,N_3997,N_3258);
or U4225 (N_4225,N_3140,N_3607);
or U4226 (N_4226,N_3819,N_3551);
nand U4227 (N_4227,N_3441,N_3294);
and U4228 (N_4228,N_3892,N_3640);
and U4229 (N_4229,N_3829,N_3596);
nand U4230 (N_4230,N_3473,N_3286);
nand U4231 (N_4231,N_3898,N_3175);
nand U4232 (N_4232,N_3330,N_3122);
nor U4233 (N_4233,N_3211,N_3035);
nor U4234 (N_4234,N_3482,N_3692);
or U4235 (N_4235,N_3610,N_3465);
or U4236 (N_4236,N_3907,N_3229);
nand U4237 (N_4237,N_3335,N_3823);
nor U4238 (N_4238,N_3539,N_3711);
and U4239 (N_4239,N_3273,N_3655);
nand U4240 (N_4240,N_3134,N_3996);
nor U4241 (N_4241,N_3344,N_3492);
nor U4242 (N_4242,N_3079,N_3902);
or U4243 (N_4243,N_3162,N_3693);
nand U4244 (N_4244,N_3169,N_3391);
nand U4245 (N_4245,N_3995,N_3093);
nor U4246 (N_4246,N_3631,N_3410);
nand U4247 (N_4247,N_3705,N_3787);
or U4248 (N_4248,N_3567,N_3680);
and U4249 (N_4249,N_3519,N_3994);
and U4250 (N_4250,N_3277,N_3305);
nand U4251 (N_4251,N_3869,N_3589);
nor U4252 (N_4252,N_3859,N_3158);
or U4253 (N_4253,N_3082,N_3510);
or U4254 (N_4254,N_3833,N_3459);
nor U4255 (N_4255,N_3173,N_3184);
or U4256 (N_4256,N_3506,N_3877);
nor U4257 (N_4257,N_3745,N_3481);
nand U4258 (N_4258,N_3301,N_3618);
nor U4259 (N_4259,N_3455,N_3698);
or U4260 (N_4260,N_3470,N_3973);
nand U4261 (N_4261,N_3580,N_3702);
or U4262 (N_4262,N_3993,N_3992);
nor U4263 (N_4263,N_3351,N_3249);
or U4264 (N_4264,N_3304,N_3413);
nor U4265 (N_4265,N_3165,N_3552);
or U4266 (N_4266,N_3978,N_3507);
nand U4267 (N_4267,N_3253,N_3531);
or U4268 (N_4268,N_3331,N_3320);
nor U4269 (N_4269,N_3085,N_3263);
and U4270 (N_4270,N_3889,N_3942);
and U4271 (N_4271,N_3233,N_3013);
and U4272 (N_4272,N_3544,N_3406);
nor U4273 (N_4273,N_3556,N_3279);
nor U4274 (N_4274,N_3780,N_3568);
nor U4275 (N_4275,N_3774,N_3792);
and U4276 (N_4276,N_3123,N_3326);
nand U4277 (N_4277,N_3773,N_3255);
or U4278 (N_4278,N_3385,N_3325);
nor U4279 (N_4279,N_3355,N_3781);
nand U4280 (N_4280,N_3154,N_3587);
nor U4281 (N_4281,N_3592,N_3656);
xnor U4282 (N_4282,N_3317,N_3449);
nor U4283 (N_4283,N_3574,N_3820);
nor U4284 (N_4284,N_3664,N_3753);
or U4285 (N_4285,N_3512,N_3915);
nand U4286 (N_4286,N_3956,N_3389);
or U4287 (N_4287,N_3145,N_3432);
and U4288 (N_4288,N_3207,N_3332);
nor U4289 (N_4289,N_3984,N_3034);
nor U4290 (N_4290,N_3179,N_3076);
and U4291 (N_4291,N_3260,N_3084);
or U4292 (N_4292,N_3643,N_3006);
nand U4293 (N_4293,N_3339,N_3937);
nand U4294 (N_4294,N_3086,N_3271);
and U4295 (N_4295,N_3953,N_3620);
nand U4296 (N_4296,N_3941,N_3658);
nand U4297 (N_4297,N_3478,N_3223);
nand U4298 (N_4298,N_3436,N_3735);
nor U4299 (N_4299,N_3971,N_3081);
or U4300 (N_4300,N_3660,N_3091);
or U4301 (N_4301,N_3189,N_3338);
and U4302 (N_4302,N_3718,N_3103);
nand U4303 (N_4303,N_3767,N_3311);
nor U4304 (N_4304,N_3751,N_3801);
nand U4305 (N_4305,N_3280,N_3053);
nand U4306 (N_4306,N_3553,N_3847);
and U4307 (N_4307,N_3701,N_3411);
nor U4308 (N_4308,N_3936,N_3030);
or U4309 (N_4309,N_3627,N_3063);
and U4310 (N_4310,N_3064,N_3975);
or U4311 (N_4311,N_3703,N_3108);
or U4312 (N_4312,N_3039,N_3181);
nand U4313 (N_4313,N_3533,N_3929);
and U4314 (N_4314,N_3967,N_3193);
nand U4315 (N_4315,N_3129,N_3969);
nor U4316 (N_4316,N_3046,N_3130);
or U4317 (N_4317,N_3856,N_3435);
or U4318 (N_4318,N_3635,N_3628);
and U4319 (N_4319,N_3616,N_3241);
and U4320 (N_4320,N_3141,N_3514);
nor U4321 (N_4321,N_3322,N_3897);
or U4322 (N_4322,N_3653,N_3509);
nand U4323 (N_4323,N_3826,N_3314);
nand U4324 (N_4324,N_3340,N_3026);
nor U4325 (N_4325,N_3841,N_3560);
or U4326 (N_4326,N_3024,N_3171);
nor U4327 (N_4327,N_3741,N_3835);
and U4328 (N_4328,N_3521,N_3388);
nand U4329 (N_4329,N_3639,N_3948);
nand U4330 (N_4330,N_3840,N_3058);
or U4331 (N_4331,N_3392,N_3788);
or U4332 (N_4332,N_3127,N_3040);
and U4333 (N_4333,N_3959,N_3244);
and U4334 (N_4334,N_3793,N_3049);
or U4335 (N_4335,N_3938,N_3900);
xnor U4336 (N_4336,N_3128,N_3649);
or U4337 (N_4337,N_3021,N_3789);
nand U4338 (N_4338,N_3468,N_3479);
nor U4339 (N_4339,N_3119,N_3803);
and U4340 (N_4340,N_3502,N_3661);
and U4341 (N_4341,N_3743,N_3597);
or U4342 (N_4342,N_3243,N_3412);
or U4343 (N_4343,N_3715,N_3398);
and U4344 (N_4344,N_3986,N_3991);
nor U4345 (N_4345,N_3608,N_3604);
nand U4346 (N_4346,N_3421,N_3472);
nor U4347 (N_4347,N_3212,N_3457);
or U4348 (N_4348,N_3454,N_3752);
nand U4349 (N_4349,N_3099,N_3381);
nand U4350 (N_4350,N_3584,N_3163);
or U4351 (N_4351,N_3606,N_3120);
nand U4352 (N_4352,N_3541,N_3142);
and U4353 (N_4353,N_3350,N_3612);
nand U4354 (N_4354,N_3434,N_3423);
and U4355 (N_4355,N_3839,N_3822);
and U4356 (N_4356,N_3044,N_3352);
nand U4357 (N_4357,N_3524,N_3234);
or U4358 (N_4358,N_3106,N_3677);
and U4359 (N_4359,N_3312,N_3872);
or U4360 (N_4360,N_3536,N_3534);
or U4361 (N_4361,N_3278,N_3732);
nand U4362 (N_4362,N_3334,N_3526);
nand U4363 (N_4363,N_3962,N_3157);
and U4364 (N_4364,N_3982,N_3957);
or U4365 (N_4365,N_3778,N_3474);
nor U4366 (N_4366,N_3156,N_3433);
or U4367 (N_4367,N_3644,N_3488);
and U4368 (N_4368,N_3066,N_3989);
nand U4369 (N_4369,N_3107,N_3368);
nand U4370 (N_4370,N_3172,N_3012);
or U4371 (N_4371,N_3857,N_3302);
and U4372 (N_4372,N_3386,N_3868);
nand U4373 (N_4373,N_3806,N_3239);
nor U4374 (N_4374,N_3266,N_3630);
and U4375 (N_4375,N_3283,N_3619);
nor U4376 (N_4376,N_3527,N_3252);
and U4377 (N_4377,N_3367,N_3251);
nor U4378 (N_4378,N_3204,N_3213);
nor U4379 (N_4379,N_3489,N_3310);
nand U4380 (N_4380,N_3666,N_3327);
nand U4381 (N_4381,N_3110,N_3216);
or U4382 (N_4382,N_3080,N_3601);
and U4383 (N_4383,N_3089,N_3009);
or U4384 (N_4384,N_3067,N_3416);
or U4385 (N_4385,N_3111,N_3731);
nor U4386 (N_4386,N_3372,N_3032);
and U4387 (N_4387,N_3494,N_3609);
or U4388 (N_4388,N_3602,N_3891);
or U4389 (N_4389,N_3033,N_3706);
or U4390 (N_4390,N_3861,N_3461);
and U4391 (N_4391,N_3548,N_3114);
nor U4392 (N_4392,N_3210,N_3756);
nor U4393 (N_4393,N_3222,N_3152);
and U4394 (N_4394,N_3750,N_3710);
or U4395 (N_4395,N_3112,N_3402);
nand U4396 (N_4396,N_3748,N_3247);
nor U4397 (N_4397,N_3068,N_3958);
nand U4398 (N_4398,N_3827,N_3729);
or U4399 (N_4399,N_3150,N_3419);
and U4400 (N_4400,N_3056,N_3117);
nand U4401 (N_4401,N_3245,N_3136);
nand U4402 (N_4402,N_3483,N_3797);
nand U4403 (N_4403,N_3057,N_3974);
nor U4404 (N_4404,N_3755,N_3719);
or U4405 (N_4405,N_3964,N_3704);
nand U4406 (N_4406,N_3115,N_3438);
nor U4407 (N_4407,N_3289,N_3825);
nand U4408 (N_4408,N_3933,N_3734);
nand U4409 (N_4409,N_3712,N_3881);
or U4410 (N_4410,N_3460,N_3194);
or U4411 (N_4411,N_3626,N_3059);
and U4412 (N_4412,N_3131,N_3250);
nor U4413 (N_4413,N_3593,N_3811);
or U4414 (N_4414,N_3672,N_3860);
and U4415 (N_4415,N_3918,N_3313);
or U4416 (N_4416,N_3016,N_3116);
or U4417 (N_4417,N_3296,N_3733);
and U4418 (N_4418,N_3714,N_3662);
nor U4419 (N_4419,N_3736,N_3863);
nor U4420 (N_4420,N_3199,N_3228);
and U4421 (N_4421,N_3200,N_3838);
or U4422 (N_4422,N_3010,N_3011);
and U4423 (N_4423,N_3262,N_3828);
and U4424 (N_4424,N_3090,N_3651);
nor U4425 (N_4425,N_3442,N_3138);
and U4426 (N_4426,N_3018,N_3226);
nand U4427 (N_4427,N_3072,N_3771);
and U4428 (N_4428,N_3543,N_3265);
and U4429 (N_4429,N_3443,N_3880);
nand U4430 (N_4430,N_3678,N_3105);
nor U4431 (N_4431,N_3668,N_3445);
nor U4432 (N_4432,N_3723,N_3405);
nor U4433 (N_4433,N_3190,N_3784);
nor U4434 (N_4434,N_3048,N_3569);
nor U4435 (N_4435,N_3815,N_3675);
nor U4436 (N_4436,N_3354,N_3147);
and U4437 (N_4437,N_3375,N_3005);
nand U4438 (N_4438,N_3707,N_3961);
or U4439 (N_4439,N_3757,N_3503);
nand U4440 (N_4440,N_3928,N_3557);
or U4441 (N_4441,N_3151,N_3078);
or U4442 (N_4442,N_3254,N_3095);
nor U4443 (N_4443,N_3866,N_3328);
or U4444 (N_4444,N_3464,N_3688);
nor U4445 (N_4445,N_3634,N_3218);
nor U4446 (N_4446,N_3542,N_3972);
and U4447 (N_4447,N_3754,N_3849);
and U4448 (N_4448,N_3132,N_3919);
nor U4449 (N_4449,N_3550,N_3764);
nor U4450 (N_4450,N_3270,N_3264);
or U4451 (N_4451,N_3096,N_3633);
nor U4452 (N_4452,N_3623,N_3170);
and U4453 (N_4453,N_3621,N_3940);
nor U4454 (N_4454,N_3888,N_3887);
and U4455 (N_4455,N_3028,N_3383);
or U4456 (N_4456,N_3528,N_3285);
nor U4457 (N_4457,N_3558,N_3810);
and U4458 (N_4458,N_3109,N_3448);
and U4459 (N_4459,N_3133,N_3201);
nand U4460 (N_4460,N_3922,N_3812);
nor U4461 (N_4461,N_3225,N_3467);
or U4462 (N_4462,N_3083,N_3846);
nand U4463 (N_4463,N_3164,N_3930);
nand U4464 (N_4464,N_3458,N_3101);
nor U4465 (N_4465,N_3380,N_3686);
nand U4466 (N_4466,N_3909,N_3523);
nand U4467 (N_4467,N_3456,N_3121);
nor U4468 (N_4468,N_3508,N_3025);
nor U4469 (N_4469,N_3530,N_3647);
or U4470 (N_4470,N_3475,N_3739);
or U4471 (N_4471,N_3679,N_3471);
nor U4472 (N_4472,N_3153,N_3396);
nor U4473 (N_4473,N_3180,N_3893);
and U4474 (N_4474,N_3670,N_3001);
nor U4475 (N_4475,N_3060,N_3400);
nor U4476 (N_4476,N_3818,N_3363);
nand U4477 (N_4477,N_3561,N_3248);
nand U4478 (N_4478,N_3036,N_3401);
and U4479 (N_4479,N_3042,N_3224);
or U4480 (N_4480,N_3740,N_3069);
and U4481 (N_4481,N_3990,N_3798);
and U4482 (N_4482,N_3983,N_3261);
nor U4483 (N_4483,N_3485,N_3373);
nand U4484 (N_4484,N_3061,N_3019);
and U4485 (N_4485,N_3786,N_3696);
nand U4486 (N_4486,N_3904,N_3850);
or U4487 (N_4487,N_3231,N_3374);
or U4488 (N_4488,N_3977,N_3905);
nand U4489 (N_4489,N_3348,N_3298);
or U4490 (N_4490,N_3765,N_3920);
nor U4491 (N_4491,N_3622,N_3404);
nand U4492 (N_4492,N_3426,N_3463);
or U4493 (N_4493,N_3831,N_3395);
or U4494 (N_4494,N_3513,N_3945);
and U4495 (N_4495,N_3876,N_3665);
nand U4496 (N_4496,N_3965,N_3912);
and U4497 (N_4497,N_3319,N_3070);
nor U4498 (N_4498,N_3137,N_3382);
or U4499 (N_4499,N_3935,N_3174);
nand U4500 (N_4500,N_3409,N_3905);
nor U4501 (N_4501,N_3739,N_3106);
or U4502 (N_4502,N_3526,N_3380);
nand U4503 (N_4503,N_3550,N_3849);
and U4504 (N_4504,N_3078,N_3930);
or U4505 (N_4505,N_3180,N_3727);
or U4506 (N_4506,N_3437,N_3074);
nand U4507 (N_4507,N_3337,N_3132);
and U4508 (N_4508,N_3819,N_3574);
or U4509 (N_4509,N_3285,N_3830);
or U4510 (N_4510,N_3644,N_3043);
or U4511 (N_4511,N_3775,N_3593);
nand U4512 (N_4512,N_3376,N_3080);
nor U4513 (N_4513,N_3943,N_3035);
nor U4514 (N_4514,N_3922,N_3194);
nor U4515 (N_4515,N_3486,N_3228);
or U4516 (N_4516,N_3521,N_3447);
nand U4517 (N_4517,N_3897,N_3723);
nand U4518 (N_4518,N_3063,N_3206);
or U4519 (N_4519,N_3328,N_3908);
nand U4520 (N_4520,N_3988,N_3899);
nor U4521 (N_4521,N_3950,N_3500);
nor U4522 (N_4522,N_3981,N_3731);
nand U4523 (N_4523,N_3467,N_3558);
and U4524 (N_4524,N_3903,N_3054);
or U4525 (N_4525,N_3160,N_3088);
nor U4526 (N_4526,N_3117,N_3333);
and U4527 (N_4527,N_3498,N_3984);
or U4528 (N_4528,N_3820,N_3589);
and U4529 (N_4529,N_3988,N_3167);
nand U4530 (N_4530,N_3375,N_3891);
or U4531 (N_4531,N_3199,N_3765);
nand U4532 (N_4532,N_3657,N_3447);
and U4533 (N_4533,N_3612,N_3450);
nand U4534 (N_4534,N_3893,N_3879);
or U4535 (N_4535,N_3274,N_3219);
and U4536 (N_4536,N_3598,N_3560);
nand U4537 (N_4537,N_3846,N_3737);
nor U4538 (N_4538,N_3861,N_3276);
nand U4539 (N_4539,N_3749,N_3502);
or U4540 (N_4540,N_3471,N_3820);
nand U4541 (N_4541,N_3127,N_3617);
or U4542 (N_4542,N_3942,N_3443);
or U4543 (N_4543,N_3552,N_3534);
nand U4544 (N_4544,N_3604,N_3338);
nor U4545 (N_4545,N_3316,N_3098);
nand U4546 (N_4546,N_3902,N_3657);
or U4547 (N_4547,N_3050,N_3227);
nand U4548 (N_4548,N_3530,N_3834);
or U4549 (N_4549,N_3485,N_3095);
and U4550 (N_4550,N_3159,N_3197);
or U4551 (N_4551,N_3247,N_3873);
nor U4552 (N_4552,N_3578,N_3675);
or U4553 (N_4553,N_3840,N_3410);
nor U4554 (N_4554,N_3256,N_3397);
nand U4555 (N_4555,N_3286,N_3047);
and U4556 (N_4556,N_3243,N_3493);
nor U4557 (N_4557,N_3830,N_3359);
or U4558 (N_4558,N_3643,N_3055);
nand U4559 (N_4559,N_3361,N_3849);
nand U4560 (N_4560,N_3886,N_3708);
or U4561 (N_4561,N_3993,N_3870);
and U4562 (N_4562,N_3323,N_3865);
nand U4563 (N_4563,N_3497,N_3972);
nand U4564 (N_4564,N_3373,N_3053);
nand U4565 (N_4565,N_3956,N_3718);
nand U4566 (N_4566,N_3446,N_3082);
nor U4567 (N_4567,N_3267,N_3211);
nand U4568 (N_4568,N_3839,N_3238);
or U4569 (N_4569,N_3356,N_3388);
nand U4570 (N_4570,N_3085,N_3791);
or U4571 (N_4571,N_3949,N_3244);
or U4572 (N_4572,N_3712,N_3937);
nor U4573 (N_4573,N_3550,N_3202);
and U4574 (N_4574,N_3977,N_3801);
nand U4575 (N_4575,N_3180,N_3579);
nand U4576 (N_4576,N_3224,N_3048);
nor U4577 (N_4577,N_3529,N_3221);
and U4578 (N_4578,N_3977,N_3601);
nand U4579 (N_4579,N_3468,N_3675);
and U4580 (N_4580,N_3902,N_3016);
nand U4581 (N_4581,N_3556,N_3069);
nor U4582 (N_4582,N_3978,N_3421);
nor U4583 (N_4583,N_3347,N_3408);
or U4584 (N_4584,N_3813,N_3598);
or U4585 (N_4585,N_3669,N_3682);
or U4586 (N_4586,N_3378,N_3164);
or U4587 (N_4587,N_3810,N_3795);
nor U4588 (N_4588,N_3453,N_3410);
nor U4589 (N_4589,N_3217,N_3437);
nor U4590 (N_4590,N_3824,N_3309);
nand U4591 (N_4591,N_3010,N_3856);
nand U4592 (N_4592,N_3079,N_3580);
and U4593 (N_4593,N_3903,N_3567);
and U4594 (N_4594,N_3735,N_3968);
and U4595 (N_4595,N_3119,N_3458);
nor U4596 (N_4596,N_3954,N_3619);
or U4597 (N_4597,N_3280,N_3342);
nand U4598 (N_4598,N_3174,N_3840);
nand U4599 (N_4599,N_3804,N_3991);
nor U4600 (N_4600,N_3982,N_3424);
nand U4601 (N_4601,N_3335,N_3334);
or U4602 (N_4602,N_3265,N_3637);
or U4603 (N_4603,N_3830,N_3846);
nand U4604 (N_4604,N_3789,N_3611);
or U4605 (N_4605,N_3381,N_3029);
and U4606 (N_4606,N_3308,N_3081);
nor U4607 (N_4607,N_3657,N_3676);
nand U4608 (N_4608,N_3549,N_3287);
nor U4609 (N_4609,N_3515,N_3685);
and U4610 (N_4610,N_3340,N_3707);
and U4611 (N_4611,N_3305,N_3568);
nand U4612 (N_4612,N_3982,N_3097);
nor U4613 (N_4613,N_3045,N_3998);
nor U4614 (N_4614,N_3904,N_3586);
nor U4615 (N_4615,N_3614,N_3962);
nor U4616 (N_4616,N_3256,N_3992);
and U4617 (N_4617,N_3989,N_3537);
and U4618 (N_4618,N_3612,N_3054);
or U4619 (N_4619,N_3598,N_3908);
nand U4620 (N_4620,N_3168,N_3573);
nand U4621 (N_4621,N_3752,N_3257);
nand U4622 (N_4622,N_3576,N_3561);
or U4623 (N_4623,N_3195,N_3957);
and U4624 (N_4624,N_3058,N_3976);
nand U4625 (N_4625,N_3524,N_3284);
nor U4626 (N_4626,N_3091,N_3018);
nand U4627 (N_4627,N_3692,N_3943);
nor U4628 (N_4628,N_3819,N_3250);
and U4629 (N_4629,N_3738,N_3715);
nor U4630 (N_4630,N_3357,N_3032);
and U4631 (N_4631,N_3789,N_3587);
and U4632 (N_4632,N_3390,N_3408);
and U4633 (N_4633,N_3828,N_3499);
nand U4634 (N_4634,N_3584,N_3730);
nand U4635 (N_4635,N_3760,N_3621);
or U4636 (N_4636,N_3002,N_3104);
or U4637 (N_4637,N_3217,N_3060);
nand U4638 (N_4638,N_3811,N_3816);
or U4639 (N_4639,N_3694,N_3101);
or U4640 (N_4640,N_3122,N_3148);
nand U4641 (N_4641,N_3080,N_3125);
nand U4642 (N_4642,N_3595,N_3493);
nand U4643 (N_4643,N_3725,N_3679);
or U4644 (N_4644,N_3697,N_3228);
nor U4645 (N_4645,N_3193,N_3349);
and U4646 (N_4646,N_3059,N_3474);
nand U4647 (N_4647,N_3039,N_3022);
and U4648 (N_4648,N_3108,N_3450);
or U4649 (N_4649,N_3067,N_3000);
nor U4650 (N_4650,N_3720,N_3185);
and U4651 (N_4651,N_3782,N_3032);
nand U4652 (N_4652,N_3404,N_3653);
and U4653 (N_4653,N_3501,N_3827);
nor U4654 (N_4654,N_3200,N_3530);
nor U4655 (N_4655,N_3867,N_3522);
and U4656 (N_4656,N_3520,N_3779);
nor U4657 (N_4657,N_3812,N_3254);
nor U4658 (N_4658,N_3724,N_3871);
and U4659 (N_4659,N_3439,N_3505);
nor U4660 (N_4660,N_3288,N_3158);
or U4661 (N_4661,N_3910,N_3664);
nand U4662 (N_4662,N_3043,N_3480);
nand U4663 (N_4663,N_3571,N_3150);
and U4664 (N_4664,N_3757,N_3993);
nand U4665 (N_4665,N_3548,N_3030);
nor U4666 (N_4666,N_3329,N_3815);
nand U4667 (N_4667,N_3674,N_3371);
nor U4668 (N_4668,N_3326,N_3134);
nand U4669 (N_4669,N_3222,N_3115);
or U4670 (N_4670,N_3467,N_3644);
and U4671 (N_4671,N_3796,N_3534);
and U4672 (N_4672,N_3334,N_3574);
and U4673 (N_4673,N_3169,N_3081);
nor U4674 (N_4674,N_3161,N_3552);
and U4675 (N_4675,N_3525,N_3095);
or U4676 (N_4676,N_3207,N_3775);
and U4677 (N_4677,N_3389,N_3274);
and U4678 (N_4678,N_3691,N_3233);
nand U4679 (N_4679,N_3158,N_3163);
or U4680 (N_4680,N_3416,N_3617);
and U4681 (N_4681,N_3062,N_3499);
and U4682 (N_4682,N_3241,N_3166);
and U4683 (N_4683,N_3793,N_3265);
nor U4684 (N_4684,N_3220,N_3706);
xnor U4685 (N_4685,N_3296,N_3508);
nand U4686 (N_4686,N_3671,N_3023);
and U4687 (N_4687,N_3084,N_3966);
nand U4688 (N_4688,N_3792,N_3883);
and U4689 (N_4689,N_3135,N_3851);
or U4690 (N_4690,N_3969,N_3026);
nand U4691 (N_4691,N_3254,N_3296);
or U4692 (N_4692,N_3699,N_3472);
nor U4693 (N_4693,N_3427,N_3975);
nor U4694 (N_4694,N_3392,N_3626);
or U4695 (N_4695,N_3309,N_3838);
nand U4696 (N_4696,N_3243,N_3518);
nand U4697 (N_4697,N_3242,N_3968);
and U4698 (N_4698,N_3562,N_3617);
nand U4699 (N_4699,N_3813,N_3748);
nand U4700 (N_4700,N_3963,N_3334);
or U4701 (N_4701,N_3299,N_3077);
nand U4702 (N_4702,N_3361,N_3489);
nand U4703 (N_4703,N_3558,N_3395);
and U4704 (N_4704,N_3608,N_3753);
nand U4705 (N_4705,N_3093,N_3147);
nor U4706 (N_4706,N_3452,N_3816);
and U4707 (N_4707,N_3917,N_3958);
and U4708 (N_4708,N_3906,N_3851);
nor U4709 (N_4709,N_3685,N_3174);
nor U4710 (N_4710,N_3998,N_3272);
and U4711 (N_4711,N_3199,N_3637);
or U4712 (N_4712,N_3311,N_3287);
or U4713 (N_4713,N_3258,N_3915);
or U4714 (N_4714,N_3973,N_3998);
and U4715 (N_4715,N_3447,N_3956);
nor U4716 (N_4716,N_3551,N_3336);
nor U4717 (N_4717,N_3459,N_3945);
or U4718 (N_4718,N_3391,N_3640);
nor U4719 (N_4719,N_3924,N_3622);
nand U4720 (N_4720,N_3551,N_3371);
nand U4721 (N_4721,N_3286,N_3193);
and U4722 (N_4722,N_3435,N_3495);
nand U4723 (N_4723,N_3762,N_3863);
nand U4724 (N_4724,N_3126,N_3218);
nand U4725 (N_4725,N_3355,N_3772);
and U4726 (N_4726,N_3193,N_3614);
or U4727 (N_4727,N_3749,N_3546);
and U4728 (N_4728,N_3078,N_3530);
or U4729 (N_4729,N_3228,N_3261);
nand U4730 (N_4730,N_3192,N_3636);
nor U4731 (N_4731,N_3984,N_3627);
nor U4732 (N_4732,N_3832,N_3615);
and U4733 (N_4733,N_3255,N_3980);
and U4734 (N_4734,N_3136,N_3326);
nor U4735 (N_4735,N_3162,N_3554);
nor U4736 (N_4736,N_3857,N_3847);
or U4737 (N_4737,N_3803,N_3714);
and U4738 (N_4738,N_3344,N_3090);
or U4739 (N_4739,N_3015,N_3580);
xnor U4740 (N_4740,N_3812,N_3207);
or U4741 (N_4741,N_3896,N_3678);
nor U4742 (N_4742,N_3246,N_3960);
or U4743 (N_4743,N_3341,N_3666);
or U4744 (N_4744,N_3890,N_3541);
nand U4745 (N_4745,N_3963,N_3673);
or U4746 (N_4746,N_3793,N_3412);
and U4747 (N_4747,N_3426,N_3334);
and U4748 (N_4748,N_3788,N_3259);
nand U4749 (N_4749,N_3752,N_3030);
nor U4750 (N_4750,N_3931,N_3179);
or U4751 (N_4751,N_3396,N_3655);
nand U4752 (N_4752,N_3908,N_3930);
or U4753 (N_4753,N_3133,N_3396);
or U4754 (N_4754,N_3561,N_3392);
nor U4755 (N_4755,N_3473,N_3285);
and U4756 (N_4756,N_3211,N_3509);
and U4757 (N_4757,N_3762,N_3264);
nand U4758 (N_4758,N_3327,N_3166);
and U4759 (N_4759,N_3903,N_3371);
or U4760 (N_4760,N_3324,N_3662);
nor U4761 (N_4761,N_3196,N_3579);
or U4762 (N_4762,N_3180,N_3103);
nor U4763 (N_4763,N_3617,N_3182);
or U4764 (N_4764,N_3486,N_3061);
xor U4765 (N_4765,N_3594,N_3489);
and U4766 (N_4766,N_3362,N_3861);
or U4767 (N_4767,N_3196,N_3321);
or U4768 (N_4768,N_3479,N_3030);
nand U4769 (N_4769,N_3009,N_3533);
nand U4770 (N_4770,N_3343,N_3698);
or U4771 (N_4771,N_3525,N_3803);
and U4772 (N_4772,N_3285,N_3578);
or U4773 (N_4773,N_3059,N_3364);
nor U4774 (N_4774,N_3178,N_3523);
and U4775 (N_4775,N_3064,N_3884);
or U4776 (N_4776,N_3219,N_3587);
and U4777 (N_4777,N_3258,N_3224);
nand U4778 (N_4778,N_3104,N_3813);
nand U4779 (N_4779,N_3862,N_3291);
and U4780 (N_4780,N_3580,N_3488);
or U4781 (N_4781,N_3238,N_3552);
nor U4782 (N_4782,N_3611,N_3943);
nand U4783 (N_4783,N_3448,N_3757);
or U4784 (N_4784,N_3460,N_3244);
nand U4785 (N_4785,N_3737,N_3948);
or U4786 (N_4786,N_3186,N_3632);
or U4787 (N_4787,N_3978,N_3014);
or U4788 (N_4788,N_3686,N_3311);
and U4789 (N_4789,N_3176,N_3371);
nand U4790 (N_4790,N_3254,N_3044);
or U4791 (N_4791,N_3541,N_3451);
nor U4792 (N_4792,N_3056,N_3422);
and U4793 (N_4793,N_3408,N_3045);
nor U4794 (N_4794,N_3872,N_3689);
or U4795 (N_4795,N_3871,N_3714);
or U4796 (N_4796,N_3152,N_3581);
and U4797 (N_4797,N_3074,N_3960);
nand U4798 (N_4798,N_3010,N_3165);
nor U4799 (N_4799,N_3645,N_3113);
nand U4800 (N_4800,N_3970,N_3585);
nand U4801 (N_4801,N_3308,N_3475);
nor U4802 (N_4802,N_3209,N_3020);
xnor U4803 (N_4803,N_3353,N_3599);
nand U4804 (N_4804,N_3535,N_3743);
or U4805 (N_4805,N_3698,N_3828);
or U4806 (N_4806,N_3863,N_3085);
and U4807 (N_4807,N_3406,N_3341);
or U4808 (N_4808,N_3330,N_3997);
nor U4809 (N_4809,N_3662,N_3561);
nand U4810 (N_4810,N_3727,N_3796);
and U4811 (N_4811,N_3482,N_3410);
or U4812 (N_4812,N_3223,N_3675);
and U4813 (N_4813,N_3212,N_3668);
nor U4814 (N_4814,N_3867,N_3982);
nor U4815 (N_4815,N_3308,N_3514);
nand U4816 (N_4816,N_3203,N_3555);
nand U4817 (N_4817,N_3018,N_3121);
and U4818 (N_4818,N_3735,N_3966);
nor U4819 (N_4819,N_3585,N_3863);
nor U4820 (N_4820,N_3412,N_3460);
nor U4821 (N_4821,N_3612,N_3055);
nand U4822 (N_4822,N_3035,N_3896);
xor U4823 (N_4823,N_3784,N_3162);
or U4824 (N_4824,N_3301,N_3060);
nand U4825 (N_4825,N_3717,N_3447);
nand U4826 (N_4826,N_3418,N_3816);
nor U4827 (N_4827,N_3465,N_3000);
or U4828 (N_4828,N_3263,N_3910);
nand U4829 (N_4829,N_3363,N_3499);
or U4830 (N_4830,N_3714,N_3740);
and U4831 (N_4831,N_3394,N_3067);
and U4832 (N_4832,N_3453,N_3028);
or U4833 (N_4833,N_3714,N_3193);
and U4834 (N_4834,N_3306,N_3195);
and U4835 (N_4835,N_3165,N_3447);
nand U4836 (N_4836,N_3371,N_3590);
or U4837 (N_4837,N_3829,N_3897);
or U4838 (N_4838,N_3028,N_3586);
and U4839 (N_4839,N_3304,N_3791);
nand U4840 (N_4840,N_3352,N_3558);
nor U4841 (N_4841,N_3514,N_3526);
nand U4842 (N_4842,N_3468,N_3834);
nor U4843 (N_4843,N_3269,N_3645);
nand U4844 (N_4844,N_3173,N_3647);
or U4845 (N_4845,N_3661,N_3482);
or U4846 (N_4846,N_3023,N_3978);
or U4847 (N_4847,N_3707,N_3133);
and U4848 (N_4848,N_3978,N_3440);
or U4849 (N_4849,N_3938,N_3962);
or U4850 (N_4850,N_3404,N_3045);
nor U4851 (N_4851,N_3220,N_3340);
nor U4852 (N_4852,N_3774,N_3781);
nand U4853 (N_4853,N_3567,N_3330);
nand U4854 (N_4854,N_3809,N_3918);
or U4855 (N_4855,N_3681,N_3893);
and U4856 (N_4856,N_3896,N_3747);
and U4857 (N_4857,N_3161,N_3500);
or U4858 (N_4858,N_3506,N_3405);
nor U4859 (N_4859,N_3689,N_3667);
nor U4860 (N_4860,N_3770,N_3381);
nor U4861 (N_4861,N_3663,N_3629);
nor U4862 (N_4862,N_3893,N_3910);
or U4863 (N_4863,N_3006,N_3854);
nand U4864 (N_4864,N_3542,N_3588);
and U4865 (N_4865,N_3169,N_3152);
or U4866 (N_4866,N_3872,N_3864);
xor U4867 (N_4867,N_3610,N_3622);
nand U4868 (N_4868,N_3659,N_3319);
or U4869 (N_4869,N_3615,N_3449);
nand U4870 (N_4870,N_3718,N_3961);
nand U4871 (N_4871,N_3294,N_3142);
nor U4872 (N_4872,N_3653,N_3438);
or U4873 (N_4873,N_3439,N_3110);
and U4874 (N_4874,N_3345,N_3082);
nor U4875 (N_4875,N_3319,N_3376);
nand U4876 (N_4876,N_3045,N_3071);
and U4877 (N_4877,N_3840,N_3994);
nor U4878 (N_4878,N_3130,N_3926);
and U4879 (N_4879,N_3158,N_3017);
and U4880 (N_4880,N_3603,N_3079);
nor U4881 (N_4881,N_3081,N_3661);
nand U4882 (N_4882,N_3556,N_3364);
nand U4883 (N_4883,N_3935,N_3992);
or U4884 (N_4884,N_3325,N_3604);
or U4885 (N_4885,N_3317,N_3272);
nand U4886 (N_4886,N_3725,N_3825);
nor U4887 (N_4887,N_3873,N_3164);
and U4888 (N_4888,N_3710,N_3225);
and U4889 (N_4889,N_3826,N_3108);
and U4890 (N_4890,N_3004,N_3218);
nor U4891 (N_4891,N_3148,N_3282);
or U4892 (N_4892,N_3577,N_3544);
nand U4893 (N_4893,N_3452,N_3214);
and U4894 (N_4894,N_3866,N_3242);
or U4895 (N_4895,N_3943,N_3402);
nand U4896 (N_4896,N_3606,N_3692);
nor U4897 (N_4897,N_3619,N_3383);
or U4898 (N_4898,N_3890,N_3853);
nand U4899 (N_4899,N_3728,N_3950);
and U4900 (N_4900,N_3916,N_3379);
nand U4901 (N_4901,N_3791,N_3545);
nor U4902 (N_4902,N_3702,N_3807);
nor U4903 (N_4903,N_3622,N_3131);
or U4904 (N_4904,N_3555,N_3604);
nand U4905 (N_4905,N_3785,N_3426);
and U4906 (N_4906,N_3273,N_3802);
and U4907 (N_4907,N_3685,N_3565);
xor U4908 (N_4908,N_3107,N_3754);
nor U4909 (N_4909,N_3156,N_3731);
nand U4910 (N_4910,N_3523,N_3011);
nor U4911 (N_4911,N_3638,N_3864);
nand U4912 (N_4912,N_3266,N_3839);
or U4913 (N_4913,N_3165,N_3732);
or U4914 (N_4914,N_3903,N_3770);
and U4915 (N_4915,N_3453,N_3475);
nor U4916 (N_4916,N_3649,N_3511);
nand U4917 (N_4917,N_3090,N_3682);
or U4918 (N_4918,N_3715,N_3634);
and U4919 (N_4919,N_3293,N_3286);
or U4920 (N_4920,N_3772,N_3412);
or U4921 (N_4921,N_3106,N_3753);
nor U4922 (N_4922,N_3852,N_3847);
and U4923 (N_4923,N_3725,N_3973);
nand U4924 (N_4924,N_3121,N_3012);
nand U4925 (N_4925,N_3686,N_3800);
and U4926 (N_4926,N_3675,N_3929);
nor U4927 (N_4927,N_3277,N_3867);
nand U4928 (N_4928,N_3467,N_3576);
nor U4929 (N_4929,N_3800,N_3990);
or U4930 (N_4930,N_3731,N_3363);
and U4931 (N_4931,N_3720,N_3438);
and U4932 (N_4932,N_3824,N_3807);
or U4933 (N_4933,N_3699,N_3164);
or U4934 (N_4934,N_3930,N_3630);
and U4935 (N_4935,N_3402,N_3394);
and U4936 (N_4936,N_3387,N_3447);
and U4937 (N_4937,N_3910,N_3700);
or U4938 (N_4938,N_3249,N_3285);
nand U4939 (N_4939,N_3245,N_3288);
nor U4940 (N_4940,N_3907,N_3515);
xor U4941 (N_4941,N_3668,N_3552);
or U4942 (N_4942,N_3735,N_3639);
nor U4943 (N_4943,N_3250,N_3828);
nor U4944 (N_4944,N_3740,N_3887);
and U4945 (N_4945,N_3501,N_3627);
or U4946 (N_4946,N_3951,N_3535);
or U4947 (N_4947,N_3677,N_3147);
and U4948 (N_4948,N_3177,N_3194);
nor U4949 (N_4949,N_3872,N_3531);
and U4950 (N_4950,N_3553,N_3831);
nand U4951 (N_4951,N_3401,N_3984);
or U4952 (N_4952,N_3636,N_3833);
or U4953 (N_4953,N_3465,N_3531);
and U4954 (N_4954,N_3210,N_3673);
nor U4955 (N_4955,N_3495,N_3182);
nor U4956 (N_4956,N_3155,N_3021);
nor U4957 (N_4957,N_3479,N_3262);
nor U4958 (N_4958,N_3963,N_3718);
and U4959 (N_4959,N_3075,N_3351);
and U4960 (N_4960,N_3203,N_3372);
nor U4961 (N_4961,N_3930,N_3343);
and U4962 (N_4962,N_3592,N_3655);
and U4963 (N_4963,N_3180,N_3487);
nor U4964 (N_4964,N_3249,N_3011);
nor U4965 (N_4965,N_3287,N_3666);
and U4966 (N_4966,N_3201,N_3508);
or U4967 (N_4967,N_3212,N_3752);
nand U4968 (N_4968,N_3809,N_3708);
and U4969 (N_4969,N_3049,N_3207);
and U4970 (N_4970,N_3409,N_3469);
or U4971 (N_4971,N_3130,N_3315);
nor U4972 (N_4972,N_3012,N_3487);
nor U4973 (N_4973,N_3857,N_3453);
nand U4974 (N_4974,N_3552,N_3695);
nor U4975 (N_4975,N_3463,N_3585);
nor U4976 (N_4976,N_3524,N_3476);
or U4977 (N_4977,N_3109,N_3902);
nor U4978 (N_4978,N_3220,N_3338);
nand U4979 (N_4979,N_3810,N_3371);
nor U4980 (N_4980,N_3502,N_3720);
nor U4981 (N_4981,N_3506,N_3299);
or U4982 (N_4982,N_3625,N_3409);
and U4983 (N_4983,N_3586,N_3652);
or U4984 (N_4984,N_3722,N_3994);
nand U4985 (N_4985,N_3442,N_3243);
nand U4986 (N_4986,N_3167,N_3031);
xnor U4987 (N_4987,N_3958,N_3844);
nor U4988 (N_4988,N_3250,N_3043);
and U4989 (N_4989,N_3322,N_3865);
nand U4990 (N_4990,N_3451,N_3806);
or U4991 (N_4991,N_3558,N_3381);
and U4992 (N_4992,N_3378,N_3561);
nor U4993 (N_4993,N_3743,N_3436);
nor U4994 (N_4994,N_3233,N_3553);
nand U4995 (N_4995,N_3251,N_3108);
and U4996 (N_4996,N_3553,N_3600);
nor U4997 (N_4997,N_3775,N_3017);
nand U4998 (N_4998,N_3381,N_3193);
nor U4999 (N_4999,N_3500,N_3125);
nand UO_0 (O_0,N_4076,N_4223);
or UO_1 (O_1,N_4669,N_4581);
or UO_2 (O_2,N_4968,N_4678);
xor UO_3 (O_3,N_4627,N_4804);
and UO_4 (O_4,N_4409,N_4272);
nand UO_5 (O_5,N_4921,N_4514);
nand UO_6 (O_6,N_4543,N_4624);
and UO_7 (O_7,N_4200,N_4722);
xnor UO_8 (O_8,N_4219,N_4760);
nor UO_9 (O_9,N_4558,N_4506);
and UO_10 (O_10,N_4779,N_4807);
and UO_11 (O_11,N_4677,N_4171);
and UO_12 (O_12,N_4960,N_4549);
and UO_13 (O_13,N_4278,N_4276);
and UO_14 (O_14,N_4464,N_4476);
nor UO_15 (O_15,N_4628,N_4946);
or UO_16 (O_16,N_4210,N_4029);
and UO_17 (O_17,N_4745,N_4397);
or UO_18 (O_18,N_4810,N_4562);
or UO_19 (O_19,N_4607,N_4295);
nand UO_20 (O_20,N_4769,N_4172);
nor UO_21 (O_21,N_4164,N_4826);
nand UO_22 (O_22,N_4268,N_4249);
nand UO_23 (O_23,N_4860,N_4613);
nor UO_24 (O_24,N_4286,N_4932);
and UO_25 (O_25,N_4495,N_4440);
nor UO_26 (O_26,N_4143,N_4371);
and UO_27 (O_27,N_4202,N_4472);
nand UO_28 (O_28,N_4261,N_4652);
or UO_29 (O_29,N_4972,N_4827);
or UO_30 (O_30,N_4351,N_4465);
nor UO_31 (O_31,N_4430,N_4701);
nor UO_32 (O_32,N_4438,N_4484);
nor UO_33 (O_33,N_4196,N_4504);
and UO_34 (O_34,N_4439,N_4648);
nand UO_35 (O_35,N_4148,N_4564);
nor UO_36 (O_36,N_4433,N_4363);
or UO_37 (O_37,N_4186,N_4608);
nor UO_38 (O_38,N_4234,N_4141);
or UO_39 (O_39,N_4181,N_4716);
and UO_40 (O_40,N_4471,N_4283);
nand UO_41 (O_41,N_4138,N_4617);
or UO_42 (O_42,N_4067,N_4887);
and UO_43 (O_43,N_4128,N_4855);
and UO_44 (O_44,N_4448,N_4612);
and UO_45 (O_45,N_4051,N_4253);
nand UO_46 (O_46,N_4541,N_4838);
nor UO_47 (O_47,N_4213,N_4707);
nand UO_48 (O_48,N_4193,N_4046);
or UO_49 (O_49,N_4184,N_4797);
or UO_50 (O_50,N_4815,N_4808);
nor UO_51 (O_51,N_4663,N_4052);
and UO_52 (O_52,N_4881,N_4729);
nand UO_53 (O_53,N_4310,N_4749);
nor UO_54 (O_54,N_4830,N_4615);
nand UO_55 (O_55,N_4401,N_4512);
or UO_56 (O_56,N_4711,N_4180);
and UO_57 (O_57,N_4653,N_4486);
nor UO_58 (O_58,N_4545,N_4157);
nand UO_59 (O_59,N_4873,N_4324);
nor UO_60 (O_60,N_4704,N_4890);
nand UO_61 (O_61,N_4415,N_4640);
and UO_62 (O_62,N_4910,N_4466);
or UO_63 (O_63,N_4657,N_4318);
nand UO_64 (O_64,N_4008,N_4799);
nand UO_65 (O_65,N_4584,N_4542);
and UO_66 (O_66,N_4328,N_4867);
or UO_67 (O_67,N_4975,N_4450);
or UO_68 (O_68,N_4053,N_4288);
and UO_69 (O_69,N_4672,N_4435);
or UO_70 (O_70,N_4990,N_4578);
and UO_71 (O_71,N_4422,N_4140);
nor UO_72 (O_72,N_4406,N_4244);
xor UO_73 (O_73,N_4367,N_4939);
and UO_74 (O_74,N_4524,N_4386);
nand UO_75 (O_75,N_4460,N_4854);
nor UO_76 (O_76,N_4851,N_4552);
nor UO_77 (O_77,N_4004,N_4935);
nand UO_78 (O_78,N_4403,N_4313);
nor UO_79 (O_79,N_4370,N_4534);
nand UO_80 (O_80,N_4049,N_4317);
or UO_81 (O_81,N_4275,N_4339);
nand UO_82 (O_82,N_4885,N_4991);
nor UO_83 (O_83,N_4000,N_4812);
or UO_84 (O_84,N_4502,N_4123);
or UO_85 (O_85,N_4727,N_4865);
and UO_86 (O_86,N_4330,N_4600);
nand UO_87 (O_87,N_4267,N_4121);
nor UO_88 (O_88,N_4548,N_4373);
or UO_89 (O_89,N_4378,N_4149);
nor UO_90 (O_90,N_4238,N_4886);
and UO_91 (O_91,N_4287,N_4894);
and UO_92 (O_92,N_4631,N_4299);
nand UO_93 (O_93,N_4952,N_4597);
or UO_94 (O_94,N_4926,N_4764);
and UO_95 (O_95,N_4513,N_4748);
nor UO_96 (O_96,N_4322,N_4679);
nand UO_97 (O_97,N_4957,N_4596);
nand UO_98 (O_98,N_4332,N_4916);
and UO_99 (O_99,N_4658,N_4353);
or UO_100 (O_100,N_4314,N_4845);
nand UO_101 (O_101,N_4226,N_4281);
nor UO_102 (O_102,N_4603,N_4126);
or UO_103 (O_103,N_4013,N_4850);
and UO_104 (O_104,N_4948,N_4966);
or UO_105 (O_105,N_4871,N_4296);
or UO_106 (O_106,N_4849,N_4791);
nand UO_107 (O_107,N_4356,N_4352);
nor UO_108 (O_108,N_4204,N_4737);
and UO_109 (O_109,N_4530,N_4614);
and UO_110 (O_110,N_4835,N_4643);
or UO_111 (O_111,N_4917,N_4576);
nand UO_112 (O_112,N_4374,N_4264);
and UO_113 (O_113,N_4980,N_4458);
nor UO_114 (O_114,N_4290,N_4011);
and UO_115 (O_115,N_4168,N_4396);
nor UO_116 (O_116,N_4787,N_4163);
and UO_117 (O_117,N_4122,N_4247);
nand UO_118 (O_118,N_4577,N_4998);
and UO_119 (O_119,N_4964,N_4803);
nor UO_120 (O_120,N_4602,N_4112);
or UO_121 (O_121,N_4015,N_4417);
and UO_122 (O_122,N_4189,N_4381);
nor UO_123 (O_123,N_4174,N_4003);
or UO_124 (O_124,N_4920,N_4416);
and UO_125 (O_125,N_4041,N_4212);
and UO_126 (O_126,N_4913,N_4647);
nor UO_127 (O_127,N_4266,N_4635);
nand UO_128 (O_128,N_4462,N_4993);
nor UO_129 (O_129,N_4104,N_4637);
nand UO_130 (O_130,N_4989,N_4096);
or UO_131 (O_131,N_4934,N_4077);
or UO_132 (O_132,N_4323,N_4194);
and UO_133 (O_133,N_4329,N_4375);
and UO_134 (O_134,N_4500,N_4733);
and UO_135 (O_135,N_4923,N_4687);
or UO_136 (O_136,N_4992,N_4644);
xor UO_137 (O_137,N_4394,N_4626);
nand UO_138 (O_138,N_4311,N_4694);
nor UO_139 (O_139,N_4840,N_4895);
nor UO_140 (O_140,N_4897,N_4661);
or UO_141 (O_141,N_4135,N_4821);
and UO_142 (O_142,N_4943,N_4216);
nor UO_143 (O_143,N_4379,N_4824);
and UO_144 (O_144,N_4765,N_4587);
nor UO_145 (O_145,N_4071,N_4805);
and UO_146 (O_146,N_4977,N_4982);
or UO_147 (O_147,N_4145,N_4270);
nor UO_148 (O_148,N_4443,N_4304);
nand UO_149 (O_149,N_4959,N_4800);
or UO_150 (O_150,N_4688,N_4254);
or UO_151 (O_151,N_4841,N_4753);
nor UO_152 (O_152,N_4823,N_4674);
nand UO_153 (O_153,N_4882,N_4540);
or UO_154 (O_154,N_4187,N_4069);
and UO_155 (O_155,N_4446,N_4525);
nand UO_156 (O_156,N_4420,N_4491);
and UO_157 (O_157,N_4047,N_4774);
nor UO_158 (O_158,N_4156,N_4349);
nand UO_159 (O_159,N_4207,N_4806);
and UO_160 (O_160,N_4695,N_4079);
and UO_161 (O_161,N_4055,N_4574);
nor UO_162 (O_162,N_4432,N_4445);
nand UO_163 (O_163,N_4241,N_4937);
nor UO_164 (O_164,N_4712,N_4451);
and UO_165 (O_165,N_4933,N_4424);
nand UO_166 (O_166,N_4362,N_4022);
and UO_167 (O_167,N_4852,N_4898);
or UO_168 (O_168,N_4719,N_4246);
nand UO_169 (O_169,N_4338,N_4211);
nor UO_170 (O_170,N_4405,N_4744);
xor UO_171 (O_171,N_4904,N_4586);
or UO_172 (O_172,N_4856,N_4444);
nand UO_173 (O_173,N_4177,N_4896);
or UO_174 (O_174,N_4582,N_4360);
and UO_175 (O_175,N_4080,N_4918);
and UO_176 (O_176,N_4366,N_4428);
or UO_177 (O_177,N_4038,N_4843);
or UO_178 (O_178,N_4588,N_4035);
nand UO_179 (O_179,N_4673,N_4343);
or UO_180 (O_180,N_4068,N_4623);
or UO_181 (O_181,N_4700,N_4818);
and UO_182 (O_182,N_4325,N_4902);
nand UO_183 (O_183,N_4198,N_4456);
nand UO_184 (O_184,N_4876,N_4889);
nand UO_185 (O_185,N_4519,N_4761);
nor UO_186 (O_186,N_4676,N_4585);
or UO_187 (O_187,N_4350,N_4978);
or UO_188 (O_188,N_4814,N_4971);
or UO_189 (O_189,N_4389,N_4593);
or UO_190 (O_190,N_4090,N_4346);
or UO_191 (O_191,N_4880,N_4538);
nor UO_192 (O_192,N_4832,N_4277);
and UO_193 (O_193,N_4134,N_4399);
nor UO_194 (O_194,N_4997,N_4962);
nand UO_195 (O_195,N_4606,N_4162);
nor UO_196 (O_196,N_4085,N_4023);
nand UO_197 (O_197,N_4054,N_4539);
nor UO_198 (O_198,N_4449,N_4706);
and UO_199 (O_199,N_4153,N_4224);
nor UO_200 (O_200,N_4218,N_4611);
nor UO_201 (O_201,N_4119,N_4083);
or UO_202 (O_202,N_4651,N_4878);
and UO_203 (O_203,N_4795,N_4221);
and UO_204 (O_204,N_4645,N_4426);
nand UO_205 (O_205,N_4258,N_4692);
nor UO_206 (O_206,N_4630,N_4892);
and UO_207 (O_207,N_4192,N_4660);
nor UO_208 (O_208,N_4175,N_4293);
or UO_209 (O_209,N_4575,N_4228);
nand UO_210 (O_210,N_4778,N_4215);
and UO_211 (O_211,N_4988,N_4736);
and UO_212 (O_212,N_4928,N_4520);
nand UO_213 (O_213,N_4685,N_4684);
or UO_214 (O_214,N_4714,N_4622);
nand UO_215 (O_215,N_4499,N_4557);
and UO_216 (O_216,N_4709,N_4217);
nand UO_217 (O_217,N_4222,N_4497);
or UO_218 (O_218,N_4167,N_4594);
nand UO_219 (O_219,N_4609,N_4730);
or UO_220 (O_220,N_4127,N_4376);
nand UO_221 (O_221,N_4831,N_4018);
nand UO_222 (O_222,N_4391,N_4559);
and UO_223 (O_223,N_4861,N_4825);
or UO_224 (O_224,N_4869,N_4361);
nor UO_225 (O_225,N_4570,N_4078);
and UO_226 (O_226,N_4477,N_4291);
nand UO_227 (O_227,N_4911,N_4649);
or UO_228 (O_228,N_4527,N_4109);
and UO_229 (O_229,N_4016,N_4750);
nor UO_230 (O_230,N_4133,N_4321);
nand UO_231 (O_231,N_4306,N_4457);
and UO_232 (O_232,N_4037,N_4509);
or UO_233 (O_233,N_4021,N_4205);
nor UO_234 (O_234,N_4877,N_4731);
nand UO_235 (O_235,N_4936,N_4066);
and UO_236 (O_236,N_4307,N_4152);
nand UO_237 (O_237,N_4984,N_4967);
nor UO_238 (O_238,N_4262,N_4014);
or UO_239 (O_239,N_4675,N_4790);
or UO_240 (O_240,N_4395,N_4087);
or UO_241 (O_241,N_4191,N_4697);
or UO_242 (O_242,N_4230,N_4473);
nand UO_243 (O_243,N_4308,N_4252);
nand UO_244 (O_244,N_4400,N_4151);
nand UO_245 (O_245,N_4829,N_4344);
nor UO_246 (O_246,N_4955,N_4620);
nor UO_247 (O_247,N_4418,N_4708);
nor UO_248 (O_248,N_4117,N_4089);
nand UO_249 (O_249,N_4702,N_4682);
nand UO_250 (O_250,N_4377,N_4494);
or UO_251 (O_251,N_4755,N_4522);
nor UO_252 (O_252,N_4533,N_4580);
nor UO_253 (O_253,N_4699,N_4475);
and UO_254 (O_254,N_4336,N_4480);
or UO_255 (O_255,N_4316,N_4488);
nand UO_256 (O_256,N_4309,N_4503);
and UO_257 (O_257,N_4099,N_4847);
nand UO_258 (O_258,N_4767,N_4691);
and UO_259 (O_259,N_4654,N_4033);
nand UO_260 (O_260,N_4801,N_4604);
nand UO_261 (O_261,N_4469,N_4155);
or UO_262 (O_262,N_4265,N_4302);
and UO_263 (O_263,N_4789,N_4728);
or UO_264 (O_264,N_4284,N_4809);
nor UO_265 (O_265,N_4185,N_4392);
or UO_266 (O_266,N_4583,N_4796);
nor UO_267 (O_267,N_4742,N_4837);
nand UO_268 (O_268,N_4772,N_4633);
or UO_269 (O_269,N_4870,N_4380);
nand UO_270 (O_270,N_4160,N_4355);
or UO_271 (O_271,N_4108,N_4632);
or UO_272 (O_272,N_4953,N_4103);
and UO_273 (O_273,N_4250,N_4528);
or UO_274 (O_274,N_4042,N_4616);
nand UO_275 (O_275,N_4650,N_4120);
nor UO_276 (O_276,N_4979,N_4908);
and UO_277 (O_277,N_4853,N_4987);
or UO_278 (O_278,N_4888,N_4834);
and UO_279 (O_279,N_4097,N_4161);
or UO_280 (O_280,N_4048,N_4754);
nor UO_281 (O_281,N_4062,N_4073);
nor UO_282 (O_282,N_4237,N_4358);
nor UO_283 (O_283,N_4065,N_4905);
and UO_284 (O_284,N_4032,N_4693);
nor UO_285 (O_285,N_4176,N_4983);
nand UO_286 (O_286,N_4280,N_4781);
or UO_287 (O_287,N_4173,N_4817);
or UO_288 (O_288,N_4340,N_4973);
or UO_289 (O_289,N_4492,N_4601);
or UO_290 (O_290,N_4482,N_4556);
and UO_291 (O_291,N_4875,N_4555);
nand UO_292 (O_292,N_4759,N_4976);
and UO_293 (O_293,N_4419,N_4107);
and UO_294 (O_294,N_4738,N_4479);
or UO_295 (O_295,N_4348,N_4402);
nor UO_296 (O_296,N_4404,N_4383);
or UO_297 (O_297,N_4822,N_4773);
nand UO_298 (O_298,N_4020,N_4546);
and UO_299 (O_299,N_4740,N_4919);
nand UO_300 (O_300,N_4214,N_4289);
or UO_301 (O_301,N_4188,N_4951);
and UO_302 (O_302,N_4146,N_4040);
nor UO_303 (O_303,N_4461,N_4002);
nand UO_304 (O_304,N_4859,N_4425);
and UO_305 (O_305,N_4592,N_4591);
nor UO_306 (O_306,N_4027,N_4220);
or UO_307 (O_307,N_4547,N_4001);
nor UO_308 (O_308,N_4434,N_4455);
and UO_309 (O_309,N_4178,N_4300);
nand UO_310 (O_310,N_4531,N_4941);
or UO_311 (O_311,N_4681,N_4866);
nand UO_312 (O_312,N_4510,N_4045);
or UO_313 (O_313,N_4165,N_4095);
nor UO_314 (O_314,N_4301,N_4413);
and UO_315 (O_315,N_4638,N_4516);
or UO_316 (O_316,N_4930,N_4408);
and UO_317 (O_317,N_4846,N_4667);
nand UO_318 (O_318,N_4182,N_4137);
or UO_319 (O_319,N_4407,N_4721);
or UO_320 (O_320,N_4084,N_4487);
nand UO_321 (O_321,N_4364,N_4891);
and UO_322 (O_322,N_4026,N_4508);
and UO_323 (O_323,N_4098,N_4092);
and UO_324 (O_324,N_4114,N_4536);
nand UO_325 (O_325,N_4024,N_4965);
nor UO_326 (O_326,N_4326,N_4357);
nor UO_327 (O_327,N_4131,N_4571);
nand UO_328 (O_328,N_4786,N_4414);
nor UO_329 (O_329,N_4197,N_4159);
nand UO_330 (O_330,N_4030,N_4431);
and UO_331 (O_331,N_4726,N_4844);
or UO_332 (O_332,N_4006,N_4044);
nor UO_333 (O_333,N_4816,N_4944);
nand UO_334 (O_334,N_4725,N_4573);
nand UO_335 (O_335,N_4111,N_4642);
nor UO_336 (O_336,N_4320,N_4715);
nand UO_337 (O_337,N_4441,N_4909);
nor UO_338 (O_338,N_4485,N_4423);
or UO_339 (O_339,N_4208,N_4981);
nand UO_340 (O_340,N_4572,N_4739);
nor UO_341 (O_341,N_4437,N_4166);
nand UO_342 (O_342,N_4190,N_4025);
and UO_343 (O_343,N_4005,N_4636);
nand UO_344 (O_344,N_4334,N_4665);
nor UO_345 (O_345,N_4124,N_4158);
nor UO_346 (O_346,N_4752,N_4907);
and UO_347 (O_347,N_4498,N_4511);
and UO_348 (O_348,N_4515,N_4100);
or UO_349 (O_349,N_4368,N_4341);
and UO_350 (O_350,N_4927,N_4255);
nand UO_351 (O_351,N_4427,N_4950);
nand UO_352 (O_352,N_4478,N_4086);
nand UO_353 (O_353,N_4879,N_4369);
nand UO_354 (O_354,N_4839,N_4147);
and UO_355 (O_355,N_4751,N_4345);
and UO_356 (O_356,N_4331,N_4996);
or UO_357 (O_357,N_4811,N_4274);
nand UO_358 (O_358,N_4010,N_4929);
or UO_359 (O_359,N_4703,N_4337);
nor UO_360 (O_360,N_4958,N_4820);
and UO_361 (O_361,N_4819,N_4836);
nand UO_362 (O_362,N_4792,N_4554);
nand UO_363 (O_363,N_4646,N_4668);
nor UO_364 (O_364,N_4619,N_4315);
and UO_365 (O_365,N_4940,N_4985);
nor UO_366 (O_366,N_4259,N_4139);
nor UO_367 (O_367,N_4914,N_4059);
nor UO_368 (O_368,N_4017,N_4771);
and UO_369 (O_369,N_4798,N_4229);
or UO_370 (O_370,N_4150,N_4347);
or UO_371 (O_371,N_4579,N_4903);
nor UO_372 (O_372,N_4741,N_4297);
or UO_373 (O_373,N_4091,N_4747);
nand UO_374 (O_374,N_4842,N_4093);
nor UO_375 (O_375,N_4793,N_4680);
nand UO_376 (O_376,N_4947,N_4075);
and UO_377 (O_377,N_4567,N_4169);
or UO_378 (O_378,N_4813,N_4243);
nand UO_379 (O_379,N_4639,N_4209);
or UO_380 (O_380,N_4470,N_4088);
nor UO_381 (O_381,N_4686,N_4129);
and UO_382 (O_382,N_4061,N_4411);
and UO_383 (O_383,N_4766,N_4938);
nor UO_384 (O_384,N_4945,N_4279);
nand UO_385 (O_385,N_4618,N_4718);
nor UO_386 (O_386,N_4012,N_4670);
and UO_387 (O_387,N_4056,N_4206);
nor UO_388 (O_388,N_4136,N_4312);
and UO_389 (O_389,N_4590,N_4863);
or UO_390 (O_390,N_4292,N_4285);
and UO_391 (O_391,N_4009,N_4452);
nor UO_392 (O_392,N_4862,N_4641);
nand UO_393 (O_393,N_4532,N_4273);
and UO_394 (O_394,N_4231,N_4036);
or UO_395 (O_395,N_4768,N_4294);
or UO_396 (O_396,N_4656,N_4746);
nor UO_397 (O_397,N_4550,N_4857);
nor UO_398 (O_398,N_4864,N_4453);
nand UO_399 (O_399,N_4101,N_4954);
or UO_400 (O_400,N_4529,N_4634);
and UO_401 (O_401,N_4717,N_4305);
nand UO_402 (O_402,N_4743,N_4248);
or UO_403 (O_403,N_4783,N_4442);
or UO_404 (O_404,N_4999,N_4621);
or UO_405 (O_405,N_4082,N_4232);
nand UO_406 (O_406,N_4788,N_4382);
and UO_407 (O_407,N_4689,N_4335);
nor UO_408 (O_408,N_4565,N_4963);
nor UO_409 (O_409,N_4154,N_4970);
nor UO_410 (O_410,N_4666,N_4388);
or UO_411 (O_411,N_4034,N_4398);
nor UO_412 (O_412,N_4116,N_4115);
or UO_413 (O_413,N_4063,N_4393);
nor UO_414 (O_414,N_4605,N_4777);
or UO_415 (O_415,N_4359,N_4130);
nand UO_416 (O_416,N_4705,N_4732);
nand UO_417 (O_417,N_4544,N_4598);
nand UO_418 (O_418,N_4995,N_4447);
xor UO_419 (O_419,N_4251,N_4235);
nor UO_420 (O_420,N_4327,N_4893);
or UO_421 (O_421,N_4459,N_4263);
nand UO_422 (O_422,N_4523,N_4481);
or UO_423 (O_423,N_4986,N_4303);
nor UO_424 (O_424,N_4553,N_4319);
nor UO_425 (O_425,N_4081,N_4956);
and UO_426 (O_426,N_4412,N_4256);
nand UO_427 (O_427,N_4526,N_4901);
nand UO_428 (O_428,N_4170,N_4659);
or UO_429 (O_429,N_4463,N_4961);
and UO_430 (O_430,N_4105,N_4125);
nor UO_431 (O_431,N_4384,N_4118);
and UO_432 (O_432,N_4713,N_4271);
or UO_433 (O_433,N_4354,N_4195);
nand UO_434 (O_434,N_4517,N_4028);
and UO_435 (O_435,N_4489,N_4610);
or UO_436 (O_436,N_4900,N_4833);
and UO_437 (O_437,N_4385,N_4925);
and UO_438 (O_438,N_4429,N_4242);
and UO_439 (O_439,N_4199,N_4734);
or UO_440 (O_440,N_4794,N_4912);
nand UO_441 (O_441,N_4183,N_4269);
nand UO_442 (O_442,N_4922,N_4257);
or UO_443 (O_443,N_4698,N_4974);
nand UO_444 (O_444,N_4072,N_4203);
or UO_445 (O_445,N_4333,N_4372);
and UO_446 (O_446,N_4671,N_4770);
and UO_447 (O_447,N_4282,N_4735);
and UO_448 (O_448,N_4240,N_4179);
and UO_449 (O_449,N_4784,N_4505);
and UO_450 (O_450,N_4690,N_4696);
and UO_451 (O_451,N_4858,N_4227);
nand UO_452 (O_452,N_4490,N_4724);
and UO_453 (O_453,N_4780,N_4915);
and UO_454 (O_454,N_4899,N_4507);
and UO_455 (O_455,N_4994,N_4058);
and UO_456 (O_456,N_4239,N_4233);
nor UO_457 (O_457,N_4102,N_4537);
nor UO_458 (O_458,N_4043,N_4201);
or UO_459 (O_459,N_4501,N_4563);
or UO_460 (O_460,N_4496,N_4756);
nor UO_461 (O_461,N_4094,N_4662);
nor UO_462 (O_462,N_4070,N_4785);
nor UO_463 (O_463,N_4454,N_4521);
or UO_464 (O_464,N_4483,N_4387);
or UO_465 (O_465,N_4763,N_4106);
and UO_466 (O_466,N_4874,N_4949);
nand UO_467 (O_467,N_4758,N_4625);
nor UO_468 (O_468,N_4629,N_4931);
or UO_469 (O_469,N_4560,N_4144);
nor UO_470 (O_470,N_4468,N_4031);
and UO_471 (O_471,N_4599,N_4236);
and UO_472 (O_472,N_4872,N_4868);
nor UO_473 (O_473,N_4225,N_4723);
nor UO_474 (O_474,N_4710,N_4906);
nor UO_475 (O_475,N_4883,N_4260);
nand UO_476 (O_476,N_4518,N_4142);
and UO_477 (O_477,N_4390,N_4884);
and UO_478 (O_478,N_4050,N_4110);
and UO_479 (O_479,N_4245,N_4074);
nand UO_480 (O_480,N_4057,N_4365);
or UO_481 (O_481,N_4782,N_4569);
nand UO_482 (O_482,N_4776,N_4467);
and UO_483 (O_483,N_4132,N_4969);
and UO_484 (O_484,N_4342,N_4064);
nand UO_485 (O_485,N_4493,N_4720);
nor UO_486 (O_486,N_4655,N_4802);
nand UO_487 (O_487,N_4410,N_4019);
nor UO_488 (O_488,N_4561,N_4060);
and UO_489 (O_489,N_4942,N_4775);
and UO_490 (O_490,N_4683,N_4828);
or UO_491 (O_491,N_4007,N_4848);
and UO_492 (O_492,N_4436,N_4589);
nand UO_493 (O_493,N_4762,N_4535);
nand UO_494 (O_494,N_4421,N_4298);
nand UO_495 (O_495,N_4595,N_4039);
nand UO_496 (O_496,N_4113,N_4664);
nand UO_497 (O_497,N_4568,N_4924);
nor UO_498 (O_498,N_4474,N_4566);
nand UO_499 (O_499,N_4757,N_4551);
nor UO_500 (O_500,N_4256,N_4343);
nand UO_501 (O_501,N_4491,N_4501);
or UO_502 (O_502,N_4624,N_4126);
or UO_503 (O_503,N_4449,N_4587);
nor UO_504 (O_504,N_4028,N_4997);
or UO_505 (O_505,N_4231,N_4795);
or UO_506 (O_506,N_4907,N_4505);
nand UO_507 (O_507,N_4698,N_4845);
or UO_508 (O_508,N_4539,N_4357);
and UO_509 (O_509,N_4396,N_4466);
nand UO_510 (O_510,N_4318,N_4601);
or UO_511 (O_511,N_4462,N_4636);
and UO_512 (O_512,N_4362,N_4506);
or UO_513 (O_513,N_4710,N_4121);
nor UO_514 (O_514,N_4590,N_4373);
nand UO_515 (O_515,N_4593,N_4613);
and UO_516 (O_516,N_4526,N_4170);
nor UO_517 (O_517,N_4158,N_4756);
and UO_518 (O_518,N_4345,N_4310);
and UO_519 (O_519,N_4176,N_4509);
nand UO_520 (O_520,N_4327,N_4909);
nor UO_521 (O_521,N_4433,N_4180);
and UO_522 (O_522,N_4765,N_4933);
nor UO_523 (O_523,N_4001,N_4273);
or UO_524 (O_524,N_4044,N_4120);
or UO_525 (O_525,N_4068,N_4598);
and UO_526 (O_526,N_4365,N_4964);
and UO_527 (O_527,N_4755,N_4409);
nor UO_528 (O_528,N_4742,N_4527);
or UO_529 (O_529,N_4784,N_4036);
or UO_530 (O_530,N_4272,N_4579);
and UO_531 (O_531,N_4788,N_4146);
or UO_532 (O_532,N_4313,N_4677);
xor UO_533 (O_533,N_4444,N_4064);
nor UO_534 (O_534,N_4956,N_4948);
nand UO_535 (O_535,N_4236,N_4462);
and UO_536 (O_536,N_4513,N_4699);
nor UO_537 (O_537,N_4377,N_4781);
nor UO_538 (O_538,N_4791,N_4533);
nor UO_539 (O_539,N_4437,N_4600);
or UO_540 (O_540,N_4058,N_4030);
nand UO_541 (O_541,N_4517,N_4381);
or UO_542 (O_542,N_4961,N_4188);
and UO_543 (O_543,N_4794,N_4571);
and UO_544 (O_544,N_4697,N_4552);
and UO_545 (O_545,N_4089,N_4425);
and UO_546 (O_546,N_4478,N_4101);
and UO_547 (O_547,N_4375,N_4386);
nor UO_548 (O_548,N_4845,N_4429);
nor UO_549 (O_549,N_4116,N_4915);
nand UO_550 (O_550,N_4903,N_4864);
nand UO_551 (O_551,N_4008,N_4083);
and UO_552 (O_552,N_4217,N_4059);
nand UO_553 (O_553,N_4603,N_4014);
or UO_554 (O_554,N_4740,N_4168);
nor UO_555 (O_555,N_4071,N_4294);
and UO_556 (O_556,N_4430,N_4345);
nor UO_557 (O_557,N_4979,N_4861);
and UO_558 (O_558,N_4998,N_4674);
nand UO_559 (O_559,N_4573,N_4537);
nand UO_560 (O_560,N_4746,N_4065);
nor UO_561 (O_561,N_4524,N_4314);
or UO_562 (O_562,N_4073,N_4440);
nand UO_563 (O_563,N_4794,N_4460);
and UO_564 (O_564,N_4997,N_4696);
nor UO_565 (O_565,N_4029,N_4098);
nand UO_566 (O_566,N_4818,N_4536);
nand UO_567 (O_567,N_4008,N_4848);
xnor UO_568 (O_568,N_4280,N_4687);
or UO_569 (O_569,N_4753,N_4097);
nor UO_570 (O_570,N_4549,N_4030);
nand UO_571 (O_571,N_4981,N_4649);
nand UO_572 (O_572,N_4643,N_4690);
nor UO_573 (O_573,N_4731,N_4995);
and UO_574 (O_574,N_4515,N_4384);
nand UO_575 (O_575,N_4510,N_4683);
nor UO_576 (O_576,N_4045,N_4080);
nand UO_577 (O_577,N_4591,N_4729);
nor UO_578 (O_578,N_4582,N_4672);
and UO_579 (O_579,N_4517,N_4367);
and UO_580 (O_580,N_4323,N_4984);
and UO_581 (O_581,N_4118,N_4993);
and UO_582 (O_582,N_4193,N_4772);
nand UO_583 (O_583,N_4792,N_4921);
nor UO_584 (O_584,N_4253,N_4152);
nand UO_585 (O_585,N_4104,N_4180);
and UO_586 (O_586,N_4429,N_4604);
or UO_587 (O_587,N_4933,N_4410);
nand UO_588 (O_588,N_4469,N_4435);
and UO_589 (O_589,N_4008,N_4004);
or UO_590 (O_590,N_4407,N_4780);
and UO_591 (O_591,N_4019,N_4699);
nand UO_592 (O_592,N_4672,N_4252);
and UO_593 (O_593,N_4073,N_4314);
nand UO_594 (O_594,N_4900,N_4529);
nand UO_595 (O_595,N_4083,N_4611);
or UO_596 (O_596,N_4833,N_4486);
nor UO_597 (O_597,N_4429,N_4187);
nand UO_598 (O_598,N_4751,N_4186);
nand UO_599 (O_599,N_4283,N_4583);
and UO_600 (O_600,N_4120,N_4228);
and UO_601 (O_601,N_4034,N_4747);
nand UO_602 (O_602,N_4171,N_4596);
nor UO_603 (O_603,N_4320,N_4235);
xnor UO_604 (O_604,N_4365,N_4394);
nor UO_605 (O_605,N_4609,N_4140);
nand UO_606 (O_606,N_4904,N_4738);
nor UO_607 (O_607,N_4432,N_4110);
nand UO_608 (O_608,N_4988,N_4304);
or UO_609 (O_609,N_4174,N_4061);
and UO_610 (O_610,N_4319,N_4528);
or UO_611 (O_611,N_4998,N_4404);
or UO_612 (O_612,N_4412,N_4963);
and UO_613 (O_613,N_4611,N_4219);
or UO_614 (O_614,N_4042,N_4193);
or UO_615 (O_615,N_4291,N_4052);
and UO_616 (O_616,N_4112,N_4888);
nor UO_617 (O_617,N_4638,N_4198);
or UO_618 (O_618,N_4739,N_4685);
nand UO_619 (O_619,N_4720,N_4203);
nor UO_620 (O_620,N_4443,N_4953);
or UO_621 (O_621,N_4058,N_4544);
nand UO_622 (O_622,N_4205,N_4563);
and UO_623 (O_623,N_4232,N_4551);
and UO_624 (O_624,N_4654,N_4685);
or UO_625 (O_625,N_4229,N_4479);
nor UO_626 (O_626,N_4749,N_4152);
and UO_627 (O_627,N_4407,N_4649);
nor UO_628 (O_628,N_4904,N_4287);
nor UO_629 (O_629,N_4054,N_4532);
nand UO_630 (O_630,N_4997,N_4908);
nand UO_631 (O_631,N_4956,N_4750);
nor UO_632 (O_632,N_4209,N_4337);
or UO_633 (O_633,N_4508,N_4539);
nor UO_634 (O_634,N_4630,N_4290);
and UO_635 (O_635,N_4427,N_4548);
nand UO_636 (O_636,N_4195,N_4091);
or UO_637 (O_637,N_4914,N_4600);
and UO_638 (O_638,N_4141,N_4653);
and UO_639 (O_639,N_4892,N_4419);
nand UO_640 (O_640,N_4497,N_4411);
nor UO_641 (O_641,N_4953,N_4852);
nor UO_642 (O_642,N_4192,N_4066);
nand UO_643 (O_643,N_4490,N_4546);
nand UO_644 (O_644,N_4039,N_4607);
and UO_645 (O_645,N_4901,N_4562);
or UO_646 (O_646,N_4146,N_4310);
nand UO_647 (O_647,N_4215,N_4551);
or UO_648 (O_648,N_4179,N_4678);
nor UO_649 (O_649,N_4616,N_4893);
nand UO_650 (O_650,N_4883,N_4769);
nand UO_651 (O_651,N_4366,N_4276);
nand UO_652 (O_652,N_4272,N_4890);
nor UO_653 (O_653,N_4242,N_4186);
or UO_654 (O_654,N_4571,N_4947);
or UO_655 (O_655,N_4090,N_4559);
xor UO_656 (O_656,N_4559,N_4265);
and UO_657 (O_657,N_4498,N_4217);
nand UO_658 (O_658,N_4862,N_4328);
or UO_659 (O_659,N_4825,N_4829);
nand UO_660 (O_660,N_4380,N_4367);
and UO_661 (O_661,N_4212,N_4748);
nor UO_662 (O_662,N_4117,N_4348);
or UO_663 (O_663,N_4170,N_4017);
or UO_664 (O_664,N_4907,N_4739);
nand UO_665 (O_665,N_4998,N_4325);
nor UO_666 (O_666,N_4567,N_4672);
or UO_667 (O_667,N_4861,N_4410);
and UO_668 (O_668,N_4934,N_4734);
or UO_669 (O_669,N_4585,N_4117);
or UO_670 (O_670,N_4257,N_4177);
nor UO_671 (O_671,N_4119,N_4821);
nand UO_672 (O_672,N_4533,N_4030);
and UO_673 (O_673,N_4705,N_4806);
and UO_674 (O_674,N_4222,N_4527);
or UO_675 (O_675,N_4737,N_4376);
nor UO_676 (O_676,N_4682,N_4373);
or UO_677 (O_677,N_4328,N_4700);
nor UO_678 (O_678,N_4742,N_4031);
nand UO_679 (O_679,N_4786,N_4658);
nor UO_680 (O_680,N_4745,N_4775);
and UO_681 (O_681,N_4641,N_4923);
or UO_682 (O_682,N_4112,N_4987);
and UO_683 (O_683,N_4482,N_4959);
and UO_684 (O_684,N_4846,N_4971);
and UO_685 (O_685,N_4081,N_4974);
nor UO_686 (O_686,N_4553,N_4969);
and UO_687 (O_687,N_4278,N_4494);
nor UO_688 (O_688,N_4205,N_4192);
nand UO_689 (O_689,N_4091,N_4207);
nand UO_690 (O_690,N_4707,N_4946);
and UO_691 (O_691,N_4957,N_4103);
nor UO_692 (O_692,N_4026,N_4334);
and UO_693 (O_693,N_4474,N_4854);
nor UO_694 (O_694,N_4470,N_4370);
and UO_695 (O_695,N_4570,N_4555);
and UO_696 (O_696,N_4868,N_4828);
or UO_697 (O_697,N_4757,N_4903);
and UO_698 (O_698,N_4993,N_4177);
and UO_699 (O_699,N_4958,N_4848);
nand UO_700 (O_700,N_4197,N_4053);
nor UO_701 (O_701,N_4864,N_4974);
and UO_702 (O_702,N_4598,N_4539);
nor UO_703 (O_703,N_4699,N_4559);
or UO_704 (O_704,N_4024,N_4413);
nand UO_705 (O_705,N_4924,N_4798);
and UO_706 (O_706,N_4309,N_4828);
and UO_707 (O_707,N_4709,N_4408);
nand UO_708 (O_708,N_4583,N_4794);
nand UO_709 (O_709,N_4268,N_4402);
or UO_710 (O_710,N_4823,N_4582);
nor UO_711 (O_711,N_4680,N_4569);
nor UO_712 (O_712,N_4610,N_4513);
nand UO_713 (O_713,N_4875,N_4181);
nand UO_714 (O_714,N_4475,N_4562);
xnor UO_715 (O_715,N_4562,N_4975);
or UO_716 (O_716,N_4837,N_4503);
or UO_717 (O_717,N_4428,N_4509);
and UO_718 (O_718,N_4890,N_4099);
nor UO_719 (O_719,N_4795,N_4326);
nor UO_720 (O_720,N_4988,N_4845);
nand UO_721 (O_721,N_4980,N_4626);
or UO_722 (O_722,N_4105,N_4729);
nand UO_723 (O_723,N_4236,N_4523);
or UO_724 (O_724,N_4960,N_4483);
or UO_725 (O_725,N_4343,N_4790);
nor UO_726 (O_726,N_4506,N_4325);
and UO_727 (O_727,N_4453,N_4523);
nor UO_728 (O_728,N_4925,N_4168);
nor UO_729 (O_729,N_4608,N_4305);
or UO_730 (O_730,N_4409,N_4797);
and UO_731 (O_731,N_4815,N_4844);
nand UO_732 (O_732,N_4160,N_4207);
nand UO_733 (O_733,N_4482,N_4971);
or UO_734 (O_734,N_4889,N_4844);
and UO_735 (O_735,N_4943,N_4860);
nand UO_736 (O_736,N_4298,N_4497);
and UO_737 (O_737,N_4439,N_4462);
or UO_738 (O_738,N_4492,N_4378);
nor UO_739 (O_739,N_4680,N_4399);
and UO_740 (O_740,N_4049,N_4693);
and UO_741 (O_741,N_4764,N_4852);
or UO_742 (O_742,N_4337,N_4725);
and UO_743 (O_743,N_4454,N_4869);
nor UO_744 (O_744,N_4353,N_4783);
or UO_745 (O_745,N_4090,N_4772);
nand UO_746 (O_746,N_4766,N_4393);
nor UO_747 (O_747,N_4316,N_4361);
nand UO_748 (O_748,N_4127,N_4969);
nor UO_749 (O_749,N_4847,N_4999);
or UO_750 (O_750,N_4679,N_4638);
and UO_751 (O_751,N_4594,N_4656);
or UO_752 (O_752,N_4088,N_4016);
nor UO_753 (O_753,N_4053,N_4139);
and UO_754 (O_754,N_4107,N_4670);
and UO_755 (O_755,N_4567,N_4693);
and UO_756 (O_756,N_4476,N_4789);
or UO_757 (O_757,N_4836,N_4911);
nor UO_758 (O_758,N_4010,N_4738);
nor UO_759 (O_759,N_4184,N_4229);
nor UO_760 (O_760,N_4594,N_4522);
and UO_761 (O_761,N_4427,N_4573);
and UO_762 (O_762,N_4398,N_4321);
nor UO_763 (O_763,N_4102,N_4131);
or UO_764 (O_764,N_4956,N_4930);
nor UO_765 (O_765,N_4216,N_4289);
nor UO_766 (O_766,N_4360,N_4288);
nor UO_767 (O_767,N_4571,N_4416);
nand UO_768 (O_768,N_4480,N_4792);
and UO_769 (O_769,N_4784,N_4597);
and UO_770 (O_770,N_4693,N_4604);
and UO_771 (O_771,N_4239,N_4612);
nor UO_772 (O_772,N_4638,N_4587);
nand UO_773 (O_773,N_4740,N_4416);
or UO_774 (O_774,N_4510,N_4443);
nor UO_775 (O_775,N_4575,N_4541);
or UO_776 (O_776,N_4977,N_4022);
or UO_777 (O_777,N_4000,N_4150);
and UO_778 (O_778,N_4940,N_4765);
or UO_779 (O_779,N_4548,N_4115);
and UO_780 (O_780,N_4346,N_4625);
nand UO_781 (O_781,N_4452,N_4086);
or UO_782 (O_782,N_4684,N_4079);
nor UO_783 (O_783,N_4269,N_4213);
nand UO_784 (O_784,N_4199,N_4024);
and UO_785 (O_785,N_4932,N_4847);
nand UO_786 (O_786,N_4516,N_4483);
or UO_787 (O_787,N_4977,N_4035);
or UO_788 (O_788,N_4271,N_4345);
or UO_789 (O_789,N_4967,N_4328);
nand UO_790 (O_790,N_4959,N_4326);
nor UO_791 (O_791,N_4357,N_4237);
and UO_792 (O_792,N_4053,N_4104);
or UO_793 (O_793,N_4908,N_4865);
nand UO_794 (O_794,N_4232,N_4660);
nor UO_795 (O_795,N_4611,N_4979);
or UO_796 (O_796,N_4283,N_4384);
nand UO_797 (O_797,N_4101,N_4220);
nand UO_798 (O_798,N_4052,N_4474);
nor UO_799 (O_799,N_4431,N_4731);
nor UO_800 (O_800,N_4583,N_4569);
or UO_801 (O_801,N_4587,N_4141);
nor UO_802 (O_802,N_4062,N_4972);
nor UO_803 (O_803,N_4750,N_4004);
and UO_804 (O_804,N_4621,N_4670);
nor UO_805 (O_805,N_4578,N_4684);
or UO_806 (O_806,N_4020,N_4966);
and UO_807 (O_807,N_4192,N_4639);
nand UO_808 (O_808,N_4851,N_4793);
or UO_809 (O_809,N_4771,N_4108);
nor UO_810 (O_810,N_4654,N_4393);
nor UO_811 (O_811,N_4060,N_4379);
nor UO_812 (O_812,N_4844,N_4303);
or UO_813 (O_813,N_4623,N_4230);
nand UO_814 (O_814,N_4600,N_4615);
nor UO_815 (O_815,N_4121,N_4357);
nor UO_816 (O_816,N_4066,N_4404);
nand UO_817 (O_817,N_4706,N_4624);
and UO_818 (O_818,N_4330,N_4823);
nor UO_819 (O_819,N_4027,N_4406);
nand UO_820 (O_820,N_4413,N_4005);
or UO_821 (O_821,N_4397,N_4466);
or UO_822 (O_822,N_4483,N_4344);
or UO_823 (O_823,N_4272,N_4371);
or UO_824 (O_824,N_4865,N_4028);
nor UO_825 (O_825,N_4468,N_4866);
or UO_826 (O_826,N_4488,N_4799);
nand UO_827 (O_827,N_4869,N_4574);
or UO_828 (O_828,N_4557,N_4295);
nand UO_829 (O_829,N_4307,N_4115);
or UO_830 (O_830,N_4656,N_4123);
and UO_831 (O_831,N_4361,N_4757);
nor UO_832 (O_832,N_4609,N_4680);
or UO_833 (O_833,N_4783,N_4261);
nor UO_834 (O_834,N_4292,N_4834);
nor UO_835 (O_835,N_4668,N_4420);
or UO_836 (O_836,N_4466,N_4394);
or UO_837 (O_837,N_4196,N_4652);
and UO_838 (O_838,N_4410,N_4151);
or UO_839 (O_839,N_4930,N_4821);
nand UO_840 (O_840,N_4695,N_4296);
or UO_841 (O_841,N_4051,N_4284);
nand UO_842 (O_842,N_4216,N_4824);
nand UO_843 (O_843,N_4054,N_4808);
nand UO_844 (O_844,N_4488,N_4117);
or UO_845 (O_845,N_4337,N_4903);
or UO_846 (O_846,N_4962,N_4661);
nor UO_847 (O_847,N_4871,N_4758);
or UO_848 (O_848,N_4389,N_4647);
or UO_849 (O_849,N_4913,N_4749);
nand UO_850 (O_850,N_4093,N_4109);
nor UO_851 (O_851,N_4345,N_4116);
nand UO_852 (O_852,N_4661,N_4078);
nor UO_853 (O_853,N_4786,N_4582);
nand UO_854 (O_854,N_4429,N_4856);
nand UO_855 (O_855,N_4001,N_4964);
nor UO_856 (O_856,N_4482,N_4503);
and UO_857 (O_857,N_4272,N_4639);
nor UO_858 (O_858,N_4868,N_4846);
nand UO_859 (O_859,N_4704,N_4010);
and UO_860 (O_860,N_4463,N_4060);
or UO_861 (O_861,N_4545,N_4538);
or UO_862 (O_862,N_4485,N_4031);
or UO_863 (O_863,N_4477,N_4115);
nand UO_864 (O_864,N_4763,N_4385);
nor UO_865 (O_865,N_4440,N_4382);
or UO_866 (O_866,N_4990,N_4472);
nor UO_867 (O_867,N_4873,N_4298);
nor UO_868 (O_868,N_4657,N_4999);
or UO_869 (O_869,N_4475,N_4871);
and UO_870 (O_870,N_4901,N_4884);
nand UO_871 (O_871,N_4126,N_4295);
or UO_872 (O_872,N_4033,N_4695);
and UO_873 (O_873,N_4886,N_4254);
nand UO_874 (O_874,N_4287,N_4510);
and UO_875 (O_875,N_4764,N_4565);
and UO_876 (O_876,N_4409,N_4150);
or UO_877 (O_877,N_4119,N_4774);
xnor UO_878 (O_878,N_4862,N_4080);
and UO_879 (O_879,N_4045,N_4481);
and UO_880 (O_880,N_4372,N_4430);
nor UO_881 (O_881,N_4064,N_4496);
nor UO_882 (O_882,N_4589,N_4957);
nand UO_883 (O_883,N_4901,N_4763);
nor UO_884 (O_884,N_4053,N_4767);
and UO_885 (O_885,N_4365,N_4536);
or UO_886 (O_886,N_4842,N_4997);
xnor UO_887 (O_887,N_4974,N_4845);
and UO_888 (O_888,N_4291,N_4596);
nand UO_889 (O_889,N_4755,N_4758);
nand UO_890 (O_890,N_4524,N_4354);
or UO_891 (O_891,N_4755,N_4044);
nor UO_892 (O_892,N_4152,N_4746);
or UO_893 (O_893,N_4649,N_4120);
or UO_894 (O_894,N_4683,N_4498);
nand UO_895 (O_895,N_4921,N_4043);
nand UO_896 (O_896,N_4790,N_4811);
or UO_897 (O_897,N_4138,N_4395);
or UO_898 (O_898,N_4876,N_4423);
and UO_899 (O_899,N_4317,N_4988);
and UO_900 (O_900,N_4444,N_4504);
and UO_901 (O_901,N_4349,N_4993);
nor UO_902 (O_902,N_4436,N_4324);
nor UO_903 (O_903,N_4035,N_4992);
and UO_904 (O_904,N_4082,N_4263);
nor UO_905 (O_905,N_4861,N_4776);
or UO_906 (O_906,N_4567,N_4202);
and UO_907 (O_907,N_4676,N_4911);
nand UO_908 (O_908,N_4264,N_4622);
and UO_909 (O_909,N_4469,N_4105);
nand UO_910 (O_910,N_4362,N_4956);
or UO_911 (O_911,N_4296,N_4039);
or UO_912 (O_912,N_4341,N_4906);
or UO_913 (O_913,N_4865,N_4645);
nor UO_914 (O_914,N_4215,N_4402);
nor UO_915 (O_915,N_4374,N_4130);
nor UO_916 (O_916,N_4284,N_4028);
nand UO_917 (O_917,N_4714,N_4320);
nand UO_918 (O_918,N_4737,N_4256);
nor UO_919 (O_919,N_4712,N_4697);
nand UO_920 (O_920,N_4373,N_4435);
nand UO_921 (O_921,N_4443,N_4027);
and UO_922 (O_922,N_4755,N_4662);
nand UO_923 (O_923,N_4789,N_4184);
nor UO_924 (O_924,N_4141,N_4863);
nor UO_925 (O_925,N_4524,N_4379);
nand UO_926 (O_926,N_4522,N_4002);
or UO_927 (O_927,N_4452,N_4673);
nor UO_928 (O_928,N_4358,N_4636);
or UO_929 (O_929,N_4950,N_4319);
or UO_930 (O_930,N_4092,N_4854);
nor UO_931 (O_931,N_4793,N_4010);
and UO_932 (O_932,N_4263,N_4794);
or UO_933 (O_933,N_4973,N_4401);
nor UO_934 (O_934,N_4368,N_4373);
nor UO_935 (O_935,N_4678,N_4841);
nand UO_936 (O_936,N_4728,N_4441);
or UO_937 (O_937,N_4219,N_4355);
nand UO_938 (O_938,N_4559,N_4778);
and UO_939 (O_939,N_4198,N_4008);
and UO_940 (O_940,N_4804,N_4571);
and UO_941 (O_941,N_4818,N_4033);
or UO_942 (O_942,N_4493,N_4192);
nor UO_943 (O_943,N_4390,N_4802);
and UO_944 (O_944,N_4312,N_4166);
nor UO_945 (O_945,N_4628,N_4110);
nor UO_946 (O_946,N_4034,N_4085);
and UO_947 (O_947,N_4447,N_4841);
nand UO_948 (O_948,N_4710,N_4303);
or UO_949 (O_949,N_4106,N_4793);
nor UO_950 (O_950,N_4863,N_4914);
nand UO_951 (O_951,N_4785,N_4025);
nand UO_952 (O_952,N_4578,N_4821);
nand UO_953 (O_953,N_4034,N_4802);
and UO_954 (O_954,N_4899,N_4104);
and UO_955 (O_955,N_4658,N_4243);
or UO_956 (O_956,N_4626,N_4681);
nor UO_957 (O_957,N_4459,N_4934);
and UO_958 (O_958,N_4283,N_4045);
nand UO_959 (O_959,N_4720,N_4419);
or UO_960 (O_960,N_4570,N_4840);
or UO_961 (O_961,N_4304,N_4276);
nor UO_962 (O_962,N_4097,N_4981);
nand UO_963 (O_963,N_4744,N_4086);
or UO_964 (O_964,N_4639,N_4195);
nor UO_965 (O_965,N_4407,N_4392);
or UO_966 (O_966,N_4076,N_4986);
nor UO_967 (O_967,N_4067,N_4476);
nor UO_968 (O_968,N_4698,N_4004);
nor UO_969 (O_969,N_4439,N_4412);
nor UO_970 (O_970,N_4910,N_4345);
nand UO_971 (O_971,N_4527,N_4892);
or UO_972 (O_972,N_4411,N_4287);
nand UO_973 (O_973,N_4167,N_4308);
nor UO_974 (O_974,N_4529,N_4727);
nand UO_975 (O_975,N_4959,N_4474);
and UO_976 (O_976,N_4532,N_4001);
and UO_977 (O_977,N_4514,N_4071);
or UO_978 (O_978,N_4329,N_4332);
nand UO_979 (O_979,N_4538,N_4179);
nor UO_980 (O_980,N_4589,N_4125);
nand UO_981 (O_981,N_4956,N_4299);
nand UO_982 (O_982,N_4686,N_4953);
and UO_983 (O_983,N_4819,N_4421);
nor UO_984 (O_984,N_4494,N_4230);
nand UO_985 (O_985,N_4580,N_4249);
or UO_986 (O_986,N_4558,N_4840);
or UO_987 (O_987,N_4604,N_4846);
nand UO_988 (O_988,N_4760,N_4045);
or UO_989 (O_989,N_4995,N_4495);
or UO_990 (O_990,N_4226,N_4481);
or UO_991 (O_991,N_4732,N_4107);
and UO_992 (O_992,N_4862,N_4534);
or UO_993 (O_993,N_4589,N_4912);
nor UO_994 (O_994,N_4423,N_4681);
and UO_995 (O_995,N_4054,N_4757);
nor UO_996 (O_996,N_4808,N_4875);
and UO_997 (O_997,N_4441,N_4039);
nand UO_998 (O_998,N_4963,N_4160);
nor UO_999 (O_999,N_4377,N_4334);
endmodule