module basic_500_3000_500_4_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_238,In_344);
xor U1 (N_1,In_29,In_169);
nor U2 (N_2,In_153,In_85);
nor U3 (N_3,In_39,In_413);
or U4 (N_4,In_218,In_480);
and U5 (N_5,In_307,In_204);
nor U6 (N_6,In_11,In_350);
nand U7 (N_7,In_15,In_224);
and U8 (N_8,In_314,In_200);
and U9 (N_9,In_320,In_405);
xnor U10 (N_10,In_410,In_117);
or U11 (N_11,In_371,In_287);
or U12 (N_12,In_354,In_68);
nor U13 (N_13,In_342,In_340);
nor U14 (N_14,In_103,In_404);
nand U15 (N_15,In_42,In_306);
nor U16 (N_16,In_156,In_245);
or U17 (N_17,In_319,In_32);
xor U18 (N_18,In_493,In_461);
and U19 (N_19,In_244,In_270);
or U20 (N_20,In_94,In_130);
or U21 (N_21,In_150,In_43);
xor U22 (N_22,In_122,In_34);
xnor U23 (N_23,In_358,In_106);
nand U24 (N_24,In_431,In_231);
nand U25 (N_25,In_330,In_72);
nand U26 (N_26,In_267,In_341);
xnor U27 (N_27,In_113,In_135);
nand U28 (N_28,In_22,In_456);
nor U29 (N_29,In_172,In_305);
or U30 (N_30,In_481,In_293);
or U31 (N_31,In_177,In_112);
and U32 (N_32,In_123,In_273);
or U33 (N_33,In_363,In_282);
or U34 (N_34,In_194,In_65);
nand U35 (N_35,In_451,In_284);
and U36 (N_36,In_274,In_47);
xnor U37 (N_37,In_375,In_151);
nand U38 (N_38,In_246,In_428);
nand U39 (N_39,In_66,In_271);
xnor U40 (N_40,In_285,In_120);
xnor U41 (N_41,In_323,In_1);
and U42 (N_42,In_18,In_230);
nor U43 (N_43,In_365,In_214);
or U44 (N_44,In_476,In_394);
nor U45 (N_45,In_91,In_116);
and U46 (N_46,In_381,In_102);
or U47 (N_47,In_191,In_392);
xnor U48 (N_48,In_118,In_168);
xor U49 (N_49,In_26,In_119);
xor U50 (N_50,In_115,In_356);
nor U51 (N_51,In_133,In_324);
xor U52 (N_52,In_260,In_304);
or U53 (N_53,In_69,In_425);
nor U54 (N_54,In_255,In_351);
nor U55 (N_55,In_455,In_128);
nand U56 (N_56,In_61,In_485);
nand U57 (N_57,In_166,In_23);
xnor U58 (N_58,In_209,In_417);
xor U59 (N_59,In_202,In_438);
nand U60 (N_60,In_373,In_429);
nand U61 (N_61,In_75,In_199);
and U62 (N_62,In_154,In_395);
and U63 (N_63,In_317,In_221);
or U64 (N_64,In_269,In_348);
and U65 (N_65,In_121,In_299);
and U66 (N_66,In_189,In_489);
xnor U67 (N_67,In_423,In_250);
or U68 (N_68,In_89,In_5);
xor U69 (N_69,In_100,In_460);
or U70 (N_70,In_334,In_328);
and U71 (N_71,In_445,In_60);
xor U72 (N_72,In_131,In_124);
xor U73 (N_73,In_316,In_25);
and U74 (N_74,In_162,In_452);
and U75 (N_75,In_170,In_297);
and U76 (N_76,In_152,In_37);
nand U77 (N_77,In_278,In_54);
nand U78 (N_78,In_12,In_275);
or U79 (N_79,In_418,In_402);
xnor U80 (N_80,In_84,In_302);
nand U81 (N_81,In_173,In_441);
nand U82 (N_82,In_474,In_242);
xnor U83 (N_83,In_176,In_80);
nand U84 (N_84,In_160,In_453);
nor U85 (N_85,In_19,In_36);
or U86 (N_86,In_276,In_74);
nand U87 (N_87,In_462,In_181);
or U88 (N_88,In_146,In_184);
and U89 (N_89,In_228,In_107);
xnor U90 (N_90,In_73,In_397);
nor U91 (N_91,In_440,In_56);
nor U92 (N_92,In_457,In_82);
or U93 (N_93,In_58,In_279);
nor U94 (N_94,In_187,In_213);
and U95 (N_95,In_303,In_175);
or U96 (N_96,In_399,In_9);
nor U97 (N_97,In_248,In_338);
and U98 (N_98,In_467,In_64);
and U99 (N_99,In_129,In_370);
or U100 (N_100,In_398,In_494);
nor U101 (N_101,In_207,In_468);
nand U102 (N_102,In_179,In_143);
xor U103 (N_103,In_497,In_163);
xnor U104 (N_104,In_157,In_300);
nor U105 (N_105,In_251,In_424);
nand U106 (N_106,In_329,In_262);
nor U107 (N_107,In_437,In_336);
xor U108 (N_108,In_450,In_111);
xnor U109 (N_109,In_24,In_290);
and U110 (N_110,In_28,In_426);
xor U111 (N_111,In_171,In_387);
nand U112 (N_112,In_70,In_27);
nand U113 (N_113,In_142,In_337);
or U114 (N_114,In_99,In_333);
nand U115 (N_115,In_280,In_235);
xor U116 (N_116,In_53,In_138);
and U117 (N_117,In_96,In_487);
xnor U118 (N_118,In_454,In_458);
or U119 (N_119,In_110,In_379);
nor U120 (N_120,In_174,In_491);
or U121 (N_121,In_471,In_7);
xor U122 (N_122,In_496,In_232);
nand U123 (N_123,In_51,In_374);
and U124 (N_124,In_478,In_436);
nand U125 (N_125,In_326,In_208);
and U126 (N_126,In_249,In_98);
or U127 (N_127,In_185,In_281);
nor U128 (N_128,In_407,In_40);
or U129 (N_129,In_132,In_470);
xor U130 (N_130,In_145,In_35);
or U131 (N_131,In_393,In_205);
xor U132 (N_132,In_109,In_352);
nor U133 (N_133,In_78,In_432);
and U134 (N_134,In_376,In_211);
nor U135 (N_135,In_186,In_97);
nand U136 (N_136,In_446,In_219);
nor U137 (N_137,In_366,In_391);
and U138 (N_138,In_400,In_155);
nand U139 (N_139,In_258,In_312);
nand U140 (N_140,In_93,In_38);
nor U141 (N_141,In_439,In_396);
xnor U142 (N_142,In_332,In_164);
nor U143 (N_143,In_222,In_447);
nand U144 (N_144,In_406,In_158);
nand U145 (N_145,In_147,In_292);
xor U146 (N_146,In_71,In_197);
or U147 (N_147,In_210,In_486);
and U148 (N_148,In_482,In_459);
and U149 (N_149,In_389,In_355);
and U150 (N_150,In_498,In_322);
xnor U151 (N_151,In_313,In_490);
xor U152 (N_152,In_20,In_144);
nand U153 (N_153,In_383,In_475);
nand U154 (N_154,In_63,In_477);
xor U155 (N_155,In_159,In_294);
or U156 (N_156,In_180,In_414);
or U157 (N_157,In_309,In_442);
nand U158 (N_158,In_412,In_443);
xor U159 (N_159,In_264,In_265);
nor U160 (N_160,In_101,In_421);
and U161 (N_161,In_263,In_335);
nor U162 (N_162,In_241,In_234);
nor U163 (N_163,In_295,In_401);
nand U164 (N_164,In_161,In_315);
or U165 (N_165,In_52,In_108);
xor U166 (N_166,In_464,In_465);
and U167 (N_167,In_268,In_422);
nand U168 (N_168,In_247,In_67);
xnor U169 (N_169,In_472,In_188);
nor U170 (N_170,In_367,In_165);
or U171 (N_171,In_45,In_237);
nand U172 (N_172,In_254,In_257);
nand U173 (N_173,In_499,In_347);
or U174 (N_174,In_83,In_41);
and U175 (N_175,In_55,In_4);
xnor U176 (N_176,In_149,In_362);
or U177 (N_177,In_349,In_484);
nand U178 (N_178,In_215,In_378);
or U179 (N_179,In_141,In_8);
nor U180 (N_180,In_140,In_372);
nor U181 (N_181,In_223,In_283);
nor U182 (N_182,In_385,In_206);
and U183 (N_183,In_88,In_291);
nand U184 (N_184,In_277,In_236);
and U185 (N_185,In_382,In_409);
and U186 (N_186,In_416,In_50);
and U187 (N_187,In_46,In_17);
or U188 (N_188,In_125,In_31);
nand U189 (N_189,In_311,In_325);
xnor U190 (N_190,In_105,In_148);
nor U191 (N_191,In_233,In_10);
nor U192 (N_192,In_427,In_220);
or U193 (N_193,In_403,In_30);
or U194 (N_194,In_377,In_380);
nand U195 (N_195,In_386,In_288);
nand U196 (N_196,In_196,In_256);
or U197 (N_197,In_448,In_167);
and U198 (N_198,In_126,In_243);
xor U199 (N_199,In_14,In_466);
nor U200 (N_200,In_227,In_79);
nor U201 (N_201,In_369,In_343);
nand U202 (N_202,In_87,In_339);
nor U203 (N_203,In_104,In_321);
and U204 (N_204,In_479,In_252);
nand U205 (N_205,In_253,In_21);
nor U206 (N_206,In_388,In_76);
nor U207 (N_207,In_361,In_81);
xor U208 (N_208,In_212,In_239);
and U209 (N_209,In_318,In_327);
nor U210 (N_210,In_137,In_48);
nor U211 (N_211,In_216,In_433);
nand U212 (N_212,In_44,In_16);
nor U213 (N_213,In_408,In_178);
nor U214 (N_214,In_259,In_198);
nand U215 (N_215,In_310,In_286);
nand U216 (N_216,In_331,In_415);
xor U217 (N_217,In_359,In_308);
nand U218 (N_218,In_33,In_0);
nand U219 (N_219,In_345,In_49);
and U220 (N_220,In_463,In_201);
nand U221 (N_221,In_59,In_420);
or U222 (N_222,In_353,In_357);
and U223 (N_223,In_217,In_2);
or U224 (N_224,In_469,In_368);
nand U225 (N_225,In_190,In_240);
nand U226 (N_226,In_13,In_272);
nand U227 (N_227,In_261,In_488);
or U228 (N_228,In_492,In_229);
or U229 (N_229,In_298,In_127);
or U230 (N_230,In_225,In_90);
and U231 (N_231,In_289,In_296);
nor U232 (N_232,In_483,In_390);
nor U233 (N_233,In_360,In_346);
and U234 (N_234,In_444,In_6);
nand U235 (N_235,In_77,In_57);
or U236 (N_236,In_495,In_193);
or U237 (N_237,In_92,In_434);
and U238 (N_238,In_203,In_136);
nand U239 (N_239,In_114,In_411);
and U240 (N_240,In_419,In_62);
or U241 (N_241,In_195,In_449);
or U242 (N_242,In_183,In_3);
xor U243 (N_243,In_134,In_192);
xor U244 (N_244,In_139,In_182);
xor U245 (N_245,In_435,In_364);
or U246 (N_246,In_430,In_301);
nand U247 (N_247,In_384,In_226);
and U248 (N_248,In_473,In_95);
nor U249 (N_249,In_266,In_86);
nor U250 (N_250,In_330,In_6);
xnor U251 (N_251,In_260,In_22);
nand U252 (N_252,In_458,In_169);
xnor U253 (N_253,In_146,In_429);
and U254 (N_254,In_453,In_490);
nor U255 (N_255,In_483,In_258);
xnor U256 (N_256,In_200,In_117);
nand U257 (N_257,In_223,In_147);
nor U258 (N_258,In_181,In_285);
or U259 (N_259,In_178,In_108);
nand U260 (N_260,In_89,In_143);
nand U261 (N_261,In_479,In_142);
or U262 (N_262,In_9,In_294);
and U263 (N_263,In_52,In_467);
nand U264 (N_264,In_1,In_84);
xnor U265 (N_265,In_386,In_188);
xnor U266 (N_266,In_386,In_366);
nand U267 (N_267,In_360,In_322);
nand U268 (N_268,In_118,In_388);
or U269 (N_269,In_405,In_312);
nor U270 (N_270,In_256,In_428);
and U271 (N_271,In_298,In_192);
xnor U272 (N_272,In_399,In_299);
or U273 (N_273,In_116,In_314);
xor U274 (N_274,In_169,In_129);
nand U275 (N_275,In_35,In_191);
xor U276 (N_276,In_482,In_282);
nor U277 (N_277,In_497,In_130);
or U278 (N_278,In_29,In_51);
nor U279 (N_279,In_295,In_337);
nand U280 (N_280,In_357,In_473);
or U281 (N_281,In_66,In_398);
nor U282 (N_282,In_435,In_233);
and U283 (N_283,In_250,In_254);
and U284 (N_284,In_448,In_146);
and U285 (N_285,In_424,In_191);
and U286 (N_286,In_203,In_439);
or U287 (N_287,In_448,In_332);
xor U288 (N_288,In_123,In_188);
nand U289 (N_289,In_228,In_231);
and U290 (N_290,In_32,In_488);
and U291 (N_291,In_465,In_98);
or U292 (N_292,In_391,In_472);
and U293 (N_293,In_130,In_123);
and U294 (N_294,In_334,In_391);
or U295 (N_295,In_428,In_475);
nand U296 (N_296,In_139,In_405);
nand U297 (N_297,In_35,In_7);
nor U298 (N_298,In_186,In_222);
nand U299 (N_299,In_43,In_459);
xor U300 (N_300,In_40,In_480);
or U301 (N_301,In_173,In_350);
and U302 (N_302,In_99,In_301);
nor U303 (N_303,In_419,In_126);
nor U304 (N_304,In_215,In_344);
xnor U305 (N_305,In_298,In_352);
nand U306 (N_306,In_140,In_157);
nand U307 (N_307,In_178,In_202);
nand U308 (N_308,In_189,In_13);
or U309 (N_309,In_180,In_424);
xor U310 (N_310,In_51,In_433);
nor U311 (N_311,In_445,In_468);
or U312 (N_312,In_204,In_358);
and U313 (N_313,In_79,In_308);
xnor U314 (N_314,In_225,In_367);
nand U315 (N_315,In_102,In_224);
or U316 (N_316,In_111,In_325);
and U317 (N_317,In_79,In_415);
or U318 (N_318,In_164,In_404);
nand U319 (N_319,In_223,In_134);
nand U320 (N_320,In_336,In_68);
xor U321 (N_321,In_243,In_90);
or U322 (N_322,In_328,In_356);
or U323 (N_323,In_60,In_400);
and U324 (N_324,In_412,In_195);
and U325 (N_325,In_256,In_438);
nor U326 (N_326,In_32,In_431);
and U327 (N_327,In_89,In_144);
or U328 (N_328,In_448,In_403);
nor U329 (N_329,In_488,In_168);
or U330 (N_330,In_498,In_321);
nand U331 (N_331,In_74,In_0);
nand U332 (N_332,In_413,In_430);
and U333 (N_333,In_29,In_415);
nand U334 (N_334,In_498,In_409);
xnor U335 (N_335,In_147,In_461);
nor U336 (N_336,In_348,In_130);
or U337 (N_337,In_490,In_483);
or U338 (N_338,In_177,In_361);
xor U339 (N_339,In_135,In_123);
or U340 (N_340,In_433,In_317);
xnor U341 (N_341,In_344,In_190);
xnor U342 (N_342,In_498,In_408);
nor U343 (N_343,In_230,In_163);
nand U344 (N_344,In_132,In_3);
xnor U345 (N_345,In_170,In_480);
and U346 (N_346,In_366,In_71);
nor U347 (N_347,In_269,In_496);
nor U348 (N_348,In_474,In_488);
nand U349 (N_349,In_192,In_498);
nor U350 (N_350,In_135,In_103);
xnor U351 (N_351,In_183,In_370);
or U352 (N_352,In_244,In_282);
xor U353 (N_353,In_373,In_70);
nor U354 (N_354,In_17,In_372);
nand U355 (N_355,In_164,In_34);
or U356 (N_356,In_257,In_285);
and U357 (N_357,In_4,In_299);
and U358 (N_358,In_52,In_242);
and U359 (N_359,In_342,In_468);
nand U360 (N_360,In_281,In_393);
or U361 (N_361,In_418,In_375);
or U362 (N_362,In_439,In_369);
or U363 (N_363,In_382,In_364);
and U364 (N_364,In_310,In_407);
and U365 (N_365,In_113,In_104);
nor U366 (N_366,In_284,In_218);
nand U367 (N_367,In_450,In_33);
or U368 (N_368,In_400,In_448);
and U369 (N_369,In_62,In_105);
xor U370 (N_370,In_460,In_83);
xnor U371 (N_371,In_435,In_52);
nand U372 (N_372,In_391,In_149);
or U373 (N_373,In_52,In_331);
or U374 (N_374,In_326,In_319);
or U375 (N_375,In_365,In_224);
nor U376 (N_376,In_153,In_335);
xnor U377 (N_377,In_212,In_96);
nor U378 (N_378,In_268,In_95);
or U379 (N_379,In_235,In_29);
xnor U380 (N_380,In_209,In_240);
nor U381 (N_381,In_73,In_268);
nand U382 (N_382,In_476,In_250);
nor U383 (N_383,In_16,In_58);
and U384 (N_384,In_274,In_183);
and U385 (N_385,In_260,In_348);
and U386 (N_386,In_456,In_232);
or U387 (N_387,In_368,In_58);
xor U388 (N_388,In_198,In_386);
xor U389 (N_389,In_380,In_381);
nor U390 (N_390,In_118,In_175);
xor U391 (N_391,In_490,In_357);
or U392 (N_392,In_370,In_1);
nor U393 (N_393,In_475,In_92);
xnor U394 (N_394,In_347,In_321);
nor U395 (N_395,In_282,In_399);
and U396 (N_396,In_320,In_341);
nor U397 (N_397,In_40,In_95);
xor U398 (N_398,In_103,In_259);
nand U399 (N_399,In_434,In_322);
nand U400 (N_400,In_91,In_499);
nand U401 (N_401,In_200,In_85);
xnor U402 (N_402,In_363,In_208);
and U403 (N_403,In_94,In_113);
nor U404 (N_404,In_266,In_416);
nor U405 (N_405,In_180,In_497);
and U406 (N_406,In_265,In_345);
xor U407 (N_407,In_100,In_98);
and U408 (N_408,In_390,In_52);
nand U409 (N_409,In_77,In_269);
nor U410 (N_410,In_101,In_345);
or U411 (N_411,In_196,In_157);
xor U412 (N_412,In_148,In_330);
nor U413 (N_413,In_272,In_197);
and U414 (N_414,In_176,In_293);
nand U415 (N_415,In_381,In_446);
nor U416 (N_416,In_268,In_430);
and U417 (N_417,In_446,In_350);
nor U418 (N_418,In_73,In_130);
nor U419 (N_419,In_401,In_224);
and U420 (N_420,In_37,In_61);
xnor U421 (N_421,In_419,In_363);
and U422 (N_422,In_493,In_388);
xor U423 (N_423,In_354,In_401);
nand U424 (N_424,In_497,In_153);
nand U425 (N_425,In_7,In_422);
xor U426 (N_426,In_156,In_3);
nand U427 (N_427,In_278,In_97);
xor U428 (N_428,In_243,In_51);
xnor U429 (N_429,In_450,In_427);
nand U430 (N_430,In_178,In_414);
or U431 (N_431,In_373,In_323);
nand U432 (N_432,In_200,In_175);
nand U433 (N_433,In_453,In_38);
nor U434 (N_434,In_8,In_496);
xnor U435 (N_435,In_33,In_20);
xnor U436 (N_436,In_232,In_199);
xnor U437 (N_437,In_342,In_366);
nand U438 (N_438,In_197,In_302);
nand U439 (N_439,In_217,In_103);
and U440 (N_440,In_443,In_441);
nand U441 (N_441,In_240,In_212);
and U442 (N_442,In_214,In_412);
nor U443 (N_443,In_49,In_147);
nand U444 (N_444,In_42,In_470);
nor U445 (N_445,In_393,In_138);
and U446 (N_446,In_292,In_421);
nor U447 (N_447,In_47,In_133);
nand U448 (N_448,In_293,In_23);
xnor U449 (N_449,In_176,In_15);
and U450 (N_450,In_195,In_339);
nand U451 (N_451,In_397,In_245);
and U452 (N_452,In_200,In_436);
nand U453 (N_453,In_107,In_241);
nand U454 (N_454,In_310,In_333);
or U455 (N_455,In_480,In_393);
or U456 (N_456,In_479,In_205);
and U457 (N_457,In_382,In_233);
or U458 (N_458,In_138,In_446);
or U459 (N_459,In_130,In_227);
nand U460 (N_460,In_352,In_475);
xnor U461 (N_461,In_413,In_142);
nor U462 (N_462,In_36,In_349);
xnor U463 (N_463,In_321,In_158);
or U464 (N_464,In_17,In_120);
xnor U465 (N_465,In_136,In_28);
nor U466 (N_466,In_84,In_307);
and U467 (N_467,In_142,In_426);
nor U468 (N_468,In_349,In_83);
nor U469 (N_469,In_394,In_3);
or U470 (N_470,In_477,In_443);
and U471 (N_471,In_55,In_184);
nor U472 (N_472,In_436,In_231);
nor U473 (N_473,In_146,In_472);
and U474 (N_474,In_285,In_91);
nor U475 (N_475,In_206,In_405);
xnor U476 (N_476,In_196,In_478);
nand U477 (N_477,In_260,In_487);
xnor U478 (N_478,In_98,In_151);
or U479 (N_479,In_272,In_67);
and U480 (N_480,In_497,In_186);
and U481 (N_481,In_188,In_92);
xnor U482 (N_482,In_259,In_123);
xor U483 (N_483,In_186,In_395);
nand U484 (N_484,In_344,In_56);
xor U485 (N_485,In_72,In_491);
nand U486 (N_486,In_465,In_11);
xor U487 (N_487,In_330,In_34);
xor U488 (N_488,In_235,In_320);
or U489 (N_489,In_452,In_83);
and U490 (N_490,In_405,In_496);
or U491 (N_491,In_385,In_247);
nor U492 (N_492,In_179,In_322);
xnor U493 (N_493,In_168,In_342);
and U494 (N_494,In_227,In_87);
nor U495 (N_495,In_200,In_154);
or U496 (N_496,In_481,In_178);
xnor U497 (N_497,In_206,In_299);
xnor U498 (N_498,In_320,In_240);
xnor U499 (N_499,In_146,In_36);
and U500 (N_500,In_104,In_305);
or U501 (N_501,In_17,In_189);
nor U502 (N_502,In_429,In_472);
xnor U503 (N_503,In_106,In_433);
nor U504 (N_504,In_497,In_139);
xnor U505 (N_505,In_287,In_318);
or U506 (N_506,In_117,In_441);
and U507 (N_507,In_487,In_405);
nor U508 (N_508,In_264,In_348);
nand U509 (N_509,In_405,In_240);
or U510 (N_510,In_309,In_18);
nor U511 (N_511,In_103,In_224);
and U512 (N_512,In_232,In_13);
nor U513 (N_513,In_372,In_492);
or U514 (N_514,In_362,In_428);
or U515 (N_515,In_430,In_443);
and U516 (N_516,In_195,In_367);
nor U517 (N_517,In_54,In_466);
xor U518 (N_518,In_379,In_369);
nand U519 (N_519,In_278,In_3);
and U520 (N_520,In_125,In_309);
nand U521 (N_521,In_241,In_365);
xnor U522 (N_522,In_205,In_125);
nand U523 (N_523,In_307,In_2);
and U524 (N_524,In_22,In_315);
nand U525 (N_525,In_267,In_100);
or U526 (N_526,In_7,In_88);
or U527 (N_527,In_179,In_45);
or U528 (N_528,In_198,In_104);
nor U529 (N_529,In_153,In_20);
and U530 (N_530,In_90,In_454);
and U531 (N_531,In_420,In_442);
nor U532 (N_532,In_384,In_391);
nand U533 (N_533,In_363,In_306);
or U534 (N_534,In_364,In_428);
xnor U535 (N_535,In_413,In_366);
or U536 (N_536,In_115,In_207);
or U537 (N_537,In_105,In_205);
and U538 (N_538,In_176,In_433);
xnor U539 (N_539,In_327,In_33);
xor U540 (N_540,In_179,In_308);
nand U541 (N_541,In_317,In_458);
or U542 (N_542,In_134,In_271);
and U543 (N_543,In_463,In_102);
xnor U544 (N_544,In_203,In_238);
nor U545 (N_545,In_409,In_167);
or U546 (N_546,In_60,In_206);
nand U547 (N_547,In_315,In_94);
xor U548 (N_548,In_227,In_40);
nor U549 (N_549,In_391,In_283);
nand U550 (N_550,In_205,In_95);
xor U551 (N_551,In_186,In_361);
or U552 (N_552,In_450,In_285);
nand U553 (N_553,In_150,In_205);
and U554 (N_554,In_51,In_173);
nand U555 (N_555,In_185,In_461);
nand U556 (N_556,In_18,In_494);
and U557 (N_557,In_354,In_378);
or U558 (N_558,In_33,In_79);
nand U559 (N_559,In_184,In_491);
or U560 (N_560,In_93,In_301);
or U561 (N_561,In_200,In_34);
nor U562 (N_562,In_95,In_400);
xnor U563 (N_563,In_206,In_366);
xor U564 (N_564,In_432,In_41);
and U565 (N_565,In_406,In_169);
and U566 (N_566,In_318,In_415);
nor U567 (N_567,In_398,In_421);
nand U568 (N_568,In_55,In_0);
xnor U569 (N_569,In_274,In_60);
nor U570 (N_570,In_290,In_82);
and U571 (N_571,In_337,In_305);
nor U572 (N_572,In_18,In_33);
xor U573 (N_573,In_105,In_444);
or U574 (N_574,In_263,In_286);
xor U575 (N_575,In_64,In_196);
nor U576 (N_576,In_80,In_218);
and U577 (N_577,In_412,In_268);
xnor U578 (N_578,In_288,In_376);
or U579 (N_579,In_245,In_197);
and U580 (N_580,In_248,In_196);
and U581 (N_581,In_317,In_257);
nor U582 (N_582,In_431,In_21);
xnor U583 (N_583,In_164,In_51);
nand U584 (N_584,In_454,In_257);
nor U585 (N_585,In_276,In_354);
and U586 (N_586,In_116,In_264);
xor U587 (N_587,In_277,In_62);
or U588 (N_588,In_304,In_401);
and U589 (N_589,In_248,In_135);
nor U590 (N_590,In_146,In_60);
xnor U591 (N_591,In_174,In_67);
and U592 (N_592,In_219,In_223);
and U593 (N_593,In_251,In_183);
xor U594 (N_594,In_324,In_179);
xor U595 (N_595,In_467,In_101);
nor U596 (N_596,In_407,In_367);
or U597 (N_597,In_366,In_138);
and U598 (N_598,In_382,In_129);
xnor U599 (N_599,In_264,In_315);
nor U600 (N_600,In_358,In_57);
nor U601 (N_601,In_257,In_325);
xnor U602 (N_602,In_143,In_49);
and U603 (N_603,In_396,In_235);
xnor U604 (N_604,In_431,In_366);
and U605 (N_605,In_457,In_473);
nand U606 (N_606,In_238,In_230);
xor U607 (N_607,In_121,In_282);
and U608 (N_608,In_345,In_58);
nor U609 (N_609,In_41,In_55);
or U610 (N_610,In_135,In_64);
and U611 (N_611,In_85,In_121);
and U612 (N_612,In_326,In_340);
and U613 (N_613,In_233,In_473);
or U614 (N_614,In_418,In_237);
nor U615 (N_615,In_282,In_390);
nand U616 (N_616,In_30,In_404);
nand U617 (N_617,In_4,In_183);
or U618 (N_618,In_266,In_143);
or U619 (N_619,In_364,In_224);
and U620 (N_620,In_496,In_142);
and U621 (N_621,In_78,In_483);
nand U622 (N_622,In_8,In_19);
nand U623 (N_623,In_370,In_10);
nand U624 (N_624,In_274,In_354);
xnor U625 (N_625,In_346,In_287);
and U626 (N_626,In_305,In_286);
and U627 (N_627,In_146,In_212);
and U628 (N_628,In_429,In_302);
nor U629 (N_629,In_102,In_419);
or U630 (N_630,In_100,In_75);
xor U631 (N_631,In_459,In_201);
xor U632 (N_632,In_456,In_406);
or U633 (N_633,In_169,In_290);
and U634 (N_634,In_378,In_364);
nor U635 (N_635,In_361,In_477);
and U636 (N_636,In_251,In_475);
or U637 (N_637,In_171,In_294);
or U638 (N_638,In_280,In_362);
or U639 (N_639,In_473,In_137);
xor U640 (N_640,In_265,In_246);
and U641 (N_641,In_356,In_441);
nand U642 (N_642,In_234,In_68);
and U643 (N_643,In_351,In_397);
xnor U644 (N_644,In_217,In_480);
and U645 (N_645,In_372,In_155);
nor U646 (N_646,In_197,In_404);
nand U647 (N_647,In_41,In_186);
nor U648 (N_648,In_387,In_428);
nand U649 (N_649,In_334,In_29);
nor U650 (N_650,In_105,In_18);
and U651 (N_651,In_388,In_308);
xor U652 (N_652,In_354,In_240);
nor U653 (N_653,In_390,In_252);
xor U654 (N_654,In_71,In_358);
nand U655 (N_655,In_79,In_27);
xnor U656 (N_656,In_152,In_41);
and U657 (N_657,In_290,In_175);
and U658 (N_658,In_274,In_146);
nand U659 (N_659,In_201,In_438);
xnor U660 (N_660,In_60,In_423);
or U661 (N_661,In_206,In_115);
nor U662 (N_662,In_270,In_59);
nor U663 (N_663,In_392,In_70);
xnor U664 (N_664,In_308,In_2);
nor U665 (N_665,In_59,In_291);
or U666 (N_666,In_380,In_121);
and U667 (N_667,In_496,In_328);
nor U668 (N_668,In_4,In_81);
and U669 (N_669,In_422,In_395);
nand U670 (N_670,In_64,In_203);
or U671 (N_671,In_313,In_86);
and U672 (N_672,In_4,In_404);
nor U673 (N_673,In_76,In_17);
nand U674 (N_674,In_241,In_482);
xor U675 (N_675,In_162,In_139);
nand U676 (N_676,In_483,In_220);
nand U677 (N_677,In_497,In_34);
or U678 (N_678,In_125,In_103);
xnor U679 (N_679,In_5,In_90);
or U680 (N_680,In_336,In_80);
nand U681 (N_681,In_430,In_120);
nand U682 (N_682,In_301,In_31);
xor U683 (N_683,In_108,In_444);
or U684 (N_684,In_298,In_249);
nor U685 (N_685,In_405,In_301);
nand U686 (N_686,In_337,In_309);
or U687 (N_687,In_125,In_377);
nand U688 (N_688,In_393,In_349);
nor U689 (N_689,In_245,In_354);
nand U690 (N_690,In_495,In_150);
nor U691 (N_691,In_220,In_332);
nand U692 (N_692,In_455,In_254);
and U693 (N_693,In_291,In_241);
xor U694 (N_694,In_68,In_493);
nor U695 (N_695,In_100,In_111);
nand U696 (N_696,In_129,In_107);
nor U697 (N_697,In_288,In_197);
nand U698 (N_698,In_478,In_445);
nor U699 (N_699,In_296,In_303);
nand U700 (N_700,In_422,In_325);
or U701 (N_701,In_269,In_67);
xor U702 (N_702,In_385,In_315);
xnor U703 (N_703,In_109,In_72);
xnor U704 (N_704,In_111,In_176);
nor U705 (N_705,In_460,In_180);
xnor U706 (N_706,In_483,In_212);
nand U707 (N_707,In_82,In_347);
nand U708 (N_708,In_137,In_335);
nor U709 (N_709,In_132,In_493);
xnor U710 (N_710,In_409,In_18);
nor U711 (N_711,In_293,In_150);
nor U712 (N_712,In_108,In_17);
or U713 (N_713,In_323,In_311);
and U714 (N_714,In_344,In_284);
nand U715 (N_715,In_356,In_393);
nand U716 (N_716,In_106,In_129);
nor U717 (N_717,In_460,In_227);
or U718 (N_718,In_373,In_24);
nor U719 (N_719,In_178,In_303);
xor U720 (N_720,In_246,In_251);
xor U721 (N_721,In_388,In_386);
or U722 (N_722,In_149,In_250);
nor U723 (N_723,In_400,In_464);
nor U724 (N_724,In_466,In_76);
nand U725 (N_725,In_318,In_400);
nand U726 (N_726,In_261,In_291);
xnor U727 (N_727,In_259,In_104);
nand U728 (N_728,In_357,In_395);
or U729 (N_729,In_494,In_24);
nand U730 (N_730,In_169,In_213);
xnor U731 (N_731,In_237,In_379);
nand U732 (N_732,In_42,In_232);
nor U733 (N_733,In_334,In_332);
nor U734 (N_734,In_165,In_414);
and U735 (N_735,In_235,In_88);
or U736 (N_736,In_103,In_132);
xnor U737 (N_737,In_266,In_57);
and U738 (N_738,In_77,In_118);
xnor U739 (N_739,In_226,In_291);
or U740 (N_740,In_197,In_279);
nand U741 (N_741,In_369,In_44);
and U742 (N_742,In_440,In_372);
nand U743 (N_743,In_178,In_52);
or U744 (N_744,In_250,In_59);
and U745 (N_745,In_494,In_161);
nor U746 (N_746,In_242,In_396);
or U747 (N_747,In_463,In_402);
xor U748 (N_748,In_106,In_105);
nand U749 (N_749,In_361,In_317);
and U750 (N_750,N_176,N_705);
xor U751 (N_751,N_174,N_560);
or U752 (N_752,N_462,N_434);
or U753 (N_753,N_335,N_652);
nand U754 (N_754,N_233,N_733);
and U755 (N_755,N_115,N_490);
or U756 (N_756,N_193,N_619);
or U757 (N_757,N_232,N_119);
xor U758 (N_758,N_295,N_410);
xor U759 (N_759,N_53,N_3);
or U760 (N_760,N_707,N_363);
nor U761 (N_761,N_469,N_573);
xor U762 (N_762,N_63,N_708);
or U763 (N_763,N_664,N_314);
and U764 (N_764,N_442,N_109);
or U765 (N_765,N_575,N_535);
xor U766 (N_766,N_268,N_431);
nand U767 (N_767,N_501,N_320);
and U768 (N_768,N_595,N_5);
or U769 (N_769,N_99,N_608);
nor U770 (N_770,N_383,N_325);
and U771 (N_771,N_220,N_148);
nor U772 (N_772,N_130,N_355);
nor U773 (N_773,N_533,N_31);
xor U774 (N_774,N_513,N_161);
and U775 (N_775,N_646,N_588);
xor U776 (N_776,N_550,N_509);
or U777 (N_777,N_321,N_379);
xor U778 (N_778,N_6,N_522);
or U779 (N_779,N_480,N_275);
and U780 (N_780,N_329,N_444);
xnor U781 (N_781,N_475,N_629);
or U782 (N_782,N_61,N_242);
xnor U783 (N_783,N_504,N_553);
or U784 (N_784,N_391,N_514);
xnor U785 (N_785,N_178,N_74);
and U786 (N_786,N_145,N_36);
or U787 (N_787,N_559,N_428);
xnor U788 (N_788,N_389,N_173);
and U789 (N_789,N_32,N_19);
or U790 (N_790,N_67,N_365);
xnor U791 (N_791,N_191,N_357);
nand U792 (N_792,N_223,N_638);
and U793 (N_793,N_582,N_603);
nand U794 (N_794,N_590,N_76);
nand U795 (N_795,N_437,N_485);
xor U796 (N_796,N_134,N_579);
and U797 (N_797,N_616,N_257);
or U798 (N_798,N_40,N_461);
nand U799 (N_799,N_517,N_286);
xor U800 (N_800,N_135,N_746);
and U801 (N_801,N_448,N_453);
nand U802 (N_802,N_584,N_373);
or U803 (N_803,N_278,N_68);
or U804 (N_804,N_88,N_250);
nand U805 (N_805,N_150,N_179);
nor U806 (N_806,N_370,N_709);
nor U807 (N_807,N_665,N_388);
and U808 (N_808,N_537,N_287);
nor U809 (N_809,N_11,N_626);
xor U810 (N_810,N_123,N_185);
and U811 (N_811,N_393,N_308);
and U812 (N_812,N_503,N_65);
and U813 (N_813,N_152,N_15);
xnor U814 (N_814,N_244,N_92);
xor U815 (N_815,N_79,N_49);
or U816 (N_816,N_228,N_613);
nand U817 (N_817,N_743,N_731);
and U818 (N_818,N_649,N_378);
nand U819 (N_819,N_341,N_104);
xnor U820 (N_820,N_112,N_467);
nor U821 (N_821,N_634,N_127);
xnor U822 (N_822,N_77,N_455);
and U823 (N_823,N_269,N_85);
or U824 (N_824,N_133,N_201);
xnor U825 (N_825,N_103,N_310);
xnor U826 (N_826,N_489,N_668);
and U827 (N_827,N_139,N_396);
nand U828 (N_828,N_24,N_345);
nand U829 (N_829,N_532,N_691);
or U830 (N_830,N_549,N_336);
nand U831 (N_831,N_449,N_422);
or U832 (N_832,N_202,N_194);
or U833 (N_833,N_471,N_238);
or U834 (N_834,N_83,N_203);
and U835 (N_835,N_254,N_234);
and U836 (N_836,N_372,N_331);
nand U837 (N_837,N_399,N_420);
or U838 (N_838,N_165,N_33);
or U839 (N_839,N_235,N_27);
nand U840 (N_840,N_439,N_62);
and U841 (N_841,N_452,N_280);
nor U842 (N_842,N_277,N_168);
and U843 (N_843,N_407,N_270);
nor U844 (N_844,N_690,N_673);
and U845 (N_845,N_657,N_474);
nor U846 (N_846,N_229,N_730);
or U847 (N_847,N_742,N_218);
nand U848 (N_848,N_23,N_720);
xor U849 (N_849,N_230,N_339);
nor U850 (N_850,N_264,N_632);
and U851 (N_851,N_326,N_231);
xnor U852 (N_852,N_481,N_576);
or U853 (N_853,N_156,N_351);
nor U854 (N_854,N_566,N_35);
nand U855 (N_855,N_398,N_546);
xor U856 (N_856,N_122,N_248);
or U857 (N_857,N_205,N_246);
nor U858 (N_858,N_618,N_368);
or U859 (N_859,N_98,N_221);
or U860 (N_860,N_574,N_728);
or U861 (N_861,N_450,N_186);
and U862 (N_862,N_492,N_682);
nor U863 (N_863,N_536,N_643);
nand U864 (N_864,N_96,N_146);
nand U865 (N_865,N_157,N_412);
xor U866 (N_866,N_95,N_506);
nand U867 (N_867,N_600,N_674);
nor U868 (N_868,N_208,N_581);
and U869 (N_869,N_713,N_463);
xor U870 (N_870,N_362,N_408);
nand U871 (N_871,N_556,N_592);
xor U872 (N_872,N_494,N_51);
xnor U873 (N_873,N_294,N_18);
nor U874 (N_874,N_531,N_188);
nand U875 (N_875,N_89,N_525);
or U876 (N_876,N_245,N_596);
and U877 (N_877,N_43,N_240);
or U878 (N_878,N_170,N_631);
xnor U879 (N_879,N_587,N_128);
and U880 (N_880,N_374,N_526);
nor U881 (N_881,N_361,N_360);
nor U882 (N_882,N_255,N_712);
or U883 (N_883,N_521,N_432);
xnor U884 (N_884,N_628,N_117);
or U885 (N_885,N_411,N_710);
nor U886 (N_886,N_554,N_344);
xor U887 (N_887,N_171,N_296);
nor U888 (N_888,N_736,N_679);
or U889 (N_889,N_583,N_349);
nor U890 (N_890,N_495,N_660);
nor U891 (N_891,N_538,N_256);
and U892 (N_892,N_266,N_721);
or U893 (N_893,N_25,N_441);
and U894 (N_894,N_624,N_675);
nand U895 (N_895,N_395,N_702);
nor U896 (N_896,N_209,N_650);
nor U897 (N_897,N_570,N_272);
xor U898 (N_898,N_153,N_327);
nand U899 (N_899,N_252,N_22);
xnor U900 (N_900,N_94,N_283);
nand U901 (N_901,N_580,N_50);
nand U902 (N_902,N_376,N_358);
xor U903 (N_903,N_493,N_100);
and U904 (N_904,N_0,N_260);
or U905 (N_905,N_10,N_507);
nor U906 (N_906,N_164,N_45);
and U907 (N_907,N_73,N_671);
xor U908 (N_908,N_540,N_367);
nor U909 (N_909,N_177,N_741);
and U910 (N_910,N_21,N_158);
and U911 (N_911,N_703,N_167);
xor U912 (N_912,N_732,N_542);
xor U913 (N_913,N_118,N_38);
nand U914 (N_914,N_593,N_9);
nand U915 (N_915,N_440,N_182);
and U916 (N_916,N_738,N_445);
or U917 (N_917,N_686,N_669);
or U918 (N_918,N_416,N_175);
nand U919 (N_919,N_488,N_384);
or U920 (N_920,N_464,N_359);
xnor U921 (N_921,N_635,N_694);
nor U922 (N_922,N_353,N_381);
or U923 (N_923,N_567,N_500);
xnor U924 (N_924,N_747,N_28);
or U925 (N_925,N_421,N_315);
xor U926 (N_926,N_371,N_54);
nor U927 (N_927,N_338,N_701);
nor U928 (N_928,N_42,N_419);
nor U929 (N_929,N_143,N_297);
nand U930 (N_930,N_217,N_267);
nor U931 (N_931,N_499,N_337);
nand U932 (N_932,N_636,N_447);
nand U933 (N_933,N_505,N_274);
xnor U934 (N_934,N_529,N_627);
nand U935 (N_935,N_71,N_400);
nand U936 (N_936,N_312,N_633);
or U937 (N_937,N_639,N_433);
xnor U938 (N_938,N_527,N_700);
or U939 (N_939,N_334,N_216);
xnor U940 (N_940,N_496,N_647);
nor U941 (N_941,N_438,N_190);
nor U942 (N_942,N_685,N_642);
and U943 (N_943,N_734,N_166);
and U944 (N_944,N_259,N_564);
nor U945 (N_945,N_594,N_75);
and U946 (N_946,N_443,N_90);
or U947 (N_947,N_313,N_317);
nand U948 (N_948,N_409,N_697);
and U949 (N_949,N_680,N_615);
nor U950 (N_950,N_102,N_215);
or U951 (N_951,N_451,N_343);
nor U952 (N_952,N_472,N_465);
xnor U953 (N_953,N_716,N_219);
and U954 (N_954,N_565,N_403);
nand U955 (N_955,N_199,N_136);
and U956 (N_956,N_387,N_693);
nand U957 (N_957,N_670,N_429);
nor U958 (N_958,N_298,N_291);
nor U959 (N_959,N_704,N_58);
nand U960 (N_960,N_249,N_107);
nor U961 (N_961,N_607,N_749);
nor U962 (N_962,N_539,N_591);
or U963 (N_963,N_124,N_160);
nor U964 (N_964,N_617,N_140);
or U965 (N_965,N_319,N_692);
xor U966 (N_966,N_159,N_460);
xor U967 (N_967,N_585,N_557);
or U968 (N_968,N_484,N_210);
nor U969 (N_969,N_423,N_604);
nand U970 (N_970,N_273,N_149);
nand U971 (N_971,N_677,N_237);
xnor U972 (N_972,N_189,N_404);
xor U973 (N_973,N_612,N_198);
xor U974 (N_974,N_477,N_645);
or U975 (N_975,N_282,N_727);
and U976 (N_976,N_470,N_436);
xor U977 (N_977,N_289,N_147);
and U978 (N_978,N_2,N_309);
and U979 (N_979,N_7,N_426);
xnor U980 (N_980,N_29,N_333);
nand U981 (N_981,N_518,N_390);
and U982 (N_982,N_302,N_108);
or U983 (N_983,N_288,N_456);
xor U984 (N_984,N_516,N_316);
nor U985 (N_985,N_578,N_551);
and U986 (N_986,N_623,N_226);
or U987 (N_987,N_224,N_508);
and U988 (N_988,N_430,N_91);
nand U989 (N_989,N_279,N_356);
or U990 (N_990,N_60,N_12);
nor U991 (N_991,N_744,N_37);
nor U992 (N_992,N_78,N_597);
xor U993 (N_993,N_719,N_724);
nand U994 (N_994,N_323,N_586);
nand U995 (N_995,N_726,N_722);
xor U996 (N_996,N_41,N_547);
xor U997 (N_997,N_459,N_487);
nand U998 (N_998,N_662,N_328);
xnor U999 (N_999,N_364,N_666);
or U1000 (N_1000,N_8,N_180);
nor U1001 (N_1001,N_654,N_16);
or U1002 (N_1002,N_394,N_142);
and U1003 (N_1003,N_200,N_81);
nor U1004 (N_1004,N_155,N_380);
or U1005 (N_1005,N_163,N_281);
xor U1006 (N_1006,N_125,N_183);
nand U1007 (N_1007,N_611,N_214);
and U1008 (N_1008,N_656,N_17);
nor U1009 (N_1009,N_305,N_402);
nor U1010 (N_1010,N_524,N_154);
nand U1011 (N_1011,N_548,N_56);
and U1012 (N_1012,N_663,N_20);
nand U1013 (N_1013,N_262,N_59);
xnor U1014 (N_1014,N_644,N_70);
nand U1015 (N_1015,N_213,N_195);
nor U1016 (N_1016,N_625,N_322);
or U1017 (N_1017,N_57,N_172);
nor U1018 (N_1018,N_552,N_300);
and U1019 (N_1019,N_110,N_290);
and U1020 (N_1020,N_285,N_737);
or U1021 (N_1021,N_46,N_385);
nor U1022 (N_1022,N_515,N_545);
nand U1023 (N_1023,N_479,N_169);
or U1024 (N_1024,N_196,N_468);
nand U1025 (N_1025,N_497,N_263);
nor U1026 (N_1026,N_52,N_86);
nor U1027 (N_1027,N_725,N_324);
and U1028 (N_1028,N_69,N_745);
xnor U1029 (N_1029,N_131,N_212);
or U1030 (N_1030,N_243,N_478);
nand U1031 (N_1031,N_523,N_251);
or U1032 (N_1032,N_640,N_427);
and U1033 (N_1033,N_332,N_599);
nand U1034 (N_1034,N_609,N_684);
nand U1035 (N_1035,N_676,N_458);
nand U1036 (N_1036,N_714,N_601);
nand U1037 (N_1037,N_589,N_241);
nand U1038 (N_1038,N_695,N_683);
xor U1039 (N_1039,N_340,N_739);
and U1040 (N_1040,N_116,N_386);
xor U1041 (N_1041,N_397,N_688);
xor U1042 (N_1042,N_706,N_543);
or U1043 (N_1043,N_413,N_101);
or U1044 (N_1044,N_621,N_648);
xnor U1045 (N_1045,N_405,N_64);
or U1046 (N_1046,N_519,N_352);
or U1047 (N_1047,N_129,N_30);
nand U1048 (N_1048,N_561,N_406);
and U1049 (N_1049,N_120,N_162);
nand U1050 (N_1050,N_658,N_126);
xnor U1051 (N_1051,N_502,N_687);
nor U1052 (N_1052,N_4,N_292);
and U1053 (N_1053,N_498,N_678);
xnor U1054 (N_1054,N_454,N_424);
xor U1055 (N_1055,N_261,N_598);
and U1056 (N_1056,N_622,N_132);
and U1057 (N_1057,N_620,N_418);
and U1058 (N_1058,N_247,N_541);
nand U1059 (N_1059,N_138,N_562);
and U1060 (N_1060,N_184,N_610);
and U1061 (N_1061,N_354,N_306);
or U1062 (N_1062,N_572,N_80);
xor U1063 (N_1063,N_511,N_39);
nand U1064 (N_1064,N_667,N_144);
xor U1065 (N_1065,N_655,N_740);
and U1066 (N_1066,N_192,N_661);
and U1067 (N_1067,N_659,N_414);
and U1068 (N_1068,N_299,N_113);
nor U1069 (N_1069,N_748,N_293);
nand U1070 (N_1070,N_630,N_415);
and U1071 (N_1071,N_653,N_563);
and U1072 (N_1072,N_510,N_258);
xor U1073 (N_1073,N_637,N_318);
nor U1074 (N_1074,N_276,N_366);
nor U1075 (N_1075,N_271,N_486);
nor U1076 (N_1076,N_555,N_55);
nor U1077 (N_1077,N_87,N_206);
xnor U1078 (N_1078,N_181,N_672);
xnor U1079 (N_1079,N_392,N_491);
and U1080 (N_1080,N_72,N_715);
xor U1081 (N_1081,N_137,N_236);
nor U1082 (N_1082,N_717,N_699);
xnor U1083 (N_1083,N_84,N_26);
nor U1084 (N_1084,N_558,N_141);
xnor U1085 (N_1085,N_605,N_114);
nand U1086 (N_1086,N_227,N_606);
nand U1087 (N_1087,N_417,N_377);
nor U1088 (N_1088,N_696,N_66);
nor U1089 (N_1089,N_568,N_106);
and U1090 (N_1090,N_577,N_253);
and U1091 (N_1091,N_681,N_482);
nor U1092 (N_1092,N_204,N_301);
nand U1093 (N_1093,N_512,N_48);
nor U1094 (N_1094,N_446,N_47);
nor U1095 (N_1095,N_265,N_520);
xor U1096 (N_1096,N_614,N_735);
or U1097 (N_1097,N_473,N_14);
nor U1098 (N_1098,N_689,N_239);
and U1099 (N_1099,N_375,N_105);
nor U1100 (N_1100,N_342,N_225);
or U1101 (N_1101,N_698,N_723);
nand U1102 (N_1102,N_457,N_44);
nor U1103 (N_1103,N_347,N_304);
xnor U1104 (N_1104,N_350,N_435);
nand U1105 (N_1105,N_651,N_207);
nand U1106 (N_1106,N_151,N_641);
xnor U1107 (N_1107,N_544,N_711);
nand U1108 (N_1108,N_1,N_476);
and U1109 (N_1109,N_466,N_483);
nand U1110 (N_1110,N_82,N_571);
xor U1111 (N_1111,N_348,N_34);
and U1112 (N_1112,N_311,N_382);
and U1113 (N_1113,N_13,N_303);
or U1114 (N_1114,N_528,N_330);
and U1115 (N_1115,N_569,N_602);
xnor U1116 (N_1116,N_284,N_729);
and U1117 (N_1117,N_111,N_222);
or U1118 (N_1118,N_97,N_530);
xnor U1119 (N_1119,N_534,N_346);
xor U1120 (N_1120,N_369,N_718);
nor U1121 (N_1121,N_197,N_121);
nor U1122 (N_1122,N_425,N_307);
xor U1123 (N_1123,N_187,N_401);
nand U1124 (N_1124,N_211,N_93);
or U1125 (N_1125,N_725,N_530);
or U1126 (N_1126,N_676,N_527);
xnor U1127 (N_1127,N_363,N_559);
or U1128 (N_1128,N_235,N_137);
nor U1129 (N_1129,N_539,N_738);
and U1130 (N_1130,N_59,N_510);
and U1131 (N_1131,N_92,N_113);
nand U1132 (N_1132,N_407,N_184);
nand U1133 (N_1133,N_311,N_697);
and U1134 (N_1134,N_499,N_495);
nor U1135 (N_1135,N_364,N_692);
xor U1136 (N_1136,N_445,N_47);
nand U1137 (N_1137,N_612,N_578);
or U1138 (N_1138,N_620,N_238);
or U1139 (N_1139,N_209,N_431);
and U1140 (N_1140,N_471,N_748);
nand U1141 (N_1141,N_518,N_391);
or U1142 (N_1142,N_722,N_73);
xnor U1143 (N_1143,N_651,N_476);
xor U1144 (N_1144,N_170,N_570);
or U1145 (N_1145,N_213,N_201);
and U1146 (N_1146,N_262,N_36);
nand U1147 (N_1147,N_121,N_620);
nor U1148 (N_1148,N_322,N_546);
nand U1149 (N_1149,N_117,N_407);
nor U1150 (N_1150,N_663,N_714);
nor U1151 (N_1151,N_97,N_499);
nand U1152 (N_1152,N_734,N_147);
and U1153 (N_1153,N_737,N_711);
or U1154 (N_1154,N_319,N_88);
xor U1155 (N_1155,N_571,N_253);
xor U1156 (N_1156,N_82,N_524);
xor U1157 (N_1157,N_204,N_666);
xor U1158 (N_1158,N_345,N_73);
or U1159 (N_1159,N_44,N_531);
nand U1160 (N_1160,N_669,N_422);
nand U1161 (N_1161,N_307,N_136);
xnor U1162 (N_1162,N_448,N_586);
nand U1163 (N_1163,N_179,N_285);
or U1164 (N_1164,N_90,N_276);
and U1165 (N_1165,N_188,N_211);
nor U1166 (N_1166,N_61,N_685);
or U1167 (N_1167,N_574,N_478);
and U1168 (N_1168,N_679,N_422);
and U1169 (N_1169,N_343,N_347);
xor U1170 (N_1170,N_73,N_136);
xnor U1171 (N_1171,N_619,N_333);
nor U1172 (N_1172,N_639,N_127);
nand U1173 (N_1173,N_655,N_414);
or U1174 (N_1174,N_731,N_159);
or U1175 (N_1175,N_41,N_112);
nor U1176 (N_1176,N_629,N_132);
xor U1177 (N_1177,N_480,N_64);
and U1178 (N_1178,N_501,N_97);
or U1179 (N_1179,N_173,N_340);
xor U1180 (N_1180,N_27,N_520);
nand U1181 (N_1181,N_547,N_227);
or U1182 (N_1182,N_578,N_402);
nand U1183 (N_1183,N_472,N_666);
xor U1184 (N_1184,N_107,N_587);
or U1185 (N_1185,N_294,N_549);
nor U1186 (N_1186,N_501,N_103);
and U1187 (N_1187,N_344,N_12);
or U1188 (N_1188,N_685,N_167);
nor U1189 (N_1189,N_258,N_75);
xnor U1190 (N_1190,N_102,N_374);
nand U1191 (N_1191,N_590,N_567);
nor U1192 (N_1192,N_23,N_337);
xor U1193 (N_1193,N_488,N_221);
nor U1194 (N_1194,N_625,N_348);
and U1195 (N_1195,N_63,N_311);
and U1196 (N_1196,N_254,N_422);
or U1197 (N_1197,N_89,N_537);
nand U1198 (N_1198,N_420,N_361);
xnor U1199 (N_1199,N_494,N_250);
xor U1200 (N_1200,N_14,N_342);
nor U1201 (N_1201,N_162,N_450);
xor U1202 (N_1202,N_540,N_654);
or U1203 (N_1203,N_415,N_667);
nand U1204 (N_1204,N_447,N_509);
or U1205 (N_1205,N_261,N_146);
nor U1206 (N_1206,N_665,N_332);
or U1207 (N_1207,N_375,N_137);
or U1208 (N_1208,N_17,N_605);
nand U1209 (N_1209,N_647,N_645);
and U1210 (N_1210,N_519,N_208);
nor U1211 (N_1211,N_692,N_376);
nand U1212 (N_1212,N_71,N_87);
or U1213 (N_1213,N_469,N_114);
nand U1214 (N_1214,N_368,N_100);
or U1215 (N_1215,N_436,N_627);
or U1216 (N_1216,N_177,N_234);
and U1217 (N_1217,N_43,N_502);
or U1218 (N_1218,N_367,N_344);
nor U1219 (N_1219,N_29,N_356);
xnor U1220 (N_1220,N_399,N_530);
and U1221 (N_1221,N_472,N_121);
or U1222 (N_1222,N_394,N_694);
and U1223 (N_1223,N_448,N_555);
and U1224 (N_1224,N_374,N_727);
or U1225 (N_1225,N_274,N_499);
or U1226 (N_1226,N_431,N_743);
xnor U1227 (N_1227,N_68,N_510);
nor U1228 (N_1228,N_519,N_710);
nor U1229 (N_1229,N_574,N_532);
nor U1230 (N_1230,N_38,N_429);
or U1231 (N_1231,N_505,N_639);
nor U1232 (N_1232,N_739,N_612);
nand U1233 (N_1233,N_515,N_615);
or U1234 (N_1234,N_390,N_517);
or U1235 (N_1235,N_147,N_298);
nand U1236 (N_1236,N_8,N_712);
and U1237 (N_1237,N_443,N_394);
nand U1238 (N_1238,N_439,N_30);
xor U1239 (N_1239,N_15,N_580);
or U1240 (N_1240,N_458,N_261);
nor U1241 (N_1241,N_128,N_176);
nor U1242 (N_1242,N_306,N_20);
nand U1243 (N_1243,N_429,N_193);
or U1244 (N_1244,N_51,N_343);
nor U1245 (N_1245,N_608,N_545);
xnor U1246 (N_1246,N_151,N_703);
nand U1247 (N_1247,N_671,N_728);
or U1248 (N_1248,N_743,N_423);
nor U1249 (N_1249,N_235,N_680);
nand U1250 (N_1250,N_83,N_676);
or U1251 (N_1251,N_196,N_283);
and U1252 (N_1252,N_71,N_666);
nand U1253 (N_1253,N_668,N_107);
or U1254 (N_1254,N_247,N_442);
nor U1255 (N_1255,N_285,N_588);
nor U1256 (N_1256,N_393,N_79);
nand U1257 (N_1257,N_597,N_158);
and U1258 (N_1258,N_363,N_39);
nor U1259 (N_1259,N_92,N_68);
nor U1260 (N_1260,N_316,N_306);
or U1261 (N_1261,N_662,N_643);
nor U1262 (N_1262,N_458,N_464);
and U1263 (N_1263,N_638,N_125);
xnor U1264 (N_1264,N_683,N_666);
and U1265 (N_1265,N_640,N_242);
and U1266 (N_1266,N_240,N_104);
xor U1267 (N_1267,N_646,N_312);
nand U1268 (N_1268,N_117,N_457);
nor U1269 (N_1269,N_372,N_659);
or U1270 (N_1270,N_53,N_508);
and U1271 (N_1271,N_538,N_218);
and U1272 (N_1272,N_633,N_279);
nor U1273 (N_1273,N_50,N_289);
nand U1274 (N_1274,N_184,N_521);
nor U1275 (N_1275,N_286,N_317);
xor U1276 (N_1276,N_275,N_114);
or U1277 (N_1277,N_219,N_715);
nand U1278 (N_1278,N_493,N_159);
nand U1279 (N_1279,N_687,N_150);
nor U1280 (N_1280,N_162,N_614);
and U1281 (N_1281,N_450,N_368);
or U1282 (N_1282,N_587,N_629);
nor U1283 (N_1283,N_183,N_498);
nand U1284 (N_1284,N_241,N_406);
nor U1285 (N_1285,N_124,N_418);
nand U1286 (N_1286,N_550,N_86);
xnor U1287 (N_1287,N_184,N_289);
nand U1288 (N_1288,N_269,N_233);
nor U1289 (N_1289,N_160,N_123);
and U1290 (N_1290,N_6,N_524);
xnor U1291 (N_1291,N_382,N_209);
and U1292 (N_1292,N_360,N_427);
or U1293 (N_1293,N_196,N_26);
and U1294 (N_1294,N_95,N_624);
and U1295 (N_1295,N_657,N_329);
nand U1296 (N_1296,N_658,N_155);
nor U1297 (N_1297,N_354,N_717);
or U1298 (N_1298,N_198,N_606);
nand U1299 (N_1299,N_46,N_535);
xnor U1300 (N_1300,N_362,N_698);
nand U1301 (N_1301,N_211,N_655);
nand U1302 (N_1302,N_655,N_154);
xnor U1303 (N_1303,N_336,N_447);
xor U1304 (N_1304,N_306,N_498);
nor U1305 (N_1305,N_509,N_247);
nor U1306 (N_1306,N_388,N_123);
nor U1307 (N_1307,N_661,N_157);
xor U1308 (N_1308,N_583,N_200);
nor U1309 (N_1309,N_570,N_728);
nor U1310 (N_1310,N_311,N_580);
and U1311 (N_1311,N_479,N_61);
nor U1312 (N_1312,N_175,N_490);
xor U1313 (N_1313,N_491,N_62);
and U1314 (N_1314,N_484,N_348);
xnor U1315 (N_1315,N_387,N_724);
xnor U1316 (N_1316,N_657,N_226);
nor U1317 (N_1317,N_417,N_424);
or U1318 (N_1318,N_731,N_695);
nand U1319 (N_1319,N_696,N_120);
xor U1320 (N_1320,N_392,N_339);
and U1321 (N_1321,N_647,N_693);
nor U1322 (N_1322,N_677,N_589);
xnor U1323 (N_1323,N_61,N_115);
nor U1324 (N_1324,N_115,N_22);
and U1325 (N_1325,N_169,N_310);
xnor U1326 (N_1326,N_110,N_670);
and U1327 (N_1327,N_691,N_455);
nand U1328 (N_1328,N_314,N_200);
and U1329 (N_1329,N_182,N_741);
nand U1330 (N_1330,N_519,N_456);
nand U1331 (N_1331,N_263,N_276);
nand U1332 (N_1332,N_669,N_482);
xor U1333 (N_1333,N_656,N_480);
nand U1334 (N_1334,N_412,N_334);
or U1335 (N_1335,N_94,N_699);
nand U1336 (N_1336,N_198,N_24);
and U1337 (N_1337,N_599,N_280);
nand U1338 (N_1338,N_265,N_527);
xor U1339 (N_1339,N_437,N_500);
or U1340 (N_1340,N_270,N_63);
and U1341 (N_1341,N_735,N_419);
nor U1342 (N_1342,N_145,N_32);
nor U1343 (N_1343,N_377,N_277);
nor U1344 (N_1344,N_512,N_671);
xor U1345 (N_1345,N_347,N_407);
nor U1346 (N_1346,N_337,N_261);
and U1347 (N_1347,N_100,N_309);
xor U1348 (N_1348,N_32,N_193);
nor U1349 (N_1349,N_647,N_660);
and U1350 (N_1350,N_641,N_542);
nor U1351 (N_1351,N_36,N_523);
or U1352 (N_1352,N_66,N_396);
xnor U1353 (N_1353,N_192,N_64);
xor U1354 (N_1354,N_239,N_712);
and U1355 (N_1355,N_8,N_705);
nand U1356 (N_1356,N_91,N_512);
xnor U1357 (N_1357,N_186,N_371);
or U1358 (N_1358,N_289,N_78);
xor U1359 (N_1359,N_34,N_473);
nand U1360 (N_1360,N_83,N_278);
nand U1361 (N_1361,N_664,N_691);
or U1362 (N_1362,N_43,N_695);
or U1363 (N_1363,N_117,N_338);
nand U1364 (N_1364,N_542,N_171);
nor U1365 (N_1365,N_550,N_586);
nor U1366 (N_1366,N_23,N_493);
nand U1367 (N_1367,N_587,N_529);
xor U1368 (N_1368,N_274,N_156);
or U1369 (N_1369,N_285,N_489);
and U1370 (N_1370,N_57,N_649);
and U1371 (N_1371,N_55,N_161);
xnor U1372 (N_1372,N_359,N_140);
nor U1373 (N_1373,N_285,N_110);
and U1374 (N_1374,N_620,N_566);
or U1375 (N_1375,N_143,N_725);
nor U1376 (N_1376,N_287,N_629);
nor U1377 (N_1377,N_354,N_449);
and U1378 (N_1378,N_549,N_327);
nor U1379 (N_1379,N_432,N_50);
or U1380 (N_1380,N_587,N_39);
or U1381 (N_1381,N_549,N_650);
nor U1382 (N_1382,N_726,N_626);
and U1383 (N_1383,N_661,N_695);
and U1384 (N_1384,N_325,N_673);
and U1385 (N_1385,N_255,N_501);
nor U1386 (N_1386,N_115,N_399);
nor U1387 (N_1387,N_547,N_485);
and U1388 (N_1388,N_316,N_367);
xor U1389 (N_1389,N_275,N_45);
nor U1390 (N_1390,N_628,N_579);
xnor U1391 (N_1391,N_503,N_371);
xor U1392 (N_1392,N_538,N_249);
or U1393 (N_1393,N_47,N_354);
or U1394 (N_1394,N_424,N_375);
and U1395 (N_1395,N_88,N_151);
or U1396 (N_1396,N_597,N_671);
nand U1397 (N_1397,N_638,N_484);
or U1398 (N_1398,N_235,N_449);
and U1399 (N_1399,N_645,N_626);
or U1400 (N_1400,N_182,N_657);
nor U1401 (N_1401,N_134,N_156);
nor U1402 (N_1402,N_716,N_587);
nor U1403 (N_1403,N_609,N_466);
nor U1404 (N_1404,N_377,N_168);
nor U1405 (N_1405,N_690,N_709);
and U1406 (N_1406,N_680,N_26);
nand U1407 (N_1407,N_677,N_317);
and U1408 (N_1408,N_503,N_223);
nor U1409 (N_1409,N_129,N_385);
xnor U1410 (N_1410,N_574,N_317);
nor U1411 (N_1411,N_547,N_477);
nand U1412 (N_1412,N_245,N_122);
or U1413 (N_1413,N_481,N_472);
nor U1414 (N_1414,N_244,N_5);
and U1415 (N_1415,N_424,N_730);
nor U1416 (N_1416,N_238,N_422);
nor U1417 (N_1417,N_405,N_209);
nor U1418 (N_1418,N_268,N_224);
nand U1419 (N_1419,N_714,N_620);
xor U1420 (N_1420,N_498,N_459);
xnor U1421 (N_1421,N_534,N_302);
nand U1422 (N_1422,N_641,N_405);
or U1423 (N_1423,N_690,N_643);
and U1424 (N_1424,N_74,N_674);
or U1425 (N_1425,N_134,N_470);
nand U1426 (N_1426,N_17,N_698);
and U1427 (N_1427,N_478,N_361);
nand U1428 (N_1428,N_733,N_335);
and U1429 (N_1429,N_380,N_62);
nor U1430 (N_1430,N_71,N_43);
nor U1431 (N_1431,N_6,N_577);
and U1432 (N_1432,N_529,N_191);
nand U1433 (N_1433,N_604,N_524);
nor U1434 (N_1434,N_558,N_421);
nor U1435 (N_1435,N_279,N_618);
xnor U1436 (N_1436,N_54,N_110);
or U1437 (N_1437,N_439,N_396);
and U1438 (N_1438,N_16,N_503);
or U1439 (N_1439,N_372,N_553);
or U1440 (N_1440,N_51,N_336);
xor U1441 (N_1441,N_192,N_221);
or U1442 (N_1442,N_513,N_223);
nor U1443 (N_1443,N_306,N_265);
xnor U1444 (N_1444,N_607,N_103);
or U1445 (N_1445,N_722,N_287);
or U1446 (N_1446,N_217,N_9);
nand U1447 (N_1447,N_41,N_581);
nor U1448 (N_1448,N_665,N_454);
nand U1449 (N_1449,N_661,N_207);
xnor U1450 (N_1450,N_520,N_478);
or U1451 (N_1451,N_151,N_122);
or U1452 (N_1452,N_11,N_134);
and U1453 (N_1453,N_291,N_58);
nand U1454 (N_1454,N_295,N_140);
or U1455 (N_1455,N_357,N_533);
xnor U1456 (N_1456,N_371,N_37);
xor U1457 (N_1457,N_249,N_315);
or U1458 (N_1458,N_448,N_60);
nor U1459 (N_1459,N_391,N_557);
and U1460 (N_1460,N_229,N_561);
nand U1461 (N_1461,N_475,N_421);
nand U1462 (N_1462,N_176,N_304);
and U1463 (N_1463,N_690,N_147);
nand U1464 (N_1464,N_568,N_608);
or U1465 (N_1465,N_599,N_248);
xnor U1466 (N_1466,N_729,N_615);
or U1467 (N_1467,N_144,N_726);
or U1468 (N_1468,N_463,N_172);
nor U1469 (N_1469,N_647,N_710);
and U1470 (N_1470,N_46,N_228);
nand U1471 (N_1471,N_75,N_154);
and U1472 (N_1472,N_372,N_356);
xnor U1473 (N_1473,N_438,N_143);
nor U1474 (N_1474,N_715,N_238);
xor U1475 (N_1475,N_82,N_356);
nand U1476 (N_1476,N_661,N_550);
xnor U1477 (N_1477,N_675,N_358);
xnor U1478 (N_1478,N_386,N_139);
xnor U1479 (N_1479,N_579,N_596);
nor U1480 (N_1480,N_144,N_165);
or U1481 (N_1481,N_181,N_508);
nor U1482 (N_1482,N_607,N_292);
nand U1483 (N_1483,N_728,N_287);
xor U1484 (N_1484,N_207,N_478);
nor U1485 (N_1485,N_193,N_211);
or U1486 (N_1486,N_690,N_575);
or U1487 (N_1487,N_229,N_508);
and U1488 (N_1488,N_45,N_257);
xor U1489 (N_1489,N_702,N_596);
nor U1490 (N_1490,N_395,N_115);
xnor U1491 (N_1491,N_470,N_618);
and U1492 (N_1492,N_589,N_171);
xor U1493 (N_1493,N_155,N_507);
nand U1494 (N_1494,N_349,N_172);
or U1495 (N_1495,N_666,N_562);
and U1496 (N_1496,N_80,N_727);
nor U1497 (N_1497,N_83,N_484);
nand U1498 (N_1498,N_463,N_284);
xor U1499 (N_1499,N_567,N_263);
nor U1500 (N_1500,N_1290,N_1178);
nor U1501 (N_1501,N_929,N_757);
nor U1502 (N_1502,N_915,N_1481);
nand U1503 (N_1503,N_809,N_802);
nor U1504 (N_1504,N_1026,N_1160);
xor U1505 (N_1505,N_1373,N_1497);
or U1506 (N_1506,N_759,N_926);
nand U1507 (N_1507,N_768,N_1341);
and U1508 (N_1508,N_790,N_1389);
nor U1509 (N_1509,N_777,N_1172);
and U1510 (N_1510,N_912,N_1169);
and U1511 (N_1511,N_1311,N_1372);
and U1512 (N_1512,N_1374,N_1384);
nand U1513 (N_1513,N_967,N_1415);
or U1514 (N_1514,N_928,N_839);
nor U1515 (N_1515,N_1204,N_966);
and U1516 (N_1516,N_1427,N_1316);
or U1517 (N_1517,N_1129,N_751);
nor U1518 (N_1518,N_1141,N_1445);
or U1519 (N_1519,N_917,N_881);
or U1520 (N_1520,N_978,N_843);
xor U1521 (N_1521,N_1358,N_1030);
and U1522 (N_1522,N_869,N_868);
or U1523 (N_1523,N_1032,N_805);
nor U1524 (N_1524,N_1492,N_1464);
xnor U1525 (N_1525,N_1288,N_1385);
xor U1526 (N_1526,N_950,N_1058);
or U1527 (N_1527,N_1121,N_1225);
or U1528 (N_1528,N_1371,N_810);
xnor U1529 (N_1529,N_1197,N_892);
xor U1530 (N_1530,N_1086,N_1043);
nor U1531 (N_1531,N_1240,N_1281);
and U1532 (N_1532,N_1291,N_984);
and U1533 (N_1533,N_945,N_1479);
xnor U1534 (N_1534,N_1262,N_1236);
nor U1535 (N_1535,N_1294,N_903);
or U1536 (N_1536,N_1274,N_865);
nand U1537 (N_1537,N_880,N_1229);
or U1538 (N_1538,N_1418,N_807);
xnor U1539 (N_1539,N_1231,N_1090);
and U1540 (N_1540,N_845,N_1496);
nor U1541 (N_1541,N_1054,N_1142);
or U1542 (N_1542,N_851,N_846);
and U1543 (N_1543,N_1200,N_789);
and U1544 (N_1544,N_960,N_1198);
xor U1545 (N_1545,N_1213,N_1089);
nand U1546 (N_1546,N_1016,N_1472);
xnor U1547 (N_1547,N_1303,N_764);
nor U1548 (N_1548,N_1345,N_977);
xnor U1549 (N_1549,N_1476,N_1180);
xor U1550 (N_1550,N_1220,N_1454);
and U1551 (N_1551,N_1255,N_1013);
nand U1552 (N_1552,N_1352,N_1401);
nor U1553 (N_1553,N_1143,N_987);
xor U1554 (N_1554,N_1264,N_904);
and U1555 (N_1555,N_1258,N_788);
nand U1556 (N_1556,N_762,N_1201);
xor U1557 (N_1557,N_1320,N_1446);
and U1558 (N_1558,N_925,N_933);
nor U1559 (N_1559,N_1117,N_1202);
and U1560 (N_1560,N_1430,N_1414);
or U1561 (N_1561,N_979,N_971);
or U1562 (N_1562,N_934,N_1301);
nand U1563 (N_1563,N_1495,N_1322);
and U1564 (N_1564,N_1191,N_801);
xnor U1565 (N_1565,N_1440,N_1078);
nor U1566 (N_1566,N_1069,N_1457);
xnor U1567 (N_1567,N_1152,N_857);
and U1568 (N_1568,N_1079,N_1353);
nor U1569 (N_1569,N_823,N_1287);
or U1570 (N_1570,N_808,N_1250);
nor U1571 (N_1571,N_932,N_905);
nor U1572 (N_1572,N_804,N_1488);
and U1573 (N_1573,N_957,N_1394);
nand U1574 (N_1574,N_1148,N_1273);
and U1575 (N_1575,N_961,N_1046);
and U1576 (N_1576,N_1421,N_1478);
or U1577 (N_1577,N_1383,N_1006);
nand U1578 (N_1578,N_923,N_1323);
xor U1579 (N_1579,N_1453,N_1092);
xor U1580 (N_1580,N_1138,N_1012);
and U1581 (N_1581,N_1381,N_847);
xor U1582 (N_1582,N_1252,N_1110);
and U1583 (N_1583,N_1195,N_792);
nand U1584 (N_1584,N_1115,N_1139);
or U1585 (N_1585,N_952,N_1159);
and U1586 (N_1586,N_1282,N_1116);
or U1587 (N_1587,N_958,N_1420);
or U1588 (N_1588,N_1182,N_1285);
nor U1589 (N_1589,N_1306,N_754);
xor U1590 (N_1590,N_1486,N_884);
xor U1591 (N_1591,N_794,N_913);
and U1592 (N_1592,N_756,N_986);
nand U1593 (N_1593,N_1120,N_780);
and U1594 (N_1594,N_838,N_849);
and U1595 (N_1595,N_861,N_872);
and U1596 (N_1596,N_993,N_1028);
xor U1597 (N_1597,N_1437,N_1151);
nand U1598 (N_1598,N_891,N_1087);
and U1599 (N_1599,N_1238,N_1470);
and U1600 (N_1600,N_1118,N_1408);
nand U1601 (N_1601,N_1266,N_972);
xor U1602 (N_1602,N_1442,N_949);
or U1603 (N_1603,N_862,N_1217);
nand U1604 (N_1604,N_1302,N_879);
xnor U1605 (N_1605,N_1475,N_755);
xor U1606 (N_1606,N_889,N_1035);
or U1607 (N_1607,N_1073,N_1256);
or U1608 (N_1608,N_899,N_948);
and U1609 (N_1609,N_822,N_1491);
nand U1610 (N_1610,N_1222,N_1188);
or U1611 (N_1611,N_1096,N_1104);
nand U1612 (N_1612,N_1356,N_1350);
nor U1613 (N_1613,N_1226,N_1330);
and U1614 (N_1614,N_753,N_1002);
and U1615 (N_1615,N_1490,N_1157);
and U1616 (N_1616,N_816,N_1154);
or U1617 (N_1617,N_820,N_1462);
and U1618 (N_1618,N_1349,N_1441);
or U1619 (N_1619,N_975,N_882);
and U1620 (N_1620,N_763,N_1216);
nand U1621 (N_1621,N_1275,N_1247);
nor U1622 (N_1622,N_1365,N_824);
or U1623 (N_1623,N_1362,N_1304);
and U1624 (N_1624,N_1315,N_1339);
and U1625 (N_1625,N_896,N_871);
or U1626 (N_1626,N_1125,N_1230);
nor U1627 (N_1627,N_1289,N_1091);
or U1628 (N_1628,N_1268,N_1249);
or U1629 (N_1629,N_911,N_1328);
and U1630 (N_1630,N_1337,N_1257);
and U1631 (N_1631,N_1082,N_752);
xnor U1632 (N_1632,N_797,N_1379);
or U1633 (N_1633,N_1245,N_1095);
xor U1634 (N_1634,N_936,N_1199);
nor U1635 (N_1635,N_1338,N_1380);
xnor U1636 (N_1636,N_1260,N_1327);
nand U1637 (N_1637,N_1033,N_1402);
xnor U1638 (N_1638,N_1136,N_1056);
nor U1639 (N_1639,N_907,N_776);
nand U1640 (N_1640,N_853,N_767);
nand U1641 (N_1641,N_1468,N_1270);
nand U1642 (N_1642,N_916,N_1321);
and U1643 (N_1643,N_1269,N_1443);
and U1644 (N_1644,N_841,N_795);
nand U1645 (N_1645,N_1444,N_963);
nor U1646 (N_1646,N_959,N_999);
and U1647 (N_1647,N_791,N_870);
xnor U1648 (N_1648,N_1098,N_1070);
or U1649 (N_1649,N_1359,N_894);
nor U1650 (N_1650,N_1094,N_766);
and U1651 (N_1651,N_1131,N_1449);
xor U1652 (N_1652,N_981,N_1037);
nand U1653 (N_1653,N_1439,N_1342);
and U1654 (N_1654,N_1161,N_1367);
and U1655 (N_1655,N_962,N_1041);
or U1656 (N_1656,N_842,N_1210);
and U1657 (N_1657,N_1387,N_1396);
or U1658 (N_1658,N_1061,N_990);
or U1659 (N_1659,N_1227,N_1280);
xor U1660 (N_1660,N_927,N_1029);
nand U1661 (N_1661,N_1018,N_941);
nand U1662 (N_1662,N_783,N_1326);
nand U1663 (N_1663,N_1065,N_887);
and U1664 (N_1664,N_968,N_1485);
nor U1665 (N_1665,N_989,N_897);
and U1666 (N_1666,N_1283,N_1325);
xnor U1667 (N_1667,N_1049,N_1466);
or U1668 (N_1668,N_1127,N_852);
nand U1669 (N_1669,N_1332,N_840);
or U1670 (N_1670,N_817,N_955);
nand U1671 (N_1671,N_1451,N_1426);
or U1672 (N_1672,N_1346,N_918);
nor U1673 (N_1673,N_856,N_819);
nand U1674 (N_1674,N_1417,N_1044);
nand U1675 (N_1675,N_1128,N_1234);
nand U1676 (N_1676,N_1007,N_1413);
or U1677 (N_1677,N_1461,N_1023);
nor U1678 (N_1678,N_1187,N_1045);
xnor U1679 (N_1679,N_1166,N_787);
and U1680 (N_1680,N_898,N_848);
or U1681 (N_1681,N_863,N_812);
or U1682 (N_1682,N_1331,N_938);
nor U1683 (N_1683,N_1119,N_1364);
and U1684 (N_1684,N_773,N_1314);
and U1685 (N_1685,N_1004,N_1233);
xor U1686 (N_1686,N_760,N_996);
xnor U1687 (N_1687,N_1375,N_910);
nand U1688 (N_1688,N_770,N_854);
xnor U1689 (N_1689,N_1147,N_860);
xnor U1690 (N_1690,N_1433,N_956);
and U1691 (N_1691,N_895,N_1022);
xor U1692 (N_1692,N_864,N_1034);
or U1693 (N_1693,N_1031,N_1319);
nor U1694 (N_1694,N_1378,N_1277);
and U1695 (N_1695,N_1067,N_1480);
xnor U1696 (N_1696,N_786,N_969);
nor U1697 (N_1697,N_1186,N_1419);
nor U1698 (N_1698,N_1493,N_799);
nand U1699 (N_1699,N_1053,N_1145);
and U1700 (N_1700,N_1153,N_798);
nor U1701 (N_1701,N_1298,N_976);
and U1702 (N_1702,N_1395,N_1171);
nor U1703 (N_1703,N_1436,N_1126);
nand U1704 (N_1704,N_1072,N_836);
and U1705 (N_1705,N_793,N_769);
nand U1706 (N_1706,N_1015,N_1447);
nand U1707 (N_1707,N_1101,N_1422);
or U1708 (N_1708,N_946,N_1036);
or U1709 (N_1709,N_1076,N_831);
xnor U1710 (N_1710,N_1235,N_1412);
nand U1711 (N_1711,N_1048,N_1218);
and U1712 (N_1712,N_1386,N_803);
nand U1713 (N_1713,N_821,N_1123);
and U1714 (N_1714,N_825,N_1060);
xnor U1715 (N_1715,N_1124,N_1471);
nand U1716 (N_1716,N_937,N_1363);
nand U1717 (N_1717,N_1062,N_1404);
or U1718 (N_1718,N_1391,N_1077);
or U1719 (N_1719,N_1164,N_1162);
or U1720 (N_1720,N_1390,N_1474);
and U1721 (N_1721,N_878,N_877);
and U1722 (N_1722,N_867,N_1050);
nand U1723 (N_1723,N_998,N_1361);
nor U1724 (N_1724,N_1080,N_997);
nor U1725 (N_1725,N_1360,N_1312);
or U1726 (N_1726,N_1122,N_1438);
xnor U1727 (N_1727,N_1010,N_1448);
and U1728 (N_1728,N_1196,N_1173);
or U1729 (N_1729,N_924,N_1206);
or U1730 (N_1730,N_835,N_1107);
xor U1731 (N_1731,N_992,N_951);
xor U1732 (N_1732,N_1071,N_761);
xnor U1733 (N_1733,N_1097,N_1211);
nor U1734 (N_1734,N_922,N_813);
xor U1735 (N_1735,N_1009,N_900);
nor U1736 (N_1736,N_1237,N_832);
and U1737 (N_1737,N_1271,N_1263);
or U1738 (N_1738,N_1203,N_779);
xnor U1739 (N_1739,N_908,N_874);
nor U1740 (N_1740,N_1297,N_1254);
xor U1741 (N_1741,N_1135,N_1005);
xor U1742 (N_1742,N_1344,N_1063);
nand U1743 (N_1743,N_1484,N_1168);
xnor U1744 (N_1744,N_942,N_1189);
or U1745 (N_1745,N_1112,N_1137);
nor U1746 (N_1746,N_1299,N_1134);
nand U1747 (N_1747,N_1055,N_1313);
or U1748 (N_1748,N_1400,N_909);
nand U1749 (N_1749,N_827,N_1165);
nand U1750 (N_1750,N_1042,N_1099);
nand U1751 (N_1751,N_1300,N_1088);
and U1752 (N_1752,N_1310,N_876);
xor U1753 (N_1753,N_1467,N_1146);
nor U1754 (N_1754,N_1064,N_980);
and U1755 (N_1755,N_1194,N_826);
nand U1756 (N_1756,N_1376,N_1158);
xnor U1757 (N_1757,N_1214,N_1347);
xor U1758 (N_1758,N_814,N_1163);
nor U1759 (N_1759,N_1108,N_1355);
or U1760 (N_1760,N_1431,N_830);
nand U1761 (N_1761,N_1409,N_873);
xor U1762 (N_1762,N_1228,N_1340);
xnor U1763 (N_1763,N_970,N_1111);
xor U1764 (N_1764,N_1405,N_785);
xor U1765 (N_1765,N_931,N_965);
nand U1766 (N_1766,N_800,N_1432);
or U1767 (N_1767,N_982,N_750);
and U1768 (N_1768,N_1286,N_1293);
or U1769 (N_1769,N_1174,N_901);
and U1770 (N_1770,N_834,N_890);
or U1771 (N_1771,N_1487,N_1469);
nand U1772 (N_1772,N_947,N_1190);
or U1773 (N_1773,N_1068,N_1155);
nor U1774 (N_1774,N_1223,N_1251);
and U1775 (N_1775,N_1292,N_1008);
and U1776 (N_1776,N_888,N_1179);
or U1777 (N_1777,N_930,N_1209);
or U1778 (N_1778,N_778,N_1105);
and U1779 (N_1779,N_1399,N_1185);
nand U1780 (N_1780,N_1144,N_765);
nor U1781 (N_1781,N_983,N_818);
xnor U1782 (N_1782,N_1424,N_1215);
nand U1783 (N_1783,N_1156,N_1348);
or U1784 (N_1784,N_906,N_1382);
or U1785 (N_1785,N_1435,N_1103);
xor U1786 (N_1786,N_1221,N_858);
nand U1787 (N_1787,N_893,N_1377);
or U1788 (N_1788,N_1208,N_1456);
and U1789 (N_1789,N_1140,N_1003);
nand U1790 (N_1790,N_1040,N_919);
nand U1791 (N_1791,N_1130,N_1403);
nor U1792 (N_1792,N_1425,N_1406);
xor U1793 (N_1793,N_781,N_772);
and U1794 (N_1794,N_1192,N_1177);
xnor U1795 (N_1795,N_883,N_1388);
nand U1796 (N_1796,N_1193,N_1429);
nor U1797 (N_1797,N_1494,N_1259);
nor U1798 (N_1798,N_1333,N_1265);
nor U1799 (N_1799,N_1232,N_943);
nor U1800 (N_1800,N_1000,N_1416);
nand U1801 (N_1801,N_1329,N_995);
nand U1802 (N_1802,N_1351,N_811);
or U1803 (N_1803,N_1113,N_855);
nand U1804 (N_1804,N_914,N_985);
xor U1805 (N_1805,N_1343,N_1463);
nand U1806 (N_1806,N_1392,N_1317);
and U1807 (N_1807,N_1370,N_1242);
and U1808 (N_1808,N_1025,N_796);
and U1809 (N_1809,N_1244,N_953);
or U1810 (N_1810,N_1369,N_1102);
and U1811 (N_1811,N_1020,N_1279);
nand U1812 (N_1812,N_1499,N_1465);
xor U1813 (N_1813,N_1428,N_1307);
nor U1814 (N_1814,N_1272,N_1324);
or U1815 (N_1815,N_1335,N_988);
nor U1816 (N_1816,N_1366,N_1150);
and U1817 (N_1817,N_1261,N_1167);
nand U1818 (N_1818,N_1407,N_1334);
nand U1819 (N_1819,N_1368,N_1024);
xor U1820 (N_1820,N_1219,N_1176);
nor U1821 (N_1821,N_935,N_1423);
or U1822 (N_1822,N_1085,N_1460);
nand U1823 (N_1823,N_1253,N_1066);
and U1824 (N_1824,N_1434,N_1170);
and U1825 (N_1825,N_1057,N_1458);
xnor U1826 (N_1826,N_885,N_1019);
nand U1827 (N_1827,N_1081,N_1309);
nor U1828 (N_1828,N_1038,N_1093);
nand U1829 (N_1829,N_902,N_944);
xor U1830 (N_1830,N_833,N_939);
or U1831 (N_1831,N_1278,N_1021);
nand U1832 (N_1832,N_1109,N_1411);
or U1833 (N_1833,N_1477,N_1489);
nand U1834 (N_1834,N_920,N_1083);
nand U1835 (N_1835,N_774,N_921);
xor U1836 (N_1836,N_875,N_1318);
nor U1837 (N_1837,N_1175,N_1393);
xnor U1838 (N_1838,N_1295,N_771);
and U1839 (N_1839,N_1410,N_991);
and U1840 (N_1840,N_1047,N_1241);
xor U1841 (N_1841,N_837,N_1305);
xor U1842 (N_1842,N_1308,N_1459);
or U1843 (N_1843,N_886,N_815);
and U1844 (N_1844,N_994,N_1114);
or U1845 (N_1845,N_1248,N_1052);
nand U1846 (N_1846,N_1014,N_1284);
and U1847 (N_1847,N_1473,N_1450);
nand U1848 (N_1848,N_1267,N_1452);
nand U1849 (N_1849,N_954,N_1357);
xor U1850 (N_1850,N_859,N_1074);
or U1851 (N_1851,N_866,N_1132);
xnor U1852 (N_1852,N_1084,N_829);
or U1853 (N_1853,N_1498,N_1243);
or U1854 (N_1854,N_1011,N_1106);
nor U1855 (N_1855,N_1296,N_1224);
nand U1856 (N_1856,N_758,N_1212);
or U1857 (N_1857,N_1205,N_1017);
or U1858 (N_1858,N_1246,N_1398);
or U1859 (N_1859,N_784,N_1207);
xnor U1860 (N_1860,N_775,N_1184);
nand U1861 (N_1861,N_1181,N_1039);
and U1862 (N_1862,N_1354,N_1239);
and U1863 (N_1863,N_1183,N_844);
and U1864 (N_1864,N_1001,N_1133);
and U1865 (N_1865,N_964,N_1482);
xnor U1866 (N_1866,N_806,N_1051);
xnor U1867 (N_1867,N_782,N_940);
or U1868 (N_1868,N_1027,N_828);
xnor U1869 (N_1869,N_1149,N_1276);
nor U1870 (N_1870,N_1336,N_1059);
nand U1871 (N_1871,N_1397,N_1075);
xor U1872 (N_1872,N_1100,N_1455);
nand U1873 (N_1873,N_1483,N_974);
or U1874 (N_1874,N_973,N_850);
nand U1875 (N_1875,N_796,N_1126);
nor U1876 (N_1876,N_1078,N_970);
and U1877 (N_1877,N_1243,N_1328);
xor U1878 (N_1878,N_860,N_1016);
and U1879 (N_1879,N_1317,N_799);
or U1880 (N_1880,N_1464,N_1291);
and U1881 (N_1881,N_752,N_1327);
nor U1882 (N_1882,N_1014,N_919);
or U1883 (N_1883,N_1213,N_995);
and U1884 (N_1884,N_1111,N_1352);
or U1885 (N_1885,N_1136,N_1268);
or U1886 (N_1886,N_939,N_1011);
and U1887 (N_1887,N_1382,N_1143);
nand U1888 (N_1888,N_1349,N_902);
or U1889 (N_1889,N_1004,N_1074);
or U1890 (N_1890,N_854,N_1335);
nand U1891 (N_1891,N_1379,N_1236);
or U1892 (N_1892,N_1331,N_1118);
xnor U1893 (N_1893,N_787,N_1190);
xnor U1894 (N_1894,N_1468,N_1388);
xnor U1895 (N_1895,N_1191,N_1361);
nor U1896 (N_1896,N_900,N_1332);
xor U1897 (N_1897,N_906,N_1282);
nand U1898 (N_1898,N_875,N_1236);
nor U1899 (N_1899,N_794,N_1390);
xor U1900 (N_1900,N_1201,N_950);
nor U1901 (N_1901,N_1297,N_750);
nor U1902 (N_1902,N_1112,N_1185);
nand U1903 (N_1903,N_1268,N_883);
nor U1904 (N_1904,N_1116,N_1181);
and U1905 (N_1905,N_1159,N_805);
and U1906 (N_1906,N_1434,N_1042);
nor U1907 (N_1907,N_1437,N_1363);
nor U1908 (N_1908,N_1466,N_1261);
nor U1909 (N_1909,N_941,N_891);
and U1910 (N_1910,N_889,N_1306);
nand U1911 (N_1911,N_904,N_1288);
xor U1912 (N_1912,N_1476,N_1197);
nor U1913 (N_1913,N_993,N_1227);
nor U1914 (N_1914,N_1460,N_980);
nand U1915 (N_1915,N_1078,N_1387);
or U1916 (N_1916,N_1086,N_1222);
xor U1917 (N_1917,N_1355,N_1008);
nor U1918 (N_1918,N_1347,N_1487);
xnor U1919 (N_1919,N_1175,N_1325);
and U1920 (N_1920,N_1471,N_1378);
nand U1921 (N_1921,N_1456,N_1387);
nand U1922 (N_1922,N_885,N_1320);
xor U1923 (N_1923,N_957,N_1297);
or U1924 (N_1924,N_1169,N_1495);
xnor U1925 (N_1925,N_1350,N_1251);
nand U1926 (N_1926,N_991,N_1090);
and U1927 (N_1927,N_950,N_1179);
or U1928 (N_1928,N_902,N_816);
or U1929 (N_1929,N_979,N_1438);
xnor U1930 (N_1930,N_1343,N_754);
and U1931 (N_1931,N_976,N_1498);
nand U1932 (N_1932,N_1113,N_1267);
nand U1933 (N_1933,N_1470,N_1147);
xor U1934 (N_1934,N_815,N_828);
or U1935 (N_1935,N_1028,N_1241);
xnor U1936 (N_1936,N_1360,N_1018);
nand U1937 (N_1937,N_1163,N_1486);
or U1938 (N_1938,N_795,N_1247);
and U1939 (N_1939,N_1489,N_908);
or U1940 (N_1940,N_1198,N_1291);
nand U1941 (N_1941,N_923,N_1172);
nor U1942 (N_1942,N_1042,N_1376);
xor U1943 (N_1943,N_1142,N_937);
nor U1944 (N_1944,N_820,N_1026);
nor U1945 (N_1945,N_854,N_906);
and U1946 (N_1946,N_925,N_908);
and U1947 (N_1947,N_1358,N_760);
and U1948 (N_1948,N_1207,N_1245);
nand U1949 (N_1949,N_1476,N_895);
and U1950 (N_1950,N_763,N_1085);
xor U1951 (N_1951,N_816,N_1205);
nand U1952 (N_1952,N_1061,N_1156);
or U1953 (N_1953,N_842,N_993);
and U1954 (N_1954,N_907,N_1360);
nor U1955 (N_1955,N_1222,N_786);
and U1956 (N_1956,N_1479,N_1394);
nor U1957 (N_1957,N_1042,N_821);
nor U1958 (N_1958,N_1045,N_815);
xnor U1959 (N_1959,N_993,N_1433);
nor U1960 (N_1960,N_1207,N_772);
nand U1961 (N_1961,N_1159,N_1075);
and U1962 (N_1962,N_1013,N_1069);
or U1963 (N_1963,N_1355,N_1363);
nor U1964 (N_1964,N_1112,N_1386);
and U1965 (N_1965,N_1291,N_888);
and U1966 (N_1966,N_763,N_1415);
xnor U1967 (N_1967,N_1274,N_1313);
or U1968 (N_1968,N_978,N_1086);
xnor U1969 (N_1969,N_1101,N_1385);
xor U1970 (N_1970,N_949,N_1417);
nand U1971 (N_1971,N_1036,N_1216);
nor U1972 (N_1972,N_939,N_986);
and U1973 (N_1973,N_1009,N_896);
and U1974 (N_1974,N_1490,N_1363);
and U1975 (N_1975,N_1346,N_963);
nor U1976 (N_1976,N_759,N_858);
and U1977 (N_1977,N_1280,N_1435);
xor U1978 (N_1978,N_1161,N_925);
xor U1979 (N_1979,N_842,N_1091);
nand U1980 (N_1980,N_1268,N_997);
nor U1981 (N_1981,N_1259,N_1353);
nand U1982 (N_1982,N_1367,N_1257);
or U1983 (N_1983,N_794,N_1308);
xnor U1984 (N_1984,N_1074,N_1311);
nor U1985 (N_1985,N_1292,N_1240);
nand U1986 (N_1986,N_970,N_940);
nand U1987 (N_1987,N_1271,N_1196);
nor U1988 (N_1988,N_770,N_1344);
nor U1989 (N_1989,N_852,N_1409);
or U1990 (N_1990,N_1008,N_1438);
or U1991 (N_1991,N_1247,N_1364);
nor U1992 (N_1992,N_1055,N_1019);
nor U1993 (N_1993,N_1010,N_1400);
or U1994 (N_1994,N_960,N_1149);
nor U1995 (N_1995,N_847,N_810);
and U1996 (N_1996,N_1183,N_1488);
xor U1997 (N_1997,N_987,N_1141);
or U1998 (N_1998,N_1375,N_783);
xor U1999 (N_1999,N_841,N_1391);
nand U2000 (N_2000,N_829,N_790);
or U2001 (N_2001,N_785,N_973);
xor U2002 (N_2002,N_766,N_937);
nand U2003 (N_2003,N_1399,N_1028);
nand U2004 (N_2004,N_898,N_904);
and U2005 (N_2005,N_1027,N_1076);
or U2006 (N_2006,N_1350,N_922);
nand U2007 (N_2007,N_1078,N_1290);
nor U2008 (N_2008,N_1054,N_1165);
nor U2009 (N_2009,N_1170,N_1183);
xnor U2010 (N_2010,N_1252,N_844);
nand U2011 (N_2011,N_1178,N_1149);
and U2012 (N_2012,N_1376,N_978);
nor U2013 (N_2013,N_951,N_1242);
and U2014 (N_2014,N_1105,N_848);
and U2015 (N_2015,N_791,N_1269);
nor U2016 (N_2016,N_949,N_1364);
nor U2017 (N_2017,N_957,N_1011);
nor U2018 (N_2018,N_1045,N_1088);
and U2019 (N_2019,N_945,N_877);
xnor U2020 (N_2020,N_1394,N_925);
nand U2021 (N_2021,N_857,N_869);
nand U2022 (N_2022,N_1153,N_1309);
nor U2023 (N_2023,N_1327,N_781);
xnor U2024 (N_2024,N_1245,N_950);
and U2025 (N_2025,N_1067,N_1074);
nand U2026 (N_2026,N_1222,N_1029);
xnor U2027 (N_2027,N_1254,N_947);
or U2028 (N_2028,N_919,N_1128);
nand U2029 (N_2029,N_882,N_1085);
nand U2030 (N_2030,N_1043,N_845);
nor U2031 (N_2031,N_1351,N_1290);
xor U2032 (N_2032,N_1480,N_1083);
nand U2033 (N_2033,N_1146,N_1250);
xor U2034 (N_2034,N_1309,N_829);
and U2035 (N_2035,N_1430,N_1435);
nand U2036 (N_2036,N_807,N_1103);
or U2037 (N_2037,N_847,N_908);
or U2038 (N_2038,N_1154,N_1016);
or U2039 (N_2039,N_770,N_1353);
xor U2040 (N_2040,N_1085,N_1336);
nand U2041 (N_2041,N_906,N_1041);
nor U2042 (N_2042,N_960,N_1284);
or U2043 (N_2043,N_1407,N_1142);
and U2044 (N_2044,N_1068,N_1139);
and U2045 (N_2045,N_1347,N_1346);
nand U2046 (N_2046,N_1176,N_936);
xor U2047 (N_2047,N_1190,N_974);
and U2048 (N_2048,N_1355,N_1388);
xnor U2049 (N_2049,N_1320,N_800);
xnor U2050 (N_2050,N_1365,N_1431);
nand U2051 (N_2051,N_1280,N_1066);
nand U2052 (N_2052,N_1019,N_1332);
nor U2053 (N_2053,N_894,N_1151);
nand U2054 (N_2054,N_917,N_965);
and U2055 (N_2055,N_1125,N_1225);
or U2056 (N_2056,N_761,N_966);
and U2057 (N_2057,N_1198,N_827);
nor U2058 (N_2058,N_773,N_1246);
xor U2059 (N_2059,N_965,N_1109);
and U2060 (N_2060,N_1082,N_951);
nand U2061 (N_2061,N_1008,N_1387);
nand U2062 (N_2062,N_945,N_1043);
xor U2063 (N_2063,N_1479,N_1340);
or U2064 (N_2064,N_1440,N_815);
and U2065 (N_2065,N_798,N_990);
and U2066 (N_2066,N_903,N_1333);
or U2067 (N_2067,N_1458,N_821);
xnor U2068 (N_2068,N_982,N_1024);
nor U2069 (N_2069,N_1026,N_804);
xnor U2070 (N_2070,N_1440,N_803);
nand U2071 (N_2071,N_1255,N_1389);
and U2072 (N_2072,N_1156,N_1078);
xnor U2073 (N_2073,N_1445,N_760);
or U2074 (N_2074,N_1287,N_929);
nor U2075 (N_2075,N_1280,N_1196);
and U2076 (N_2076,N_1186,N_1124);
xor U2077 (N_2077,N_836,N_1307);
nand U2078 (N_2078,N_825,N_1417);
and U2079 (N_2079,N_1446,N_1441);
xnor U2080 (N_2080,N_1289,N_902);
and U2081 (N_2081,N_1129,N_803);
nor U2082 (N_2082,N_840,N_1340);
and U2083 (N_2083,N_888,N_1129);
nor U2084 (N_2084,N_1420,N_836);
and U2085 (N_2085,N_1264,N_1148);
and U2086 (N_2086,N_1117,N_1484);
nor U2087 (N_2087,N_866,N_1028);
nor U2088 (N_2088,N_871,N_992);
xor U2089 (N_2089,N_947,N_1360);
or U2090 (N_2090,N_1131,N_1284);
nand U2091 (N_2091,N_1428,N_1226);
nor U2092 (N_2092,N_1058,N_939);
nand U2093 (N_2093,N_1416,N_987);
nand U2094 (N_2094,N_899,N_1082);
nor U2095 (N_2095,N_1094,N_1038);
nor U2096 (N_2096,N_1406,N_1191);
or U2097 (N_2097,N_827,N_1046);
xnor U2098 (N_2098,N_1293,N_1478);
or U2099 (N_2099,N_1436,N_969);
nand U2100 (N_2100,N_1430,N_894);
nand U2101 (N_2101,N_1014,N_819);
or U2102 (N_2102,N_1053,N_1434);
nand U2103 (N_2103,N_1303,N_993);
or U2104 (N_2104,N_1299,N_1359);
xnor U2105 (N_2105,N_880,N_1317);
and U2106 (N_2106,N_1048,N_1082);
nor U2107 (N_2107,N_818,N_868);
nand U2108 (N_2108,N_839,N_995);
or U2109 (N_2109,N_752,N_1268);
or U2110 (N_2110,N_953,N_1334);
nand U2111 (N_2111,N_1252,N_810);
or U2112 (N_2112,N_1287,N_1163);
or U2113 (N_2113,N_1382,N_1125);
or U2114 (N_2114,N_1388,N_807);
xor U2115 (N_2115,N_897,N_1170);
and U2116 (N_2116,N_1180,N_1446);
xor U2117 (N_2117,N_1225,N_1473);
nor U2118 (N_2118,N_873,N_1236);
nor U2119 (N_2119,N_876,N_799);
nor U2120 (N_2120,N_1197,N_1491);
and U2121 (N_2121,N_1345,N_1230);
xnor U2122 (N_2122,N_1049,N_883);
and U2123 (N_2123,N_1174,N_875);
xor U2124 (N_2124,N_942,N_885);
or U2125 (N_2125,N_1346,N_815);
nor U2126 (N_2126,N_1467,N_1220);
or U2127 (N_2127,N_829,N_1404);
or U2128 (N_2128,N_981,N_986);
nor U2129 (N_2129,N_1400,N_905);
xor U2130 (N_2130,N_1152,N_819);
or U2131 (N_2131,N_1436,N_1469);
or U2132 (N_2132,N_1001,N_1310);
nor U2133 (N_2133,N_972,N_898);
nand U2134 (N_2134,N_1466,N_1189);
xnor U2135 (N_2135,N_1301,N_1085);
nor U2136 (N_2136,N_999,N_1207);
or U2137 (N_2137,N_1199,N_1228);
nor U2138 (N_2138,N_914,N_812);
xor U2139 (N_2139,N_915,N_773);
and U2140 (N_2140,N_1110,N_1097);
nor U2141 (N_2141,N_1277,N_1440);
nand U2142 (N_2142,N_1328,N_1260);
xnor U2143 (N_2143,N_920,N_778);
and U2144 (N_2144,N_1279,N_1118);
nand U2145 (N_2145,N_1161,N_1035);
xor U2146 (N_2146,N_804,N_1098);
and U2147 (N_2147,N_930,N_1055);
or U2148 (N_2148,N_1263,N_1232);
and U2149 (N_2149,N_1340,N_817);
xor U2150 (N_2150,N_1400,N_1175);
xnor U2151 (N_2151,N_1379,N_1389);
xor U2152 (N_2152,N_955,N_1300);
xor U2153 (N_2153,N_778,N_1191);
nor U2154 (N_2154,N_832,N_1176);
xor U2155 (N_2155,N_1253,N_1086);
nor U2156 (N_2156,N_1038,N_1430);
or U2157 (N_2157,N_956,N_1243);
or U2158 (N_2158,N_1071,N_1156);
nor U2159 (N_2159,N_1003,N_1122);
xor U2160 (N_2160,N_1452,N_1475);
nor U2161 (N_2161,N_1288,N_1375);
nor U2162 (N_2162,N_1248,N_1090);
xnor U2163 (N_2163,N_1276,N_889);
xor U2164 (N_2164,N_1384,N_1033);
or U2165 (N_2165,N_1254,N_850);
xnor U2166 (N_2166,N_852,N_1429);
nand U2167 (N_2167,N_969,N_1015);
nor U2168 (N_2168,N_947,N_928);
nand U2169 (N_2169,N_1147,N_1225);
or U2170 (N_2170,N_1074,N_1347);
nand U2171 (N_2171,N_1258,N_1179);
or U2172 (N_2172,N_1015,N_1376);
or U2173 (N_2173,N_1401,N_1356);
nand U2174 (N_2174,N_1018,N_1178);
or U2175 (N_2175,N_1082,N_784);
or U2176 (N_2176,N_1318,N_1279);
or U2177 (N_2177,N_985,N_1433);
xnor U2178 (N_2178,N_1075,N_1128);
and U2179 (N_2179,N_1127,N_1000);
nor U2180 (N_2180,N_1409,N_1289);
nor U2181 (N_2181,N_1345,N_807);
nand U2182 (N_2182,N_1478,N_966);
and U2183 (N_2183,N_1422,N_1218);
nor U2184 (N_2184,N_971,N_904);
and U2185 (N_2185,N_1478,N_1180);
or U2186 (N_2186,N_1067,N_1259);
and U2187 (N_2187,N_1005,N_805);
nand U2188 (N_2188,N_1336,N_1009);
nor U2189 (N_2189,N_1280,N_1121);
nand U2190 (N_2190,N_1319,N_1169);
xnor U2191 (N_2191,N_1052,N_1476);
and U2192 (N_2192,N_870,N_1497);
xor U2193 (N_2193,N_953,N_1365);
nand U2194 (N_2194,N_1299,N_1468);
xnor U2195 (N_2195,N_1109,N_1125);
nand U2196 (N_2196,N_893,N_1255);
or U2197 (N_2197,N_1408,N_919);
xor U2198 (N_2198,N_939,N_913);
or U2199 (N_2199,N_893,N_1208);
xor U2200 (N_2200,N_878,N_1093);
or U2201 (N_2201,N_963,N_835);
or U2202 (N_2202,N_840,N_1336);
or U2203 (N_2203,N_1068,N_1015);
xor U2204 (N_2204,N_793,N_1461);
nor U2205 (N_2205,N_1151,N_1485);
and U2206 (N_2206,N_1419,N_813);
or U2207 (N_2207,N_1073,N_1341);
xnor U2208 (N_2208,N_1103,N_1151);
or U2209 (N_2209,N_993,N_899);
nor U2210 (N_2210,N_792,N_1359);
xnor U2211 (N_2211,N_1090,N_1475);
and U2212 (N_2212,N_1412,N_1003);
and U2213 (N_2213,N_1128,N_844);
and U2214 (N_2214,N_1463,N_1305);
or U2215 (N_2215,N_839,N_967);
xnor U2216 (N_2216,N_928,N_1424);
or U2217 (N_2217,N_916,N_1130);
nor U2218 (N_2218,N_934,N_1078);
nor U2219 (N_2219,N_1340,N_1269);
xnor U2220 (N_2220,N_848,N_1301);
or U2221 (N_2221,N_981,N_1021);
nand U2222 (N_2222,N_1257,N_1427);
or U2223 (N_2223,N_753,N_1427);
nand U2224 (N_2224,N_1084,N_768);
nand U2225 (N_2225,N_1344,N_942);
or U2226 (N_2226,N_1469,N_1441);
nor U2227 (N_2227,N_1178,N_1163);
nand U2228 (N_2228,N_1278,N_798);
and U2229 (N_2229,N_922,N_1484);
nand U2230 (N_2230,N_1329,N_1324);
xor U2231 (N_2231,N_906,N_1455);
and U2232 (N_2232,N_1296,N_1269);
or U2233 (N_2233,N_1444,N_1102);
nor U2234 (N_2234,N_1404,N_1052);
xnor U2235 (N_2235,N_779,N_941);
nand U2236 (N_2236,N_785,N_1158);
nand U2237 (N_2237,N_1282,N_918);
and U2238 (N_2238,N_988,N_914);
nand U2239 (N_2239,N_811,N_958);
or U2240 (N_2240,N_1071,N_1153);
nand U2241 (N_2241,N_1211,N_1049);
nor U2242 (N_2242,N_1068,N_1175);
and U2243 (N_2243,N_805,N_1141);
nand U2244 (N_2244,N_1362,N_1239);
nor U2245 (N_2245,N_1299,N_955);
nor U2246 (N_2246,N_1318,N_977);
xnor U2247 (N_2247,N_845,N_1094);
and U2248 (N_2248,N_1028,N_755);
nand U2249 (N_2249,N_1046,N_1289);
nand U2250 (N_2250,N_2076,N_1650);
nand U2251 (N_2251,N_1624,N_2058);
xnor U2252 (N_2252,N_1774,N_1952);
nand U2253 (N_2253,N_1981,N_1793);
or U2254 (N_2254,N_1810,N_1946);
nand U2255 (N_2255,N_1564,N_1849);
nand U2256 (N_2256,N_1853,N_2116);
nor U2257 (N_2257,N_1872,N_2079);
and U2258 (N_2258,N_2091,N_1530);
nor U2259 (N_2259,N_1591,N_1799);
nor U2260 (N_2260,N_2161,N_1533);
xor U2261 (N_2261,N_2033,N_1995);
nand U2262 (N_2262,N_1769,N_1549);
xnor U2263 (N_2263,N_1871,N_1722);
or U2264 (N_2264,N_1802,N_2151);
or U2265 (N_2265,N_2142,N_2128);
and U2266 (N_2266,N_1512,N_1760);
and U2267 (N_2267,N_1667,N_2111);
or U2268 (N_2268,N_1688,N_1898);
nor U2269 (N_2269,N_1526,N_2208);
and U2270 (N_2270,N_1921,N_1525);
nand U2271 (N_2271,N_2190,N_1546);
xnor U2272 (N_2272,N_2085,N_1778);
nor U2273 (N_2273,N_1666,N_1971);
nor U2274 (N_2274,N_1974,N_2083);
xor U2275 (N_2275,N_1587,N_2172);
nand U2276 (N_2276,N_2082,N_1836);
and U2277 (N_2277,N_1879,N_2201);
and U2278 (N_2278,N_2038,N_1531);
and U2279 (N_2279,N_1814,N_1585);
nor U2280 (N_2280,N_2248,N_1606);
and U2281 (N_2281,N_1963,N_2048);
or U2282 (N_2282,N_1955,N_1939);
xor U2283 (N_2283,N_1708,N_1966);
nor U2284 (N_2284,N_1729,N_2112);
xnor U2285 (N_2285,N_1867,N_1588);
xnor U2286 (N_2286,N_1837,N_1592);
nor U2287 (N_2287,N_1596,N_1862);
or U2288 (N_2288,N_1753,N_1577);
and U2289 (N_2289,N_1692,N_1684);
nand U2290 (N_2290,N_1603,N_2149);
xor U2291 (N_2291,N_1851,N_2163);
and U2292 (N_2292,N_1611,N_1870);
xnor U2293 (N_2293,N_1795,N_1701);
xor U2294 (N_2294,N_1714,N_1718);
or U2295 (N_2295,N_1831,N_1846);
nand U2296 (N_2296,N_1682,N_2146);
nand U2297 (N_2297,N_1741,N_1863);
nor U2298 (N_2298,N_1675,N_2185);
or U2299 (N_2299,N_2003,N_2053);
and U2300 (N_2300,N_1510,N_1731);
and U2301 (N_2301,N_1744,N_1809);
or U2302 (N_2302,N_1518,N_2102);
and U2303 (N_2303,N_1940,N_1792);
or U2304 (N_2304,N_1516,N_1706);
or U2305 (N_2305,N_1768,N_2013);
nand U2306 (N_2306,N_2122,N_2051);
xor U2307 (N_2307,N_1913,N_1960);
xor U2308 (N_2308,N_1922,N_2064);
nor U2309 (N_2309,N_1780,N_1626);
nand U2310 (N_2310,N_1545,N_1888);
nor U2311 (N_2311,N_2200,N_2097);
nand U2312 (N_2312,N_1647,N_1557);
nor U2313 (N_2313,N_1961,N_1779);
and U2314 (N_2314,N_1926,N_1983);
nor U2315 (N_2315,N_2216,N_1556);
or U2316 (N_2316,N_2054,N_2007);
and U2317 (N_2317,N_1878,N_1555);
xor U2318 (N_2318,N_1899,N_1785);
nand U2319 (N_2319,N_1916,N_1674);
or U2320 (N_2320,N_1565,N_1664);
nor U2321 (N_2321,N_2059,N_1751);
nor U2322 (N_2322,N_1991,N_2095);
and U2323 (N_2323,N_1873,N_1844);
xnor U2324 (N_2324,N_1571,N_1665);
or U2325 (N_2325,N_1835,N_1820);
nor U2326 (N_2326,N_1761,N_1796);
and U2327 (N_2327,N_2158,N_1987);
nor U2328 (N_2328,N_1568,N_2042);
or U2329 (N_2329,N_2093,N_2075);
nor U2330 (N_2330,N_2171,N_1906);
nand U2331 (N_2331,N_1947,N_1797);
xnor U2332 (N_2332,N_2067,N_2119);
xor U2333 (N_2333,N_2100,N_1941);
nand U2334 (N_2334,N_2150,N_1747);
nand U2335 (N_2335,N_1515,N_1874);
and U2336 (N_2336,N_1736,N_2098);
nor U2337 (N_2337,N_2104,N_1543);
nand U2338 (N_2338,N_2004,N_1724);
or U2339 (N_2339,N_1663,N_1788);
and U2340 (N_2340,N_1629,N_1639);
and U2341 (N_2341,N_1806,N_1601);
nor U2342 (N_2342,N_1958,N_1959);
nand U2343 (N_2343,N_1553,N_1640);
and U2344 (N_2344,N_1819,N_1656);
and U2345 (N_2345,N_1746,N_2164);
and U2346 (N_2346,N_2065,N_2213);
or U2347 (N_2347,N_2162,N_1977);
xor U2348 (N_2348,N_1965,N_1576);
and U2349 (N_2349,N_2189,N_2219);
nand U2350 (N_2350,N_1877,N_1956);
nor U2351 (N_2351,N_1670,N_1843);
or U2352 (N_2352,N_1693,N_2245);
or U2353 (N_2353,N_1679,N_1969);
xor U2354 (N_2354,N_2140,N_1506);
and U2355 (N_2355,N_2180,N_1570);
xnor U2356 (N_2356,N_1643,N_1550);
nor U2357 (N_2357,N_2237,N_2176);
and U2358 (N_2358,N_2022,N_2160);
nor U2359 (N_2359,N_1756,N_2125);
or U2360 (N_2360,N_1999,N_1602);
or U2361 (N_2361,N_2030,N_2069);
and U2362 (N_2362,N_2139,N_1794);
and U2363 (N_2363,N_1558,N_2019);
nand U2364 (N_2364,N_1676,N_1535);
nor U2365 (N_2365,N_1786,N_1772);
xor U2366 (N_2366,N_2221,N_2192);
nand U2367 (N_2367,N_2061,N_1979);
xnor U2368 (N_2368,N_1850,N_2239);
xnor U2369 (N_2369,N_1798,N_1860);
nor U2370 (N_2370,N_1962,N_1604);
or U2371 (N_2371,N_1903,N_1929);
and U2372 (N_2372,N_1887,N_1749);
and U2373 (N_2373,N_1928,N_2089);
xnor U2374 (N_2374,N_2209,N_2127);
nand U2375 (N_2375,N_2035,N_2047);
nand U2376 (N_2376,N_2143,N_1694);
or U2377 (N_2377,N_2238,N_1509);
nor U2378 (N_2378,N_1856,N_1996);
xor U2379 (N_2379,N_1644,N_1598);
nand U2380 (N_2380,N_2233,N_2194);
xor U2381 (N_2381,N_1990,N_2105);
and U2382 (N_2382,N_1582,N_1934);
and U2383 (N_2383,N_1909,N_1513);
nor U2384 (N_2384,N_2010,N_1919);
and U2385 (N_2385,N_1847,N_1538);
and U2386 (N_2386,N_2141,N_1935);
or U2387 (N_2387,N_1813,N_1583);
nor U2388 (N_2388,N_1998,N_2231);
xor U2389 (N_2389,N_1918,N_2080);
and U2390 (N_2390,N_1700,N_2060);
or U2391 (N_2391,N_1646,N_2009);
or U2392 (N_2392,N_1561,N_2099);
nor U2393 (N_2393,N_1619,N_1889);
nand U2394 (N_2394,N_2152,N_2134);
nand U2395 (N_2395,N_2199,N_1876);
nor U2396 (N_2396,N_1567,N_1677);
and U2397 (N_2397,N_2036,N_1933);
nor U2398 (N_2398,N_2206,N_1719);
or U2399 (N_2399,N_1901,N_2191);
nand U2400 (N_2400,N_2230,N_1704);
and U2401 (N_2401,N_1637,N_1953);
nor U2402 (N_2402,N_2137,N_2074);
and U2403 (N_2403,N_1972,N_2197);
and U2404 (N_2404,N_2016,N_2148);
nor U2405 (N_2405,N_1709,N_1711);
and U2406 (N_2406,N_1816,N_1655);
and U2407 (N_2407,N_1978,N_2052);
nor U2408 (N_2408,N_2008,N_1771);
xor U2409 (N_2409,N_1949,N_1770);
nor U2410 (N_2410,N_1743,N_1707);
and U2411 (N_2411,N_2057,N_1528);
or U2412 (N_2412,N_2202,N_1757);
xnor U2413 (N_2413,N_1520,N_1652);
nand U2414 (N_2414,N_1766,N_2113);
nor U2415 (N_2415,N_2120,N_1623);
nand U2416 (N_2416,N_1855,N_1593);
or U2417 (N_2417,N_2168,N_1866);
and U2418 (N_2418,N_2068,N_1580);
nand U2419 (N_2419,N_1748,N_1578);
nand U2420 (N_2420,N_2027,N_1735);
nand U2421 (N_2421,N_2050,N_2228);
xnor U2422 (N_2422,N_1628,N_1575);
or U2423 (N_2423,N_2002,N_2039);
nand U2424 (N_2424,N_1517,N_2012);
nand U2425 (N_2425,N_1875,N_2108);
xnor U2426 (N_2426,N_1800,N_1521);
and U2427 (N_2427,N_1739,N_1861);
nor U2428 (N_2428,N_1884,N_1833);
or U2429 (N_2429,N_1503,N_2032);
nor U2430 (N_2430,N_2026,N_1857);
and U2431 (N_2431,N_1698,N_2044);
and U2432 (N_2432,N_2196,N_2001);
nand U2433 (N_2433,N_1572,N_1631);
nand U2434 (N_2434,N_1653,N_1609);
or U2435 (N_2435,N_1508,N_2103);
nor U2436 (N_2436,N_1830,N_1989);
and U2437 (N_2437,N_2155,N_1671);
or U2438 (N_2438,N_1566,N_1697);
nor U2439 (N_2439,N_2118,N_1865);
and U2440 (N_2440,N_1573,N_2045);
nand U2441 (N_2441,N_2123,N_1773);
xnor U2442 (N_2442,N_2218,N_2188);
nand U2443 (N_2443,N_1973,N_1529);
xnor U2444 (N_2444,N_1937,N_1801);
nor U2445 (N_2445,N_1712,N_2145);
nor U2446 (N_2446,N_1811,N_1829);
or U2447 (N_2447,N_1662,N_1752);
xnor U2448 (N_2448,N_1992,N_2204);
xnor U2449 (N_2449,N_1762,N_2167);
xnor U2450 (N_2450,N_1777,N_1661);
nor U2451 (N_2451,N_2070,N_2138);
nand U2452 (N_2452,N_1548,N_2130);
nand U2453 (N_2453,N_1594,N_2198);
xor U2454 (N_2454,N_2225,N_1902);
and U2455 (N_2455,N_1673,N_1791);
and U2456 (N_2456,N_1840,N_1890);
and U2457 (N_2457,N_2017,N_2159);
nor U2458 (N_2458,N_2014,N_1911);
xor U2459 (N_2459,N_1822,N_2041);
nor U2460 (N_2460,N_1938,N_1915);
or U2461 (N_2461,N_2087,N_2242);
xnor U2462 (N_2462,N_1783,N_1642);
and U2463 (N_2463,N_1554,N_2217);
nor U2464 (N_2464,N_1621,N_1635);
nand U2465 (N_2465,N_1616,N_2210);
and U2466 (N_2466,N_2124,N_1534);
nor U2467 (N_2467,N_2028,N_1514);
nand U2468 (N_2468,N_1563,N_1982);
nand U2469 (N_2469,N_1808,N_1597);
nand U2470 (N_2470,N_1608,N_2110);
nand U2471 (N_2471,N_1931,N_1805);
nor U2472 (N_2472,N_1910,N_1511);
xnor U2473 (N_2473,N_1532,N_2147);
xor U2474 (N_2474,N_2055,N_1854);
and U2475 (N_2475,N_1713,N_2072);
nand U2476 (N_2476,N_1569,N_2165);
and U2477 (N_2477,N_1574,N_2182);
nand U2478 (N_2478,N_1895,N_2144);
nor U2479 (N_2479,N_1765,N_1638);
xnor U2480 (N_2480,N_1614,N_1925);
nor U2481 (N_2481,N_2115,N_2183);
or U2482 (N_2482,N_1505,N_1993);
nor U2483 (N_2483,N_1680,N_2203);
nand U2484 (N_2484,N_1845,N_2181);
and U2485 (N_2485,N_2227,N_2094);
or U2486 (N_2486,N_1552,N_1970);
xnor U2487 (N_2487,N_1522,N_2157);
nor U2488 (N_2488,N_2056,N_1834);
or U2489 (N_2489,N_1636,N_1590);
or U2490 (N_2490,N_1527,N_2226);
and U2491 (N_2491,N_1904,N_1559);
or U2492 (N_2492,N_1524,N_2177);
or U2493 (N_2493,N_1660,N_1579);
nor U2494 (N_2494,N_2133,N_1787);
or U2495 (N_2495,N_2235,N_2066);
or U2496 (N_2496,N_2187,N_1767);
nand U2497 (N_2497,N_1702,N_1723);
and U2498 (N_2498,N_1657,N_2049);
xnor U2499 (N_2499,N_2234,N_1562);
and U2500 (N_2500,N_1672,N_1584);
and U2501 (N_2501,N_1804,N_1838);
or U2502 (N_2502,N_1897,N_1886);
xnor U2503 (N_2503,N_1907,N_1618);
xor U2504 (N_2504,N_2121,N_1504);
xnor U2505 (N_2505,N_1868,N_2131);
nand U2506 (N_2506,N_1980,N_1669);
and U2507 (N_2507,N_1852,N_2246);
nand U2508 (N_2508,N_2015,N_2090);
nand U2509 (N_2509,N_1730,N_1790);
xnor U2510 (N_2510,N_2166,N_1900);
nand U2511 (N_2511,N_2247,N_1542);
xnor U2512 (N_2512,N_2106,N_2153);
xnor U2513 (N_2513,N_1612,N_1658);
or U2514 (N_2514,N_1882,N_2109);
nor U2515 (N_2515,N_1763,N_1968);
and U2516 (N_2516,N_1745,N_1826);
xnor U2517 (N_2517,N_1781,N_1930);
or U2518 (N_2518,N_2078,N_1893);
and U2519 (N_2519,N_1633,N_1710);
xnor U2520 (N_2520,N_1738,N_1825);
or U2521 (N_2521,N_2062,N_2046);
nor U2522 (N_2522,N_1881,N_1627);
xnor U2523 (N_2523,N_2249,N_2214);
and U2524 (N_2524,N_1950,N_1696);
or U2525 (N_2525,N_1817,N_2136);
nand U2526 (N_2526,N_1776,N_2086);
nand U2527 (N_2527,N_1645,N_1914);
nor U2528 (N_2528,N_1595,N_1892);
nor U2529 (N_2529,N_1678,N_1848);
nand U2530 (N_2530,N_2174,N_1858);
xor U2531 (N_2531,N_1964,N_2034);
xor U2532 (N_2532,N_1905,N_1832);
or U2533 (N_2533,N_1734,N_2195);
xnor U2534 (N_2534,N_2173,N_1944);
and U2535 (N_2535,N_2229,N_1932);
and U2536 (N_2536,N_1648,N_1641);
nand U2537 (N_2537,N_1540,N_1758);
nor U2538 (N_2538,N_2241,N_2005);
nor U2539 (N_2539,N_1803,N_2175);
nor U2540 (N_2540,N_1782,N_1740);
nand U2541 (N_2541,N_1581,N_1685);
or U2542 (N_2542,N_2244,N_1859);
xnor U2543 (N_2543,N_1519,N_1622);
nor U2544 (N_2544,N_2169,N_1755);
or U2545 (N_2545,N_1589,N_1997);
nor U2546 (N_2546,N_1703,N_2040);
nor U2547 (N_2547,N_1732,N_1537);
nor U2548 (N_2548,N_2063,N_2071);
nor U2549 (N_2549,N_1927,N_1942);
or U2550 (N_2550,N_1764,N_2232);
xnor U2551 (N_2551,N_1617,N_2211);
and U2552 (N_2552,N_1824,N_1507);
and U2553 (N_2553,N_2215,N_1668);
nor U2554 (N_2554,N_1541,N_2031);
or U2555 (N_2555,N_1721,N_2212);
and U2556 (N_2556,N_1632,N_2184);
or U2557 (N_2557,N_2205,N_1924);
xnor U2558 (N_2558,N_1985,N_2156);
nor U2559 (N_2559,N_1691,N_1737);
and U2560 (N_2560,N_2193,N_1705);
nand U2561 (N_2561,N_2170,N_2077);
or U2562 (N_2562,N_1954,N_1894);
xor U2563 (N_2563,N_1500,N_1984);
nand U2564 (N_2564,N_1716,N_1994);
nand U2565 (N_2565,N_1759,N_2025);
or U2566 (N_2566,N_2224,N_2207);
nand U2567 (N_2567,N_2043,N_1539);
and U2568 (N_2568,N_1726,N_1864);
or U2569 (N_2569,N_2243,N_2006);
xor U2570 (N_2570,N_1908,N_1630);
and U2571 (N_2571,N_1742,N_2021);
or U2572 (N_2572,N_1986,N_1920);
or U2573 (N_2573,N_1586,N_2129);
and U2574 (N_2574,N_1689,N_1536);
nand U2575 (N_2575,N_1615,N_1605);
or U2576 (N_2576,N_2037,N_1883);
or U2577 (N_2577,N_2114,N_2081);
or U2578 (N_2578,N_1815,N_1789);
nor U2579 (N_2579,N_1625,N_1839);
and U2580 (N_2580,N_1613,N_1501);
or U2581 (N_2581,N_1727,N_2220);
nor U2582 (N_2582,N_1891,N_1975);
or U2583 (N_2583,N_1560,N_1957);
and U2584 (N_2584,N_1649,N_1917);
or U2585 (N_2585,N_2084,N_2179);
nand U2586 (N_2586,N_1715,N_1943);
and U2587 (N_2587,N_1885,N_2092);
xor U2588 (N_2588,N_2107,N_1923);
nor U2589 (N_2589,N_2178,N_1607);
nor U2590 (N_2590,N_2101,N_2088);
and U2591 (N_2591,N_2011,N_2186);
or U2592 (N_2592,N_1720,N_1717);
nand U2593 (N_2593,N_1733,N_1775);
and U2594 (N_2594,N_2132,N_1620);
and U2595 (N_2595,N_2236,N_1690);
xor U2596 (N_2596,N_1823,N_1821);
or U2597 (N_2597,N_1599,N_2073);
nor U2598 (N_2598,N_1725,N_1610);
xnor U2599 (N_2599,N_2135,N_1551);
or U2600 (N_2600,N_1828,N_1686);
or U2601 (N_2601,N_2154,N_1896);
xnor U2602 (N_2602,N_1754,N_1681);
nand U2603 (N_2603,N_1976,N_1842);
nand U2604 (N_2604,N_1699,N_2096);
nand U2605 (N_2605,N_1728,N_2126);
nor U2606 (N_2606,N_1967,N_2117);
or U2607 (N_2607,N_1687,N_1880);
or U2608 (N_2608,N_1544,N_1750);
nor U2609 (N_2609,N_2018,N_1651);
xnor U2610 (N_2610,N_1936,N_2024);
nand U2611 (N_2611,N_1600,N_1841);
nor U2612 (N_2612,N_2023,N_1988);
or U2613 (N_2613,N_1654,N_1547);
xnor U2614 (N_2614,N_1695,N_1807);
nor U2615 (N_2615,N_2240,N_1951);
or U2616 (N_2616,N_1827,N_2029);
nand U2617 (N_2617,N_2000,N_1523);
and U2618 (N_2618,N_1659,N_1948);
or U2619 (N_2619,N_1784,N_2223);
or U2620 (N_2620,N_1812,N_1818);
nand U2621 (N_2621,N_2222,N_1502);
nand U2622 (N_2622,N_1634,N_1683);
and U2623 (N_2623,N_1869,N_2020);
nor U2624 (N_2624,N_1912,N_1945);
nand U2625 (N_2625,N_1831,N_2108);
and U2626 (N_2626,N_1820,N_2167);
or U2627 (N_2627,N_1905,N_1860);
and U2628 (N_2628,N_1506,N_1646);
xnor U2629 (N_2629,N_1901,N_1600);
nor U2630 (N_2630,N_1823,N_2045);
and U2631 (N_2631,N_1692,N_1568);
and U2632 (N_2632,N_1954,N_2182);
and U2633 (N_2633,N_2118,N_1908);
and U2634 (N_2634,N_1625,N_1833);
xnor U2635 (N_2635,N_1842,N_1847);
nand U2636 (N_2636,N_1847,N_2204);
or U2637 (N_2637,N_1651,N_1642);
xor U2638 (N_2638,N_1793,N_1751);
or U2639 (N_2639,N_2045,N_1811);
and U2640 (N_2640,N_2049,N_1763);
or U2641 (N_2641,N_1643,N_1895);
nor U2642 (N_2642,N_1789,N_1930);
or U2643 (N_2643,N_1867,N_1831);
nor U2644 (N_2644,N_2025,N_2237);
and U2645 (N_2645,N_2146,N_1940);
nand U2646 (N_2646,N_1811,N_1650);
nor U2647 (N_2647,N_2228,N_1523);
xor U2648 (N_2648,N_1674,N_2110);
xor U2649 (N_2649,N_1944,N_2104);
nor U2650 (N_2650,N_1553,N_1509);
nand U2651 (N_2651,N_1814,N_1765);
and U2652 (N_2652,N_1835,N_2207);
nand U2653 (N_2653,N_2119,N_1577);
xnor U2654 (N_2654,N_1699,N_1879);
nand U2655 (N_2655,N_2051,N_2114);
xnor U2656 (N_2656,N_2205,N_2233);
nand U2657 (N_2657,N_1540,N_1768);
xnor U2658 (N_2658,N_2066,N_2227);
nor U2659 (N_2659,N_1571,N_1982);
or U2660 (N_2660,N_1971,N_2221);
and U2661 (N_2661,N_2222,N_2216);
xor U2662 (N_2662,N_2063,N_2166);
nor U2663 (N_2663,N_1696,N_2210);
nor U2664 (N_2664,N_2089,N_1689);
nand U2665 (N_2665,N_2188,N_2087);
nand U2666 (N_2666,N_1764,N_1894);
and U2667 (N_2667,N_1886,N_1856);
or U2668 (N_2668,N_1697,N_1910);
or U2669 (N_2669,N_1837,N_1724);
nand U2670 (N_2670,N_1860,N_2131);
or U2671 (N_2671,N_2103,N_2017);
and U2672 (N_2672,N_1765,N_1622);
nor U2673 (N_2673,N_1628,N_2072);
xor U2674 (N_2674,N_1836,N_2108);
nor U2675 (N_2675,N_1591,N_2244);
nor U2676 (N_2676,N_2075,N_1553);
nand U2677 (N_2677,N_2122,N_1754);
or U2678 (N_2678,N_1859,N_1616);
nor U2679 (N_2679,N_2083,N_2207);
xor U2680 (N_2680,N_2101,N_2230);
xnor U2681 (N_2681,N_2146,N_1628);
nand U2682 (N_2682,N_2008,N_1554);
xnor U2683 (N_2683,N_2112,N_2204);
nor U2684 (N_2684,N_1759,N_2022);
xor U2685 (N_2685,N_2088,N_1687);
or U2686 (N_2686,N_1937,N_2123);
or U2687 (N_2687,N_1602,N_1622);
and U2688 (N_2688,N_1512,N_1878);
xor U2689 (N_2689,N_1930,N_2170);
nand U2690 (N_2690,N_1961,N_1630);
or U2691 (N_2691,N_2240,N_1588);
and U2692 (N_2692,N_1815,N_1787);
nor U2693 (N_2693,N_1732,N_2236);
or U2694 (N_2694,N_1855,N_2058);
and U2695 (N_2695,N_1559,N_1510);
xnor U2696 (N_2696,N_1732,N_1750);
xnor U2697 (N_2697,N_2082,N_1658);
or U2698 (N_2698,N_1809,N_1575);
xor U2699 (N_2699,N_1963,N_2123);
nand U2700 (N_2700,N_1837,N_1554);
nand U2701 (N_2701,N_1536,N_2054);
and U2702 (N_2702,N_1675,N_1540);
nand U2703 (N_2703,N_1795,N_2242);
xor U2704 (N_2704,N_1518,N_1602);
nand U2705 (N_2705,N_1628,N_1860);
or U2706 (N_2706,N_1916,N_1540);
xnor U2707 (N_2707,N_1677,N_1650);
nor U2708 (N_2708,N_1554,N_1562);
or U2709 (N_2709,N_1646,N_2108);
and U2710 (N_2710,N_2055,N_2192);
nand U2711 (N_2711,N_2144,N_1516);
nor U2712 (N_2712,N_1610,N_1707);
nand U2713 (N_2713,N_1643,N_1844);
and U2714 (N_2714,N_2214,N_1796);
or U2715 (N_2715,N_2174,N_1828);
and U2716 (N_2716,N_1892,N_1666);
xor U2717 (N_2717,N_2014,N_1879);
and U2718 (N_2718,N_2087,N_2123);
xnor U2719 (N_2719,N_1870,N_1751);
nand U2720 (N_2720,N_2168,N_1693);
nor U2721 (N_2721,N_1610,N_2145);
or U2722 (N_2722,N_1942,N_2226);
nor U2723 (N_2723,N_2227,N_2078);
nor U2724 (N_2724,N_1937,N_2214);
nand U2725 (N_2725,N_1983,N_1891);
nand U2726 (N_2726,N_1906,N_2213);
nand U2727 (N_2727,N_1827,N_1676);
and U2728 (N_2728,N_1839,N_1852);
nand U2729 (N_2729,N_1617,N_1791);
or U2730 (N_2730,N_1648,N_1677);
xnor U2731 (N_2731,N_1637,N_2025);
nor U2732 (N_2732,N_1955,N_2045);
nor U2733 (N_2733,N_1754,N_2097);
or U2734 (N_2734,N_1608,N_2154);
nor U2735 (N_2735,N_1705,N_2065);
nor U2736 (N_2736,N_2205,N_1868);
and U2737 (N_2737,N_1813,N_1745);
nand U2738 (N_2738,N_1629,N_1830);
xor U2739 (N_2739,N_2070,N_1717);
nand U2740 (N_2740,N_1605,N_1856);
or U2741 (N_2741,N_2186,N_1817);
nor U2742 (N_2742,N_1801,N_1840);
xnor U2743 (N_2743,N_1831,N_2140);
xor U2744 (N_2744,N_1588,N_2095);
xnor U2745 (N_2745,N_1669,N_1672);
or U2746 (N_2746,N_1625,N_1945);
and U2747 (N_2747,N_1923,N_1628);
and U2748 (N_2748,N_1679,N_1716);
nand U2749 (N_2749,N_1997,N_1641);
nand U2750 (N_2750,N_2050,N_1653);
or U2751 (N_2751,N_1928,N_1745);
or U2752 (N_2752,N_2060,N_1988);
or U2753 (N_2753,N_1616,N_1806);
xor U2754 (N_2754,N_2158,N_2089);
nand U2755 (N_2755,N_1681,N_1805);
nor U2756 (N_2756,N_1698,N_2123);
or U2757 (N_2757,N_1763,N_2030);
nand U2758 (N_2758,N_1596,N_2208);
xor U2759 (N_2759,N_1716,N_1558);
and U2760 (N_2760,N_1784,N_1984);
nand U2761 (N_2761,N_1964,N_2246);
nor U2762 (N_2762,N_2099,N_1857);
nand U2763 (N_2763,N_1682,N_2056);
nor U2764 (N_2764,N_1983,N_1583);
nor U2765 (N_2765,N_1760,N_1942);
and U2766 (N_2766,N_1830,N_2188);
nand U2767 (N_2767,N_1561,N_1907);
xor U2768 (N_2768,N_1638,N_1779);
xor U2769 (N_2769,N_2071,N_1705);
xnor U2770 (N_2770,N_2059,N_1988);
and U2771 (N_2771,N_2173,N_1704);
nand U2772 (N_2772,N_1723,N_2040);
nor U2773 (N_2773,N_2224,N_2010);
xor U2774 (N_2774,N_2099,N_2087);
nor U2775 (N_2775,N_1914,N_1660);
xor U2776 (N_2776,N_1987,N_1684);
nand U2777 (N_2777,N_1594,N_1993);
nor U2778 (N_2778,N_1655,N_2083);
nor U2779 (N_2779,N_1522,N_2028);
nand U2780 (N_2780,N_2188,N_2079);
xor U2781 (N_2781,N_1729,N_1773);
nand U2782 (N_2782,N_1929,N_1700);
xnor U2783 (N_2783,N_2210,N_1531);
or U2784 (N_2784,N_2031,N_2112);
nand U2785 (N_2785,N_1915,N_1742);
xnor U2786 (N_2786,N_1566,N_1955);
nand U2787 (N_2787,N_1833,N_1871);
xnor U2788 (N_2788,N_1754,N_1901);
and U2789 (N_2789,N_1837,N_2189);
or U2790 (N_2790,N_1809,N_2098);
nor U2791 (N_2791,N_1833,N_2178);
or U2792 (N_2792,N_1675,N_2071);
or U2793 (N_2793,N_1795,N_1504);
nor U2794 (N_2794,N_1523,N_2240);
or U2795 (N_2795,N_2160,N_2175);
xor U2796 (N_2796,N_1765,N_1780);
nor U2797 (N_2797,N_2123,N_1545);
and U2798 (N_2798,N_2102,N_1567);
and U2799 (N_2799,N_2015,N_2246);
nor U2800 (N_2800,N_1870,N_1614);
xnor U2801 (N_2801,N_1659,N_2029);
or U2802 (N_2802,N_1999,N_2157);
and U2803 (N_2803,N_2213,N_1615);
or U2804 (N_2804,N_1854,N_1658);
nor U2805 (N_2805,N_1662,N_2221);
xor U2806 (N_2806,N_1522,N_2060);
and U2807 (N_2807,N_2047,N_2177);
nor U2808 (N_2808,N_2142,N_1580);
or U2809 (N_2809,N_2195,N_1708);
and U2810 (N_2810,N_1688,N_1617);
nand U2811 (N_2811,N_1517,N_2188);
or U2812 (N_2812,N_1886,N_1740);
nor U2813 (N_2813,N_1904,N_1517);
nor U2814 (N_2814,N_2207,N_1972);
or U2815 (N_2815,N_2112,N_2136);
or U2816 (N_2816,N_1717,N_2199);
nor U2817 (N_2817,N_2022,N_1966);
nand U2818 (N_2818,N_1836,N_1681);
or U2819 (N_2819,N_1500,N_1935);
or U2820 (N_2820,N_2139,N_2036);
nand U2821 (N_2821,N_2244,N_1775);
or U2822 (N_2822,N_1555,N_2055);
and U2823 (N_2823,N_1778,N_2125);
and U2824 (N_2824,N_1510,N_1607);
xor U2825 (N_2825,N_1870,N_1837);
xor U2826 (N_2826,N_2096,N_1771);
or U2827 (N_2827,N_2104,N_1691);
xnor U2828 (N_2828,N_1705,N_2222);
nand U2829 (N_2829,N_1702,N_1920);
or U2830 (N_2830,N_1920,N_1530);
nand U2831 (N_2831,N_1861,N_2192);
nor U2832 (N_2832,N_2046,N_2175);
xnor U2833 (N_2833,N_1507,N_1775);
xnor U2834 (N_2834,N_1942,N_2048);
and U2835 (N_2835,N_1722,N_1901);
nor U2836 (N_2836,N_1718,N_1818);
or U2837 (N_2837,N_1840,N_2061);
xor U2838 (N_2838,N_1567,N_1837);
xnor U2839 (N_2839,N_1975,N_1565);
xor U2840 (N_2840,N_1990,N_1779);
nor U2841 (N_2841,N_2052,N_1988);
and U2842 (N_2842,N_1998,N_2113);
and U2843 (N_2843,N_2097,N_1572);
xnor U2844 (N_2844,N_1971,N_1931);
nand U2845 (N_2845,N_2168,N_1772);
and U2846 (N_2846,N_1625,N_1867);
xor U2847 (N_2847,N_1924,N_1955);
nand U2848 (N_2848,N_1770,N_2129);
nor U2849 (N_2849,N_1731,N_1865);
and U2850 (N_2850,N_2038,N_1649);
xor U2851 (N_2851,N_1954,N_1560);
nand U2852 (N_2852,N_2116,N_2018);
or U2853 (N_2853,N_1880,N_1910);
and U2854 (N_2854,N_1595,N_1519);
and U2855 (N_2855,N_1738,N_1667);
nand U2856 (N_2856,N_1550,N_1933);
nor U2857 (N_2857,N_1542,N_1556);
and U2858 (N_2858,N_1736,N_2142);
and U2859 (N_2859,N_2011,N_1850);
xnor U2860 (N_2860,N_2142,N_1537);
xnor U2861 (N_2861,N_1534,N_1999);
nor U2862 (N_2862,N_2151,N_1721);
xnor U2863 (N_2863,N_1762,N_2077);
nand U2864 (N_2864,N_2070,N_1912);
xnor U2865 (N_2865,N_1832,N_2149);
nor U2866 (N_2866,N_1679,N_1683);
xnor U2867 (N_2867,N_2146,N_2179);
xor U2868 (N_2868,N_2018,N_1546);
xor U2869 (N_2869,N_2104,N_2244);
xor U2870 (N_2870,N_1930,N_1806);
and U2871 (N_2871,N_1864,N_1951);
nand U2872 (N_2872,N_1778,N_2090);
or U2873 (N_2873,N_1735,N_2061);
nand U2874 (N_2874,N_1845,N_1642);
and U2875 (N_2875,N_1876,N_2112);
and U2876 (N_2876,N_1934,N_1640);
nor U2877 (N_2877,N_1678,N_1856);
or U2878 (N_2878,N_1536,N_2167);
xor U2879 (N_2879,N_1697,N_1572);
and U2880 (N_2880,N_1603,N_2111);
and U2881 (N_2881,N_1604,N_2100);
or U2882 (N_2882,N_1612,N_1946);
nand U2883 (N_2883,N_1827,N_2248);
and U2884 (N_2884,N_2219,N_1975);
xnor U2885 (N_2885,N_2066,N_1855);
xor U2886 (N_2886,N_2134,N_1509);
and U2887 (N_2887,N_1905,N_1805);
and U2888 (N_2888,N_2068,N_2089);
nand U2889 (N_2889,N_2064,N_2118);
or U2890 (N_2890,N_2048,N_1801);
nor U2891 (N_2891,N_2169,N_2057);
or U2892 (N_2892,N_1822,N_1862);
xor U2893 (N_2893,N_1735,N_1585);
nor U2894 (N_2894,N_2070,N_2120);
nand U2895 (N_2895,N_1989,N_1913);
and U2896 (N_2896,N_1817,N_1588);
nand U2897 (N_2897,N_1904,N_2019);
or U2898 (N_2898,N_1974,N_1758);
or U2899 (N_2899,N_2178,N_1581);
nand U2900 (N_2900,N_1903,N_2144);
nor U2901 (N_2901,N_2096,N_2144);
nor U2902 (N_2902,N_1817,N_2126);
nor U2903 (N_2903,N_2128,N_1903);
nand U2904 (N_2904,N_1834,N_2071);
and U2905 (N_2905,N_1605,N_1553);
or U2906 (N_2906,N_1992,N_1621);
or U2907 (N_2907,N_1884,N_2000);
xnor U2908 (N_2908,N_1705,N_2066);
nor U2909 (N_2909,N_2026,N_2035);
or U2910 (N_2910,N_1819,N_1594);
nand U2911 (N_2911,N_2248,N_1577);
or U2912 (N_2912,N_1758,N_2019);
and U2913 (N_2913,N_2118,N_2167);
and U2914 (N_2914,N_2122,N_2049);
nor U2915 (N_2915,N_1716,N_1906);
xor U2916 (N_2916,N_1996,N_1730);
xnor U2917 (N_2917,N_1881,N_1707);
xor U2918 (N_2918,N_2031,N_1711);
nor U2919 (N_2919,N_1669,N_1640);
xor U2920 (N_2920,N_1702,N_1587);
nor U2921 (N_2921,N_1590,N_1686);
nand U2922 (N_2922,N_2060,N_1521);
nor U2923 (N_2923,N_1561,N_1655);
xnor U2924 (N_2924,N_1771,N_2225);
xor U2925 (N_2925,N_2241,N_2169);
nand U2926 (N_2926,N_2238,N_1584);
nand U2927 (N_2927,N_1961,N_2071);
or U2928 (N_2928,N_2133,N_1543);
or U2929 (N_2929,N_2220,N_2227);
xnor U2930 (N_2930,N_1940,N_2049);
or U2931 (N_2931,N_1538,N_2155);
nor U2932 (N_2932,N_2044,N_2085);
or U2933 (N_2933,N_2165,N_1689);
nor U2934 (N_2934,N_2174,N_2002);
and U2935 (N_2935,N_1723,N_1649);
nand U2936 (N_2936,N_1576,N_1749);
nor U2937 (N_2937,N_1656,N_1861);
xor U2938 (N_2938,N_1819,N_1846);
nand U2939 (N_2939,N_2214,N_1966);
or U2940 (N_2940,N_1940,N_1522);
or U2941 (N_2941,N_1988,N_1647);
nor U2942 (N_2942,N_1947,N_1574);
or U2943 (N_2943,N_2247,N_1759);
or U2944 (N_2944,N_2191,N_2128);
and U2945 (N_2945,N_2221,N_1557);
and U2946 (N_2946,N_2155,N_1563);
nand U2947 (N_2947,N_1722,N_1541);
and U2948 (N_2948,N_1836,N_2243);
and U2949 (N_2949,N_1966,N_2242);
and U2950 (N_2950,N_2073,N_2198);
xor U2951 (N_2951,N_1500,N_2161);
xnor U2952 (N_2952,N_2120,N_1685);
or U2953 (N_2953,N_1639,N_2231);
nand U2954 (N_2954,N_1975,N_1985);
or U2955 (N_2955,N_2173,N_1749);
nor U2956 (N_2956,N_1937,N_1916);
nor U2957 (N_2957,N_1773,N_2218);
or U2958 (N_2958,N_2248,N_1869);
nand U2959 (N_2959,N_1735,N_1921);
nand U2960 (N_2960,N_2055,N_2153);
nand U2961 (N_2961,N_1752,N_1824);
nor U2962 (N_2962,N_1952,N_1556);
nand U2963 (N_2963,N_1674,N_1624);
and U2964 (N_2964,N_2079,N_1698);
nand U2965 (N_2965,N_1930,N_1892);
nand U2966 (N_2966,N_2058,N_2153);
or U2967 (N_2967,N_2073,N_2010);
or U2968 (N_2968,N_2214,N_2177);
and U2969 (N_2969,N_2125,N_2058);
nor U2970 (N_2970,N_1661,N_2208);
nor U2971 (N_2971,N_1517,N_1847);
nor U2972 (N_2972,N_2161,N_1819);
nor U2973 (N_2973,N_1711,N_1978);
and U2974 (N_2974,N_1881,N_1703);
nor U2975 (N_2975,N_1972,N_1967);
xnor U2976 (N_2976,N_2222,N_1583);
or U2977 (N_2977,N_1910,N_1973);
nand U2978 (N_2978,N_1577,N_2186);
and U2979 (N_2979,N_1619,N_1672);
and U2980 (N_2980,N_1657,N_2102);
and U2981 (N_2981,N_1831,N_2221);
or U2982 (N_2982,N_1761,N_1936);
xnor U2983 (N_2983,N_1919,N_1973);
or U2984 (N_2984,N_1641,N_2126);
nand U2985 (N_2985,N_1695,N_1956);
and U2986 (N_2986,N_1592,N_1502);
nand U2987 (N_2987,N_1865,N_1853);
or U2988 (N_2988,N_1956,N_2013);
nor U2989 (N_2989,N_1745,N_1792);
and U2990 (N_2990,N_1746,N_1822);
xor U2991 (N_2991,N_1511,N_2115);
xor U2992 (N_2992,N_2064,N_1714);
nand U2993 (N_2993,N_1951,N_1703);
nand U2994 (N_2994,N_2120,N_2060);
xnor U2995 (N_2995,N_1997,N_1504);
and U2996 (N_2996,N_1839,N_1546);
xor U2997 (N_2997,N_1900,N_1831);
nor U2998 (N_2998,N_1599,N_1809);
and U2999 (N_2999,N_1917,N_1694);
xor UO_0 (O_0,N_2259,N_2331);
xor UO_1 (O_1,N_2535,N_2948);
nand UO_2 (O_2,N_2341,N_2662);
nand UO_3 (O_3,N_2916,N_2870);
or UO_4 (O_4,N_2792,N_2348);
xnor UO_5 (O_5,N_2598,N_2364);
xnor UO_6 (O_6,N_2761,N_2497);
or UO_7 (O_7,N_2506,N_2635);
xnor UO_8 (O_8,N_2597,N_2834);
xor UO_9 (O_9,N_2596,N_2633);
or UO_10 (O_10,N_2504,N_2265);
or UO_11 (O_11,N_2936,N_2647);
xor UO_12 (O_12,N_2789,N_2886);
or UO_13 (O_13,N_2583,N_2460);
and UO_14 (O_14,N_2723,N_2977);
nand UO_15 (O_15,N_2577,N_2283);
nor UO_16 (O_16,N_2405,N_2315);
and UO_17 (O_17,N_2841,N_2314);
or UO_18 (O_18,N_2437,N_2652);
nor UO_19 (O_19,N_2940,N_2755);
nor UO_20 (O_20,N_2260,N_2367);
xnor UO_21 (O_21,N_2725,N_2857);
or UO_22 (O_22,N_2706,N_2892);
nand UO_23 (O_23,N_2880,N_2564);
nand UO_24 (O_24,N_2756,N_2396);
xnor UO_25 (O_25,N_2584,N_2909);
nand UO_26 (O_26,N_2398,N_2743);
and UO_27 (O_27,N_2994,N_2316);
nand UO_28 (O_28,N_2608,N_2907);
xnor UO_29 (O_29,N_2650,N_2842);
or UO_30 (O_30,N_2619,N_2956);
nand UO_31 (O_31,N_2753,N_2860);
and UO_32 (O_32,N_2530,N_2809);
or UO_33 (O_33,N_2879,N_2567);
nor UO_34 (O_34,N_2592,N_2637);
nor UO_35 (O_35,N_2589,N_2313);
or UO_36 (O_36,N_2551,N_2812);
nand UO_37 (O_37,N_2252,N_2636);
nor UO_38 (O_38,N_2421,N_2914);
nand UO_39 (O_39,N_2988,N_2675);
nor UO_40 (O_40,N_2747,N_2441);
nand UO_41 (O_41,N_2394,N_2849);
or UO_42 (O_42,N_2918,N_2453);
and UO_43 (O_43,N_2431,N_2721);
nand UO_44 (O_44,N_2972,N_2778);
nand UO_45 (O_45,N_2447,N_2470);
or UO_46 (O_46,N_2526,N_2872);
and UO_47 (O_47,N_2974,N_2534);
xor UO_48 (O_48,N_2978,N_2830);
xor UO_49 (O_49,N_2660,N_2281);
and UO_50 (O_50,N_2933,N_2762);
and UO_51 (O_51,N_2754,N_2997);
and UO_52 (O_52,N_2739,N_2986);
and UO_53 (O_53,N_2544,N_2646);
nand UO_54 (O_54,N_2590,N_2305);
and UO_55 (O_55,N_2649,N_2628);
or UO_56 (O_56,N_2268,N_2850);
or UO_57 (O_57,N_2278,N_2802);
xnor UO_58 (O_58,N_2772,N_2665);
xnor UO_59 (O_59,N_2319,N_2429);
and UO_60 (O_60,N_2851,N_2536);
and UO_61 (O_61,N_2345,N_2670);
nor UO_62 (O_62,N_2552,N_2444);
or UO_63 (O_63,N_2381,N_2286);
nand UO_64 (O_64,N_2903,N_2528);
and UO_65 (O_65,N_2449,N_2611);
and UO_66 (O_66,N_2482,N_2338);
nor UO_67 (O_67,N_2365,N_2712);
nand UO_68 (O_68,N_2794,N_2703);
and UO_69 (O_69,N_2784,N_2507);
or UO_70 (O_70,N_2919,N_2737);
nor UO_71 (O_71,N_2443,N_2539);
and UO_72 (O_72,N_2959,N_2266);
nand UO_73 (O_73,N_2912,N_2563);
xor UO_74 (O_74,N_2688,N_2687);
xnor UO_75 (O_75,N_2780,N_2658);
and UO_76 (O_76,N_2831,N_2284);
nand UO_77 (O_77,N_2478,N_2663);
and UO_78 (O_78,N_2622,N_2485);
xor UO_79 (O_79,N_2942,N_2648);
xor UO_80 (O_80,N_2454,N_2632);
and UO_81 (O_81,N_2964,N_2764);
nand UO_82 (O_82,N_2736,N_2751);
and UO_83 (O_83,N_2492,N_2407);
nand UO_84 (O_84,N_2791,N_2807);
nand UO_85 (O_85,N_2932,N_2783);
and UO_86 (O_86,N_2822,N_2966);
nand UO_87 (O_87,N_2895,N_2640);
nand UO_88 (O_88,N_2771,N_2846);
and UO_89 (O_89,N_2533,N_2351);
nor UO_90 (O_90,N_2624,N_2818);
nand UO_91 (O_91,N_2490,N_2343);
nand UO_92 (O_92,N_2484,N_2430);
nand UO_93 (O_93,N_2885,N_2613);
nand UO_94 (O_94,N_2621,N_2397);
nor UO_95 (O_95,N_2576,N_2825);
nand UO_96 (O_96,N_2935,N_2913);
nand UO_97 (O_97,N_2678,N_2815);
nor UO_98 (O_98,N_2340,N_2385);
and UO_99 (O_99,N_2273,N_2603);
and UO_100 (O_100,N_2927,N_2710);
nand UO_101 (O_101,N_2973,N_2990);
or UO_102 (O_102,N_2776,N_2604);
nand UO_103 (O_103,N_2414,N_2373);
and UO_104 (O_104,N_2760,N_2420);
or UO_105 (O_105,N_2828,N_2954);
xor UO_106 (O_106,N_2573,N_2735);
and UO_107 (O_107,N_2814,N_2399);
and UO_108 (O_108,N_2602,N_2882);
xor UO_109 (O_109,N_2806,N_2446);
or UO_110 (O_110,N_2740,N_2963);
and UO_111 (O_111,N_2730,N_2386);
xnor UO_112 (O_112,N_2984,N_2354);
and UO_113 (O_113,N_2661,N_2701);
and UO_114 (O_114,N_2749,N_2931);
or UO_115 (O_115,N_2889,N_2525);
xnor UO_116 (O_116,N_2861,N_2821);
or UO_117 (O_117,N_2673,N_2685);
nand UO_118 (O_118,N_2450,N_2411);
xnor UO_119 (O_119,N_2768,N_2378);
nand UO_120 (O_120,N_2826,N_2541);
or UO_121 (O_121,N_2989,N_2323);
xnor UO_122 (O_122,N_2500,N_2915);
nor UO_123 (O_123,N_2334,N_2926);
nand UO_124 (O_124,N_2804,N_2677);
nand UO_125 (O_125,N_2837,N_2819);
xor UO_126 (O_126,N_2312,N_2298);
xor UO_127 (O_127,N_2516,N_2352);
or UO_128 (O_128,N_2930,N_2587);
nor UO_129 (O_129,N_2529,N_2473);
and UO_130 (O_130,N_2422,N_2554);
or UO_131 (O_131,N_2594,N_2499);
xnor UO_132 (O_132,N_2545,N_2466);
or UO_133 (O_133,N_2409,N_2339);
and UO_134 (O_134,N_2494,N_2958);
nor UO_135 (O_135,N_2741,N_2356);
nor UO_136 (O_136,N_2433,N_2408);
nor UO_137 (O_137,N_2653,N_2700);
xor UO_138 (O_138,N_2540,N_2944);
and UO_139 (O_139,N_2871,N_2757);
or UO_140 (O_140,N_2616,N_2342);
and UO_141 (O_141,N_2777,N_2642);
nor UO_142 (O_142,N_2669,N_2383);
nand UO_143 (O_143,N_2403,N_2404);
and UO_144 (O_144,N_2998,N_2838);
nand UO_145 (O_145,N_2332,N_2401);
or UO_146 (O_146,N_2855,N_2766);
xnor UO_147 (O_147,N_2579,N_2750);
and UO_148 (O_148,N_2434,N_2863);
nand UO_149 (O_149,N_2271,N_2439);
nor UO_150 (O_150,N_2881,N_2412);
xnor UO_151 (O_151,N_2392,N_2575);
xor UO_152 (O_152,N_2538,N_2615);
nand UO_153 (O_153,N_2694,N_2377);
nand UO_154 (O_154,N_2867,N_2620);
and UO_155 (O_155,N_2558,N_2543);
or UO_156 (O_156,N_2793,N_2276);
nor UO_157 (O_157,N_2417,N_2774);
or UO_158 (O_158,N_2285,N_2690);
xnor UO_159 (O_159,N_2329,N_2897);
or UO_160 (O_160,N_2371,N_2258);
xor UO_161 (O_161,N_2854,N_2318);
nand UO_162 (O_162,N_2264,N_2537);
or UO_163 (O_163,N_2501,N_2522);
xnor UO_164 (O_164,N_2709,N_2696);
xnor UO_165 (O_165,N_2455,N_2512);
and UO_166 (O_166,N_2303,N_2742);
or UO_167 (O_167,N_2843,N_2614);
nor UO_168 (O_168,N_2436,N_2428);
and UO_169 (O_169,N_2302,N_2968);
xnor UO_170 (O_170,N_2350,N_2362);
and UO_171 (O_171,N_2718,N_2773);
xor UO_172 (O_172,N_2574,N_2983);
or UO_173 (O_173,N_2910,N_2560);
xor UO_174 (O_174,N_2686,N_2487);
and UO_175 (O_175,N_2711,N_2297);
or UO_176 (O_176,N_2874,N_2659);
or UO_177 (O_177,N_2427,N_2758);
nand UO_178 (O_178,N_2257,N_2581);
and UO_179 (O_179,N_2811,N_2901);
xor UO_180 (O_180,N_2275,N_2508);
and UO_181 (O_181,N_2705,N_2287);
or UO_182 (O_182,N_2625,N_2906);
or UO_183 (O_183,N_2905,N_2423);
nand UO_184 (O_184,N_2566,N_2631);
and UO_185 (O_185,N_2941,N_2971);
nor UO_186 (O_186,N_2985,N_2698);
xnor UO_187 (O_187,N_2513,N_2790);
or UO_188 (O_188,N_2402,N_2309);
nand UO_189 (O_189,N_2839,N_2668);
or UO_190 (O_190,N_2785,N_2716);
nor UO_191 (O_191,N_2600,N_2481);
nand UO_192 (O_192,N_2713,N_2496);
and UO_193 (O_193,N_2335,N_2992);
and UO_194 (O_194,N_2645,N_2468);
nand UO_195 (O_195,N_2923,N_2883);
or UO_196 (O_196,N_2813,N_2588);
xor UO_197 (O_197,N_2488,N_2559);
and UO_198 (O_198,N_2426,N_2925);
or UO_199 (O_199,N_2267,N_2389);
nor UO_200 (O_200,N_2719,N_2456);
nand UO_201 (O_201,N_2462,N_2418);
xor UO_202 (O_202,N_2320,N_2578);
xor UO_203 (O_203,N_2279,N_2734);
or UO_204 (O_204,N_2786,N_2961);
xnor UO_205 (O_205,N_2435,N_2483);
and UO_206 (O_206,N_2571,N_2432);
xor UO_207 (O_207,N_2502,N_2726);
or UO_208 (O_208,N_2795,N_2556);
nor UO_209 (O_209,N_2480,N_2752);
nor UO_210 (O_210,N_2656,N_2952);
nand UO_211 (O_211,N_2946,N_2651);
or UO_212 (O_212,N_2689,N_2363);
or UO_213 (O_213,N_2550,N_2442);
nor UO_214 (O_214,N_2250,N_2410);
and UO_215 (O_215,N_2474,N_2347);
xor UO_216 (O_216,N_2947,N_2708);
xnor UO_217 (O_217,N_2519,N_2894);
nor UO_218 (O_218,N_2609,N_2937);
or UO_219 (O_219,N_2585,N_2326);
nand UO_220 (O_220,N_2951,N_2344);
xor UO_221 (O_221,N_2962,N_2748);
and UO_222 (O_222,N_2369,N_2333);
nor UO_223 (O_223,N_2699,N_2955);
nor UO_224 (O_224,N_2294,N_2469);
nand UO_225 (O_225,N_2505,N_2511);
and UO_226 (O_226,N_2251,N_2461);
and UO_227 (O_227,N_2835,N_2666);
nand UO_228 (O_228,N_2531,N_2920);
xor UO_229 (O_229,N_2565,N_2898);
nor UO_230 (O_230,N_2452,N_2738);
nand UO_231 (O_231,N_2641,N_2293);
or UO_232 (O_232,N_2532,N_2727);
nor UO_233 (O_233,N_2805,N_2865);
xor UO_234 (O_234,N_2569,N_2729);
or UO_235 (O_235,N_2272,N_2262);
or UO_236 (O_236,N_2400,N_2981);
nor UO_237 (O_237,N_2891,N_2606);
xnor UO_238 (O_238,N_2707,N_2489);
nor UO_239 (O_239,N_2680,N_2800);
xor UO_240 (O_240,N_2714,N_2382);
and UO_241 (O_241,N_2254,N_2953);
nor UO_242 (O_242,N_2840,N_2495);
and UO_243 (O_243,N_2349,N_2355);
xor UO_244 (O_244,N_2803,N_2384);
nor UO_245 (O_245,N_2987,N_2358);
or UO_246 (O_246,N_2939,N_2928);
nor UO_247 (O_247,N_2817,N_2884);
nor UO_248 (O_248,N_2899,N_2848);
or UO_249 (O_249,N_2976,N_2965);
or UO_250 (O_250,N_2921,N_2859);
nor UO_251 (O_251,N_2852,N_2368);
nand UO_252 (O_252,N_2390,N_2671);
nor UO_253 (O_253,N_2869,N_2887);
or UO_254 (O_254,N_2862,N_2996);
nand UO_255 (O_255,N_2844,N_2463);
or UO_256 (O_256,N_2995,N_2722);
or UO_257 (O_257,N_2498,N_2610);
and UO_258 (O_258,N_2683,N_2324);
or UO_259 (O_259,N_2810,N_2982);
nor UO_260 (O_260,N_2547,N_2280);
nor UO_261 (O_261,N_2292,N_2361);
and UO_262 (O_262,N_2509,N_2877);
nand UO_263 (O_263,N_2634,N_2679);
xor UO_264 (O_264,N_2797,N_2731);
xor UO_265 (O_265,N_2289,N_2304);
or UO_266 (O_266,N_2704,N_2288);
and UO_267 (O_267,N_2514,N_2801);
xor UO_268 (O_268,N_2424,N_2299);
and UO_269 (O_269,N_2527,N_2425);
nand UO_270 (O_270,N_2263,N_2975);
xor UO_271 (O_271,N_2391,N_2582);
or UO_272 (O_272,N_2518,N_2759);
xnor UO_273 (O_273,N_2943,N_2676);
nand UO_274 (O_274,N_2360,N_2465);
xnor UO_275 (O_275,N_2546,N_2770);
or UO_276 (O_276,N_2542,N_2684);
xor UO_277 (O_277,N_2639,N_2562);
or UO_278 (O_278,N_2440,N_2599);
or UO_279 (O_279,N_2779,N_2568);
or UO_280 (O_280,N_2993,N_2799);
xor UO_281 (O_281,N_2732,N_2827);
nor UO_282 (O_282,N_2864,N_2503);
nor UO_283 (O_283,N_2969,N_2457);
or UO_284 (O_284,N_2655,N_2824);
or UO_285 (O_285,N_2798,N_2379);
or UO_286 (O_286,N_2702,N_2823);
nand UO_287 (O_287,N_2256,N_2717);
or UO_288 (O_288,N_2957,N_2617);
nor UO_289 (O_289,N_2471,N_2682);
nor UO_290 (O_290,N_2847,N_2787);
xor UO_291 (O_291,N_2380,N_2724);
nand UO_292 (O_292,N_2261,N_2376);
or UO_293 (O_293,N_2691,N_2464);
and UO_294 (O_294,N_2630,N_2307);
nor UO_295 (O_295,N_2322,N_2458);
nand UO_296 (O_296,N_2715,N_2856);
xor UO_297 (O_297,N_2832,N_2908);
nand UO_298 (O_298,N_2548,N_2664);
or UO_299 (O_299,N_2623,N_2853);
nand UO_300 (O_300,N_2336,N_2595);
or UO_301 (O_301,N_2359,N_2366);
and UO_302 (O_302,N_2517,N_2306);
nor UO_303 (O_303,N_2999,N_2255);
xor UO_304 (O_304,N_2561,N_2667);
and UO_305 (O_305,N_2605,N_2745);
and UO_306 (O_306,N_2521,N_2681);
or UO_307 (O_307,N_2419,N_2555);
xnor UO_308 (O_308,N_2720,N_2310);
nand UO_309 (O_309,N_2782,N_2438);
nor UO_310 (O_310,N_2896,N_2788);
and UO_311 (O_311,N_2393,N_2644);
xor UO_312 (O_312,N_2922,N_2970);
nand UO_313 (O_313,N_2878,N_2627);
or UO_314 (O_314,N_2416,N_2820);
or UO_315 (O_315,N_2586,N_2866);
nor UO_316 (O_316,N_2744,N_2672);
xor UO_317 (O_317,N_2888,N_2949);
or UO_318 (O_318,N_2321,N_2697);
nor UO_319 (O_319,N_2290,N_2991);
xor UO_320 (O_320,N_2570,N_2733);
xnor UO_321 (O_321,N_2638,N_2626);
and UO_322 (O_322,N_2911,N_2467);
or UO_323 (O_323,N_2893,N_2524);
nor UO_324 (O_324,N_2728,N_2346);
nand UO_325 (O_325,N_2451,N_2924);
nor UO_326 (O_326,N_2295,N_2308);
and UO_327 (O_327,N_2960,N_2693);
or UO_328 (O_328,N_2375,N_2612);
nand UO_329 (O_329,N_2291,N_2591);
xnor UO_330 (O_330,N_2479,N_2775);
and UO_331 (O_331,N_2767,N_2607);
nand UO_332 (O_332,N_2282,N_2328);
nor UO_333 (O_333,N_2520,N_2868);
xor UO_334 (O_334,N_2269,N_2808);
or UO_335 (O_335,N_2388,N_2938);
and UO_336 (O_336,N_2395,N_2274);
xor UO_337 (O_337,N_2674,N_2934);
nand UO_338 (O_338,N_2557,N_2876);
nand UO_339 (O_339,N_2781,N_2657);
nor UO_340 (O_340,N_2459,N_2327);
or UO_341 (O_341,N_2337,N_2270);
nand UO_342 (O_342,N_2406,N_2572);
or UO_343 (O_343,N_2593,N_2510);
or UO_344 (O_344,N_2580,N_2765);
nand UO_345 (O_345,N_2387,N_2374);
nand UO_346 (O_346,N_2300,N_2372);
nor UO_347 (O_347,N_2301,N_2904);
nand UO_348 (O_348,N_2253,N_2763);
and UO_349 (O_349,N_2601,N_2448);
xnor UO_350 (O_350,N_2929,N_2875);
and UO_351 (O_351,N_2415,N_2353);
nor UO_352 (O_352,N_2477,N_2796);
and UO_353 (O_353,N_2950,N_2979);
or UO_354 (O_354,N_2816,N_2523);
nand UO_355 (O_355,N_2917,N_2845);
xor UO_356 (O_356,N_2486,N_2858);
xor UO_357 (O_357,N_2654,N_2829);
xnor UO_358 (O_358,N_2873,N_2695);
or UO_359 (O_359,N_2553,N_2900);
xor UO_360 (O_360,N_2618,N_2475);
xnor UO_361 (O_361,N_2330,N_2515);
nor UO_362 (O_362,N_2833,N_2357);
xor UO_363 (O_363,N_2445,N_2472);
nor UO_364 (O_364,N_2413,N_2277);
or UO_365 (O_365,N_2890,N_2945);
xor UO_366 (O_366,N_2967,N_2549);
nor UO_367 (O_367,N_2836,N_2980);
nor UO_368 (O_368,N_2325,N_2643);
and UO_369 (O_369,N_2629,N_2491);
nor UO_370 (O_370,N_2692,N_2493);
nor UO_371 (O_371,N_2370,N_2476);
or UO_372 (O_372,N_2311,N_2317);
and UO_373 (O_373,N_2769,N_2296);
xnor UO_374 (O_374,N_2746,N_2902);
xor UO_375 (O_375,N_2369,N_2811);
xnor UO_376 (O_376,N_2932,N_2717);
or UO_377 (O_377,N_2940,N_2952);
or UO_378 (O_378,N_2524,N_2747);
or UO_379 (O_379,N_2274,N_2328);
nor UO_380 (O_380,N_2874,N_2944);
nor UO_381 (O_381,N_2448,N_2387);
nand UO_382 (O_382,N_2367,N_2823);
nand UO_383 (O_383,N_2678,N_2493);
or UO_384 (O_384,N_2787,N_2724);
nand UO_385 (O_385,N_2971,N_2718);
nor UO_386 (O_386,N_2482,N_2973);
and UO_387 (O_387,N_2804,N_2624);
nand UO_388 (O_388,N_2320,N_2647);
and UO_389 (O_389,N_2435,N_2992);
nand UO_390 (O_390,N_2280,N_2982);
nand UO_391 (O_391,N_2348,N_2529);
or UO_392 (O_392,N_2959,N_2769);
xor UO_393 (O_393,N_2987,N_2483);
or UO_394 (O_394,N_2400,N_2620);
or UO_395 (O_395,N_2328,N_2497);
or UO_396 (O_396,N_2898,N_2968);
nor UO_397 (O_397,N_2574,N_2343);
and UO_398 (O_398,N_2350,N_2794);
xnor UO_399 (O_399,N_2683,N_2511);
and UO_400 (O_400,N_2648,N_2769);
nand UO_401 (O_401,N_2741,N_2436);
nand UO_402 (O_402,N_2777,N_2608);
nand UO_403 (O_403,N_2571,N_2840);
xnor UO_404 (O_404,N_2843,N_2579);
nand UO_405 (O_405,N_2909,N_2452);
nand UO_406 (O_406,N_2897,N_2769);
nand UO_407 (O_407,N_2802,N_2940);
and UO_408 (O_408,N_2348,N_2257);
xnor UO_409 (O_409,N_2486,N_2646);
or UO_410 (O_410,N_2320,N_2430);
or UO_411 (O_411,N_2606,N_2292);
nor UO_412 (O_412,N_2641,N_2580);
and UO_413 (O_413,N_2937,N_2780);
and UO_414 (O_414,N_2784,N_2577);
xor UO_415 (O_415,N_2339,N_2470);
nor UO_416 (O_416,N_2797,N_2307);
nor UO_417 (O_417,N_2469,N_2907);
nor UO_418 (O_418,N_2680,N_2913);
or UO_419 (O_419,N_2479,N_2854);
or UO_420 (O_420,N_2955,N_2717);
or UO_421 (O_421,N_2561,N_2814);
nand UO_422 (O_422,N_2559,N_2526);
or UO_423 (O_423,N_2586,N_2322);
xnor UO_424 (O_424,N_2689,N_2383);
and UO_425 (O_425,N_2703,N_2690);
and UO_426 (O_426,N_2278,N_2585);
and UO_427 (O_427,N_2484,N_2929);
and UO_428 (O_428,N_2804,N_2987);
nor UO_429 (O_429,N_2379,N_2481);
nor UO_430 (O_430,N_2373,N_2509);
nor UO_431 (O_431,N_2609,N_2808);
nand UO_432 (O_432,N_2421,N_2804);
nand UO_433 (O_433,N_2293,N_2930);
nand UO_434 (O_434,N_2589,N_2872);
and UO_435 (O_435,N_2955,N_2324);
xor UO_436 (O_436,N_2517,N_2745);
and UO_437 (O_437,N_2278,N_2259);
and UO_438 (O_438,N_2710,N_2820);
nand UO_439 (O_439,N_2437,N_2826);
nor UO_440 (O_440,N_2487,N_2460);
xnor UO_441 (O_441,N_2708,N_2372);
or UO_442 (O_442,N_2607,N_2595);
nor UO_443 (O_443,N_2803,N_2900);
or UO_444 (O_444,N_2297,N_2417);
or UO_445 (O_445,N_2351,N_2685);
or UO_446 (O_446,N_2727,N_2831);
xnor UO_447 (O_447,N_2719,N_2746);
and UO_448 (O_448,N_2812,N_2549);
and UO_449 (O_449,N_2508,N_2356);
nor UO_450 (O_450,N_2671,N_2453);
or UO_451 (O_451,N_2658,N_2278);
nor UO_452 (O_452,N_2714,N_2796);
xnor UO_453 (O_453,N_2733,N_2762);
nor UO_454 (O_454,N_2960,N_2965);
nor UO_455 (O_455,N_2255,N_2537);
and UO_456 (O_456,N_2791,N_2838);
nand UO_457 (O_457,N_2554,N_2274);
and UO_458 (O_458,N_2914,N_2929);
or UO_459 (O_459,N_2754,N_2823);
or UO_460 (O_460,N_2362,N_2728);
nor UO_461 (O_461,N_2448,N_2655);
or UO_462 (O_462,N_2726,N_2711);
nand UO_463 (O_463,N_2839,N_2258);
nand UO_464 (O_464,N_2381,N_2913);
xnor UO_465 (O_465,N_2684,N_2268);
nand UO_466 (O_466,N_2503,N_2418);
or UO_467 (O_467,N_2842,N_2838);
or UO_468 (O_468,N_2250,N_2557);
xnor UO_469 (O_469,N_2920,N_2683);
nor UO_470 (O_470,N_2545,N_2949);
xnor UO_471 (O_471,N_2501,N_2921);
xor UO_472 (O_472,N_2945,N_2451);
and UO_473 (O_473,N_2933,N_2676);
nand UO_474 (O_474,N_2666,N_2285);
xnor UO_475 (O_475,N_2271,N_2997);
or UO_476 (O_476,N_2884,N_2796);
and UO_477 (O_477,N_2544,N_2449);
xor UO_478 (O_478,N_2654,N_2586);
and UO_479 (O_479,N_2386,N_2850);
and UO_480 (O_480,N_2675,N_2623);
and UO_481 (O_481,N_2985,N_2413);
xnor UO_482 (O_482,N_2337,N_2362);
nor UO_483 (O_483,N_2277,N_2454);
xor UO_484 (O_484,N_2387,N_2807);
xor UO_485 (O_485,N_2678,N_2845);
nor UO_486 (O_486,N_2621,N_2991);
and UO_487 (O_487,N_2897,N_2954);
nand UO_488 (O_488,N_2899,N_2465);
or UO_489 (O_489,N_2638,N_2463);
xnor UO_490 (O_490,N_2408,N_2627);
xor UO_491 (O_491,N_2483,N_2665);
nand UO_492 (O_492,N_2595,N_2304);
nor UO_493 (O_493,N_2887,N_2505);
nor UO_494 (O_494,N_2292,N_2425);
xor UO_495 (O_495,N_2549,N_2393);
nor UO_496 (O_496,N_2545,N_2565);
or UO_497 (O_497,N_2375,N_2358);
nand UO_498 (O_498,N_2942,N_2407);
or UO_499 (O_499,N_2800,N_2889);
endmodule