module basic_500_3000_500_5_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_248,In_71);
or U1 (N_1,In_418,In_433);
nand U2 (N_2,In_67,In_470);
nand U3 (N_3,In_360,In_320);
or U4 (N_4,In_337,In_472);
and U5 (N_5,In_366,In_180);
nor U6 (N_6,In_175,In_440);
nand U7 (N_7,In_200,In_16);
or U8 (N_8,In_377,In_24);
nor U9 (N_9,In_93,In_140);
and U10 (N_10,In_295,In_454);
nand U11 (N_11,In_88,In_239);
nor U12 (N_12,In_261,In_282);
and U13 (N_13,In_263,In_374);
or U14 (N_14,In_460,In_149);
or U15 (N_15,In_9,In_475);
and U16 (N_16,In_420,In_403);
and U17 (N_17,In_43,In_449);
or U18 (N_18,In_354,In_498);
and U19 (N_19,In_342,In_307);
or U20 (N_20,In_206,In_353);
and U21 (N_21,In_400,In_404);
nand U22 (N_22,In_183,In_283);
nor U23 (N_23,In_350,In_123);
or U24 (N_24,In_170,In_486);
or U25 (N_25,In_333,In_61);
nor U26 (N_26,In_119,In_101);
nand U27 (N_27,In_151,In_284);
nand U28 (N_28,In_301,In_122);
nor U29 (N_29,In_227,In_421);
or U30 (N_30,In_18,In_458);
nand U31 (N_31,In_96,In_330);
and U32 (N_32,In_461,In_201);
nor U33 (N_33,In_316,In_436);
nand U34 (N_34,In_304,In_429);
nand U35 (N_35,In_121,In_255);
or U36 (N_36,In_424,In_469);
or U37 (N_37,In_174,In_62);
and U38 (N_38,In_51,In_185);
nand U39 (N_39,In_318,In_172);
or U40 (N_40,In_91,In_252);
or U41 (N_41,In_192,In_438);
nand U42 (N_42,In_467,In_484);
xor U43 (N_43,In_89,In_463);
nand U44 (N_44,In_146,In_285);
nor U45 (N_45,In_4,In_395);
or U46 (N_46,In_387,In_173);
and U47 (N_47,In_102,In_265);
nor U48 (N_48,In_323,In_362);
or U49 (N_49,In_321,In_226);
nor U50 (N_50,In_439,In_124);
or U51 (N_51,In_390,In_292);
or U52 (N_52,In_363,In_343);
nand U53 (N_53,In_215,In_459);
and U54 (N_54,In_311,In_225);
nor U55 (N_55,In_234,In_299);
or U56 (N_56,In_340,In_15);
nor U57 (N_57,In_270,In_468);
or U58 (N_58,In_237,In_69);
nor U59 (N_59,In_254,In_46);
and U60 (N_60,In_312,In_29);
or U61 (N_61,In_138,In_55);
and U62 (N_62,In_257,In_245);
and U63 (N_63,In_189,In_352);
nor U64 (N_64,In_148,In_481);
nand U65 (N_65,In_332,In_150);
nor U66 (N_66,In_266,In_0);
nor U67 (N_67,In_157,In_359);
nand U68 (N_68,In_488,In_203);
nor U69 (N_69,In_313,In_40);
and U70 (N_70,In_217,In_75);
nand U71 (N_71,In_346,In_73);
nand U72 (N_72,In_218,In_52);
nand U73 (N_73,In_106,In_479);
and U74 (N_74,In_5,In_464);
or U75 (N_75,In_166,In_11);
or U76 (N_76,In_159,In_267);
and U77 (N_77,In_129,In_365);
or U78 (N_78,In_153,In_385);
nor U79 (N_79,In_202,In_405);
nor U80 (N_80,In_378,In_494);
nand U81 (N_81,In_489,In_394);
nand U82 (N_82,In_358,In_383);
nor U83 (N_83,In_347,In_31);
nand U84 (N_84,In_128,In_45);
and U85 (N_85,In_289,In_407);
and U86 (N_86,In_372,In_81);
or U87 (N_87,In_274,In_431);
nand U88 (N_88,In_36,In_286);
or U89 (N_89,In_115,In_13);
nor U90 (N_90,In_238,In_413);
nand U91 (N_91,In_462,In_416);
nand U92 (N_92,In_490,In_72);
nand U93 (N_93,In_209,In_57);
xor U94 (N_94,In_341,In_240);
and U95 (N_95,In_262,In_97);
nand U96 (N_96,In_275,In_210);
nand U97 (N_97,In_497,In_94);
or U98 (N_98,In_432,In_406);
nand U99 (N_99,In_14,In_367);
nor U100 (N_100,In_241,In_145);
or U101 (N_101,In_477,In_41);
nor U102 (N_102,In_34,In_117);
and U103 (N_103,In_103,In_398);
and U104 (N_104,In_6,In_39);
nor U105 (N_105,In_434,In_345);
nand U106 (N_106,In_92,In_393);
nand U107 (N_107,In_22,In_132);
nor U108 (N_108,In_338,In_483);
nand U109 (N_109,In_49,In_308);
or U110 (N_110,In_130,In_325);
or U111 (N_111,In_373,In_348);
or U112 (N_112,In_59,In_380);
nand U113 (N_113,In_277,In_253);
or U114 (N_114,In_496,In_471);
or U115 (N_115,In_356,In_164);
and U116 (N_116,In_491,In_379);
and U117 (N_117,In_44,In_12);
nand U118 (N_118,In_281,In_8);
nor U119 (N_119,In_453,In_176);
nand U120 (N_120,In_137,In_2);
or U121 (N_121,In_17,In_370);
nand U122 (N_122,In_371,In_120);
or U123 (N_123,In_99,In_474);
nor U124 (N_124,In_317,In_30);
nand U125 (N_125,In_473,In_271);
or U126 (N_126,In_198,In_273);
and U127 (N_127,In_264,In_194);
nor U128 (N_128,In_376,In_455);
or U129 (N_129,In_127,In_53);
nor U130 (N_130,In_391,In_162);
xor U131 (N_131,In_205,In_80);
or U132 (N_132,In_452,In_351);
or U133 (N_133,In_110,In_314);
and U134 (N_134,In_178,In_139);
and U135 (N_135,In_408,In_77);
or U136 (N_136,In_169,In_65);
or U137 (N_137,In_384,In_3);
or U138 (N_138,In_446,In_50);
nor U139 (N_139,In_193,In_269);
nor U140 (N_140,In_278,In_95);
or U141 (N_141,In_165,In_293);
nand U142 (N_142,In_20,In_48);
nor U143 (N_143,In_224,In_279);
or U144 (N_144,In_154,In_242);
nand U145 (N_145,In_415,In_231);
nor U146 (N_146,In_297,In_256);
xor U147 (N_147,In_287,In_179);
or U148 (N_148,In_76,In_211);
nand U149 (N_149,In_63,In_331);
nor U150 (N_150,In_168,In_381);
and U151 (N_151,In_250,In_195);
nand U152 (N_152,In_223,In_186);
nand U153 (N_153,In_339,In_156);
or U154 (N_154,In_136,In_221);
and U155 (N_155,In_199,In_143);
nor U156 (N_156,In_290,In_485);
and U157 (N_157,In_228,In_357);
nor U158 (N_158,In_329,In_147);
nand U159 (N_159,In_98,In_422);
or U160 (N_160,In_300,In_399);
and U161 (N_161,In_430,In_161);
or U162 (N_162,In_104,In_260);
or U163 (N_163,In_495,In_19);
or U164 (N_164,In_60,In_303);
or U165 (N_165,In_204,In_197);
nand U166 (N_166,In_326,In_451);
nand U167 (N_167,In_155,In_111);
and U168 (N_168,In_216,In_448);
and U169 (N_169,In_276,In_410);
or U170 (N_170,In_447,In_492);
or U171 (N_171,In_84,In_435);
or U172 (N_172,In_369,In_37);
nor U173 (N_173,In_389,In_327);
nand U174 (N_174,In_82,In_392);
and U175 (N_175,In_427,In_133);
nor U176 (N_176,In_58,In_291);
or U177 (N_177,In_465,In_114);
or U178 (N_178,In_280,In_296);
or U179 (N_179,In_401,In_414);
nand U180 (N_180,In_184,In_361);
nor U181 (N_181,In_268,In_107);
nand U182 (N_182,In_334,In_412);
nor U183 (N_183,In_74,In_220);
and U184 (N_184,In_397,In_78);
nor U185 (N_185,In_409,In_402);
or U186 (N_186,In_87,In_417);
nor U187 (N_187,In_294,In_190);
nor U188 (N_188,In_426,In_466);
or U189 (N_189,In_131,In_244);
xor U190 (N_190,In_368,In_382);
or U191 (N_191,In_437,In_444);
nand U192 (N_192,In_152,In_324);
nor U193 (N_193,In_336,In_26);
nand U194 (N_194,In_315,In_142);
or U195 (N_195,In_236,In_79);
nor U196 (N_196,In_457,In_298);
nand U197 (N_197,In_83,In_135);
nand U198 (N_198,In_476,In_27);
nor U199 (N_199,In_158,In_28);
or U200 (N_200,In_355,In_134);
or U201 (N_201,In_493,In_70);
or U202 (N_202,In_441,In_112);
nand U203 (N_203,In_456,In_181);
nor U204 (N_204,In_232,In_419);
nand U205 (N_205,In_42,In_196);
xnor U206 (N_206,In_126,In_310);
and U207 (N_207,In_25,In_23);
xor U208 (N_208,In_125,In_33);
nor U209 (N_209,In_246,In_251);
nor U210 (N_210,In_349,In_212);
or U211 (N_211,In_482,In_259);
nand U212 (N_212,In_233,In_10);
or U213 (N_213,In_109,In_38);
nor U214 (N_214,In_105,In_375);
nand U215 (N_215,In_425,In_66);
nand U216 (N_216,In_100,In_163);
and U217 (N_217,In_208,In_35);
nor U218 (N_218,In_272,In_423);
nor U219 (N_219,In_54,In_480);
or U220 (N_220,In_249,In_86);
nand U221 (N_221,In_396,In_56);
and U222 (N_222,In_305,In_230);
nand U223 (N_223,In_428,In_344);
or U224 (N_224,In_214,In_411);
nand U225 (N_225,In_116,In_443);
nor U226 (N_226,In_328,In_187);
nand U227 (N_227,In_177,In_335);
nor U228 (N_228,In_302,In_213);
nor U229 (N_229,In_90,In_118);
nor U230 (N_230,In_182,In_188);
nor U231 (N_231,In_364,In_309);
and U232 (N_232,In_167,In_499);
nor U233 (N_233,In_21,In_442);
and U234 (N_234,In_319,In_113);
nor U235 (N_235,In_306,In_386);
or U236 (N_236,In_32,In_235);
nand U237 (N_237,In_1,In_322);
xnor U238 (N_238,In_207,In_258);
or U239 (N_239,In_288,In_7);
nand U240 (N_240,In_68,In_108);
nor U241 (N_241,In_144,In_478);
nor U242 (N_242,In_487,In_243);
and U243 (N_243,In_219,In_229);
nor U244 (N_244,In_222,In_160);
or U245 (N_245,In_388,In_64);
nor U246 (N_246,In_450,In_445);
and U247 (N_247,In_85,In_247);
or U248 (N_248,In_141,In_171);
or U249 (N_249,In_191,In_47);
or U250 (N_250,In_288,In_272);
and U251 (N_251,In_423,In_46);
nand U252 (N_252,In_104,In_413);
nand U253 (N_253,In_466,In_414);
or U254 (N_254,In_419,In_426);
and U255 (N_255,In_73,In_65);
or U256 (N_256,In_145,In_30);
nor U257 (N_257,In_398,In_471);
and U258 (N_258,In_14,In_208);
and U259 (N_259,In_68,In_224);
nor U260 (N_260,In_262,In_114);
or U261 (N_261,In_374,In_63);
or U262 (N_262,In_80,In_7);
nand U263 (N_263,In_400,In_484);
nand U264 (N_264,In_205,In_229);
or U265 (N_265,In_452,In_364);
nand U266 (N_266,In_286,In_206);
nor U267 (N_267,In_120,In_476);
and U268 (N_268,In_27,In_65);
or U269 (N_269,In_256,In_72);
or U270 (N_270,In_188,In_353);
and U271 (N_271,In_399,In_229);
or U272 (N_272,In_321,In_363);
nor U273 (N_273,In_222,In_152);
or U274 (N_274,In_211,In_312);
nand U275 (N_275,In_81,In_114);
nand U276 (N_276,In_79,In_275);
or U277 (N_277,In_120,In_366);
nor U278 (N_278,In_301,In_344);
nand U279 (N_279,In_393,In_428);
nand U280 (N_280,In_419,In_284);
or U281 (N_281,In_364,In_449);
and U282 (N_282,In_217,In_339);
nor U283 (N_283,In_293,In_250);
or U284 (N_284,In_311,In_430);
nor U285 (N_285,In_298,In_211);
nor U286 (N_286,In_223,In_91);
nor U287 (N_287,In_388,In_254);
or U288 (N_288,In_161,In_203);
nand U289 (N_289,In_368,In_80);
nand U290 (N_290,In_88,In_437);
or U291 (N_291,In_258,In_166);
nand U292 (N_292,In_392,In_487);
nand U293 (N_293,In_338,In_496);
or U294 (N_294,In_310,In_271);
nand U295 (N_295,In_178,In_382);
and U296 (N_296,In_204,In_157);
nor U297 (N_297,In_63,In_22);
nand U298 (N_298,In_432,In_463);
or U299 (N_299,In_47,In_412);
nand U300 (N_300,In_68,In_5);
or U301 (N_301,In_251,In_51);
or U302 (N_302,In_56,In_267);
and U303 (N_303,In_244,In_409);
and U304 (N_304,In_393,In_98);
nor U305 (N_305,In_30,In_148);
nand U306 (N_306,In_190,In_168);
or U307 (N_307,In_212,In_163);
and U308 (N_308,In_82,In_132);
nor U309 (N_309,In_301,In_328);
or U310 (N_310,In_400,In_470);
nand U311 (N_311,In_17,In_193);
xor U312 (N_312,In_440,In_138);
and U313 (N_313,In_385,In_216);
nand U314 (N_314,In_493,In_320);
and U315 (N_315,In_136,In_53);
or U316 (N_316,In_493,In_162);
and U317 (N_317,In_23,In_282);
or U318 (N_318,In_27,In_14);
and U319 (N_319,In_237,In_267);
nor U320 (N_320,In_385,In_104);
or U321 (N_321,In_93,In_480);
nand U322 (N_322,In_147,In_446);
and U323 (N_323,In_434,In_290);
and U324 (N_324,In_491,In_372);
and U325 (N_325,In_458,In_272);
or U326 (N_326,In_270,In_268);
and U327 (N_327,In_184,In_308);
or U328 (N_328,In_458,In_286);
and U329 (N_329,In_71,In_196);
nand U330 (N_330,In_493,In_311);
and U331 (N_331,In_82,In_127);
nand U332 (N_332,In_323,In_144);
or U333 (N_333,In_299,In_270);
and U334 (N_334,In_349,In_389);
nand U335 (N_335,In_414,In_15);
nor U336 (N_336,In_92,In_351);
nor U337 (N_337,In_302,In_470);
and U338 (N_338,In_163,In_127);
nand U339 (N_339,In_383,In_136);
nor U340 (N_340,In_31,In_279);
nand U341 (N_341,In_299,In_272);
and U342 (N_342,In_213,In_381);
nor U343 (N_343,In_312,In_174);
nand U344 (N_344,In_300,In_277);
nand U345 (N_345,In_262,In_271);
nor U346 (N_346,In_489,In_434);
or U347 (N_347,In_240,In_340);
and U348 (N_348,In_81,In_343);
nor U349 (N_349,In_129,In_340);
nand U350 (N_350,In_146,In_3);
nand U351 (N_351,In_436,In_435);
and U352 (N_352,In_219,In_33);
nand U353 (N_353,In_307,In_68);
or U354 (N_354,In_279,In_302);
nor U355 (N_355,In_363,In_257);
or U356 (N_356,In_449,In_356);
or U357 (N_357,In_375,In_368);
and U358 (N_358,In_107,In_412);
or U359 (N_359,In_453,In_218);
nor U360 (N_360,In_413,In_308);
and U361 (N_361,In_440,In_80);
or U362 (N_362,In_62,In_153);
and U363 (N_363,In_157,In_297);
or U364 (N_364,In_85,In_232);
nor U365 (N_365,In_320,In_103);
and U366 (N_366,In_360,In_333);
or U367 (N_367,In_416,In_108);
nand U368 (N_368,In_50,In_475);
and U369 (N_369,In_244,In_382);
nand U370 (N_370,In_195,In_494);
nor U371 (N_371,In_331,In_329);
or U372 (N_372,In_50,In_443);
and U373 (N_373,In_309,In_477);
nand U374 (N_374,In_213,In_161);
nor U375 (N_375,In_296,In_407);
xor U376 (N_376,In_349,In_191);
nor U377 (N_377,In_304,In_351);
xor U378 (N_378,In_24,In_172);
nor U379 (N_379,In_392,In_254);
and U380 (N_380,In_167,In_416);
and U381 (N_381,In_371,In_354);
or U382 (N_382,In_448,In_232);
and U383 (N_383,In_126,In_141);
nand U384 (N_384,In_383,In_379);
nor U385 (N_385,In_351,In_212);
nor U386 (N_386,In_75,In_260);
nor U387 (N_387,In_247,In_300);
and U388 (N_388,In_430,In_485);
nor U389 (N_389,In_418,In_274);
nand U390 (N_390,In_361,In_76);
and U391 (N_391,In_162,In_89);
nand U392 (N_392,In_140,In_328);
nand U393 (N_393,In_106,In_402);
nor U394 (N_394,In_426,In_69);
nor U395 (N_395,In_96,In_179);
nand U396 (N_396,In_33,In_205);
xor U397 (N_397,In_134,In_294);
nor U398 (N_398,In_128,In_211);
or U399 (N_399,In_490,In_485);
nor U400 (N_400,In_424,In_68);
or U401 (N_401,In_261,In_415);
nand U402 (N_402,In_491,In_187);
or U403 (N_403,In_266,In_120);
nand U404 (N_404,In_61,In_88);
or U405 (N_405,In_15,In_168);
nand U406 (N_406,In_238,In_16);
nand U407 (N_407,In_79,In_191);
nand U408 (N_408,In_327,In_204);
and U409 (N_409,In_189,In_162);
and U410 (N_410,In_333,In_75);
nor U411 (N_411,In_14,In_393);
xor U412 (N_412,In_7,In_69);
and U413 (N_413,In_381,In_282);
nand U414 (N_414,In_368,In_267);
nor U415 (N_415,In_465,In_276);
or U416 (N_416,In_419,In_255);
and U417 (N_417,In_295,In_185);
nor U418 (N_418,In_466,In_105);
nor U419 (N_419,In_399,In_129);
and U420 (N_420,In_315,In_125);
nand U421 (N_421,In_101,In_283);
or U422 (N_422,In_171,In_10);
nor U423 (N_423,In_159,In_162);
or U424 (N_424,In_328,In_289);
and U425 (N_425,In_392,In_459);
nor U426 (N_426,In_293,In_15);
nand U427 (N_427,In_384,In_219);
and U428 (N_428,In_88,In_184);
nor U429 (N_429,In_38,In_344);
nor U430 (N_430,In_456,In_445);
or U431 (N_431,In_312,In_299);
and U432 (N_432,In_64,In_185);
nor U433 (N_433,In_8,In_187);
xor U434 (N_434,In_182,In_366);
nand U435 (N_435,In_439,In_307);
and U436 (N_436,In_19,In_493);
nor U437 (N_437,In_9,In_256);
and U438 (N_438,In_497,In_407);
nand U439 (N_439,In_497,In_273);
or U440 (N_440,In_2,In_173);
nand U441 (N_441,In_193,In_397);
or U442 (N_442,In_482,In_475);
nand U443 (N_443,In_279,In_23);
nand U444 (N_444,In_224,In_223);
and U445 (N_445,In_353,In_493);
and U446 (N_446,In_244,In_203);
or U447 (N_447,In_90,In_174);
or U448 (N_448,In_126,In_111);
and U449 (N_449,In_50,In_144);
nor U450 (N_450,In_480,In_132);
nand U451 (N_451,In_324,In_468);
nor U452 (N_452,In_489,In_456);
nand U453 (N_453,In_272,In_211);
nor U454 (N_454,In_387,In_323);
or U455 (N_455,In_31,In_422);
or U456 (N_456,In_455,In_124);
or U457 (N_457,In_422,In_43);
or U458 (N_458,In_283,In_80);
and U459 (N_459,In_233,In_397);
and U460 (N_460,In_448,In_480);
or U461 (N_461,In_52,In_350);
or U462 (N_462,In_120,In_82);
and U463 (N_463,In_413,In_117);
nand U464 (N_464,In_22,In_230);
and U465 (N_465,In_460,In_466);
nor U466 (N_466,In_439,In_152);
or U467 (N_467,In_149,In_432);
nor U468 (N_468,In_384,In_137);
or U469 (N_469,In_448,In_329);
or U470 (N_470,In_191,In_320);
and U471 (N_471,In_230,In_346);
or U472 (N_472,In_449,In_434);
and U473 (N_473,In_454,In_18);
or U474 (N_474,In_108,In_181);
nor U475 (N_475,In_282,In_129);
and U476 (N_476,In_456,In_110);
nand U477 (N_477,In_164,In_129);
or U478 (N_478,In_54,In_5);
xnor U479 (N_479,In_433,In_150);
nor U480 (N_480,In_352,In_365);
and U481 (N_481,In_424,In_100);
nor U482 (N_482,In_240,In_401);
nand U483 (N_483,In_443,In_282);
and U484 (N_484,In_462,In_181);
nor U485 (N_485,In_90,In_230);
nand U486 (N_486,In_323,In_104);
nor U487 (N_487,In_36,In_231);
and U488 (N_488,In_49,In_383);
nand U489 (N_489,In_116,In_338);
nand U490 (N_490,In_368,In_221);
nor U491 (N_491,In_360,In_17);
and U492 (N_492,In_275,In_135);
nor U493 (N_493,In_86,In_300);
or U494 (N_494,In_59,In_200);
nor U495 (N_495,In_149,In_317);
nor U496 (N_496,In_178,In_458);
or U497 (N_497,In_364,In_155);
nor U498 (N_498,In_233,In_268);
nor U499 (N_499,In_456,In_299);
or U500 (N_500,In_172,In_144);
or U501 (N_501,In_405,In_300);
and U502 (N_502,In_222,In_253);
nand U503 (N_503,In_329,In_60);
nand U504 (N_504,In_124,In_461);
or U505 (N_505,In_64,In_130);
or U506 (N_506,In_431,In_403);
and U507 (N_507,In_468,In_195);
or U508 (N_508,In_347,In_344);
and U509 (N_509,In_103,In_288);
or U510 (N_510,In_458,In_329);
xor U511 (N_511,In_283,In_299);
nand U512 (N_512,In_323,In_40);
nand U513 (N_513,In_197,In_356);
and U514 (N_514,In_98,In_161);
or U515 (N_515,In_371,In_411);
nand U516 (N_516,In_23,In_37);
nor U517 (N_517,In_84,In_54);
or U518 (N_518,In_259,In_229);
nor U519 (N_519,In_244,In_472);
or U520 (N_520,In_434,In_363);
or U521 (N_521,In_50,In_311);
nor U522 (N_522,In_121,In_320);
nand U523 (N_523,In_394,In_134);
nand U524 (N_524,In_414,In_120);
nand U525 (N_525,In_136,In_140);
and U526 (N_526,In_125,In_396);
nand U527 (N_527,In_206,In_31);
xor U528 (N_528,In_2,In_206);
nand U529 (N_529,In_329,In_6);
nor U530 (N_530,In_192,In_380);
and U531 (N_531,In_198,In_497);
and U532 (N_532,In_157,In_198);
or U533 (N_533,In_208,In_238);
and U534 (N_534,In_136,In_199);
and U535 (N_535,In_491,In_172);
nand U536 (N_536,In_365,In_404);
nand U537 (N_537,In_51,In_336);
or U538 (N_538,In_296,In_251);
or U539 (N_539,In_113,In_39);
nor U540 (N_540,In_168,In_77);
nand U541 (N_541,In_287,In_358);
nand U542 (N_542,In_74,In_12);
or U543 (N_543,In_113,In_488);
and U544 (N_544,In_321,In_326);
or U545 (N_545,In_239,In_337);
or U546 (N_546,In_465,In_218);
or U547 (N_547,In_31,In_33);
or U548 (N_548,In_273,In_329);
or U549 (N_549,In_188,In_372);
nand U550 (N_550,In_408,In_130);
and U551 (N_551,In_181,In_255);
and U552 (N_552,In_237,In_357);
and U553 (N_553,In_328,In_337);
and U554 (N_554,In_135,In_43);
or U555 (N_555,In_280,In_83);
nand U556 (N_556,In_318,In_129);
nor U557 (N_557,In_109,In_197);
nand U558 (N_558,In_347,In_238);
and U559 (N_559,In_304,In_19);
nor U560 (N_560,In_207,In_181);
nor U561 (N_561,In_300,In_486);
or U562 (N_562,In_118,In_388);
or U563 (N_563,In_378,In_200);
nand U564 (N_564,In_54,In_57);
or U565 (N_565,In_241,In_489);
or U566 (N_566,In_145,In_194);
or U567 (N_567,In_14,In_370);
and U568 (N_568,In_235,In_319);
or U569 (N_569,In_390,In_342);
or U570 (N_570,In_300,In_210);
nor U571 (N_571,In_401,In_324);
or U572 (N_572,In_347,In_196);
and U573 (N_573,In_246,In_267);
nand U574 (N_574,In_471,In_26);
nor U575 (N_575,In_46,In_387);
nand U576 (N_576,In_85,In_435);
nor U577 (N_577,In_142,In_379);
and U578 (N_578,In_167,In_498);
nor U579 (N_579,In_124,In_107);
and U580 (N_580,In_86,In_351);
or U581 (N_581,In_475,In_27);
nor U582 (N_582,In_108,In_312);
and U583 (N_583,In_244,In_5);
and U584 (N_584,In_314,In_354);
and U585 (N_585,In_238,In_53);
nand U586 (N_586,In_40,In_248);
and U587 (N_587,In_264,In_222);
or U588 (N_588,In_406,In_322);
nand U589 (N_589,In_145,In_84);
nor U590 (N_590,In_97,In_118);
nand U591 (N_591,In_455,In_106);
nor U592 (N_592,In_321,In_173);
and U593 (N_593,In_304,In_242);
and U594 (N_594,In_23,In_222);
and U595 (N_595,In_299,In_317);
xor U596 (N_596,In_83,In_62);
and U597 (N_597,In_222,In_134);
nor U598 (N_598,In_207,In_17);
nand U599 (N_599,In_11,In_367);
and U600 (N_600,N_72,N_467);
or U601 (N_601,N_594,N_169);
and U602 (N_602,N_228,N_272);
or U603 (N_603,N_57,N_273);
nor U604 (N_604,N_490,N_581);
nor U605 (N_605,N_363,N_444);
nand U606 (N_606,N_91,N_203);
nand U607 (N_607,N_542,N_144);
or U608 (N_608,N_351,N_449);
nor U609 (N_609,N_428,N_156);
or U610 (N_610,N_382,N_567);
nor U611 (N_611,N_450,N_580);
or U612 (N_612,N_284,N_410);
nand U613 (N_613,N_385,N_9);
and U614 (N_614,N_310,N_359);
nor U615 (N_615,N_174,N_298);
nor U616 (N_616,N_507,N_308);
nor U617 (N_617,N_239,N_141);
nand U618 (N_618,N_333,N_213);
or U619 (N_619,N_271,N_160);
or U620 (N_620,N_69,N_297);
and U621 (N_621,N_430,N_122);
nor U622 (N_622,N_397,N_421);
nor U623 (N_623,N_199,N_570);
xor U624 (N_624,N_353,N_51);
and U625 (N_625,N_322,N_586);
nand U626 (N_626,N_488,N_223);
or U627 (N_627,N_220,N_42);
and U628 (N_628,N_14,N_23);
nand U629 (N_629,N_13,N_90);
and U630 (N_630,N_403,N_126);
nand U631 (N_631,N_264,N_167);
nor U632 (N_632,N_435,N_139);
nor U633 (N_633,N_320,N_202);
and U634 (N_634,N_509,N_423);
or U635 (N_635,N_283,N_473);
and U636 (N_636,N_43,N_548);
and U637 (N_637,N_99,N_103);
xor U638 (N_638,N_577,N_270);
or U639 (N_639,N_74,N_439);
nand U640 (N_640,N_562,N_536);
nor U641 (N_641,N_288,N_335);
nand U642 (N_642,N_15,N_392);
and U643 (N_643,N_313,N_304);
nand U644 (N_644,N_314,N_242);
nor U645 (N_645,N_268,N_471);
or U646 (N_646,N_376,N_131);
nand U647 (N_647,N_62,N_215);
or U648 (N_648,N_412,N_218);
or U649 (N_649,N_535,N_157);
nor U650 (N_650,N_550,N_521);
or U651 (N_651,N_360,N_495);
nand U652 (N_652,N_528,N_425);
and U653 (N_653,N_316,N_94);
nand U654 (N_654,N_433,N_390);
and U655 (N_655,N_575,N_455);
nand U656 (N_656,N_135,N_451);
and U657 (N_657,N_16,N_311);
nor U658 (N_658,N_501,N_492);
nor U659 (N_659,N_484,N_250);
or U660 (N_660,N_201,N_188);
nor U661 (N_661,N_422,N_491);
nand U662 (N_662,N_357,N_7);
nand U663 (N_663,N_34,N_315);
and U664 (N_664,N_513,N_192);
nand U665 (N_665,N_365,N_306);
nor U666 (N_666,N_50,N_463);
nor U667 (N_667,N_367,N_378);
nand U668 (N_668,N_416,N_545);
and U669 (N_669,N_185,N_325);
nor U670 (N_670,N_35,N_456);
nor U671 (N_671,N_443,N_517);
nor U672 (N_672,N_248,N_373);
and U673 (N_673,N_532,N_583);
nand U674 (N_674,N_190,N_401);
or U675 (N_675,N_398,N_53);
or U676 (N_676,N_66,N_393);
or U677 (N_677,N_33,N_279);
nand U678 (N_678,N_476,N_10);
and U679 (N_679,N_565,N_596);
nor U680 (N_680,N_136,N_205);
nor U681 (N_681,N_132,N_123);
nor U682 (N_682,N_25,N_415);
or U683 (N_683,N_65,N_183);
nand U684 (N_684,N_175,N_510);
or U685 (N_685,N_159,N_41);
nand U686 (N_686,N_151,N_511);
and U687 (N_687,N_252,N_529);
nor U688 (N_688,N_564,N_38);
nor U689 (N_689,N_82,N_275);
nand U690 (N_690,N_24,N_28);
nor U691 (N_691,N_278,N_245);
nor U692 (N_692,N_453,N_55);
nor U693 (N_693,N_481,N_193);
and U694 (N_694,N_194,N_552);
nor U695 (N_695,N_478,N_85);
or U696 (N_696,N_520,N_262);
nor U697 (N_697,N_303,N_299);
and U698 (N_698,N_461,N_39);
nor U699 (N_699,N_436,N_219);
nand U700 (N_700,N_572,N_114);
and U701 (N_701,N_234,N_502);
and U702 (N_702,N_8,N_258);
nor U703 (N_703,N_230,N_447);
nand U704 (N_704,N_457,N_187);
or U705 (N_705,N_4,N_196);
nor U706 (N_706,N_296,N_568);
nand U707 (N_707,N_249,N_500);
nor U708 (N_708,N_533,N_130);
and U709 (N_709,N_247,N_89);
nand U710 (N_710,N_599,N_485);
or U711 (N_711,N_374,N_327);
or U712 (N_712,N_379,N_76);
nand U713 (N_713,N_530,N_543);
nor U714 (N_714,N_56,N_197);
nor U715 (N_715,N_79,N_20);
nor U716 (N_716,N_343,N_493);
nor U717 (N_717,N_186,N_224);
and U718 (N_718,N_285,N_368);
and U719 (N_719,N_98,N_445);
and U720 (N_720,N_526,N_408);
or U721 (N_721,N_387,N_380);
nand U722 (N_722,N_150,N_300);
or U723 (N_723,N_503,N_30);
or U724 (N_724,N_576,N_420);
nor U725 (N_725,N_579,N_255);
nand U726 (N_726,N_221,N_515);
nand U727 (N_727,N_217,N_358);
nor U728 (N_728,N_554,N_229);
nor U729 (N_729,N_340,N_329);
or U730 (N_730,N_138,N_319);
nand U731 (N_731,N_177,N_95);
nand U732 (N_732,N_287,N_514);
nand U733 (N_733,N_102,N_163);
nor U734 (N_734,N_483,N_466);
nor U735 (N_735,N_330,N_556);
and U736 (N_736,N_180,N_96);
nor U737 (N_737,N_231,N_563);
or U738 (N_738,N_469,N_555);
or U739 (N_739,N_71,N_290);
nor U740 (N_740,N_505,N_46);
nand U741 (N_741,N_411,N_566);
nand U742 (N_742,N_326,N_595);
nor U743 (N_743,N_384,N_291);
or U744 (N_744,N_464,N_208);
nand U745 (N_745,N_178,N_107);
and U746 (N_746,N_154,N_116);
nor U747 (N_747,N_1,N_539);
nor U748 (N_748,N_40,N_588);
nor U749 (N_749,N_371,N_352);
or U750 (N_750,N_585,N_31);
nand U751 (N_751,N_64,N_386);
nor U752 (N_752,N_155,N_369);
or U753 (N_753,N_170,N_269);
nor U754 (N_754,N_328,N_274);
and U755 (N_755,N_293,N_171);
or U756 (N_756,N_312,N_342);
or U757 (N_757,N_332,N_182);
nand U758 (N_758,N_350,N_537);
nand U759 (N_759,N_149,N_336);
and U760 (N_760,N_119,N_477);
and U761 (N_761,N_260,N_204);
and U762 (N_762,N_582,N_244);
or U763 (N_763,N_84,N_60);
nor U764 (N_764,N_142,N_121);
or U765 (N_765,N_222,N_210);
nor U766 (N_766,N_519,N_525);
or U767 (N_767,N_59,N_452);
and U768 (N_768,N_26,N_446);
nand U769 (N_769,N_323,N_573);
and U770 (N_770,N_97,N_482);
and U771 (N_771,N_129,N_292);
nand U772 (N_772,N_191,N_117);
nor U773 (N_773,N_294,N_541);
nand U774 (N_774,N_338,N_251);
nand U775 (N_775,N_404,N_337);
nand U776 (N_776,N_152,N_118);
nor U777 (N_777,N_47,N_302);
nor U778 (N_778,N_459,N_189);
and U779 (N_779,N_597,N_240);
or U780 (N_780,N_557,N_354);
nor U781 (N_781,N_276,N_394);
nand U782 (N_782,N_124,N_140);
or U783 (N_783,N_516,N_77);
and U784 (N_784,N_465,N_238);
or U785 (N_785,N_93,N_441);
and U786 (N_786,N_402,N_61);
and U787 (N_787,N_17,N_438);
nor U788 (N_788,N_396,N_364);
or U789 (N_789,N_437,N_105);
nand U790 (N_790,N_518,N_113);
or U791 (N_791,N_591,N_207);
nor U792 (N_792,N_560,N_27);
nand U793 (N_793,N_589,N_499);
or U794 (N_794,N_19,N_246);
nor U795 (N_795,N_417,N_143);
nor U796 (N_796,N_468,N_317);
nand U797 (N_797,N_256,N_389);
nand U798 (N_798,N_558,N_106);
nor U799 (N_799,N_486,N_263);
nor U800 (N_800,N_128,N_508);
or U801 (N_801,N_146,N_318);
or U802 (N_802,N_243,N_432);
or U803 (N_803,N_161,N_559);
nand U804 (N_804,N_399,N_561);
nand U805 (N_805,N_348,N_214);
and U806 (N_806,N_361,N_334);
nor U807 (N_807,N_22,N_67);
and U808 (N_808,N_475,N_165);
or U809 (N_809,N_198,N_429);
nand U810 (N_810,N_295,N_496);
nand U811 (N_811,N_406,N_73);
or U812 (N_812,N_166,N_349);
or U813 (N_813,N_454,N_32);
or U814 (N_814,N_236,N_321);
nand U815 (N_815,N_58,N_241);
nand U816 (N_816,N_216,N_101);
and U817 (N_817,N_409,N_574);
nand U818 (N_818,N_227,N_587);
or U819 (N_819,N_83,N_538);
or U820 (N_820,N_504,N_200);
and U821 (N_821,N_286,N_120);
or U822 (N_822,N_512,N_233);
or U823 (N_823,N_524,N_181);
nor U824 (N_824,N_184,N_18);
and U825 (N_825,N_225,N_346);
or U826 (N_826,N_544,N_212);
and U827 (N_827,N_80,N_472);
nor U828 (N_828,N_172,N_489);
nand U829 (N_829,N_158,N_100);
nor U830 (N_830,N_362,N_134);
and U831 (N_831,N_506,N_12);
or U832 (N_832,N_145,N_108);
nand U833 (N_833,N_419,N_49);
and U834 (N_834,N_115,N_54);
nand U835 (N_835,N_179,N_259);
nand U836 (N_836,N_11,N_281);
or U837 (N_837,N_86,N_527);
or U838 (N_838,N_460,N_133);
or U839 (N_839,N_78,N_88);
and U840 (N_840,N_571,N_540);
and U841 (N_841,N_104,N_395);
nand U842 (N_842,N_70,N_289);
nor U843 (N_843,N_305,N_81);
and U844 (N_844,N_209,N_52);
nor U845 (N_845,N_92,N_3);
nor U846 (N_846,N_153,N_6);
nor U847 (N_847,N_109,N_522);
or U848 (N_848,N_0,N_590);
or U849 (N_849,N_366,N_301);
and U850 (N_850,N_168,N_344);
and U851 (N_851,N_494,N_400);
and U852 (N_852,N_75,N_164);
and U853 (N_853,N_355,N_206);
and U854 (N_854,N_63,N_226);
nand U855 (N_855,N_267,N_211);
or U856 (N_856,N_462,N_21);
xnor U857 (N_857,N_546,N_45);
nor U858 (N_858,N_195,N_266);
or U859 (N_859,N_405,N_427);
nor U860 (N_860,N_498,N_127);
nor U861 (N_861,N_111,N_383);
and U862 (N_862,N_37,N_2);
nor U863 (N_863,N_547,N_148);
and U864 (N_864,N_29,N_112);
nor U865 (N_865,N_356,N_36);
nor U866 (N_866,N_125,N_331);
nor U867 (N_867,N_474,N_282);
nand U868 (N_868,N_324,N_569);
nor U869 (N_869,N_592,N_309);
and U870 (N_870,N_593,N_280);
and U871 (N_871,N_551,N_370);
nor U872 (N_872,N_448,N_375);
nor U873 (N_873,N_87,N_377);
nor U874 (N_874,N_458,N_235);
nand U875 (N_875,N_347,N_237);
nor U876 (N_876,N_442,N_265);
or U877 (N_877,N_497,N_534);
nand U878 (N_878,N_173,N_391);
nand U879 (N_879,N_253,N_531);
and U880 (N_880,N_553,N_48);
and U881 (N_881,N_388,N_341);
or U882 (N_882,N_414,N_277);
and U883 (N_883,N_434,N_523);
or U884 (N_884,N_339,N_480);
nand U885 (N_885,N_137,N_254);
or U886 (N_886,N_5,N_549);
and U887 (N_887,N_44,N_345);
nor U888 (N_888,N_257,N_162);
and U889 (N_889,N_470,N_578);
nand U890 (N_890,N_147,N_407);
or U891 (N_891,N_487,N_598);
nand U892 (N_892,N_110,N_307);
nor U893 (N_893,N_68,N_413);
nand U894 (N_894,N_381,N_176);
and U895 (N_895,N_584,N_440);
or U896 (N_896,N_431,N_479);
nor U897 (N_897,N_232,N_261);
or U898 (N_898,N_426,N_424);
nand U899 (N_899,N_418,N_372);
and U900 (N_900,N_303,N_2);
and U901 (N_901,N_445,N_580);
nand U902 (N_902,N_360,N_468);
xor U903 (N_903,N_163,N_35);
nor U904 (N_904,N_315,N_384);
and U905 (N_905,N_436,N_484);
or U906 (N_906,N_272,N_200);
xnor U907 (N_907,N_126,N_339);
nand U908 (N_908,N_396,N_588);
nand U909 (N_909,N_19,N_365);
nand U910 (N_910,N_126,N_91);
or U911 (N_911,N_507,N_417);
nand U912 (N_912,N_108,N_334);
and U913 (N_913,N_130,N_256);
nand U914 (N_914,N_81,N_595);
and U915 (N_915,N_411,N_433);
xnor U916 (N_916,N_35,N_464);
nand U917 (N_917,N_265,N_65);
and U918 (N_918,N_5,N_385);
nand U919 (N_919,N_149,N_269);
nor U920 (N_920,N_37,N_266);
or U921 (N_921,N_448,N_402);
nor U922 (N_922,N_406,N_554);
nor U923 (N_923,N_594,N_78);
nand U924 (N_924,N_386,N_498);
nor U925 (N_925,N_463,N_202);
or U926 (N_926,N_225,N_330);
and U927 (N_927,N_471,N_451);
nand U928 (N_928,N_327,N_491);
nor U929 (N_929,N_109,N_17);
and U930 (N_930,N_17,N_400);
nand U931 (N_931,N_351,N_536);
and U932 (N_932,N_258,N_219);
nor U933 (N_933,N_508,N_306);
nand U934 (N_934,N_14,N_284);
nand U935 (N_935,N_339,N_224);
nor U936 (N_936,N_359,N_573);
or U937 (N_937,N_48,N_23);
nand U938 (N_938,N_104,N_130);
nand U939 (N_939,N_243,N_427);
nor U940 (N_940,N_520,N_42);
and U941 (N_941,N_365,N_107);
and U942 (N_942,N_199,N_320);
nor U943 (N_943,N_495,N_295);
nor U944 (N_944,N_241,N_306);
nand U945 (N_945,N_245,N_579);
nor U946 (N_946,N_414,N_252);
or U947 (N_947,N_443,N_372);
nor U948 (N_948,N_586,N_470);
nand U949 (N_949,N_335,N_441);
and U950 (N_950,N_458,N_463);
nor U951 (N_951,N_440,N_513);
nand U952 (N_952,N_107,N_526);
nor U953 (N_953,N_237,N_222);
and U954 (N_954,N_59,N_192);
nor U955 (N_955,N_29,N_411);
nand U956 (N_956,N_148,N_244);
and U957 (N_957,N_473,N_256);
nand U958 (N_958,N_577,N_127);
or U959 (N_959,N_261,N_7);
nor U960 (N_960,N_277,N_587);
nor U961 (N_961,N_554,N_169);
and U962 (N_962,N_2,N_281);
or U963 (N_963,N_425,N_489);
nand U964 (N_964,N_218,N_372);
nor U965 (N_965,N_482,N_549);
and U966 (N_966,N_130,N_593);
or U967 (N_967,N_143,N_564);
nand U968 (N_968,N_88,N_105);
and U969 (N_969,N_476,N_349);
or U970 (N_970,N_526,N_48);
xnor U971 (N_971,N_91,N_581);
and U972 (N_972,N_598,N_399);
nand U973 (N_973,N_548,N_257);
or U974 (N_974,N_152,N_195);
xnor U975 (N_975,N_426,N_242);
nor U976 (N_976,N_424,N_1);
or U977 (N_977,N_467,N_272);
or U978 (N_978,N_519,N_284);
nor U979 (N_979,N_139,N_259);
nor U980 (N_980,N_412,N_36);
nand U981 (N_981,N_171,N_422);
nor U982 (N_982,N_149,N_584);
and U983 (N_983,N_68,N_71);
or U984 (N_984,N_478,N_288);
nor U985 (N_985,N_196,N_237);
or U986 (N_986,N_402,N_268);
nand U987 (N_987,N_168,N_146);
nand U988 (N_988,N_75,N_112);
nor U989 (N_989,N_287,N_463);
nor U990 (N_990,N_43,N_565);
and U991 (N_991,N_596,N_93);
or U992 (N_992,N_2,N_570);
nand U993 (N_993,N_177,N_308);
or U994 (N_994,N_140,N_59);
nor U995 (N_995,N_151,N_234);
nor U996 (N_996,N_322,N_271);
and U997 (N_997,N_500,N_175);
nor U998 (N_998,N_22,N_96);
nor U999 (N_999,N_191,N_455);
nand U1000 (N_1000,N_178,N_506);
and U1001 (N_1001,N_262,N_324);
nand U1002 (N_1002,N_171,N_423);
and U1003 (N_1003,N_374,N_321);
and U1004 (N_1004,N_306,N_533);
nand U1005 (N_1005,N_341,N_303);
or U1006 (N_1006,N_478,N_251);
and U1007 (N_1007,N_224,N_256);
nand U1008 (N_1008,N_596,N_396);
nor U1009 (N_1009,N_197,N_591);
nand U1010 (N_1010,N_157,N_410);
or U1011 (N_1011,N_262,N_309);
and U1012 (N_1012,N_171,N_122);
and U1013 (N_1013,N_24,N_145);
or U1014 (N_1014,N_164,N_346);
nand U1015 (N_1015,N_76,N_329);
and U1016 (N_1016,N_71,N_111);
and U1017 (N_1017,N_56,N_162);
nand U1018 (N_1018,N_516,N_99);
nand U1019 (N_1019,N_5,N_541);
and U1020 (N_1020,N_397,N_411);
and U1021 (N_1021,N_541,N_500);
nand U1022 (N_1022,N_41,N_140);
and U1023 (N_1023,N_289,N_0);
nor U1024 (N_1024,N_168,N_508);
nor U1025 (N_1025,N_231,N_225);
nand U1026 (N_1026,N_6,N_557);
nor U1027 (N_1027,N_22,N_135);
and U1028 (N_1028,N_317,N_248);
nor U1029 (N_1029,N_13,N_97);
or U1030 (N_1030,N_57,N_586);
nand U1031 (N_1031,N_234,N_20);
nor U1032 (N_1032,N_542,N_550);
or U1033 (N_1033,N_202,N_51);
nor U1034 (N_1034,N_401,N_23);
and U1035 (N_1035,N_191,N_76);
nor U1036 (N_1036,N_432,N_543);
or U1037 (N_1037,N_323,N_488);
nand U1038 (N_1038,N_585,N_456);
nand U1039 (N_1039,N_254,N_316);
nor U1040 (N_1040,N_199,N_140);
and U1041 (N_1041,N_134,N_136);
nand U1042 (N_1042,N_245,N_425);
nand U1043 (N_1043,N_97,N_74);
nor U1044 (N_1044,N_421,N_580);
nor U1045 (N_1045,N_380,N_568);
and U1046 (N_1046,N_545,N_142);
nor U1047 (N_1047,N_120,N_455);
and U1048 (N_1048,N_378,N_554);
nand U1049 (N_1049,N_249,N_472);
nand U1050 (N_1050,N_280,N_300);
nor U1051 (N_1051,N_310,N_55);
or U1052 (N_1052,N_467,N_351);
or U1053 (N_1053,N_403,N_42);
nor U1054 (N_1054,N_105,N_431);
or U1055 (N_1055,N_521,N_106);
nor U1056 (N_1056,N_544,N_452);
or U1057 (N_1057,N_438,N_206);
and U1058 (N_1058,N_484,N_162);
and U1059 (N_1059,N_541,N_64);
nand U1060 (N_1060,N_563,N_569);
nor U1061 (N_1061,N_276,N_400);
and U1062 (N_1062,N_216,N_27);
and U1063 (N_1063,N_89,N_54);
and U1064 (N_1064,N_36,N_147);
and U1065 (N_1065,N_393,N_293);
or U1066 (N_1066,N_504,N_255);
nand U1067 (N_1067,N_140,N_314);
or U1068 (N_1068,N_172,N_310);
nand U1069 (N_1069,N_393,N_290);
or U1070 (N_1070,N_529,N_25);
and U1071 (N_1071,N_197,N_490);
or U1072 (N_1072,N_309,N_236);
or U1073 (N_1073,N_221,N_509);
nor U1074 (N_1074,N_506,N_268);
nand U1075 (N_1075,N_370,N_114);
nor U1076 (N_1076,N_103,N_434);
or U1077 (N_1077,N_587,N_426);
or U1078 (N_1078,N_19,N_518);
nor U1079 (N_1079,N_83,N_397);
or U1080 (N_1080,N_366,N_199);
or U1081 (N_1081,N_482,N_312);
or U1082 (N_1082,N_432,N_422);
nor U1083 (N_1083,N_463,N_393);
or U1084 (N_1084,N_75,N_570);
and U1085 (N_1085,N_285,N_172);
or U1086 (N_1086,N_143,N_361);
nand U1087 (N_1087,N_426,N_122);
nand U1088 (N_1088,N_189,N_550);
nor U1089 (N_1089,N_306,N_257);
or U1090 (N_1090,N_76,N_503);
nand U1091 (N_1091,N_211,N_119);
nand U1092 (N_1092,N_133,N_356);
nand U1093 (N_1093,N_307,N_239);
and U1094 (N_1094,N_156,N_343);
and U1095 (N_1095,N_237,N_303);
nor U1096 (N_1096,N_303,N_55);
and U1097 (N_1097,N_252,N_437);
or U1098 (N_1098,N_395,N_116);
nand U1099 (N_1099,N_241,N_296);
nand U1100 (N_1100,N_31,N_360);
xnor U1101 (N_1101,N_313,N_102);
nand U1102 (N_1102,N_206,N_389);
and U1103 (N_1103,N_416,N_557);
and U1104 (N_1104,N_346,N_209);
nand U1105 (N_1105,N_329,N_214);
nor U1106 (N_1106,N_498,N_63);
or U1107 (N_1107,N_244,N_431);
or U1108 (N_1108,N_284,N_5);
nor U1109 (N_1109,N_150,N_216);
and U1110 (N_1110,N_298,N_523);
nor U1111 (N_1111,N_329,N_479);
nor U1112 (N_1112,N_348,N_202);
xor U1113 (N_1113,N_509,N_417);
or U1114 (N_1114,N_372,N_390);
nand U1115 (N_1115,N_320,N_111);
nand U1116 (N_1116,N_10,N_42);
nor U1117 (N_1117,N_585,N_355);
or U1118 (N_1118,N_15,N_470);
nand U1119 (N_1119,N_468,N_460);
nand U1120 (N_1120,N_31,N_89);
or U1121 (N_1121,N_548,N_230);
nand U1122 (N_1122,N_368,N_291);
nand U1123 (N_1123,N_331,N_439);
nand U1124 (N_1124,N_247,N_395);
nor U1125 (N_1125,N_238,N_17);
and U1126 (N_1126,N_449,N_525);
nand U1127 (N_1127,N_287,N_281);
nand U1128 (N_1128,N_264,N_270);
nand U1129 (N_1129,N_25,N_435);
nand U1130 (N_1130,N_245,N_318);
or U1131 (N_1131,N_193,N_488);
nand U1132 (N_1132,N_220,N_479);
nand U1133 (N_1133,N_249,N_499);
and U1134 (N_1134,N_329,N_465);
and U1135 (N_1135,N_226,N_585);
nand U1136 (N_1136,N_568,N_159);
nor U1137 (N_1137,N_327,N_524);
nor U1138 (N_1138,N_130,N_265);
and U1139 (N_1139,N_193,N_333);
nor U1140 (N_1140,N_446,N_265);
and U1141 (N_1141,N_71,N_545);
nand U1142 (N_1142,N_368,N_197);
or U1143 (N_1143,N_14,N_229);
xor U1144 (N_1144,N_428,N_475);
and U1145 (N_1145,N_149,N_188);
and U1146 (N_1146,N_84,N_472);
or U1147 (N_1147,N_404,N_108);
and U1148 (N_1148,N_32,N_299);
nor U1149 (N_1149,N_269,N_507);
nor U1150 (N_1150,N_28,N_477);
and U1151 (N_1151,N_323,N_75);
or U1152 (N_1152,N_223,N_25);
or U1153 (N_1153,N_157,N_118);
and U1154 (N_1154,N_5,N_60);
nor U1155 (N_1155,N_194,N_158);
nand U1156 (N_1156,N_526,N_411);
and U1157 (N_1157,N_551,N_52);
nand U1158 (N_1158,N_525,N_133);
and U1159 (N_1159,N_108,N_32);
or U1160 (N_1160,N_308,N_305);
nor U1161 (N_1161,N_111,N_488);
or U1162 (N_1162,N_327,N_163);
or U1163 (N_1163,N_35,N_593);
or U1164 (N_1164,N_560,N_177);
nor U1165 (N_1165,N_339,N_508);
nor U1166 (N_1166,N_419,N_563);
or U1167 (N_1167,N_423,N_568);
and U1168 (N_1168,N_119,N_354);
or U1169 (N_1169,N_530,N_111);
or U1170 (N_1170,N_243,N_493);
nor U1171 (N_1171,N_151,N_273);
nor U1172 (N_1172,N_532,N_397);
or U1173 (N_1173,N_16,N_475);
and U1174 (N_1174,N_172,N_594);
nor U1175 (N_1175,N_519,N_15);
nand U1176 (N_1176,N_100,N_125);
or U1177 (N_1177,N_466,N_253);
or U1178 (N_1178,N_476,N_141);
and U1179 (N_1179,N_505,N_288);
nand U1180 (N_1180,N_73,N_525);
and U1181 (N_1181,N_598,N_18);
nor U1182 (N_1182,N_495,N_569);
or U1183 (N_1183,N_240,N_224);
nand U1184 (N_1184,N_331,N_491);
nor U1185 (N_1185,N_471,N_525);
nor U1186 (N_1186,N_193,N_344);
or U1187 (N_1187,N_439,N_343);
nor U1188 (N_1188,N_285,N_349);
nor U1189 (N_1189,N_499,N_541);
nand U1190 (N_1190,N_60,N_451);
nand U1191 (N_1191,N_254,N_85);
nor U1192 (N_1192,N_388,N_549);
and U1193 (N_1193,N_209,N_115);
and U1194 (N_1194,N_145,N_289);
and U1195 (N_1195,N_40,N_194);
and U1196 (N_1196,N_477,N_597);
nor U1197 (N_1197,N_441,N_578);
and U1198 (N_1198,N_110,N_77);
or U1199 (N_1199,N_218,N_360);
nor U1200 (N_1200,N_908,N_672);
nor U1201 (N_1201,N_718,N_1077);
nand U1202 (N_1202,N_1185,N_1093);
nor U1203 (N_1203,N_889,N_1101);
and U1204 (N_1204,N_902,N_639);
nor U1205 (N_1205,N_1021,N_755);
nor U1206 (N_1206,N_1156,N_1134);
and U1207 (N_1207,N_995,N_1023);
nand U1208 (N_1208,N_967,N_1102);
nor U1209 (N_1209,N_1193,N_1033);
nor U1210 (N_1210,N_609,N_957);
nor U1211 (N_1211,N_863,N_694);
nand U1212 (N_1212,N_941,N_797);
or U1213 (N_1213,N_956,N_666);
xor U1214 (N_1214,N_775,N_971);
and U1215 (N_1215,N_799,N_1196);
nor U1216 (N_1216,N_859,N_1012);
nor U1217 (N_1217,N_1135,N_1067);
nand U1218 (N_1218,N_1079,N_1031);
and U1219 (N_1219,N_879,N_1032);
or U1220 (N_1220,N_660,N_691);
nand U1221 (N_1221,N_959,N_838);
nor U1222 (N_1222,N_1174,N_835);
nand U1223 (N_1223,N_1051,N_638);
or U1224 (N_1224,N_826,N_876);
nand U1225 (N_1225,N_686,N_1087);
and U1226 (N_1226,N_724,N_630);
or U1227 (N_1227,N_720,N_669);
nand U1228 (N_1228,N_858,N_896);
nor U1229 (N_1229,N_1078,N_920);
and U1230 (N_1230,N_823,N_973);
nand U1231 (N_1231,N_1131,N_1030);
or U1232 (N_1232,N_703,N_757);
nor U1233 (N_1233,N_642,N_831);
nand U1234 (N_1234,N_647,N_1133);
and U1235 (N_1235,N_1144,N_680);
or U1236 (N_1236,N_994,N_982);
and U1237 (N_1237,N_1153,N_1029);
or U1238 (N_1238,N_751,N_731);
and U1239 (N_1239,N_878,N_1019);
and U1240 (N_1240,N_1114,N_884);
nand U1241 (N_1241,N_1167,N_911);
and U1242 (N_1242,N_632,N_766);
nand U1243 (N_1243,N_1122,N_1076);
nand U1244 (N_1244,N_1084,N_899);
xnor U1245 (N_1245,N_1081,N_933);
nor U1246 (N_1246,N_948,N_931);
nand U1247 (N_1247,N_937,N_1117);
or U1248 (N_1248,N_641,N_1178);
or U1249 (N_1249,N_1177,N_992);
nand U1250 (N_1250,N_893,N_1095);
nand U1251 (N_1251,N_998,N_1001);
nor U1252 (N_1252,N_830,N_781);
xnor U1253 (N_1253,N_617,N_658);
nand U1254 (N_1254,N_778,N_722);
or U1255 (N_1255,N_942,N_1128);
nor U1256 (N_1256,N_1037,N_1161);
and U1257 (N_1257,N_1020,N_739);
nor U1258 (N_1258,N_880,N_1042);
or U1259 (N_1259,N_1017,N_1013);
and U1260 (N_1260,N_1108,N_843);
and U1261 (N_1261,N_626,N_704);
nor U1262 (N_1262,N_729,N_980);
or U1263 (N_1263,N_857,N_986);
and U1264 (N_1264,N_954,N_825);
and U1265 (N_1265,N_758,N_1034);
or U1266 (N_1266,N_610,N_763);
or U1267 (N_1267,N_1035,N_1024);
or U1268 (N_1268,N_1136,N_780);
nand U1269 (N_1269,N_1151,N_900);
and U1270 (N_1270,N_915,N_795);
and U1271 (N_1271,N_719,N_1058);
nor U1272 (N_1272,N_1073,N_892);
or U1273 (N_1273,N_1062,N_921);
nand U1274 (N_1274,N_983,N_634);
and U1275 (N_1275,N_1104,N_807);
nor U1276 (N_1276,N_916,N_675);
nor U1277 (N_1277,N_640,N_978);
or U1278 (N_1278,N_1119,N_635);
or U1279 (N_1279,N_949,N_1146);
nor U1280 (N_1280,N_913,N_988);
and U1281 (N_1281,N_1159,N_1008);
nand U1282 (N_1282,N_1063,N_645);
nand U1283 (N_1283,N_1150,N_714);
xor U1284 (N_1284,N_1006,N_800);
nor U1285 (N_1285,N_699,N_733);
or U1286 (N_1286,N_721,N_681);
or U1287 (N_1287,N_782,N_1145);
nor U1288 (N_1288,N_656,N_1155);
or U1289 (N_1289,N_636,N_643);
or U1290 (N_1290,N_732,N_1057);
nand U1291 (N_1291,N_919,N_926);
nor U1292 (N_1292,N_796,N_760);
nand U1293 (N_1293,N_845,N_793);
nand U1294 (N_1294,N_1169,N_813);
nand U1295 (N_1295,N_789,N_667);
nor U1296 (N_1296,N_670,N_708);
and U1297 (N_1297,N_1036,N_1115);
nand U1298 (N_1298,N_1074,N_770);
nand U1299 (N_1299,N_690,N_1061);
nand U1300 (N_1300,N_1045,N_1195);
or U1301 (N_1301,N_673,N_717);
and U1302 (N_1302,N_895,N_907);
nor U1303 (N_1303,N_692,N_882);
nor U1304 (N_1304,N_827,N_804);
nor U1305 (N_1305,N_1164,N_996);
xnor U1306 (N_1306,N_687,N_776);
and U1307 (N_1307,N_1168,N_898);
or U1308 (N_1308,N_984,N_897);
or U1309 (N_1309,N_657,N_1189);
and U1310 (N_1310,N_664,N_890);
and U1311 (N_1311,N_1147,N_702);
nor U1312 (N_1312,N_1184,N_1011);
and U1313 (N_1313,N_1171,N_820);
nand U1314 (N_1314,N_1130,N_964);
nor U1315 (N_1315,N_874,N_1197);
nor U1316 (N_1316,N_1094,N_1086);
or U1317 (N_1317,N_761,N_1047);
nor U1318 (N_1318,N_979,N_794);
nor U1319 (N_1319,N_904,N_842);
nor U1320 (N_1320,N_1052,N_1046);
nand U1321 (N_1321,N_628,N_940);
or U1322 (N_1322,N_841,N_1091);
nand U1323 (N_1323,N_754,N_625);
and U1324 (N_1324,N_762,N_999);
nand U1325 (N_1325,N_1187,N_867);
or U1326 (N_1326,N_706,N_816);
and U1327 (N_1327,N_1009,N_950);
nand U1328 (N_1328,N_749,N_834);
and U1329 (N_1329,N_737,N_932);
nor U1330 (N_1330,N_1106,N_912);
nand U1331 (N_1331,N_611,N_847);
and U1332 (N_1332,N_1148,N_877);
and U1333 (N_1333,N_1142,N_872);
nand U1334 (N_1334,N_786,N_946);
and U1335 (N_1335,N_844,N_1129);
nor U1336 (N_1336,N_987,N_1066);
and U1337 (N_1337,N_990,N_1089);
nor U1338 (N_1338,N_738,N_1099);
nand U1339 (N_1339,N_934,N_1048);
nor U1340 (N_1340,N_849,N_1162);
or U1341 (N_1341,N_1010,N_852);
nor U1342 (N_1342,N_1107,N_759);
and U1343 (N_1343,N_1172,N_871);
nand U1344 (N_1344,N_792,N_1085);
nor U1345 (N_1345,N_616,N_752);
and U1346 (N_1346,N_1025,N_1163);
and U1347 (N_1347,N_618,N_608);
or U1348 (N_1348,N_685,N_707);
nor U1349 (N_1349,N_828,N_661);
nand U1350 (N_1350,N_1072,N_651);
nand U1351 (N_1351,N_928,N_869);
nand U1352 (N_1352,N_765,N_637);
or U1353 (N_1353,N_993,N_972);
and U1354 (N_1354,N_976,N_1180);
nor U1355 (N_1355,N_866,N_1103);
nor U1356 (N_1356,N_1109,N_802);
nand U1357 (N_1357,N_945,N_1040);
xnor U1358 (N_1358,N_1199,N_710);
or U1359 (N_1359,N_1152,N_909);
or U1360 (N_1360,N_1140,N_1186);
and U1361 (N_1361,N_850,N_822);
or U1362 (N_1362,N_924,N_679);
or U1363 (N_1363,N_832,N_963);
nand U1364 (N_1364,N_929,N_1138);
or U1365 (N_1365,N_772,N_1139);
and U1366 (N_1366,N_1158,N_1132);
or U1367 (N_1367,N_1088,N_712);
nor U1368 (N_1368,N_701,N_974);
nor U1369 (N_1369,N_705,N_1166);
nand U1370 (N_1370,N_1065,N_1126);
or U1371 (N_1371,N_955,N_709);
nand U1372 (N_1372,N_854,N_684);
nand U1373 (N_1373,N_756,N_966);
and U1374 (N_1374,N_1041,N_881);
and U1375 (N_1375,N_695,N_734);
nand U1376 (N_1376,N_649,N_894);
and U1377 (N_1377,N_633,N_862);
or U1378 (N_1378,N_1082,N_981);
or U1379 (N_1379,N_612,N_989);
nor U1380 (N_1380,N_1149,N_870);
and U1381 (N_1381,N_1005,N_747);
nand U1382 (N_1382,N_905,N_698);
and U1383 (N_1383,N_774,N_1069);
nor U1384 (N_1384,N_677,N_935);
or U1385 (N_1385,N_1022,N_764);
or U1386 (N_1386,N_619,N_997);
nor U1387 (N_1387,N_696,N_1050);
or U1388 (N_1388,N_991,N_1026);
or U1389 (N_1389,N_925,N_650);
nand U1390 (N_1390,N_1190,N_1179);
and U1391 (N_1391,N_644,N_740);
and U1392 (N_1392,N_829,N_906);
nand U1393 (N_1393,N_631,N_953);
or U1394 (N_1394,N_605,N_812);
and U1395 (N_1395,N_1124,N_1173);
and U1396 (N_1396,N_746,N_1125);
or U1397 (N_1397,N_910,N_663);
nand U1398 (N_1398,N_697,N_1118);
and U1399 (N_1399,N_1143,N_629);
nand U1400 (N_1400,N_1110,N_723);
or U1401 (N_1401,N_1004,N_744);
nor U1402 (N_1402,N_965,N_865);
nor U1403 (N_1403,N_1038,N_1055);
or U1404 (N_1404,N_700,N_676);
nor U1405 (N_1405,N_961,N_603);
or U1406 (N_1406,N_741,N_736);
or U1407 (N_1407,N_969,N_839);
nand U1408 (N_1408,N_840,N_769);
nor U1409 (N_1409,N_1183,N_665);
or U1410 (N_1410,N_1014,N_1027);
nor U1411 (N_1411,N_668,N_883);
and U1412 (N_1412,N_604,N_1015);
and U1413 (N_1413,N_1121,N_1068);
nor U1414 (N_1414,N_715,N_1141);
or U1415 (N_1415,N_622,N_1056);
xor U1416 (N_1416,N_1176,N_1096);
nand U1417 (N_1417,N_817,N_623);
nor U1418 (N_1418,N_1043,N_1002);
or U1419 (N_1419,N_726,N_671);
nand U1420 (N_1420,N_951,N_975);
and U1421 (N_1421,N_788,N_803);
nor U1422 (N_1422,N_683,N_1154);
and U1423 (N_1423,N_868,N_783);
and U1424 (N_1424,N_1007,N_1112);
and U1425 (N_1425,N_1060,N_1105);
nand U1426 (N_1426,N_798,N_1097);
nor U1427 (N_1427,N_1044,N_748);
nand U1428 (N_1428,N_960,N_624);
or U1429 (N_1429,N_922,N_943);
and U1430 (N_1430,N_837,N_962);
nor U1431 (N_1431,N_627,N_923);
and U1432 (N_1432,N_1198,N_903);
and U1433 (N_1433,N_735,N_1080);
nor U1434 (N_1434,N_856,N_725);
nand U1435 (N_1435,N_1000,N_716);
and U1436 (N_1436,N_1192,N_654);
and U1437 (N_1437,N_1083,N_674);
and U1438 (N_1438,N_601,N_659);
and U1439 (N_1439,N_713,N_1028);
and U1440 (N_1440,N_891,N_918);
and U1441 (N_1441,N_768,N_753);
nand U1442 (N_1442,N_767,N_930);
and U1443 (N_1443,N_1182,N_824);
nand U1444 (N_1444,N_648,N_806);
and U1445 (N_1445,N_688,N_833);
or U1446 (N_1446,N_809,N_864);
nor U1447 (N_1447,N_655,N_1175);
or U1448 (N_1448,N_888,N_801);
or U1449 (N_1449,N_1016,N_808);
nor U1450 (N_1450,N_1160,N_1137);
nand U1451 (N_1451,N_901,N_821);
nor U1452 (N_1452,N_607,N_711);
nor U1453 (N_1453,N_1188,N_958);
nor U1454 (N_1454,N_1071,N_678);
and U1455 (N_1455,N_970,N_1092);
nand U1456 (N_1456,N_936,N_771);
and U1457 (N_1457,N_653,N_791);
nor U1458 (N_1458,N_1075,N_728);
and U1459 (N_1459,N_621,N_861);
nand U1460 (N_1460,N_952,N_1098);
and U1461 (N_1461,N_811,N_853);
or U1462 (N_1462,N_836,N_620);
nand U1463 (N_1463,N_927,N_745);
nand U1464 (N_1464,N_875,N_1157);
and U1465 (N_1465,N_848,N_815);
nand U1466 (N_1466,N_846,N_1194);
and U1467 (N_1467,N_939,N_682);
and U1468 (N_1468,N_1165,N_790);
or U1469 (N_1469,N_1170,N_1049);
nor U1470 (N_1470,N_1018,N_947);
nand U1471 (N_1471,N_968,N_602);
nand U1472 (N_1472,N_606,N_1064);
and U1473 (N_1473,N_693,N_1127);
or U1474 (N_1474,N_662,N_646);
or U1475 (N_1475,N_750,N_614);
nand U1476 (N_1476,N_819,N_785);
and U1477 (N_1477,N_773,N_917);
or U1478 (N_1478,N_600,N_887);
nor U1479 (N_1479,N_652,N_977);
or U1480 (N_1480,N_886,N_1039);
and U1481 (N_1481,N_860,N_851);
nand U1482 (N_1482,N_787,N_1090);
nor U1483 (N_1483,N_615,N_1054);
or U1484 (N_1484,N_1123,N_743);
nand U1485 (N_1485,N_805,N_613);
and U1486 (N_1486,N_914,N_1070);
or U1487 (N_1487,N_944,N_742);
nand U1488 (N_1488,N_1120,N_1116);
xnor U1489 (N_1489,N_689,N_1113);
and U1490 (N_1490,N_1181,N_855);
nand U1491 (N_1491,N_810,N_938);
nand U1492 (N_1492,N_784,N_1191);
nor U1493 (N_1493,N_985,N_779);
nand U1494 (N_1494,N_1059,N_777);
or U1495 (N_1495,N_1100,N_873);
nand U1496 (N_1496,N_885,N_1111);
nor U1497 (N_1497,N_818,N_814);
and U1498 (N_1498,N_1003,N_730);
or U1499 (N_1499,N_727,N_1053);
and U1500 (N_1500,N_1016,N_1198);
nor U1501 (N_1501,N_817,N_811);
nor U1502 (N_1502,N_1177,N_725);
and U1503 (N_1503,N_773,N_737);
and U1504 (N_1504,N_1018,N_698);
and U1505 (N_1505,N_1187,N_1075);
and U1506 (N_1506,N_966,N_905);
and U1507 (N_1507,N_1057,N_1027);
and U1508 (N_1508,N_756,N_1170);
and U1509 (N_1509,N_773,N_911);
nor U1510 (N_1510,N_814,N_906);
and U1511 (N_1511,N_997,N_1070);
and U1512 (N_1512,N_1192,N_676);
xor U1513 (N_1513,N_609,N_897);
and U1514 (N_1514,N_1136,N_697);
and U1515 (N_1515,N_909,N_955);
and U1516 (N_1516,N_749,N_939);
nand U1517 (N_1517,N_1005,N_1070);
nor U1518 (N_1518,N_1150,N_853);
nand U1519 (N_1519,N_931,N_1101);
nor U1520 (N_1520,N_714,N_948);
and U1521 (N_1521,N_704,N_603);
nand U1522 (N_1522,N_1085,N_1061);
and U1523 (N_1523,N_1167,N_627);
or U1524 (N_1524,N_871,N_1088);
and U1525 (N_1525,N_626,N_743);
and U1526 (N_1526,N_1109,N_1082);
nand U1527 (N_1527,N_609,N_621);
or U1528 (N_1528,N_873,N_740);
and U1529 (N_1529,N_827,N_777);
nand U1530 (N_1530,N_806,N_856);
nand U1531 (N_1531,N_993,N_1082);
xnor U1532 (N_1532,N_1105,N_1089);
nor U1533 (N_1533,N_979,N_1089);
or U1534 (N_1534,N_834,N_1028);
nand U1535 (N_1535,N_1000,N_956);
nor U1536 (N_1536,N_915,N_764);
and U1537 (N_1537,N_830,N_625);
nand U1538 (N_1538,N_749,N_1125);
nand U1539 (N_1539,N_993,N_840);
or U1540 (N_1540,N_1071,N_648);
nand U1541 (N_1541,N_957,N_690);
nand U1542 (N_1542,N_1194,N_957);
nand U1543 (N_1543,N_860,N_713);
nor U1544 (N_1544,N_1151,N_676);
or U1545 (N_1545,N_1065,N_1036);
and U1546 (N_1546,N_712,N_1065);
nor U1547 (N_1547,N_830,N_853);
nor U1548 (N_1548,N_701,N_1055);
nor U1549 (N_1549,N_1139,N_1182);
nor U1550 (N_1550,N_681,N_612);
nand U1551 (N_1551,N_786,N_1006);
nand U1552 (N_1552,N_1017,N_1125);
nand U1553 (N_1553,N_1071,N_977);
nand U1554 (N_1554,N_748,N_755);
and U1555 (N_1555,N_1119,N_1140);
and U1556 (N_1556,N_641,N_921);
or U1557 (N_1557,N_1080,N_1083);
nand U1558 (N_1558,N_1125,N_825);
and U1559 (N_1559,N_865,N_660);
and U1560 (N_1560,N_1127,N_1004);
nor U1561 (N_1561,N_1119,N_799);
xor U1562 (N_1562,N_1164,N_664);
nor U1563 (N_1563,N_1157,N_1070);
and U1564 (N_1564,N_730,N_1172);
nor U1565 (N_1565,N_774,N_1033);
and U1566 (N_1566,N_1108,N_1102);
nand U1567 (N_1567,N_684,N_835);
nor U1568 (N_1568,N_644,N_743);
or U1569 (N_1569,N_1001,N_822);
nand U1570 (N_1570,N_839,N_1162);
and U1571 (N_1571,N_926,N_971);
or U1572 (N_1572,N_745,N_1068);
or U1573 (N_1573,N_1190,N_1145);
nand U1574 (N_1574,N_1055,N_1026);
or U1575 (N_1575,N_812,N_1180);
and U1576 (N_1576,N_1024,N_905);
nor U1577 (N_1577,N_987,N_1157);
nand U1578 (N_1578,N_1172,N_963);
nand U1579 (N_1579,N_892,N_698);
or U1580 (N_1580,N_709,N_604);
and U1581 (N_1581,N_851,N_974);
or U1582 (N_1582,N_711,N_728);
nor U1583 (N_1583,N_1116,N_1103);
nor U1584 (N_1584,N_917,N_953);
nor U1585 (N_1585,N_1076,N_878);
nand U1586 (N_1586,N_1164,N_793);
nand U1587 (N_1587,N_869,N_1180);
and U1588 (N_1588,N_735,N_1006);
nor U1589 (N_1589,N_850,N_983);
nor U1590 (N_1590,N_845,N_1113);
or U1591 (N_1591,N_651,N_825);
or U1592 (N_1592,N_1092,N_871);
nand U1593 (N_1593,N_896,N_922);
nand U1594 (N_1594,N_1062,N_648);
nand U1595 (N_1595,N_883,N_1162);
and U1596 (N_1596,N_1101,N_934);
or U1597 (N_1597,N_1190,N_861);
and U1598 (N_1598,N_1165,N_681);
nand U1599 (N_1599,N_876,N_1061);
nand U1600 (N_1600,N_1148,N_969);
or U1601 (N_1601,N_1140,N_1035);
nor U1602 (N_1602,N_1118,N_1049);
xor U1603 (N_1603,N_631,N_742);
nor U1604 (N_1604,N_944,N_706);
nor U1605 (N_1605,N_801,N_610);
or U1606 (N_1606,N_1064,N_727);
nor U1607 (N_1607,N_795,N_657);
and U1608 (N_1608,N_620,N_754);
nor U1609 (N_1609,N_795,N_1197);
and U1610 (N_1610,N_952,N_767);
nand U1611 (N_1611,N_741,N_645);
nand U1612 (N_1612,N_1007,N_1127);
nand U1613 (N_1613,N_983,N_1101);
and U1614 (N_1614,N_688,N_1169);
nor U1615 (N_1615,N_718,N_1064);
or U1616 (N_1616,N_873,N_1103);
and U1617 (N_1617,N_930,N_757);
xor U1618 (N_1618,N_1042,N_688);
or U1619 (N_1619,N_753,N_878);
nor U1620 (N_1620,N_924,N_931);
and U1621 (N_1621,N_820,N_934);
nor U1622 (N_1622,N_994,N_1160);
and U1623 (N_1623,N_851,N_1083);
or U1624 (N_1624,N_1193,N_1157);
nor U1625 (N_1625,N_799,N_861);
nor U1626 (N_1626,N_779,N_782);
nand U1627 (N_1627,N_668,N_889);
nor U1628 (N_1628,N_1053,N_998);
nand U1629 (N_1629,N_1097,N_785);
nand U1630 (N_1630,N_826,N_763);
or U1631 (N_1631,N_986,N_879);
nor U1632 (N_1632,N_807,N_1141);
nor U1633 (N_1633,N_1058,N_690);
or U1634 (N_1634,N_1029,N_1146);
nand U1635 (N_1635,N_642,N_932);
and U1636 (N_1636,N_996,N_964);
or U1637 (N_1637,N_632,N_925);
and U1638 (N_1638,N_1091,N_893);
and U1639 (N_1639,N_1145,N_707);
or U1640 (N_1640,N_834,N_632);
nand U1641 (N_1641,N_1172,N_673);
and U1642 (N_1642,N_978,N_653);
or U1643 (N_1643,N_623,N_704);
and U1644 (N_1644,N_907,N_1007);
or U1645 (N_1645,N_717,N_982);
xor U1646 (N_1646,N_681,N_1109);
or U1647 (N_1647,N_1190,N_722);
nor U1648 (N_1648,N_1078,N_668);
nor U1649 (N_1649,N_892,N_1039);
and U1650 (N_1650,N_736,N_1191);
or U1651 (N_1651,N_1006,N_768);
nor U1652 (N_1652,N_621,N_884);
or U1653 (N_1653,N_1154,N_941);
nor U1654 (N_1654,N_654,N_790);
nand U1655 (N_1655,N_766,N_1123);
nand U1656 (N_1656,N_977,N_1040);
and U1657 (N_1657,N_621,N_749);
xnor U1658 (N_1658,N_741,N_839);
or U1659 (N_1659,N_989,N_777);
nor U1660 (N_1660,N_744,N_834);
nor U1661 (N_1661,N_1171,N_1017);
nor U1662 (N_1662,N_715,N_865);
and U1663 (N_1663,N_975,N_701);
nor U1664 (N_1664,N_741,N_689);
or U1665 (N_1665,N_1081,N_1058);
and U1666 (N_1666,N_1131,N_1118);
nand U1667 (N_1667,N_753,N_1048);
or U1668 (N_1668,N_944,N_791);
or U1669 (N_1669,N_1027,N_1117);
nand U1670 (N_1670,N_920,N_1051);
nand U1671 (N_1671,N_1196,N_1092);
nor U1672 (N_1672,N_712,N_693);
nor U1673 (N_1673,N_1124,N_822);
and U1674 (N_1674,N_742,N_860);
xor U1675 (N_1675,N_699,N_1009);
and U1676 (N_1676,N_1066,N_762);
or U1677 (N_1677,N_1000,N_981);
nor U1678 (N_1678,N_1041,N_684);
nor U1679 (N_1679,N_650,N_982);
or U1680 (N_1680,N_946,N_1123);
nor U1681 (N_1681,N_1160,N_826);
and U1682 (N_1682,N_946,N_875);
xor U1683 (N_1683,N_1076,N_990);
nor U1684 (N_1684,N_716,N_707);
nor U1685 (N_1685,N_1156,N_946);
nor U1686 (N_1686,N_1164,N_997);
or U1687 (N_1687,N_803,N_1185);
and U1688 (N_1688,N_1172,N_1029);
nand U1689 (N_1689,N_949,N_1195);
nor U1690 (N_1690,N_653,N_825);
or U1691 (N_1691,N_979,N_641);
and U1692 (N_1692,N_950,N_888);
or U1693 (N_1693,N_684,N_682);
nand U1694 (N_1694,N_794,N_618);
or U1695 (N_1695,N_907,N_998);
and U1696 (N_1696,N_828,N_1104);
nand U1697 (N_1697,N_743,N_1175);
or U1698 (N_1698,N_959,N_714);
or U1699 (N_1699,N_774,N_909);
nor U1700 (N_1700,N_851,N_915);
and U1701 (N_1701,N_758,N_981);
or U1702 (N_1702,N_1074,N_1159);
nor U1703 (N_1703,N_1092,N_696);
nand U1704 (N_1704,N_644,N_661);
and U1705 (N_1705,N_1016,N_1111);
nor U1706 (N_1706,N_750,N_882);
nor U1707 (N_1707,N_661,N_1026);
nor U1708 (N_1708,N_1112,N_1031);
nand U1709 (N_1709,N_1009,N_719);
and U1710 (N_1710,N_1107,N_677);
or U1711 (N_1711,N_763,N_701);
nor U1712 (N_1712,N_1157,N_1163);
and U1713 (N_1713,N_935,N_703);
and U1714 (N_1714,N_1010,N_1187);
nor U1715 (N_1715,N_777,N_996);
or U1716 (N_1716,N_1181,N_886);
or U1717 (N_1717,N_799,N_667);
nor U1718 (N_1718,N_690,N_782);
and U1719 (N_1719,N_1138,N_652);
or U1720 (N_1720,N_745,N_1076);
nor U1721 (N_1721,N_680,N_616);
nand U1722 (N_1722,N_857,N_818);
nor U1723 (N_1723,N_715,N_638);
nor U1724 (N_1724,N_835,N_896);
nor U1725 (N_1725,N_809,N_1019);
or U1726 (N_1726,N_938,N_1026);
and U1727 (N_1727,N_959,N_892);
or U1728 (N_1728,N_749,N_832);
or U1729 (N_1729,N_963,N_893);
nor U1730 (N_1730,N_1106,N_1190);
nor U1731 (N_1731,N_971,N_992);
and U1732 (N_1732,N_808,N_792);
or U1733 (N_1733,N_1017,N_1010);
or U1734 (N_1734,N_863,N_891);
or U1735 (N_1735,N_790,N_820);
nor U1736 (N_1736,N_924,N_601);
nand U1737 (N_1737,N_772,N_770);
or U1738 (N_1738,N_846,N_1078);
nand U1739 (N_1739,N_600,N_1190);
nand U1740 (N_1740,N_959,N_911);
nor U1741 (N_1741,N_654,N_697);
nand U1742 (N_1742,N_904,N_885);
or U1743 (N_1743,N_842,N_927);
nand U1744 (N_1744,N_603,N_831);
nand U1745 (N_1745,N_1111,N_900);
nor U1746 (N_1746,N_675,N_655);
and U1747 (N_1747,N_722,N_1194);
or U1748 (N_1748,N_812,N_1159);
or U1749 (N_1749,N_987,N_912);
or U1750 (N_1750,N_1119,N_823);
nand U1751 (N_1751,N_974,N_702);
and U1752 (N_1752,N_854,N_885);
nand U1753 (N_1753,N_866,N_851);
nor U1754 (N_1754,N_887,N_962);
xnor U1755 (N_1755,N_879,N_617);
nor U1756 (N_1756,N_709,N_693);
and U1757 (N_1757,N_1067,N_623);
nor U1758 (N_1758,N_1005,N_783);
nor U1759 (N_1759,N_682,N_651);
nand U1760 (N_1760,N_687,N_710);
and U1761 (N_1761,N_1042,N_771);
nor U1762 (N_1762,N_673,N_691);
xor U1763 (N_1763,N_941,N_1162);
nand U1764 (N_1764,N_780,N_1186);
nand U1765 (N_1765,N_921,N_1104);
or U1766 (N_1766,N_1120,N_876);
nor U1767 (N_1767,N_628,N_855);
nor U1768 (N_1768,N_1131,N_1188);
nor U1769 (N_1769,N_773,N_1051);
nand U1770 (N_1770,N_643,N_803);
nand U1771 (N_1771,N_1134,N_889);
nor U1772 (N_1772,N_1134,N_1192);
or U1773 (N_1773,N_767,N_1014);
nand U1774 (N_1774,N_977,N_896);
nor U1775 (N_1775,N_704,N_948);
nand U1776 (N_1776,N_886,N_978);
and U1777 (N_1777,N_673,N_936);
or U1778 (N_1778,N_947,N_712);
or U1779 (N_1779,N_1115,N_1042);
or U1780 (N_1780,N_772,N_848);
or U1781 (N_1781,N_915,N_991);
nor U1782 (N_1782,N_889,N_1123);
nand U1783 (N_1783,N_924,N_1058);
or U1784 (N_1784,N_1177,N_629);
nand U1785 (N_1785,N_978,N_804);
nand U1786 (N_1786,N_804,N_977);
nor U1787 (N_1787,N_1161,N_986);
xor U1788 (N_1788,N_918,N_1147);
nor U1789 (N_1789,N_1081,N_1169);
nor U1790 (N_1790,N_804,N_936);
nor U1791 (N_1791,N_764,N_615);
nor U1792 (N_1792,N_1175,N_1065);
or U1793 (N_1793,N_817,N_890);
and U1794 (N_1794,N_1046,N_830);
xnor U1795 (N_1795,N_817,N_1178);
and U1796 (N_1796,N_760,N_931);
or U1797 (N_1797,N_1157,N_1158);
or U1798 (N_1798,N_749,N_1140);
and U1799 (N_1799,N_751,N_1108);
nor U1800 (N_1800,N_1418,N_1785);
and U1801 (N_1801,N_1411,N_1400);
or U1802 (N_1802,N_1635,N_1748);
nor U1803 (N_1803,N_1603,N_1641);
and U1804 (N_1804,N_1611,N_1541);
nand U1805 (N_1805,N_1780,N_1728);
nor U1806 (N_1806,N_1204,N_1619);
nor U1807 (N_1807,N_1661,N_1290);
or U1808 (N_1808,N_1225,N_1300);
nor U1809 (N_1809,N_1386,N_1244);
nor U1810 (N_1810,N_1508,N_1348);
and U1811 (N_1811,N_1500,N_1586);
and U1812 (N_1812,N_1520,N_1387);
nor U1813 (N_1813,N_1401,N_1471);
nand U1814 (N_1814,N_1605,N_1773);
or U1815 (N_1815,N_1797,N_1629);
nor U1816 (N_1816,N_1336,N_1534);
nand U1817 (N_1817,N_1596,N_1454);
or U1818 (N_1818,N_1683,N_1590);
and U1819 (N_1819,N_1342,N_1364);
or U1820 (N_1820,N_1309,N_1388);
or U1821 (N_1821,N_1432,N_1578);
nand U1822 (N_1822,N_1742,N_1535);
and U1823 (N_1823,N_1567,N_1207);
nand U1824 (N_1824,N_1221,N_1550);
and U1825 (N_1825,N_1260,N_1781);
nor U1826 (N_1826,N_1558,N_1798);
nand U1827 (N_1827,N_1750,N_1408);
or U1828 (N_1828,N_1227,N_1493);
and U1829 (N_1829,N_1465,N_1673);
and U1830 (N_1830,N_1371,N_1580);
nor U1831 (N_1831,N_1701,N_1599);
nor U1832 (N_1832,N_1627,N_1369);
nor U1833 (N_1833,N_1698,N_1726);
and U1834 (N_1834,N_1690,N_1390);
nor U1835 (N_1835,N_1623,N_1437);
nand U1836 (N_1836,N_1756,N_1582);
and U1837 (N_1837,N_1251,N_1425);
nor U1838 (N_1838,N_1604,N_1243);
or U1839 (N_1839,N_1575,N_1306);
and U1840 (N_1840,N_1659,N_1211);
or U1841 (N_1841,N_1694,N_1380);
nor U1842 (N_1842,N_1600,N_1555);
or U1843 (N_1843,N_1431,N_1275);
nor U1844 (N_1844,N_1654,N_1291);
and U1845 (N_1845,N_1542,N_1759);
or U1846 (N_1846,N_1624,N_1526);
nor U1847 (N_1847,N_1305,N_1710);
nand U1848 (N_1848,N_1258,N_1311);
nand U1849 (N_1849,N_1469,N_1206);
or U1850 (N_1850,N_1328,N_1723);
or U1851 (N_1851,N_1315,N_1532);
and U1852 (N_1852,N_1621,N_1419);
and U1853 (N_1853,N_1547,N_1761);
or U1854 (N_1854,N_1446,N_1436);
nor U1855 (N_1855,N_1791,N_1491);
or U1856 (N_1856,N_1396,N_1378);
nand U1857 (N_1857,N_1598,N_1265);
or U1858 (N_1858,N_1571,N_1499);
or U1859 (N_1859,N_1770,N_1540);
nand U1860 (N_1860,N_1398,N_1583);
nor U1861 (N_1861,N_1686,N_1415);
nand U1862 (N_1862,N_1638,N_1358);
nand U1863 (N_1863,N_1664,N_1402);
and U1864 (N_1864,N_1769,N_1682);
or U1865 (N_1865,N_1608,N_1472);
and U1866 (N_1866,N_1261,N_1650);
and U1867 (N_1867,N_1434,N_1671);
nor U1868 (N_1868,N_1556,N_1457);
or U1869 (N_1869,N_1395,N_1721);
nand U1870 (N_1870,N_1767,N_1361);
nand U1871 (N_1871,N_1569,N_1745);
nor U1872 (N_1872,N_1539,N_1775);
and U1873 (N_1873,N_1612,N_1692);
nand U1874 (N_1874,N_1743,N_1372);
or U1875 (N_1875,N_1444,N_1697);
and U1876 (N_1876,N_1696,N_1771);
nor U1877 (N_1877,N_1518,N_1318);
and U1878 (N_1878,N_1549,N_1533);
or U1879 (N_1879,N_1463,N_1787);
or U1880 (N_1880,N_1732,N_1570);
and U1881 (N_1881,N_1676,N_1393);
nand U1882 (N_1882,N_1262,N_1294);
or U1883 (N_1883,N_1588,N_1512);
and U1884 (N_1884,N_1259,N_1482);
or U1885 (N_1885,N_1385,N_1660);
and U1886 (N_1886,N_1579,N_1622);
or U1887 (N_1887,N_1651,N_1210);
and U1888 (N_1888,N_1462,N_1288);
nand U1889 (N_1889,N_1617,N_1447);
and U1890 (N_1890,N_1779,N_1216);
or U1891 (N_1891,N_1452,N_1413);
and U1892 (N_1892,N_1642,N_1296);
or U1893 (N_1893,N_1354,N_1248);
and U1894 (N_1894,N_1223,N_1610);
or U1895 (N_1895,N_1403,N_1502);
nand U1896 (N_1896,N_1422,N_1272);
and U1897 (N_1897,N_1584,N_1559);
and U1898 (N_1898,N_1631,N_1341);
and U1899 (N_1899,N_1509,N_1215);
or U1900 (N_1900,N_1752,N_1504);
nand U1901 (N_1901,N_1793,N_1203);
or U1902 (N_1902,N_1766,N_1657);
or U1903 (N_1903,N_1407,N_1636);
or U1904 (N_1904,N_1691,N_1298);
nand U1905 (N_1905,N_1427,N_1323);
and U1906 (N_1906,N_1331,N_1332);
and U1907 (N_1907,N_1230,N_1524);
nor U1908 (N_1908,N_1634,N_1320);
nor U1909 (N_1909,N_1490,N_1201);
nand U1910 (N_1910,N_1317,N_1740);
and U1911 (N_1911,N_1428,N_1576);
nor U1912 (N_1912,N_1370,N_1647);
or U1913 (N_1913,N_1754,N_1438);
and U1914 (N_1914,N_1392,N_1784);
nand U1915 (N_1915,N_1652,N_1351);
and U1916 (N_1916,N_1238,N_1565);
or U1917 (N_1917,N_1523,N_1783);
nor U1918 (N_1918,N_1794,N_1764);
nor U1919 (N_1919,N_1553,N_1321);
nand U1920 (N_1920,N_1356,N_1618);
nand U1921 (N_1921,N_1768,N_1441);
or U1922 (N_1922,N_1365,N_1552);
nor U1923 (N_1923,N_1782,N_1377);
nor U1924 (N_1924,N_1443,N_1246);
and U1925 (N_1925,N_1391,N_1359);
or U1926 (N_1926,N_1355,N_1234);
nor U1927 (N_1927,N_1276,N_1573);
or U1928 (N_1928,N_1645,N_1360);
and U1929 (N_1929,N_1405,N_1267);
nand U1930 (N_1930,N_1412,N_1464);
nand U1931 (N_1931,N_1712,N_1724);
or U1932 (N_1932,N_1346,N_1551);
or U1933 (N_1933,N_1734,N_1302);
nor U1934 (N_1934,N_1406,N_1247);
nand U1935 (N_1935,N_1731,N_1497);
nor U1936 (N_1936,N_1480,N_1477);
or U1937 (N_1937,N_1777,N_1527);
nor U1938 (N_1938,N_1439,N_1442);
and U1939 (N_1939,N_1677,N_1574);
and U1940 (N_1940,N_1733,N_1467);
or U1941 (N_1941,N_1585,N_1543);
nor U1942 (N_1942,N_1609,N_1488);
or U1943 (N_1943,N_1648,N_1330);
nor U1944 (N_1944,N_1269,N_1685);
nor U1945 (N_1945,N_1277,N_1455);
and U1946 (N_1946,N_1693,N_1268);
nor U1947 (N_1947,N_1202,N_1772);
nor U1948 (N_1948,N_1792,N_1343);
or U1949 (N_1949,N_1283,N_1708);
and U1950 (N_1950,N_1278,N_1233);
or U1951 (N_1951,N_1451,N_1626);
or U1952 (N_1952,N_1738,N_1562);
nand U1953 (N_1953,N_1284,N_1394);
nand U1954 (N_1954,N_1257,N_1758);
and U1955 (N_1955,N_1461,N_1709);
and U1956 (N_1956,N_1459,N_1719);
and U1957 (N_1957,N_1445,N_1466);
or U1958 (N_1958,N_1531,N_1630);
nor U1959 (N_1959,N_1414,N_1749);
nand U1960 (N_1960,N_1592,N_1568);
nor U1961 (N_1961,N_1319,N_1666);
nor U1962 (N_1962,N_1560,N_1478);
nor U1963 (N_1963,N_1591,N_1699);
and U1964 (N_1964,N_1790,N_1270);
or U1965 (N_1965,N_1663,N_1473);
and U1966 (N_1966,N_1633,N_1389);
or U1967 (N_1967,N_1453,N_1614);
nand U1968 (N_1968,N_1561,N_1684);
or U1969 (N_1969,N_1236,N_1668);
or U1970 (N_1970,N_1587,N_1498);
nor U1971 (N_1971,N_1707,N_1301);
nand U1972 (N_1972,N_1308,N_1566);
or U1973 (N_1973,N_1513,N_1607);
nand U1974 (N_1974,N_1212,N_1514);
and U1975 (N_1975,N_1433,N_1313);
nor U1976 (N_1976,N_1546,N_1384);
or U1977 (N_1977,N_1687,N_1220);
or U1978 (N_1978,N_1640,N_1487);
or U1979 (N_1979,N_1322,N_1544);
nand U1980 (N_1980,N_1572,N_1620);
or U1981 (N_1981,N_1339,N_1688);
and U1982 (N_1982,N_1352,N_1510);
or U1983 (N_1983,N_1327,N_1448);
nor U1984 (N_1984,N_1727,N_1675);
nand U1985 (N_1985,N_1333,N_1702);
nand U1986 (N_1986,N_1737,N_1324);
nor U1987 (N_1987,N_1705,N_1674);
nand U1988 (N_1988,N_1450,N_1314);
xnor U1989 (N_1989,N_1435,N_1746);
nand U1990 (N_1990,N_1337,N_1706);
and U1991 (N_1991,N_1209,N_1410);
or U1992 (N_1992,N_1736,N_1237);
and U1993 (N_1993,N_1286,N_1280);
or U1994 (N_1994,N_1762,N_1700);
or U1995 (N_1995,N_1293,N_1672);
or U1996 (N_1996,N_1242,N_1379);
or U1997 (N_1997,N_1338,N_1226);
xor U1998 (N_1998,N_1200,N_1397);
nor U1999 (N_1999,N_1557,N_1577);
or U2000 (N_2000,N_1789,N_1429);
or U2001 (N_2001,N_1501,N_1335);
nor U2002 (N_2002,N_1765,N_1751);
nor U2003 (N_2003,N_1409,N_1417);
nand U2004 (N_2004,N_1213,N_1366);
and U2005 (N_2005,N_1628,N_1208);
and U2006 (N_2006,N_1639,N_1615);
nand U2007 (N_2007,N_1521,N_1279);
or U2008 (N_2008,N_1720,N_1519);
nand U2009 (N_2009,N_1704,N_1597);
or U2010 (N_2010,N_1649,N_1753);
and U2011 (N_2011,N_1416,N_1744);
nor U2012 (N_2012,N_1662,N_1474);
nor U2013 (N_2013,N_1430,N_1292);
and U2014 (N_2014,N_1739,N_1374);
or U2015 (N_2015,N_1424,N_1481);
nand U2016 (N_2016,N_1722,N_1678);
or U2017 (N_2017,N_1287,N_1515);
nand U2018 (N_2018,N_1581,N_1589);
nand U2019 (N_2019,N_1646,N_1282);
and U2020 (N_2020,N_1755,N_1741);
and U2021 (N_2021,N_1266,N_1363);
nor U2022 (N_2022,N_1484,N_1730);
or U2023 (N_2023,N_1367,N_1228);
and U2024 (N_2024,N_1456,N_1274);
nand U2025 (N_2025,N_1214,N_1725);
nor U2026 (N_2026,N_1253,N_1256);
and U2027 (N_2027,N_1511,N_1423);
or U2028 (N_2028,N_1667,N_1517);
or U2029 (N_2029,N_1538,N_1217);
nor U2030 (N_2030,N_1316,N_1613);
nor U2031 (N_2031,N_1285,N_1537);
nor U2032 (N_2032,N_1658,N_1289);
or U2033 (N_2033,N_1264,N_1495);
nor U2034 (N_2034,N_1205,N_1329);
nand U2035 (N_2035,N_1345,N_1757);
or U2036 (N_2036,N_1679,N_1334);
and U2037 (N_2037,N_1326,N_1426);
nand U2038 (N_2038,N_1670,N_1601);
or U2039 (N_2039,N_1476,N_1563);
nand U2040 (N_2040,N_1494,N_1479);
nand U2041 (N_2041,N_1249,N_1516);
or U2042 (N_2042,N_1254,N_1713);
or U2043 (N_2043,N_1564,N_1353);
and U2044 (N_2044,N_1774,N_1350);
nand U2045 (N_2045,N_1763,N_1503);
and U2046 (N_2046,N_1470,N_1241);
or U2047 (N_2047,N_1376,N_1554);
or U2048 (N_2048,N_1536,N_1747);
nand U2049 (N_2049,N_1304,N_1310);
nor U2050 (N_2050,N_1729,N_1606);
nand U2051 (N_2051,N_1344,N_1485);
and U2052 (N_2052,N_1695,N_1460);
and U2053 (N_2053,N_1522,N_1506);
and U2054 (N_2054,N_1224,N_1656);
or U2055 (N_2055,N_1449,N_1643);
nand U2056 (N_2056,N_1593,N_1669);
nand U2057 (N_2057,N_1382,N_1625);
nand U2058 (N_2058,N_1475,N_1735);
nand U2059 (N_2059,N_1637,N_1680);
or U2060 (N_2060,N_1786,N_1528);
or U2061 (N_2061,N_1548,N_1689);
or U2062 (N_2062,N_1507,N_1489);
nor U2063 (N_2063,N_1245,N_1232);
nand U2064 (N_2064,N_1594,N_1229);
nor U2065 (N_2065,N_1525,N_1250);
nor U2066 (N_2066,N_1715,N_1357);
nor U2067 (N_2067,N_1255,N_1231);
and U2068 (N_2068,N_1760,N_1349);
nand U2069 (N_2069,N_1340,N_1716);
or U2070 (N_2070,N_1440,N_1530);
nand U2071 (N_2071,N_1799,N_1235);
nor U2072 (N_2072,N_1653,N_1239);
or U2073 (N_2073,N_1263,N_1222);
nor U2074 (N_2074,N_1703,N_1795);
nand U2075 (N_2075,N_1655,N_1404);
nand U2076 (N_2076,N_1545,N_1219);
nand U2077 (N_2077,N_1468,N_1496);
and U2078 (N_2078,N_1632,N_1796);
nand U2079 (N_2079,N_1297,N_1644);
or U2080 (N_2080,N_1325,N_1616);
or U2081 (N_2081,N_1240,N_1373);
or U2082 (N_2082,N_1665,N_1375);
and U2083 (N_2083,N_1362,N_1486);
and U2084 (N_2084,N_1273,N_1505);
or U2085 (N_2085,N_1312,N_1303);
nand U2086 (N_2086,N_1788,N_1714);
and U2087 (N_2087,N_1271,N_1383);
nand U2088 (N_2088,N_1252,N_1421);
and U2089 (N_2089,N_1778,N_1681);
nand U2090 (N_2090,N_1483,N_1381);
and U2091 (N_2091,N_1218,N_1602);
and U2092 (N_2092,N_1458,N_1492);
nor U2093 (N_2093,N_1307,N_1776);
and U2094 (N_2094,N_1718,N_1368);
nor U2095 (N_2095,N_1420,N_1717);
or U2096 (N_2096,N_1295,N_1595);
and U2097 (N_2097,N_1529,N_1711);
nor U2098 (N_2098,N_1299,N_1347);
and U2099 (N_2099,N_1399,N_1281);
and U2100 (N_2100,N_1238,N_1604);
nand U2101 (N_2101,N_1702,N_1701);
or U2102 (N_2102,N_1434,N_1428);
or U2103 (N_2103,N_1377,N_1314);
nand U2104 (N_2104,N_1719,N_1501);
nor U2105 (N_2105,N_1714,N_1772);
nor U2106 (N_2106,N_1728,N_1267);
or U2107 (N_2107,N_1484,N_1388);
nand U2108 (N_2108,N_1574,N_1245);
nand U2109 (N_2109,N_1448,N_1481);
nor U2110 (N_2110,N_1733,N_1221);
nor U2111 (N_2111,N_1345,N_1315);
nand U2112 (N_2112,N_1471,N_1513);
and U2113 (N_2113,N_1744,N_1684);
nand U2114 (N_2114,N_1709,N_1652);
nand U2115 (N_2115,N_1557,N_1716);
and U2116 (N_2116,N_1374,N_1799);
or U2117 (N_2117,N_1349,N_1748);
nor U2118 (N_2118,N_1553,N_1347);
nand U2119 (N_2119,N_1556,N_1745);
nor U2120 (N_2120,N_1332,N_1658);
nand U2121 (N_2121,N_1475,N_1215);
nand U2122 (N_2122,N_1727,N_1738);
or U2123 (N_2123,N_1480,N_1343);
nand U2124 (N_2124,N_1761,N_1731);
nand U2125 (N_2125,N_1226,N_1735);
and U2126 (N_2126,N_1214,N_1349);
nor U2127 (N_2127,N_1410,N_1227);
nand U2128 (N_2128,N_1569,N_1403);
and U2129 (N_2129,N_1511,N_1572);
nor U2130 (N_2130,N_1779,N_1268);
xnor U2131 (N_2131,N_1347,N_1615);
and U2132 (N_2132,N_1364,N_1224);
nand U2133 (N_2133,N_1677,N_1329);
nand U2134 (N_2134,N_1383,N_1671);
nor U2135 (N_2135,N_1463,N_1404);
nand U2136 (N_2136,N_1400,N_1377);
nor U2137 (N_2137,N_1755,N_1442);
or U2138 (N_2138,N_1590,N_1212);
nor U2139 (N_2139,N_1263,N_1743);
or U2140 (N_2140,N_1239,N_1435);
nor U2141 (N_2141,N_1776,N_1409);
nor U2142 (N_2142,N_1343,N_1766);
nand U2143 (N_2143,N_1486,N_1494);
nand U2144 (N_2144,N_1220,N_1554);
nand U2145 (N_2145,N_1487,N_1455);
or U2146 (N_2146,N_1598,N_1309);
nand U2147 (N_2147,N_1673,N_1597);
and U2148 (N_2148,N_1785,N_1348);
nor U2149 (N_2149,N_1392,N_1211);
nand U2150 (N_2150,N_1300,N_1555);
nor U2151 (N_2151,N_1797,N_1311);
and U2152 (N_2152,N_1776,N_1752);
nand U2153 (N_2153,N_1283,N_1200);
nand U2154 (N_2154,N_1527,N_1794);
or U2155 (N_2155,N_1265,N_1576);
nor U2156 (N_2156,N_1608,N_1659);
or U2157 (N_2157,N_1683,N_1514);
nand U2158 (N_2158,N_1422,N_1493);
nand U2159 (N_2159,N_1768,N_1259);
and U2160 (N_2160,N_1272,N_1796);
and U2161 (N_2161,N_1345,N_1634);
nand U2162 (N_2162,N_1753,N_1378);
nand U2163 (N_2163,N_1569,N_1454);
or U2164 (N_2164,N_1431,N_1704);
and U2165 (N_2165,N_1376,N_1301);
nand U2166 (N_2166,N_1483,N_1541);
nand U2167 (N_2167,N_1353,N_1510);
nor U2168 (N_2168,N_1509,N_1514);
nand U2169 (N_2169,N_1780,N_1785);
nand U2170 (N_2170,N_1304,N_1706);
or U2171 (N_2171,N_1695,N_1766);
and U2172 (N_2172,N_1463,N_1319);
and U2173 (N_2173,N_1596,N_1681);
nor U2174 (N_2174,N_1377,N_1348);
and U2175 (N_2175,N_1309,N_1627);
or U2176 (N_2176,N_1312,N_1423);
or U2177 (N_2177,N_1622,N_1485);
or U2178 (N_2178,N_1403,N_1621);
nand U2179 (N_2179,N_1777,N_1618);
and U2180 (N_2180,N_1771,N_1758);
and U2181 (N_2181,N_1511,N_1670);
and U2182 (N_2182,N_1497,N_1676);
nand U2183 (N_2183,N_1579,N_1605);
nand U2184 (N_2184,N_1767,N_1267);
nand U2185 (N_2185,N_1618,N_1720);
nor U2186 (N_2186,N_1208,N_1653);
nand U2187 (N_2187,N_1493,N_1356);
and U2188 (N_2188,N_1397,N_1376);
or U2189 (N_2189,N_1628,N_1430);
nor U2190 (N_2190,N_1382,N_1303);
nand U2191 (N_2191,N_1379,N_1677);
or U2192 (N_2192,N_1606,N_1550);
and U2193 (N_2193,N_1205,N_1282);
nand U2194 (N_2194,N_1534,N_1586);
nor U2195 (N_2195,N_1391,N_1541);
and U2196 (N_2196,N_1604,N_1690);
nor U2197 (N_2197,N_1770,N_1720);
or U2198 (N_2198,N_1697,N_1474);
or U2199 (N_2199,N_1237,N_1436);
and U2200 (N_2200,N_1305,N_1452);
nor U2201 (N_2201,N_1579,N_1469);
and U2202 (N_2202,N_1494,N_1606);
or U2203 (N_2203,N_1579,N_1684);
xnor U2204 (N_2204,N_1642,N_1611);
and U2205 (N_2205,N_1791,N_1621);
nand U2206 (N_2206,N_1670,N_1735);
nor U2207 (N_2207,N_1639,N_1701);
or U2208 (N_2208,N_1785,N_1796);
or U2209 (N_2209,N_1659,N_1751);
and U2210 (N_2210,N_1489,N_1647);
nor U2211 (N_2211,N_1664,N_1617);
or U2212 (N_2212,N_1790,N_1597);
and U2213 (N_2213,N_1326,N_1667);
nor U2214 (N_2214,N_1539,N_1723);
nor U2215 (N_2215,N_1455,N_1630);
or U2216 (N_2216,N_1452,N_1595);
nor U2217 (N_2217,N_1274,N_1399);
nand U2218 (N_2218,N_1553,N_1307);
or U2219 (N_2219,N_1435,N_1389);
and U2220 (N_2220,N_1563,N_1266);
or U2221 (N_2221,N_1344,N_1527);
nor U2222 (N_2222,N_1404,N_1764);
nand U2223 (N_2223,N_1599,N_1579);
and U2224 (N_2224,N_1771,N_1205);
or U2225 (N_2225,N_1270,N_1351);
or U2226 (N_2226,N_1351,N_1280);
and U2227 (N_2227,N_1388,N_1757);
and U2228 (N_2228,N_1408,N_1326);
or U2229 (N_2229,N_1685,N_1347);
nor U2230 (N_2230,N_1586,N_1299);
nand U2231 (N_2231,N_1435,N_1636);
and U2232 (N_2232,N_1494,N_1322);
nor U2233 (N_2233,N_1567,N_1431);
or U2234 (N_2234,N_1782,N_1205);
nand U2235 (N_2235,N_1334,N_1794);
nand U2236 (N_2236,N_1429,N_1339);
or U2237 (N_2237,N_1693,N_1370);
nor U2238 (N_2238,N_1421,N_1316);
or U2239 (N_2239,N_1406,N_1525);
nor U2240 (N_2240,N_1397,N_1485);
nor U2241 (N_2241,N_1279,N_1423);
and U2242 (N_2242,N_1790,N_1771);
nand U2243 (N_2243,N_1706,N_1682);
nand U2244 (N_2244,N_1353,N_1606);
nor U2245 (N_2245,N_1686,N_1460);
nand U2246 (N_2246,N_1761,N_1680);
xor U2247 (N_2247,N_1529,N_1475);
and U2248 (N_2248,N_1501,N_1517);
nand U2249 (N_2249,N_1276,N_1483);
nor U2250 (N_2250,N_1562,N_1284);
nor U2251 (N_2251,N_1451,N_1220);
and U2252 (N_2252,N_1738,N_1435);
nor U2253 (N_2253,N_1294,N_1793);
or U2254 (N_2254,N_1313,N_1407);
nand U2255 (N_2255,N_1777,N_1454);
nor U2256 (N_2256,N_1696,N_1552);
nand U2257 (N_2257,N_1585,N_1400);
nor U2258 (N_2258,N_1600,N_1205);
nor U2259 (N_2259,N_1394,N_1685);
nor U2260 (N_2260,N_1559,N_1547);
nor U2261 (N_2261,N_1281,N_1359);
nand U2262 (N_2262,N_1618,N_1667);
nor U2263 (N_2263,N_1482,N_1556);
nor U2264 (N_2264,N_1415,N_1202);
nand U2265 (N_2265,N_1249,N_1709);
or U2266 (N_2266,N_1476,N_1582);
nand U2267 (N_2267,N_1688,N_1704);
nor U2268 (N_2268,N_1202,N_1740);
nor U2269 (N_2269,N_1557,N_1614);
and U2270 (N_2270,N_1497,N_1331);
nor U2271 (N_2271,N_1642,N_1567);
nor U2272 (N_2272,N_1420,N_1310);
or U2273 (N_2273,N_1308,N_1794);
nor U2274 (N_2274,N_1694,N_1652);
nor U2275 (N_2275,N_1438,N_1394);
nand U2276 (N_2276,N_1797,N_1765);
and U2277 (N_2277,N_1787,N_1720);
or U2278 (N_2278,N_1568,N_1248);
or U2279 (N_2279,N_1740,N_1264);
nand U2280 (N_2280,N_1300,N_1653);
and U2281 (N_2281,N_1609,N_1627);
nor U2282 (N_2282,N_1731,N_1496);
xnor U2283 (N_2283,N_1663,N_1304);
nor U2284 (N_2284,N_1308,N_1483);
or U2285 (N_2285,N_1247,N_1671);
and U2286 (N_2286,N_1311,N_1649);
and U2287 (N_2287,N_1462,N_1660);
nand U2288 (N_2288,N_1315,N_1464);
or U2289 (N_2289,N_1765,N_1246);
nor U2290 (N_2290,N_1769,N_1587);
nand U2291 (N_2291,N_1584,N_1556);
nor U2292 (N_2292,N_1767,N_1339);
and U2293 (N_2293,N_1632,N_1533);
nand U2294 (N_2294,N_1560,N_1269);
and U2295 (N_2295,N_1426,N_1670);
or U2296 (N_2296,N_1567,N_1797);
and U2297 (N_2297,N_1216,N_1435);
and U2298 (N_2298,N_1477,N_1326);
and U2299 (N_2299,N_1415,N_1782);
and U2300 (N_2300,N_1614,N_1420);
or U2301 (N_2301,N_1532,N_1784);
and U2302 (N_2302,N_1620,N_1540);
nor U2303 (N_2303,N_1446,N_1693);
or U2304 (N_2304,N_1734,N_1500);
and U2305 (N_2305,N_1331,N_1287);
and U2306 (N_2306,N_1473,N_1612);
or U2307 (N_2307,N_1565,N_1275);
nand U2308 (N_2308,N_1679,N_1543);
nand U2309 (N_2309,N_1428,N_1325);
and U2310 (N_2310,N_1439,N_1543);
and U2311 (N_2311,N_1284,N_1710);
xnor U2312 (N_2312,N_1437,N_1442);
or U2313 (N_2313,N_1305,N_1499);
and U2314 (N_2314,N_1700,N_1769);
xor U2315 (N_2315,N_1723,N_1612);
nor U2316 (N_2316,N_1785,N_1545);
nor U2317 (N_2317,N_1562,N_1221);
or U2318 (N_2318,N_1247,N_1473);
nand U2319 (N_2319,N_1797,N_1747);
nand U2320 (N_2320,N_1782,N_1423);
and U2321 (N_2321,N_1730,N_1770);
nor U2322 (N_2322,N_1617,N_1713);
and U2323 (N_2323,N_1531,N_1236);
nand U2324 (N_2324,N_1725,N_1215);
nand U2325 (N_2325,N_1566,N_1372);
nor U2326 (N_2326,N_1687,N_1733);
nor U2327 (N_2327,N_1409,N_1783);
nor U2328 (N_2328,N_1383,N_1425);
or U2329 (N_2329,N_1479,N_1618);
or U2330 (N_2330,N_1740,N_1339);
and U2331 (N_2331,N_1388,N_1356);
xnor U2332 (N_2332,N_1318,N_1411);
nor U2333 (N_2333,N_1219,N_1561);
or U2334 (N_2334,N_1251,N_1755);
and U2335 (N_2335,N_1655,N_1284);
nand U2336 (N_2336,N_1659,N_1525);
nand U2337 (N_2337,N_1321,N_1613);
or U2338 (N_2338,N_1755,N_1353);
nand U2339 (N_2339,N_1771,N_1665);
nand U2340 (N_2340,N_1477,N_1332);
or U2341 (N_2341,N_1477,N_1722);
and U2342 (N_2342,N_1771,N_1217);
nand U2343 (N_2343,N_1281,N_1696);
nor U2344 (N_2344,N_1688,N_1221);
or U2345 (N_2345,N_1649,N_1354);
nor U2346 (N_2346,N_1394,N_1471);
nor U2347 (N_2347,N_1715,N_1415);
and U2348 (N_2348,N_1296,N_1401);
nand U2349 (N_2349,N_1697,N_1341);
or U2350 (N_2350,N_1736,N_1548);
or U2351 (N_2351,N_1646,N_1523);
nor U2352 (N_2352,N_1699,N_1624);
nand U2353 (N_2353,N_1288,N_1724);
nor U2354 (N_2354,N_1665,N_1590);
or U2355 (N_2355,N_1397,N_1550);
nand U2356 (N_2356,N_1258,N_1267);
and U2357 (N_2357,N_1588,N_1749);
nor U2358 (N_2358,N_1466,N_1685);
nand U2359 (N_2359,N_1247,N_1391);
nand U2360 (N_2360,N_1622,N_1627);
and U2361 (N_2361,N_1481,N_1345);
or U2362 (N_2362,N_1250,N_1385);
nand U2363 (N_2363,N_1519,N_1516);
nand U2364 (N_2364,N_1219,N_1711);
or U2365 (N_2365,N_1713,N_1755);
or U2366 (N_2366,N_1548,N_1200);
or U2367 (N_2367,N_1537,N_1403);
and U2368 (N_2368,N_1286,N_1520);
nor U2369 (N_2369,N_1364,N_1331);
and U2370 (N_2370,N_1472,N_1597);
nand U2371 (N_2371,N_1467,N_1712);
nor U2372 (N_2372,N_1404,N_1367);
or U2373 (N_2373,N_1258,N_1388);
and U2374 (N_2374,N_1578,N_1698);
nand U2375 (N_2375,N_1241,N_1503);
and U2376 (N_2376,N_1379,N_1237);
and U2377 (N_2377,N_1331,N_1469);
nor U2378 (N_2378,N_1282,N_1609);
or U2379 (N_2379,N_1586,N_1552);
nor U2380 (N_2380,N_1348,N_1418);
and U2381 (N_2381,N_1427,N_1514);
nand U2382 (N_2382,N_1649,N_1719);
nor U2383 (N_2383,N_1221,N_1464);
or U2384 (N_2384,N_1222,N_1614);
and U2385 (N_2385,N_1415,N_1410);
or U2386 (N_2386,N_1342,N_1295);
nand U2387 (N_2387,N_1304,N_1495);
nor U2388 (N_2388,N_1672,N_1565);
and U2389 (N_2389,N_1208,N_1523);
xnor U2390 (N_2390,N_1449,N_1431);
or U2391 (N_2391,N_1477,N_1604);
xor U2392 (N_2392,N_1602,N_1727);
and U2393 (N_2393,N_1327,N_1759);
or U2394 (N_2394,N_1542,N_1620);
and U2395 (N_2395,N_1203,N_1303);
nand U2396 (N_2396,N_1750,N_1603);
and U2397 (N_2397,N_1361,N_1639);
and U2398 (N_2398,N_1430,N_1319);
nor U2399 (N_2399,N_1640,N_1336);
and U2400 (N_2400,N_2071,N_1914);
nor U2401 (N_2401,N_2101,N_2173);
nor U2402 (N_2402,N_2135,N_2192);
nor U2403 (N_2403,N_1846,N_1887);
and U2404 (N_2404,N_1835,N_2337);
nor U2405 (N_2405,N_2289,N_2222);
nand U2406 (N_2406,N_2338,N_2002);
nor U2407 (N_2407,N_2371,N_2282);
and U2408 (N_2408,N_1948,N_1903);
or U2409 (N_2409,N_2179,N_2311);
nor U2410 (N_2410,N_1837,N_2017);
nand U2411 (N_2411,N_1998,N_1985);
and U2412 (N_2412,N_2156,N_2115);
nand U2413 (N_2413,N_1889,N_2004);
or U2414 (N_2414,N_2062,N_2044);
and U2415 (N_2415,N_1978,N_2176);
or U2416 (N_2416,N_2155,N_2328);
nand U2417 (N_2417,N_2309,N_2237);
or U2418 (N_2418,N_2157,N_2164);
or U2419 (N_2419,N_2194,N_2057);
nor U2420 (N_2420,N_1994,N_2011);
and U2421 (N_2421,N_2379,N_2297);
nor U2422 (N_2422,N_1969,N_2375);
or U2423 (N_2423,N_2386,N_2060);
or U2424 (N_2424,N_1920,N_2049);
nor U2425 (N_2425,N_1809,N_1943);
nand U2426 (N_2426,N_2113,N_2267);
and U2427 (N_2427,N_2263,N_2242);
nor U2428 (N_2428,N_2254,N_2315);
nor U2429 (N_2429,N_2239,N_2108);
or U2430 (N_2430,N_2147,N_2170);
or U2431 (N_2431,N_2109,N_2260);
and U2432 (N_2432,N_1944,N_2078);
nand U2433 (N_2433,N_1840,N_2354);
and U2434 (N_2434,N_2075,N_2358);
nand U2435 (N_2435,N_2080,N_2180);
or U2436 (N_2436,N_2066,N_1947);
and U2437 (N_2437,N_2266,N_1866);
or U2438 (N_2438,N_2177,N_2185);
and U2439 (N_2439,N_1960,N_2050);
and U2440 (N_2440,N_2208,N_2046);
or U2441 (N_2441,N_2035,N_1908);
nor U2442 (N_2442,N_1891,N_2143);
nor U2443 (N_2443,N_1935,N_2335);
and U2444 (N_2444,N_2212,N_2387);
nor U2445 (N_2445,N_2224,N_1800);
or U2446 (N_2446,N_1828,N_2161);
nand U2447 (N_2447,N_2376,N_1855);
nand U2448 (N_2448,N_2174,N_2305);
nor U2449 (N_2449,N_2366,N_2076);
and U2450 (N_2450,N_1818,N_1955);
nor U2451 (N_2451,N_1839,N_1951);
nand U2452 (N_2452,N_2111,N_1897);
and U2453 (N_2453,N_2356,N_2063);
and U2454 (N_2454,N_2023,N_1876);
nand U2455 (N_2455,N_1885,N_2107);
nor U2456 (N_2456,N_2265,N_1805);
or U2457 (N_2457,N_1848,N_2350);
and U2458 (N_2458,N_1850,N_2130);
nor U2459 (N_2459,N_2284,N_1962);
nand U2460 (N_2460,N_1958,N_2392);
and U2461 (N_2461,N_1932,N_1827);
nand U2462 (N_2462,N_1918,N_1817);
and U2463 (N_2463,N_2093,N_1814);
nor U2464 (N_2464,N_1857,N_2318);
nand U2465 (N_2465,N_1851,N_2285);
and U2466 (N_2466,N_1934,N_2127);
and U2467 (N_2467,N_1841,N_2132);
and U2468 (N_2468,N_2280,N_2074);
nand U2469 (N_2469,N_2020,N_1931);
and U2470 (N_2470,N_2040,N_1939);
or U2471 (N_2471,N_2148,N_2008);
or U2472 (N_2472,N_2259,N_1825);
nor U2473 (N_2473,N_1813,N_2162);
nand U2474 (N_2474,N_2165,N_1988);
and U2475 (N_2475,N_1956,N_1957);
and U2476 (N_2476,N_1886,N_2277);
nand U2477 (N_2477,N_1912,N_2047);
nand U2478 (N_2478,N_1976,N_2056);
and U2479 (N_2479,N_1815,N_2045);
or U2480 (N_2480,N_2152,N_2058);
nand U2481 (N_2481,N_2088,N_1870);
or U2482 (N_2482,N_2031,N_2333);
or U2483 (N_2483,N_2121,N_2264);
nand U2484 (N_2484,N_2306,N_2225);
nor U2485 (N_2485,N_2012,N_1804);
or U2486 (N_2486,N_2229,N_2244);
or U2487 (N_2487,N_2330,N_2106);
or U2488 (N_2488,N_2013,N_2251);
or U2489 (N_2489,N_2268,N_2191);
nor U2490 (N_2490,N_1895,N_2167);
and U2491 (N_2491,N_1854,N_1911);
and U2492 (N_2492,N_2153,N_2054);
nor U2493 (N_2493,N_2223,N_2238);
nor U2494 (N_2494,N_2043,N_1875);
nand U2495 (N_2495,N_2279,N_2367);
nor U2496 (N_2496,N_2114,N_2384);
nand U2497 (N_2497,N_2334,N_2016);
nand U2498 (N_2498,N_1829,N_2015);
or U2499 (N_2499,N_2287,N_1880);
nor U2500 (N_2500,N_1992,N_2083);
or U2501 (N_2501,N_1922,N_2186);
and U2502 (N_2502,N_2304,N_2316);
or U2503 (N_2503,N_2131,N_2068);
nor U2504 (N_2504,N_1884,N_2144);
nor U2505 (N_2505,N_2141,N_1989);
nor U2506 (N_2506,N_2018,N_1819);
and U2507 (N_2507,N_2373,N_2134);
or U2508 (N_2508,N_2308,N_2369);
or U2509 (N_2509,N_2301,N_1861);
nand U2510 (N_2510,N_2230,N_2150);
and U2511 (N_2511,N_2325,N_1975);
or U2512 (N_2512,N_2110,N_1982);
nand U2513 (N_2513,N_2365,N_2032);
and U2514 (N_2514,N_2278,N_2341);
nor U2515 (N_2515,N_1890,N_1919);
nand U2516 (N_2516,N_2118,N_1831);
and U2517 (N_2517,N_2184,N_1898);
and U2518 (N_2518,N_2061,N_2104);
or U2519 (N_2519,N_1970,N_2357);
nor U2520 (N_2520,N_1842,N_2105);
nor U2521 (N_2521,N_2295,N_1987);
and U2522 (N_2522,N_2323,N_2202);
and U2523 (N_2523,N_1984,N_2321);
nor U2524 (N_2524,N_2226,N_2204);
or U2525 (N_2525,N_2030,N_1983);
or U2526 (N_2526,N_2236,N_2089);
or U2527 (N_2527,N_1968,N_1858);
nand U2528 (N_2528,N_2175,N_1961);
nand U2529 (N_2529,N_1972,N_2188);
nand U2530 (N_2530,N_1964,N_1959);
nor U2531 (N_2531,N_2073,N_2235);
nand U2532 (N_2532,N_2378,N_2055);
nand U2533 (N_2533,N_2160,N_2228);
and U2534 (N_2534,N_1971,N_2122);
or U2535 (N_2535,N_2079,N_2261);
nor U2536 (N_2536,N_2381,N_1833);
and U2537 (N_2537,N_2178,N_2036);
nand U2538 (N_2538,N_1926,N_1990);
and U2539 (N_2539,N_2291,N_2019);
nor U2540 (N_2540,N_1917,N_2048);
nand U2541 (N_2541,N_2293,N_2125);
xor U2542 (N_2542,N_2273,N_2317);
and U2543 (N_2543,N_2014,N_2352);
or U2544 (N_2544,N_2219,N_2041);
xnor U2545 (N_2545,N_1869,N_1907);
nor U2546 (N_2546,N_1965,N_1810);
and U2547 (N_2547,N_2339,N_2097);
and U2548 (N_2548,N_2025,N_2158);
nand U2549 (N_2549,N_1882,N_2037);
and U2550 (N_2550,N_2103,N_1945);
and U2551 (N_2551,N_2344,N_2374);
and U2552 (N_2552,N_1963,N_1999);
or U2553 (N_2553,N_2099,N_1834);
or U2554 (N_2554,N_2138,N_1967);
and U2555 (N_2555,N_1879,N_2190);
nor U2556 (N_2556,N_1946,N_1801);
or U2557 (N_2557,N_1995,N_2027);
nor U2558 (N_2558,N_2053,N_2253);
nand U2559 (N_2559,N_2052,N_2154);
or U2560 (N_2560,N_2021,N_2003);
nor U2561 (N_2561,N_2213,N_1977);
nor U2562 (N_2562,N_2022,N_1916);
nor U2563 (N_2563,N_2329,N_2388);
or U2564 (N_2564,N_2345,N_2391);
and U2565 (N_2565,N_2355,N_2248);
nor U2566 (N_2566,N_1865,N_2241);
nand U2567 (N_2567,N_2166,N_1868);
nand U2568 (N_2568,N_1832,N_2322);
or U2569 (N_2569,N_2262,N_2258);
nor U2570 (N_2570,N_2171,N_2303);
or U2571 (N_2571,N_1808,N_2302);
or U2572 (N_2572,N_2064,N_1823);
nand U2573 (N_2573,N_1996,N_1940);
and U2574 (N_2574,N_1864,N_1930);
nor U2575 (N_2575,N_1923,N_2240);
or U2576 (N_2576,N_2051,N_2163);
and U2577 (N_2577,N_1873,N_1860);
xor U2578 (N_2578,N_2327,N_1816);
or U2579 (N_2579,N_1847,N_1973);
and U2580 (N_2580,N_1921,N_2142);
nor U2581 (N_2581,N_2007,N_2187);
or U2582 (N_2582,N_2065,N_2368);
or U2583 (N_2583,N_2296,N_2136);
and U2584 (N_2584,N_1980,N_2256);
nor U2585 (N_2585,N_2126,N_2360);
and U2586 (N_2586,N_2059,N_1905);
nand U2587 (N_2587,N_2169,N_2397);
and U2588 (N_2588,N_2340,N_2332);
nand U2589 (N_2589,N_1812,N_2077);
nand U2590 (N_2590,N_1991,N_2086);
nand U2591 (N_2591,N_2133,N_2209);
and U2592 (N_2592,N_2197,N_1937);
or U2593 (N_2593,N_2276,N_1802);
and U2594 (N_2594,N_2070,N_2182);
nor U2595 (N_2595,N_2314,N_2000);
or U2596 (N_2596,N_2232,N_2390);
or U2597 (N_2597,N_2348,N_1900);
and U2598 (N_2598,N_2139,N_1953);
or U2599 (N_2599,N_1830,N_2140);
nand U2600 (N_2600,N_2290,N_1974);
and U2601 (N_2601,N_1899,N_1928);
nor U2602 (N_2602,N_1806,N_1979);
nand U2603 (N_2603,N_2200,N_2146);
nor U2604 (N_2604,N_1942,N_2310);
nand U2605 (N_2605,N_2382,N_2149);
nand U2606 (N_2606,N_1936,N_1993);
or U2607 (N_2607,N_2399,N_2269);
and U2608 (N_2608,N_1852,N_1986);
or U2609 (N_2609,N_2010,N_1938);
nand U2610 (N_2610,N_1896,N_2181);
nand U2611 (N_2611,N_1925,N_2094);
and U2612 (N_2612,N_2199,N_1913);
and U2613 (N_2613,N_2275,N_2361);
and U2614 (N_2614,N_1853,N_2005);
nand U2615 (N_2615,N_2359,N_1849);
or U2616 (N_2616,N_2283,N_2353);
or U2617 (N_2617,N_1803,N_2201);
nand U2618 (N_2618,N_2298,N_1892);
nor U2619 (N_2619,N_2081,N_2385);
nand U2620 (N_2620,N_1954,N_2028);
and U2621 (N_2621,N_2084,N_2039);
nor U2622 (N_2622,N_2172,N_2336);
nor U2623 (N_2623,N_2319,N_2343);
or U2624 (N_2624,N_1821,N_2255);
and U2625 (N_2625,N_2299,N_2286);
and U2626 (N_2626,N_2393,N_2196);
nor U2627 (N_2627,N_2072,N_2270);
and U2628 (N_2628,N_2009,N_2029);
and U2629 (N_2629,N_1893,N_2120);
or U2630 (N_2630,N_1867,N_2294);
or U2631 (N_2631,N_2362,N_2096);
nand U2632 (N_2632,N_2288,N_1872);
nor U2633 (N_2633,N_2117,N_2234);
nand U2634 (N_2634,N_2091,N_1874);
or U2635 (N_2635,N_2300,N_1878);
nand U2636 (N_2636,N_1881,N_2001);
or U2637 (N_2637,N_1904,N_2067);
nor U2638 (N_2638,N_1981,N_2324);
nor U2639 (N_2639,N_2349,N_2250);
and U2640 (N_2640,N_1838,N_2069);
and U2641 (N_2641,N_1966,N_1894);
or U2642 (N_2642,N_2312,N_1871);
nand U2643 (N_2643,N_2098,N_1924);
nand U2644 (N_2644,N_1856,N_2231);
and U2645 (N_2645,N_1811,N_2313);
or U2646 (N_2646,N_2217,N_1836);
nor U2647 (N_2647,N_1820,N_2189);
nand U2648 (N_2648,N_2128,N_2006);
and U2649 (N_2649,N_2129,N_1910);
nor U2650 (N_2650,N_2124,N_2233);
and U2651 (N_2651,N_2112,N_2207);
and U2652 (N_2652,N_2271,N_2252);
and U2653 (N_2653,N_1843,N_2151);
nor U2654 (N_2654,N_2218,N_2363);
nor U2655 (N_2655,N_2220,N_2307);
or U2656 (N_2656,N_2249,N_2100);
nand U2657 (N_2657,N_2168,N_1877);
or U2658 (N_2658,N_2380,N_2042);
nand U2659 (N_2659,N_1933,N_1906);
nand U2660 (N_2660,N_1863,N_2095);
nand U2661 (N_2661,N_2210,N_2342);
nor U2662 (N_2662,N_2159,N_2085);
and U2663 (N_2663,N_2274,N_1949);
nor U2664 (N_2664,N_2090,N_1950);
nor U2665 (N_2665,N_2257,N_2394);
or U2666 (N_2666,N_1822,N_2216);
nand U2667 (N_2667,N_1927,N_2351);
or U2668 (N_2668,N_2183,N_2038);
and U2669 (N_2669,N_2246,N_1888);
or U2670 (N_2670,N_1909,N_2119);
xor U2671 (N_2671,N_2383,N_2247);
nand U2672 (N_2672,N_1997,N_2205);
nand U2673 (N_2673,N_2292,N_2372);
nand U2674 (N_2674,N_1845,N_2377);
or U2675 (N_2675,N_1862,N_1941);
nand U2676 (N_2676,N_2145,N_2203);
or U2677 (N_2677,N_2193,N_1902);
and U2678 (N_2678,N_1807,N_2221);
nand U2679 (N_2679,N_2227,N_2326);
or U2680 (N_2680,N_2082,N_2395);
and U2681 (N_2681,N_2026,N_2137);
nand U2682 (N_2682,N_1826,N_2211);
nor U2683 (N_2683,N_1915,N_2389);
nor U2684 (N_2684,N_2102,N_2024);
nor U2685 (N_2685,N_1952,N_2215);
nand U2686 (N_2686,N_2272,N_2087);
nor U2687 (N_2687,N_2245,N_2034);
nor U2688 (N_2688,N_1883,N_2331);
nor U2689 (N_2689,N_2320,N_2198);
nand U2690 (N_2690,N_1929,N_2123);
and U2691 (N_2691,N_2195,N_2398);
or U2692 (N_2692,N_2092,N_2346);
and U2693 (N_2693,N_2033,N_2370);
and U2694 (N_2694,N_2396,N_2364);
or U2695 (N_2695,N_2281,N_2347);
and U2696 (N_2696,N_2243,N_1901);
nor U2697 (N_2697,N_1859,N_2206);
nand U2698 (N_2698,N_1844,N_2214);
and U2699 (N_2699,N_1824,N_2116);
nor U2700 (N_2700,N_2317,N_2198);
and U2701 (N_2701,N_2212,N_2382);
nand U2702 (N_2702,N_1808,N_1891);
and U2703 (N_2703,N_2364,N_1902);
nand U2704 (N_2704,N_2366,N_2242);
nand U2705 (N_2705,N_2036,N_2352);
and U2706 (N_2706,N_2370,N_1958);
nor U2707 (N_2707,N_2233,N_2379);
nand U2708 (N_2708,N_2348,N_1830);
nor U2709 (N_2709,N_1851,N_2299);
or U2710 (N_2710,N_2188,N_2169);
nor U2711 (N_2711,N_2152,N_2300);
nand U2712 (N_2712,N_2379,N_2345);
and U2713 (N_2713,N_2325,N_1920);
nand U2714 (N_2714,N_2218,N_1885);
nand U2715 (N_2715,N_2124,N_2011);
and U2716 (N_2716,N_2151,N_2365);
and U2717 (N_2717,N_2197,N_1952);
nor U2718 (N_2718,N_2184,N_1909);
or U2719 (N_2719,N_1934,N_2223);
and U2720 (N_2720,N_2065,N_2179);
and U2721 (N_2721,N_2113,N_2298);
nor U2722 (N_2722,N_2334,N_1974);
and U2723 (N_2723,N_2311,N_1965);
nor U2724 (N_2724,N_1902,N_2320);
or U2725 (N_2725,N_2297,N_2097);
and U2726 (N_2726,N_1881,N_2302);
and U2727 (N_2727,N_2020,N_2161);
or U2728 (N_2728,N_1889,N_1972);
nor U2729 (N_2729,N_2237,N_2230);
and U2730 (N_2730,N_2378,N_2034);
nor U2731 (N_2731,N_2225,N_2114);
and U2732 (N_2732,N_2394,N_2131);
nor U2733 (N_2733,N_1855,N_2039);
nor U2734 (N_2734,N_2394,N_2343);
nand U2735 (N_2735,N_2358,N_2073);
nor U2736 (N_2736,N_1836,N_2014);
or U2737 (N_2737,N_1939,N_2330);
nand U2738 (N_2738,N_2272,N_2249);
nand U2739 (N_2739,N_2307,N_1814);
nand U2740 (N_2740,N_1865,N_1964);
nand U2741 (N_2741,N_2301,N_1829);
and U2742 (N_2742,N_1850,N_1821);
and U2743 (N_2743,N_2222,N_2378);
and U2744 (N_2744,N_1940,N_2399);
nor U2745 (N_2745,N_2259,N_2047);
and U2746 (N_2746,N_1928,N_2159);
nand U2747 (N_2747,N_1993,N_1894);
and U2748 (N_2748,N_1811,N_1993);
nor U2749 (N_2749,N_2367,N_1942);
and U2750 (N_2750,N_2254,N_1864);
nor U2751 (N_2751,N_2274,N_1857);
nor U2752 (N_2752,N_1985,N_1856);
nor U2753 (N_2753,N_2203,N_2380);
or U2754 (N_2754,N_2020,N_1848);
nor U2755 (N_2755,N_2399,N_1896);
or U2756 (N_2756,N_2302,N_2280);
and U2757 (N_2757,N_2348,N_2327);
or U2758 (N_2758,N_2036,N_2300);
or U2759 (N_2759,N_1944,N_2008);
or U2760 (N_2760,N_2182,N_2121);
nor U2761 (N_2761,N_1916,N_2268);
nor U2762 (N_2762,N_2194,N_1916);
nand U2763 (N_2763,N_1886,N_2335);
and U2764 (N_2764,N_2240,N_2261);
or U2765 (N_2765,N_1939,N_1935);
or U2766 (N_2766,N_1864,N_2334);
nand U2767 (N_2767,N_1953,N_2136);
xnor U2768 (N_2768,N_2326,N_2078);
and U2769 (N_2769,N_2096,N_2038);
or U2770 (N_2770,N_2251,N_1815);
or U2771 (N_2771,N_2066,N_1814);
nor U2772 (N_2772,N_2143,N_1974);
or U2773 (N_2773,N_2378,N_2096);
nor U2774 (N_2774,N_2005,N_2065);
or U2775 (N_2775,N_2368,N_2364);
nand U2776 (N_2776,N_2262,N_2131);
nor U2777 (N_2777,N_1956,N_2321);
or U2778 (N_2778,N_1960,N_2255);
nor U2779 (N_2779,N_1977,N_1846);
and U2780 (N_2780,N_1887,N_1975);
nor U2781 (N_2781,N_2338,N_2081);
and U2782 (N_2782,N_2288,N_2191);
or U2783 (N_2783,N_2399,N_1974);
nor U2784 (N_2784,N_1916,N_2053);
nor U2785 (N_2785,N_2243,N_2315);
or U2786 (N_2786,N_2336,N_2151);
nor U2787 (N_2787,N_1814,N_1974);
xnor U2788 (N_2788,N_2263,N_2205);
and U2789 (N_2789,N_2346,N_1948);
nor U2790 (N_2790,N_1945,N_2031);
and U2791 (N_2791,N_1971,N_2320);
nor U2792 (N_2792,N_2235,N_2140);
and U2793 (N_2793,N_2389,N_2240);
and U2794 (N_2794,N_2247,N_1919);
nand U2795 (N_2795,N_2248,N_1940);
nor U2796 (N_2796,N_1967,N_2067);
nand U2797 (N_2797,N_1882,N_2171);
and U2798 (N_2798,N_1902,N_2251);
and U2799 (N_2799,N_2016,N_2190);
or U2800 (N_2800,N_1903,N_1803);
xnor U2801 (N_2801,N_2361,N_2396);
nor U2802 (N_2802,N_1933,N_1816);
and U2803 (N_2803,N_2114,N_2279);
nor U2804 (N_2804,N_2130,N_2280);
nor U2805 (N_2805,N_2253,N_2381);
and U2806 (N_2806,N_2178,N_2293);
and U2807 (N_2807,N_2142,N_2258);
or U2808 (N_2808,N_1995,N_2121);
or U2809 (N_2809,N_2264,N_1801);
nor U2810 (N_2810,N_2045,N_2331);
or U2811 (N_2811,N_1803,N_2023);
nand U2812 (N_2812,N_1931,N_2077);
nand U2813 (N_2813,N_2035,N_2278);
and U2814 (N_2814,N_2235,N_2219);
or U2815 (N_2815,N_1910,N_2215);
and U2816 (N_2816,N_1951,N_1962);
nor U2817 (N_2817,N_2132,N_1837);
and U2818 (N_2818,N_2269,N_2198);
or U2819 (N_2819,N_2110,N_2146);
and U2820 (N_2820,N_2011,N_2346);
or U2821 (N_2821,N_2390,N_1985);
nor U2822 (N_2822,N_2304,N_2072);
nor U2823 (N_2823,N_1848,N_2080);
nand U2824 (N_2824,N_1989,N_2327);
nand U2825 (N_2825,N_1968,N_2190);
nor U2826 (N_2826,N_2372,N_1982);
and U2827 (N_2827,N_2228,N_2390);
nor U2828 (N_2828,N_2342,N_2191);
or U2829 (N_2829,N_1904,N_2396);
or U2830 (N_2830,N_2045,N_1962);
nor U2831 (N_2831,N_2369,N_2193);
nor U2832 (N_2832,N_1889,N_1823);
or U2833 (N_2833,N_1977,N_2099);
and U2834 (N_2834,N_2140,N_2237);
nand U2835 (N_2835,N_2385,N_2342);
nor U2836 (N_2836,N_2334,N_2340);
or U2837 (N_2837,N_2167,N_2256);
nor U2838 (N_2838,N_2207,N_2066);
and U2839 (N_2839,N_2132,N_2042);
or U2840 (N_2840,N_1817,N_2207);
and U2841 (N_2841,N_1960,N_1893);
or U2842 (N_2842,N_2000,N_2350);
or U2843 (N_2843,N_2011,N_1953);
nor U2844 (N_2844,N_1808,N_2030);
nor U2845 (N_2845,N_2171,N_2321);
nand U2846 (N_2846,N_2079,N_2121);
nand U2847 (N_2847,N_2275,N_2212);
nand U2848 (N_2848,N_2289,N_1873);
and U2849 (N_2849,N_2089,N_1904);
or U2850 (N_2850,N_2185,N_2341);
or U2851 (N_2851,N_1909,N_2182);
or U2852 (N_2852,N_1946,N_2201);
nand U2853 (N_2853,N_1978,N_1950);
and U2854 (N_2854,N_1818,N_2049);
and U2855 (N_2855,N_2167,N_2298);
or U2856 (N_2856,N_2160,N_2351);
nand U2857 (N_2857,N_2284,N_2252);
and U2858 (N_2858,N_2277,N_2358);
or U2859 (N_2859,N_1947,N_2198);
nand U2860 (N_2860,N_2096,N_2154);
nor U2861 (N_2861,N_1956,N_2250);
nand U2862 (N_2862,N_1838,N_2281);
nor U2863 (N_2863,N_1815,N_2060);
nor U2864 (N_2864,N_1905,N_1902);
nand U2865 (N_2865,N_2080,N_2040);
nor U2866 (N_2866,N_2112,N_2275);
nand U2867 (N_2867,N_2052,N_2225);
nand U2868 (N_2868,N_2026,N_1962);
nor U2869 (N_2869,N_2080,N_2329);
and U2870 (N_2870,N_2019,N_2013);
or U2871 (N_2871,N_2369,N_2299);
nor U2872 (N_2872,N_2208,N_2142);
nor U2873 (N_2873,N_2348,N_1958);
or U2874 (N_2874,N_2131,N_2144);
nor U2875 (N_2875,N_1937,N_2055);
nand U2876 (N_2876,N_2391,N_2290);
xnor U2877 (N_2877,N_2132,N_2167);
nand U2878 (N_2878,N_2182,N_2276);
nand U2879 (N_2879,N_2162,N_1988);
nor U2880 (N_2880,N_2005,N_2018);
or U2881 (N_2881,N_1837,N_1968);
nand U2882 (N_2882,N_2131,N_2024);
or U2883 (N_2883,N_2006,N_1848);
nor U2884 (N_2884,N_1910,N_2200);
nand U2885 (N_2885,N_2392,N_2191);
and U2886 (N_2886,N_2236,N_1853);
nand U2887 (N_2887,N_2028,N_1876);
or U2888 (N_2888,N_2351,N_2238);
or U2889 (N_2889,N_2349,N_2127);
nor U2890 (N_2890,N_2257,N_2265);
and U2891 (N_2891,N_2126,N_2324);
nor U2892 (N_2892,N_2026,N_1991);
and U2893 (N_2893,N_1959,N_1889);
or U2894 (N_2894,N_2308,N_1872);
nand U2895 (N_2895,N_1995,N_2351);
nor U2896 (N_2896,N_2112,N_2297);
nand U2897 (N_2897,N_2287,N_2237);
nor U2898 (N_2898,N_2122,N_1982);
or U2899 (N_2899,N_1959,N_1975);
and U2900 (N_2900,N_1886,N_1923);
or U2901 (N_2901,N_1911,N_2346);
nor U2902 (N_2902,N_2356,N_2341);
nand U2903 (N_2903,N_2163,N_2244);
xor U2904 (N_2904,N_2144,N_2275);
or U2905 (N_2905,N_2175,N_2286);
or U2906 (N_2906,N_1954,N_2194);
nand U2907 (N_2907,N_1859,N_1879);
and U2908 (N_2908,N_2284,N_2214);
and U2909 (N_2909,N_1984,N_1875);
or U2910 (N_2910,N_1971,N_1897);
and U2911 (N_2911,N_2212,N_2011);
nand U2912 (N_2912,N_2124,N_2327);
and U2913 (N_2913,N_1976,N_1945);
and U2914 (N_2914,N_1877,N_1824);
and U2915 (N_2915,N_2196,N_2021);
and U2916 (N_2916,N_1928,N_2135);
and U2917 (N_2917,N_2371,N_2331);
and U2918 (N_2918,N_1887,N_2193);
nand U2919 (N_2919,N_1864,N_2078);
xor U2920 (N_2920,N_2121,N_2194);
or U2921 (N_2921,N_1990,N_1991);
and U2922 (N_2922,N_2351,N_1942);
nand U2923 (N_2923,N_2249,N_2317);
nor U2924 (N_2924,N_1867,N_2069);
nand U2925 (N_2925,N_2055,N_1953);
nand U2926 (N_2926,N_2270,N_2056);
nor U2927 (N_2927,N_1854,N_2181);
nor U2928 (N_2928,N_2280,N_1939);
nor U2929 (N_2929,N_1913,N_1828);
nand U2930 (N_2930,N_2095,N_2310);
and U2931 (N_2931,N_2171,N_1975);
nand U2932 (N_2932,N_2229,N_1958);
or U2933 (N_2933,N_1937,N_1924);
or U2934 (N_2934,N_2348,N_2289);
nand U2935 (N_2935,N_1838,N_2060);
or U2936 (N_2936,N_1951,N_2396);
nor U2937 (N_2937,N_2005,N_2009);
and U2938 (N_2938,N_1916,N_2141);
nor U2939 (N_2939,N_1929,N_2371);
nor U2940 (N_2940,N_2232,N_2253);
nor U2941 (N_2941,N_1893,N_2142);
nand U2942 (N_2942,N_1901,N_2213);
and U2943 (N_2943,N_2339,N_1832);
nor U2944 (N_2944,N_2108,N_1883);
or U2945 (N_2945,N_2027,N_2174);
or U2946 (N_2946,N_2227,N_1970);
nor U2947 (N_2947,N_1908,N_2381);
nand U2948 (N_2948,N_1876,N_1896);
or U2949 (N_2949,N_1890,N_1982);
and U2950 (N_2950,N_2311,N_2011);
nor U2951 (N_2951,N_2224,N_1827);
nor U2952 (N_2952,N_1817,N_2092);
nand U2953 (N_2953,N_1877,N_1825);
and U2954 (N_2954,N_2288,N_2219);
or U2955 (N_2955,N_2267,N_1878);
or U2956 (N_2956,N_2350,N_2267);
nand U2957 (N_2957,N_1942,N_2164);
or U2958 (N_2958,N_2074,N_1800);
nor U2959 (N_2959,N_1842,N_2290);
or U2960 (N_2960,N_2251,N_2370);
nor U2961 (N_2961,N_2256,N_1837);
or U2962 (N_2962,N_2258,N_2257);
nand U2963 (N_2963,N_2113,N_2066);
nand U2964 (N_2964,N_2318,N_1925);
nor U2965 (N_2965,N_1894,N_2326);
nor U2966 (N_2966,N_1911,N_2303);
nor U2967 (N_2967,N_2057,N_2355);
xor U2968 (N_2968,N_1909,N_2227);
or U2969 (N_2969,N_1808,N_1835);
or U2970 (N_2970,N_1816,N_2209);
or U2971 (N_2971,N_2313,N_2195);
nand U2972 (N_2972,N_1897,N_1992);
xor U2973 (N_2973,N_2025,N_2368);
nor U2974 (N_2974,N_2037,N_2277);
or U2975 (N_2975,N_2328,N_2026);
or U2976 (N_2976,N_2201,N_2035);
or U2977 (N_2977,N_2239,N_2134);
nand U2978 (N_2978,N_2144,N_2337);
and U2979 (N_2979,N_2071,N_2080);
or U2980 (N_2980,N_2390,N_2122);
nor U2981 (N_2981,N_2202,N_2339);
and U2982 (N_2982,N_2191,N_1879);
or U2983 (N_2983,N_2041,N_2313);
nor U2984 (N_2984,N_2022,N_1975);
or U2985 (N_2985,N_1971,N_2143);
or U2986 (N_2986,N_2295,N_1818);
or U2987 (N_2987,N_2204,N_2295);
and U2988 (N_2988,N_2027,N_2338);
and U2989 (N_2989,N_2015,N_2225);
and U2990 (N_2990,N_2307,N_2308);
nor U2991 (N_2991,N_2305,N_2333);
and U2992 (N_2992,N_2005,N_1893);
nand U2993 (N_2993,N_1884,N_1869);
nor U2994 (N_2994,N_2103,N_2275);
and U2995 (N_2995,N_1994,N_2350);
and U2996 (N_2996,N_1913,N_2397);
nand U2997 (N_2997,N_2297,N_2323);
and U2998 (N_2998,N_2300,N_1989);
or U2999 (N_2999,N_2247,N_2049);
or UO_0 (O_0,N_2510,N_2995);
nand UO_1 (O_1,N_2984,N_2896);
nand UO_2 (O_2,N_2581,N_2849);
and UO_3 (O_3,N_2658,N_2686);
and UO_4 (O_4,N_2470,N_2821);
and UO_5 (O_5,N_2925,N_2950);
and UO_6 (O_6,N_2722,N_2983);
and UO_7 (O_7,N_2608,N_2412);
or UO_8 (O_8,N_2498,N_2794);
or UO_9 (O_9,N_2446,N_2939);
or UO_10 (O_10,N_2723,N_2952);
or UO_11 (O_11,N_2780,N_2753);
or UO_12 (O_12,N_2543,N_2555);
and UO_13 (O_13,N_2963,N_2974);
and UO_14 (O_14,N_2530,N_2484);
or UO_15 (O_15,N_2724,N_2876);
nand UO_16 (O_16,N_2497,N_2444);
and UO_17 (O_17,N_2519,N_2451);
and UO_18 (O_18,N_2758,N_2852);
or UO_19 (O_19,N_2430,N_2557);
and UO_20 (O_20,N_2871,N_2752);
nand UO_21 (O_21,N_2973,N_2710);
or UO_22 (O_22,N_2874,N_2458);
and UO_23 (O_23,N_2690,N_2568);
or UO_24 (O_24,N_2701,N_2884);
nand UO_25 (O_25,N_2808,N_2540);
nor UO_26 (O_26,N_2728,N_2433);
and UO_27 (O_27,N_2797,N_2570);
or UO_28 (O_28,N_2825,N_2492);
nand UO_29 (O_29,N_2580,N_2861);
and UO_30 (O_30,N_2601,N_2514);
nand UO_31 (O_31,N_2733,N_2404);
or UO_32 (O_32,N_2661,N_2585);
nand UO_33 (O_33,N_2831,N_2979);
and UO_34 (O_34,N_2777,N_2864);
or UO_35 (O_35,N_2562,N_2439);
nand UO_36 (O_36,N_2588,N_2885);
nor UO_37 (O_37,N_2487,N_2746);
nor UO_38 (O_38,N_2897,N_2668);
nand UO_39 (O_39,N_2757,N_2785);
nand UO_40 (O_40,N_2428,N_2842);
nand UO_41 (O_41,N_2857,N_2994);
or UO_42 (O_42,N_2878,N_2517);
nand UO_43 (O_43,N_2845,N_2731);
nand UO_44 (O_44,N_2700,N_2594);
or UO_45 (O_45,N_2415,N_2771);
nor UO_46 (O_46,N_2953,N_2678);
nor UO_47 (O_47,N_2694,N_2649);
and UO_48 (O_48,N_2596,N_2919);
nor UO_49 (O_49,N_2591,N_2932);
nand UO_50 (O_50,N_2991,N_2798);
nor UO_51 (O_51,N_2822,N_2703);
nand UO_52 (O_52,N_2491,N_2511);
and UO_53 (O_53,N_2719,N_2804);
and UO_54 (O_54,N_2559,N_2784);
or UO_55 (O_55,N_2566,N_2403);
nand UO_56 (O_56,N_2469,N_2604);
or UO_57 (O_57,N_2419,N_2704);
or UO_58 (O_58,N_2882,N_2429);
nand UO_59 (O_59,N_2619,N_2706);
nand UO_60 (O_60,N_2781,N_2664);
nor UO_61 (O_61,N_2677,N_2602);
or UO_62 (O_62,N_2667,N_2579);
nand UO_63 (O_63,N_2793,N_2572);
and UO_64 (O_64,N_2740,N_2506);
nand UO_65 (O_65,N_2747,N_2717);
nor UO_66 (O_66,N_2824,N_2598);
nand UO_67 (O_67,N_2900,N_2989);
nand UO_68 (O_68,N_2475,N_2966);
or UO_69 (O_69,N_2502,N_2906);
and UO_70 (O_70,N_2891,N_2676);
or UO_71 (O_71,N_2967,N_2726);
nand UO_72 (O_72,N_2810,N_2448);
nand UO_73 (O_73,N_2571,N_2751);
and UO_74 (O_74,N_2660,N_2818);
and UO_75 (O_75,N_2923,N_2625);
nor UO_76 (O_76,N_2872,N_2956);
or UO_77 (O_77,N_2955,N_2437);
nand UO_78 (O_78,N_2901,N_2600);
or UO_79 (O_79,N_2426,N_2560);
nor UO_80 (O_80,N_2980,N_2858);
nor UO_81 (O_81,N_2563,N_2941);
nand UO_82 (O_82,N_2424,N_2578);
and UO_83 (O_83,N_2464,N_2958);
nor UO_84 (O_84,N_2501,N_2832);
and UO_85 (O_85,N_2815,N_2607);
nor UO_86 (O_86,N_2739,N_2924);
nand UO_87 (O_87,N_2682,N_2637);
and UO_88 (O_88,N_2413,N_2732);
or UO_89 (O_89,N_2800,N_2862);
nand UO_90 (O_90,N_2836,N_2957);
or UO_91 (O_91,N_2536,N_2621);
or UO_92 (O_92,N_2729,N_2802);
and UO_93 (O_93,N_2528,N_2554);
nor UO_94 (O_94,N_2809,N_2453);
nor UO_95 (O_95,N_2814,N_2524);
and UO_96 (O_96,N_2567,N_2406);
and UO_97 (O_97,N_2883,N_2636);
and UO_98 (O_98,N_2848,N_2679);
nor UO_99 (O_99,N_2903,N_2829);
nand UO_100 (O_100,N_2407,N_2480);
or UO_101 (O_101,N_2503,N_2485);
or UO_102 (O_102,N_2665,N_2899);
nand UO_103 (O_103,N_2927,N_2949);
or UO_104 (O_104,N_2541,N_2930);
nand UO_105 (O_105,N_2805,N_2438);
nor UO_106 (O_106,N_2748,N_2975);
or UO_107 (O_107,N_2551,N_2410);
or UO_108 (O_108,N_2811,N_2730);
nand UO_109 (O_109,N_2441,N_2471);
or UO_110 (O_110,N_2847,N_2499);
or UO_111 (O_111,N_2762,N_2855);
nor UO_112 (O_112,N_2655,N_2539);
and UO_113 (O_113,N_2422,N_2614);
or UO_114 (O_114,N_2968,N_2881);
nor UO_115 (O_115,N_2473,N_2945);
xor UO_116 (O_116,N_2738,N_2807);
nand UO_117 (O_117,N_2854,N_2505);
and UO_118 (O_118,N_2529,N_2913);
or UO_119 (O_119,N_2875,N_2918);
or UO_120 (O_120,N_2612,N_2978);
and UO_121 (O_121,N_2662,N_2767);
nor UO_122 (O_122,N_2638,N_2860);
nor UO_123 (O_123,N_2414,N_2546);
and UO_124 (O_124,N_2783,N_2763);
nor UO_125 (O_125,N_2859,N_2709);
or UO_126 (O_126,N_2460,N_2856);
nand UO_127 (O_127,N_2532,N_2666);
or UO_128 (O_128,N_2435,N_2915);
nand UO_129 (O_129,N_2615,N_2795);
nand UO_130 (O_130,N_2477,N_2586);
xor UO_131 (O_131,N_2518,N_2789);
or UO_132 (O_132,N_2630,N_2741);
nor UO_133 (O_133,N_2650,N_2495);
nor UO_134 (O_134,N_2760,N_2486);
or UO_135 (O_135,N_2877,N_2756);
nand UO_136 (O_136,N_2516,N_2909);
nor UO_137 (O_137,N_2712,N_2674);
nand UO_138 (O_138,N_2917,N_2421);
and UO_139 (O_139,N_2489,N_2613);
nor UO_140 (O_140,N_2617,N_2827);
or UO_141 (O_141,N_2961,N_2605);
nand UO_142 (O_142,N_2715,N_2409);
nor UO_143 (O_143,N_2640,N_2670);
nor UO_144 (O_144,N_2669,N_2645);
or UO_145 (O_145,N_2744,N_2773);
and UO_146 (O_146,N_2713,N_2936);
and UO_147 (O_147,N_2754,N_2556);
nand UO_148 (O_148,N_2427,N_2863);
and UO_149 (O_149,N_2445,N_2454);
or UO_150 (O_150,N_2971,N_2931);
or UO_151 (O_151,N_2692,N_2623);
nor UO_152 (O_152,N_2935,N_2500);
or UO_153 (O_153,N_2577,N_2698);
nand UO_154 (O_154,N_2663,N_2902);
nor UO_155 (O_155,N_2592,N_2643);
or UO_156 (O_156,N_2987,N_2998);
or UO_157 (O_157,N_2791,N_2488);
and UO_158 (O_158,N_2926,N_2972);
nor UO_159 (O_159,N_2479,N_2648);
nand UO_160 (O_160,N_2442,N_2766);
nand UO_161 (O_161,N_2436,N_2507);
nand UO_162 (O_162,N_2449,N_2574);
and UO_163 (O_163,N_2622,N_2838);
or UO_164 (O_164,N_2776,N_2887);
or UO_165 (O_165,N_2736,N_2721);
and UO_166 (O_166,N_2850,N_2790);
nor UO_167 (O_167,N_2796,N_2707);
and UO_168 (O_168,N_2764,N_2819);
and UO_169 (O_169,N_2916,N_2558);
nor UO_170 (O_170,N_2472,N_2513);
or UO_171 (O_171,N_2970,N_2779);
nor UO_172 (O_172,N_2531,N_2632);
and UO_173 (O_173,N_2687,N_2944);
and UO_174 (O_174,N_2711,N_2584);
nor UO_175 (O_175,N_2702,N_2631);
or UO_176 (O_176,N_2928,N_2959);
or UO_177 (O_177,N_2914,N_2496);
or UO_178 (O_178,N_2526,N_2629);
nand UO_179 (O_179,N_2801,N_2642);
or UO_180 (O_180,N_2889,N_2985);
and UO_181 (O_181,N_2937,N_2898);
nand UO_182 (O_182,N_2735,N_2583);
or UO_183 (O_183,N_2725,N_2490);
and UO_184 (O_184,N_2634,N_2922);
nor UO_185 (O_185,N_2626,N_2840);
or UO_186 (O_186,N_2737,N_2405);
or UO_187 (O_187,N_2992,N_2853);
and UO_188 (O_188,N_2846,N_2873);
or UO_189 (O_189,N_2569,N_2705);
and UO_190 (O_190,N_2512,N_2755);
nor UO_191 (O_191,N_2651,N_2894);
or UO_192 (O_192,N_2646,N_2673);
or UO_193 (O_193,N_2684,N_2938);
or UO_194 (O_194,N_2675,N_2934);
and UO_195 (O_195,N_2770,N_2504);
nor UO_196 (O_196,N_2590,N_2423);
or UO_197 (O_197,N_2525,N_2474);
or UO_198 (O_198,N_2943,N_2693);
nor UO_199 (O_199,N_2954,N_2450);
and UO_200 (O_200,N_2683,N_2483);
and UO_201 (O_201,N_2467,N_2982);
or UO_202 (O_202,N_2720,N_2522);
nor UO_203 (O_203,N_2787,N_2947);
and UO_204 (O_204,N_2948,N_2830);
or UO_205 (O_205,N_2907,N_2401);
or UO_206 (O_206,N_2879,N_2459);
and UO_207 (O_207,N_2812,N_2549);
nand UO_208 (O_208,N_2657,N_2521);
or UO_209 (O_209,N_2835,N_2716);
nor UO_210 (O_210,N_2465,N_2672);
or UO_211 (O_211,N_2960,N_2988);
nand UO_212 (O_212,N_2603,N_2432);
nand UO_213 (O_213,N_2652,N_2921);
nand UO_214 (O_214,N_2452,N_2759);
nor UO_215 (O_215,N_2624,N_2680);
nor UO_216 (O_216,N_2564,N_2933);
and UO_217 (O_217,N_2886,N_2742);
or UO_218 (O_218,N_2418,N_2696);
nor UO_219 (O_219,N_2527,N_2482);
or UO_220 (O_220,N_2641,N_2494);
and UO_221 (O_221,N_2537,N_2806);
nand UO_222 (O_222,N_2553,N_2695);
nor UO_223 (O_223,N_2476,N_2786);
nand UO_224 (O_224,N_2841,N_2792);
nand UO_225 (O_225,N_2408,N_2691);
and UO_226 (O_226,N_2447,N_2548);
and UO_227 (O_227,N_2538,N_2654);
nand UO_228 (O_228,N_2561,N_2456);
nand UO_229 (O_229,N_2440,N_2964);
and UO_230 (O_230,N_2888,N_2400);
nor UO_231 (O_231,N_2851,N_2828);
or UO_232 (O_232,N_2618,N_2576);
or UO_233 (O_233,N_2969,N_2462);
nand UO_234 (O_234,N_2443,N_2799);
nor UO_235 (O_235,N_2816,N_2813);
nor UO_236 (O_236,N_2547,N_2893);
nor UO_237 (O_237,N_2595,N_2599);
and UO_238 (O_238,N_2425,N_2772);
nor UO_239 (O_239,N_2908,N_2688);
and UO_240 (O_240,N_2761,N_2417);
and UO_241 (O_241,N_2820,N_2627);
and UO_242 (O_242,N_2788,N_2644);
nand UO_243 (O_243,N_2455,N_2823);
nor UO_244 (O_244,N_2544,N_2468);
nor UO_245 (O_245,N_2734,N_2609);
nor UO_246 (O_246,N_2905,N_2911);
and UO_247 (O_247,N_2635,N_2550);
nand UO_248 (O_248,N_2867,N_2671);
nand UO_249 (O_249,N_2610,N_2833);
or UO_250 (O_250,N_2515,N_2545);
nand UO_251 (O_251,N_2466,N_2589);
or UO_252 (O_252,N_2778,N_2892);
or UO_253 (O_253,N_2708,N_2866);
or UO_254 (O_254,N_2699,N_2946);
and UO_255 (O_255,N_2587,N_2996);
nand UO_256 (O_256,N_2434,N_2689);
nor UO_257 (O_257,N_2750,N_2765);
nor UO_258 (O_258,N_2461,N_2837);
and UO_259 (O_259,N_2942,N_2977);
nor UO_260 (O_260,N_2639,N_2880);
nand UO_261 (O_261,N_2951,N_2768);
or UO_262 (O_262,N_2535,N_2520);
or UO_263 (O_263,N_2910,N_2727);
nor UO_264 (O_264,N_2997,N_2993);
or UO_265 (O_265,N_2962,N_2826);
or UO_266 (O_266,N_2478,N_2534);
nor UO_267 (O_267,N_2628,N_2647);
or UO_268 (O_268,N_2573,N_2493);
nor UO_269 (O_269,N_2606,N_2912);
or UO_270 (O_270,N_2745,N_2920);
and UO_271 (O_271,N_2411,N_2775);
nand UO_272 (O_272,N_2714,N_2620);
and UO_273 (O_273,N_2523,N_2633);
or UO_274 (O_274,N_2817,N_2659);
and UO_275 (O_275,N_2681,N_2940);
nand UO_276 (O_276,N_2990,N_2508);
nand UO_277 (O_277,N_2895,N_2769);
nor UO_278 (O_278,N_2976,N_2718);
nor UO_279 (O_279,N_2839,N_2904);
nand UO_280 (O_280,N_2749,N_2774);
or UO_281 (O_281,N_2870,N_2616);
and UO_282 (O_282,N_2868,N_2981);
nand UO_283 (O_283,N_2743,N_2463);
or UO_284 (O_284,N_2533,N_2402);
and UO_285 (O_285,N_2929,N_2843);
nor UO_286 (O_286,N_2431,N_2782);
nand UO_287 (O_287,N_2582,N_2685);
nor UO_288 (O_288,N_2834,N_2965);
nor UO_289 (O_289,N_2697,N_2986);
and UO_290 (O_290,N_2552,N_2416);
or UO_291 (O_291,N_2803,N_2481);
or UO_292 (O_292,N_2656,N_2509);
nand UO_293 (O_293,N_2869,N_2457);
xnor UO_294 (O_294,N_2611,N_2565);
nor UO_295 (O_295,N_2542,N_2844);
and UO_296 (O_296,N_2593,N_2653);
and UO_297 (O_297,N_2575,N_2890);
or UO_298 (O_298,N_2999,N_2420);
nor UO_299 (O_299,N_2597,N_2865);
nand UO_300 (O_300,N_2900,N_2531);
or UO_301 (O_301,N_2406,N_2603);
nor UO_302 (O_302,N_2548,N_2722);
and UO_303 (O_303,N_2654,N_2970);
and UO_304 (O_304,N_2655,N_2473);
nand UO_305 (O_305,N_2643,N_2535);
or UO_306 (O_306,N_2902,N_2830);
nor UO_307 (O_307,N_2568,N_2672);
nor UO_308 (O_308,N_2751,N_2888);
and UO_309 (O_309,N_2815,N_2960);
and UO_310 (O_310,N_2557,N_2597);
and UO_311 (O_311,N_2932,N_2748);
nand UO_312 (O_312,N_2579,N_2643);
or UO_313 (O_313,N_2880,N_2830);
or UO_314 (O_314,N_2402,N_2555);
nand UO_315 (O_315,N_2483,N_2654);
or UO_316 (O_316,N_2894,N_2696);
nand UO_317 (O_317,N_2473,N_2803);
and UO_318 (O_318,N_2936,N_2757);
or UO_319 (O_319,N_2652,N_2419);
nor UO_320 (O_320,N_2498,N_2510);
nor UO_321 (O_321,N_2950,N_2966);
or UO_322 (O_322,N_2904,N_2721);
or UO_323 (O_323,N_2869,N_2463);
xnor UO_324 (O_324,N_2966,N_2946);
nor UO_325 (O_325,N_2485,N_2460);
nand UO_326 (O_326,N_2530,N_2820);
nand UO_327 (O_327,N_2717,N_2550);
nand UO_328 (O_328,N_2521,N_2545);
and UO_329 (O_329,N_2510,N_2872);
nor UO_330 (O_330,N_2594,N_2628);
or UO_331 (O_331,N_2578,N_2439);
nor UO_332 (O_332,N_2822,N_2963);
and UO_333 (O_333,N_2940,N_2961);
nor UO_334 (O_334,N_2604,N_2654);
and UO_335 (O_335,N_2943,N_2771);
nand UO_336 (O_336,N_2683,N_2702);
and UO_337 (O_337,N_2864,N_2836);
and UO_338 (O_338,N_2725,N_2759);
xnor UO_339 (O_339,N_2479,N_2712);
nor UO_340 (O_340,N_2703,N_2893);
and UO_341 (O_341,N_2494,N_2673);
nand UO_342 (O_342,N_2438,N_2753);
nor UO_343 (O_343,N_2727,N_2778);
or UO_344 (O_344,N_2939,N_2807);
or UO_345 (O_345,N_2824,N_2739);
nor UO_346 (O_346,N_2727,N_2546);
nand UO_347 (O_347,N_2598,N_2730);
nand UO_348 (O_348,N_2560,N_2562);
nand UO_349 (O_349,N_2568,N_2505);
nand UO_350 (O_350,N_2751,N_2473);
nor UO_351 (O_351,N_2928,N_2892);
and UO_352 (O_352,N_2465,N_2705);
nand UO_353 (O_353,N_2623,N_2907);
and UO_354 (O_354,N_2483,N_2865);
and UO_355 (O_355,N_2783,N_2507);
and UO_356 (O_356,N_2809,N_2802);
nand UO_357 (O_357,N_2806,N_2714);
nor UO_358 (O_358,N_2429,N_2853);
nand UO_359 (O_359,N_2683,N_2804);
or UO_360 (O_360,N_2424,N_2995);
or UO_361 (O_361,N_2688,N_2964);
or UO_362 (O_362,N_2514,N_2875);
or UO_363 (O_363,N_2516,N_2680);
and UO_364 (O_364,N_2446,N_2403);
or UO_365 (O_365,N_2623,N_2405);
or UO_366 (O_366,N_2857,N_2425);
or UO_367 (O_367,N_2448,N_2983);
nand UO_368 (O_368,N_2849,N_2906);
and UO_369 (O_369,N_2416,N_2640);
nand UO_370 (O_370,N_2784,N_2933);
or UO_371 (O_371,N_2784,N_2807);
nor UO_372 (O_372,N_2714,N_2728);
and UO_373 (O_373,N_2951,N_2771);
or UO_374 (O_374,N_2914,N_2769);
nor UO_375 (O_375,N_2563,N_2918);
nor UO_376 (O_376,N_2522,N_2985);
or UO_377 (O_377,N_2648,N_2466);
nor UO_378 (O_378,N_2533,N_2634);
and UO_379 (O_379,N_2588,N_2967);
and UO_380 (O_380,N_2840,N_2763);
nand UO_381 (O_381,N_2476,N_2986);
or UO_382 (O_382,N_2723,N_2493);
nor UO_383 (O_383,N_2749,N_2631);
nand UO_384 (O_384,N_2800,N_2812);
xor UO_385 (O_385,N_2468,N_2490);
or UO_386 (O_386,N_2853,N_2929);
or UO_387 (O_387,N_2835,N_2552);
nor UO_388 (O_388,N_2836,N_2639);
nor UO_389 (O_389,N_2760,N_2679);
nor UO_390 (O_390,N_2764,N_2922);
nor UO_391 (O_391,N_2879,N_2892);
and UO_392 (O_392,N_2577,N_2883);
nor UO_393 (O_393,N_2794,N_2644);
or UO_394 (O_394,N_2434,N_2479);
nand UO_395 (O_395,N_2736,N_2448);
and UO_396 (O_396,N_2571,N_2688);
and UO_397 (O_397,N_2426,N_2934);
nor UO_398 (O_398,N_2586,N_2442);
nand UO_399 (O_399,N_2657,N_2945);
xor UO_400 (O_400,N_2648,N_2671);
or UO_401 (O_401,N_2574,N_2942);
nand UO_402 (O_402,N_2873,N_2906);
or UO_403 (O_403,N_2746,N_2879);
and UO_404 (O_404,N_2969,N_2817);
nand UO_405 (O_405,N_2696,N_2622);
and UO_406 (O_406,N_2887,N_2655);
nand UO_407 (O_407,N_2547,N_2482);
nand UO_408 (O_408,N_2471,N_2468);
nand UO_409 (O_409,N_2922,N_2864);
nand UO_410 (O_410,N_2465,N_2981);
or UO_411 (O_411,N_2627,N_2562);
nand UO_412 (O_412,N_2443,N_2694);
nand UO_413 (O_413,N_2761,N_2815);
nand UO_414 (O_414,N_2595,N_2802);
or UO_415 (O_415,N_2420,N_2574);
or UO_416 (O_416,N_2726,N_2581);
or UO_417 (O_417,N_2463,N_2518);
or UO_418 (O_418,N_2489,N_2850);
nor UO_419 (O_419,N_2411,N_2625);
or UO_420 (O_420,N_2732,N_2862);
or UO_421 (O_421,N_2959,N_2796);
nand UO_422 (O_422,N_2932,N_2552);
xor UO_423 (O_423,N_2971,N_2417);
or UO_424 (O_424,N_2578,N_2626);
and UO_425 (O_425,N_2919,N_2673);
or UO_426 (O_426,N_2941,N_2686);
or UO_427 (O_427,N_2739,N_2575);
nor UO_428 (O_428,N_2997,N_2649);
nand UO_429 (O_429,N_2948,N_2973);
nand UO_430 (O_430,N_2818,N_2657);
nor UO_431 (O_431,N_2719,N_2575);
or UO_432 (O_432,N_2637,N_2696);
and UO_433 (O_433,N_2862,N_2457);
and UO_434 (O_434,N_2713,N_2673);
nor UO_435 (O_435,N_2772,N_2909);
nor UO_436 (O_436,N_2682,N_2898);
and UO_437 (O_437,N_2506,N_2973);
or UO_438 (O_438,N_2793,N_2960);
or UO_439 (O_439,N_2953,N_2471);
and UO_440 (O_440,N_2426,N_2992);
or UO_441 (O_441,N_2660,N_2604);
nor UO_442 (O_442,N_2664,N_2465);
and UO_443 (O_443,N_2626,N_2765);
nor UO_444 (O_444,N_2407,N_2637);
nor UO_445 (O_445,N_2517,N_2505);
nand UO_446 (O_446,N_2536,N_2681);
nand UO_447 (O_447,N_2463,N_2907);
nor UO_448 (O_448,N_2437,N_2480);
or UO_449 (O_449,N_2924,N_2441);
and UO_450 (O_450,N_2962,N_2516);
nor UO_451 (O_451,N_2475,N_2657);
or UO_452 (O_452,N_2750,N_2824);
nand UO_453 (O_453,N_2838,N_2885);
nand UO_454 (O_454,N_2804,N_2619);
or UO_455 (O_455,N_2532,N_2531);
and UO_456 (O_456,N_2601,N_2528);
or UO_457 (O_457,N_2922,N_2841);
nor UO_458 (O_458,N_2921,N_2697);
nand UO_459 (O_459,N_2480,N_2944);
nor UO_460 (O_460,N_2757,N_2401);
and UO_461 (O_461,N_2638,N_2645);
nor UO_462 (O_462,N_2608,N_2821);
or UO_463 (O_463,N_2990,N_2853);
nand UO_464 (O_464,N_2462,N_2860);
and UO_465 (O_465,N_2687,N_2666);
or UO_466 (O_466,N_2473,N_2949);
nor UO_467 (O_467,N_2590,N_2966);
nor UO_468 (O_468,N_2633,N_2518);
and UO_469 (O_469,N_2628,N_2676);
or UO_470 (O_470,N_2483,N_2760);
or UO_471 (O_471,N_2447,N_2430);
nand UO_472 (O_472,N_2406,N_2878);
and UO_473 (O_473,N_2560,N_2961);
or UO_474 (O_474,N_2939,N_2753);
nand UO_475 (O_475,N_2544,N_2927);
or UO_476 (O_476,N_2563,N_2932);
and UO_477 (O_477,N_2687,N_2657);
and UO_478 (O_478,N_2878,N_2783);
and UO_479 (O_479,N_2657,N_2996);
or UO_480 (O_480,N_2660,N_2866);
nand UO_481 (O_481,N_2455,N_2948);
nor UO_482 (O_482,N_2803,N_2754);
or UO_483 (O_483,N_2732,N_2685);
nor UO_484 (O_484,N_2495,N_2403);
or UO_485 (O_485,N_2426,N_2631);
nand UO_486 (O_486,N_2764,N_2457);
and UO_487 (O_487,N_2756,N_2715);
or UO_488 (O_488,N_2739,N_2756);
nor UO_489 (O_489,N_2862,N_2936);
nand UO_490 (O_490,N_2988,N_2841);
nand UO_491 (O_491,N_2636,N_2474);
nand UO_492 (O_492,N_2668,N_2975);
or UO_493 (O_493,N_2708,N_2486);
nand UO_494 (O_494,N_2482,N_2880);
nor UO_495 (O_495,N_2966,N_2647);
nand UO_496 (O_496,N_2647,N_2676);
and UO_497 (O_497,N_2512,N_2696);
and UO_498 (O_498,N_2508,N_2805);
and UO_499 (O_499,N_2487,N_2433);
endmodule