module basic_1000_10000_1500_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_293,In_865);
xor U1 (N_1,In_366,In_664);
nor U2 (N_2,In_626,In_41);
nand U3 (N_3,In_992,In_152);
nand U4 (N_4,In_808,In_734);
nor U5 (N_5,In_785,In_776);
nor U6 (N_6,In_116,In_662);
nand U7 (N_7,In_264,In_475);
nor U8 (N_8,In_290,In_336);
nand U9 (N_9,In_685,In_476);
nand U10 (N_10,In_781,In_146);
nor U11 (N_11,In_724,In_582);
or U12 (N_12,In_614,In_747);
or U13 (N_13,In_148,In_256);
or U14 (N_14,In_520,In_84);
nand U15 (N_15,In_732,In_139);
xnor U16 (N_16,In_454,In_166);
and U17 (N_17,In_481,In_483);
xor U18 (N_18,In_935,In_187);
nand U19 (N_19,In_10,In_228);
xor U20 (N_20,In_874,In_742);
and U21 (N_21,In_389,In_676);
or U22 (N_22,In_671,In_886);
and U23 (N_23,In_160,In_206);
or U24 (N_24,In_348,In_118);
nand U25 (N_25,In_986,In_912);
xor U26 (N_26,In_119,In_44);
and U27 (N_27,In_409,In_134);
or U28 (N_28,In_815,In_677);
xor U29 (N_29,In_611,In_926);
xnor U30 (N_30,In_461,In_564);
nor U31 (N_31,In_243,In_971);
nor U32 (N_32,In_233,In_385);
xnor U33 (N_33,In_943,In_496);
or U34 (N_34,In_247,In_88);
xnor U35 (N_35,In_4,In_360);
nand U36 (N_36,In_684,In_589);
xor U37 (N_37,In_430,In_32);
and U38 (N_38,In_831,In_258);
xnor U39 (N_39,In_124,In_940);
or U40 (N_40,In_334,In_898);
nand U41 (N_41,In_132,In_601);
nand U42 (N_42,In_39,In_110);
nor U43 (N_43,In_314,In_749);
xor U44 (N_44,In_423,In_996);
xnor U45 (N_45,In_52,In_800);
nand U46 (N_46,In_858,In_463);
and U47 (N_47,In_603,In_79);
or U48 (N_48,In_567,In_445);
or U49 (N_49,In_592,In_566);
or U50 (N_50,In_340,In_809);
or U51 (N_51,In_916,In_449);
nor U52 (N_52,In_299,In_978);
nand U53 (N_53,In_844,In_668);
and U54 (N_54,In_920,In_543);
and U55 (N_55,In_377,In_770);
or U56 (N_56,In_534,In_536);
and U57 (N_57,In_472,In_591);
xnor U58 (N_58,In_94,In_801);
nand U59 (N_59,In_876,In_194);
or U60 (N_60,In_437,In_99);
nand U61 (N_61,In_200,In_939);
and U62 (N_62,In_38,In_261);
or U63 (N_63,In_300,In_530);
nor U64 (N_64,In_689,In_833);
nand U65 (N_65,In_414,In_165);
nand U66 (N_66,In_362,In_140);
or U67 (N_67,In_594,In_549);
xor U68 (N_68,In_904,In_917);
or U69 (N_69,In_87,In_954);
nor U70 (N_70,In_524,In_315);
and U71 (N_71,In_238,In_184);
nand U72 (N_72,In_251,In_861);
nand U73 (N_73,In_688,In_379);
nand U74 (N_74,In_304,In_620);
xor U75 (N_75,In_108,In_448);
nand U76 (N_76,In_806,In_307);
or U77 (N_77,In_205,In_55);
and U78 (N_78,In_846,In_380);
nand U79 (N_79,In_548,In_95);
nand U80 (N_80,In_777,In_623);
nand U81 (N_81,In_695,In_827);
nor U82 (N_82,In_398,In_284);
xnor U83 (N_83,In_637,In_85);
and U84 (N_84,In_973,In_487);
and U85 (N_85,In_521,In_835);
or U86 (N_86,In_97,In_525);
and U87 (N_87,In_422,In_590);
nand U88 (N_88,In_696,In_608);
or U89 (N_89,In_753,In_186);
or U90 (N_90,In_675,In_965);
nand U91 (N_91,In_416,In_242);
nand U92 (N_92,In_378,In_817);
and U93 (N_93,In_367,In_830);
or U94 (N_94,In_425,In_149);
nor U95 (N_95,In_743,In_927);
or U96 (N_96,In_999,In_646);
nand U97 (N_97,In_259,In_473);
nor U98 (N_98,In_80,In_26);
or U99 (N_99,In_498,In_225);
nand U100 (N_100,In_829,In_931);
or U101 (N_101,In_474,In_232);
and U102 (N_102,In_673,In_308);
or U103 (N_103,In_640,In_419);
or U104 (N_104,In_75,In_432);
or U105 (N_105,In_453,In_945);
xnor U106 (N_106,In_539,In_136);
or U107 (N_107,In_352,In_23);
xor U108 (N_108,In_174,In_182);
and U109 (N_109,In_899,In_459);
or U110 (N_110,In_62,In_515);
or U111 (N_111,In_370,In_579);
xor U112 (N_112,In_735,In_224);
xor U113 (N_113,In_36,In_762);
xnor U114 (N_114,In_153,In_993);
or U115 (N_115,In_410,In_504);
and U116 (N_116,In_848,In_460);
nand U117 (N_117,In_491,In_540);
nand U118 (N_118,In_550,In_244);
and U119 (N_119,In_654,In_83);
xor U120 (N_120,In_201,In_330);
nand U121 (N_121,In_68,In_934);
nand U122 (N_122,In_114,In_871);
or U123 (N_123,In_960,In_823);
nand U124 (N_124,In_514,In_435);
and U125 (N_125,In_740,In_839);
nor U126 (N_126,In_207,In_665);
nor U127 (N_127,In_127,In_910);
nand U128 (N_128,In_17,In_404);
nand U129 (N_129,In_782,In_131);
and U130 (N_130,In_57,In_292);
or U131 (N_131,In_164,In_928);
and U132 (N_132,In_130,In_730);
xnor U133 (N_133,In_546,In_138);
and U134 (N_134,In_947,In_885);
or U135 (N_135,In_209,In_884);
xnor U136 (N_136,In_101,In_325);
nand U137 (N_137,In_451,In_249);
nor U138 (N_138,In_587,In_621);
nand U139 (N_139,In_499,In_368);
and U140 (N_140,In_911,In_576);
or U141 (N_141,In_107,In_253);
xor U142 (N_142,In_531,In_226);
xor U143 (N_143,In_826,In_706);
or U144 (N_144,In_528,In_652);
nor U145 (N_145,In_275,In_157);
nor U146 (N_146,In_838,In_317);
nand U147 (N_147,In_558,In_485);
xnor U148 (N_148,In_736,In_63);
and U149 (N_149,In_755,In_778);
nand U150 (N_150,In_220,In_758);
nor U151 (N_151,In_70,In_78);
or U152 (N_152,In_533,In_418);
xor U153 (N_153,In_89,In_252);
xnor U154 (N_154,In_512,In_875);
xor U155 (N_155,In_745,In_272);
nand U156 (N_156,In_22,In_371);
xor U157 (N_157,In_807,In_399);
and U158 (N_158,In_143,In_958);
nor U159 (N_159,In_922,In_6);
xnor U160 (N_160,In_738,In_37);
xor U161 (N_161,In_211,In_704);
nor U162 (N_162,In_909,In_105);
or U163 (N_163,In_480,In_431);
xnor U164 (N_164,In_163,In_634);
nor U165 (N_165,In_698,In_810);
nor U166 (N_166,In_599,In_343);
nand U167 (N_167,In_661,In_267);
or U168 (N_168,In_401,In_386);
nor U169 (N_169,In_56,In_310);
nor U170 (N_170,In_741,In_277);
xor U171 (N_171,In_622,In_507);
nand U172 (N_172,In_218,In_667);
or U173 (N_173,In_705,In_361);
nor U174 (N_174,In_772,In_718);
and U175 (N_175,In_168,In_880);
or U176 (N_176,In_649,In_250);
nand U177 (N_177,In_725,In_557);
or U178 (N_178,In_11,In_245);
nand U179 (N_179,In_113,In_702);
nand U180 (N_180,In_175,In_337);
xnor U181 (N_181,In_50,In_853);
or U182 (N_182,In_509,In_321);
nor U183 (N_183,In_683,In_632);
and U184 (N_184,In_586,In_851);
and U185 (N_185,In_612,In_331);
nand U186 (N_186,In_535,In_638);
or U187 (N_187,In_906,In_873);
nor U188 (N_188,In_471,In_279);
or U189 (N_189,In_301,In_902);
nor U190 (N_190,In_703,In_998);
or U191 (N_191,In_881,In_584);
xnor U192 (N_192,In_47,In_426);
xnor U193 (N_193,In_952,In_135);
nor U194 (N_194,In_505,In_574);
nor U195 (N_195,In_411,In_71);
xnor U196 (N_196,In_191,In_221);
or U197 (N_197,In_774,In_417);
or U198 (N_198,In_752,In_790);
nor U199 (N_199,In_767,In_276);
nand U200 (N_200,In_494,In_890);
xnor U201 (N_201,In_151,In_670);
and U202 (N_202,In_964,In_158);
or U203 (N_203,In_439,In_568);
and U204 (N_204,In_651,In_588);
nand U205 (N_205,In_322,In_511);
xor U206 (N_206,In_7,In_571);
or U207 (N_207,In_493,In_298);
and U208 (N_208,In_400,In_388);
nand U209 (N_209,In_222,In_856);
and U210 (N_210,In_270,In_636);
nor U211 (N_211,In_722,In_102);
xor U212 (N_212,In_553,In_30);
and U213 (N_213,In_181,In_193);
xnor U214 (N_214,In_488,In_605);
nor U215 (N_215,In_365,In_983);
xnor U216 (N_216,In_721,In_763);
nor U217 (N_217,In_440,In_77);
nor U218 (N_218,In_679,In_8);
nand U219 (N_219,In_223,In_739);
or U220 (N_220,In_561,In_748);
and U221 (N_221,In_953,In_374);
nor U222 (N_222,In_674,In_639);
and U223 (N_223,In_1,In_822);
nor U224 (N_224,In_771,In_708);
and U225 (N_225,In_345,In_74);
nand U226 (N_226,In_754,In_396);
nor U227 (N_227,In_92,In_759);
nand U228 (N_228,In_756,In_457);
nand U229 (N_229,In_66,In_645);
or U230 (N_230,In_484,In_342);
or U231 (N_231,In_901,In_968);
and U232 (N_232,In_860,In_693);
nand U233 (N_233,In_936,In_537);
and U234 (N_234,In_797,In_845);
and U235 (N_235,In_358,In_659);
nand U236 (N_236,In_470,In_58);
and U237 (N_237,In_982,In_333);
nor U238 (N_238,In_492,In_610);
nand U239 (N_239,In_268,In_692);
nand U240 (N_240,In_593,In_699);
and U241 (N_241,In_779,In_580);
xnor U242 (N_242,In_13,In_327);
and U243 (N_243,In_849,In_145);
nor U244 (N_244,In_604,In_289);
nor U245 (N_245,In_510,In_828);
or U246 (N_246,In_554,In_857);
and U247 (N_247,In_644,In_231);
or U248 (N_248,In_443,In_282);
nand U249 (N_249,In_569,In_522);
nor U250 (N_250,In_794,In_274);
and U251 (N_251,In_892,In_918);
and U252 (N_252,In_286,In_517);
xnor U253 (N_253,In_20,In_64);
and U254 (N_254,In_96,In_323);
nor U255 (N_255,In_204,In_29);
xor U256 (N_256,In_458,In_691);
nand U257 (N_257,In_598,In_43);
and U258 (N_258,In_196,In_183);
xor U259 (N_259,In_479,In_864);
nand U260 (N_260,In_951,In_281);
nor U261 (N_261,In_962,In_847);
or U262 (N_262,In_981,In_93);
or U263 (N_263,In_650,In_570);
nand U264 (N_264,In_188,In_316);
nor U265 (N_265,In_328,In_681);
or U266 (N_266,In_82,In_229);
and U267 (N_267,In_320,In_585);
xnor U268 (N_268,In_424,In_375);
or U269 (N_269,In_834,In_489);
nor U270 (N_270,In_16,In_643);
or U271 (N_271,In_825,In_841);
xnor U272 (N_272,In_803,In_869);
xor U273 (N_273,In_581,In_477);
nand U274 (N_274,In_719,In_545);
or U275 (N_275,In_295,In_761);
or U276 (N_276,In_556,In_987);
or U277 (N_277,In_497,In_2);
xnor U278 (N_278,In_628,In_609);
or U279 (N_279,In_773,In_508);
or U280 (N_280,In_59,In_867);
or U281 (N_281,In_167,In_98);
xor U282 (N_282,In_359,In_516);
and U283 (N_283,In_429,In_957);
nor U284 (N_284,In_805,In_120);
xor U285 (N_285,In_527,In_271);
nor U286 (N_286,In_210,In_905);
xnor U287 (N_287,In_583,In_816);
and U288 (N_288,In_929,In_769);
xnor U289 (N_289,In_544,In_121);
nand U290 (N_290,In_248,In_783);
or U291 (N_291,In_112,In_67);
nor U292 (N_292,In_596,In_789);
xor U293 (N_293,In_387,In_811);
or U294 (N_294,In_446,In_467);
xor U295 (N_295,In_888,In_879);
xnor U296 (N_296,In_40,In_538);
nor U297 (N_297,In_280,In_0);
nand U298 (N_298,In_447,In_560);
and U299 (N_299,In_859,In_933);
nand U300 (N_300,In_788,In_716);
or U301 (N_301,In_91,In_324);
and U302 (N_302,In_117,In_441);
or U303 (N_303,In_393,In_737);
or U304 (N_304,In_214,In_103);
nand U305 (N_305,In_176,In_697);
nor U306 (N_306,In_278,In_390);
nand U307 (N_307,In_713,In_791);
xnor U308 (N_308,In_296,In_921);
nor U309 (N_309,In_73,In_21);
xnor U310 (N_310,In_764,In_995);
or U311 (N_311,In_802,In_12);
or U312 (N_312,In_969,In_14);
nor U313 (N_313,In_642,In_893);
and U314 (N_314,In_9,In_565);
xor U315 (N_315,In_500,In_372);
nor U316 (N_316,In_989,In_376);
xnor U317 (N_317,In_635,In_624);
nor U318 (N_318,In_452,In_555);
and U319 (N_319,In_616,In_208);
nand U320 (N_320,In_395,In_33);
nand U321 (N_321,In_700,In_701);
nand U322 (N_322,In_519,In_819);
or U323 (N_323,In_990,In_541);
xnor U324 (N_324,In_949,In_887);
or U325 (N_325,In_24,In_924);
nand U326 (N_326,In_751,In_364);
or U327 (N_327,In_775,In_518);
nor U328 (N_328,In_963,In_547);
nor U329 (N_329,In_273,In_154);
or U330 (N_330,In_302,In_818);
nand U331 (N_331,In_311,In_227);
nand U332 (N_332,In_144,In_728);
nor U333 (N_333,In_100,In_469);
nor U334 (N_334,In_180,In_746);
nand U335 (N_335,In_678,In_353);
xor U336 (N_336,In_397,In_607);
xor U337 (N_337,In_656,In_950);
or U338 (N_338,In_723,In_903);
or U339 (N_339,In_234,In_559);
and U340 (N_340,In_69,In_572);
xor U341 (N_341,In_263,In_687);
xnor U342 (N_342,In_850,In_796);
nor U343 (N_343,In_382,In_217);
and U344 (N_344,In_680,In_198);
nor U345 (N_345,In_672,In_54);
xnor U346 (N_346,In_402,In_313);
nand U347 (N_347,In_919,In_914);
xnor U348 (N_348,In_595,In_147);
nor U349 (N_349,In_717,In_798);
nor U350 (N_350,In_821,In_991);
xor U351 (N_351,In_551,In_937);
or U352 (N_352,In_161,In_897);
and U353 (N_353,In_31,In_303);
or U354 (N_354,In_562,In_465);
or U355 (N_355,In_578,In_765);
or U356 (N_356,In_141,In_563);
and U357 (N_357,In_197,In_820);
nand U358 (N_358,In_237,In_655);
nor U359 (N_359,In_294,In_177);
nand U360 (N_360,In_466,In_339);
xnor U361 (N_361,In_363,In_335);
nand U362 (N_362,In_240,In_959);
and U363 (N_363,In_970,In_369);
or U364 (N_364,In_173,In_438);
and U365 (N_365,In_529,In_72);
nand U366 (N_366,In_215,In_955);
nand U367 (N_367,In_686,In_883);
nor U368 (N_368,In_889,In_600);
xor U369 (N_369,In_49,In_666);
xnor U370 (N_370,In_941,In_486);
nand U371 (N_371,In_795,In_577);
or U372 (N_372,In_641,In_625);
or U373 (N_373,In_285,In_236);
xnor U374 (N_374,In_5,In_915);
nor U375 (N_375,In_442,In_766);
and U376 (N_376,In_552,In_450);
nand U377 (N_377,In_944,In_854);
nand U378 (N_378,In_878,In_35);
and U379 (N_379,In_254,In_150);
xnor U380 (N_380,In_908,In_757);
and U381 (N_381,In_413,In_109);
and U382 (N_382,In_506,In_750);
nand U383 (N_383,In_162,In_309);
or U384 (N_384,In_428,In_61);
or U385 (N_385,In_46,In_977);
or U386 (N_386,In_42,In_714);
or U387 (N_387,In_51,In_633);
nor U388 (N_388,In_824,In_48);
or U389 (N_389,In_630,In_495);
nor U390 (N_390,In_606,In_235);
or U391 (N_391,In_265,In_669);
nor U392 (N_392,In_171,In_357);
nor U393 (N_393,In_354,In_255);
xnor U394 (N_394,In_356,In_690);
nand U395 (N_395,In_142,In_925);
xnor U396 (N_396,In_532,In_111);
nor U397 (N_397,In_203,In_573);
xnor U398 (N_398,In_329,In_408);
nor U399 (N_399,In_349,In_710);
and U400 (N_400,In_351,In_852);
nand U401 (N_401,In_170,In_122);
nor U402 (N_402,In_870,In_60);
and U403 (N_403,In_384,In_837);
or U404 (N_404,In_726,In_976);
xnor U405 (N_405,In_287,In_169);
and U406 (N_406,In_974,In_312);
or U407 (N_407,In_597,In_305);
or U408 (N_408,In_25,In_421);
or U409 (N_409,In_988,In_799);
nor U410 (N_410,In_90,In_895);
nor U411 (N_411,In_502,In_219);
nor U412 (N_412,In_381,In_863);
nor U413 (N_413,In_709,In_104);
xor U414 (N_414,In_15,In_985);
xor U415 (N_415,In_694,In_731);
and U416 (N_416,In_478,In_972);
and U417 (N_417,In_464,In_729);
nand U418 (N_418,In_900,In_266);
nand U419 (N_419,In_980,In_288);
nand U420 (N_420,In_283,In_629);
or U421 (N_421,In_787,In_383);
xor U422 (N_422,In_185,In_786);
nor U423 (N_423,In_436,In_456);
and U424 (N_424,In_882,In_123);
and U425 (N_425,In_602,In_804);
and U426 (N_426,In_179,In_427);
and U427 (N_427,In_760,In_269);
xor U428 (N_428,In_202,In_979);
xnor U429 (N_429,In_462,In_866);
nand U430 (N_430,In_3,In_523);
nand U431 (N_431,In_45,In_468);
or U432 (N_432,In_840,In_246);
nor U433 (N_433,In_613,In_923);
nor U434 (N_434,In_542,In_780);
nor U435 (N_435,In_19,In_326);
and U436 (N_436,In_894,In_28);
nand U437 (N_437,In_913,In_297);
nor U438 (N_438,In_18,In_793);
xnor U439 (N_439,In_712,In_407);
xnor U440 (N_440,In_813,In_733);
and U441 (N_441,In_347,In_199);
and U442 (N_442,In_355,In_997);
xnor U443 (N_443,In_619,In_129);
or U444 (N_444,In_420,In_501);
and U445 (N_445,In_872,In_156);
nand U446 (N_446,In_86,In_34);
or U447 (N_447,In_27,In_930);
nor U448 (N_448,In_373,In_412);
nor U449 (N_449,In_455,In_291);
or U450 (N_450,In_956,In_653);
nor U451 (N_451,In_812,In_53);
or U452 (N_452,In_126,In_482);
nor U453 (N_453,In_332,In_306);
xor U454 (N_454,In_444,In_192);
or U455 (N_455,In_260,In_338);
xnor U456 (N_456,In_946,In_784);
nor U457 (N_457,In_896,In_115);
xor U458 (N_458,In_216,In_682);
nand U459 (N_459,In_125,In_526);
nor U460 (N_460,In_832,In_189);
xor U461 (N_461,In_257,In_647);
nand U462 (N_462,In_660,In_907);
or U463 (N_463,In_975,In_575);
xnor U464 (N_464,In_615,In_212);
nor U465 (N_465,In_618,In_137);
nand U466 (N_466,In_262,In_513);
nand U467 (N_467,In_942,In_961);
nand U468 (N_468,In_391,In_344);
or U469 (N_469,In_346,In_938);
xnor U470 (N_470,In_877,In_155);
nand U471 (N_471,In_843,In_792);
or U472 (N_472,In_648,In_631);
xnor U473 (N_473,In_241,In_128);
nand U474 (N_474,In_862,In_663);
nor U475 (N_475,In_403,In_213);
xor U476 (N_476,In_172,In_842);
and U477 (N_477,In_868,In_503);
and U478 (N_478,In_727,In_658);
and U479 (N_479,In_392,In_178);
nor U480 (N_480,In_190,In_715);
and U481 (N_481,In_627,In_490);
nand U482 (N_482,In_984,In_350);
nor U483 (N_483,In_707,In_891);
xor U484 (N_484,In_967,In_81);
nand U485 (N_485,In_768,In_433);
or U486 (N_486,In_711,In_814);
nand U487 (N_487,In_133,In_239);
and U488 (N_488,In_394,In_434);
or U489 (N_489,In_159,In_966);
xor U490 (N_490,In_836,In_318);
xor U491 (N_491,In_341,In_319);
nor U492 (N_492,In_106,In_195);
nand U493 (N_493,In_415,In_932);
xnor U494 (N_494,In_855,In_720);
and U495 (N_495,In_406,In_65);
and U496 (N_496,In_948,In_617);
or U497 (N_497,In_230,In_76);
xnor U498 (N_498,In_744,In_994);
nand U499 (N_499,In_657,In_405);
or U500 (N_500,N_165,N_310);
nand U501 (N_501,N_155,N_283);
nor U502 (N_502,N_59,N_352);
nand U503 (N_503,N_280,N_487);
nor U504 (N_504,N_403,N_319);
and U505 (N_505,N_435,N_169);
nor U506 (N_506,N_253,N_323);
xnor U507 (N_507,N_249,N_190);
nor U508 (N_508,N_57,N_274);
and U509 (N_509,N_410,N_95);
nand U510 (N_510,N_245,N_206);
xnor U511 (N_511,N_121,N_246);
xor U512 (N_512,N_90,N_474);
nor U513 (N_513,N_378,N_259);
nand U514 (N_514,N_480,N_45);
nor U515 (N_515,N_127,N_458);
nand U516 (N_516,N_63,N_294);
or U517 (N_517,N_203,N_463);
xnor U518 (N_518,N_252,N_176);
and U519 (N_519,N_147,N_402);
and U520 (N_520,N_178,N_390);
and U521 (N_521,N_193,N_198);
nand U522 (N_522,N_207,N_51);
or U523 (N_523,N_243,N_142);
nor U524 (N_524,N_264,N_483);
nand U525 (N_525,N_247,N_391);
xor U526 (N_526,N_301,N_67);
or U527 (N_527,N_419,N_236);
and U528 (N_528,N_71,N_156);
or U529 (N_529,N_369,N_132);
and U530 (N_530,N_96,N_192);
and U531 (N_531,N_314,N_5);
or U532 (N_532,N_262,N_111);
xor U533 (N_533,N_332,N_489);
xnor U534 (N_534,N_9,N_381);
xnor U535 (N_535,N_20,N_105);
nor U536 (N_536,N_337,N_285);
xor U537 (N_537,N_490,N_197);
or U538 (N_538,N_358,N_226);
and U539 (N_539,N_414,N_467);
or U540 (N_540,N_231,N_129);
and U541 (N_541,N_189,N_360);
nand U542 (N_542,N_37,N_106);
nand U543 (N_543,N_290,N_154);
xor U544 (N_544,N_386,N_224);
nand U545 (N_545,N_89,N_72);
nor U546 (N_546,N_284,N_309);
xnor U547 (N_547,N_327,N_199);
xnor U548 (N_548,N_44,N_49);
or U549 (N_549,N_135,N_196);
or U550 (N_550,N_346,N_240);
nand U551 (N_551,N_65,N_394);
nor U552 (N_552,N_366,N_424);
and U553 (N_553,N_216,N_422);
or U554 (N_554,N_218,N_3);
nor U555 (N_555,N_19,N_244);
and U556 (N_556,N_382,N_70);
xnor U557 (N_557,N_279,N_343);
nand U558 (N_558,N_449,N_174);
and U559 (N_559,N_282,N_82);
xor U560 (N_560,N_40,N_361);
or U561 (N_561,N_173,N_324);
nand U562 (N_562,N_87,N_433);
or U563 (N_563,N_325,N_357);
nor U564 (N_564,N_320,N_136);
nand U565 (N_565,N_408,N_377);
or U566 (N_566,N_116,N_184);
nor U567 (N_567,N_98,N_450);
nand U568 (N_568,N_340,N_81);
and U569 (N_569,N_229,N_370);
and U570 (N_570,N_263,N_373);
nand U571 (N_571,N_148,N_80);
xnor U572 (N_572,N_304,N_493);
and U573 (N_573,N_462,N_146);
and U574 (N_574,N_430,N_34);
nand U575 (N_575,N_115,N_163);
nand U576 (N_576,N_302,N_441);
nand U577 (N_577,N_478,N_428);
or U578 (N_578,N_261,N_36);
nor U579 (N_579,N_125,N_268);
or U580 (N_580,N_260,N_112);
nand U581 (N_581,N_418,N_191);
nand U582 (N_582,N_464,N_482);
or U583 (N_583,N_102,N_440);
xnor U584 (N_584,N_238,N_496);
and U585 (N_585,N_141,N_210);
xor U586 (N_586,N_251,N_123);
nor U587 (N_587,N_398,N_442);
nand U588 (N_588,N_322,N_257);
nor U589 (N_589,N_367,N_446);
or U590 (N_590,N_383,N_103);
nand U591 (N_591,N_432,N_14);
xor U592 (N_592,N_33,N_491);
nand U593 (N_593,N_300,N_421);
xor U594 (N_594,N_56,N_328);
nand U595 (N_595,N_372,N_120);
or U596 (N_596,N_177,N_131);
xor U597 (N_597,N_270,N_88);
nand U598 (N_598,N_488,N_312);
or U599 (N_599,N_25,N_341);
and U600 (N_600,N_338,N_269);
and U601 (N_601,N_273,N_35);
and U602 (N_602,N_461,N_393);
xor U603 (N_603,N_318,N_472);
or U604 (N_604,N_291,N_27);
or U605 (N_605,N_371,N_17);
and U606 (N_606,N_50,N_151);
and U607 (N_607,N_456,N_93);
or U608 (N_608,N_139,N_75);
nand U609 (N_609,N_21,N_172);
xnor U610 (N_610,N_401,N_94);
nand U611 (N_611,N_362,N_99);
nor U612 (N_612,N_448,N_62);
xor U613 (N_613,N_454,N_91);
xnor U614 (N_614,N_438,N_437);
and U615 (N_615,N_219,N_230);
nor U616 (N_616,N_481,N_215);
nor U617 (N_617,N_277,N_466);
nor U618 (N_618,N_321,N_473);
xor U619 (N_619,N_188,N_335);
nor U620 (N_620,N_258,N_355);
or U621 (N_621,N_256,N_363);
xor U622 (N_622,N_375,N_315);
xor U623 (N_623,N_234,N_134);
nor U624 (N_624,N_468,N_73);
and U625 (N_625,N_159,N_168);
xor U626 (N_626,N_164,N_39);
or U627 (N_627,N_232,N_429);
or U628 (N_628,N_186,N_201);
or U629 (N_629,N_347,N_162);
or U630 (N_630,N_133,N_104);
or U631 (N_631,N_223,N_225);
or U632 (N_632,N_417,N_109);
and U633 (N_633,N_306,N_113);
or U634 (N_634,N_145,N_143);
nand U635 (N_635,N_356,N_431);
or U636 (N_636,N_167,N_166);
or U637 (N_637,N_118,N_475);
xor U638 (N_638,N_406,N_157);
and U639 (N_639,N_101,N_384);
nand U640 (N_640,N_353,N_329);
xor U641 (N_641,N_298,N_160);
nand U642 (N_642,N_439,N_110);
nor U643 (N_643,N_211,N_122);
nor U644 (N_644,N_497,N_470);
nor U645 (N_645,N_11,N_15);
and U646 (N_646,N_344,N_60);
or U647 (N_647,N_333,N_30);
xor U648 (N_648,N_426,N_427);
nor U649 (N_649,N_77,N_465);
nor U650 (N_650,N_107,N_479);
xnor U651 (N_651,N_239,N_492);
and U652 (N_652,N_313,N_179);
or U653 (N_653,N_425,N_46);
nor U654 (N_654,N_486,N_287);
nor U655 (N_655,N_235,N_7);
and U656 (N_656,N_255,N_214);
nand U657 (N_657,N_4,N_183);
or U658 (N_658,N_52,N_222);
nor U659 (N_659,N_237,N_451);
nor U660 (N_660,N_365,N_228);
nor U661 (N_661,N_220,N_434);
nor U662 (N_662,N_185,N_68);
and U663 (N_663,N_275,N_117);
or U664 (N_664,N_387,N_296);
or U665 (N_665,N_350,N_175);
and U666 (N_666,N_209,N_108);
nor U667 (N_667,N_385,N_217);
nor U668 (N_668,N_477,N_484);
nor U669 (N_669,N_409,N_376);
and U670 (N_670,N_18,N_368);
xnor U671 (N_671,N_396,N_295);
or U672 (N_672,N_364,N_158);
or U673 (N_673,N_92,N_303);
nor U674 (N_674,N_420,N_380);
xnor U675 (N_675,N_171,N_140);
or U676 (N_676,N_42,N_86);
or U677 (N_677,N_1,N_399);
and U678 (N_678,N_161,N_276);
xnor U679 (N_679,N_307,N_311);
and U680 (N_680,N_359,N_374);
nor U681 (N_681,N_130,N_289);
and U682 (N_682,N_61,N_221);
xor U683 (N_683,N_6,N_316);
nor U684 (N_684,N_28,N_469);
nand U685 (N_685,N_202,N_308);
or U686 (N_686,N_31,N_345);
and U687 (N_687,N_12,N_348);
xor U688 (N_688,N_476,N_413);
or U689 (N_689,N_455,N_248);
xor U690 (N_690,N_153,N_227);
nand U691 (N_691,N_305,N_389);
nand U692 (N_692,N_137,N_55);
or U693 (N_693,N_459,N_293);
nor U694 (N_694,N_411,N_85);
nand U695 (N_695,N_242,N_397);
and U696 (N_696,N_471,N_64);
or U697 (N_697,N_292,N_299);
nand U698 (N_698,N_445,N_460);
or U699 (N_699,N_286,N_412);
xor U700 (N_700,N_495,N_187);
nand U701 (N_701,N_79,N_330);
nor U702 (N_702,N_498,N_213);
or U703 (N_703,N_22,N_0);
or U704 (N_704,N_48,N_233);
xor U705 (N_705,N_41,N_443);
nand U706 (N_706,N_392,N_97);
nand U707 (N_707,N_78,N_76);
nor U708 (N_708,N_388,N_204);
nor U709 (N_709,N_212,N_26);
or U710 (N_710,N_181,N_485);
nand U711 (N_711,N_453,N_317);
and U712 (N_712,N_271,N_278);
nand U713 (N_713,N_200,N_24);
or U714 (N_714,N_250,N_334);
or U715 (N_715,N_288,N_114);
and U716 (N_716,N_152,N_342);
or U717 (N_717,N_195,N_66);
and U718 (N_718,N_53,N_10);
nor U719 (N_719,N_241,N_128);
xor U720 (N_720,N_8,N_349);
and U721 (N_721,N_336,N_43);
xnor U722 (N_722,N_119,N_149);
and U723 (N_723,N_170,N_180);
nand U724 (N_724,N_54,N_23);
and U725 (N_725,N_150,N_272);
nand U726 (N_726,N_416,N_400);
and U727 (N_727,N_144,N_379);
xnor U728 (N_728,N_124,N_208);
or U729 (N_729,N_84,N_447);
xor U730 (N_730,N_205,N_407);
xnor U731 (N_731,N_13,N_58);
nor U732 (N_732,N_297,N_100);
or U733 (N_733,N_405,N_444);
and U734 (N_734,N_47,N_326);
or U735 (N_735,N_404,N_16);
xor U736 (N_736,N_83,N_499);
xnor U737 (N_737,N_452,N_194);
and U738 (N_738,N_415,N_69);
nor U739 (N_739,N_182,N_423);
nand U740 (N_740,N_138,N_29);
nand U741 (N_741,N_126,N_331);
nand U742 (N_742,N_436,N_267);
or U743 (N_743,N_351,N_281);
xnor U744 (N_744,N_354,N_254);
nand U745 (N_745,N_339,N_32);
nand U746 (N_746,N_266,N_494);
nand U747 (N_747,N_395,N_2);
nor U748 (N_748,N_38,N_457);
nand U749 (N_749,N_265,N_74);
and U750 (N_750,N_489,N_316);
and U751 (N_751,N_315,N_402);
or U752 (N_752,N_398,N_452);
nand U753 (N_753,N_14,N_35);
nor U754 (N_754,N_23,N_450);
and U755 (N_755,N_137,N_179);
nand U756 (N_756,N_325,N_59);
xor U757 (N_757,N_138,N_170);
xor U758 (N_758,N_22,N_157);
and U759 (N_759,N_303,N_78);
nand U760 (N_760,N_417,N_75);
nand U761 (N_761,N_420,N_361);
or U762 (N_762,N_428,N_239);
nor U763 (N_763,N_144,N_185);
or U764 (N_764,N_93,N_183);
nand U765 (N_765,N_144,N_417);
xor U766 (N_766,N_351,N_496);
nand U767 (N_767,N_494,N_91);
nor U768 (N_768,N_493,N_51);
nand U769 (N_769,N_133,N_470);
xnor U770 (N_770,N_446,N_183);
nand U771 (N_771,N_45,N_215);
nand U772 (N_772,N_108,N_25);
xnor U773 (N_773,N_27,N_115);
nand U774 (N_774,N_72,N_462);
xor U775 (N_775,N_426,N_447);
xnor U776 (N_776,N_283,N_224);
and U777 (N_777,N_107,N_429);
xnor U778 (N_778,N_307,N_334);
nor U779 (N_779,N_465,N_336);
nand U780 (N_780,N_304,N_61);
and U781 (N_781,N_230,N_162);
xor U782 (N_782,N_276,N_318);
or U783 (N_783,N_430,N_444);
nand U784 (N_784,N_354,N_301);
xnor U785 (N_785,N_227,N_176);
nor U786 (N_786,N_309,N_266);
and U787 (N_787,N_103,N_2);
or U788 (N_788,N_137,N_276);
nand U789 (N_789,N_4,N_82);
or U790 (N_790,N_354,N_31);
or U791 (N_791,N_408,N_4);
nor U792 (N_792,N_68,N_450);
nor U793 (N_793,N_201,N_406);
and U794 (N_794,N_176,N_43);
nor U795 (N_795,N_363,N_466);
xor U796 (N_796,N_235,N_25);
or U797 (N_797,N_379,N_182);
nor U798 (N_798,N_269,N_188);
and U799 (N_799,N_277,N_257);
nor U800 (N_800,N_225,N_289);
nor U801 (N_801,N_286,N_146);
xor U802 (N_802,N_453,N_48);
or U803 (N_803,N_418,N_239);
nand U804 (N_804,N_104,N_198);
nor U805 (N_805,N_482,N_461);
or U806 (N_806,N_201,N_160);
nor U807 (N_807,N_365,N_247);
nor U808 (N_808,N_404,N_200);
nor U809 (N_809,N_312,N_144);
and U810 (N_810,N_7,N_101);
or U811 (N_811,N_359,N_12);
and U812 (N_812,N_330,N_408);
or U813 (N_813,N_427,N_72);
xnor U814 (N_814,N_49,N_397);
or U815 (N_815,N_36,N_302);
nand U816 (N_816,N_51,N_82);
nor U817 (N_817,N_138,N_410);
nor U818 (N_818,N_388,N_11);
nor U819 (N_819,N_67,N_150);
xor U820 (N_820,N_224,N_464);
nor U821 (N_821,N_376,N_454);
xor U822 (N_822,N_27,N_387);
or U823 (N_823,N_116,N_281);
nand U824 (N_824,N_136,N_408);
or U825 (N_825,N_180,N_33);
xnor U826 (N_826,N_179,N_1);
and U827 (N_827,N_261,N_67);
nor U828 (N_828,N_152,N_221);
or U829 (N_829,N_374,N_11);
or U830 (N_830,N_181,N_499);
nor U831 (N_831,N_244,N_136);
nor U832 (N_832,N_239,N_126);
nor U833 (N_833,N_382,N_150);
nand U834 (N_834,N_118,N_304);
nand U835 (N_835,N_183,N_42);
nor U836 (N_836,N_296,N_42);
nor U837 (N_837,N_56,N_276);
or U838 (N_838,N_421,N_65);
nor U839 (N_839,N_114,N_128);
nand U840 (N_840,N_146,N_444);
nand U841 (N_841,N_286,N_88);
or U842 (N_842,N_413,N_279);
and U843 (N_843,N_325,N_321);
and U844 (N_844,N_69,N_93);
nand U845 (N_845,N_270,N_196);
and U846 (N_846,N_121,N_92);
nand U847 (N_847,N_65,N_322);
xnor U848 (N_848,N_196,N_423);
nor U849 (N_849,N_360,N_104);
or U850 (N_850,N_95,N_246);
nand U851 (N_851,N_392,N_123);
nand U852 (N_852,N_390,N_449);
or U853 (N_853,N_446,N_311);
nand U854 (N_854,N_266,N_3);
nand U855 (N_855,N_208,N_226);
nor U856 (N_856,N_305,N_79);
nand U857 (N_857,N_47,N_57);
xnor U858 (N_858,N_439,N_4);
nor U859 (N_859,N_421,N_471);
nor U860 (N_860,N_337,N_338);
xnor U861 (N_861,N_289,N_161);
xor U862 (N_862,N_473,N_37);
nor U863 (N_863,N_2,N_214);
and U864 (N_864,N_310,N_366);
and U865 (N_865,N_372,N_380);
or U866 (N_866,N_434,N_148);
xor U867 (N_867,N_426,N_303);
nor U868 (N_868,N_389,N_418);
nor U869 (N_869,N_466,N_413);
nor U870 (N_870,N_161,N_1);
xnor U871 (N_871,N_433,N_303);
or U872 (N_872,N_236,N_0);
xor U873 (N_873,N_81,N_388);
or U874 (N_874,N_377,N_485);
nor U875 (N_875,N_220,N_379);
nand U876 (N_876,N_129,N_187);
and U877 (N_877,N_35,N_309);
or U878 (N_878,N_311,N_395);
and U879 (N_879,N_95,N_198);
and U880 (N_880,N_224,N_405);
nand U881 (N_881,N_167,N_302);
nand U882 (N_882,N_94,N_82);
nor U883 (N_883,N_137,N_78);
xor U884 (N_884,N_473,N_475);
nand U885 (N_885,N_297,N_279);
or U886 (N_886,N_226,N_252);
xnor U887 (N_887,N_75,N_183);
nand U888 (N_888,N_16,N_405);
xor U889 (N_889,N_14,N_55);
nand U890 (N_890,N_364,N_231);
or U891 (N_891,N_293,N_311);
xor U892 (N_892,N_231,N_149);
or U893 (N_893,N_495,N_123);
nor U894 (N_894,N_428,N_240);
nand U895 (N_895,N_477,N_397);
xnor U896 (N_896,N_63,N_495);
or U897 (N_897,N_458,N_190);
and U898 (N_898,N_294,N_375);
or U899 (N_899,N_198,N_386);
and U900 (N_900,N_268,N_202);
nand U901 (N_901,N_247,N_107);
nand U902 (N_902,N_272,N_82);
xnor U903 (N_903,N_346,N_499);
nand U904 (N_904,N_201,N_172);
nand U905 (N_905,N_84,N_140);
nand U906 (N_906,N_202,N_78);
xnor U907 (N_907,N_279,N_291);
or U908 (N_908,N_288,N_471);
and U909 (N_909,N_238,N_239);
and U910 (N_910,N_411,N_415);
nor U911 (N_911,N_34,N_180);
xnor U912 (N_912,N_185,N_36);
nand U913 (N_913,N_47,N_81);
nor U914 (N_914,N_459,N_152);
nor U915 (N_915,N_409,N_17);
xnor U916 (N_916,N_21,N_30);
nor U917 (N_917,N_243,N_93);
nor U918 (N_918,N_284,N_239);
and U919 (N_919,N_117,N_360);
and U920 (N_920,N_134,N_239);
or U921 (N_921,N_241,N_323);
nor U922 (N_922,N_466,N_327);
or U923 (N_923,N_193,N_419);
nand U924 (N_924,N_325,N_419);
nor U925 (N_925,N_103,N_321);
nand U926 (N_926,N_338,N_432);
nand U927 (N_927,N_252,N_195);
nand U928 (N_928,N_475,N_33);
nor U929 (N_929,N_94,N_120);
and U930 (N_930,N_177,N_268);
xor U931 (N_931,N_448,N_222);
nand U932 (N_932,N_407,N_364);
nor U933 (N_933,N_77,N_46);
xnor U934 (N_934,N_224,N_280);
and U935 (N_935,N_109,N_130);
nand U936 (N_936,N_85,N_492);
and U937 (N_937,N_135,N_462);
nand U938 (N_938,N_279,N_376);
nor U939 (N_939,N_164,N_365);
xnor U940 (N_940,N_334,N_398);
and U941 (N_941,N_354,N_156);
nor U942 (N_942,N_12,N_267);
nand U943 (N_943,N_249,N_344);
nor U944 (N_944,N_359,N_379);
and U945 (N_945,N_253,N_444);
and U946 (N_946,N_364,N_224);
nand U947 (N_947,N_79,N_427);
xor U948 (N_948,N_440,N_422);
nor U949 (N_949,N_66,N_305);
nand U950 (N_950,N_248,N_368);
and U951 (N_951,N_242,N_363);
or U952 (N_952,N_38,N_278);
nand U953 (N_953,N_321,N_246);
xor U954 (N_954,N_233,N_272);
xor U955 (N_955,N_81,N_216);
xnor U956 (N_956,N_230,N_54);
or U957 (N_957,N_133,N_50);
nor U958 (N_958,N_459,N_150);
nand U959 (N_959,N_177,N_193);
nor U960 (N_960,N_1,N_259);
xnor U961 (N_961,N_193,N_68);
and U962 (N_962,N_447,N_421);
xor U963 (N_963,N_150,N_142);
and U964 (N_964,N_411,N_413);
xnor U965 (N_965,N_386,N_480);
and U966 (N_966,N_444,N_402);
xnor U967 (N_967,N_85,N_78);
and U968 (N_968,N_155,N_74);
or U969 (N_969,N_432,N_286);
or U970 (N_970,N_20,N_399);
xor U971 (N_971,N_137,N_70);
and U972 (N_972,N_341,N_219);
nor U973 (N_973,N_492,N_236);
nor U974 (N_974,N_174,N_267);
nor U975 (N_975,N_316,N_448);
xnor U976 (N_976,N_494,N_281);
nand U977 (N_977,N_276,N_197);
nor U978 (N_978,N_411,N_17);
or U979 (N_979,N_79,N_340);
nand U980 (N_980,N_472,N_145);
xnor U981 (N_981,N_102,N_244);
or U982 (N_982,N_8,N_207);
nand U983 (N_983,N_252,N_453);
or U984 (N_984,N_61,N_134);
nand U985 (N_985,N_194,N_266);
or U986 (N_986,N_323,N_88);
nor U987 (N_987,N_207,N_61);
and U988 (N_988,N_416,N_325);
xnor U989 (N_989,N_403,N_275);
and U990 (N_990,N_206,N_489);
and U991 (N_991,N_159,N_344);
nand U992 (N_992,N_440,N_53);
or U993 (N_993,N_343,N_311);
and U994 (N_994,N_387,N_117);
xnor U995 (N_995,N_482,N_419);
and U996 (N_996,N_67,N_139);
nor U997 (N_997,N_175,N_291);
nor U998 (N_998,N_34,N_488);
nand U999 (N_999,N_58,N_344);
xor U1000 (N_1000,N_644,N_786);
nor U1001 (N_1001,N_757,N_646);
and U1002 (N_1002,N_558,N_660);
nand U1003 (N_1003,N_874,N_563);
and U1004 (N_1004,N_622,N_752);
xor U1005 (N_1005,N_546,N_908);
nor U1006 (N_1006,N_948,N_989);
nand U1007 (N_1007,N_535,N_674);
nand U1008 (N_1008,N_781,N_549);
nand U1009 (N_1009,N_946,N_821);
nand U1010 (N_1010,N_987,N_921);
xor U1011 (N_1011,N_667,N_709);
and U1012 (N_1012,N_841,N_689);
xnor U1013 (N_1013,N_716,N_918);
xor U1014 (N_1014,N_993,N_554);
nor U1015 (N_1015,N_606,N_832);
or U1016 (N_1016,N_574,N_528);
and U1017 (N_1017,N_695,N_883);
nor U1018 (N_1018,N_762,N_794);
or U1019 (N_1019,N_710,N_933);
nor U1020 (N_1020,N_871,N_766);
nor U1021 (N_1021,N_715,N_631);
or U1022 (N_1022,N_595,N_515);
and U1023 (N_1023,N_979,N_659);
nand U1024 (N_1024,N_550,N_553);
xor U1025 (N_1025,N_712,N_584);
and U1026 (N_1026,N_639,N_517);
and U1027 (N_1027,N_976,N_647);
nor U1028 (N_1028,N_912,N_530);
nor U1029 (N_1029,N_573,N_893);
nor U1030 (N_1030,N_888,N_729);
and U1031 (N_1031,N_610,N_842);
or U1032 (N_1032,N_889,N_787);
xor U1033 (N_1033,N_759,N_527);
or U1034 (N_1034,N_688,N_742);
or U1035 (N_1035,N_941,N_512);
xnor U1036 (N_1036,N_945,N_697);
and U1037 (N_1037,N_625,N_561);
nand U1038 (N_1038,N_902,N_592);
and U1039 (N_1039,N_605,N_840);
or U1040 (N_1040,N_788,N_895);
xor U1041 (N_1041,N_833,N_925);
xnor U1042 (N_1042,N_800,N_763);
and U1043 (N_1043,N_702,N_614);
nor U1044 (N_1044,N_663,N_732);
nor U1045 (N_1045,N_621,N_814);
or U1046 (N_1046,N_679,N_881);
xor U1047 (N_1047,N_858,N_939);
xor U1048 (N_1048,N_940,N_543);
nand U1049 (N_1049,N_966,N_990);
nor U1050 (N_1050,N_739,N_831);
nand U1051 (N_1051,N_538,N_587);
and U1052 (N_1052,N_637,N_579);
xnor U1053 (N_1053,N_765,N_506);
xnor U1054 (N_1054,N_919,N_819);
xnor U1055 (N_1055,N_636,N_648);
nand U1056 (N_1056,N_728,N_552);
nor U1057 (N_1057,N_932,N_632);
and U1058 (N_1058,N_582,N_534);
nand U1059 (N_1059,N_964,N_661);
or U1060 (N_1060,N_928,N_731);
nor U1061 (N_1061,N_854,N_656);
xor U1062 (N_1062,N_827,N_686);
and U1063 (N_1063,N_980,N_746);
and U1064 (N_1064,N_655,N_607);
or U1065 (N_1065,N_892,N_718);
and U1066 (N_1066,N_780,N_801);
xnor U1067 (N_1067,N_782,N_594);
nor U1068 (N_1068,N_880,N_789);
and U1069 (N_1069,N_523,N_521);
nand U1070 (N_1070,N_922,N_968);
nor U1071 (N_1071,N_913,N_577);
nand U1072 (N_1072,N_982,N_873);
nand U1073 (N_1073,N_749,N_770);
xnor U1074 (N_1074,N_704,N_955);
nand U1075 (N_1075,N_693,N_872);
or U1076 (N_1076,N_572,N_745);
xor U1077 (N_1077,N_511,N_862);
and U1078 (N_1078,N_935,N_950);
or U1079 (N_1079,N_896,N_949);
nand U1080 (N_1080,N_779,N_985);
and U1081 (N_1081,N_815,N_600);
and U1082 (N_1082,N_568,N_743);
nor U1083 (N_1083,N_834,N_609);
nand U1084 (N_1084,N_901,N_744);
or U1085 (N_1085,N_641,N_843);
nand U1086 (N_1086,N_685,N_876);
xor U1087 (N_1087,N_967,N_856);
or U1088 (N_1088,N_531,N_929);
xnor U1089 (N_1089,N_585,N_599);
nor U1090 (N_1090,N_683,N_981);
nor U1091 (N_1091,N_545,N_720);
nor U1092 (N_1092,N_920,N_691);
and U1093 (N_1093,N_516,N_645);
xor U1094 (N_1094,N_707,N_542);
nor U1095 (N_1095,N_662,N_962);
and U1096 (N_1096,N_867,N_975);
nand U1097 (N_1097,N_995,N_520);
and U1098 (N_1098,N_774,N_775);
or U1099 (N_1099,N_690,N_589);
nand U1100 (N_1100,N_899,N_954);
nand U1101 (N_1101,N_978,N_750);
nor U1102 (N_1102,N_785,N_591);
and U1103 (N_1103,N_986,N_996);
or U1104 (N_1104,N_510,N_806);
nor U1105 (N_1105,N_803,N_758);
or U1106 (N_1106,N_708,N_548);
nor U1107 (N_1107,N_608,N_866);
nor U1108 (N_1108,N_851,N_910);
nand U1109 (N_1109,N_570,N_713);
or U1110 (N_1110,N_664,N_926);
nor U1111 (N_1111,N_882,N_529);
and U1112 (N_1112,N_556,N_813);
nor U1113 (N_1113,N_942,N_859);
nand U1114 (N_1114,N_738,N_673);
and U1115 (N_1115,N_924,N_958);
nor U1116 (N_1116,N_615,N_723);
nor U1117 (N_1117,N_703,N_783);
xor U1118 (N_1118,N_701,N_879);
nand U1119 (N_1119,N_736,N_658);
nand U1120 (N_1120,N_604,N_635);
or U1121 (N_1121,N_751,N_578);
nand U1122 (N_1122,N_848,N_860);
or U1123 (N_1123,N_952,N_937);
and U1124 (N_1124,N_825,N_914);
nand U1125 (N_1125,N_822,N_828);
and U1126 (N_1126,N_657,N_740);
nand U1127 (N_1127,N_972,N_977);
nand U1128 (N_1128,N_559,N_923);
or U1129 (N_1129,N_726,N_551);
and U1130 (N_1130,N_875,N_557);
and U1131 (N_1131,N_569,N_590);
nor U1132 (N_1132,N_830,N_628);
nand U1133 (N_1133,N_500,N_887);
xnor U1134 (N_1134,N_798,N_602);
nor U1135 (N_1135,N_878,N_974);
nand U1136 (N_1136,N_760,N_863);
nor U1137 (N_1137,N_620,N_983);
nand U1138 (N_1138,N_727,N_812);
xnor U1139 (N_1139,N_586,N_884);
xor U1140 (N_1140,N_906,N_818);
and U1141 (N_1141,N_643,N_838);
nor U1142 (N_1142,N_717,N_885);
xnor U1143 (N_1143,N_654,N_761);
nor U1144 (N_1144,N_817,N_963);
nor U1145 (N_1145,N_810,N_583);
or U1146 (N_1146,N_769,N_507);
and U1147 (N_1147,N_501,N_777);
and U1148 (N_1148,N_518,N_820);
nand U1149 (N_1149,N_877,N_824);
nand U1150 (N_1150,N_675,N_796);
nand U1151 (N_1151,N_665,N_504);
and U1152 (N_1152,N_960,N_634);
nand U1153 (N_1153,N_730,N_539);
nor U1154 (N_1154,N_541,N_651);
and U1155 (N_1155,N_677,N_555);
nor U1156 (N_1156,N_865,N_580);
xor U1157 (N_1157,N_532,N_997);
nand U1158 (N_1158,N_505,N_536);
nor U1159 (N_1159,N_640,N_544);
or U1160 (N_1160,N_627,N_698);
nor U1161 (N_1161,N_957,N_984);
or U1162 (N_1162,N_721,N_560);
or U1163 (N_1163,N_694,N_951);
nand U1164 (N_1164,N_617,N_747);
xor U1165 (N_1165,N_998,N_891);
xor U1166 (N_1166,N_959,N_671);
nand U1167 (N_1167,N_524,N_619);
xor U1168 (N_1168,N_791,N_588);
nor U1169 (N_1169,N_965,N_936);
or U1170 (N_1170,N_633,N_714);
or U1171 (N_1171,N_927,N_649);
nand U1172 (N_1172,N_755,N_894);
or U1173 (N_1173,N_650,N_537);
nand U1174 (N_1174,N_735,N_795);
nor U1175 (N_1175,N_823,N_680);
nor U1176 (N_1176,N_696,N_564);
and U1177 (N_1177,N_508,N_826);
xor U1178 (N_1178,N_670,N_699);
nand U1179 (N_1179,N_849,N_700);
nand U1180 (N_1180,N_567,N_853);
nand U1181 (N_1181,N_915,N_784);
or U1182 (N_1182,N_869,N_597);
or U1183 (N_1183,N_756,N_630);
nand U1184 (N_1184,N_846,N_971);
nor U1185 (N_1185,N_845,N_711);
nor U1186 (N_1186,N_611,N_930);
or U1187 (N_1187,N_581,N_857);
nand U1188 (N_1188,N_861,N_672);
xnor U1189 (N_1189,N_575,N_768);
and U1190 (N_1190,N_669,N_754);
or U1191 (N_1191,N_705,N_999);
xor U1192 (N_1192,N_626,N_519);
or U1193 (N_1193,N_776,N_953);
nor U1194 (N_1194,N_904,N_870);
nor U1195 (N_1195,N_733,N_684);
and U1196 (N_1196,N_767,N_753);
nand U1197 (N_1197,N_601,N_829);
and U1198 (N_1198,N_562,N_947);
and U1199 (N_1199,N_804,N_623);
nand U1200 (N_1200,N_808,N_844);
xor U1201 (N_1201,N_847,N_502);
xor U1202 (N_1202,N_917,N_973);
nor U1203 (N_1203,N_682,N_816);
nand U1204 (N_1204,N_836,N_513);
or U1205 (N_1205,N_916,N_944);
or U1206 (N_1206,N_612,N_722);
and U1207 (N_1207,N_835,N_681);
nor U1208 (N_1208,N_503,N_687);
nand U1209 (N_1209,N_719,N_864);
xnor U1210 (N_1210,N_629,N_961);
xnor U1211 (N_1211,N_725,N_850);
nand U1212 (N_1212,N_900,N_692);
nand U1213 (N_1213,N_593,N_613);
nor U1214 (N_1214,N_596,N_571);
nor U1215 (N_1215,N_565,N_943);
nor U1216 (N_1216,N_852,N_907);
nor U1217 (N_1217,N_676,N_956);
nand U1218 (N_1218,N_652,N_526);
and U1219 (N_1219,N_547,N_793);
xnor U1220 (N_1220,N_764,N_603);
and U1221 (N_1221,N_666,N_799);
and U1222 (N_1222,N_741,N_991);
and U1223 (N_1223,N_802,N_624);
nand U1224 (N_1224,N_938,N_790);
nor U1225 (N_1225,N_992,N_778);
nor U1226 (N_1226,N_734,N_737);
nor U1227 (N_1227,N_706,N_540);
nor U1228 (N_1228,N_638,N_886);
nor U1229 (N_1229,N_797,N_970);
and U1230 (N_1230,N_839,N_855);
and U1231 (N_1231,N_653,N_837);
nor U1232 (N_1232,N_911,N_522);
or U1233 (N_1233,N_724,N_931);
xnor U1234 (N_1234,N_811,N_566);
or U1235 (N_1235,N_748,N_805);
or U1236 (N_1236,N_807,N_618);
nor U1237 (N_1237,N_772,N_533);
xor U1238 (N_1238,N_668,N_868);
nand U1239 (N_1239,N_909,N_598);
nand U1240 (N_1240,N_514,N_773);
nor U1241 (N_1241,N_771,N_792);
nor U1242 (N_1242,N_897,N_809);
nand U1243 (N_1243,N_934,N_678);
nand U1244 (N_1244,N_525,N_642);
xnor U1245 (N_1245,N_898,N_903);
nand U1246 (N_1246,N_905,N_576);
xnor U1247 (N_1247,N_890,N_988);
and U1248 (N_1248,N_969,N_509);
or U1249 (N_1249,N_616,N_994);
nor U1250 (N_1250,N_914,N_765);
or U1251 (N_1251,N_776,N_682);
or U1252 (N_1252,N_510,N_753);
or U1253 (N_1253,N_757,N_725);
nand U1254 (N_1254,N_639,N_622);
nor U1255 (N_1255,N_905,N_558);
or U1256 (N_1256,N_814,N_697);
nor U1257 (N_1257,N_818,N_554);
xor U1258 (N_1258,N_730,N_772);
or U1259 (N_1259,N_643,N_922);
nand U1260 (N_1260,N_755,N_884);
nor U1261 (N_1261,N_734,N_524);
xor U1262 (N_1262,N_556,N_603);
nand U1263 (N_1263,N_764,N_843);
xnor U1264 (N_1264,N_582,N_846);
nor U1265 (N_1265,N_935,N_760);
nand U1266 (N_1266,N_968,N_500);
nor U1267 (N_1267,N_600,N_552);
and U1268 (N_1268,N_947,N_523);
nor U1269 (N_1269,N_958,N_609);
or U1270 (N_1270,N_922,N_702);
xnor U1271 (N_1271,N_697,N_745);
nand U1272 (N_1272,N_704,N_647);
nor U1273 (N_1273,N_629,N_805);
nor U1274 (N_1274,N_772,N_517);
xnor U1275 (N_1275,N_953,N_654);
nor U1276 (N_1276,N_877,N_614);
xor U1277 (N_1277,N_890,N_750);
nand U1278 (N_1278,N_711,N_540);
xnor U1279 (N_1279,N_697,N_683);
nand U1280 (N_1280,N_627,N_757);
xnor U1281 (N_1281,N_598,N_575);
and U1282 (N_1282,N_782,N_924);
or U1283 (N_1283,N_663,N_751);
xnor U1284 (N_1284,N_581,N_675);
nand U1285 (N_1285,N_918,N_507);
xnor U1286 (N_1286,N_841,N_552);
or U1287 (N_1287,N_774,N_591);
xor U1288 (N_1288,N_598,N_844);
nor U1289 (N_1289,N_621,N_944);
and U1290 (N_1290,N_515,N_510);
or U1291 (N_1291,N_820,N_696);
nor U1292 (N_1292,N_695,N_676);
or U1293 (N_1293,N_745,N_652);
or U1294 (N_1294,N_760,N_577);
nor U1295 (N_1295,N_943,N_553);
and U1296 (N_1296,N_688,N_960);
or U1297 (N_1297,N_749,N_786);
nand U1298 (N_1298,N_624,N_668);
and U1299 (N_1299,N_800,N_882);
nand U1300 (N_1300,N_712,N_975);
or U1301 (N_1301,N_516,N_958);
nor U1302 (N_1302,N_690,N_536);
xor U1303 (N_1303,N_560,N_742);
nand U1304 (N_1304,N_749,N_603);
xnor U1305 (N_1305,N_983,N_624);
and U1306 (N_1306,N_745,N_536);
xor U1307 (N_1307,N_932,N_520);
and U1308 (N_1308,N_626,N_980);
nor U1309 (N_1309,N_763,N_560);
and U1310 (N_1310,N_556,N_527);
nand U1311 (N_1311,N_957,N_718);
nor U1312 (N_1312,N_836,N_896);
or U1313 (N_1313,N_626,N_801);
nor U1314 (N_1314,N_560,N_720);
nor U1315 (N_1315,N_529,N_553);
or U1316 (N_1316,N_553,N_957);
and U1317 (N_1317,N_634,N_970);
or U1318 (N_1318,N_860,N_671);
nor U1319 (N_1319,N_849,N_933);
and U1320 (N_1320,N_787,N_660);
and U1321 (N_1321,N_800,N_583);
and U1322 (N_1322,N_547,N_597);
and U1323 (N_1323,N_895,N_801);
nand U1324 (N_1324,N_747,N_573);
and U1325 (N_1325,N_783,N_950);
nand U1326 (N_1326,N_570,N_804);
nand U1327 (N_1327,N_780,N_788);
xor U1328 (N_1328,N_962,N_658);
nor U1329 (N_1329,N_948,N_670);
nand U1330 (N_1330,N_632,N_902);
xnor U1331 (N_1331,N_983,N_651);
xor U1332 (N_1332,N_900,N_802);
or U1333 (N_1333,N_727,N_751);
and U1334 (N_1334,N_724,N_752);
xnor U1335 (N_1335,N_580,N_625);
nand U1336 (N_1336,N_557,N_568);
xor U1337 (N_1337,N_798,N_539);
or U1338 (N_1338,N_546,N_599);
nand U1339 (N_1339,N_709,N_830);
nor U1340 (N_1340,N_965,N_916);
and U1341 (N_1341,N_766,N_773);
nor U1342 (N_1342,N_648,N_707);
nor U1343 (N_1343,N_802,N_625);
nand U1344 (N_1344,N_560,N_615);
nand U1345 (N_1345,N_675,N_503);
xor U1346 (N_1346,N_521,N_997);
nor U1347 (N_1347,N_601,N_756);
or U1348 (N_1348,N_583,N_874);
xor U1349 (N_1349,N_757,N_590);
nor U1350 (N_1350,N_793,N_543);
xnor U1351 (N_1351,N_769,N_724);
xor U1352 (N_1352,N_704,N_867);
nor U1353 (N_1353,N_762,N_714);
nand U1354 (N_1354,N_826,N_582);
nand U1355 (N_1355,N_746,N_644);
and U1356 (N_1356,N_633,N_768);
nor U1357 (N_1357,N_606,N_721);
nor U1358 (N_1358,N_710,N_871);
nor U1359 (N_1359,N_628,N_661);
nor U1360 (N_1360,N_735,N_744);
nand U1361 (N_1361,N_527,N_830);
xnor U1362 (N_1362,N_651,N_984);
and U1363 (N_1363,N_621,N_590);
or U1364 (N_1364,N_627,N_640);
xnor U1365 (N_1365,N_877,N_930);
and U1366 (N_1366,N_587,N_561);
nor U1367 (N_1367,N_709,N_811);
nand U1368 (N_1368,N_656,N_640);
xor U1369 (N_1369,N_648,N_943);
xnor U1370 (N_1370,N_892,N_596);
xnor U1371 (N_1371,N_753,N_722);
or U1372 (N_1372,N_941,N_848);
nand U1373 (N_1373,N_540,N_951);
or U1374 (N_1374,N_982,N_875);
or U1375 (N_1375,N_569,N_824);
and U1376 (N_1376,N_848,N_791);
xnor U1377 (N_1377,N_845,N_950);
nand U1378 (N_1378,N_733,N_712);
nand U1379 (N_1379,N_618,N_799);
and U1380 (N_1380,N_738,N_953);
nand U1381 (N_1381,N_551,N_772);
or U1382 (N_1382,N_914,N_550);
and U1383 (N_1383,N_527,N_780);
or U1384 (N_1384,N_749,N_768);
or U1385 (N_1385,N_771,N_834);
and U1386 (N_1386,N_574,N_836);
and U1387 (N_1387,N_594,N_692);
or U1388 (N_1388,N_870,N_582);
and U1389 (N_1389,N_937,N_715);
or U1390 (N_1390,N_867,N_512);
xnor U1391 (N_1391,N_640,N_558);
or U1392 (N_1392,N_936,N_747);
nor U1393 (N_1393,N_822,N_839);
xor U1394 (N_1394,N_550,N_830);
and U1395 (N_1395,N_910,N_549);
or U1396 (N_1396,N_781,N_701);
and U1397 (N_1397,N_867,N_841);
nand U1398 (N_1398,N_832,N_924);
xnor U1399 (N_1399,N_665,N_967);
xnor U1400 (N_1400,N_661,N_887);
nor U1401 (N_1401,N_771,N_703);
xnor U1402 (N_1402,N_521,N_839);
nor U1403 (N_1403,N_978,N_764);
and U1404 (N_1404,N_796,N_633);
xor U1405 (N_1405,N_914,N_788);
nor U1406 (N_1406,N_799,N_915);
nand U1407 (N_1407,N_869,N_662);
nor U1408 (N_1408,N_918,N_513);
nand U1409 (N_1409,N_636,N_595);
nand U1410 (N_1410,N_985,N_738);
xnor U1411 (N_1411,N_733,N_982);
or U1412 (N_1412,N_628,N_522);
xor U1413 (N_1413,N_816,N_942);
nor U1414 (N_1414,N_563,N_535);
or U1415 (N_1415,N_814,N_785);
nor U1416 (N_1416,N_800,N_983);
or U1417 (N_1417,N_996,N_656);
and U1418 (N_1418,N_647,N_561);
nor U1419 (N_1419,N_567,N_965);
and U1420 (N_1420,N_732,N_965);
and U1421 (N_1421,N_952,N_713);
and U1422 (N_1422,N_801,N_576);
or U1423 (N_1423,N_711,N_767);
xor U1424 (N_1424,N_963,N_874);
and U1425 (N_1425,N_724,N_708);
or U1426 (N_1426,N_968,N_747);
xnor U1427 (N_1427,N_884,N_912);
nor U1428 (N_1428,N_521,N_594);
or U1429 (N_1429,N_824,N_655);
nor U1430 (N_1430,N_505,N_767);
nand U1431 (N_1431,N_564,N_654);
nand U1432 (N_1432,N_500,N_597);
nor U1433 (N_1433,N_694,N_958);
xnor U1434 (N_1434,N_929,N_848);
and U1435 (N_1435,N_552,N_589);
nand U1436 (N_1436,N_812,N_832);
or U1437 (N_1437,N_511,N_727);
nand U1438 (N_1438,N_684,N_968);
and U1439 (N_1439,N_953,N_917);
nor U1440 (N_1440,N_984,N_975);
nand U1441 (N_1441,N_886,N_874);
nand U1442 (N_1442,N_865,N_967);
or U1443 (N_1443,N_795,N_733);
nand U1444 (N_1444,N_861,N_602);
nand U1445 (N_1445,N_908,N_929);
xor U1446 (N_1446,N_633,N_596);
nor U1447 (N_1447,N_980,N_973);
nand U1448 (N_1448,N_904,N_740);
xnor U1449 (N_1449,N_983,N_952);
or U1450 (N_1450,N_758,N_764);
or U1451 (N_1451,N_941,N_811);
xor U1452 (N_1452,N_835,N_777);
xnor U1453 (N_1453,N_704,N_633);
or U1454 (N_1454,N_655,N_739);
nor U1455 (N_1455,N_606,N_682);
nor U1456 (N_1456,N_994,N_829);
nor U1457 (N_1457,N_684,N_946);
and U1458 (N_1458,N_955,N_823);
xnor U1459 (N_1459,N_552,N_954);
xnor U1460 (N_1460,N_933,N_851);
nand U1461 (N_1461,N_524,N_692);
nor U1462 (N_1462,N_705,N_845);
xnor U1463 (N_1463,N_733,N_620);
xnor U1464 (N_1464,N_630,N_635);
or U1465 (N_1465,N_805,N_817);
and U1466 (N_1466,N_691,N_630);
nor U1467 (N_1467,N_560,N_893);
nor U1468 (N_1468,N_540,N_673);
nand U1469 (N_1469,N_662,N_535);
and U1470 (N_1470,N_568,N_966);
nand U1471 (N_1471,N_927,N_994);
nand U1472 (N_1472,N_654,N_730);
and U1473 (N_1473,N_508,N_848);
nor U1474 (N_1474,N_524,N_873);
nor U1475 (N_1475,N_771,N_621);
nand U1476 (N_1476,N_933,N_690);
nor U1477 (N_1477,N_917,N_730);
nor U1478 (N_1478,N_552,N_903);
nor U1479 (N_1479,N_922,N_865);
nand U1480 (N_1480,N_936,N_924);
nand U1481 (N_1481,N_527,N_710);
or U1482 (N_1482,N_817,N_540);
nand U1483 (N_1483,N_970,N_920);
nor U1484 (N_1484,N_936,N_605);
xnor U1485 (N_1485,N_836,N_916);
or U1486 (N_1486,N_699,N_606);
xor U1487 (N_1487,N_717,N_827);
nor U1488 (N_1488,N_694,N_574);
and U1489 (N_1489,N_679,N_597);
nand U1490 (N_1490,N_819,N_902);
nand U1491 (N_1491,N_672,N_884);
nand U1492 (N_1492,N_742,N_630);
and U1493 (N_1493,N_632,N_924);
and U1494 (N_1494,N_657,N_508);
or U1495 (N_1495,N_775,N_510);
nand U1496 (N_1496,N_573,N_512);
or U1497 (N_1497,N_701,N_586);
nand U1498 (N_1498,N_800,N_940);
nand U1499 (N_1499,N_863,N_773);
and U1500 (N_1500,N_1462,N_1349);
nor U1501 (N_1501,N_1356,N_1407);
nor U1502 (N_1502,N_1438,N_1090);
and U1503 (N_1503,N_1359,N_1254);
nor U1504 (N_1504,N_1123,N_1456);
nand U1505 (N_1505,N_1103,N_1242);
nand U1506 (N_1506,N_1178,N_1129);
xnor U1507 (N_1507,N_1382,N_1189);
or U1508 (N_1508,N_1116,N_1088);
or U1509 (N_1509,N_1460,N_1468);
nor U1510 (N_1510,N_1112,N_1117);
xor U1511 (N_1511,N_1311,N_1362);
nand U1512 (N_1512,N_1134,N_1445);
nand U1513 (N_1513,N_1338,N_1160);
xnor U1514 (N_1514,N_1008,N_1387);
xnor U1515 (N_1515,N_1007,N_1040);
or U1516 (N_1516,N_1035,N_1137);
xor U1517 (N_1517,N_1094,N_1432);
nand U1518 (N_1518,N_1493,N_1290);
nand U1519 (N_1519,N_1175,N_1425);
nor U1520 (N_1520,N_1062,N_1264);
xnor U1521 (N_1521,N_1163,N_1195);
or U1522 (N_1522,N_1437,N_1193);
nand U1523 (N_1523,N_1279,N_1442);
and U1524 (N_1524,N_1474,N_1249);
nor U1525 (N_1525,N_1216,N_1325);
xnor U1526 (N_1526,N_1471,N_1488);
nand U1527 (N_1527,N_1145,N_1065);
and U1528 (N_1528,N_1370,N_1310);
nor U1529 (N_1529,N_1330,N_1089);
and U1530 (N_1530,N_1095,N_1033);
and U1531 (N_1531,N_1139,N_1306);
nand U1532 (N_1532,N_1102,N_1473);
nand U1533 (N_1533,N_1034,N_1205);
nand U1534 (N_1534,N_1157,N_1141);
nor U1535 (N_1535,N_1384,N_1245);
or U1536 (N_1536,N_1379,N_1267);
xor U1537 (N_1537,N_1326,N_1128);
xor U1538 (N_1538,N_1053,N_1498);
and U1539 (N_1539,N_1410,N_1466);
or U1540 (N_1540,N_1050,N_1101);
nand U1541 (N_1541,N_1074,N_1204);
nand U1542 (N_1542,N_1272,N_1332);
xnor U1543 (N_1543,N_1239,N_1111);
xor U1544 (N_1544,N_1457,N_1293);
or U1545 (N_1545,N_1212,N_1097);
nand U1546 (N_1546,N_1105,N_1336);
nor U1547 (N_1547,N_1274,N_1415);
and U1548 (N_1548,N_1217,N_1182);
xnor U1549 (N_1549,N_1023,N_1361);
or U1550 (N_1550,N_1435,N_1452);
nand U1551 (N_1551,N_1122,N_1342);
and U1552 (N_1552,N_1098,N_1060);
xnor U1553 (N_1553,N_1283,N_1397);
xnor U1554 (N_1554,N_1100,N_1164);
nand U1555 (N_1555,N_1312,N_1269);
nor U1556 (N_1556,N_1411,N_1433);
or U1557 (N_1557,N_1369,N_1064);
nor U1558 (N_1558,N_1403,N_1333);
nand U1559 (N_1559,N_1177,N_1377);
and U1560 (N_1560,N_1467,N_1078);
nor U1561 (N_1561,N_1258,N_1373);
or U1562 (N_1562,N_1434,N_1131);
and U1563 (N_1563,N_1358,N_1307);
nand U1564 (N_1564,N_1109,N_1191);
nand U1565 (N_1565,N_1146,N_1346);
or U1566 (N_1566,N_1124,N_1126);
xnor U1567 (N_1567,N_1091,N_1421);
nand U1568 (N_1568,N_1199,N_1067);
and U1569 (N_1569,N_1138,N_1280);
nand U1570 (N_1570,N_1380,N_1207);
xnor U1571 (N_1571,N_1263,N_1057);
nor U1572 (N_1572,N_1276,N_1453);
nand U1573 (N_1573,N_1213,N_1464);
xnor U1574 (N_1574,N_1142,N_1357);
xnor U1575 (N_1575,N_1083,N_1448);
xor U1576 (N_1576,N_1299,N_1130);
nand U1577 (N_1577,N_1255,N_1496);
or U1578 (N_1578,N_1196,N_1499);
nor U1579 (N_1579,N_1005,N_1028);
nor U1580 (N_1580,N_1451,N_1444);
or U1581 (N_1581,N_1268,N_1019);
and U1582 (N_1582,N_1260,N_1472);
xor U1583 (N_1583,N_1270,N_1406);
and U1584 (N_1584,N_1198,N_1208);
or U1585 (N_1585,N_1278,N_1221);
or U1586 (N_1586,N_1398,N_1085);
xnor U1587 (N_1587,N_1291,N_1032);
nor U1588 (N_1588,N_1353,N_1354);
or U1589 (N_1589,N_1262,N_1069);
or U1590 (N_1590,N_1009,N_1055);
or U1591 (N_1591,N_1165,N_1381);
or U1592 (N_1592,N_1147,N_1121);
or U1593 (N_1593,N_1430,N_1324);
xnor U1594 (N_1594,N_1409,N_1450);
or U1595 (N_1595,N_1282,N_1001);
nor U1596 (N_1596,N_1487,N_1423);
and U1597 (N_1597,N_1174,N_1389);
nand U1598 (N_1598,N_1081,N_1153);
xor U1599 (N_1599,N_1003,N_1427);
xor U1600 (N_1600,N_1092,N_1171);
and U1601 (N_1601,N_1294,N_1486);
nand U1602 (N_1602,N_1393,N_1224);
and U1603 (N_1603,N_1017,N_1203);
nand U1604 (N_1604,N_1211,N_1015);
nand U1605 (N_1605,N_1314,N_1148);
nor U1606 (N_1606,N_1368,N_1316);
and U1607 (N_1607,N_1162,N_1351);
xor U1608 (N_1608,N_1226,N_1093);
nor U1609 (N_1609,N_1428,N_1475);
or U1610 (N_1610,N_1237,N_1495);
xor U1611 (N_1611,N_1289,N_1233);
xnor U1612 (N_1612,N_1419,N_1219);
nand U1613 (N_1613,N_1202,N_1363);
or U1614 (N_1614,N_1340,N_1039);
or U1615 (N_1615,N_1395,N_1072);
or U1616 (N_1616,N_1455,N_1386);
xnor U1617 (N_1617,N_1234,N_1176);
xor U1618 (N_1618,N_1253,N_1096);
and U1619 (N_1619,N_1244,N_1151);
or U1620 (N_1620,N_1303,N_1011);
or U1621 (N_1621,N_1315,N_1076);
nor U1622 (N_1622,N_1296,N_1113);
xnor U1623 (N_1623,N_1284,N_1155);
nor U1624 (N_1624,N_1227,N_1075);
or U1625 (N_1625,N_1149,N_1477);
or U1626 (N_1626,N_1000,N_1429);
xnor U1627 (N_1627,N_1396,N_1230);
and U1628 (N_1628,N_1218,N_1048);
or U1629 (N_1629,N_1073,N_1158);
nand U1630 (N_1630,N_1288,N_1002);
or U1631 (N_1631,N_1250,N_1412);
nand U1632 (N_1632,N_1115,N_1490);
or U1633 (N_1633,N_1214,N_1376);
nor U1634 (N_1634,N_1480,N_1236);
or U1635 (N_1635,N_1166,N_1181);
and U1636 (N_1636,N_1248,N_1232);
and U1637 (N_1637,N_1300,N_1084);
nand U1638 (N_1638,N_1059,N_1080);
or U1639 (N_1639,N_1309,N_1461);
nand U1640 (N_1640,N_1443,N_1063);
nor U1641 (N_1641,N_1018,N_1179);
nor U1642 (N_1642,N_1420,N_1172);
and U1643 (N_1643,N_1012,N_1401);
xnor U1644 (N_1644,N_1273,N_1335);
xor U1645 (N_1645,N_1385,N_1352);
or U1646 (N_1646,N_1099,N_1029);
nand U1647 (N_1647,N_1402,N_1365);
nor U1648 (N_1648,N_1271,N_1476);
and U1649 (N_1649,N_1238,N_1114);
or U1650 (N_1650,N_1156,N_1140);
xor U1651 (N_1651,N_1483,N_1405);
and U1652 (N_1652,N_1322,N_1038);
nor U1653 (N_1653,N_1305,N_1136);
xor U1654 (N_1654,N_1259,N_1025);
nand U1655 (N_1655,N_1378,N_1231);
nor U1656 (N_1656,N_1341,N_1133);
or U1657 (N_1657,N_1043,N_1167);
and U1658 (N_1658,N_1399,N_1068);
or U1659 (N_1659,N_1256,N_1187);
nor U1660 (N_1660,N_1497,N_1297);
xor U1661 (N_1661,N_1321,N_1209);
nand U1662 (N_1662,N_1388,N_1006);
or U1663 (N_1663,N_1004,N_1194);
or U1664 (N_1664,N_1491,N_1329);
and U1665 (N_1665,N_1235,N_1281);
or U1666 (N_1666,N_1334,N_1478);
xor U1667 (N_1667,N_1266,N_1215);
or U1668 (N_1668,N_1021,N_1049);
xnor U1669 (N_1669,N_1404,N_1037);
nor U1670 (N_1670,N_1454,N_1184);
nand U1671 (N_1671,N_1107,N_1173);
nand U1672 (N_1672,N_1127,N_1257);
xor U1673 (N_1673,N_1036,N_1304);
xnor U1674 (N_1674,N_1119,N_1343);
nand U1675 (N_1675,N_1228,N_1374);
and U1676 (N_1676,N_1247,N_1143);
and U1677 (N_1677,N_1417,N_1056);
or U1678 (N_1678,N_1344,N_1013);
nand U1679 (N_1679,N_1240,N_1459);
or U1680 (N_1680,N_1366,N_1408);
xor U1681 (N_1681,N_1328,N_1125);
nand U1682 (N_1682,N_1392,N_1106);
nand U1683 (N_1683,N_1070,N_1355);
or U1684 (N_1684,N_1022,N_1225);
and U1685 (N_1685,N_1104,N_1180);
nor U1686 (N_1686,N_1479,N_1440);
nor U1687 (N_1687,N_1161,N_1120);
nor U1688 (N_1688,N_1030,N_1313);
or U1689 (N_1689,N_1243,N_1422);
nor U1690 (N_1690,N_1337,N_1168);
or U1691 (N_1691,N_1044,N_1446);
nor U1692 (N_1692,N_1295,N_1016);
nand U1693 (N_1693,N_1319,N_1251);
nor U1694 (N_1694,N_1371,N_1223);
or U1695 (N_1695,N_1375,N_1170);
xnor U1696 (N_1696,N_1339,N_1027);
and U1697 (N_1697,N_1169,N_1087);
nand U1698 (N_1698,N_1327,N_1287);
and U1699 (N_1699,N_1086,N_1241);
and U1700 (N_1700,N_1183,N_1154);
nor U1701 (N_1701,N_1229,N_1082);
or U1702 (N_1702,N_1391,N_1046);
or U1703 (N_1703,N_1317,N_1484);
and U1704 (N_1704,N_1058,N_1220);
or U1705 (N_1705,N_1345,N_1144);
and U1706 (N_1706,N_1159,N_1348);
and U1707 (N_1707,N_1400,N_1277);
xor U1708 (N_1708,N_1426,N_1201);
nor U1709 (N_1709,N_1054,N_1265);
nand U1710 (N_1710,N_1135,N_1469);
xor U1711 (N_1711,N_1190,N_1458);
nand U1712 (N_1712,N_1470,N_1347);
and U1713 (N_1713,N_1108,N_1047);
nand U1714 (N_1714,N_1200,N_1424);
or U1715 (N_1715,N_1077,N_1041);
or U1716 (N_1716,N_1350,N_1323);
nor U1717 (N_1717,N_1360,N_1026);
or U1718 (N_1718,N_1489,N_1061);
nor U1719 (N_1719,N_1431,N_1416);
or U1720 (N_1720,N_1246,N_1418);
nor U1721 (N_1721,N_1051,N_1465);
and U1722 (N_1722,N_1372,N_1031);
nor U1723 (N_1723,N_1320,N_1110);
nor U1724 (N_1724,N_1042,N_1020);
nand U1725 (N_1725,N_1118,N_1186);
nand U1726 (N_1726,N_1441,N_1188);
xor U1727 (N_1727,N_1185,N_1482);
xnor U1728 (N_1728,N_1298,N_1079);
nand U1729 (N_1729,N_1413,N_1152);
nor U1730 (N_1730,N_1066,N_1301);
xor U1731 (N_1731,N_1052,N_1390);
nand U1732 (N_1732,N_1447,N_1308);
and U1733 (N_1733,N_1414,N_1318);
and U1734 (N_1734,N_1439,N_1285);
or U1735 (N_1735,N_1024,N_1481);
nor U1736 (N_1736,N_1364,N_1367);
nand U1737 (N_1737,N_1292,N_1485);
and U1738 (N_1738,N_1286,N_1494);
or U1739 (N_1739,N_1275,N_1436);
or U1740 (N_1740,N_1331,N_1302);
and U1741 (N_1741,N_1197,N_1210);
nor U1742 (N_1742,N_1222,N_1192);
nand U1743 (N_1743,N_1071,N_1463);
xnor U1744 (N_1744,N_1150,N_1014);
and U1745 (N_1745,N_1252,N_1206);
nor U1746 (N_1746,N_1394,N_1045);
or U1747 (N_1747,N_1261,N_1449);
or U1748 (N_1748,N_1010,N_1492);
or U1749 (N_1749,N_1383,N_1132);
and U1750 (N_1750,N_1377,N_1318);
nand U1751 (N_1751,N_1361,N_1433);
nor U1752 (N_1752,N_1434,N_1013);
and U1753 (N_1753,N_1384,N_1202);
xnor U1754 (N_1754,N_1271,N_1255);
nor U1755 (N_1755,N_1087,N_1329);
and U1756 (N_1756,N_1425,N_1331);
nor U1757 (N_1757,N_1016,N_1182);
or U1758 (N_1758,N_1154,N_1430);
and U1759 (N_1759,N_1066,N_1225);
or U1760 (N_1760,N_1432,N_1402);
or U1761 (N_1761,N_1025,N_1364);
nand U1762 (N_1762,N_1248,N_1342);
nand U1763 (N_1763,N_1009,N_1285);
nor U1764 (N_1764,N_1360,N_1271);
nor U1765 (N_1765,N_1422,N_1274);
and U1766 (N_1766,N_1367,N_1382);
nand U1767 (N_1767,N_1366,N_1006);
nor U1768 (N_1768,N_1243,N_1077);
nand U1769 (N_1769,N_1097,N_1084);
nor U1770 (N_1770,N_1051,N_1306);
nand U1771 (N_1771,N_1260,N_1056);
nor U1772 (N_1772,N_1168,N_1205);
nor U1773 (N_1773,N_1120,N_1484);
or U1774 (N_1774,N_1399,N_1413);
nor U1775 (N_1775,N_1413,N_1069);
or U1776 (N_1776,N_1346,N_1304);
nand U1777 (N_1777,N_1101,N_1424);
nand U1778 (N_1778,N_1026,N_1253);
or U1779 (N_1779,N_1478,N_1243);
nor U1780 (N_1780,N_1318,N_1049);
and U1781 (N_1781,N_1054,N_1077);
xor U1782 (N_1782,N_1340,N_1177);
xor U1783 (N_1783,N_1435,N_1496);
nand U1784 (N_1784,N_1320,N_1497);
or U1785 (N_1785,N_1401,N_1108);
nand U1786 (N_1786,N_1261,N_1457);
and U1787 (N_1787,N_1096,N_1149);
and U1788 (N_1788,N_1389,N_1265);
or U1789 (N_1789,N_1311,N_1371);
and U1790 (N_1790,N_1163,N_1330);
nor U1791 (N_1791,N_1467,N_1136);
or U1792 (N_1792,N_1027,N_1402);
nand U1793 (N_1793,N_1251,N_1273);
and U1794 (N_1794,N_1349,N_1099);
nand U1795 (N_1795,N_1352,N_1388);
nand U1796 (N_1796,N_1352,N_1219);
nor U1797 (N_1797,N_1134,N_1026);
or U1798 (N_1798,N_1449,N_1479);
xor U1799 (N_1799,N_1391,N_1459);
and U1800 (N_1800,N_1484,N_1063);
and U1801 (N_1801,N_1354,N_1096);
nor U1802 (N_1802,N_1443,N_1439);
and U1803 (N_1803,N_1185,N_1192);
nor U1804 (N_1804,N_1271,N_1353);
and U1805 (N_1805,N_1463,N_1085);
nand U1806 (N_1806,N_1182,N_1100);
or U1807 (N_1807,N_1056,N_1049);
and U1808 (N_1808,N_1228,N_1302);
nand U1809 (N_1809,N_1388,N_1273);
and U1810 (N_1810,N_1366,N_1081);
nor U1811 (N_1811,N_1290,N_1256);
or U1812 (N_1812,N_1157,N_1435);
nor U1813 (N_1813,N_1472,N_1284);
or U1814 (N_1814,N_1433,N_1382);
nand U1815 (N_1815,N_1172,N_1250);
and U1816 (N_1816,N_1196,N_1320);
or U1817 (N_1817,N_1451,N_1381);
xnor U1818 (N_1818,N_1276,N_1347);
nor U1819 (N_1819,N_1332,N_1135);
and U1820 (N_1820,N_1470,N_1272);
nor U1821 (N_1821,N_1032,N_1159);
nand U1822 (N_1822,N_1463,N_1141);
and U1823 (N_1823,N_1211,N_1452);
or U1824 (N_1824,N_1106,N_1009);
xnor U1825 (N_1825,N_1455,N_1385);
nand U1826 (N_1826,N_1205,N_1184);
and U1827 (N_1827,N_1488,N_1322);
or U1828 (N_1828,N_1337,N_1063);
or U1829 (N_1829,N_1484,N_1070);
xor U1830 (N_1830,N_1111,N_1458);
and U1831 (N_1831,N_1386,N_1184);
nand U1832 (N_1832,N_1348,N_1174);
or U1833 (N_1833,N_1490,N_1291);
nand U1834 (N_1834,N_1247,N_1185);
nand U1835 (N_1835,N_1276,N_1245);
and U1836 (N_1836,N_1451,N_1293);
nand U1837 (N_1837,N_1104,N_1413);
or U1838 (N_1838,N_1406,N_1481);
nor U1839 (N_1839,N_1178,N_1124);
xor U1840 (N_1840,N_1097,N_1026);
and U1841 (N_1841,N_1204,N_1017);
xnor U1842 (N_1842,N_1388,N_1204);
xor U1843 (N_1843,N_1459,N_1244);
or U1844 (N_1844,N_1472,N_1133);
nand U1845 (N_1845,N_1107,N_1475);
or U1846 (N_1846,N_1361,N_1178);
or U1847 (N_1847,N_1128,N_1370);
and U1848 (N_1848,N_1456,N_1448);
or U1849 (N_1849,N_1377,N_1388);
and U1850 (N_1850,N_1281,N_1246);
and U1851 (N_1851,N_1317,N_1476);
or U1852 (N_1852,N_1427,N_1343);
xor U1853 (N_1853,N_1065,N_1311);
and U1854 (N_1854,N_1185,N_1009);
and U1855 (N_1855,N_1168,N_1469);
nor U1856 (N_1856,N_1113,N_1344);
nand U1857 (N_1857,N_1414,N_1198);
nand U1858 (N_1858,N_1199,N_1417);
xnor U1859 (N_1859,N_1323,N_1106);
and U1860 (N_1860,N_1180,N_1244);
and U1861 (N_1861,N_1207,N_1069);
xnor U1862 (N_1862,N_1284,N_1096);
nor U1863 (N_1863,N_1132,N_1043);
or U1864 (N_1864,N_1489,N_1352);
xnor U1865 (N_1865,N_1172,N_1070);
xnor U1866 (N_1866,N_1242,N_1290);
and U1867 (N_1867,N_1184,N_1309);
and U1868 (N_1868,N_1212,N_1125);
or U1869 (N_1869,N_1108,N_1338);
and U1870 (N_1870,N_1222,N_1308);
nor U1871 (N_1871,N_1155,N_1413);
nor U1872 (N_1872,N_1414,N_1135);
nor U1873 (N_1873,N_1354,N_1001);
and U1874 (N_1874,N_1121,N_1342);
nand U1875 (N_1875,N_1319,N_1414);
nand U1876 (N_1876,N_1028,N_1407);
xor U1877 (N_1877,N_1057,N_1087);
nor U1878 (N_1878,N_1249,N_1343);
or U1879 (N_1879,N_1161,N_1235);
and U1880 (N_1880,N_1380,N_1119);
nor U1881 (N_1881,N_1472,N_1198);
xor U1882 (N_1882,N_1448,N_1363);
nand U1883 (N_1883,N_1473,N_1427);
nor U1884 (N_1884,N_1221,N_1204);
xor U1885 (N_1885,N_1077,N_1140);
or U1886 (N_1886,N_1415,N_1210);
xnor U1887 (N_1887,N_1459,N_1069);
nor U1888 (N_1888,N_1396,N_1159);
xnor U1889 (N_1889,N_1062,N_1236);
and U1890 (N_1890,N_1071,N_1073);
nor U1891 (N_1891,N_1148,N_1137);
xor U1892 (N_1892,N_1109,N_1453);
xor U1893 (N_1893,N_1064,N_1028);
nand U1894 (N_1894,N_1082,N_1485);
and U1895 (N_1895,N_1350,N_1389);
and U1896 (N_1896,N_1172,N_1185);
xor U1897 (N_1897,N_1081,N_1001);
nand U1898 (N_1898,N_1339,N_1401);
or U1899 (N_1899,N_1169,N_1060);
nor U1900 (N_1900,N_1260,N_1334);
nor U1901 (N_1901,N_1453,N_1402);
nand U1902 (N_1902,N_1012,N_1476);
or U1903 (N_1903,N_1180,N_1234);
nand U1904 (N_1904,N_1277,N_1480);
nor U1905 (N_1905,N_1236,N_1150);
or U1906 (N_1906,N_1217,N_1122);
and U1907 (N_1907,N_1137,N_1205);
or U1908 (N_1908,N_1001,N_1384);
nand U1909 (N_1909,N_1378,N_1008);
nor U1910 (N_1910,N_1186,N_1248);
nor U1911 (N_1911,N_1488,N_1008);
xor U1912 (N_1912,N_1312,N_1019);
nand U1913 (N_1913,N_1060,N_1254);
nor U1914 (N_1914,N_1137,N_1418);
xor U1915 (N_1915,N_1134,N_1017);
or U1916 (N_1916,N_1238,N_1015);
or U1917 (N_1917,N_1389,N_1033);
xnor U1918 (N_1918,N_1303,N_1358);
or U1919 (N_1919,N_1378,N_1135);
or U1920 (N_1920,N_1483,N_1231);
nor U1921 (N_1921,N_1021,N_1455);
nand U1922 (N_1922,N_1268,N_1031);
nand U1923 (N_1923,N_1282,N_1353);
nor U1924 (N_1924,N_1231,N_1306);
or U1925 (N_1925,N_1381,N_1423);
nand U1926 (N_1926,N_1275,N_1029);
or U1927 (N_1927,N_1468,N_1122);
xor U1928 (N_1928,N_1045,N_1211);
and U1929 (N_1929,N_1324,N_1078);
and U1930 (N_1930,N_1491,N_1470);
xnor U1931 (N_1931,N_1163,N_1328);
xor U1932 (N_1932,N_1318,N_1462);
xnor U1933 (N_1933,N_1049,N_1360);
and U1934 (N_1934,N_1275,N_1450);
or U1935 (N_1935,N_1086,N_1037);
or U1936 (N_1936,N_1187,N_1232);
nand U1937 (N_1937,N_1027,N_1139);
xnor U1938 (N_1938,N_1114,N_1153);
and U1939 (N_1939,N_1225,N_1290);
nor U1940 (N_1940,N_1131,N_1067);
and U1941 (N_1941,N_1286,N_1128);
and U1942 (N_1942,N_1344,N_1269);
nor U1943 (N_1943,N_1352,N_1459);
nor U1944 (N_1944,N_1212,N_1184);
or U1945 (N_1945,N_1351,N_1384);
xnor U1946 (N_1946,N_1191,N_1277);
nor U1947 (N_1947,N_1304,N_1077);
and U1948 (N_1948,N_1063,N_1085);
and U1949 (N_1949,N_1422,N_1363);
nand U1950 (N_1950,N_1383,N_1255);
nand U1951 (N_1951,N_1055,N_1334);
and U1952 (N_1952,N_1498,N_1060);
nand U1953 (N_1953,N_1200,N_1459);
or U1954 (N_1954,N_1297,N_1160);
nor U1955 (N_1955,N_1056,N_1064);
nand U1956 (N_1956,N_1270,N_1277);
nor U1957 (N_1957,N_1195,N_1162);
nand U1958 (N_1958,N_1482,N_1224);
nand U1959 (N_1959,N_1119,N_1298);
xnor U1960 (N_1960,N_1310,N_1300);
or U1961 (N_1961,N_1202,N_1358);
xnor U1962 (N_1962,N_1370,N_1204);
or U1963 (N_1963,N_1498,N_1027);
nor U1964 (N_1964,N_1314,N_1180);
xor U1965 (N_1965,N_1340,N_1150);
xnor U1966 (N_1966,N_1320,N_1239);
and U1967 (N_1967,N_1385,N_1180);
xor U1968 (N_1968,N_1499,N_1314);
or U1969 (N_1969,N_1418,N_1358);
nand U1970 (N_1970,N_1316,N_1243);
and U1971 (N_1971,N_1172,N_1308);
nor U1972 (N_1972,N_1049,N_1281);
or U1973 (N_1973,N_1484,N_1005);
xor U1974 (N_1974,N_1119,N_1181);
and U1975 (N_1975,N_1463,N_1163);
xor U1976 (N_1976,N_1137,N_1151);
nand U1977 (N_1977,N_1265,N_1397);
or U1978 (N_1978,N_1330,N_1005);
xor U1979 (N_1979,N_1210,N_1275);
nand U1980 (N_1980,N_1448,N_1085);
nand U1981 (N_1981,N_1383,N_1281);
xnor U1982 (N_1982,N_1156,N_1375);
xnor U1983 (N_1983,N_1293,N_1197);
and U1984 (N_1984,N_1110,N_1054);
and U1985 (N_1985,N_1113,N_1372);
or U1986 (N_1986,N_1082,N_1025);
nand U1987 (N_1987,N_1481,N_1215);
and U1988 (N_1988,N_1364,N_1276);
and U1989 (N_1989,N_1033,N_1212);
nand U1990 (N_1990,N_1326,N_1076);
xnor U1991 (N_1991,N_1217,N_1496);
or U1992 (N_1992,N_1456,N_1263);
or U1993 (N_1993,N_1406,N_1010);
and U1994 (N_1994,N_1449,N_1415);
xor U1995 (N_1995,N_1418,N_1344);
nand U1996 (N_1996,N_1216,N_1158);
or U1997 (N_1997,N_1401,N_1016);
nor U1998 (N_1998,N_1437,N_1201);
and U1999 (N_1999,N_1369,N_1312);
and U2000 (N_2000,N_1590,N_1531);
nand U2001 (N_2001,N_1581,N_1714);
xnor U2002 (N_2002,N_1579,N_1616);
or U2003 (N_2003,N_1549,N_1625);
xor U2004 (N_2004,N_1606,N_1920);
or U2005 (N_2005,N_1709,N_1659);
xnor U2006 (N_2006,N_1612,N_1726);
nand U2007 (N_2007,N_1749,N_1545);
nor U2008 (N_2008,N_1993,N_1793);
nand U2009 (N_2009,N_1780,N_1570);
or U2010 (N_2010,N_1639,N_1679);
nand U2011 (N_2011,N_1552,N_1913);
nand U2012 (N_2012,N_1719,N_1928);
nor U2013 (N_2013,N_1621,N_1853);
and U2014 (N_2014,N_1995,N_1643);
and U2015 (N_2015,N_1897,N_1828);
and U2016 (N_2016,N_1566,N_1624);
or U2017 (N_2017,N_1597,N_1670);
and U2018 (N_2018,N_1628,N_1630);
xnor U2019 (N_2019,N_1845,N_1955);
nor U2020 (N_2020,N_1971,N_1953);
or U2021 (N_2021,N_1645,N_1684);
and U2022 (N_2022,N_1803,N_1868);
xor U2023 (N_2023,N_1692,N_1596);
xor U2024 (N_2024,N_1786,N_1617);
or U2025 (N_2025,N_1686,N_1833);
and U2026 (N_2026,N_1790,N_1905);
or U2027 (N_2027,N_1843,N_1556);
and U2028 (N_2028,N_1841,N_1945);
nor U2029 (N_2029,N_1926,N_1664);
and U2030 (N_2030,N_1830,N_1798);
nor U2031 (N_2031,N_1771,N_1613);
nand U2032 (N_2032,N_1737,N_1848);
and U2033 (N_2033,N_1513,N_1998);
nand U2034 (N_2034,N_1578,N_1705);
nand U2035 (N_2035,N_1773,N_1947);
nand U2036 (N_2036,N_1862,N_1875);
and U2037 (N_2037,N_1656,N_1687);
and U2038 (N_2038,N_1846,N_1829);
nand U2039 (N_2039,N_1521,N_1909);
nor U2040 (N_2040,N_1879,N_1574);
nand U2041 (N_2041,N_1523,N_1565);
xor U2042 (N_2042,N_1535,N_1819);
xnor U2043 (N_2043,N_1682,N_1776);
nor U2044 (N_2044,N_1964,N_1525);
nor U2045 (N_2045,N_1760,N_1637);
xnor U2046 (N_2046,N_1688,N_1575);
xnor U2047 (N_2047,N_1541,N_1778);
and U2048 (N_2048,N_1915,N_1595);
nand U2049 (N_2049,N_1623,N_1599);
nor U2050 (N_2050,N_1745,N_1674);
nand U2051 (N_2051,N_1954,N_1547);
xnor U2052 (N_2052,N_1904,N_1658);
xor U2053 (N_2053,N_1816,N_1936);
nor U2054 (N_2054,N_1815,N_1660);
nand U2055 (N_2055,N_1729,N_1834);
or U2056 (N_2056,N_1885,N_1799);
and U2057 (N_2057,N_1666,N_1818);
nor U2058 (N_2058,N_1806,N_1600);
nor U2059 (N_2059,N_1896,N_1756);
nor U2060 (N_2060,N_1938,N_1584);
xnor U2061 (N_2061,N_1743,N_1580);
and U2062 (N_2062,N_1717,N_1907);
nor U2063 (N_2063,N_1949,N_1532);
xor U2064 (N_2064,N_1812,N_1638);
nor U2065 (N_2065,N_1591,N_1857);
xnor U2066 (N_2066,N_1860,N_1956);
or U2067 (N_2067,N_1622,N_1608);
xor U2068 (N_2068,N_1738,N_1943);
nand U2069 (N_2069,N_1657,N_1654);
and U2070 (N_2070,N_1510,N_1842);
xor U2071 (N_2071,N_1902,N_1516);
nor U2072 (N_2072,N_1941,N_1605);
or U2073 (N_2073,N_1859,N_1540);
nand U2074 (N_2074,N_1651,N_1661);
nand U2075 (N_2075,N_1882,N_1877);
nor U2076 (N_2076,N_1967,N_1614);
xnor U2077 (N_2077,N_1831,N_1730);
nand U2078 (N_2078,N_1937,N_1663);
xor U2079 (N_2079,N_1792,N_1800);
and U2080 (N_2080,N_1741,N_1689);
nor U2081 (N_2081,N_1539,N_1672);
and U2082 (N_2082,N_1988,N_1631);
nor U2083 (N_2083,N_1512,N_1876);
or U2084 (N_2084,N_1784,N_1935);
nor U2085 (N_2085,N_1675,N_1804);
or U2086 (N_2086,N_1867,N_1808);
nor U2087 (N_2087,N_1888,N_1986);
and U2088 (N_2088,N_1711,N_1871);
xor U2089 (N_2089,N_1783,N_1923);
or U2090 (N_2090,N_1946,N_1940);
xnor U2091 (N_2091,N_1589,N_1921);
and U2092 (N_2092,N_1872,N_1568);
xnor U2093 (N_2093,N_1603,N_1914);
and U2094 (N_2094,N_1824,N_1980);
nor U2095 (N_2095,N_1996,N_1891);
xnor U2096 (N_2096,N_1615,N_1640);
or U2097 (N_2097,N_1973,N_1823);
or U2098 (N_2098,N_1899,N_1735);
and U2099 (N_2099,N_1634,N_1985);
or U2100 (N_2100,N_1524,N_1744);
nor U2101 (N_2101,N_1644,N_1633);
xor U2102 (N_2102,N_1901,N_1538);
or U2103 (N_2103,N_1752,N_1894);
nor U2104 (N_2104,N_1536,N_1677);
and U2105 (N_2105,N_1856,N_1832);
nand U2106 (N_2106,N_1777,N_1759);
nand U2107 (N_2107,N_1567,N_1765);
or U2108 (N_2108,N_1895,N_1713);
or U2109 (N_2109,N_1557,N_1981);
nand U2110 (N_2110,N_1725,N_1917);
and U2111 (N_2111,N_1683,N_1821);
and U2112 (N_2112,N_1836,N_1855);
xnor U2113 (N_2113,N_1721,N_1802);
nand U2114 (N_2114,N_1609,N_1788);
and U2115 (N_2115,N_1933,N_1839);
or U2116 (N_2116,N_1647,N_1911);
nand U2117 (N_2117,N_1572,N_1553);
and U2118 (N_2118,N_1963,N_1690);
and U2119 (N_2119,N_1602,N_1969);
nand U2120 (N_2120,N_1555,N_1662);
nor U2121 (N_2121,N_1811,N_1626);
and U2122 (N_2122,N_1794,N_1700);
xnor U2123 (N_2123,N_1585,N_1671);
nand U2124 (N_2124,N_1970,N_1766);
nand U2125 (N_2125,N_1515,N_1518);
nor U2126 (N_2126,N_1542,N_1910);
nor U2127 (N_2127,N_1680,N_1850);
nand U2128 (N_2128,N_1734,N_1870);
and U2129 (N_2129,N_1837,N_1987);
and U2130 (N_2130,N_1789,N_1653);
or U2131 (N_2131,N_1546,N_1912);
nand U2132 (N_2132,N_1560,N_1931);
nand U2133 (N_2133,N_1736,N_1758);
or U2134 (N_2134,N_1797,N_1810);
xor U2135 (N_2135,N_1762,N_1880);
xor U2136 (N_2136,N_1708,N_1866);
and U2137 (N_2137,N_1695,N_1724);
nor U2138 (N_2138,N_1696,N_1618);
xor U2139 (N_2139,N_1932,N_1764);
nor U2140 (N_2140,N_1983,N_1611);
nand U2141 (N_2141,N_1503,N_1972);
xnor U2142 (N_2142,N_1874,N_1667);
nor U2143 (N_2143,N_1976,N_1534);
and U2144 (N_2144,N_1573,N_1959);
and U2145 (N_2145,N_1785,N_1727);
nor U2146 (N_2146,N_1522,N_1991);
or U2147 (N_2147,N_1903,N_1883);
xnor U2148 (N_2148,N_1769,N_1801);
and U2149 (N_2149,N_1500,N_1641);
nor U2150 (N_2150,N_1962,N_1728);
or U2151 (N_2151,N_1636,N_1607);
xor U2152 (N_2152,N_1648,N_1997);
xnor U2153 (N_2153,N_1893,N_1886);
xor U2154 (N_2154,N_1772,N_1509);
nor U2155 (N_2155,N_1506,N_1554);
nor U2156 (N_2156,N_1873,N_1982);
nand U2157 (N_2157,N_1994,N_1968);
and U2158 (N_2158,N_1582,N_1533);
or U2159 (N_2159,N_1739,N_1588);
xor U2160 (N_2160,N_1564,N_1770);
and U2161 (N_2161,N_1517,N_1558);
and U2162 (N_2162,N_1961,N_1592);
nor U2163 (N_2163,N_1809,N_1577);
and U2164 (N_2164,N_1852,N_1586);
or U2165 (N_2165,N_1977,N_1748);
xnor U2166 (N_2166,N_1703,N_1723);
xnor U2167 (N_2167,N_1960,N_1782);
nand U2168 (N_2168,N_1571,N_1520);
nor U2169 (N_2169,N_1537,N_1864);
nand U2170 (N_2170,N_1889,N_1665);
nand U2171 (N_2171,N_1733,N_1863);
nor U2172 (N_2172,N_1732,N_1712);
or U2173 (N_2173,N_1508,N_1747);
xnor U2174 (N_2174,N_1598,N_1898);
xor U2175 (N_2175,N_1668,N_1562);
xor U2176 (N_2176,N_1501,N_1918);
and U2177 (N_2177,N_1827,N_1858);
nor U2178 (N_2178,N_1559,N_1774);
and U2179 (N_2179,N_1543,N_1502);
nand U2180 (N_2180,N_1551,N_1822);
nand U2181 (N_2181,N_1881,N_1906);
nand U2182 (N_2182,N_1849,N_1763);
and U2183 (N_2183,N_1865,N_1563);
nand U2184 (N_2184,N_1924,N_1927);
or U2185 (N_2185,N_1706,N_1887);
and U2186 (N_2186,N_1978,N_1673);
xnor U2187 (N_2187,N_1740,N_1681);
nor U2188 (N_2188,N_1781,N_1957);
nor U2189 (N_2189,N_1699,N_1878);
xor U2190 (N_2190,N_1929,N_1805);
nand U2191 (N_2191,N_1835,N_1627);
or U2192 (N_2192,N_1975,N_1505);
or U2193 (N_2193,N_1755,N_1576);
or U2194 (N_2194,N_1948,N_1847);
nand U2195 (N_2195,N_1807,N_1750);
xor U2196 (N_2196,N_1796,N_1610);
or U2197 (N_2197,N_1594,N_1814);
and U2198 (N_2198,N_1619,N_1820);
and U2199 (N_2199,N_1925,N_1694);
xor U2200 (N_2200,N_1916,N_1840);
or U2201 (N_2201,N_1649,N_1958);
nand U2202 (N_2202,N_1685,N_1569);
nand U2203 (N_2203,N_1722,N_1702);
xor U2204 (N_2204,N_1838,N_1950);
nor U2205 (N_2205,N_1952,N_1791);
nand U2206 (N_2206,N_1544,N_1951);
and U2207 (N_2207,N_1718,N_1742);
or U2208 (N_2208,N_1751,N_1731);
nor U2209 (N_2209,N_1892,N_1922);
or U2210 (N_2210,N_1691,N_1698);
or U2211 (N_2211,N_1635,N_1548);
nor U2212 (N_2212,N_1825,N_1908);
nand U2213 (N_2213,N_1519,N_1966);
or U2214 (N_2214,N_1795,N_1530);
nand U2215 (N_2215,N_1919,N_1704);
or U2216 (N_2216,N_1990,N_1779);
nor U2217 (N_2217,N_1989,N_1707);
nand U2218 (N_2218,N_1620,N_1817);
or U2219 (N_2219,N_1854,N_1550);
xnor U2220 (N_2220,N_1561,N_1720);
nor U2221 (N_2221,N_1944,N_1884);
and U2222 (N_2222,N_1753,N_1642);
and U2223 (N_2223,N_1851,N_1527);
xnor U2224 (N_2224,N_1604,N_1593);
xor U2225 (N_2225,N_1992,N_1930);
xor U2226 (N_2226,N_1526,N_1676);
nor U2227 (N_2227,N_1775,N_1601);
nor U2228 (N_2228,N_1746,N_1701);
nor U2229 (N_2229,N_1629,N_1869);
nand U2230 (N_2230,N_1984,N_1979);
nand U2231 (N_2231,N_1787,N_1826);
or U2232 (N_2232,N_1890,N_1767);
xor U2233 (N_2233,N_1999,N_1965);
nand U2234 (N_2234,N_1710,N_1761);
and U2235 (N_2235,N_1583,N_1646);
nand U2236 (N_2236,N_1504,N_1697);
or U2237 (N_2237,N_1813,N_1900);
xnor U2238 (N_2238,N_1844,N_1528);
xor U2239 (N_2239,N_1511,N_1715);
xor U2240 (N_2240,N_1587,N_1974);
xor U2241 (N_2241,N_1716,N_1678);
or U2242 (N_2242,N_1754,N_1669);
and U2243 (N_2243,N_1514,N_1507);
and U2244 (N_2244,N_1652,N_1934);
nor U2245 (N_2245,N_1768,N_1861);
or U2246 (N_2246,N_1655,N_1632);
nor U2247 (N_2247,N_1693,N_1939);
or U2248 (N_2248,N_1529,N_1942);
xor U2249 (N_2249,N_1757,N_1650);
or U2250 (N_2250,N_1800,N_1505);
xnor U2251 (N_2251,N_1552,N_1894);
and U2252 (N_2252,N_1781,N_1580);
and U2253 (N_2253,N_1890,N_1776);
or U2254 (N_2254,N_1921,N_1532);
xor U2255 (N_2255,N_1839,N_1791);
nor U2256 (N_2256,N_1544,N_1514);
xnor U2257 (N_2257,N_1813,N_1669);
or U2258 (N_2258,N_1758,N_1917);
xor U2259 (N_2259,N_1689,N_1966);
nand U2260 (N_2260,N_1880,N_1640);
nand U2261 (N_2261,N_1894,N_1976);
xnor U2262 (N_2262,N_1513,N_1826);
nand U2263 (N_2263,N_1655,N_1843);
xor U2264 (N_2264,N_1513,N_1681);
nand U2265 (N_2265,N_1924,N_1874);
xor U2266 (N_2266,N_1690,N_1589);
nand U2267 (N_2267,N_1614,N_1679);
and U2268 (N_2268,N_1971,N_1649);
nand U2269 (N_2269,N_1611,N_1675);
and U2270 (N_2270,N_1539,N_1608);
nor U2271 (N_2271,N_1903,N_1660);
or U2272 (N_2272,N_1946,N_1774);
and U2273 (N_2273,N_1960,N_1542);
xnor U2274 (N_2274,N_1664,N_1546);
nor U2275 (N_2275,N_1880,N_1969);
or U2276 (N_2276,N_1895,N_1727);
nand U2277 (N_2277,N_1987,N_1963);
nand U2278 (N_2278,N_1885,N_1626);
nand U2279 (N_2279,N_1870,N_1997);
xor U2280 (N_2280,N_1629,N_1825);
nand U2281 (N_2281,N_1855,N_1528);
nor U2282 (N_2282,N_1660,N_1936);
nor U2283 (N_2283,N_1543,N_1998);
or U2284 (N_2284,N_1928,N_1545);
nand U2285 (N_2285,N_1784,N_1592);
and U2286 (N_2286,N_1562,N_1630);
xor U2287 (N_2287,N_1554,N_1827);
xor U2288 (N_2288,N_1677,N_1990);
or U2289 (N_2289,N_1996,N_1838);
nor U2290 (N_2290,N_1909,N_1547);
nand U2291 (N_2291,N_1844,N_1912);
and U2292 (N_2292,N_1880,N_1643);
and U2293 (N_2293,N_1665,N_1626);
nor U2294 (N_2294,N_1914,N_1583);
and U2295 (N_2295,N_1665,N_1633);
or U2296 (N_2296,N_1781,N_1796);
nor U2297 (N_2297,N_1689,N_1828);
xnor U2298 (N_2298,N_1567,N_1611);
nand U2299 (N_2299,N_1848,N_1630);
and U2300 (N_2300,N_1728,N_1970);
or U2301 (N_2301,N_1964,N_1609);
and U2302 (N_2302,N_1786,N_1917);
or U2303 (N_2303,N_1966,N_1642);
nand U2304 (N_2304,N_1641,N_1502);
or U2305 (N_2305,N_1511,N_1927);
nor U2306 (N_2306,N_1567,N_1755);
nor U2307 (N_2307,N_1983,N_1845);
xor U2308 (N_2308,N_1786,N_1559);
nor U2309 (N_2309,N_1884,N_1770);
nand U2310 (N_2310,N_1720,N_1732);
or U2311 (N_2311,N_1586,N_1743);
nor U2312 (N_2312,N_1904,N_1764);
or U2313 (N_2313,N_1867,N_1761);
nor U2314 (N_2314,N_1771,N_1986);
nor U2315 (N_2315,N_1816,N_1970);
and U2316 (N_2316,N_1978,N_1876);
nor U2317 (N_2317,N_1739,N_1655);
and U2318 (N_2318,N_1651,N_1749);
or U2319 (N_2319,N_1716,N_1858);
xor U2320 (N_2320,N_1519,N_1704);
xnor U2321 (N_2321,N_1830,N_1802);
and U2322 (N_2322,N_1563,N_1961);
and U2323 (N_2323,N_1747,N_1517);
xnor U2324 (N_2324,N_1552,N_1891);
nand U2325 (N_2325,N_1663,N_1853);
nor U2326 (N_2326,N_1901,N_1676);
nand U2327 (N_2327,N_1964,N_1565);
or U2328 (N_2328,N_1643,N_1554);
or U2329 (N_2329,N_1521,N_1605);
nand U2330 (N_2330,N_1724,N_1950);
or U2331 (N_2331,N_1848,N_1869);
nand U2332 (N_2332,N_1543,N_1828);
nor U2333 (N_2333,N_1588,N_1810);
nand U2334 (N_2334,N_1830,N_1912);
or U2335 (N_2335,N_1553,N_1591);
and U2336 (N_2336,N_1669,N_1824);
or U2337 (N_2337,N_1582,N_1975);
or U2338 (N_2338,N_1838,N_1676);
and U2339 (N_2339,N_1893,N_1950);
nor U2340 (N_2340,N_1916,N_1599);
or U2341 (N_2341,N_1876,N_1867);
and U2342 (N_2342,N_1936,N_1652);
and U2343 (N_2343,N_1516,N_1852);
or U2344 (N_2344,N_1927,N_1507);
nand U2345 (N_2345,N_1595,N_1783);
and U2346 (N_2346,N_1849,N_1624);
and U2347 (N_2347,N_1886,N_1791);
or U2348 (N_2348,N_1571,N_1518);
and U2349 (N_2349,N_1792,N_1909);
and U2350 (N_2350,N_1751,N_1770);
or U2351 (N_2351,N_1925,N_1870);
xor U2352 (N_2352,N_1739,N_1820);
or U2353 (N_2353,N_1925,N_1837);
xnor U2354 (N_2354,N_1593,N_1818);
nand U2355 (N_2355,N_1580,N_1947);
nand U2356 (N_2356,N_1649,N_1892);
or U2357 (N_2357,N_1923,N_1805);
nor U2358 (N_2358,N_1842,N_1831);
and U2359 (N_2359,N_1878,N_1943);
nor U2360 (N_2360,N_1612,N_1505);
and U2361 (N_2361,N_1832,N_1890);
nor U2362 (N_2362,N_1630,N_1808);
and U2363 (N_2363,N_1933,N_1538);
nor U2364 (N_2364,N_1699,N_1961);
nor U2365 (N_2365,N_1848,N_1999);
and U2366 (N_2366,N_1957,N_1519);
nand U2367 (N_2367,N_1720,N_1661);
or U2368 (N_2368,N_1779,N_1516);
xor U2369 (N_2369,N_1871,N_1601);
xor U2370 (N_2370,N_1928,N_1933);
nor U2371 (N_2371,N_1757,N_1880);
or U2372 (N_2372,N_1589,N_1883);
nor U2373 (N_2373,N_1910,N_1921);
nor U2374 (N_2374,N_1725,N_1743);
and U2375 (N_2375,N_1986,N_1556);
and U2376 (N_2376,N_1860,N_1644);
nor U2377 (N_2377,N_1736,N_1869);
nor U2378 (N_2378,N_1728,N_1556);
nand U2379 (N_2379,N_1961,N_1534);
or U2380 (N_2380,N_1834,N_1568);
xor U2381 (N_2381,N_1945,N_1623);
xnor U2382 (N_2382,N_1624,N_1857);
nand U2383 (N_2383,N_1689,N_1808);
nor U2384 (N_2384,N_1549,N_1680);
nand U2385 (N_2385,N_1877,N_1786);
nor U2386 (N_2386,N_1845,N_1924);
nand U2387 (N_2387,N_1537,N_1996);
and U2388 (N_2388,N_1510,N_1893);
nor U2389 (N_2389,N_1536,N_1643);
and U2390 (N_2390,N_1872,N_1847);
nor U2391 (N_2391,N_1652,N_1536);
nor U2392 (N_2392,N_1914,N_1968);
and U2393 (N_2393,N_1870,N_1809);
nor U2394 (N_2394,N_1710,N_1774);
xnor U2395 (N_2395,N_1853,N_1682);
or U2396 (N_2396,N_1592,N_1770);
or U2397 (N_2397,N_1547,N_1688);
or U2398 (N_2398,N_1649,N_1682);
and U2399 (N_2399,N_1971,N_1681);
nor U2400 (N_2400,N_1733,N_1621);
nor U2401 (N_2401,N_1832,N_1969);
nor U2402 (N_2402,N_1655,N_1963);
nor U2403 (N_2403,N_1964,N_1607);
xnor U2404 (N_2404,N_1834,N_1790);
or U2405 (N_2405,N_1734,N_1772);
or U2406 (N_2406,N_1823,N_1507);
xnor U2407 (N_2407,N_1906,N_1827);
and U2408 (N_2408,N_1895,N_1629);
or U2409 (N_2409,N_1860,N_1841);
xnor U2410 (N_2410,N_1554,N_1994);
nor U2411 (N_2411,N_1823,N_1675);
nand U2412 (N_2412,N_1857,N_1759);
or U2413 (N_2413,N_1682,N_1832);
and U2414 (N_2414,N_1818,N_1589);
nand U2415 (N_2415,N_1882,N_1988);
or U2416 (N_2416,N_1903,N_1811);
nand U2417 (N_2417,N_1821,N_1904);
nand U2418 (N_2418,N_1618,N_1990);
xor U2419 (N_2419,N_1667,N_1811);
and U2420 (N_2420,N_1635,N_1717);
or U2421 (N_2421,N_1872,N_1586);
or U2422 (N_2422,N_1895,N_1953);
xor U2423 (N_2423,N_1570,N_1601);
nor U2424 (N_2424,N_1924,N_1613);
nor U2425 (N_2425,N_1583,N_1864);
or U2426 (N_2426,N_1929,N_1920);
nand U2427 (N_2427,N_1833,N_1838);
nor U2428 (N_2428,N_1973,N_1539);
nand U2429 (N_2429,N_1976,N_1822);
and U2430 (N_2430,N_1628,N_1814);
xor U2431 (N_2431,N_1991,N_1754);
and U2432 (N_2432,N_1669,N_1656);
nand U2433 (N_2433,N_1851,N_1712);
and U2434 (N_2434,N_1673,N_1509);
or U2435 (N_2435,N_1893,N_1734);
or U2436 (N_2436,N_1900,N_1525);
xor U2437 (N_2437,N_1674,N_1857);
or U2438 (N_2438,N_1883,N_1906);
nor U2439 (N_2439,N_1582,N_1585);
xor U2440 (N_2440,N_1510,N_1931);
or U2441 (N_2441,N_1953,N_1962);
xor U2442 (N_2442,N_1685,N_1519);
nor U2443 (N_2443,N_1706,N_1805);
nor U2444 (N_2444,N_1784,N_1516);
or U2445 (N_2445,N_1735,N_1834);
nand U2446 (N_2446,N_1512,N_1743);
or U2447 (N_2447,N_1978,N_1989);
or U2448 (N_2448,N_1675,N_1581);
nand U2449 (N_2449,N_1542,N_1626);
or U2450 (N_2450,N_1805,N_1815);
or U2451 (N_2451,N_1643,N_1953);
and U2452 (N_2452,N_1852,N_1538);
and U2453 (N_2453,N_1822,N_1579);
xnor U2454 (N_2454,N_1841,N_1983);
xnor U2455 (N_2455,N_1999,N_1917);
and U2456 (N_2456,N_1842,N_1678);
and U2457 (N_2457,N_1726,N_1757);
and U2458 (N_2458,N_1802,N_1926);
nand U2459 (N_2459,N_1983,N_1507);
and U2460 (N_2460,N_1578,N_1814);
and U2461 (N_2461,N_1893,N_1773);
nand U2462 (N_2462,N_1696,N_1867);
xnor U2463 (N_2463,N_1538,N_1771);
nand U2464 (N_2464,N_1861,N_1701);
nand U2465 (N_2465,N_1836,N_1503);
nand U2466 (N_2466,N_1747,N_1704);
or U2467 (N_2467,N_1949,N_1587);
xor U2468 (N_2468,N_1785,N_1804);
xnor U2469 (N_2469,N_1544,N_1537);
or U2470 (N_2470,N_1603,N_1859);
and U2471 (N_2471,N_1682,N_1756);
or U2472 (N_2472,N_1605,N_1569);
xor U2473 (N_2473,N_1803,N_1520);
nor U2474 (N_2474,N_1812,N_1800);
nand U2475 (N_2475,N_1610,N_1812);
xor U2476 (N_2476,N_1606,N_1767);
and U2477 (N_2477,N_1954,N_1949);
xnor U2478 (N_2478,N_1587,N_1709);
xnor U2479 (N_2479,N_1966,N_1896);
nor U2480 (N_2480,N_1843,N_1937);
and U2481 (N_2481,N_1621,N_1551);
nor U2482 (N_2482,N_1972,N_1940);
nand U2483 (N_2483,N_1810,N_1547);
and U2484 (N_2484,N_1576,N_1599);
nand U2485 (N_2485,N_1816,N_1508);
nor U2486 (N_2486,N_1941,N_1643);
nand U2487 (N_2487,N_1973,N_1860);
xor U2488 (N_2488,N_1875,N_1941);
xor U2489 (N_2489,N_1716,N_1996);
nand U2490 (N_2490,N_1772,N_1808);
xnor U2491 (N_2491,N_1889,N_1556);
nand U2492 (N_2492,N_1839,N_1948);
nand U2493 (N_2493,N_1901,N_1925);
nand U2494 (N_2494,N_1656,N_1751);
nand U2495 (N_2495,N_1670,N_1777);
nor U2496 (N_2496,N_1640,N_1507);
or U2497 (N_2497,N_1547,N_1686);
xor U2498 (N_2498,N_1919,N_1645);
nor U2499 (N_2499,N_1536,N_1602);
and U2500 (N_2500,N_2397,N_2322);
and U2501 (N_2501,N_2245,N_2039);
nand U2502 (N_2502,N_2361,N_2035);
and U2503 (N_2503,N_2020,N_2115);
nand U2504 (N_2504,N_2244,N_2295);
or U2505 (N_2505,N_2183,N_2284);
xnor U2506 (N_2506,N_2427,N_2433);
nand U2507 (N_2507,N_2242,N_2168);
or U2508 (N_2508,N_2184,N_2356);
nor U2509 (N_2509,N_2089,N_2112);
xor U2510 (N_2510,N_2457,N_2252);
nand U2511 (N_2511,N_2493,N_2166);
and U2512 (N_2512,N_2359,N_2179);
nor U2513 (N_2513,N_2008,N_2111);
and U2514 (N_2514,N_2419,N_2446);
nor U2515 (N_2515,N_2213,N_2299);
or U2516 (N_2516,N_2309,N_2262);
nand U2517 (N_2517,N_2297,N_2260);
and U2518 (N_2518,N_2498,N_2456);
and U2519 (N_2519,N_2234,N_2033);
xor U2520 (N_2520,N_2018,N_2449);
nor U2521 (N_2521,N_2411,N_2134);
or U2522 (N_2522,N_2474,N_2060);
nand U2523 (N_2523,N_2492,N_2478);
nor U2524 (N_2524,N_2384,N_2014);
and U2525 (N_2525,N_2116,N_2318);
nor U2526 (N_2526,N_2348,N_2197);
xor U2527 (N_2527,N_2317,N_2365);
nand U2528 (N_2528,N_2142,N_2338);
xor U2529 (N_2529,N_2231,N_2430);
or U2530 (N_2530,N_2432,N_2188);
or U2531 (N_2531,N_2203,N_2319);
nor U2532 (N_2532,N_2403,N_2340);
nor U2533 (N_2533,N_2472,N_2378);
nand U2534 (N_2534,N_2047,N_2294);
or U2535 (N_2535,N_2323,N_2335);
nor U2536 (N_2536,N_2311,N_2256);
or U2537 (N_2537,N_2199,N_2337);
and U2538 (N_2538,N_2350,N_2225);
and U2539 (N_2539,N_2095,N_2010);
nor U2540 (N_2540,N_2494,N_2296);
or U2541 (N_2541,N_2125,N_2367);
nor U2542 (N_2542,N_2431,N_2212);
nor U2543 (N_2543,N_2172,N_2285);
xnor U2544 (N_2544,N_2450,N_2394);
nand U2545 (N_2545,N_2163,N_2391);
xor U2546 (N_2546,N_2438,N_2281);
and U2547 (N_2547,N_2036,N_2000);
nor U2548 (N_2548,N_2117,N_2380);
nand U2549 (N_2549,N_2287,N_2342);
nor U2550 (N_2550,N_2255,N_2050);
xnor U2551 (N_2551,N_2436,N_2371);
and U2552 (N_2552,N_2270,N_2028);
nand U2553 (N_2553,N_2088,N_2085);
or U2554 (N_2554,N_2370,N_2488);
or U2555 (N_2555,N_2237,N_2227);
nand U2556 (N_2556,N_2043,N_2171);
xor U2557 (N_2557,N_2402,N_2407);
xor U2558 (N_2558,N_2150,N_2071);
and U2559 (N_2559,N_2290,N_2249);
xnor U2560 (N_2560,N_2375,N_2462);
and U2561 (N_2561,N_2004,N_2248);
nor U2562 (N_2562,N_2169,N_2413);
xnor U2563 (N_2563,N_2268,N_2235);
nor U2564 (N_2564,N_2420,N_2229);
nor U2565 (N_2565,N_2025,N_2329);
xor U2566 (N_2566,N_2289,N_2392);
xnor U2567 (N_2567,N_2483,N_2122);
nor U2568 (N_2568,N_2360,N_2209);
xor U2569 (N_2569,N_2276,N_2222);
xnor U2570 (N_2570,N_2239,N_2190);
xnor U2571 (N_2571,N_2351,N_2224);
nor U2572 (N_2572,N_2137,N_2343);
xor U2573 (N_2573,N_2286,N_2045);
nor U2574 (N_2574,N_2062,N_2021);
nor U2575 (N_2575,N_2486,N_2046);
nor U2576 (N_2576,N_2410,N_2448);
or U2577 (N_2577,N_2321,N_2455);
nor U2578 (N_2578,N_2056,N_2019);
nor U2579 (N_2579,N_2186,N_2477);
and U2580 (N_2580,N_2135,N_2292);
nand U2581 (N_2581,N_2463,N_2110);
or U2582 (N_2582,N_2422,N_2073);
xnor U2583 (N_2583,N_2029,N_2086);
nand U2584 (N_2584,N_2167,N_2467);
nand U2585 (N_2585,N_2324,N_2133);
or U2586 (N_2586,N_2230,N_2312);
xnor U2587 (N_2587,N_2158,N_2013);
or U2588 (N_2588,N_2087,N_2444);
nand U2589 (N_2589,N_2083,N_2246);
and U2590 (N_2590,N_2121,N_2288);
nand U2591 (N_2591,N_2228,N_2310);
nor U2592 (N_2592,N_2194,N_2416);
xnor U2593 (N_2593,N_2044,N_2423);
xnor U2594 (N_2594,N_2373,N_2017);
or U2595 (N_2595,N_2193,N_2070);
nand U2596 (N_2596,N_2182,N_2064);
nand U2597 (N_2597,N_2489,N_2440);
xor U2598 (N_2598,N_2024,N_2108);
or U2599 (N_2599,N_2173,N_2068);
nand U2600 (N_2600,N_2041,N_2439);
nand U2601 (N_2601,N_2481,N_2156);
nand U2602 (N_2602,N_2105,N_2215);
nor U2603 (N_2603,N_2057,N_2098);
xor U2604 (N_2604,N_2100,N_2140);
nor U2605 (N_2605,N_2253,N_2065);
and U2606 (N_2606,N_2376,N_2031);
or U2607 (N_2607,N_2325,N_2495);
xor U2608 (N_2608,N_2153,N_2139);
xor U2609 (N_2609,N_2442,N_2251);
or U2610 (N_2610,N_2372,N_2366);
nor U2611 (N_2611,N_2097,N_2174);
or U2612 (N_2612,N_2464,N_2302);
and U2613 (N_2613,N_2145,N_2077);
nor U2614 (N_2614,N_2265,N_2141);
xnor U2615 (N_2615,N_2460,N_2195);
nor U2616 (N_2616,N_2303,N_2447);
or U2617 (N_2617,N_2126,N_2395);
xnor U2618 (N_2618,N_2192,N_2272);
xnor U2619 (N_2619,N_2331,N_2084);
and U2620 (N_2620,N_2434,N_2369);
nor U2621 (N_2621,N_2119,N_2149);
or U2622 (N_2622,N_2226,N_2345);
nand U2623 (N_2623,N_2067,N_2362);
xnor U2624 (N_2624,N_2114,N_2473);
or U2625 (N_2625,N_2469,N_2206);
and U2626 (N_2626,N_2291,N_2408);
nand U2627 (N_2627,N_2424,N_2468);
and U2628 (N_2628,N_2154,N_2274);
xor U2629 (N_2629,N_2401,N_2279);
and U2630 (N_2630,N_2232,N_2339);
nand U2631 (N_2631,N_2214,N_2298);
or U2632 (N_2632,N_2128,N_2006);
nor U2633 (N_2633,N_2189,N_2336);
nor U2634 (N_2634,N_2211,N_2470);
and U2635 (N_2635,N_2306,N_2143);
nor U2636 (N_2636,N_2264,N_2208);
nand U2637 (N_2637,N_2104,N_2418);
and U2638 (N_2638,N_2081,N_2353);
nor U2639 (N_2639,N_2146,N_2103);
nand U2640 (N_2640,N_2058,N_2344);
and U2641 (N_2641,N_2417,N_2405);
and U2642 (N_2642,N_2012,N_2181);
and U2643 (N_2643,N_2162,N_2451);
or U2644 (N_2644,N_2147,N_2130);
xnor U2645 (N_2645,N_2155,N_2328);
xor U2646 (N_2646,N_2106,N_2038);
or U2647 (N_2647,N_2437,N_2254);
or U2648 (N_2648,N_2053,N_2009);
and U2649 (N_2649,N_2175,N_2374);
and U2650 (N_2650,N_2113,N_2091);
nor U2651 (N_2651,N_2461,N_2412);
nor U2652 (N_2652,N_2385,N_2015);
or U2653 (N_2653,N_2129,N_2198);
xnor U2654 (N_2654,N_2003,N_2051);
nor U2655 (N_2655,N_2352,N_2393);
xnor U2656 (N_2656,N_2032,N_2377);
nor U2657 (N_2657,N_2148,N_2123);
nand U2658 (N_2658,N_2280,N_2426);
xor U2659 (N_2659,N_2157,N_2210);
and U2660 (N_2660,N_2204,N_2334);
nand U2661 (N_2661,N_2102,N_2421);
or U2662 (N_2662,N_2136,N_2487);
and U2663 (N_2663,N_2454,N_2005);
xor U2664 (N_2664,N_2308,N_2409);
nand U2665 (N_2665,N_2435,N_2497);
and U2666 (N_2666,N_2466,N_2109);
xor U2667 (N_2667,N_2452,N_2459);
nand U2668 (N_2668,N_2042,N_2026);
nor U2669 (N_2669,N_2072,N_2159);
xor U2670 (N_2670,N_2207,N_2316);
nand U2671 (N_2671,N_2482,N_2066);
nand U2672 (N_2672,N_2022,N_2161);
nand U2673 (N_2673,N_2002,N_2074);
and U2674 (N_2674,N_2093,N_2263);
or U2675 (N_2675,N_2250,N_2386);
or U2676 (N_2676,N_2282,N_2273);
and U2677 (N_2677,N_2034,N_2101);
and U2678 (N_2678,N_2221,N_2120);
and U2679 (N_2679,N_2082,N_2180);
and U2680 (N_2680,N_2277,N_2379);
xnor U2681 (N_2681,N_2247,N_2138);
and U2682 (N_2682,N_2382,N_2202);
xor U2683 (N_2683,N_2445,N_2368);
or U2684 (N_2684,N_2011,N_2096);
nor U2685 (N_2685,N_2388,N_2076);
or U2686 (N_2686,N_2132,N_2267);
nor U2687 (N_2687,N_2314,N_2381);
and U2688 (N_2688,N_2383,N_2363);
xor U2689 (N_2689,N_2040,N_2326);
nand U2690 (N_2690,N_2216,N_2052);
nor U2691 (N_2691,N_2293,N_2355);
xor U2692 (N_2692,N_2200,N_2001);
nand U2693 (N_2693,N_2443,N_2164);
and U2694 (N_2694,N_2075,N_2217);
nand U2695 (N_2695,N_2429,N_2465);
xnor U2696 (N_2696,N_2398,N_2332);
or U2697 (N_2697,N_2485,N_2305);
and U2698 (N_2698,N_2107,N_2220);
nand U2699 (N_2699,N_2400,N_2484);
nor U2700 (N_2700,N_2144,N_2257);
xor U2701 (N_2701,N_2307,N_2118);
nand U2702 (N_2702,N_2030,N_2389);
or U2703 (N_2703,N_2069,N_2349);
or U2704 (N_2704,N_2358,N_2201);
nand U2705 (N_2705,N_2387,N_2300);
or U2706 (N_2706,N_2415,N_2238);
and U2707 (N_2707,N_2491,N_2414);
nor U2708 (N_2708,N_2425,N_2177);
nor U2709 (N_2709,N_2357,N_2079);
nor U2710 (N_2710,N_2131,N_2261);
nor U2711 (N_2711,N_2341,N_2480);
nor U2712 (N_2712,N_2490,N_2266);
or U2713 (N_2713,N_2278,N_2048);
nor U2714 (N_2714,N_2320,N_2259);
nor U2715 (N_2715,N_2016,N_2094);
nor U2716 (N_2716,N_2218,N_2269);
and U2717 (N_2717,N_2205,N_2037);
nor U2718 (N_2718,N_2099,N_2406);
and U2719 (N_2719,N_2313,N_2476);
and U2720 (N_2720,N_2327,N_2223);
and U2721 (N_2721,N_2152,N_2428);
and U2722 (N_2722,N_2023,N_2258);
and U2723 (N_2723,N_2007,N_2176);
and U2724 (N_2724,N_2301,N_2347);
nand U2725 (N_2725,N_2055,N_2499);
and U2726 (N_2726,N_2364,N_2054);
nor U2727 (N_2727,N_2092,N_2160);
and U2728 (N_2728,N_2049,N_2346);
nand U2729 (N_2729,N_2191,N_2304);
nand U2730 (N_2730,N_2441,N_2453);
or U2731 (N_2731,N_2127,N_2275);
or U2732 (N_2732,N_2315,N_2271);
xor U2733 (N_2733,N_2399,N_2185);
xor U2734 (N_2734,N_2187,N_2063);
xnor U2735 (N_2735,N_2458,N_2061);
and U2736 (N_2736,N_2496,N_2390);
or U2737 (N_2737,N_2027,N_2233);
or U2738 (N_2738,N_2471,N_2078);
nor U2739 (N_2739,N_2165,N_2475);
nor U2740 (N_2740,N_2170,N_2241);
nor U2741 (N_2741,N_2396,N_2243);
and U2742 (N_2742,N_2404,N_2059);
xnor U2743 (N_2743,N_2354,N_2219);
nand U2744 (N_2744,N_2479,N_2090);
xnor U2745 (N_2745,N_2080,N_2196);
and U2746 (N_2746,N_2240,N_2333);
xnor U2747 (N_2747,N_2330,N_2283);
nor U2748 (N_2748,N_2178,N_2124);
nor U2749 (N_2749,N_2151,N_2236);
nor U2750 (N_2750,N_2064,N_2149);
xnor U2751 (N_2751,N_2489,N_2038);
or U2752 (N_2752,N_2224,N_2049);
nand U2753 (N_2753,N_2415,N_2180);
xor U2754 (N_2754,N_2249,N_2342);
or U2755 (N_2755,N_2487,N_2029);
xnor U2756 (N_2756,N_2214,N_2100);
nand U2757 (N_2757,N_2493,N_2467);
or U2758 (N_2758,N_2042,N_2359);
and U2759 (N_2759,N_2100,N_2422);
nor U2760 (N_2760,N_2133,N_2055);
and U2761 (N_2761,N_2104,N_2357);
nand U2762 (N_2762,N_2488,N_2007);
nor U2763 (N_2763,N_2029,N_2270);
and U2764 (N_2764,N_2351,N_2105);
xor U2765 (N_2765,N_2215,N_2172);
nor U2766 (N_2766,N_2079,N_2156);
and U2767 (N_2767,N_2077,N_2198);
or U2768 (N_2768,N_2234,N_2249);
or U2769 (N_2769,N_2168,N_2273);
and U2770 (N_2770,N_2281,N_2277);
and U2771 (N_2771,N_2029,N_2122);
or U2772 (N_2772,N_2038,N_2209);
xor U2773 (N_2773,N_2290,N_2363);
nand U2774 (N_2774,N_2415,N_2323);
xor U2775 (N_2775,N_2423,N_2147);
and U2776 (N_2776,N_2352,N_2260);
and U2777 (N_2777,N_2292,N_2111);
xor U2778 (N_2778,N_2152,N_2146);
or U2779 (N_2779,N_2378,N_2295);
and U2780 (N_2780,N_2119,N_2344);
xnor U2781 (N_2781,N_2164,N_2109);
xor U2782 (N_2782,N_2149,N_2315);
nor U2783 (N_2783,N_2042,N_2040);
nand U2784 (N_2784,N_2388,N_2179);
xnor U2785 (N_2785,N_2238,N_2452);
or U2786 (N_2786,N_2417,N_2482);
nor U2787 (N_2787,N_2258,N_2115);
or U2788 (N_2788,N_2152,N_2489);
or U2789 (N_2789,N_2010,N_2258);
or U2790 (N_2790,N_2050,N_2210);
xor U2791 (N_2791,N_2309,N_2059);
or U2792 (N_2792,N_2487,N_2363);
xnor U2793 (N_2793,N_2390,N_2441);
nand U2794 (N_2794,N_2420,N_2446);
nand U2795 (N_2795,N_2494,N_2106);
nor U2796 (N_2796,N_2158,N_2412);
and U2797 (N_2797,N_2079,N_2118);
xnor U2798 (N_2798,N_2481,N_2002);
or U2799 (N_2799,N_2354,N_2491);
xnor U2800 (N_2800,N_2214,N_2242);
or U2801 (N_2801,N_2462,N_2448);
nor U2802 (N_2802,N_2410,N_2014);
xor U2803 (N_2803,N_2047,N_2328);
and U2804 (N_2804,N_2130,N_2292);
xnor U2805 (N_2805,N_2017,N_2164);
xnor U2806 (N_2806,N_2100,N_2239);
nand U2807 (N_2807,N_2095,N_2289);
nor U2808 (N_2808,N_2000,N_2195);
nor U2809 (N_2809,N_2401,N_2499);
xnor U2810 (N_2810,N_2445,N_2186);
nor U2811 (N_2811,N_2069,N_2027);
xnor U2812 (N_2812,N_2492,N_2417);
or U2813 (N_2813,N_2406,N_2334);
nor U2814 (N_2814,N_2011,N_2332);
nor U2815 (N_2815,N_2174,N_2373);
nand U2816 (N_2816,N_2294,N_2005);
nor U2817 (N_2817,N_2348,N_2411);
or U2818 (N_2818,N_2169,N_2390);
xnor U2819 (N_2819,N_2059,N_2238);
or U2820 (N_2820,N_2042,N_2392);
nor U2821 (N_2821,N_2292,N_2092);
xor U2822 (N_2822,N_2053,N_2453);
nand U2823 (N_2823,N_2343,N_2195);
or U2824 (N_2824,N_2136,N_2062);
or U2825 (N_2825,N_2354,N_2278);
nor U2826 (N_2826,N_2495,N_2288);
or U2827 (N_2827,N_2198,N_2333);
and U2828 (N_2828,N_2467,N_2209);
xor U2829 (N_2829,N_2297,N_2403);
xnor U2830 (N_2830,N_2204,N_2292);
xnor U2831 (N_2831,N_2067,N_2287);
nand U2832 (N_2832,N_2027,N_2348);
and U2833 (N_2833,N_2002,N_2252);
and U2834 (N_2834,N_2494,N_2050);
xnor U2835 (N_2835,N_2450,N_2391);
nor U2836 (N_2836,N_2499,N_2309);
nor U2837 (N_2837,N_2481,N_2137);
or U2838 (N_2838,N_2126,N_2006);
or U2839 (N_2839,N_2176,N_2459);
nor U2840 (N_2840,N_2171,N_2106);
nor U2841 (N_2841,N_2497,N_2011);
and U2842 (N_2842,N_2243,N_2177);
xor U2843 (N_2843,N_2350,N_2314);
xnor U2844 (N_2844,N_2364,N_2220);
nand U2845 (N_2845,N_2237,N_2090);
and U2846 (N_2846,N_2148,N_2305);
xnor U2847 (N_2847,N_2021,N_2089);
and U2848 (N_2848,N_2462,N_2312);
xor U2849 (N_2849,N_2355,N_2206);
nand U2850 (N_2850,N_2402,N_2231);
nor U2851 (N_2851,N_2157,N_2161);
nand U2852 (N_2852,N_2402,N_2252);
nor U2853 (N_2853,N_2120,N_2395);
xor U2854 (N_2854,N_2439,N_2246);
xor U2855 (N_2855,N_2024,N_2049);
and U2856 (N_2856,N_2116,N_2079);
and U2857 (N_2857,N_2173,N_2061);
or U2858 (N_2858,N_2443,N_2418);
nor U2859 (N_2859,N_2034,N_2120);
or U2860 (N_2860,N_2263,N_2016);
xnor U2861 (N_2861,N_2001,N_2350);
nand U2862 (N_2862,N_2439,N_2467);
and U2863 (N_2863,N_2400,N_2029);
or U2864 (N_2864,N_2053,N_2449);
and U2865 (N_2865,N_2257,N_2329);
nor U2866 (N_2866,N_2135,N_2419);
nand U2867 (N_2867,N_2406,N_2104);
nor U2868 (N_2868,N_2380,N_2433);
xor U2869 (N_2869,N_2053,N_2417);
nor U2870 (N_2870,N_2257,N_2321);
nand U2871 (N_2871,N_2031,N_2045);
nor U2872 (N_2872,N_2370,N_2233);
or U2873 (N_2873,N_2202,N_2131);
nand U2874 (N_2874,N_2235,N_2142);
nor U2875 (N_2875,N_2318,N_2066);
and U2876 (N_2876,N_2159,N_2092);
nand U2877 (N_2877,N_2432,N_2493);
and U2878 (N_2878,N_2415,N_2302);
nor U2879 (N_2879,N_2246,N_2407);
nor U2880 (N_2880,N_2079,N_2251);
nand U2881 (N_2881,N_2369,N_2273);
or U2882 (N_2882,N_2322,N_2158);
or U2883 (N_2883,N_2051,N_2002);
nor U2884 (N_2884,N_2136,N_2468);
xor U2885 (N_2885,N_2261,N_2219);
xor U2886 (N_2886,N_2267,N_2372);
or U2887 (N_2887,N_2156,N_2306);
nand U2888 (N_2888,N_2202,N_2072);
nor U2889 (N_2889,N_2223,N_2390);
or U2890 (N_2890,N_2201,N_2098);
and U2891 (N_2891,N_2030,N_2120);
and U2892 (N_2892,N_2376,N_2235);
and U2893 (N_2893,N_2282,N_2492);
nor U2894 (N_2894,N_2185,N_2314);
nor U2895 (N_2895,N_2359,N_2432);
nand U2896 (N_2896,N_2106,N_2242);
nand U2897 (N_2897,N_2261,N_2107);
nand U2898 (N_2898,N_2118,N_2456);
xor U2899 (N_2899,N_2264,N_2128);
or U2900 (N_2900,N_2385,N_2137);
xnor U2901 (N_2901,N_2093,N_2194);
xor U2902 (N_2902,N_2148,N_2452);
nor U2903 (N_2903,N_2455,N_2057);
xnor U2904 (N_2904,N_2052,N_2176);
or U2905 (N_2905,N_2353,N_2247);
nand U2906 (N_2906,N_2034,N_2307);
or U2907 (N_2907,N_2453,N_2089);
and U2908 (N_2908,N_2440,N_2022);
or U2909 (N_2909,N_2051,N_2346);
and U2910 (N_2910,N_2167,N_2476);
xnor U2911 (N_2911,N_2295,N_2413);
or U2912 (N_2912,N_2214,N_2422);
nor U2913 (N_2913,N_2491,N_2289);
xnor U2914 (N_2914,N_2136,N_2112);
or U2915 (N_2915,N_2051,N_2153);
xnor U2916 (N_2916,N_2361,N_2262);
and U2917 (N_2917,N_2303,N_2291);
or U2918 (N_2918,N_2175,N_2310);
and U2919 (N_2919,N_2263,N_2383);
and U2920 (N_2920,N_2398,N_2416);
xnor U2921 (N_2921,N_2107,N_2455);
xnor U2922 (N_2922,N_2100,N_2366);
nor U2923 (N_2923,N_2450,N_2170);
xor U2924 (N_2924,N_2228,N_2408);
nor U2925 (N_2925,N_2329,N_2008);
and U2926 (N_2926,N_2436,N_2281);
or U2927 (N_2927,N_2307,N_2270);
xnor U2928 (N_2928,N_2038,N_2425);
or U2929 (N_2929,N_2456,N_2469);
nor U2930 (N_2930,N_2000,N_2449);
xor U2931 (N_2931,N_2317,N_2231);
nand U2932 (N_2932,N_2307,N_2470);
nor U2933 (N_2933,N_2086,N_2215);
xnor U2934 (N_2934,N_2245,N_2024);
nor U2935 (N_2935,N_2128,N_2416);
and U2936 (N_2936,N_2426,N_2014);
nand U2937 (N_2937,N_2156,N_2119);
and U2938 (N_2938,N_2203,N_2218);
nor U2939 (N_2939,N_2338,N_2195);
and U2940 (N_2940,N_2443,N_2332);
or U2941 (N_2941,N_2163,N_2384);
nand U2942 (N_2942,N_2042,N_2407);
nor U2943 (N_2943,N_2077,N_2264);
or U2944 (N_2944,N_2055,N_2152);
nand U2945 (N_2945,N_2021,N_2483);
xor U2946 (N_2946,N_2414,N_2168);
or U2947 (N_2947,N_2025,N_2348);
xnor U2948 (N_2948,N_2410,N_2381);
nor U2949 (N_2949,N_2149,N_2059);
xor U2950 (N_2950,N_2161,N_2217);
or U2951 (N_2951,N_2447,N_2384);
nor U2952 (N_2952,N_2423,N_2394);
or U2953 (N_2953,N_2102,N_2498);
and U2954 (N_2954,N_2326,N_2237);
xnor U2955 (N_2955,N_2301,N_2107);
xnor U2956 (N_2956,N_2201,N_2360);
xor U2957 (N_2957,N_2492,N_2132);
nand U2958 (N_2958,N_2221,N_2461);
nor U2959 (N_2959,N_2011,N_2458);
nand U2960 (N_2960,N_2323,N_2247);
or U2961 (N_2961,N_2415,N_2066);
or U2962 (N_2962,N_2179,N_2123);
nand U2963 (N_2963,N_2085,N_2357);
and U2964 (N_2964,N_2040,N_2153);
xnor U2965 (N_2965,N_2069,N_2137);
or U2966 (N_2966,N_2454,N_2289);
xor U2967 (N_2967,N_2340,N_2423);
and U2968 (N_2968,N_2474,N_2438);
and U2969 (N_2969,N_2095,N_2313);
and U2970 (N_2970,N_2095,N_2263);
xor U2971 (N_2971,N_2484,N_2470);
or U2972 (N_2972,N_2091,N_2464);
nand U2973 (N_2973,N_2471,N_2069);
or U2974 (N_2974,N_2272,N_2454);
xor U2975 (N_2975,N_2197,N_2317);
nand U2976 (N_2976,N_2045,N_2120);
xor U2977 (N_2977,N_2114,N_2156);
nand U2978 (N_2978,N_2139,N_2389);
xor U2979 (N_2979,N_2342,N_2086);
nand U2980 (N_2980,N_2448,N_2013);
xnor U2981 (N_2981,N_2349,N_2351);
nand U2982 (N_2982,N_2350,N_2421);
xnor U2983 (N_2983,N_2200,N_2382);
nand U2984 (N_2984,N_2252,N_2262);
and U2985 (N_2985,N_2300,N_2414);
or U2986 (N_2986,N_2360,N_2210);
nand U2987 (N_2987,N_2333,N_2125);
nand U2988 (N_2988,N_2149,N_2293);
nand U2989 (N_2989,N_2416,N_2062);
nor U2990 (N_2990,N_2116,N_2432);
or U2991 (N_2991,N_2452,N_2335);
xor U2992 (N_2992,N_2227,N_2472);
or U2993 (N_2993,N_2246,N_2299);
nor U2994 (N_2994,N_2470,N_2456);
xor U2995 (N_2995,N_2340,N_2285);
and U2996 (N_2996,N_2145,N_2371);
nor U2997 (N_2997,N_2049,N_2354);
xnor U2998 (N_2998,N_2421,N_2162);
and U2999 (N_2999,N_2423,N_2411);
xor U3000 (N_3000,N_2858,N_2522);
nor U3001 (N_3001,N_2826,N_2805);
nand U3002 (N_3002,N_2927,N_2770);
or U3003 (N_3003,N_2725,N_2845);
nor U3004 (N_3004,N_2658,N_2681);
nand U3005 (N_3005,N_2780,N_2769);
and U3006 (N_3006,N_2582,N_2850);
or U3007 (N_3007,N_2961,N_2797);
and U3008 (N_3008,N_2650,N_2536);
and U3009 (N_3009,N_2840,N_2617);
nand U3010 (N_3010,N_2559,N_2603);
nand U3011 (N_3011,N_2854,N_2706);
xnor U3012 (N_3012,N_2970,N_2788);
nand U3013 (N_3013,N_2527,N_2873);
xor U3014 (N_3014,N_2995,N_2879);
xnor U3015 (N_3015,N_2763,N_2510);
nor U3016 (N_3016,N_2885,N_2920);
xnor U3017 (N_3017,N_2673,N_2701);
nand U3018 (N_3018,N_2570,N_2669);
nand U3019 (N_3019,N_2657,N_2550);
and U3020 (N_3020,N_2734,N_2985);
nor U3021 (N_3021,N_2859,N_2781);
nand U3022 (N_3022,N_2990,N_2719);
nor U3023 (N_3023,N_2878,N_2910);
xnor U3024 (N_3024,N_2965,N_2688);
and U3025 (N_3025,N_2670,N_2933);
or U3026 (N_3026,N_2899,N_2543);
xnor U3027 (N_3027,N_2590,N_2634);
nand U3028 (N_3028,N_2684,N_2857);
xor U3029 (N_3029,N_2666,N_2690);
nor U3030 (N_3030,N_2622,N_2908);
nand U3031 (N_3031,N_2856,N_2555);
nand U3032 (N_3032,N_2735,N_2904);
nor U3033 (N_3033,N_2612,N_2976);
nand U3034 (N_3034,N_2632,N_2938);
and U3035 (N_3035,N_2546,N_2714);
xnor U3036 (N_3036,N_2647,N_2786);
xnor U3037 (N_3037,N_2761,N_2676);
nor U3038 (N_3038,N_2790,N_2838);
and U3039 (N_3039,N_2989,N_2697);
and U3040 (N_3040,N_2515,N_2872);
nor U3041 (N_3041,N_2951,N_2796);
xor U3042 (N_3042,N_2942,N_2604);
or U3043 (N_3043,N_2553,N_2560);
and U3044 (N_3044,N_2554,N_2695);
and U3045 (N_3045,N_2984,N_2762);
or U3046 (N_3046,N_2668,N_2837);
xor U3047 (N_3047,N_2831,N_2649);
nand U3048 (N_3048,N_2778,N_2909);
nor U3049 (N_3049,N_2549,N_2860);
or U3050 (N_3050,N_2548,N_2758);
nand U3051 (N_3051,N_2694,N_2947);
nor U3052 (N_3052,N_2664,N_2918);
nor U3053 (N_3053,N_2744,N_2700);
nand U3054 (N_3054,N_2902,N_2924);
and U3055 (N_3055,N_2974,N_2847);
xor U3056 (N_3056,N_2577,N_2644);
and U3057 (N_3057,N_2584,N_2538);
or U3058 (N_3058,N_2834,N_2730);
nor U3059 (N_3059,N_2643,N_2846);
and U3060 (N_3060,N_2573,N_2642);
and U3061 (N_3061,N_2640,N_2791);
or U3062 (N_3062,N_2898,N_2978);
nand U3063 (N_3063,N_2988,N_2880);
and U3064 (N_3064,N_2993,N_2547);
or U3065 (N_3065,N_2811,N_2637);
nand U3066 (N_3066,N_2614,N_2591);
xor U3067 (N_3067,N_2520,N_2896);
xnor U3068 (N_3068,N_2599,N_2506);
and U3069 (N_3069,N_2660,N_2819);
nor U3070 (N_3070,N_2756,N_2720);
and U3071 (N_3071,N_2930,N_2530);
or U3072 (N_3072,N_2956,N_2539);
nor U3073 (N_3073,N_2906,N_2566);
or U3074 (N_3074,N_2563,N_2957);
or U3075 (N_3075,N_2708,N_2944);
or U3076 (N_3076,N_2602,N_2994);
or U3077 (N_3077,N_2803,N_2870);
or U3078 (N_3078,N_2979,N_2749);
nand U3079 (N_3079,N_2516,N_2844);
or U3080 (N_3080,N_2864,N_2512);
nor U3081 (N_3081,N_2972,N_2691);
nor U3082 (N_3082,N_2799,N_2958);
nor U3083 (N_3083,N_2661,N_2656);
nand U3084 (N_3084,N_2542,N_2912);
nand U3085 (N_3085,N_2954,N_2812);
nand U3086 (N_3086,N_2501,N_2508);
xor U3087 (N_3087,N_2534,N_2528);
nor U3088 (N_3088,N_2897,N_2894);
xnor U3089 (N_3089,N_2800,N_2905);
nor U3090 (N_3090,N_2816,N_2729);
or U3091 (N_3091,N_2948,N_2773);
and U3092 (N_3092,N_2741,N_2615);
or U3093 (N_3093,N_2783,N_2699);
nor U3094 (N_3094,N_2784,N_2757);
nand U3095 (N_3095,N_2986,N_2609);
and U3096 (N_3096,N_2710,N_2728);
nor U3097 (N_3097,N_2541,N_2765);
or U3098 (N_3098,N_2675,N_2771);
nand U3099 (N_3099,N_2925,N_2500);
nand U3100 (N_3100,N_2960,N_2991);
or U3101 (N_3101,N_2628,N_2895);
or U3102 (N_3102,N_2815,N_2524);
nor U3103 (N_3103,N_2809,N_2638);
nand U3104 (N_3104,N_2853,N_2975);
xor U3105 (N_3105,N_2705,N_2968);
and U3106 (N_3106,N_2513,N_2716);
nor U3107 (N_3107,N_2843,N_2750);
or U3108 (N_3108,N_2674,N_2959);
nand U3109 (N_3109,N_2597,N_2552);
xnor U3110 (N_3110,N_2693,N_2667);
nor U3111 (N_3111,N_2869,N_2672);
or U3112 (N_3112,N_2682,N_2955);
nor U3113 (N_3113,N_2997,N_2832);
nand U3114 (N_3114,N_2569,N_2608);
nand U3115 (N_3115,N_2813,N_2683);
nor U3116 (N_3116,N_2935,N_2767);
xor U3117 (N_3117,N_2718,N_2868);
nor U3118 (N_3118,N_2629,N_2753);
and U3119 (N_3119,N_2601,N_2889);
or U3120 (N_3120,N_2561,N_2564);
or U3121 (N_3121,N_2631,N_2915);
nand U3122 (N_3122,N_2523,N_2923);
xor U3123 (N_3123,N_2653,N_2882);
nand U3124 (N_3124,N_2579,N_2619);
xor U3125 (N_3125,N_2545,N_2852);
or U3126 (N_3126,N_2928,N_2588);
nand U3127 (N_3127,N_2849,N_2806);
xnor U3128 (N_3128,N_2759,N_2651);
and U3129 (N_3129,N_2967,N_2863);
nor U3130 (N_3130,N_2807,N_2817);
nor U3131 (N_3131,N_2711,N_2887);
nand U3132 (N_3132,N_2941,N_2848);
nand U3133 (N_3133,N_2698,N_2921);
xnor U3134 (N_3134,N_2940,N_2823);
or U3135 (N_3135,N_2821,N_2911);
nand U3136 (N_3136,N_2535,N_2917);
or U3137 (N_3137,N_2862,N_2825);
nor U3138 (N_3138,N_2521,N_2525);
nand U3139 (N_3139,N_2736,N_2829);
nand U3140 (N_3140,N_2943,N_2743);
xor U3141 (N_3141,N_2893,N_2966);
or U3142 (N_3142,N_2861,N_2739);
or U3143 (N_3143,N_2576,N_2727);
nor U3144 (N_3144,N_2685,N_2914);
and U3145 (N_3145,N_2611,N_2818);
xnor U3146 (N_3146,N_2594,N_2916);
xor U3147 (N_3147,N_2686,N_2953);
xnor U3148 (N_3148,N_2931,N_2999);
nand U3149 (N_3149,N_2625,N_2575);
nand U3150 (N_3150,N_2503,N_2977);
xnor U3151 (N_3151,N_2866,N_2782);
or U3152 (N_3152,N_2529,N_2574);
nand U3153 (N_3153,N_2883,N_2751);
nand U3154 (N_3154,N_2822,N_2937);
nor U3155 (N_3155,N_2874,N_2963);
or U3156 (N_3156,N_2738,N_2648);
nand U3157 (N_3157,N_2600,N_2903);
and U3158 (N_3158,N_2692,N_2892);
xnor U3159 (N_3159,N_2726,N_2772);
nand U3160 (N_3160,N_2867,N_2624);
xnor U3161 (N_3161,N_2774,N_2777);
and U3162 (N_3162,N_2830,N_2981);
xor U3163 (N_3163,N_2680,N_2626);
or U3164 (N_3164,N_2721,N_2572);
or U3165 (N_3165,N_2881,N_2715);
or U3166 (N_3166,N_2665,N_2540);
xor U3167 (N_3167,N_2630,N_2531);
nor U3168 (N_3168,N_2519,N_2704);
xor U3169 (N_3169,N_2936,N_2639);
and U3170 (N_3170,N_2724,N_2747);
nor U3171 (N_3171,N_2980,N_2679);
or U3172 (N_3172,N_2973,N_2802);
xnor U3173 (N_3173,N_2571,N_2587);
nor U3174 (N_3174,N_2969,N_2713);
xnor U3175 (N_3175,N_2616,N_2623);
nand U3176 (N_3176,N_2851,N_2787);
or U3177 (N_3177,N_2717,N_2946);
or U3178 (N_3178,N_2659,N_2745);
nor U3179 (N_3179,N_2998,N_2703);
nand U3180 (N_3180,N_2755,N_2907);
nand U3181 (N_3181,N_2952,N_2775);
or U3182 (N_3182,N_2792,N_2776);
or U3183 (N_3183,N_2833,N_2919);
nand U3184 (N_3184,N_2645,N_2886);
xnor U3185 (N_3185,N_2733,N_2610);
xnor U3186 (N_3186,N_2779,N_2824);
nor U3187 (N_3187,N_2511,N_2865);
and U3188 (N_3188,N_2641,N_2592);
nand U3189 (N_3189,N_2731,N_2732);
xor U3190 (N_3190,N_2502,N_2996);
nor U3191 (N_3191,N_2633,N_2804);
nor U3192 (N_3192,N_2752,N_2890);
and U3193 (N_3193,N_2593,N_2607);
xor U3194 (N_3194,N_2652,N_2504);
and U3195 (N_3195,N_2537,N_2696);
nor U3196 (N_3196,N_2557,N_2526);
or U3197 (N_3197,N_2983,N_2891);
nor U3198 (N_3198,N_2841,N_2971);
nor U3199 (N_3199,N_2509,N_2962);
nand U3200 (N_3200,N_2583,N_2835);
or U3201 (N_3201,N_2926,N_2627);
and U3202 (N_3202,N_2798,N_2635);
nor U3203 (N_3203,N_2514,N_2934);
nor U3204 (N_3204,N_2875,N_2544);
or U3205 (N_3205,N_2598,N_2689);
nand U3206 (N_3206,N_2662,N_2949);
or U3207 (N_3207,N_2518,N_2808);
or U3208 (N_3208,N_2589,N_2562);
and U3209 (N_3209,N_2795,N_2746);
nand U3210 (N_3210,N_2654,N_2888);
nor U3211 (N_3211,N_2663,N_2606);
xnor U3212 (N_3212,N_2922,N_2793);
and U3213 (N_3213,N_2842,N_2855);
nand U3214 (N_3214,N_2581,N_2655);
xnor U3215 (N_3215,N_2722,N_2742);
xnor U3216 (N_3216,N_2964,N_2586);
xnor U3217 (N_3217,N_2801,N_2982);
and U3218 (N_3218,N_2621,N_2754);
nor U3219 (N_3219,N_2687,N_2618);
or U3220 (N_3220,N_2556,N_2507);
nand U3221 (N_3221,N_2595,N_2871);
xnor U3222 (N_3222,N_2620,N_2877);
nand U3223 (N_3223,N_2900,N_2737);
and U3224 (N_3224,N_2764,N_2533);
xor U3225 (N_3225,N_2768,N_2876);
xnor U3226 (N_3226,N_2677,N_2884);
and U3227 (N_3227,N_2810,N_2596);
or U3228 (N_3228,N_2712,N_2517);
and U3229 (N_3229,N_2568,N_2814);
nand U3230 (N_3230,N_2794,N_2702);
nor U3231 (N_3231,N_2578,N_2740);
and U3232 (N_3232,N_2567,N_2839);
or U3233 (N_3233,N_2558,N_2913);
and U3234 (N_3234,N_2565,N_2785);
xor U3235 (N_3235,N_2932,N_2992);
nand U3236 (N_3236,N_2636,N_2950);
or U3237 (N_3237,N_2532,N_2827);
nand U3238 (N_3238,N_2709,N_2580);
xor U3239 (N_3239,N_2987,N_2585);
and U3240 (N_3240,N_2723,N_2551);
nor U3241 (N_3241,N_2945,N_2929);
or U3242 (N_3242,N_2671,N_2678);
or U3243 (N_3243,N_2505,N_2828);
nor U3244 (N_3244,N_2707,N_2901);
nor U3245 (N_3245,N_2646,N_2820);
nand U3246 (N_3246,N_2766,N_2789);
and U3247 (N_3247,N_2760,N_2605);
nor U3248 (N_3248,N_2939,N_2748);
nor U3249 (N_3249,N_2613,N_2836);
nand U3250 (N_3250,N_2562,N_2938);
xnor U3251 (N_3251,N_2578,N_2546);
and U3252 (N_3252,N_2675,N_2612);
or U3253 (N_3253,N_2995,N_2559);
nor U3254 (N_3254,N_2832,N_2887);
xnor U3255 (N_3255,N_2707,N_2670);
and U3256 (N_3256,N_2891,N_2913);
nor U3257 (N_3257,N_2665,N_2646);
or U3258 (N_3258,N_2696,N_2576);
nor U3259 (N_3259,N_2538,N_2753);
and U3260 (N_3260,N_2981,N_2810);
nand U3261 (N_3261,N_2879,N_2559);
nand U3262 (N_3262,N_2693,N_2908);
and U3263 (N_3263,N_2505,N_2831);
nand U3264 (N_3264,N_2514,N_2563);
xor U3265 (N_3265,N_2759,N_2850);
xnor U3266 (N_3266,N_2501,N_2830);
xor U3267 (N_3267,N_2513,N_2507);
or U3268 (N_3268,N_2528,N_2529);
and U3269 (N_3269,N_2502,N_2853);
xor U3270 (N_3270,N_2747,N_2581);
or U3271 (N_3271,N_2870,N_2778);
or U3272 (N_3272,N_2853,N_2892);
and U3273 (N_3273,N_2584,N_2596);
or U3274 (N_3274,N_2746,N_2554);
xor U3275 (N_3275,N_2536,N_2852);
nor U3276 (N_3276,N_2829,N_2817);
nand U3277 (N_3277,N_2946,N_2703);
nor U3278 (N_3278,N_2936,N_2632);
or U3279 (N_3279,N_2502,N_2523);
and U3280 (N_3280,N_2650,N_2867);
and U3281 (N_3281,N_2752,N_2560);
and U3282 (N_3282,N_2544,N_2537);
nand U3283 (N_3283,N_2717,N_2981);
xnor U3284 (N_3284,N_2591,N_2850);
and U3285 (N_3285,N_2607,N_2969);
nor U3286 (N_3286,N_2732,N_2937);
xnor U3287 (N_3287,N_2930,N_2535);
or U3288 (N_3288,N_2519,N_2741);
and U3289 (N_3289,N_2507,N_2720);
and U3290 (N_3290,N_2900,N_2634);
and U3291 (N_3291,N_2518,N_2528);
nand U3292 (N_3292,N_2697,N_2592);
and U3293 (N_3293,N_2573,N_2703);
nor U3294 (N_3294,N_2948,N_2822);
xnor U3295 (N_3295,N_2559,N_2859);
xor U3296 (N_3296,N_2877,N_2652);
nor U3297 (N_3297,N_2699,N_2859);
nor U3298 (N_3298,N_2848,N_2707);
xnor U3299 (N_3299,N_2810,N_2663);
nand U3300 (N_3300,N_2615,N_2924);
nand U3301 (N_3301,N_2955,N_2661);
or U3302 (N_3302,N_2800,N_2615);
xnor U3303 (N_3303,N_2922,N_2693);
nand U3304 (N_3304,N_2819,N_2543);
or U3305 (N_3305,N_2572,N_2577);
and U3306 (N_3306,N_2645,N_2630);
nand U3307 (N_3307,N_2629,N_2502);
xnor U3308 (N_3308,N_2560,N_2985);
nor U3309 (N_3309,N_2885,N_2776);
and U3310 (N_3310,N_2928,N_2976);
nand U3311 (N_3311,N_2657,N_2759);
nor U3312 (N_3312,N_2737,N_2993);
and U3313 (N_3313,N_2929,N_2916);
nor U3314 (N_3314,N_2977,N_2955);
or U3315 (N_3315,N_2982,N_2996);
xnor U3316 (N_3316,N_2558,N_2928);
or U3317 (N_3317,N_2689,N_2596);
and U3318 (N_3318,N_2901,N_2851);
xor U3319 (N_3319,N_2702,N_2946);
nor U3320 (N_3320,N_2811,N_2721);
and U3321 (N_3321,N_2727,N_2510);
or U3322 (N_3322,N_2946,N_2794);
nand U3323 (N_3323,N_2863,N_2853);
nand U3324 (N_3324,N_2634,N_2678);
xor U3325 (N_3325,N_2689,N_2587);
or U3326 (N_3326,N_2568,N_2734);
or U3327 (N_3327,N_2932,N_2981);
or U3328 (N_3328,N_2790,N_2694);
nor U3329 (N_3329,N_2545,N_2700);
nor U3330 (N_3330,N_2671,N_2595);
and U3331 (N_3331,N_2735,N_2758);
xor U3332 (N_3332,N_2939,N_2535);
or U3333 (N_3333,N_2516,N_2876);
nand U3334 (N_3334,N_2590,N_2870);
xor U3335 (N_3335,N_2812,N_2588);
nand U3336 (N_3336,N_2912,N_2966);
or U3337 (N_3337,N_2964,N_2532);
or U3338 (N_3338,N_2511,N_2811);
and U3339 (N_3339,N_2706,N_2670);
nor U3340 (N_3340,N_2562,N_2984);
nor U3341 (N_3341,N_2971,N_2544);
nor U3342 (N_3342,N_2838,N_2658);
or U3343 (N_3343,N_2906,N_2589);
nand U3344 (N_3344,N_2855,N_2749);
xor U3345 (N_3345,N_2775,N_2947);
xnor U3346 (N_3346,N_2658,N_2908);
and U3347 (N_3347,N_2789,N_2525);
and U3348 (N_3348,N_2783,N_2649);
nand U3349 (N_3349,N_2693,N_2830);
xor U3350 (N_3350,N_2703,N_2770);
nor U3351 (N_3351,N_2877,N_2883);
xor U3352 (N_3352,N_2874,N_2616);
or U3353 (N_3353,N_2980,N_2997);
or U3354 (N_3354,N_2527,N_2682);
or U3355 (N_3355,N_2574,N_2734);
nor U3356 (N_3356,N_2678,N_2977);
and U3357 (N_3357,N_2818,N_2991);
nor U3358 (N_3358,N_2548,N_2875);
or U3359 (N_3359,N_2708,N_2500);
or U3360 (N_3360,N_2596,N_2528);
nor U3361 (N_3361,N_2899,N_2549);
or U3362 (N_3362,N_2594,N_2884);
xor U3363 (N_3363,N_2961,N_2823);
and U3364 (N_3364,N_2821,N_2959);
nor U3365 (N_3365,N_2942,N_2997);
and U3366 (N_3366,N_2519,N_2928);
nand U3367 (N_3367,N_2992,N_2757);
nor U3368 (N_3368,N_2684,N_2527);
and U3369 (N_3369,N_2744,N_2995);
nand U3370 (N_3370,N_2561,N_2724);
xnor U3371 (N_3371,N_2946,N_2983);
nor U3372 (N_3372,N_2845,N_2727);
and U3373 (N_3373,N_2665,N_2609);
nor U3374 (N_3374,N_2678,N_2826);
and U3375 (N_3375,N_2826,N_2648);
nor U3376 (N_3376,N_2715,N_2836);
and U3377 (N_3377,N_2678,N_2643);
and U3378 (N_3378,N_2925,N_2614);
nand U3379 (N_3379,N_2775,N_2725);
xnor U3380 (N_3380,N_2837,N_2933);
nor U3381 (N_3381,N_2692,N_2846);
or U3382 (N_3382,N_2838,N_2680);
and U3383 (N_3383,N_2843,N_2945);
nand U3384 (N_3384,N_2700,N_2725);
nand U3385 (N_3385,N_2909,N_2762);
xor U3386 (N_3386,N_2531,N_2788);
xnor U3387 (N_3387,N_2625,N_2801);
or U3388 (N_3388,N_2906,N_2812);
nand U3389 (N_3389,N_2659,N_2970);
or U3390 (N_3390,N_2865,N_2796);
or U3391 (N_3391,N_2892,N_2902);
nor U3392 (N_3392,N_2912,N_2755);
nand U3393 (N_3393,N_2933,N_2920);
and U3394 (N_3394,N_2566,N_2640);
and U3395 (N_3395,N_2514,N_2710);
or U3396 (N_3396,N_2603,N_2815);
nor U3397 (N_3397,N_2800,N_2570);
nand U3398 (N_3398,N_2927,N_2537);
xnor U3399 (N_3399,N_2579,N_2544);
and U3400 (N_3400,N_2912,N_2972);
or U3401 (N_3401,N_2923,N_2665);
xnor U3402 (N_3402,N_2909,N_2788);
nor U3403 (N_3403,N_2828,N_2950);
nand U3404 (N_3404,N_2603,N_2948);
or U3405 (N_3405,N_2651,N_2815);
nor U3406 (N_3406,N_2671,N_2941);
or U3407 (N_3407,N_2838,N_2716);
or U3408 (N_3408,N_2680,N_2757);
or U3409 (N_3409,N_2937,N_2870);
nor U3410 (N_3410,N_2580,N_2579);
xor U3411 (N_3411,N_2528,N_2778);
or U3412 (N_3412,N_2838,N_2778);
or U3413 (N_3413,N_2677,N_2909);
and U3414 (N_3414,N_2570,N_2563);
nand U3415 (N_3415,N_2965,N_2881);
nor U3416 (N_3416,N_2958,N_2529);
xor U3417 (N_3417,N_2601,N_2521);
or U3418 (N_3418,N_2916,N_2528);
xor U3419 (N_3419,N_2627,N_2934);
and U3420 (N_3420,N_2756,N_2551);
xnor U3421 (N_3421,N_2928,N_2912);
xnor U3422 (N_3422,N_2525,N_2540);
nor U3423 (N_3423,N_2939,N_2785);
and U3424 (N_3424,N_2759,N_2637);
nor U3425 (N_3425,N_2623,N_2524);
nand U3426 (N_3426,N_2874,N_2634);
xnor U3427 (N_3427,N_2937,N_2611);
nor U3428 (N_3428,N_2963,N_2641);
xnor U3429 (N_3429,N_2991,N_2663);
xnor U3430 (N_3430,N_2672,N_2596);
nor U3431 (N_3431,N_2750,N_2839);
or U3432 (N_3432,N_2843,N_2508);
nor U3433 (N_3433,N_2558,N_2580);
or U3434 (N_3434,N_2819,N_2700);
or U3435 (N_3435,N_2993,N_2985);
and U3436 (N_3436,N_2626,N_2797);
nand U3437 (N_3437,N_2949,N_2960);
and U3438 (N_3438,N_2586,N_2703);
and U3439 (N_3439,N_2680,N_2910);
xnor U3440 (N_3440,N_2979,N_2818);
or U3441 (N_3441,N_2651,N_2690);
xor U3442 (N_3442,N_2678,N_2648);
nand U3443 (N_3443,N_2656,N_2864);
and U3444 (N_3444,N_2916,N_2836);
and U3445 (N_3445,N_2935,N_2558);
and U3446 (N_3446,N_2668,N_2829);
or U3447 (N_3447,N_2562,N_2732);
or U3448 (N_3448,N_2505,N_2575);
xor U3449 (N_3449,N_2594,N_2740);
nand U3450 (N_3450,N_2975,N_2990);
or U3451 (N_3451,N_2912,N_2949);
nand U3452 (N_3452,N_2722,N_2633);
nor U3453 (N_3453,N_2618,N_2519);
nor U3454 (N_3454,N_2566,N_2759);
or U3455 (N_3455,N_2967,N_2911);
xor U3456 (N_3456,N_2524,N_2798);
nor U3457 (N_3457,N_2589,N_2930);
nor U3458 (N_3458,N_2638,N_2532);
or U3459 (N_3459,N_2552,N_2717);
or U3460 (N_3460,N_2663,N_2660);
xor U3461 (N_3461,N_2611,N_2942);
nand U3462 (N_3462,N_2874,N_2905);
or U3463 (N_3463,N_2967,N_2702);
or U3464 (N_3464,N_2995,N_2500);
and U3465 (N_3465,N_2755,N_2674);
and U3466 (N_3466,N_2921,N_2858);
nor U3467 (N_3467,N_2539,N_2523);
or U3468 (N_3468,N_2791,N_2910);
nor U3469 (N_3469,N_2806,N_2958);
xnor U3470 (N_3470,N_2543,N_2752);
xnor U3471 (N_3471,N_2730,N_2755);
nor U3472 (N_3472,N_2550,N_2931);
or U3473 (N_3473,N_2849,N_2770);
nand U3474 (N_3474,N_2577,N_2595);
and U3475 (N_3475,N_2524,N_2778);
nand U3476 (N_3476,N_2831,N_2548);
xor U3477 (N_3477,N_2607,N_2861);
xor U3478 (N_3478,N_2536,N_2990);
nor U3479 (N_3479,N_2851,N_2560);
and U3480 (N_3480,N_2679,N_2943);
nand U3481 (N_3481,N_2768,N_2647);
xnor U3482 (N_3482,N_2640,N_2516);
or U3483 (N_3483,N_2740,N_2907);
or U3484 (N_3484,N_2514,N_2949);
or U3485 (N_3485,N_2749,N_2688);
and U3486 (N_3486,N_2619,N_2903);
and U3487 (N_3487,N_2924,N_2538);
xnor U3488 (N_3488,N_2861,N_2578);
nand U3489 (N_3489,N_2705,N_2578);
nand U3490 (N_3490,N_2651,N_2686);
or U3491 (N_3491,N_2850,N_2884);
or U3492 (N_3492,N_2642,N_2647);
nor U3493 (N_3493,N_2875,N_2961);
nor U3494 (N_3494,N_2582,N_2542);
and U3495 (N_3495,N_2603,N_2619);
nand U3496 (N_3496,N_2836,N_2565);
xnor U3497 (N_3497,N_2899,N_2735);
and U3498 (N_3498,N_2585,N_2693);
xor U3499 (N_3499,N_2714,N_2550);
xnor U3500 (N_3500,N_3020,N_3191);
xnor U3501 (N_3501,N_3226,N_3162);
or U3502 (N_3502,N_3276,N_3135);
nor U3503 (N_3503,N_3401,N_3475);
nor U3504 (N_3504,N_3242,N_3407);
and U3505 (N_3505,N_3152,N_3057);
nor U3506 (N_3506,N_3261,N_3246);
or U3507 (N_3507,N_3027,N_3255);
nand U3508 (N_3508,N_3081,N_3237);
nand U3509 (N_3509,N_3428,N_3084);
and U3510 (N_3510,N_3159,N_3447);
and U3511 (N_3511,N_3254,N_3239);
and U3512 (N_3512,N_3129,N_3157);
or U3513 (N_3513,N_3161,N_3438);
and U3514 (N_3514,N_3153,N_3422);
or U3515 (N_3515,N_3453,N_3414);
nor U3516 (N_3516,N_3105,N_3173);
or U3517 (N_3517,N_3429,N_3283);
nor U3518 (N_3518,N_3091,N_3053);
and U3519 (N_3519,N_3298,N_3096);
nand U3520 (N_3520,N_3369,N_3037);
xor U3521 (N_3521,N_3028,N_3035);
nor U3522 (N_3522,N_3209,N_3364);
xnor U3523 (N_3523,N_3275,N_3311);
nor U3524 (N_3524,N_3287,N_3183);
nor U3525 (N_3525,N_3188,N_3079);
nand U3526 (N_3526,N_3021,N_3212);
or U3527 (N_3527,N_3274,N_3430);
xor U3528 (N_3528,N_3123,N_3415);
nor U3529 (N_3529,N_3030,N_3342);
and U3530 (N_3530,N_3359,N_3221);
or U3531 (N_3531,N_3256,N_3354);
xor U3532 (N_3532,N_3385,N_3337);
nand U3533 (N_3533,N_3405,N_3263);
nor U3534 (N_3534,N_3233,N_3493);
and U3535 (N_3535,N_3076,N_3134);
and U3536 (N_3536,N_3033,N_3420);
or U3537 (N_3537,N_3379,N_3392);
and U3538 (N_3538,N_3497,N_3358);
nand U3539 (N_3539,N_3333,N_3264);
xor U3540 (N_3540,N_3106,N_3217);
and U3541 (N_3541,N_3499,N_3299);
xnor U3542 (N_3542,N_3085,N_3269);
nor U3543 (N_3543,N_3160,N_3349);
or U3544 (N_3544,N_3114,N_3381);
or U3545 (N_3545,N_3334,N_3127);
or U3546 (N_3546,N_3348,N_3278);
and U3547 (N_3547,N_3351,N_3412);
xnor U3548 (N_3548,N_3046,N_3155);
xnor U3549 (N_3549,N_3145,N_3366);
or U3550 (N_3550,N_3286,N_3456);
nand U3551 (N_3551,N_3017,N_3446);
xor U3552 (N_3552,N_3010,N_3386);
nand U3553 (N_3553,N_3198,N_3055);
or U3554 (N_3554,N_3330,N_3075);
and U3555 (N_3555,N_3262,N_3180);
or U3556 (N_3556,N_3419,N_3302);
nand U3557 (N_3557,N_3174,N_3067);
nor U3558 (N_3558,N_3095,N_3062);
xnor U3559 (N_3559,N_3203,N_3316);
and U3560 (N_3560,N_3448,N_3346);
xnor U3561 (N_3561,N_3368,N_3058);
or U3562 (N_3562,N_3408,N_3471);
xnor U3563 (N_3563,N_3063,N_3249);
or U3564 (N_3564,N_3459,N_3380);
nand U3565 (N_3565,N_3088,N_3181);
xnor U3566 (N_3566,N_3109,N_3111);
or U3567 (N_3567,N_3102,N_3393);
nor U3568 (N_3568,N_3151,N_3389);
or U3569 (N_3569,N_3252,N_3306);
or U3570 (N_3570,N_3464,N_3433);
nor U3571 (N_3571,N_3170,N_3011);
xor U3572 (N_3572,N_3418,N_3018);
and U3573 (N_3573,N_3344,N_3400);
or U3574 (N_3574,N_3003,N_3394);
nor U3575 (N_3575,N_3353,N_3116);
xnor U3576 (N_3576,N_3495,N_3189);
nand U3577 (N_3577,N_3310,N_3051);
or U3578 (N_3578,N_3352,N_3399);
nor U3579 (N_3579,N_3089,N_3373);
or U3580 (N_3580,N_3049,N_3317);
nand U3581 (N_3581,N_3194,N_3176);
nand U3582 (N_3582,N_3083,N_3402);
nand U3583 (N_3583,N_3068,N_3455);
nand U3584 (N_3584,N_3434,N_3031);
or U3585 (N_3585,N_3016,N_3466);
nand U3586 (N_3586,N_3074,N_3207);
nor U3587 (N_3587,N_3234,N_3034);
nand U3588 (N_3588,N_3013,N_3492);
nor U3589 (N_3589,N_3376,N_3069);
and U3590 (N_3590,N_3006,N_3103);
nor U3591 (N_3591,N_3340,N_3266);
or U3592 (N_3592,N_3375,N_3000);
xor U3593 (N_3593,N_3427,N_3440);
xnor U3594 (N_3594,N_3222,N_3086);
or U3595 (N_3595,N_3245,N_3431);
or U3596 (N_3596,N_3240,N_3338);
xnor U3597 (N_3597,N_3213,N_3056);
nor U3598 (N_3598,N_3320,N_3332);
nand U3599 (N_3599,N_3099,N_3219);
and U3600 (N_3600,N_3195,N_3048);
xnor U3601 (N_3601,N_3026,N_3060);
xnor U3602 (N_3602,N_3029,N_3087);
nor U3603 (N_3603,N_3100,N_3211);
nor U3604 (N_3604,N_3248,N_3167);
nor U3605 (N_3605,N_3361,N_3235);
xnor U3606 (N_3606,N_3295,N_3175);
or U3607 (N_3607,N_3477,N_3474);
and U3608 (N_3608,N_3479,N_3271);
nand U3609 (N_3609,N_3118,N_3166);
or U3610 (N_3610,N_3260,N_3491);
nor U3611 (N_3611,N_3268,N_3498);
or U3612 (N_3612,N_3168,N_3259);
nor U3613 (N_3613,N_3371,N_3257);
nand U3614 (N_3614,N_3122,N_3054);
nor U3615 (N_3615,N_3487,N_3098);
nor U3616 (N_3616,N_3097,N_3179);
nand U3617 (N_3617,N_3232,N_3357);
nand U3618 (N_3618,N_3241,N_3101);
nor U3619 (N_3619,N_3132,N_3403);
nand U3620 (N_3620,N_3472,N_3112);
nor U3621 (N_3621,N_3409,N_3312);
nor U3622 (N_3622,N_3315,N_3478);
xor U3623 (N_3623,N_3082,N_3215);
nor U3624 (N_3624,N_3164,N_3163);
nor U3625 (N_3625,N_3465,N_3150);
or U3626 (N_3626,N_3469,N_3193);
nand U3627 (N_3627,N_3064,N_3172);
nand U3628 (N_3628,N_3496,N_3149);
or U3629 (N_3629,N_3300,N_3121);
nand U3630 (N_3630,N_3273,N_3244);
xor U3631 (N_3631,N_3439,N_3186);
nor U3632 (N_3632,N_3314,N_3243);
nor U3633 (N_3633,N_3313,N_3279);
xnor U3634 (N_3634,N_3490,N_3050);
or U3635 (N_3635,N_3094,N_3367);
and U3636 (N_3636,N_3220,N_3297);
xnor U3637 (N_3637,N_3301,N_3025);
nand U3638 (N_3638,N_3238,N_3210);
or U3639 (N_3639,N_3139,N_3457);
and U3640 (N_3640,N_3202,N_3432);
xor U3641 (N_3641,N_3383,N_3481);
xnor U3642 (N_3642,N_3372,N_3125);
or U3643 (N_3643,N_3382,N_3015);
and U3644 (N_3644,N_3200,N_3486);
nor U3645 (N_3645,N_3458,N_3108);
nand U3646 (N_3646,N_3126,N_3324);
nor U3647 (N_3647,N_3285,N_3061);
and U3648 (N_3648,N_3090,N_3258);
or U3649 (N_3649,N_3148,N_3187);
or U3650 (N_3650,N_3229,N_3206);
nand U3651 (N_3651,N_3253,N_3047);
or U3652 (N_3652,N_3467,N_3347);
nor U3653 (N_3653,N_3045,N_3304);
and U3654 (N_3654,N_3441,N_3377);
and U3655 (N_3655,N_3454,N_3321);
and U3656 (N_3656,N_3370,N_3303);
or U3657 (N_3657,N_3120,N_3328);
or U3658 (N_3658,N_3444,N_3230);
nand U3659 (N_3659,N_3443,N_3398);
nand U3660 (N_3660,N_3071,N_3146);
or U3661 (N_3661,N_3231,N_3406);
and U3662 (N_3662,N_3282,N_3072);
nor U3663 (N_3663,N_3305,N_3436);
nor U3664 (N_3664,N_3133,N_3204);
and U3665 (N_3665,N_3073,N_3468);
or U3666 (N_3666,N_3093,N_3201);
xor U3667 (N_3667,N_3002,N_3374);
nand U3668 (N_3668,N_3451,N_3323);
nor U3669 (N_3669,N_3442,N_3463);
nand U3670 (N_3670,N_3007,N_3169);
or U3671 (N_3671,N_3318,N_3250);
xnor U3672 (N_3672,N_3343,N_3391);
nand U3673 (N_3673,N_3115,N_3308);
nand U3674 (N_3674,N_3396,N_3480);
or U3675 (N_3675,N_3325,N_3041);
nor U3676 (N_3676,N_3450,N_3397);
or U3677 (N_3677,N_3294,N_3184);
and U3678 (N_3678,N_3008,N_3395);
and U3679 (N_3679,N_3205,N_3042);
and U3680 (N_3680,N_3485,N_3363);
and U3681 (N_3681,N_3066,N_3272);
xnor U3682 (N_3682,N_3199,N_3178);
nor U3683 (N_3683,N_3390,N_3411);
or U3684 (N_3684,N_3336,N_3156);
xor U3685 (N_3685,N_3104,N_3012);
xnor U3686 (N_3686,N_3043,N_3326);
xor U3687 (N_3687,N_3052,N_3197);
and U3688 (N_3688,N_3384,N_3192);
and U3689 (N_3689,N_3331,N_3019);
xor U3690 (N_3690,N_3130,N_3117);
or U3691 (N_3691,N_3425,N_3280);
nor U3692 (N_3692,N_3158,N_3437);
xor U3693 (N_3693,N_3165,N_3296);
xnor U3694 (N_3694,N_3154,N_3309);
nand U3695 (N_3695,N_3119,N_3005);
or U3696 (N_3696,N_3218,N_3277);
and U3697 (N_3697,N_3424,N_3208);
and U3698 (N_3698,N_3247,N_3417);
nor U3699 (N_3699,N_3378,N_3177);
nand U3700 (N_3700,N_3489,N_3004);
and U3701 (N_3701,N_3236,N_3092);
xnor U3702 (N_3702,N_3227,N_3022);
or U3703 (N_3703,N_3270,N_3410);
or U3704 (N_3704,N_3107,N_3423);
or U3705 (N_3705,N_3251,N_3488);
nand U3706 (N_3706,N_3038,N_3341);
and U3707 (N_3707,N_3141,N_3142);
nor U3708 (N_3708,N_3322,N_3143);
or U3709 (N_3709,N_3327,N_3335);
nand U3710 (N_3710,N_3024,N_3144);
or U3711 (N_3711,N_3426,N_3360);
or U3712 (N_3712,N_3001,N_3185);
nor U3713 (N_3713,N_3267,N_3483);
xnor U3714 (N_3714,N_3059,N_3413);
or U3715 (N_3715,N_3350,N_3032);
and U3716 (N_3716,N_3040,N_3388);
and U3717 (N_3717,N_3339,N_3077);
and U3718 (N_3718,N_3136,N_3140);
and U3719 (N_3719,N_3445,N_3473);
nand U3720 (N_3720,N_3291,N_3289);
or U3721 (N_3721,N_3009,N_3044);
and U3722 (N_3722,N_3080,N_3070);
or U3723 (N_3723,N_3228,N_3036);
nand U3724 (N_3724,N_3288,N_3292);
or U3725 (N_3725,N_3307,N_3462);
nand U3726 (N_3726,N_3113,N_3023);
nor U3727 (N_3727,N_3065,N_3265);
xnor U3728 (N_3728,N_3196,N_3014);
xor U3729 (N_3729,N_3387,N_3449);
nand U3730 (N_3730,N_3362,N_3147);
or U3731 (N_3731,N_3404,N_3345);
and U3732 (N_3732,N_3416,N_3484);
and U3733 (N_3733,N_3290,N_3329);
nand U3734 (N_3734,N_3171,N_3128);
and U3735 (N_3735,N_3138,N_3319);
and U3736 (N_3736,N_3223,N_3190);
nand U3737 (N_3737,N_3482,N_3124);
xnor U3738 (N_3738,N_3137,N_3460);
nand U3739 (N_3739,N_3365,N_3461);
nand U3740 (N_3740,N_3355,N_3421);
nand U3741 (N_3741,N_3182,N_3435);
nand U3742 (N_3742,N_3225,N_3293);
and U3743 (N_3743,N_3078,N_3284);
xor U3744 (N_3744,N_3039,N_3224);
nand U3745 (N_3745,N_3281,N_3452);
and U3746 (N_3746,N_3356,N_3476);
xor U3747 (N_3747,N_3470,N_3494);
and U3748 (N_3748,N_3110,N_3131);
xor U3749 (N_3749,N_3214,N_3216);
xnor U3750 (N_3750,N_3192,N_3228);
and U3751 (N_3751,N_3389,N_3405);
xnor U3752 (N_3752,N_3012,N_3114);
nor U3753 (N_3753,N_3399,N_3416);
or U3754 (N_3754,N_3094,N_3234);
nor U3755 (N_3755,N_3393,N_3473);
xor U3756 (N_3756,N_3376,N_3354);
and U3757 (N_3757,N_3135,N_3491);
nand U3758 (N_3758,N_3458,N_3435);
nor U3759 (N_3759,N_3347,N_3435);
nand U3760 (N_3760,N_3258,N_3400);
and U3761 (N_3761,N_3464,N_3121);
and U3762 (N_3762,N_3060,N_3374);
nand U3763 (N_3763,N_3072,N_3191);
or U3764 (N_3764,N_3106,N_3274);
xnor U3765 (N_3765,N_3268,N_3267);
xor U3766 (N_3766,N_3482,N_3446);
or U3767 (N_3767,N_3328,N_3457);
nand U3768 (N_3768,N_3238,N_3064);
xor U3769 (N_3769,N_3283,N_3452);
nand U3770 (N_3770,N_3459,N_3086);
nand U3771 (N_3771,N_3277,N_3165);
xor U3772 (N_3772,N_3347,N_3379);
xnor U3773 (N_3773,N_3463,N_3486);
nor U3774 (N_3774,N_3471,N_3378);
or U3775 (N_3775,N_3086,N_3207);
nor U3776 (N_3776,N_3039,N_3381);
or U3777 (N_3777,N_3289,N_3047);
and U3778 (N_3778,N_3393,N_3410);
nand U3779 (N_3779,N_3050,N_3148);
and U3780 (N_3780,N_3399,N_3238);
nand U3781 (N_3781,N_3201,N_3132);
and U3782 (N_3782,N_3159,N_3005);
and U3783 (N_3783,N_3241,N_3267);
and U3784 (N_3784,N_3437,N_3257);
or U3785 (N_3785,N_3181,N_3204);
nand U3786 (N_3786,N_3442,N_3346);
xnor U3787 (N_3787,N_3304,N_3240);
nand U3788 (N_3788,N_3296,N_3181);
and U3789 (N_3789,N_3023,N_3351);
or U3790 (N_3790,N_3147,N_3328);
nand U3791 (N_3791,N_3272,N_3299);
xnor U3792 (N_3792,N_3313,N_3014);
nor U3793 (N_3793,N_3378,N_3035);
or U3794 (N_3794,N_3454,N_3433);
nand U3795 (N_3795,N_3181,N_3455);
xnor U3796 (N_3796,N_3316,N_3383);
or U3797 (N_3797,N_3125,N_3160);
and U3798 (N_3798,N_3296,N_3192);
or U3799 (N_3799,N_3297,N_3298);
or U3800 (N_3800,N_3270,N_3380);
and U3801 (N_3801,N_3328,N_3378);
nand U3802 (N_3802,N_3183,N_3397);
nor U3803 (N_3803,N_3368,N_3434);
xor U3804 (N_3804,N_3038,N_3100);
nand U3805 (N_3805,N_3233,N_3039);
xnor U3806 (N_3806,N_3450,N_3161);
and U3807 (N_3807,N_3455,N_3276);
or U3808 (N_3808,N_3455,N_3077);
nor U3809 (N_3809,N_3352,N_3299);
nand U3810 (N_3810,N_3193,N_3270);
nand U3811 (N_3811,N_3203,N_3263);
xor U3812 (N_3812,N_3173,N_3360);
nand U3813 (N_3813,N_3253,N_3240);
and U3814 (N_3814,N_3297,N_3440);
or U3815 (N_3815,N_3468,N_3406);
xor U3816 (N_3816,N_3490,N_3321);
xor U3817 (N_3817,N_3079,N_3174);
nor U3818 (N_3818,N_3172,N_3315);
xor U3819 (N_3819,N_3442,N_3322);
and U3820 (N_3820,N_3222,N_3238);
or U3821 (N_3821,N_3313,N_3420);
and U3822 (N_3822,N_3321,N_3419);
xnor U3823 (N_3823,N_3140,N_3465);
or U3824 (N_3824,N_3158,N_3084);
or U3825 (N_3825,N_3350,N_3163);
nor U3826 (N_3826,N_3256,N_3282);
and U3827 (N_3827,N_3338,N_3347);
or U3828 (N_3828,N_3258,N_3155);
nand U3829 (N_3829,N_3032,N_3060);
or U3830 (N_3830,N_3157,N_3114);
nor U3831 (N_3831,N_3246,N_3397);
nand U3832 (N_3832,N_3430,N_3482);
and U3833 (N_3833,N_3019,N_3230);
or U3834 (N_3834,N_3027,N_3349);
xor U3835 (N_3835,N_3197,N_3206);
or U3836 (N_3836,N_3110,N_3497);
xnor U3837 (N_3837,N_3415,N_3033);
nor U3838 (N_3838,N_3475,N_3022);
or U3839 (N_3839,N_3049,N_3220);
nand U3840 (N_3840,N_3146,N_3461);
or U3841 (N_3841,N_3392,N_3228);
nor U3842 (N_3842,N_3447,N_3371);
nand U3843 (N_3843,N_3306,N_3262);
or U3844 (N_3844,N_3095,N_3491);
and U3845 (N_3845,N_3126,N_3478);
nand U3846 (N_3846,N_3063,N_3266);
xor U3847 (N_3847,N_3356,N_3061);
nand U3848 (N_3848,N_3477,N_3287);
nor U3849 (N_3849,N_3027,N_3199);
nor U3850 (N_3850,N_3365,N_3307);
nand U3851 (N_3851,N_3415,N_3320);
xor U3852 (N_3852,N_3426,N_3029);
and U3853 (N_3853,N_3223,N_3228);
and U3854 (N_3854,N_3321,N_3359);
nand U3855 (N_3855,N_3069,N_3361);
or U3856 (N_3856,N_3063,N_3494);
and U3857 (N_3857,N_3122,N_3410);
and U3858 (N_3858,N_3337,N_3317);
nand U3859 (N_3859,N_3071,N_3020);
or U3860 (N_3860,N_3259,N_3306);
xnor U3861 (N_3861,N_3000,N_3322);
and U3862 (N_3862,N_3018,N_3049);
xor U3863 (N_3863,N_3060,N_3178);
nand U3864 (N_3864,N_3331,N_3199);
nand U3865 (N_3865,N_3095,N_3168);
xor U3866 (N_3866,N_3063,N_3282);
and U3867 (N_3867,N_3235,N_3468);
and U3868 (N_3868,N_3144,N_3097);
and U3869 (N_3869,N_3308,N_3338);
xnor U3870 (N_3870,N_3325,N_3294);
nor U3871 (N_3871,N_3488,N_3409);
xnor U3872 (N_3872,N_3069,N_3451);
xor U3873 (N_3873,N_3221,N_3060);
or U3874 (N_3874,N_3314,N_3269);
or U3875 (N_3875,N_3135,N_3073);
or U3876 (N_3876,N_3060,N_3421);
xor U3877 (N_3877,N_3104,N_3300);
and U3878 (N_3878,N_3021,N_3018);
nand U3879 (N_3879,N_3284,N_3262);
or U3880 (N_3880,N_3302,N_3070);
and U3881 (N_3881,N_3024,N_3087);
or U3882 (N_3882,N_3355,N_3452);
or U3883 (N_3883,N_3345,N_3168);
nand U3884 (N_3884,N_3059,N_3357);
nand U3885 (N_3885,N_3415,N_3012);
and U3886 (N_3886,N_3218,N_3358);
and U3887 (N_3887,N_3402,N_3277);
nand U3888 (N_3888,N_3226,N_3475);
xor U3889 (N_3889,N_3074,N_3228);
and U3890 (N_3890,N_3088,N_3119);
nand U3891 (N_3891,N_3418,N_3320);
nor U3892 (N_3892,N_3363,N_3400);
xnor U3893 (N_3893,N_3484,N_3113);
nor U3894 (N_3894,N_3458,N_3248);
or U3895 (N_3895,N_3018,N_3065);
or U3896 (N_3896,N_3077,N_3142);
nand U3897 (N_3897,N_3264,N_3358);
nor U3898 (N_3898,N_3157,N_3146);
nand U3899 (N_3899,N_3318,N_3131);
nor U3900 (N_3900,N_3263,N_3184);
nand U3901 (N_3901,N_3108,N_3102);
or U3902 (N_3902,N_3057,N_3039);
nand U3903 (N_3903,N_3324,N_3110);
nor U3904 (N_3904,N_3093,N_3013);
nor U3905 (N_3905,N_3162,N_3138);
or U3906 (N_3906,N_3394,N_3015);
and U3907 (N_3907,N_3175,N_3445);
nor U3908 (N_3908,N_3327,N_3239);
xnor U3909 (N_3909,N_3051,N_3038);
and U3910 (N_3910,N_3263,N_3226);
or U3911 (N_3911,N_3332,N_3052);
nor U3912 (N_3912,N_3184,N_3361);
or U3913 (N_3913,N_3423,N_3085);
nor U3914 (N_3914,N_3097,N_3356);
and U3915 (N_3915,N_3082,N_3302);
nand U3916 (N_3916,N_3037,N_3489);
or U3917 (N_3917,N_3276,N_3402);
or U3918 (N_3918,N_3426,N_3345);
xor U3919 (N_3919,N_3460,N_3344);
nand U3920 (N_3920,N_3353,N_3103);
nand U3921 (N_3921,N_3340,N_3099);
nand U3922 (N_3922,N_3491,N_3186);
nor U3923 (N_3923,N_3220,N_3218);
or U3924 (N_3924,N_3400,N_3407);
xor U3925 (N_3925,N_3275,N_3066);
and U3926 (N_3926,N_3116,N_3321);
xnor U3927 (N_3927,N_3245,N_3119);
or U3928 (N_3928,N_3031,N_3415);
or U3929 (N_3929,N_3070,N_3365);
or U3930 (N_3930,N_3455,N_3066);
or U3931 (N_3931,N_3290,N_3324);
and U3932 (N_3932,N_3142,N_3380);
and U3933 (N_3933,N_3017,N_3238);
nand U3934 (N_3934,N_3496,N_3376);
xor U3935 (N_3935,N_3289,N_3076);
or U3936 (N_3936,N_3394,N_3100);
or U3937 (N_3937,N_3424,N_3163);
and U3938 (N_3938,N_3275,N_3276);
nand U3939 (N_3939,N_3120,N_3384);
nand U3940 (N_3940,N_3442,N_3399);
and U3941 (N_3941,N_3090,N_3041);
nor U3942 (N_3942,N_3277,N_3132);
nor U3943 (N_3943,N_3137,N_3023);
xnor U3944 (N_3944,N_3224,N_3408);
and U3945 (N_3945,N_3124,N_3461);
nor U3946 (N_3946,N_3374,N_3093);
nor U3947 (N_3947,N_3348,N_3461);
nand U3948 (N_3948,N_3129,N_3405);
xor U3949 (N_3949,N_3202,N_3427);
and U3950 (N_3950,N_3404,N_3027);
nand U3951 (N_3951,N_3053,N_3454);
and U3952 (N_3952,N_3358,N_3291);
nor U3953 (N_3953,N_3031,N_3368);
nor U3954 (N_3954,N_3377,N_3001);
nor U3955 (N_3955,N_3044,N_3438);
xnor U3956 (N_3956,N_3248,N_3082);
nand U3957 (N_3957,N_3463,N_3254);
nor U3958 (N_3958,N_3369,N_3396);
xor U3959 (N_3959,N_3495,N_3192);
and U3960 (N_3960,N_3428,N_3198);
or U3961 (N_3961,N_3467,N_3201);
and U3962 (N_3962,N_3184,N_3412);
or U3963 (N_3963,N_3480,N_3443);
xor U3964 (N_3964,N_3169,N_3416);
xnor U3965 (N_3965,N_3087,N_3454);
xnor U3966 (N_3966,N_3299,N_3070);
and U3967 (N_3967,N_3294,N_3164);
and U3968 (N_3968,N_3332,N_3244);
nand U3969 (N_3969,N_3100,N_3095);
nand U3970 (N_3970,N_3114,N_3140);
or U3971 (N_3971,N_3148,N_3024);
nand U3972 (N_3972,N_3396,N_3166);
nand U3973 (N_3973,N_3106,N_3424);
and U3974 (N_3974,N_3194,N_3299);
or U3975 (N_3975,N_3217,N_3422);
nor U3976 (N_3976,N_3293,N_3335);
nor U3977 (N_3977,N_3111,N_3374);
and U3978 (N_3978,N_3461,N_3476);
xnor U3979 (N_3979,N_3238,N_3167);
and U3980 (N_3980,N_3170,N_3449);
nor U3981 (N_3981,N_3456,N_3437);
nor U3982 (N_3982,N_3311,N_3207);
xnor U3983 (N_3983,N_3289,N_3152);
xnor U3984 (N_3984,N_3084,N_3124);
or U3985 (N_3985,N_3341,N_3145);
nand U3986 (N_3986,N_3354,N_3114);
and U3987 (N_3987,N_3402,N_3383);
nand U3988 (N_3988,N_3161,N_3235);
nor U3989 (N_3989,N_3023,N_3366);
nand U3990 (N_3990,N_3098,N_3443);
and U3991 (N_3991,N_3083,N_3397);
nand U3992 (N_3992,N_3294,N_3414);
nor U3993 (N_3993,N_3454,N_3209);
or U3994 (N_3994,N_3425,N_3215);
nor U3995 (N_3995,N_3205,N_3307);
or U3996 (N_3996,N_3310,N_3485);
nor U3997 (N_3997,N_3065,N_3257);
xnor U3998 (N_3998,N_3461,N_3222);
xor U3999 (N_3999,N_3472,N_3382);
xnor U4000 (N_4000,N_3645,N_3643);
xor U4001 (N_4001,N_3752,N_3728);
xor U4002 (N_4002,N_3859,N_3541);
or U4003 (N_4003,N_3780,N_3990);
xor U4004 (N_4004,N_3914,N_3705);
or U4005 (N_4005,N_3825,N_3678);
nand U4006 (N_4006,N_3816,N_3900);
nand U4007 (N_4007,N_3945,N_3547);
and U4008 (N_4008,N_3763,N_3776);
nand U4009 (N_4009,N_3996,N_3946);
nor U4010 (N_4010,N_3543,N_3591);
and U4011 (N_4011,N_3867,N_3978);
nor U4012 (N_4012,N_3896,N_3762);
xnor U4013 (N_4013,N_3759,N_3821);
nor U4014 (N_4014,N_3999,N_3722);
nand U4015 (N_4015,N_3516,N_3976);
nor U4016 (N_4016,N_3842,N_3784);
and U4017 (N_4017,N_3607,N_3693);
nor U4018 (N_4018,N_3672,N_3659);
xnor U4019 (N_4019,N_3875,N_3570);
nor U4020 (N_4020,N_3950,N_3932);
and U4021 (N_4021,N_3868,N_3563);
xor U4022 (N_4022,N_3593,N_3831);
and U4023 (N_4023,N_3505,N_3519);
nand U4024 (N_4024,N_3699,N_3847);
nor U4025 (N_4025,N_3841,N_3796);
and U4026 (N_4026,N_3617,N_3998);
xor U4027 (N_4027,N_3974,N_3857);
xnor U4028 (N_4028,N_3530,N_3740);
nor U4029 (N_4029,N_3665,N_3807);
nor U4030 (N_4030,N_3908,N_3749);
nand U4031 (N_4031,N_3524,N_3626);
nor U4032 (N_4032,N_3971,N_3551);
nand U4033 (N_4033,N_3818,N_3734);
and U4034 (N_4034,N_3791,N_3986);
nand U4035 (N_4035,N_3627,N_3721);
nand U4036 (N_4036,N_3619,N_3692);
xor U4037 (N_4037,N_3545,N_3904);
or U4038 (N_4038,N_3700,N_3797);
and U4039 (N_4039,N_3603,N_3711);
xor U4040 (N_4040,N_3792,N_3891);
and U4041 (N_4041,N_3755,N_3624);
or U4042 (N_4042,N_3641,N_3544);
xnor U4043 (N_4043,N_3913,N_3997);
xor U4044 (N_4044,N_3980,N_3592);
xor U4045 (N_4045,N_3751,N_3909);
nand U4046 (N_4046,N_3778,N_3512);
nand U4047 (N_4047,N_3561,N_3725);
nand U4048 (N_4048,N_3528,N_3680);
nor U4049 (N_4049,N_3892,N_3515);
xnor U4050 (N_4050,N_3565,N_3871);
xor U4051 (N_4051,N_3719,N_3685);
or U4052 (N_4052,N_3869,N_3691);
xnor U4053 (N_4053,N_3742,N_3992);
and U4054 (N_4054,N_3853,N_3511);
nand U4055 (N_4055,N_3523,N_3884);
xor U4056 (N_4056,N_3761,N_3596);
nand U4057 (N_4057,N_3750,N_3723);
nor U4058 (N_4058,N_3798,N_3712);
and U4059 (N_4059,N_3707,N_3564);
nand U4060 (N_4060,N_3736,N_3915);
nor U4061 (N_4061,N_3845,N_3687);
nand U4062 (N_4062,N_3850,N_3625);
nor U4063 (N_4063,N_3985,N_3872);
or U4064 (N_4064,N_3575,N_3925);
nand U4065 (N_4065,N_3959,N_3704);
and U4066 (N_4066,N_3927,N_3767);
nand U4067 (N_4067,N_3739,N_3788);
nor U4068 (N_4068,N_3956,N_3832);
nand U4069 (N_4069,N_3538,N_3890);
and U4070 (N_4070,N_3566,N_3741);
nor U4071 (N_4071,N_3569,N_3953);
nand U4072 (N_4072,N_3888,N_3826);
nor U4073 (N_4073,N_3638,N_3907);
nor U4074 (N_4074,N_3531,N_3688);
xnor U4075 (N_4075,N_3866,N_3506);
nand U4076 (N_4076,N_3865,N_3929);
or U4077 (N_4077,N_3588,N_3982);
xnor U4078 (N_4078,N_3880,N_3783);
and U4079 (N_4079,N_3676,N_3558);
xnor U4080 (N_4080,N_3955,N_3681);
and U4081 (N_4081,N_3962,N_3585);
or U4082 (N_4082,N_3604,N_3620);
xor U4083 (N_4083,N_3537,N_3616);
nand U4084 (N_4084,N_3924,N_3514);
or U4085 (N_4085,N_3942,N_3785);
nand U4086 (N_4086,N_3631,N_3597);
nand U4087 (N_4087,N_3799,N_3735);
and U4088 (N_4088,N_3636,N_3557);
xnor U4089 (N_4089,N_3768,N_3964);
nand U4090 (N_4090,N_3656,N_3658);
nand U4091 (N_4091,N_3600,N_3910);
nand U4092 (N_4092,N_3652,N_3937);
nand U4093 (N_4093,N_3614,N_3833);
and U4094 (N_4094,N_3640,N_3876);
xnor U4095 (N_4095,N_3567,N_3805);
and U4096 (N_4096,N_3520,N_3727);
nand U4097 (N_4097,N_3782,N_3529);
nor U4098 (N_4098,N_3777,N_3500);
xor U4099 (N_4099,N_3916,N_3969);
and U4100 (N_4100,N_3510,N_3527);
and U4101 (N_4101,N_3670,N_3877);
nand U4102 (N_4102,N_3606,N_3525);
xor U4103 (N_4103,N_3613,N_3917);
xor U4104 (N_4104,N_3760,N_3503);
and U4105 (N_4105,N_3828,N_3772);
and U4106 (N_4106,N_3758,N_3695);
xor U4107 (N_4107,N_3773,N_3562);
or U4108 (N_4108,N_3864,N_3651);
and U4109 (N_4109,N_3765,N_3581);
and U4110 (N_4110,N_3926,N_3897);
nand U4111 (N_4111,N_3729,N_3663);
nor U4112 (N_4112,N_3809,N_3838);
or U4113 (N_4113,N_3682,N_3786);
xnor U4114 (N_4114,N_3673,N_3854);
and U4115 (N_4115,N_3852,N_3851);
or U4116 (N_4116,N_3817,N_3931);
and U4117 (N_4117,N_3815,N_3630);
nand U4118 (N_4118,N_3963,N_3689);
xor U4119 (N_4119,N_3844,N_3883);
xor U4120 (N_4120,N_3993,N_3919);
xnor U4121 (N_4121,N_3770,N_3814);
nand U4122 (N_4122,N_3612,N_3846);
and U4123 (N_4123,N_3595,N_3889);
or U4124 (N_4124,N_3733,N_3660);
nand U4125 (N_4125,N_3881,N_3552);
nand U4126 (N_4126,N_3899,N_3666);
nand U4127 (N_4127,N_3677,N_3608);
nand U4128 (N_4128,N_3771,N_3517);
and U4129 (N_4129,N_3579,N_3732);
xnor U4130 (N_4130,N_3646,N_3582);
or U4131 (N_4131,N_3995,N_3981);
or U4132 (N_4132,N_3820,N_3701);
nor U4133 (N_4133,N_3860,N_3745);
xnor U4134 (N_4134,N_3720,N_3615);
nand U4135 (N_4135,N_3674,N_3983);
nand U4136 (N_4136,N_3954,N_3921);
nand U4137 (N_4137,N_3922,N_3573);
or U4138 (N_4138,N_3709,N_3873);
or U4139 (N_4139,N_3977,N_3539);
or U4140 (N_4140,N_3715,N_3975);
xnor U4141 (N_4141,N_3835,N_3827);
nand U4142 (N_4142,N_3843,N_3710);
nor U4143 (N_4143,N_3605,N_3787);
nand U4144 (N_4144,N_3560,N_3632);
xor U4145 (N_4145,N_3572,N_3518);
or U4146 (N_4146,N_3858,N_3936);
and U4147 (N_4147,N_3882,N_3789);
nand U4148 (N_4148,N_3795,N_3639);
and U4149 (N_4149,N_3637,N_3634);
nor U4150 (N_4150,N_3994,N_3583);
nor U4151 (N_4151,N_3513,N_3848);
and U4152 (N_4152,N_3804,N_3928);
nor U4153 (N_4153,N_3895,N_3703);
nor U4154 (N_4154,N_3911,N_3716);
nand U4155 (N_4155,N_3933,N_3781);
or U4156 (N_4156,N_3568,N_3584);
xnor U4157 (N_4157,N_3669,N_3708);
and U4158 (N_4158,N_3526,N_3675);
or U4159 (N_4159,N_3961,N_3822);
xor U4160 (N_4160,N_3879,N_3930);
nor U4161 (N_4161,N_3856,N_3939);
and U4162 (N_4162,N_3629,N_3793);
nor U4163 (N_4163,N_3935,N_3702);
nand U4164 (N_4164,N_3878,N_3988);
or U4165 (N_4165,N_3943,N_3991);
nor U4166 (N_4166,N_3553,N_3802);
xor U4167 (N_4167,N_3574,N_3813);
nor U4168 (N_4168,N_3863,N_3548);
and U4169 (N_4169,N_3586,N_3958);
or U4170 (N_4170,N_3622,N_3714);
and U4171 (N_4171,N_3902,N_3775);
and U4172 (N_4172,N_3746,N_3849);
nand U4173 (N_4173,N_3657,N_3599);
and U4174 (N_4174,N_3987,N_3536);
or U4175 (N_4175,N_3790,N_3801);
xor U4176 (N_4176,N_3508,N_3509);
nor U4177 (N_4177,N_3559,N_3979);
xnor U4178 (N_4178,N_3960,N_3923);
nor U4179 (N_4179,N_3706,N_3803);
nand U4180 (N_4180,N_3973,N_3912);
and U4181 (N_4181,N_3502,N_3812);
or U4182 (N_4182,N_3920,N_3968);
xnor U4183 (N_4183,N_3521,N_3686);
nand U4184 (N_4184,N_3903,N_3578);
or U4185 (N_4185,N_3941,N_3829);
xor U4186 (N_4186,N_3522,N_3717);
and U4187 (N_4187,N_3940,N_3535);
nor U4188 (N_4188,N_3984,N_3808);
xnor U4189 (N_4189,N_3683,N_3748);
and U4190 (N_4190,N_3664,N_3696);
xor U4191 (N_4191,N_3794,N_3504);
nand U4192 (N_4192,N_3747,N_3671);
nand U4193 (N_4193,N_3555,N_3800);
and U4194 (N_4194,N_3662,N_3824);
xor U4195 (N_4195,N_3901,N_3743);
and U4196 (N_4196,N_3764,N_3769);
xor U4197 (N_4197,N_3823,N_3577);
and U4198 (N_4198,N_3886,N_3546);
xor U4199 (N_4199,N_3730,N_3655);
xnor U4200 (N_4200,N_3554,N_3757);
nand U4201 (N_4201,N_3806,N_3906);
nor U4202 (N_4202,N_3837,N_3944);
xor U4203 (N_4203,N_3744,N_3724);
nor U4204 (N_4204,N_3644,N_3861);
or U4205 (N_4205,N_3590,N_3726);
or U4206 (N_4206,N_3507,N_3811);
and U4207 (N_4207,N_3628,N_3623);
xor U4208 (N_4208,N_3779,N_3839);
or U4209 (N_4209,N_3947,N_3810);
nor U4210 (N_4210,N_3874,N_3753);
or U4211 (N_4211,N_3949,N_3556);
nor U4212 (N_4212,N_3952,N_3594);
nand U4213 (N_4213,N_3649,N_3967);
nor U4214 (N_4214,N_3836,N_3862);
nand U4215 (N_4215,N_3690,N_3642);
xor U4216 (N_4216,N_3948,N_3766);
xor U4217 (N_4217,N_3965,N_3855);
nand U4218 (N_4218,N_3601,N_3635);
or U4219 (N_4219,N_3576,N_3887);
nor U4220 (N_4220,N_3972,N_3679);
or U4221 (N_4221,N_3542,N_3870);
or U4222 (N_4222,N_3737,N_3534);
or U4223 (N_4223,N_3694,N_3905);
xor U4224 (N_4224,N_3830,N_3938);
and U4225 (N_4225,N_3587,N_3501);
xnor U4226 (N_4226,N_3571,N_3934);
nor U4227 (N_4227,N_3667,N_3540);
nand U4228 (N_4228,N_3738,N_3648);
nor U4229 (N_4229,N_3610,N_3633);
or U4230 (N_4230,N_3653,N_3650);
nor U4231 (N_4231,N_3754,N_3698);
or U4232 (N_4232,N_3621,N_3598);
or U4233 (N_4233,N_3951,N_3966);
nor U4234 (N_4234,N_3731,N_3989);
nor U4235 (N_4235,N_3894,N_3893);
or U4236 (N_4236,N_3618,N_3549);
nor U4237 (N_4237,N_3654,N_3713);
nand U4238 (N_4238,N_3602,N_3589);
nor U4239 (N_4239,N_3647,N_3611);
nor U4240 (N_4240,N_3533,N_3898);
or U4241 (N_4241,N_3957,N_3774);
nor U4242 (N_4242,N_3668,N_3834);
or U4243 (N_4243,N_3609,N_3580);
nand U4244 (N_4244,N_3970,N_3756);
nor U4245 (N_4245,N_3819,N_3718);
nor U4246 (N_4246,N_3532,N_3684);
or U4247 (N_4247,N_3697,N_3840);
nand U4248 (N_4248,N_3661,N_3550);
nand U4249 (N_4249,N_3918,N_3885);
and U4250 (N_4250,N_3502,N_3815);
or U4251 (N_4251,N_3658,N_3580);
xor U4252 (N_4252,N_3546,N_3656);
or U4253 (N_4253,N_3622,N_3728);
or U4254 (N_4254,N_3737,N_3920);
xnor U4255 (N_4255,N_3561,N_3744);
xor U4256 (N_4256,N_3570,N_3709);
nand U4257 (N_4257,N_3963,N_3741);
or U4258 (N_4258,N_3542,N_3729);
xnor U4259 (N_4259,N_3827,N_3843);
xor U4260 (N_4260,N_3852,N_3983);
and U4261 (N_4261,N_3856,N_3671);
nor U4262 (N_4262,N_3779,N_3509);
nor U4263 (N_4263,N_3654,N_3639);
nor U4264 (N_4264,N_3903,N_3717);
xor U4265 (N_4265,N_3566,N_3767);
and U4266 (N_4266,N_3901,N_3523);
xor U4267 (N_4267,N_3707,N_3680);
nor U4268 (N_4268,N_3507,N_3566);
nor U4269 (N_4269,N_3690,N_3522);
xnor U4270 (N_4270,N_3539,N_3880);
and U4271 (N_4271,N_3611,N_3961);
xnor U4272 (N_4272,N_3960,N_3517);
xor U4273 (N_4273,N_3534,N_3673);
and U4274 (N_4274,N_3678,N_3883);
or U4275 (N_4275,N_3666,N_3737);
or U4276 (N_4276,N_3808,N_3871);
xor U4277 (N_4277,N_3700,N_3710);
and U4278 (N_4278,N_3987,N_3861);
nor U4279 (N_4279,N_3748,N_3853);
xnor U4280 (N_4280,N_3737,N_3719);
or U4281 (N_4281,N_3766,N_3527);
or U4282 (N_4282,N_3750,N_3641);
nor U4283 (N_4283,N_3889,N_3846);
nand U4284 (N_4284,N_3801,N_3898);
nand U4285 (N_4285,N_3792,N_3635);
and U4286 (N_4286,N_3867,N_3822);
nor U4287 (N_4287,N_3821,N_3995);
nand U4288 (N_4288,N_3604,N_3808);
xor U4289 (N_4289,N_3942,N_3531);
and U4290 (N_4290,N_3762,N_3717);
nand U4291 (N_4291,N_3722,N_3949);
nand U4292 (N_4292,N_3711,N_3508);
nand U4293 (N_4293,N_3906,N_3509);
xnor U4294 (N_4294,N_3635,N_3818);
and U4295 (N_4295,N_3932,N_3937);
or U4296 (N_4296,N_3690,N_3550);
and U4297 (N_4297,N_3633,N_3688);
nor U4298 (N_4298,N_3729,N_3905);
or U4299 (N_4299,N_3859,N_3513);
or U4300 (N_4300,N_3694,N_3681);
or U4301 (N_4301,N_3768,N_3624);
or U4302 (N_4302,N_3716,N_3908);
or U4303 (N_4303,N_3845,N_3980);
nand U4304 (N_4304,N_3867,N_3926);
xnor U4305 (N_4305,N_3508,N_3922);
xor U4306 (N_4306,N_3749,N_3568);
nand U4307 (N_4307,N_3722,N_3836);
nor U4308 (N_4308,N_3696,N_3978);
nand U4309 (N_4309,N_3731,N_3601);
or U4310 (N_4310,N_3821,N_3620);
xnor U4311 (N_4311,N_3754,N_3703);
or U4312 (N_4312,N_3580,N_3858);
and U4313 (N_4313,N_3874,N_3804);
nand U4314 (N_4314,N_3574,N_3828);
xnor U4315 (N_4315,N_3809,N_3589);
or U4316 (N_4316,N_3708,N_3945);
and U4317 (N_4317,N_3769,N_3923);
xor U4318 (N_4318,N_3611,N_3613);
xor U4319 (N_4319,N_3556,N_3939);
xnor U4320 (N_4320,N_3713,N_3990);
or U4321 (N_4321,N_3799,N_3738);
nor U4322 (N_4322,N_3773,N_3830);
or U4323 (N_4323,N_3829,N_3921);
and U4324 (N_4324,N_3791,N_3807);
nand U4325 (N_4325,N_3730,N_3783);
xnor U4326 (N_4326,N_3615,N_3574);
nand U4327 (N_4327,N_3717,N_3993);
nand U4328 (N_4328,N_3962,N_3611);
or U4329 (N_4329,N_3953,N_3962);
nor U4330 (N_4330,N_3923,N_3971);
or U4331 (N_4331,N_3914,N_3827);
or U4332 (N_4332,N_3795,N_3859);
nand U4333 (N_4333,N_3835,N_3852);
nand U4334 (N_4334,N_3800,N_3759);
nand U4335 (N_4335,N_3954,N_3995);
and U4336 (N_4336,N_3614,N_3862);
xnor U4337 (N_4337,N_3602,N_3630);
xnor U4338 (N_4338,N_3684,N_3689);
and U4339 (N_4339,N_3584,N_3963);
or U4340 (N_4340,N_3808,N_3506);
and U4341 (N_4341,N_3982,N_3728);
nand U4342 (N_4342,N_3639,N_3660);
nand U4343 (N_4343,N_3519,N_3847);
nor U4344 (N_4344,N_3701,N_3707);
and U4345 (N_4345,N_3720,N_3505);
nand U4346 (N_4346,N_3941,N_3813);
xor U4347 (N_4347,N_3614,N_3660);
and U4348 (N_4348,N_3504,N_3882);
nand U4349 (N_4349,N_3694,N_3944);
or U4350 (N_4350,N_3760,N_3881);
xnor U4351 (N_4351,N_3501,N_3675);
nor U4352 (N_4352,N_3843,N_3553);
and U4353 (N_4353,N_3640,N_3938);
nor U4354 (N_4354,N_3657,N_3600);
nand U4355 (N_4355,N_3550,N_3804);
nand U4356 (N_4356,N_3612,N_3989);
nor U4357 (N_4357,N_3610,N_3662);
or U4358 (N_4358,N_3973,N_3547);
xnor U4359 (N_4359,N_3703,N_3598);
nand U4360 (N_4360,N_3547,N_3743);
or U4361 (N_4361,N_3792,N_3706);
or U4362 (N_4362,N_3596,N_3911);
and U4363 (N_4363,N_3679,N_3784);
and U4364 (N_4364,N_3592,N_3822);
xnor U4365 (N_4365,N_3746,N_3588);
nand U4366 (N_4366,N_3934,N_3522);
xor U4367 (N_4367,N_3620,N_3873);
nor U4368 (N_4368,N_3563,N_3798);
nor U4369 (N_4369,N_3744,N_3810);
and U4370 (N_4370,N_3905,N_3636);
xor U4371 (N_4371,N_3568,N_3937);
and U4372 (N_4372,N_3728,N_3717);
nor U4373 (N_4373,N_3770,N_3508);
and U4374 (N_4374,N_3844,N_3531);
or U4375 (N_4375,N_3553,N_3885);
and U4376 (N_4376,N_3836,N_3679);
nand U4377 (N_4377,N_3838,N_3570);
xor U4378 (N_4378,N_3747,N_3880);
or U4379 (N_4379,N_3677,N_3727);
nor U4380 (N_4380,N_3806,N_3637);
and U4381 (N_4381,N_3758,N_3741);
and U4382 (N_4382,N_3824,N_3550);
nand U4383 (N_4383,N_3939,N_3836);
or U4384 (N_4384,N_3592,N_3728);
nor U4385 (N_4385,N_3691,N_3758);
or U4386 (N_4386,N_3960,N_3650);
nor U4387 (N_4387,N_3899,N_3596);
nand U4388 (N_4388,N_3591,N_3910);
nand U4389 (N_4389,N_3803,N_3641);
and U4390 (N_4390,N_3683,N_3558);
nand U4391 (N_4391,N_3869,N_3998);
nor U4392 (N_4392,N_3678,N_3663);
nand U4393 (N_4393,N_3732,N_3516);
or U4394 (N_4394,N_3914,N_3527);
xor U4395 (N_4395,N_3667,N_3998);
and U4396 (N_4396,N_3707,N_3827);
or U4397 (N_4397,N_3800,N_3997);
xnor U4398 (N_4398,N_3969,N_3890);
or U4399 (N_4399,N_3926,N_3741);
xor U4400 (N_4400,N_3914,N_3609);
nand U4401 (N_4401,N_3735,N_3542);
nor U4402 (N_4402,N_3752,N_3716);
nand U4403 (N_4403,N_3620,N_3639);
nand U4404 (N_4404,N_3714,N_3825);
and U4405 (N_4405,N_3750,N_3698);
and U4406 (N_4406,N_3932,N_3609);
xnor U4407 (N_4407,N_3862,N_3870);
nor U4408 (N_4408,N_3984,N_3959);
and U4409 (N_4409,N_3789,N_3634);
and U4410 (N_4410,N_3786,N_3577);
nor U4411 (N_4411,N_3842,N_3712);
nand U4412 (N_4412,N_3936,N_3745);
nor U4413 (N_4413,N_3751,N_3797);
xnor U4414 (N_4414,N_3929,N_3969);
nor U4415 (N_4415,N_3519,N_3718);
xor U4416 (N_4416,N_3529,N_3527);
nand U4417 (N_4417,N_3601,N_3543);
nor U4418 (N_4418,N_3878,N_3766);
nor U4419 (N_4419,N_3891,N_3564);
xor U4420 (N_4420,N_3659,N_3547);
nand U4421 (N_4421,N_3566,N_3563);
xor U4422 (N_4422,N_3977,N_3671);
nor U4423 (N_4423,N_3876,N_3539);
and U4424 (N_4424,N_3934,N_3955);
nand U4425 (N_4425,N_3793,N_3807);
and U4426 (N_4426,N_3764,N_3521);
nor U4427 (N_4427,N_3957,N_3942);
nand U4428 (N_4428,N_3647,N_3674);
and U4429 (N_4429,N_3607,N_3743);
xnor U4430 (N_4430,N_3947,N_3901);
and U4431 (N_4431,N_3770,N_3609);
nand U4432 (N_4432,N_3563,N_3668);
or U4433 (N_4433,N_3650,N_3870);
and U4434 (N_4434,N_3690,N_3787);
and U4435 (N_4435,N_3595,N_3764);
or U4436 (N_4436,N_3660,N_3579);
nor U4437 (N_4437,N_3614,N_3603);
and U4438 (N_4438,N_3784,N_3686);
and U4439 (N_4439,N_3796,N_3544);
and U4440 (N_4440,N_3619,N_3613);
nor U4441 (N_4441,N_3966,N_3624);
or U4442 (N_4442,N_3819,N_3587);
nor U4443 (N_4443,N_3854,N_3917);
nor U4444 (N_4444,N_3851,N_3819);
xor U4445 (N_4445,N_3934,N_3815);
nand U4446 (N_4446,N_3930,N_3714);
nor U4447 (N_4447,N_3626,N_3614);
or U4448 (N_4448,N_3556,N_3960);
xor U4449 (N_4449,N_3620,N_3510);
or U4450 (N_4450,N_3760,N_3903);
nand U4451 (N_4451,N_3641,N_3672);
or U4452 (N_4452,N_3684,N_3573);
nor U4453 (N_4453,N_3603,N_3595);
nand U4454 (N_4454,N_3859,N_3931);
xnor U4455 (N_4455,N_3716,N_3628);
xor U4456 (N_4456,N_3929,N_3800);
nor U4457 (N_4457,N_3568,N_3880);
and U4458 (N_4458,N_3600,N_3740);
xor U4459 (N_4459,N_3695,N_3820);
and U4460 (N_4460,N_3658,N_3961);
nand U4461 (N_4461,N_3964,N_3946);
nor U4462 (N_4462,N_3985,N_3725);
nor U4463 (N_4463,N_3766,N_3787);
xnor U4464 (N_4464,N_3839,N_3772);
xor U4465 (N_4465,N_3737,N_3764);
and U4466 (N_4466,N_3828,N_3645);
or U4467 (N_4467,N_3694,N_3855);
nand U4468 (N_4468,N_3716,N_3909);
nor U4469 (N_4469,N_3845,N_3924);
nand U4470 (N_4470,N_3954,N_3508);
and U4471 (N_4471,N_3954,N_3774);
nand U4472 (N_4472,N_3637,N_3959);
xnor U4473 (N_4473,N_3915,N_3651);
nand U4474 (N_4474,N_3892,N_3889);
or U4475 (N_4475,N_3550,N_3739);
xnor U4476 (N_4476,N_3954,N_3700);
nor U4477 (N_4477,N_3873,N_3515);
xnor U4478 (N_4478,N_3869,N_3669);
nand U4479 (N_4479,N_3759,N_3854);
nand U4480 (N_4480,N_3675,N_3518);
nand U4481 (N_4481,N_3532,N_3528);
nor U4482 (N_4482,N_3722,N_3657);
nor U4483 (N_4483,N_3963,N_3919);
xor U4484 (N_4484,N_3999,N_3935);
or U4485 (N_4485,N_3848,N_3706);
nand U4486 (N_4486,N_3525,N_3637);
xor U4487 (N_4487,N_3641,N_3606);
xnor U4488 (N_4488,N_3690,N_3921);
or U4489 (N_4489,N_3731,N_3910);
nand U4490 (N_4490,N_3899,N_3779);
xnor U4491 (N_4491,N_3535,N_3662);
nand U4492 (N_4492,N_3815,N_3729);
and U4493 (N_4493,N_3696,N_3538);
or U4494 (N_4494,N_3860,N_3764);
nand U4495 (N_4495,N_3643,N_3960);
and U4496 (N_4496,N_3701,N_3573);
or U4497 (N_4497,N_3936,N_3917);
or U4498 (N_4498,N_3591,N_3991);
and U4499 (N_4499,N_3568,N_3816);
nor U4500 (N_4500,N_4064,N_4202);
and U4501 (N_4501,N_4407,N_4375);
nand U4502 (N_4502,N_4044,N_4179);
and U4503 (N_4503,N_4317,N_4242);
nand U4504 (N_4504,N_4409,N_4394);
nand U4505 (N_4505,N_4494,N_4476);
or U4506 (N_4506,N_4014,N_4303);
xor U4507 (N_4507,N_4445,N_4269);
nor U4508 (N_4508,N_4092,N_4116);
nor U4509 (N_4509,N_4049,N_4389);
and U4510 (N_4510,N_4336,N_4109);
nand U4511 (N_4511,N_4368,N_4361);
nor U4512 (N_4512,N_4231,N_4395);
and U4513 (N_4513,N_4381,N_4369);
and U4514 (N_4514,N_4308,N_4316);
and U4515 (N_4515,N_4186,N_4021);
or U4516 (N_4516,N_4459,N_4222);
nand U4517 (N_4517,N_4278,N_4335);
nor U4518 (N_4518,N_4319,N_4047);
and U4519 (N_4519,N_4396,N_4161);
nand U4520 (N_4520,N_4059,N_4280);
nor U4521 (N_4521,N_4226,N_4441);
or U4522 (N_4522,N_4305,N_4166);
xor U4523 (N_4523,N_4119,N_4456);
xnor U4524 (N_4524,N_4432,N_4066);
nand U4525 (N_4525,N_4003,N_4374);
and U4526 (N_4526,N_4204,N_4053);
or U4527 (N_4527,N_4073,N_4302);
nor U4528 (N_4528,N_4209,N_4127);
and U4529 (N_4529,N_4069,N_4031);
nand U4530 (N_4530,N_4098,N_4344);
and U4531 (N_4531,N_4100,N_4266);
xnor U4532 (N_4532,N_4193,N_4417);
nand U4533 (N_4533,N_4214,N_4356);
or U4534 (N_4534,N_4249,N_4210);
xnor U4535 (N_4535,N_4435,N_4194);
xor U4536 (N_4536,N_4474,N_4181);
nand U4537 (N_4537,N_4144,N_4176);
nor U4538 (N_4538,N_4485,N_4399);
or U4539 (N_4539,N_4279,N_4205);
nor U4540 (N_4540,N_4165,N_4036);
nor U4541 (N_4541,N_4220,N_4271);
or U4542 (N_4542,N_4172,N_4486);
xnor U4543 (N_4543,N_4248,N_4182);
xor U4544 (N_4544,N_4203,N_4253);
nor U4545 (N_4545,N_4262,N_4246);
xor U4546 (N_4546,N_4338,N_4065);
nor U4547 (N_4547,N_4255,N_4217);
nor U4548 (N_4548,N_4174,N_4081);
and U4549 (N_4549,N_4112,N_4102);
and U4550 (N_4550,N_4461,N_4232);
nor U4551 (N_4551,N_4083,N_4184);
nor U4552 (N_4552,N_4314,N_4015);
and U4553 (N_4553,N_4243,N_4267);
nand U4554 (N_4554,N_4121,N_4043);
nand U4555 (N_4555,N_4228,N_4283);
or U4556 (N_4556,N_4439,N_4364);
xor U4557 (N_4557,N_4434,N_4345);
nand U4558 (N_4558,N_4088,N_4062);
xnor U4559 (N_4559,N_4078,N_4117);
xnor U4560 (N_4560,N_4240,N_4216);
nand U4561 (N_4561,N_4151,N_4192);
or U4562 (N_4562,N_4340,N_4051);
nand U4563 (N_4563,N_4200,N_4114);
and U4564 (N_4564,N_4334,N_4311);
nor U4565 (N_4565,N_4061,N_4351);
and U4566 (N_4566,N_4348,N_4390);
xnor U4567 (N_4567,N_4157,N_4056);
nand U4568 (N_4568,N_4199,N_4449);
nor U4569 (N_4569,N_4089,N_4006);
nand U4570 (N_4570,N_4341,N_4067);
and U4571 (N_4571,N_4022,N_4004);
nor U4572 (N_4572,N_4481,N_4190);
nand U4573 (N_4573,N_4388,N_4495);
nor U4574 (N_4574,N_4385,N_4413);
and U4575 (N_4575,N_4325,N_4008);
nand U4576 (N_4576,N_4419,N_4373);
and U4577 (N_4577,N_4086,N_4471);
nand U4578 (N_4578,N_4162,N_4294);
or U4579 (N_4579,N_4484,N_4028);
nand U4580 (N_4580,N_4163,N_4468);
nor U4581 (N_4581,N_4300,N_4422);
xnor U4582 (N_4582,N_4158,N_4141);
and U4583 (N_4583,N_4401,N_4378);
or U4584 (N_4584,N_4025,N_4017);
and U4585 (N_4585,N_4082,N_4332);
nor U4586 (N_4586,N_4213,N_4196);
and U4587 (N_4587,N_4387,N_4357);
nor U4588 (N_4588,N_4264,N_4403);
xnor U4589 (N_4589,N_4129,N_4398);
xnor U4590 (N_4590,N_4223,N_4307);
nand U4591 (N_4591,N_4175,N_4324);
nand U4592 (N_4592,N_4463,N_4482);
nand U4593 (N_4593,N_4293,N_4133);
or U4594 (N_4594,N_4415,N_4406);
nor U4595 (N_4595,N_4189,N_4230);
xor U4596 (N_4596,N_4152,N_4490);
nor U4597 (N_4597,N_4421,N_4339);
or U4598 (N_4598,N_4450,N_4171);
and U4599 (N_4599,N_4315,N_4355);
nand U4600 (N_4600,N_4383,N_4460);
xnor U4601 (N_4601,N_4104,N_4297);
and U4602 (N_4602,N_4273,N_4328);
or U4603 (N_4603,N_4270,N_4070);
nand U4604 (N_4604,N_4148,N_4370);
xnor U4605 (N_4605,N_4237,N_4411);
xor U4606 (N_4606,N_4147,N_4054);
and U4607 (N_4607,N_4333,N_4290);
or U4608 (N_4608,N_4020,N_4350);
and U4609 (N_4609,N_4447,N_4198);
xnor U4610 (N_4610,N_4052,N_4000);
or U4611 (N_4611,N_4349,N_4236);
xor U4612 (N_4612,N_4298,N_4386);
nor U4613 (N_4613,N_4030,N_4160);
or U4614 (N_4614,N_4026,N_4252);
and U4615 (N_4615,N_4466,N_4420);
nor U4616 (N_4616,N_4058,N_4397);
and U4617 (N_4617,N_4306,N_4090);
xnor U4618 (N_4618,N_4212,N_4009);
or U4619 (N_4619,N_4483,N_4238);
and U4620 (N_4620,N_4042,N_4312);
nor U4621 (N_4621,N_4405,N_4096);
xor U4622 (N_4622,N_4208,N_4080);
xor U4623 (N_4623,N_4060,N_4299);
xor U4624 (N_4624,N_4363,N_4288);
nand U4625 (N_4625,N_4124,N_4478);
nand U4626 (N_4626,N_4256,N_4140);
xor U4627 (N_4627,N_4095,N_4110);
xnor U4628 (N_4628,N_4154,N_4408);
and U4629 (N_4629,N_4097,N_4472);
xor U4630 (N_4630,N_4277,N_4392);
and U4631 (N_4631,N_4296,N_4219);
and U4632 (N_4632,N_4428,N_4019);
nor U4633 (N_4633,N_4491,N_4126);
and U4634 (N_4634,N_4477,N_4170);
xnor U4635 (N_4635,N_4427,N_4135);
nor U4636 (N_4636,N_4146,N_4499);
nor U4637 (N_4637,N_4108,N_4120);
or U4638 (N_4638,N_4470,N_4446);
xor U4639 (N_4639,N_4313,N_4412);
nor U4640 (N_4640,N_4462,N_4101);
and U4641 (N_4641,N_4139,N_4115);
and U4642 (N_4642,N_4143,N_4286);
and U4643 (N_4643,N_4429,N_4444);
and U4644 (N_4644,N_4010,N_4035);
xor U4645 (N_4645,N_4431,N_4099);
nand U4646 (N_4646,N_4045,N_4048);
nand U4647 (N_4647,N_4016,N_4041);
nor U4648 (N_4648,N_4259,N_4057);
or U4649 (N_4649,N_4234,N_4034);
xnor U4650 (N_4650,N_4012,N_4379);
or U4651 (N_4651,N_4168,N_4454);
or U4652 (N_4652,N_4177,N_4467);
nor U4653 (N_4653,N_4245,N_4261);
xnor U4654 (N_4654,N_4346,N_4365);
and U4655 (N_4655,N_4377,N_4440);
xnor U4656 (N_4656,N_4111,N_4107);
nand U4657 (N_4657,N_4072,N_4155);
xor U4658 (N_4658,N_4138,N_4360);
or U4659 (N_4659,N_4282,N_4137);
and U4660 (N_4660,N_4367,N_4169);
or U4661 (N_4661,N_4153,N_4076);
xnor U4662 (N_4662,N_4159,N_4487);
or U4663 (N_4663,N_4426,N_4024);
xor U4664 (N_4664,N_4023,N_4458);
nor U4665 (N_4665,N_4007,N_4465);
or U4666 (N_4666,N_4268,N_4448);
or U4667 (N_4667,N_4391,N_4173);
xor U4668 (N_4668,N_4241,N_4233);
or U4669 (N_4669,N_4145,N_4229);
and U4670 (N_4670,N_4105,N_4063);
and U4671 (N_4671,N_4106,N_4272);
and U4672 (N_4672,N_4206,N_4275);
or U4673 (N_4673,N_4301,N_4156);
or U4674 (N_4674,N_4164,N_4480);
nand U4675 (N_4675,N_4018,N_4257);
nor U4676 (N_4676,N_4260,N_4074);
or U4677 (N_4677,N_4352,N_4443);
xnor U4678 (N_4678,N_4221,N_4050);
xor U4679 (N_4679,N_4414,N_4284);
or U4680 (N_4680,N_4320,N_4195);
nand U4681 (N_4681,N_4211,N_4055);
xor U4682 (N_4682,N_4005,N_4416);
xor U4683 (N_4683,N_4473,N_4442);
nor U4684 (N_4684,N_4436,N_4464);
nand U4685 (N_4685,N_4038,N_4492);
or U4686 (N_4686,N_4091,N_4469);
nand U4687 (N_4687,N_4359,N_4289);
nand U4688 (N_4688,N_4027,N_4455);
xnor U4689 (N_4689,N_4430,N_4488);
nor U4690 (N_4690,N_4292,N_4437);
nor U4691 (N_4691,N_4479,N_4453);
and U4692 (N_4692,N_4384,N_4225);
nor U4693 (N_4693,N_4358,N_4281);
nor U4694 (N_4694,N_4489,N_4207);
nor U4695 (N_4695,N_4250,N_4029);
nand U4696 (N_4696,N_4244,N_4167);
and U4697 (N_4697,N_4239,N_4497);
nand U4698 (N_4698,N_4258,N_4118);
or U4699 (N_4699,N_4039,N_4263);
nor U4700 (N_4700,N_4400,N_4093);
nor U4701 (N_4701,N_4149,N_4180);
and U4702 (N_4702,N_4404,N_4410);
and U4703 (N_4703,N_4295,N_4329);
and U4704 (N_4704,N_4011,N_4046);
or U4705 (N_4705,N_4376,N_4457);
and U4706 (N_4706,N_4493,N_4254);
nand U4707 (N_4707,N_4122,N_4321);
and U4708 (N_4708,N_4496,N_4188);
nor U4709 (N_4709,N_4276,N_4247);
xor U4710 (N_4710,N_4347,N_4433);
nor U4711 (N_4711,N_4310,N_4094);
and U4712 (N_4712,N_4274,N_4071);
and U4713 (N_4713,N_4326,N_4224);
and U4714 (N_4714,N_4132,N_4185);
or U4715 (N_4715,N_4150,N_4013);
and U4716 (N_4716,N_4451,N_4418);
or U4717 (N_4717,N_4113,N_4131);
nor U4718 (N_4718,N_4130,N_4309);
nor U4719 (N_4719,N_4372,N_4291);
or U4720 (N_4720,N_4123,N_4380);
or U4721 (N_4721,N_4475,N_4215);
nor U4722 (N_4722,N_4218,N_4285);
or U4723 (N_4723,N_4342,N_4498);
xnor U4724 (N_4724,N_4197,N_4323);
nor U4725 (N_4725,N_4187,N_4134);
nand U4726 (N_4726,N_4075,N_4235);
nand U4727 (N_4727,N_4085,N_4304);
nand U4728 (N_4728,N_4002,N_4354);
or U4729 (N_4729,N_4327,N_4318);
and U4730 (N_4730,N_4183,N_4201);
xor U4731 (N_4731,N_4125,N_4079);
or U4732 (N_4732,N_4068,N_4424);
nand U4733 (N_4733,N_4251,N_4191);
and U4734 (N_4734,N_4371,N_4084);
nor U4735 (N_4735,N_4362,N_4337);
nand U4736 (N_4736,N_4438,N_4402);
xnor U4737 (N_4737,N_4382,N_4033);
or U4738 (N_4738,N_4322,N_4425);
nor U4739 (N_4739,N_4330,N_4142);
xnor U4740 (N_4740,N_4178,N_4032);
nor U4741 (N_4741,N_4040,N_4001);
nor U4742 (N_4742,N_4452,N_4366);
xor U4743 (N_4743,N_4077,N_4265);
nor U4744 (N_4744,N_4353,N_4128);
nor U4745 (N_4745,N_4227,N_4343);
nand U4746 (N_4746,N_4331,N_4103);
and U4747 (N_4747,N_4037,N_4423);
nand U4748 (N_4748,N_4393,N_4087);
or U4749 (N_4749,N_4136,N_4287);
and U4750 (N_4750,N_4000,N_4144);
or U4751 (N_4751,N_4247,N_4413);
xor U4752 (N_4752,N_4098,N_4391);
nand U4753 (N_4753,N_4304,N_4136);
and U4754 (N_4754,N_4236,N_4278);
xor U4755 (N_4755,N_4063,N_4228);
nor U4756 (N_4756,N_4306,N_4473);
xnor U4757 (N_4757,N_4368,N_4193);
nor U4758 (N_4758,N_4459,N_4294);
nand U4759 (N_4759,N_4447,N_4452);
xnor U4760 (N_4760,N_4148,N_4351);
nor U4761 (N_4761,N_4017,N_4151);
nand U4762 (N_4762,N_4062,N_4051);
or U4763 (N_4763,N_4234,N_4088);
xor U4764 (N_4764,N_4171,N_4193);
and U4765 (N_4765,N_4177,N_4484);
xnor U4766 (N_4766,N_4359,N_4104);
xnor U4767 (N_4767,N_4109,N_4356);
xnor U4768 (N_4768,N_4170,N_4463);
xor U4769 (N_4769,N_4130,N_4028);
or U4770 (N_4770,N_4071,N_4304);
or U4771 (N_4771,N_4314,N_4398);
nand U4772 (N_4772,N_4463,N_4039);
and U4773 (N_4773,N_4043,N_4352);
or U4774 (N_4774,N_4006,N_4339);
and U4775 (N_4775,N_4120,N_4099);
or U4776 (N_4776,N_4259,N_4211);
xnor U4777 (N_4777,N_4046,N_4258);
or U4778 (N_4778,N_4449,N_4270);
or U4779 (N_4779,N_4320,N_4001);
nand U4780 (N_4780,N_4194,N_4316);
or U4781 (N_4781,N_4478,N_4463);
nand U4782 (N_4782,N_4438,N_4259);
nand U4783 (N_4783,N_4353,N_4002);
nor U4784 (N_4784,N_4082,N_4268);
nor U4785 (N_4785,N_4310,N_4308);
xnor U4786 (N_4786,N_4367,N_4174);
xor U4787 (N_4787,N_4379,N_4056);
xor U4788 (N_4788,N_4251,N_4313);
or U4789 (N_4789,N_4467,N_4158);
xnor U4790 (N_4790,N_4386,N_4013);
nor U4791 (N_4791,N_4418,N_4098);
xor U4792 (N_4792,N_4418,N_4072);
xnor U4793 (N_4793,N_4002,N_4088);
nand U4794 (N_4794,N_4006,N_4184);
nor U4795 (N_4795,N_4261,N_4195);
and U4796 (N_4796,N_4030,N_4456);
nor U4797 (N_4797,N_4144,N_4368);
or U4798 (N_4798,N_4328,N_4164);
nand U4799 (N_4799,N_4186,N_4382);
or U4800 (N_4800,N_4157,N_4437);
or U4801 (N_4801,N_4062,N_4150);
or U4802 (N_4802,N_4033,N_4362);
or U4803 (N_4803,N_4342,N_4448);
and U4804 (N_4804,N_4460,N_4320);
xor U4805 (N_4805,N_4081,N_4328);
or U4806 (N_4806,N_4264,N_4174);
nor U4807 (N_4807,N_4103,N_4037);
nor U4808 (N_4808,N_4057,N_4255);
nor U4809 (N_4809,N_4323,N_4340);
xnor U4810 (N_4810,N_4399,N_4210);
xnor U4811 (N_4811,N_4378,N_4282);
xor U4812 (N_4812,N_4102,N_4354);
nand U4813 (N_4813,N_4145,N_4425);
and U4814 (N_4814,N_4055,N_4428);
and U4815 (N_4815,N_4061,N_4101);
xnor U4816 (N_4816,N_4035,N_4497);
nand U4817 (N_4817,N_4301,N_4247);
xor U4818 (N_4818,N_4315,N_4232);
xor U4819 (N_4819,N_4422,N_4455);
xor U4820 (N_4820,N_4364,N_4426);
or U4821 (N_4821,N_4384,N_4282);
or U4822 (N_4822,N_4057,N_4406);
and U4823 (N_4823,N_4446,N_4034);
nor U4824 (N_4824,N_4211,N_4407);
nor U4825 (N_4825,N_4011,N_4107);
nor U4826 (N_4826,N_4374,N_4115);
or U4827 (N_4827,N_4080,N_4387);
or U4828 (N_4828,N_4333,N_4010);
nor U4829 (N_4829,N_4422,N_4254);
nand U4830 (N_4830,N_4199,N_4411);
nor U4831 (N_4831,N_4003,N_4261);
and U4832 (N_4832,N_4438,N_4140);
and U4833 (N_4833,N_4047,N_4343);
nor U4834 (N_4834,N_4449,N_4031);
or U4835 (N_4835,N_4271,N_4341);
or U4836 (N_4836,N_4410,N_4320);
xnor U4837 (N_4837,N_4470,N_4365);
nand U4838 (N_4838,N_4092,N_4128);
nand U4839 (N_4839,N_4115,N_4474);
or U4840 (N_4840,N_4255,N_4332);
nand U4841 (N_4841,N_4301,N_4395);
xor U4842 (N_4842,N_4339,N_4168);
nor U4843 (N_4843,N_4467,N_4421);
or U4844 (N_4844,N_4348,N_4467);
xor U4845 (N_4845,N_4251,N_4493);
nand U4846 (N_4846,N_4283,N_4303);
nor U4847 (N_4847,N_4180,N_4035);
or U4848 (N_4848,N_4227,N_4463);
nor U4849 (N_4849,N_4066,N_4368);
nor U4850 (N_4850,N_4355,N_4323);
nand U4851 (N_4851,N_4373,N_4366);
xor U4852 (N_4852,N_4237,N_4287);
nor U4853 (N_4853,N_4390,N_4221);
nand U4854 (N_4854,N_4205,N_4389);
or U4855 (N_4855,N_4068,N_4314);
or U4856 (N_4856,N_4290,N_4154);
and U4857 (N_4857,N_4040,N_4200);
nor U4858 (N_4858,N_4308,N_4346);
xnor U4859 (N_4859,N_4312,N_4015);
xnor U4860 (N_4860,N_4350,N_4461);
or U4861 (N_4861,N_4425,N_4035);
nand U4862 (N_4862,N_4422,N_4240);
or U4863 (N_4863,N_4198,N_4190);
nand U4864 (N_4864,N_4496,N_4290);
or U4865 (N_4865,N_4184,N_4357);
xnor U4866 (N_4866,N_4415,N_4157);
nand U4867 (N_4867,N_4181,N_4411);
and U4868 (N_4868,N_4445,N_4162);
or U4869 (N_4869,N_4021,N_4304);
nor U4870 (N_4870,N_4094,N_4237);
and U4871 (N_4871,N_4377,N_4159);
nand U4872 (N_4872,N_4339,N_4211);
and U4873 (N_4873,N_4259,N_4386);
nor U4874 (N_4874,N_4005,N_4175);
and U4875 (N_4875,N_4457,N_4322);
or U4876 (N_4876,N_4166,N_4090);
or U4877 (N_4877,N_4067,N_4143);
or U4878 (N_4878,N_4387,N_4050);
and U4879 (N_4879,N_4211,N_4133);
xor U4880 (N_4880,N_4493,N_4484);
xnor U4881 (N_4881,N_4327,N_4101);
nand U4882 (N_4882,N_4229,N_4151);
and U4883 (N_4883,N_4267,N_4351);
xnor U4884 (N_4884,N_4467,N_4451);
xnor U4885 (N_4885,N_4360,N_4271);
nand U4886 (N_4886,N_4422,N_4465);
or U4887 (N_4887,N_4197,N_4283);
and U4888 (N_4888,N_4105,N_4147);
or U4889 (N_4889,N_4403,N_4229);
nand U4890 (N_4890,N_4043,N_4133);
nor U4891 (N_4891,N_4380,N_4473);
xnor U4892 (N_4892,N_4488,N_4448);
nand U4893 (N_4893,N_4203,N_4367);
or U4894 (N_4894,N_4110,N_4274);
xor U4895 (N_4895,N_4035,N_4424);
xnor U4896 (N_4896,N_4250,N_4099);
xor U4897 (N_4897,N_4318,N_4484);
xor U4898 (N_4898,N_4002,N_4367);
and U4899 (N_4899,N_4024,N_4030);
xor U4900 (N_4900,N_4049,N_4106);
nor U4901 (N_4901,N_4474,N_4272);
xnor U4902 (N_4902,N_4121,N_4184);
nand U4903 (N_4903,N_4338,N_4070);
or U4904 (N_4904,N_4420,N_4011);
nor U4905 (N_4905,N_4496,N_4001);
nor U4906 (N_4906,N_4224,N_4413);
xor U4907 (N_4907,N_4027,N_4306);
nor U4908 (N_4908,N_4137,N_4466);
xor U4909 (N_4909,N_4496,N_4193);
or U4910 (N_4910,N_4452,N_4266);
and U4911 (N_4911,N_4133,N_4396);
and U4912 (N_4912,N_4337,N_4479);
nand U4913 (N_4913,N_4301,N_4359);
or U4914 (N_4914,N_4126,N_4470);
nand U4915 (N_4915,N_4265,N_4043);
nor U4916 (N_4916,N_4137,N_4140);
nand U4917 (N_4917,N_4037,N_4144);
nand U4918 (N_4918,N_4227,N_4299);
nand U4919 (N_4919,N_4218,N_4226);
xor U4920 (N_4920,N_4039,N_4139);
or U4921 (N_4921,N_4166,N_4360);
nor U4922 (N_4922,N_4359,N_4012);
nor U4923 (N_4923,N_4394,N_4418);
nand U4924 (N_4924,N_4268,N_4436);
xor U4925 (N_4925,N_4205,N_4192);
and U4926 (N_4926,N_4123,N_4339);
nor U4927 (N_4927,N_4132,N_4495);
nor U4928 (N_4928,N_4269,N_4432);
xnor U4929 (N_4929,N_4428,N_4298);
nor U4930 (N_4930,N_4239,N_4318);
xnor U4931 (N_4931,N_4013,N_4320);
or U4932 (N_4932,N_4433,N_4451);
and U4933 (N_4933,N_4389,N_4089);
nand U4934 (N_4934,N_4174,N_4496);
and U4935 (N_4935,N_4009,N_4285);
xnor U4936 (N_4936,N_4350,N_4367);
nand U4937 (N_4937,N_4237,N_4218);
nor U4938 (N_4938,N_4313,N_4464);
xor U4939 (N_4939,N_4399,N_4217);
xnor U4940 (N_4940,N_4458,N_4326);
or U4941 (N_4941,N_4215,N_4123);
nand U4942 (N_4942,N_4414,N_4259);
or U4943 (N_4943,N_4430,N_4274);
nand U4944 (N_4944,N_4493,N_4280);
or U4945 (N_4945,N_4410,N_4450);
or U4946 (N_4946,N_4181,N_4448);
or U4947 (N_4947,N_4002,N_4390);
nand U4948 (N_4948,N_4026,N_4195);
and U4949 (N_4949,N_4031,N_4077);
xnor U4950 (N_4950,N_4395,N_4089);
nor U4951 (N_4951,N_4187,N_4277);
or U4952 (N_4952,N_4307,N_4194);
nand U4953 (N_4953,N_4323,N_4189);
and U4954 (N_4954,N_4329,N_4294);
nand U4955 (N_4955,N_4467,N_4385);
nand U4956 (N_4956,N_4155,N_4428);
nor U4957 (N_4957,N_4188,N_4030);
or U4958 (N_4958,N_4039,N_4325);
xnor U4959 (N_4959,N_4386,N_4304);
nor U4960 (N_4960,N_4251,N_4405);
and U4961 (N_4961,N_4185,N_4245);
nor U4962 (N_4962,N_4210,N_4466);
or U4963 (N_4963,N_4485,N_4157);
nor U4964 (N_4964,N_4437,N_4469);
and U4965 (N_4965,N_4450,N_4441);
and U4966 (N_4966,N_4058,N_4435);
or U4967 (N_4967,N_4328,N_4056);
or U4968 (N_4968,N_4010,N_4412);
xor U4969 (N_4969,N_4022,N_4445);
or U4970 (N_4970,N_4188,N_4148);
nand U4971 (N_4971,N_4150,N_4081);
xor U4972 (N_4972,N_4142,N_4073);
nand U4973 (N_4973,N_4450,N_4354);
or U4974 (N_4974,N_4447,N_4407);
nor U4975 (N_4975,N_4499,N_4217);
and U4976 (N_4976,N_4083,N_4390);
nor U4977 (N_4977,N_4053,N_4127);
and U4978 (N_4978,N_4222,N_4261);
xor U4979 (N_4979,N_4023,N_4457);
nor U4980 (N_4980,N_4348,N_4317);
or U4981 (N_4981,N_4361,N_4024);
nor U4982 (N_4982,N_4355,N_4402);
and U4983 (N_4983,N_4325,N_4311);
or U4984 (N_4984,N_4132,N_4027);
and U4985 (N_4985,N_4112,N_4276);
xnor U4986 (N_4986,N_4364,N_4149);
xnor U4987 (N_4987,N_4224,N_4060);
nor U4988 (N_4988,N_4301,N_4109);
nor U4989 (N_4989,N_4121,N_4050);
nor U4990 (N_4990,N_4407,N_4143);
xor U4991 (N_4991,N_4214,N_4052);
nand U4992 (N_4992,N_4043,N_4491);
nand U4993 (N_4993,N_4248,N_4264);
xor U4994 (N_4994,N_4107,N_4389);
xnor U4995 (N_4995,N_4422,N_4068);
and U4996 (N_4996,N_4355,N_4424);
or U4997 (N_4997,N_4393,N_4124);
and U4998 (N_4998,N_4400,N_4217);
xnor U4999 (N_4999,N_4178,N_4390);
and U5000 (N_5000,N_4705,N_4715);
nor U5001 (N_5001,N_4773,N_4893);
nand U5002 (N_5002,N_4993,N_4583);
or U5003 (N_5003,N_4915,N_4709);
or U5004 (N_5004,N_4854,N_4521);
nand U5005 (N_5005,N_4779,N_4607);
xor U5006 (N_5006,N_4562,N_4937);
xnor U5007 (N_5007,N_4615,N_4728);
and U5008 (N_5008,N_4957,N_4807);
xor U5009 (N_5009,N_4656,N_4929);
xor U5010 (N_5010,N_4727,N_4618);
nand U5011 (N_5011,N_4841,N_4590);
and U5012 (N_5012,N_4916,N_4701);
nor U5013 (N_5013,N_4850,N_4970);
or U5014 (N_5014,N_4644,N_4909);
and U5015 (N_5015,N_4611,N_4991);
nor U5016 (N_5016,N_4510,N_4710);
and U5017 (N_5017,N_4560,N_4787);
nand U5018 (N_5018,N_4878,N_4693);
and U5019 (N_5019,N_4828,N_4889);
xnor U5020 (N_5020,N_4913,N_4941);
nor U5021 (N_5021,N_4886,N_4997);
or U5022 (N_5022,N_4623,N_4758);
xnor U5023 (N_5023,N_4870,N_4509);
or U5024 (N_5024,N_4775,N_4637);
nor U5025 (N_5025,N_4872,N_4737);
xor U5026 (N_5026,N_4821,N_4795);
or U5027 (N_5027,N_4754,N_4662);
nand U5028 (N_5028,N_4565,N_4990);
xor U5029 (N_5029,N_4672,N_4899);
and U5030 (N_5030,N_4598,N_4516);
nand U5031 (N_5031,N_4620,N_4668);
nand U5032 (N_5032,N_4755,N_4926);
and U5033 (N_5033,N_4631,N_4684);
or U5034 (N_5034,N_4630,N_4740);
or U5035 (N_5035,N_4632,N_4679);
xnor U5036 (N_5036,N_4759,N_4503);
nand U5037 (N_5037,N_4624,N_4638);
nor U5038 (N_5038,N_4894,N_4603);
xor U5039 (N_5039,N_4946,N_4592);
xor U5040 (N_5040,N_4543,N_4525);
nand U5041 (N_5041,N_4535,N_4778);
nor U5042 (N_5042,N_4774,N_4702);
nand U5043 (N_5043,N_4971,N_4848);
xor U5044 (N_5044,N_4811,N_4805);
and U5045 (N_5045,N_4783,N_4829);
xor U5046 (N_5046,N_4748,N_4762);
nor U5047 (N_5047,N_4676,N_4548);
nand U5048 (N_5048,N_4515,N_4860);
and U5049 (N_5049,N_4981,N_4594);
nand U5050 (N_5050,N_4674,N_4648);
or U5051 (N_5051,N_4506,N_4746);
or U5052 (N_5052,N_4606,N_4939);
and U5053 (N_5053,N_4704,N_4985);
xor U5054 (N_5054,N_4921,N_4826);
nand U5055 (N_5055,N_4725,N_4585);
nand U5056 (N_5056,N_4742,N_4651);
xnor U5057 (N_5057,N_4905,N_4526);
and U5058 (N_5058,N_4852,N_4660);
or U5059 (N_5059,N_4661,N_4863);
and U5060 (N_5060,N_4527,N_4987);
and U5061 (N_5061,N_4643,N_4972);
and U5062 (N_5062,N_4599,N_4874);
xor U5063 (N_5063,N_4735,N_4883);
and U5064 (N_5064,N_4745,N_4726);
nand U5065 (N_5065,N_4875,N_4869);
nand U5066 (N_5066,N_4830,N_4782);
and U5067 (N_5067,N_4539,N_4804);
and U5068 (N_5068,N_4586,N_4511);
xor U5069 (N_5069,N_4865,N_4809);
nor U5070 (N_5070,N_4658,N_4540);
and U5071 (N_5071,N_4670,N_4563);
nand U5072 (N_5072,N_4791,N_4605);
nand U5073 (N_5073,N_4958,N_4923);
or U5074 (N_5074,N_4989,N_4906);
and U5075 (N_5075,N_4531,N_4880);
nor U5076 (N_5076,N_4538,N_4706);
and U5077 (N_5077,N_4723,N_4736);
nor U5078 (N_5078,N_4653,N_4743);
xor U5079 (N_5079,N_4873,N_4501);
nand U5080 (N_5080,N_4979,N_4690);
or U5081 (N_5081,N_4707,N_4956);
nand U5082 (N_5082,N_4943,N_4952);
and U5083 (N_5083,N_4823,N_4861);
nor U5084 (N_5084,N_4696,N_4980);
xnor U5085 (N_5085,N_4593,N_4918);
nor U5086 (N_5086,N_4832,N_4568);
nand U5087 (N_5087,N_4790,N_4776);
nor U5088 (N_5088,N_4581,N_4537);
and U5089 (N_5089,N_4756,N_4532);
or U5090 (N_5090,N_4671,N_4639);
nor U5091 (N_5091,N_4802,N_4842);
xor U5092 (N_5092,N_4810,N_4895);
nand U5093 (N_5093,N_4514,N_4719);
nor U5094 (N_5094,N_4757,N_4902);
nand U5095 (N_5095,N_4633,N_4851);
or U5096 (N_5096,N_4505,N_4798);
nor U5097 (N_5097,N_4720,N_4744);
and U5098 (N_5098,N_4610,N_4763);
and U5099 (N_5099,N_4819,N_4714);
nor U5100 (N_5100,N_4724,N_4984);
nor U5101 (N_5101,N_4730,N_4938);
and U5102 (N_5102,N_4688,N_4876);
nand U5103 (N_5103,N_4547,N_4645);
and U5104 (N_5104,N_4512,N_4888);
or U5105 (N_5105,N_4673,N_4945);
or U5106 (N_5106,N_4738,N_4846);
or U5107 (N_5107,N_4911,N_4621);
nor U5108 (N_5108,N_4649,N_4627);
and U5109 (N_5109,N_4556,N_4600);
nand U5110 (N_5110,N_4597,N_4867);
xnor U5111 (N_5111,N_4587,N_4817);
xor U5112 (N_5112,N_4544,N_4761);
nand U5113 (N_5113,N_4940,N_4733);
and U5114 (N_5114,N_4822,N_4617);
nor U5115 (N_5115,N_4741,N_4856);
or U5116 (N_5116,N_4732,N_4998);
and U5117 (N_5117,N_4519,N_4698);
nand U5118 (N_5118,N_4518,N_4978);
nand U5119 (N_5119,N_4849,N_4517);
xor U5120 (N_5120,N_4948,N_4584);
or U5121 (N_5121,N_4771,N_4847);
nand U5122 (N_5122,N_4625,N_4634);
nor U5123 (N_5123,N_4803,N_4764);
or U5124 (N_5124,N_4664,N_4609);
nor U5125 (N_5125,N_4930,N_4808);
nor U5126 (N_5126,N_4814,N_4781);
nor U5127 (N_5127,N_4654,N_4835);
nand U5128 (N_5128,N_4685,N_4722);
or U5129 (N_5129,N_4986,N_4784);
nand U5130 (N_5130,N_4932,N_4812);
or U5131 (N_5131,N_4753,N_4954);
nor U5132 (N_5132,N_4694,N_4749);
nand U5133 (N_5133,N_4833,N_4675);
and U5134 (N_5134,N_4965,N_4572);
nand U5135 (N_5135,N_4536,N_4504);
nand U5136 (N_5136,N_4928,N_4596);
xor U5137 (N_5137,N_4950,N_4765);
nor U5138 (N_5138,N_4949,N_4588);
nand U5139 (N_5139,N_4845,N_4569);
nand U5140 (N_5140,N_4574,N_4718);
and U5141 (N_5141,N_4642,N_4557);
or U5142 (N_5142,N_4864,N_4545);
and U5143 (N_5143,N_4935,N_4682);
nor U5144 (N_5144,N_4616,N_4549);
nand U5145 (N_5145,N_4602,N_4647);
nand U5146 (N_5146,N_4942,N_4799);
xor U5147 (N_5147,N_4667,N_4919);
xor U5148 (N_5148,N_4522,N_4559);
nor U5149 (N_5149,N_4831,N_4666);
xor U5150 (N_5150,N_4922,N_4968);
xor U5151 (N_5151,N_4751,N_4840);
and U5152 (N_5152,N_4962,N_4853);
nand U5153 (N_5153,N_4555,N_4579);
or U5154 (N_5154,N_4542,N_4974);
and U5155 (N_5155,N_4766,N_4975);
nor U5156 (N_5156,N_4750,N_4713);
nor U5157 (N_5157,N_4955,N_4772);
or U5158 (N_5158,N_4561,N_4691);
nor U5159 (N_5159,N_4961,N_4550);
or U5160 (N_5160,N_4862,N_4818);
and U5161 (N_5161,N_4825,N_4797);
nor U5162 (N_5162,N_4882,N_4747);
nand U5163 (N_5163,N_4612,N_4868);
or U5164 (N_5164,N_4892,N_4708);
nor U5165 (N_5165,N_4604,N_4580);
nand U5166 (N_5166,N_4881,N_4520);
and U5167 (N_5167,N_4683,N_4925);
and U5168 (N_5168,N_4964,N_4839);
nand U5169 (N_5169,N_4794,N_4793);
or U5170 (N_5170,N_4575,N_4796);
nor U5171 (N_5171,N_4900,N_4912);
nand U5172 (N_5172,N_4959,N_4677);
nor U5173 (N_5173,N_4837,N_4813);
or U5174 (N_5174,N_4988,N_4843);
nand U5175 (N_5175,N_4591,N_4785);
or U5176 (N_5176,N_4652,N_4657);
nor U5177 (N_5177,N_4871,N_4866);
xor U5178 (N_5178,N_4717,N_4689);
and U5179 (N_5179,N_4622,N_4554);
nand U5180 (N_5180,N_4760,N_4635);
xor U5181 (N_5181,N_4904,N_4963);
and U5182 (N_5182,N_4650,N_4801);
xnor U5183 (N_5183,N_4777,N_4951);
and U5184 (N_5184,N_4636,N_4884);
and U5185 (N_5185,N_4903,N_4663);
and U5186 (N_5186,N_4855,N_4827);
or U5187 (N_5187,N_4788,N_4995);
nor U5188 (N_5188,N_4992,N_4681);
xnor U5189 (N_5189,N_4578,N_4780);
nor U5190 (N_5190,N_4716,N_4769);
or U5191 (N_5191,N_4665,N_4834);
nor U5192 (N_5192,N_4524,N_4816);
xnor U5193 (N_5193,N_4699,N_4530);
xnor U5194 (N_5194,N_4815,N_4500);
nand U5195 (N_5195,N_4836,N_4507);
nand U5196 (N_5196,N_4541,N_4680);
and U5197 (N_5197,N_4570,N_4626);
xnor U5198 (N_5198,N_4857,N_4887);
nand U5199 (N_5199,N_4711,N_4721);
xor U5200 (N_5200,N_4973,N_4977);
nor U5201 (N_5201,N_4729,N_4891);
nor U5202 (N_5202,N_4695,N_4877);
nor U5203 (N_5203,N_4552,N_4901);
xor U5204 (N_5204,N_4933,N_4640);
nand U5205 (N_5205,N_4697,N_4551);
xor U5206 (N_5206,N_4800,N_4824);
or U5207 (N_5207,N_4792,N_4960);
xor U5208 (N_5208,N_4558,N_4924);
xor U5209 (N_5209,N_4994,N_4619);
and U5210 (N_5210,N_4983,N_4770);
and U5211 (N_5211,N_4908,N_4534);
and U5212 (N_5212,N_4885,N_4646);
xnor U5213 (N_5213,N_4969,N_4523);
nor U5214 (N_5214,N_4982,N_4687);
or U5215 (N_5215,N_4686,N_4898);
or U5216 (N_5216,N_4931,N_4576);
nor U5217 (N_5217,N_4573,N_4838);
xnor U5218 (N_5218,N_4659,N_4927);
nand U5219 (N_5219,N_4629,N_4655);
or U5220 (N_5220,N_4566,N_4999);
xnor U5221 (N_5221,N_4910,N_4897);
nand U5222 (N_5222,N_4508,N_4976);
nor U5223 (N_5223,N_4731,N_4553);
nor U5224 (N_5224,N_4669,N_4944);
xnor U5225 (N_5225,N_4734,N_4767);
and U5226 (N_5226,N_4582,N_4589);
or U5227 (N_5227,N_4934,N_4789);
nand U5228 (N_5228,N_4739,N_4936);
or U5229 (N_5229,N_4947,N_4608);
and U5230 (N_5230,N_4953,N_4712);
nor U5231 (N_5231,N_4879,N_4967);
nand U5232 (N_5232,N_4641,N_4678);
and U5233 (N_5233,N_4571,N_4628);
and U5234 (N_5234,N_4601,N_4703);
xnor U5235 (N_5235,N_4595,N_4996);
nor U5236 (N_5236,N_4920,N_4513);
or U5237 (N_5237,N_4966,N_4890);
nand U5238 (N_5238,N_4700,N_4546);
nor U5239 (N_5239,N_4613,N_4806);
xnor U5240 (N_5240,N_4692,N_4820);
and U5241 (N_5241,N_4533,N_4858);
nand U5242 (N_5242,N_4502,N_4529);
and U5243 (N_5243,N_4567,N_4752);
and U5244 (N_5244,N_4768,N_4917);
or U5245 (N_5245,N_4786,N_4907);
or U5246 (N_5246,N_4844,N_4528);
nor U5247 (N_5247,N_4914,N_4896);
and U5248 (N_5248,N_4859,N_4564);
nor U5249 (N_5249,N_4614,N_4577);
and U5250 (N_5250,N_4821,N_4939);
nand U5251 (N_5251,N_4642,N_4932);
nand U5252 (N_5252,N_4839,N_4719);
and U5253 (N_5253,N_4828,N_4871);
or U5254 (N_5254,N_4642,N_4653);
or U5255 (N_5255,N_4795,N_4947);
xor U5256 (N_5256,N_4908,N_4603);
or U5257 (N_5257,N_4559,N_4634);
or U5258 (N_5258,N_4678,N_4836);
nand U5259 (N_5259,N_4622,N_4914);
nor U5260 (N_5260,N_4735,N_4854);
and U5261 (N_5261,N_4595,N_4881);
nand U5262 (N_5262,N_4789,N_4801);
xor U5263 (N_5263,N_4747,N_4961);
and U5264 (N_5264,N_4929,N_4966);
xor U5265 (N_5265,N_4527,N_4985);
or U5266 (N_5266,N_4730,N_4979);
nor U5267 (N_5267,N_4648,N_4740);
nor U5268 (N_5268,N_4509,N_4616);
nor U5269 (N_5269,N_4841,N_4630);
nor U5270 (N_5270,N_4747,N_4797);
and U5271 (N_5271,N_4647,N_4535);
xor U5272 (N_5272,N_4976,N_4644);
nand U5273 (N_5273,N_4591,N_4994);
and U5274 (N_5274,N_4904,N_4573);
xor U5275 (N_5275,N_4938,N_4785);
and U5276 (N_5276,N_4959,N_4829);
nand U5277 (N_5277,N_4887,N_4636);
and U5278 (N_5278,N_4673,N_4530);
xor U5279 (N_5279,N_4845,N_4825);
nor U5280 (N_5280,N_4731,N_4512);
nor U5281 (N_5281,N_4870,N_4865);
nand U5282 (N_5282,N_4730,N_4709);
nor U5283 (N_5283,N_4764,N_4644);
nand U5284 (N_5284,N_4621,N_4647);
xor U5285 (N_5285,N_4675,N_4659);
xnor U5286 (N_5286,N_4697,N_4703);
nor U5287 (N_5287,N_4997,N_4870);
or U5288 (N_5288,N_4926,N_4640);
xnor U5289 (N_5289,N_4996,N_4511);
and U5290 (N_5290,N_4568,N_4771);
xor U5291 (N_5291,N_4791,N_4536);
nand U5292 (N_5292,N_4896,N_4681);
nor U5293 (N_5293,N_4546,N_4867);
or U5294 (N_5294,N_4637,N_4777);
nor U5295 (N_5295,N_4507,N_4847);
and U5296 (N_5296,N_4533,N_4887);
or U5297 (N_5297,N_4730,N_4803);
or U5298 (N_5298,N_4523,N_4549);
nand U5299 (N_5299,N_4952,N_4805);
nand U5300 (N_5300,N_4949,N_4968);
xor U5301 (N_5301,N_4535,N_4872);
xor U5302 (N_5302,N_4503,N_4942);
nor U5303 (N_5303,N_4999,N_4633);
and U5304 (N_5304,N_4826,N_4970);
nand U5305 (N_5305,N_4802,N_4934);
nor U5306 (N_5306,N_4659,N_4565);
or U5307 (N_5307,N_4616,N_4831);
nor U5308 (N_5308,N_4758,N_4582);
nor U5309 (N_5309,N_4709,N_4785);
nand U5310 (N_5310,N_4619,N_4799);
nor U5311 (N_5311,N_4595,N_4876);
xor U5312 (N_5312,N_4655,N_4926);
nor U5313 (N_5313,N_4697,N_4755);
xor U5314 (N_5314,N_4965,N_4677);
nand U5315 (N_5315,N_4694,N_4963);
nand U5316 (N_5316,N_4544,N_4668);
nand U5317 (N_5317,N_4886,N_4959);
nor U5318 (N_5318,N_4777,N_4882);
nand U5319 (N_5319,N_4881,N_4521);
nand U5320 (N_5320,N_4656,N_4936);
and U5321 (N_5321,N_4687,N_4641);
nor U5322 (N_5322,N_4802,N_4861);
and U5323 (N_5323,N_4883,N_4586);
xnor U5324 (N_5324,N_4899,N_4771);
nor U5325 (N_5325,N_4861,N_4682);
nand U5326 (N_5326,N_4735,N_4762);
nor U5327 (N_5327,N_4940,N_4779);
nor U5328 (N_5328,N_4500,N_4731);
nand U5329 (N_5329,N_4723,N_4511);
or U5330 (N_5330,N_4881,N_4923);
nand U5331 (N_5331,N_4659,N_4763);
or U5332 (N_5332,N_4780,N_4535);
or U5333 (N_5333,N_4987,N_4680);
or U5334 (N_5334,N_4554,N_4997);
xnor U5335 (N_5335,N_4503,N_4633);
nand U5336 (N_5336,N_4680,N_4670);
and U5337 (N_5337,N_4777,N_4914);
nor U5338 (N_5338,N_4839,N_4718);
nand U5339 (N_5339,N_4519,N_4537);
nand U5340 (N_5340,N_4850,N_4995);
or U5341 (N_5341,N_4989,N_4808);
nor U5342 (N_5342,N_4662,N_4881);
and U5343 (N_5343,N_4566,N_4935);
and U5344 (N_5344,N_4737,N_4619);
and U5345 (N_5345,N_4928,N_4958);
nand U5346 (N_5346,N_4576,N_4898);
or U5347 (N_5347,N_4744,N_4638);
nand U5348 (N_5348,N_4565,N_4765);
or U5349 (N_5349,N_4679,N_4515);
and U5350 (N_5350,N_4939,N_4624);
xnor U5351 (N_5351,N_4845,N_4896);
or U5352 (N_5352,N_4913,N_4535);
nor U5353 (N_5353,N_4603,N_4858);
nand U5354 (N_5354,N_4634,N_4852);
or U5355 (N_5355,N_4840,N_4866);
xnor U5356 (N_5356,N_4946,N_4731);
nor U5357 (N_5357,N_4927,N_4712);
and U5358 (N_5358,N_4670,N_4823);
or U5359 (N_5359,N_4544,N_4905);
nand U5360 (N_5360,N_4512,N_4525);
nor U5361 (N_5361,N_4692,N_4810);
and U5362 (N_5362,N_4831,N_4578);
nand U5363 (N_5363,N_4580,N_4854);
or U5364 (N_5364,N_4697,N_4930);
or U5365 (N_5365,N_4946,N_4656);
nor U5366 (N_5366,N_4725,N_4722);
nand U5367 (N_5367,N_4660,N_4982);
nor U5368 (N_5368,N_4818,N_4690);
or U5369 (N_5369,N_4617,N_4531);
or U5370 (N_5370,N_4893,N_4991);
nand U5371 (N_5371,N_4662,N_4639);
or U5372 (N_5372,N_4704,N_4524);
xor U5373 (N_5373,N_4918,N_4506);
xnor U5374 (N_5374,N_4955,N_4603);
nand U5375 (N_5375,N_4588,N_4616);
and U5376 (N_5376,N_4944,N_4686);
xor U5377 (N_5377,N_4982,N_4680);
nand U5378 (N_5378,N_4504,N_4928);
or U5379 (N_5379,N_4904,N_4691);
and U5380 (N_5380,N_4927,N_4851);
or U5381 (N_5381,N_4897,N_4919);
nor U5382 (N_5382,N_4713,N_4824);
or U5383 (N_5383,N_4638,N_4646);
xor U5384 (N_5384,N_4835,N_4655);
xor U5385 (N_5385,N_4509,N_4655);
or U5386 (N_5386,N_4958,N_4569);
or U5387 (N_5387,N_4735,N_4745);
nand U5388 (N_5388,N_4594,N_4777);
or U5389 (N_5389,N_4725,N_4541);
xor U5390 (N_5390,N_4674,N_4728);
and U5391 (N_5391,N_4865,N_4540);
xor U5392 (N_5392,N_4982,N_4565);
nor U5393 (N_5393,N_4889,N_4519);
nor U5394 (N_5394,N_4575,N_4623);
xnor U5395 (N_5395,N_4938,N_4802);
nand U5396 (N_5396,N_4630,N_4942);
or U5397 (N_5397,N_4563,N_4680);
and U5398 (N_5398,N_4935,N_4574);
xor U5399 (N_5399,N_4627,N_4586);
xor U5400 (N_5400,N_4680,N_4923);
nor U5401 (N_5401,N_4812,N_4988);
nor U5402 (N_5402,N_4508,N_4703);
xor U5403 (N_5403,N_4526,N_4585);
or U5404 (N_5404,N_4741,N_4761);
and U5405 (N_5405,N_4808,N_4867);
and U5406 (N_5406,N_4588,N_4842);
nor U5407 (N_5407,N_4914,N_4508);
or U5408 (N_5408,N_4648,N_4690);
and U5409 (N_5409,N_4766,N_4708);
xnor U5410 (N_5410,N_4572,N_4807);
and U5411 (N_5411,N_4537,N_4804);
or U5412 (N_5412,N_4574,N_4600);
xor U5413 (N_5413,N_4609,N_4598);
nor U5414 (N_5414,N_4690,N_4778);
nor U5415 (N_5415,N_4607,N_4753);
or U5416 (N_5416,N_4597,N_4516);
nand U5417 (N_5417,N_4660,N_4784);
xnor U5418 (N_5418,N_4717,N_4931);
or U5419 (N_5419,N_4644,N_4505);
nand U5420 (N_5420,N_4831,N_4585);
xnor U5421 (N_5421,N_4730,N_4992);
nand U5422 (N_5422,N_4534,N_4544);
nor U5423 (N_5423,N_4862,N_4712);
xor U5424 (N_5424,N_4803,N_4509);
or U5425 (N_5425,N_4651,N_4522);
and U5426 (N_5426,N_4728,N_4969);
nor U5427 (N_5427,N_4821,N_4811);
and U5428 (N_5428,N_4788,N_4972);
and U5429 (N_5429,N_4762,N_4569);
nor U5430 (N_5430,N_4669,N_4828);
nor U5431 (N_5431,N_4726,N_4619);
xor U5432 (N_5432,N_4715,N_4988);
nand U5433 (N_5433,N_4663,N_4722);
and U5434 (N_5434,N_4851,N_4537);
or U5435 (N_5435,N_4746,N_4782);
nor U5436 (N_5436,N_4856,N_4750);
nand U5437 (N_5437,N_4745,N_4684);
and U5438 (N_5438,N_4590,N_4582);
or U5439 (N_5439,N_4964,N_4613);
nor U5440 (N_5440,N_4850,N_4569);
xnor U5441 (N_5441,N_4521,N_4908);
nand U5442 (N_5442,N_4982,N_4856);
or U5443 (N_5443,N_4585,N_4506);
and U5444 (N_5444,N_4714,N_4981);
or U5445 (N_5445,N_4639,N_4894);
xnor U5446 (N_5446,N_4657,N_4588);
nor U5447 (N_5447,N_4932,N_4934);
nor U5448 (N_5448,N_4881,N_4887);
nand U5449 (N_5449,N_4621,N_4546);
and U5450 (N_5450,N_4888,N_4805);
nand U5451 (N_5451,N_4618,N_4647);
xor U5452 (N_5452,N_4873,N_4607);
and U5453 (N_5453,N_4923,N_4769);
and U5454 (N_5454,N_4659,N_4667);
xnor U5455 (N_5455,N_4887,N_4627);
or U5456 (N_5456,N_4527,N_4901);
or U5457 (N_5457,N_4632,N_4541);
nor U5458 (N_5458,N_4641,N_4565);
nand U5459 (N_5459,N_4709,N_4682);
xnor U5460 (N_5460,N_4503,N_4690);
and U5461 (N_5461,N_4975,N_4555);
or U5462 (N_5462,N_4515,N_4898);
nor U5463 (N_5463,N_4538,N_4844);
nand U5464 (N_5464,N_4942,N_4833);
xnor U5465 (N_5465,N_4808,N_4842);
and U5466 (N_5466,N_4506,N_4945);
xor U5467 (N_5467,N_4797,N_4927);
and U5468 (N_5468,N_4940,N_4686);
xor U5469 (N_5469,N_4897,N_4887);
xnor U5470 (N_5470,N_4523,N_4620);
and U5471 (N_5471,N_4861,N_4574);
or U5472 (N_5472,N_4562,N_4867);
nand U5473 (N_5473,N_4991,N_4974);
nor U5474 (N_5474,N_4951,N_4771);
and U5475 (N_5475,N_4838,N_4615);
or U5476 (N_5476,N_4908,N_4682);
nor U5477 (N_5477,N_4676,N_4949);
xor U5478 (N_5478,N_4743,N_4920);
xor U5479 (N_5479,N_4808,N_4667);
nor U5480 (N_5480,N_4904,N_4633);
or U5481 (N_5481,N_4959,N_4973);
nand U5482 (N_5482,N_4713,N_4737);
or U5483 (N_5483,N_4582,N_4967);
or U5484 (N_5484,N_4648,N_4506);
and U5485 (N_5485,N_4778,N_4813);
or U5486 (N_5486,N_4946,N_4882);
nand U5487 (N_5487,N_4930,N_4668);
nor U5488 (N_5488,N_4971,N_4932);
xnor U5489 (N_5489,N_4895,N_4723);
nand U5490 (N_5490,N_4931,N_4853);
and U5491 (N_5491,N_4969,N_4642);
xor U5492 (N_5492,N_4735,N_4965);
xnor U5493 (N_5493,N_4909,N_4755);
nor U5494 (N_5494,N_4798,N_4709);
or U5495 (N_5495,N_4796,N_4506);
nand U5496 (N_5496,N_4604,N_4710);
xnor U5497 (N_5497,N_4954,N_4577);
nor U5498 (N_5498,N_4602,N_4664);
nand U5499 (N_5499,N_4529,N_4638);
or U5500 (N_5500,N_5219,N_5270);
xor U5501 (N_5501,N_5413,N_5263);
or U5502 (N_5502,N_5124,N_5029);
xor U5503 (N_5503,N_5387,N_5330);
xnor U5504 (N_5504,N_5483,N_5318);
or U5505 (N_5505,N_5246,N_5295);
nand U5506 (N_5506,N_5205,N_5097);
xor U5507 (N_5507,N_5333,N_5166);
nor U5508 (N_5508,N_5232,N_5481);
or U5509 (N_5509,N_5396,N_5137);
nor U5510 (N_5510,N_5085,N_5266);
and U5511 (N_5511,N_5123,N_5288);
nand U5512 (N_5512,N_5499,N_5426);
and U5513 (N_5513,N_5168,N_5464);
and U5514 (N_5514,N_5132,N_5022);
xnor U5515 (N_5515,N_5379,N_5080);
or U5516 (N_5516,N_5460,N_5144);
nand U5517 (N_5517,N_5250,N_5408);
nand U5518 (N_5518,N_5202,N_5222);
and U5519 (N_5519,N_5013,N_5487);
and U5520 (N_5520,N_5200,N_5196);
or U5521 (N_5521,N_5345,N_5173);
nand U5522 (N_5522,N_5390,N_5319);
and U5523 (N_5523,N_5368,N_5428);
nand U5524 (N_5524,N_5462,N_5053);
nor U5525 (N_5525,N_5399,N_5087);
xnor U5526 (N_5526,N_5444,N_5175);
nor U5527 (N_5527,N_5465,N_5164);
nand U5528 (N_5528,N_5286,N_5057);
or U5529 (N_5529,N_5498,N_5241);
nand U5530 (N_5530,N_5195,N_5229);
nand U5531 (N_5531,N_5279,N_5313);
nor U5532 (N_5532,N_5290,N_5328);
xor U5533 (N_5533,N_5445,N_5093);
xor U5534 (N_5534,N_5435,N_5287);
and U5535 (N_5535,N_5441,N_5404);
xnor U5536 (N_5536,N_5277,N_5334);
nand U5537 (N_5537,N_5478,N_5296);
or U5538 (N_5538,N_5079,N_5257);
or U5539 (N_5539,N_5412,N_5410);
and U5540 (N_5540,N_5358,N_5044);
nor U5541 (N_5541,N_5008,N_5204);
or U5542 (N_5542,N_5361,N_5094);
and U5543 (N_5543,N_5249,N_5273);
nor U5544 (N_5544,N_5349,N_5304);
or U5545 (N_5545,N_5431,N_5443);
nor U5546 (N_5546,N_5032,N_5389);
and U5547 (N_5547,N_5161,N_5235);
or U5548 (N_5548,N_5129,N_5398);
xnor U5549 (N_5549,N_5457,N_5109);
nor U5550 (N_5550,N_5225,N_5212);
or U5551 (N_5551,N_5206,N_5010);
nand U5552 (N_5552,N_5242,N_5074);
and U5553 (N_5553,N_5201,N_5363);
or U5554 (N_5554,N_5076,N_5036);
xnor U5555 (N_5555,N_5397,N_5141);
nand U5556 (N_5556,N_5006,N_5118);
and U5557 (N_5557,N_5350,N_5121);
nor U5558 (N_5558,N_5267,N_5377);
and U5559 (N_5559,N_5421,N_5468);
or U5560 (N_5560,N_5309,N_5488);
and U5561 (N_5561,N_5223,N_5226);
nor U5562 (N_5562,N_5128,N_5491);
xnor U5563 (N_5563,N_5433,N_5068);
or U5564 (N_5564,N_5278,N_5332);
and U5565 (N_5565,N_5108,N_5459);
nor U5566 (N_5566,N_5240,N_5451);
and U5567 (N_5567,N_5213,N_5327);
nor U5568 (N_5568,N_5471,N_5024);
nor U5569 (N_5569,N_5385,N_5089);
or U5570 (N_5570,N_5496,N_5414);
nor U5571 (N_5571,N_5209,N_5180);
nand U5572 (N_5572,N_5417,N_5045);
nor U5573 (N_5573,N_5392,N_5001);
xor U5574 (N_5574,N_5217,N_5055);
nand U5575 (N_5575,N_5185,N_5194);
nor U5576 (N_5576,N_5075,N_5030);
and U5577 (N_5577,N_5113,N_5293);
nor U5578 (N_5578,N_5364,N_5071);
and U5579 (N_5579,N_5382,N_5251);
xor U5580 (N_5580,N_5002,N_5064);
nand U5581 (N_5581,N_5122,N_5082);
or U5582 (N_5582,N_5494,N_5455);
and U5583 (N_5583,N_5103,N_5186);
or U5584 (N_5584,N_5434,N_5305);
xor U5585 (N_5585,N_5126,N_5157);
nor U5586 (N_5586,N_5009,N_5004);
nor U5587 (N_5587,N_5051,N_5424);
nor U5588 (N_5588,N_5106,N_5237);
and U5589 (N_5589,N_5291,N_5130);
nand U5590 (N_5590,N_5321,N_5395);
or U5591 (N_5591,N_5475,N_5178);
xor U5592 (N_5592,N_5493,N_5102);
nand U5593 (N_5593,N_5221,N_5376);
nor U5594 (N_5594,N_5325,N_5125);
nand U5595 (N_5595,N_5469,N_5153);
nor U5596 (N_5596,N_5170,N_5127);
and U5597 (N_5597,N_5429,N_5189);
nor U5598 (N_5598,N_5381,N_5301);
nor U5599 (N_5599,N_5294,N_5422);
nand U5600 (N_5600,N_5234,N_5256);
and U5601 (N_5601,N_5098,N_5084);
or U5602 (N_5602,N_5210,N_5190);
and U5603 (N_5603,N_5322,N_5149);
and U5604 (N_5604,N_5188,N_5155);
nand U5605 (N_5605,N_5037,N_5070);
xnor U5606 (N_5606,N_5131,N_5061);
and U5607 (N_5607,N_5484,N_5261);
xnor U5608 (N_5608,N_5003,N_5238);
nor U5609 (N_5609,N_5370,N_5409);
nor U5610 (N_5610,N_5114,N_5252);
and U5611 (N_5611,N_5169,N_5477);
nor U5612 (N_5612,N_5380,N_5104);
xor U5613 (N_5613,N_5351,N_5069);
nand U5614 (N_5614,N_5083,N_5394);
xnor U5615 (N_5615,N_5049,N_5386);
xor U5616 (N_5616,N_5224,N_5208);
or U5617 (N_5617,N_5298,N_5174);
nand U5618 (N_5618,N_5449,N_5181);
or U5619 (N_5619,N_5017,N_5437);
or U5620 (N_5620,N_5147,N_5356);
and U5621 (N_5621,N_5337,N_5306);
nor U5622 (N_5622,N_5480,N_5450);
or U5623 (N_5623,N_5310,N_5214);
nor U5624 (N_5624,N_5066,N_5043);
xnor U5625 (N_5625,N_5405,N_5336);
xnor U5626 (N_5626,N_5362,N_5492);
xor U5627 (N_5627,N_5470,N_5021);
or U5628 (N_5628,N_5474,N_5182);
or U5629 (N_5629,N_5497,N_5312);
nor U5630 (N_5630,N_5211,N_5067);
nor U5631 (N_5631,N_5039,N_5150);
nand U5632 (N_5632,N_5138,N_5308);
nor U5633 (N_5633,N_5472,N_5145);
nand U5634 (N_5634,N_5183,N_5366);
and U5635 (N_5635,N_5136,N_5353);
or U5636 (N_5636,N_5116,N_5231);
nor U5637 (N_5637,N_5485,N_5090);
nand U5638 (N_5638,N_5236,N_5438);
or U5639 (N_5639,N_5193,N_5340);
nor U5640 (N_5640,N_5060,N_5315);
or U5641 (N_5641,N_5134,N_5281);
nand U5642 (N_5642,N_5244,N_5323);
nand U5643 (N_5643,N_5447,N_5099);
and U5644 (N_5644,N_5052,N_5119);
xor U5645 (N_5645,N_5248,N_5040);
nor U5646 (N_5646,N_5111,N_5343);
and U5647 (N_5647,N_5063,N_5365);
nand U5648 (N_5648,N_5357,N_5262);
xor U5649 (N_5649,N_5371,N_5299);
or U5650 (N_5650,N_5314,N_5275);
and U5651 (N_5651,N_5341,N_5375);
nor U5652 (N_5652,N_5007,N_5177);
and U5653 (N_5653,N_5442,N_5253);
or U5654 (N_5654,N_5282,N_5197);
nor U5655 (N_5655,N_5276,N_5054);
xor U5656 (N_5656,N_5415,N_5284);
or U5657 (N_5657,N_5359,N_5454);
or U5658 (N_5658,N_5378,N_5160);
nor U5659 (N_5659,N_5112,N_5207);
xnor U5660 (N_5660,N_5479,N_5014);
nor U5661 (N_5661,N_5420,N_5269);
nand U5662 (N_5662,N_5335,N_5388);
nand U5663 (N_5663,N_5259,N_5425);
nand U5664 (N_5664,N_5272,N_5401);
or U5665 (N_5665,N_5078,N_5384);
or U5666 (N_5666,N_5107,N_5203);
xnor U5667 (N_5667,N_5355,N_5360);
nand U5668 (N_5668,N_5383,N_5430);
and U5669 (N_5669,N_5041,N_5215);
nand U5670 (N_5670,N_5117,N_5011);
or U5671 (N_5671,N_5391,N_5096);
xor U5672 (N_5672,N_5440,N_5148);
nand U5673 (N_5673,N_5452,N_5218);
or U5674 (N_5674,N_5059,N_5254);
and U5675 (N_5675,N_5473,N_5020);
nand U5676 (N_5676,N_5026,N_5031);
or U5677 (N_5677,N_5342,N_5458);
or U5678 (N_5678,N_5151,N_5176);
or U5679 (N_5679,N_5005,N_5135);
and U5680 (N_5680,N_5264,N_5495);
or U5681 (N_5681,N_5320,N_5019);
nand U5682 (N_5682,N_5110,N_5033);
xnor U5683 (N_5683,N_5105,N_5165);
and U5684 (N_5684,N_5139,N_5035);
nand U5685 (N_5685,N_5461,N_5367);
or U5686 (N_5686,N_5289,N_5283);
xor U5687 (N_5687,N_5423,N_5255);
and U5688 (N_5688,N_5016,N_5432);
nand U5689 (N_5689,N_5239,N_5427);
xnor U5690 (N_5690,N_5402,N_5352);
xnor U5691 (N_5691,N_5140,N_5056);
and U5692 (N_5692,N_5091,N_5418);
and U5693 (N_5693,N_5227,N_5403);
or U5694 (N_5694,N_5354,N_5324);
xor U5695 (N_5695,N_5191,N_5326);
nor U5696 (N_5696,N_5400,N_5048);
and U5697 (N_5697,N_5015,N_5271);
xnor U5698 (N_5698,N_5265,N_5303);
nand U5699 (N_5699,N_5292,N_5120);
nor U5700 (N_5700,N_5448,N_5167);
or U5701 (N_5701,N_5439,N_5042);
nand U5702 (N_5702,N_5339,N_5274);
nand U5703 (N_5703,N_5344,N_5369);
and U5704 (N_5704,N_5489,N_5453);
or U5705 (N_5705,N_5058,N_5000);
nor U5706 (N_5706,N_5065,N_5163);
or U5707 (N_5707,N_5088,N_5316);
nor U5708 (N_5708,N_5374,N_5486);
xor U5709 (N_5709,N_5233,N_5228);
nand U5710 (N_5710,N_5086,N_5338);
xnor U5711 (N_5711,N_5025,N_5373);
nor U5712 (N_5712,N_5490,N_5172);
nor U5713 (N_5713,N_5268,N_5050);
nand U5714 (N_5714,N_5192,N_5436);
or U5715 (N_5715,N_5028,N_5467);
nor U5716 (N_5716,N_5179,N_5280);
or U5717 (N_5717,N_5154,N_5411);
or U5718 (N_5718,N_5101,N_5419);
xor U5719 (N_5719,N_5393,N_5482);
nand U5720 (N_5720,N_5152,N_5311);
or U5721 (N_5721,N_5216,N_5372);
nand U5722 (N_5722,N_5142,N_5047);
nor U5723 (N_5723,N_5199,N_5346);
nor U5724 (N_5724,N_5143,N_5156);
xnor U5725 (N_5725,N_5034,N_5300);
and U5726 (N_5726,N_5092,N_5407);
and U5727 (N_5727,N_5158,N_5115);
nand U5728 (N_5728,N_5258,N_5243);
nand U5729 (N_5729,N_5187,N_5077);
nor U5730 (N_5730,N_5162,N_5245);
and U5731 (N_5731,N_5302,N_5466);
and U5732 (N_5732,N_5446,N_5133);
nand U5733 (N_5733,N_5027,N_5100);
nor U5734 (N_5734,N_5171,N_5247);
xnor U5735 (N_5735,N_5285,N_5347);
xor U5736 (N_5736,N_5146,N_5406);
nand U5737 (N_5737,N_5159,N_5348);
nor U5738 (N_5738,N_5329,N_5230);
or U5739 (N_5739,N_5081,N_5198);
or U5740 (N_5740,N_5012,N_5463);
and U5741 (N_5741,N_5023,N_5297);
nand U5742 (N_5742,N_5062,N_5046);
xnor U5743 (N_5743,N_5038,N_5184);
and U5744 (N_5744,N_5331,N_5307);
or U5745 (N_5745,N_5416,N_5073);
nand U5746 (N_5746,N_5260,N_5220);
and U5747 (N_5747,N_5095,N_5317);
xor U5748 (N_5748,N_5072,N_5018);
or U5749 (N_5749,N_5476,N_5456);
and U5750 (N_5750,N_5094,N_5494);
xor U5751 (N_5751,N_5474,N_5230);
nor U5752 (N_5752,N_5210,N_5134);
nand U5753 (N_5753,N_5295,N_5167);
nor U5754 (N_5754,N_5347,N_5363);
nor U5755 (N_5755,N_5426,N_5218);
nand U5756 (N_5756,N_5160,N_5218);
or U5757 (N_5757,N_5371,N_5390);
and U5758 (N_5758,N_5118,N_5346);
nor U5759 (N_5759,N_5278,N_5386);
and U5760 (N_5760,N_5253,N_5414);
or U5761 (N_5761,N_5481,N_5159);
or U5762 (N_5762,N_5333,N_5305);
and U5763 (N_5763,N_5050,N_5253);
or U5764 (N_5764,N_5423,N_5007);
xor U5765 (N_5765,N_5363,N_5253);
xnor U5766 (N_5766,N_5216,N_5205);
and U5767 (N_5767,N_5250,N_5237);
nand U5768 (N_5768,N_5395,N_5089);
nor U5769 (N_5769,N_5039,N_5063);
and U5770 (N_5770,N_5101,N_5004);
xor U5771 (N_5771,N_5396,N_5213);
nor U5772 (N_5772,N_5322,N_5136);
and U5773 (N_5773,N_5411,N_5248);
xor U5774 (N_5774,N_5323,N_5264);
nand U5775 (N_5775,N_5206,N_5095);
or U5776 (N_5776,N_5133,N_5313);
nand U5777 (N_5777,N_5097,N_5352);
or U5778 (N_5778,N_5048,N_5047);
xnor U5779 (N_5779,N_5323,N_5457);
nand U5780 (N_5780,N_5432,N_5495);
and U5781 (N_5781,N_5403,N_5096);
or U5782 (N_5782,N_5497,N_5328);
xnor U5783 (N_5783,N_5332,N_5172);
or U5784 (N_5784,N_5326,N_5260);
and U5785 (N_5785,N_5337,N_5050);
or U5786 (N_5786,N_5291,N_5258);
or U5787 (N_5787,N_5122,N_5197);
and U5788 (N_5788,N_5052,N_5087);
xor U5789 (N_5789,N_5330,N_5175);
xnor U5790 (N_5790,N_5105,N_5417);
xnor U5791 (N_5791,N_5289,N_5431);
nor U5792 (N_5792,N_5161,N_5011);
nand U5793 (N_5793,N_5030,N_5469);
and U5794 (N_5794,N_5481,N_5056);
or U5795 (N_5795,N_5236,N_5461);
nand U5796 (N_5796,N_5251,N_5202);
xor U5797 (N_5797,N_5205,N_5035);
xor U5798 (N_5798,N_5265,N_5308);
nand U5799 (N_5799,N_5049,N_5094);
nor U5800 (N_5800,N_5473,N_5127);
xnor U5801 (N_5801,N_5419,N_5167);
nand U5802 (N_5802,N_5441,N_5357);
and U5803 (N_5803,N_5384,N_5188);
nand U5804 (N_5804,N_5120,N_5472);
xnor U5805 (N_5805,N_5478,N_5463);
nor U5806 (N_5806,N_5463,N_5003);
or U5807 (N_5807,N_5172,N_5390);
nor U5808 (N_5808,N_5423,N_5066);
nand U5809 (N_5809,N_5365,N_5467);
nand U5810 (N_5810,N_5428,N_5267);
and U5811 (N_5811,N_5434,N_5447);
nor U5812 (N_5812,N_5199,N_5469);
or U5813 (N_5813,N_5216,N_5156);
nor U5814 (N_5814,N_5464,N_5228);
and U5815 (N_5815,N_5106,N_5356);
nand U5816 (N_5816,N_5403,N_5205);
xor U5817 (N_5817,N_5378,N_5357);
nand U5818 (N_5818,N_5326,N_5160);
or U5819 (N_5819,N_5167,N_5290);
nand U5820 (N_5820,N_5206,N_5128);
nor U5821 (N_5821,N_5315,N_5161);
nand U5822 (N_5822,N_5290,N_5326);
xnor U5823 (N_5823,N_5435,N_5209);
xnor U5824 (N_5824,N_5490,N_5045);
or U5825 (N_5825,N_5185,N_5305);
or U5826 (N_5826,N_5177,N_5038);
xor U5827 (N_5827,N_5053,N_5300);
nand U5828 (N_5828,N_5172,N_5413);
and U5829 (N_5829,N_5432,N_5174);
xnor U5830 (N_5830,N_5083,N_5375);
nor U5831 (N_5831,N_5208,N_5198);
or U5832 (N_5832,N_5294,N_5494);
nand U5833 (N_5833,N_5098,N_5353);
xnor U5834 (N_5834,N_5088,N_5301);
nor U5835 (N_5835,N_5401,N_5365);
or U5836 (N_5836,N_5318,N_5269);
xnor U5837 (N_5837,N_5351,N_5425);
nand U5838 (N_5838,N_5426,N_5292);
nor U5839 (N_5839,N_5132,N_5206);
nand U5840 (N_5840,N_5124,N_5221);
or U5841 (N_5841,N_5167,N_5128);
or U5842 (N_5842,N_5042,N_5306);
and U5843 (N_5843,N_5492,N_5301);
nor U5844 (N_5844,N_5201,N_5223);
nor U5845 (N_5845,N_5472,N_5403);
xor U5846 (N_5846,N_5126,N_5145);
or U5847 (N_5847,N_5133,N_5123);
nor U5848 (N_5848,N_5223,N_5066);
xnor U5849 (N_5849,N_5245,N_5122);
or U5850 (N_5850,N_5335,N_5059);
or U5851 (N_5851,N_5183,N_5368);
nor U5852 (N_5852,N_5119,N_5342);
nor U5853 (N_5853,N_5009,N_5192);
nand U5854 (N_5854,N_5057,N_5130);
nor U5855 (N_5855,N_5472,N_5212);
and U5856 (N_5856,N_5219,N_5481);
nand U5857 (N_5857,N_5133,N_5221);
xnor U5858 (N_5858,N_5259,N_5365);
nand U5859 (N_5859,N_5447,N_5239);
nor U5860 (N_5860,N_5484,N_5491);
nand U5861 (N_5861,N_5259,N_5094);
and U5862 (N_5862,N_5127,N_5209);
nand U5863 (N_5863,N_5406,N_5093);
and U5864 (N_5864,N_5218,N_5400);
nand U5865 (N_5865,N_5015,N_5480);
or U5866 (N_5866,N_5001,N_5446);
and U5867 (N_5867,N_5191,N_5498);
xnor U5868 (N_5868,N_5214,N_5065);
and U5869 (N_5869,N_5350,N_5276);
nor U5870 (N_5870,N_5163,N_5354);
nor U5871 (N_5871,N_5008,N_5163);
nand U5872 (N_5872,N_5077,N_5109);
or U5873 (N_5873,N_5382,N_5440);
nand U5874 (N_5874,N_5056,N_5049);
nor U5875 (N_5875,N_5449,N_5184);
nor U5876 (N_5876,N_5420,N_5245);
nand U5877 (N_5877,N_5426,N_5202);
and U5878 (N_5878,N_5005,N_5427);
nand U5879 (N_5879,N_5147,N_5323);
or U5880 (N_5880,N_5344,N_5495);
or U5881 (N_5881,N_5413,N_5307);
xor U5882 (N_5882,N_5293,N_5462);
and U5883 (N_5883,N_5312,N_5206);
nand U5884 (N_5884,N_5122,N_5370);
or U5885 (N_5885,N_5351,N_5412);
nand U5886 (N_5886,N_5362,N_5474);
or U5887 (N_5887,N_5115,N_5253);
xnor U5888 (N_5888,N_5440,N_5454);
nand U5889 (N_5889,N_5070,N_5158);
nand U5890 (N_5890,N_5391,N_5222);
and U5891 (N_5891,N_5123,N_5327);
and U5892 (N_5892,N_5032,N_5287);
nor U5893 (N_5893,N_5120,N_5478);
nor U5894 (N_5894,N_5388,N_5154);
nand U5895 (N_5895,N_5259,N_5139);
nor U5896 (N_5896,N_5064,N_5082);
nand U5897 (N_5897,N_5179,N_5162);
xor U5898 (N_5898,N_5359,N_5461);
nor U5899 (N_5899,N_5203,N_5435);
nor U5900 (N_5900,N_5049,N_5015);
nand U5901 (N_5901,N_5413,N_5074);
or U5902 (N_5902,N_5269,N_5006);
and U5903 (N_5903,N_5014,N_5142);
and U5904 (N_5904,N_5312,N_5475);
or U5905 (N_5905,N_5309,N_5189);
and U5906 (N_5906,N_5294,N_5175);
and U5907 (N_5907,N_5365,N_5399);
or U5908 (N_5908,N_5382,N_5286);
or U5909 (N_5909,N_5369,N_5060);
nand U5910 (N_5910,N_5181,N_5240);
xor U5911 (N_5911,N_5029,N_5309);
nand U5912 (N_5912,N_5493,N_5094);
nor U5913 (N_5913,N_5132,N_5349);
and U5914 (N_5914,N_5372,N_5428);
or U5915 (N_5915,N_5098,N_5458);
and U5916 (N_5916,N_5221,N_5454);
xnor U5917 (N_5917,N_5031,N_5449);
nand U5918 (N_5918,N_5352,N_5035);
and U5919 (N_5919,N_5071,N_5445);
nand U5920 (N_5920,N_5327,N_5159);
xor U5921 (N_5921,N_5159,N_5482);
and U5922 (N_5922,N_5173,N_5251);
nor U5923 (N_5923,N_5402,N_5124);
xor U5924 (N_5924,N_5086,N_5487);
nor U5925 (N_5925,N_5084,N_5457);
nor U5926 (N_5926,N_5080,N_5138);
xnor U5927 (N_5927,N_5312,N_5374);
or U5928 (N_5928,N_5269,N_5250);
or U5929 (N_5929,N_5036,N_5145);
nor U5930 (N_5930,N_5176,N_5327);
xnor U5931 (N_5931,N_5459,N_5168);
xnor U5932 (N_5932,N_5056,N_5338);
xor U5933 (N_5933,N_5372,N_5170);
nor U5934 (N_5934,N_5363,N_5265);
nor U5935 (N_5935,N_5459,N_5262);
and U5936 (N_5936,N_5325,N_5047);
xnor U5937 (N_5937,N_5398,N_5397);
and U5938 (N_5938,N_5395,N_5131);
nand U5939 (N_5939,N_5457,N_5326);
nor U5940 (N_5940,N_5110,N_5218);
and U5941 (N_5941,N_5423,N_5409);
nor U5942 (N_5942,N_5080,N_5449);
or U5943 (N_5943,N_5201,N_5043);
nor U5944 (N_5944,N_5246,N_5488);
nand U5945 (N_5945,N_5491,N_5448);
and U5946 (N_5946,N_5106,N_5044);
xor U5947 (N_5947,N_5103,N_5302);
nand U5948 (N_5948,N_5078,N_5104);
and U5949 (N_5949,N_5026,N_5367);
nand U5950 (N_5950,N_5280,N_5101);
nand U5951 (N_5951,N_5331,N_5233);
or U5952 (N_5952,N_5472,N_5035);
and U5953 (N_5953,N_5398,N_5164);
or U5954 (N_5954,N_5021,N_5008);
or U5955 (N_5955,N_5277,N_5387);
xnor U5956 (N_5956,N_5419,N_5236);
or U5957 (N_5957,N_5195,N_5329);
nor U5958 (N_5958,N_5348,N_5306);
nand U5959 (N_5959,N_5064,N_5469);
or U5960 (N_5960,N_5466,N_5340);
nor U5961 (N_5961,N_5242,N_5035);
nand U5962 (N_5962,N_5184,N_5474);
xor U5963 (N_5963,N_5181,N_5075);
or U5964 (N_5964,N_5137,N_5164);
xnor U5965 (N_5965,N_5181,N_5177);
nand U5966 (N_5966,N_5498,N_5039);
and U5967 (N_5967,N_5470,N_5361);
nand U5968 (N_5968,N_5279,N_5250);
or U5969 (N_5969,N_5015,N_5205);
and U5970 (N_5970,N_5038,N_5391);
xnor U5971 (N_5971,N_5327,N_5491);
and U5972 (N_5972,N_5250,N_5448);
nor U5973 (N_5973,N_5269,N_5160);
or U5974 (N_5974,N_5200,N_5116);
nand U5975 (N_5975,N_5296,N_5291);
nor U5976 (N_5976,N_5059,N_5160);
nand U5977 (N_5977,N_5151,N_5028);
or U5978 (N_5978,N_5301,N_5491);
nor U5979 (N_5979,N_5342,N_5440);
nand U5980 (N_5980,N_5125,N_5014);
xor U5981 (N_5981,N_5351,N_5168);
or U5982 (N_5982,N_5073,N_5439);
or U5983 (N_5983,N_5308,N_5352);
and U5984 (N_5984,N_5231,N_5201);
nor U5985 (N_5985,N_5407,N_5491);
nand U5986 (N_5986,N_5371,N_5411);
nor U5987 (N_5987,N_5337,N_5079);
and U5988 (N_5988,N_5017,N_5273);
or U5989 (N_5989,N_5138,N_5162);
xnor U5990 (N_5990,N_5288,N_5157);
nand U5991 (N_5991,N_5379,N_5456);
nand U5992 (N_5992,N_5185,N_5375);
nor U5993 (N_5993,N_5255,N_5041);
or U5994 (N_5994,N_5032,N_5406);
or U5995 (N_5995,N_5462,N_5142);
nor U5996 (N_5996,N_5067,N_5327);
or U5997 (N_5997,N_5470,N_5308);
xor U5998 (N_5998,N_5108,N_5366);
and U5999 (N_5999,N_5396,N_5125);
xor U6000 (N_6000,N_5681,N_5795);
nor U6001 (N_6001,N_5987,N_5820);
nand U6002 (N_6002,N_5758,N_5660);
or U6003 (N_6003,N_5573,N_5624);
nor U6004 (N_6004,N_5603,N_5914);
xor U6005 (N_6005,N_5546,N_5583);
or U6006 (N_6006,N_5705,N_5727);
nor U6007 (N_6007,N_5604,N_5676);
or U6008 (N_6008,N_5719,N_5993);
nand U6009 (N_6009,N_5922,N_5895);
xor U6010 (N_6010,N_5958,N_5946);
and U6011 (N_6011,N_5668,N_5636);
xnor U6012 (N_6012,N_5571,N_5974);
nand U6013 (N_6013,N_5970,N_5582);
xnor U6014 (N_6014,N_5627,N_5834);
xor U6015 (N_6015,N_5770,N_5568);
nor U6016 (N_6016,N_5803,N_5728);
xnor U6017 (N_6017,N_5665,N_5606);
xnor U6018 (N_6018,N_5519,N_5680);
nand U6019 (N_6019,N_5733,N_5817);
nand U6020 (N_6020,N_5672,N_5923);
xor U6021 (N_6021,N_5677,N_5578);
nand U6022 (N_6022,N_5514,N_5642);
xnor U6023 (N_6023,N_5601,N_5917);
nor U6024 (N_6024,N_5701,N_5826);
nand U6025 (N_6025,N_5945,N_5543);
nand U6026 (N_6026,N_5520,N_5679);
nor U6027 (N_6027,N_5761,N_5745);
or U6028 (N_6028,N_5663,N_5581);
and U6029 (N_6029,N_5845,N_5882);
or U6030 (N_6030,N_5542,N_5830);
xnor U6031 (N_6031,N_5666,N_5975);
and U6032 (N_6032,N_5717,N_5539);
nand U6033 (N_6033,N_5551,N_5731);
xnor U6034 (N_6034,N_5777,N_5916);
and U6035 (N_6035,N_5708,N_5842);
and U6036 (N_6036,N_5599,N_5956);
or U6037 (N_6037,N_5775,N_5620);
xor U6038 (N_6038,N_5595,N_5545);
xor U6039 (N_6039,N_5819,N_5691);
nor U6040 (N_6040,N_5686,N_5739);
and U6041 (N_6041,N_5889,N_5871);
nand U6042 (N_6042,N_5779,N_5644);
and U6043 (N_6043,N_5645,N_5813);
nand U6044 (N_6044,N_5517,N_5983);
nand U6045 (N_6045,N_5751,N_5589);
or U6046 (N_6046,N_5857,N_5839);
xor U6047 (N_6047,N_5698,N_5920);
nand U6048 (N_6048,N_5629,N_5893);
nand U6049 (N_6049,N_5657,N_5593);
or U6050 (N_6050,N_5781,N_5936);
xnor U6051 (N_6051,N_5768,N_5626);
xnor U6052 (N_6052,N_5836,N_5506);
xnor U6053 (N_6053,N_5750,N_5843);
or U6054 (N_6054,N_5821,N_5904);
nand U6055 (N_6055,N_5855,N_5658);
nor U6056 (N_6056,N_5902,N_5726);
or U6057 (N_6057,N_5518,N_5961);
and U6058 (N_6058,N_5921,N_5748);
or U6059 (N_6059,N_5702,N_5858);
nand U6060 (N_6060,N_5872,N_5963);
nor U6061 (N_6061,N_5877,N_5793);
nor U6062 (N_6062,N_5553,N_5976);
nand U6063 (N_6063,N_5856,N_5554);
and U6064 (N_6064,N_5841,N_5513);
nor U6065 (N_6065,N_5764,N_5847);
xor U6066 (N_6066,N_5865,N_5704);
nor U6067 (N_6067,N_5787,N_5939);
xnor U6068 (N_6068,N_5564,N_5639);
nand U6069 (N_6069,N_5827,N_5935);
xor U6070 (N_6070,N_5547,N_5861);
and U6071 (N_6071,N_5584,N_5875);
nor U6072 (N_6072,N_5789,N_5960);
or U6073 (N_6073,N_5550,N_5722);
or U6074 (N_6074,N_5887,N_5586);
nor U6075 (N_6075,N_5971,N_5614);
xnor U6076 (N_6076,N_5576,N_5712);
nand U6077 (N_6077,N_5912,N_5918);
xor U6078 (N_6078,N_5716,N_5590);
and U6079 (N_6079,N_5757,N_5860);
nand U6080 (N_6080,N_5791,N_5972);
nand U6081 (N_6081,N_5682,N_5693);
nand U6082 (N_6082,N_5968,N_5560);
nand U6083 (N_6083,N_5510,N_5744);
and U6084 (N_6084,N_5684,N_5754);
and U6085 (N_6085,N_5585,N_5846);
or U6086 (N_6086,N_5790,N_5621);
and U6087 (N_6087,N_5531,N_5714);
and U6088 (N_6088,N_5591,N_5903);
and U6089 (N_6089,N_5610,N_5874);
and U6090 (N_6090,N_5756,N_5628);
nand U6091 (N_6091,N_5619,N_5954);
or U6092 (N_6092,N_5558,N_5730);
xor U6093 (N_6093,N_5673,N_5650);
or U6094 (N_6094,N_5773,N_5617);
xor U6095 (N_6095,N_5713,N_5955);
and U6096 (N_6096,N_5613,N_5723);
and U6097 (N_6097,N_5502,N_5869);
xnor U6098 (N_6098,N_5907,N_5715);
nand U6099 (N_6099,N_5800,N_5537);
and U6100 (N_6100,N_5931,N_5563);
nand U6101 (N_6101,N_5616,N_5671);
nor U6102 (N_6102,N_5835,N_5966);
and U6103 (N_6103,N_5598,N_5840);
and U6104 (N_6104,N_5894,N_5635);
nor U6105 (N_6105,N_5771,N_5504);
or U6106 (N_6106,N_5982,N_5964);
and U6107 (N_6107,N_5749,N_5664);
xor U6108 (N_6108,N_5804,N_5500);
or U6109 (N_6109,N_5659,N_5505);
nand U6110 (N_6110,N_5556,N_5862);
and U6111 (N_6111,N_5981,N_5809);
or U6112 (N_6112,N_5801,N_5979);
or U6113 (N_6113,N_5577,N_5957);
and U6114 (N_6114,N_5509,N_5527);
and U6115 (N_6115,N_5710,N_5930);
or U6116 (N_6116,N_5605,N_5900);
and U6117 (N_6117,N_5528,N_5609);
and U6118 (N_6118,N_5938,N_5909);
nand U6119 (N_6119,N_5868,N_5759);
xor U6120 (N_6120,N_5525,N_5711);
or U6121 (N_6121,N_5695,N_5988);
nand U6122 (N_6122,N_5765,N_5600);
xnor U6123 (N_6123,N_5780,N_5953);
nand U6124 (N_6124,N_5611,N_5588);
xor U6125 (N_6125,N_5511,N_5538);
or U6126 (N_6126,N_5608,N_5667);
nand U6127 (N_6127,N_5552,N_5998);
or U6128 (N_6128,N_5678,N_5876);
nor U6129 (N_6129,N_5625,N_5818);
nand U6130 (N_6130,N_5825,N_5829);
nor U6131 (N_6131,N_5986,N_5767);
nor U6132 (N_6132,N_5524,N_5833);
nor U6133 (N_6133,N_5752,N_5973);
nand U6134 (N_6134,N_5735,N_5880);
nand U6135 (N_6135,N_5926,N_5885);
xnor U6136 (N_6136,N_5596,N_5859);
and U6137 (N_6137,N_5724,N_5661);
and U6138 (N_6138,N_5823,N_5890);
or U6139 (N_6139,N_5990,N_5898);
nor U6140 (N_6140,N_5854,N_5892);
xnor U6141 (N_6141,N_5631,N_5995);
and U6142 (N_6142,N_5737,N_5741);
nor U6143 (N_6143,N_5721,N_5747);
xnor U6144 (N_6144,N_5574,N_5928);
or U6145 (N_6145,N_5655,N_5808);
xnor U6146 (N_6146,N_5703,N_5534);
nand U6147 (N_6147,N_5763,N_5798);
and U6148 (N_6148,N_5648,N_5521);
and U6149 (N_6149,N_5888,N_5740);
or U6150 (N_6150,N_5906,N_5788);
nand U6151 (N_6151,N_5797,N_5852);
or U6152 (N_6152,N_5812,N_5736);
nor U6153 (N_6153,N_5565,N_5996);
and U6154 (N_6154,N_5526,N_5951);
nor U6155 (N_6155,N_5508,N_5653);
nand U6156 (N_6156,N_5637,N_5783);
nor U6157 (N_6157,N_5607,N_5994);
nand U6158 (N_6158,N_5943,N_5533);
xor U6159 (N_6159,N_5561,N_5962);
and U6160 (N_6160,N_5699,N_5612);
and U6161 (N_6161,N_5883,N_5932);
nand U6162 (N_6162,N_5866,N_5844);
and U6163 (N_6163,N_5940,N_5572);
and U6164 (N_6164,N_5814,N_5718);
nand U6165 (N_6165,N_5646,N_5549);
xor U6166 (N_6166,N_5815,N_5557);
or U6167 (N_6167,N_5949,N_5670);
xnor U6168 (N_6168,N_5555,N_5592);
xor U6169 (N_6169,N_5516,N_5615);
or U6170 (N_6170,N_5562,N_5760);
or U6171 (N_6171,N_5630,N_5769);
and U6172 (N_6172,N_5662,N_5579);
or U6173 (N_6173,N_5811,N_5729);
nor U6174 (N_6174,N_5884,N_5950);
and U6175 (N_6175,N_5649,N_5734);
nand U6176 (N_6176,N_5706,N_5725);
and U6177 (N_6177,N_5700,N_5683);
or U6178 (N_6178,N_5929,N_5632);
nor U6179 (N_6179,N_5806,N_5991);
nor U6180 (N_6180,N_5908,N_5873);
and U6181 (N_6181,N_5848,N_5965);
nor U6182 (N_6182,N_5762,N_5794);
nand U6183 (N_6183,N_5540,N_5515);
and U6184 (N_6184,N_5782,N_5831);
or U6185 (N_6185,N_5503,N_5618);
and U6186 (N_6186,N_5947,N_5742);
and U6187 (N_6187,N_5566,N_5837);
and U6188 (N_6188,N_5785,N_5915);
and U6189 (N_6189,N_5934,N_5707);
nor U6190 (N_6190,N_5977,N_5822);
and U6191 (N_6191,N_5863,N_5901);
xor U6192 (N_6192,N_5697,N_5541);
and U6193 (N_6193,N_5807,N_5559);
xnor U6194 (N_6194,N_5984,N_5640);
or U6195 (N_6195,N_5999,N_5774);
or U6196 (N_6196,N_5910,N_5623);
or U6197 (N_6197,N_5886,N_5656);
or U6198 (N_6198,N_5891,N_5720);
or U6199 (N_6199,N_5512,N_5948);
xor U6200 (N_6200,N_5905,N_5523);
nor U6201 (N_6201,N_5980,N_5870);
nand U6202 (N_6202,N_5776,N_5738);
or U6203 (N_6203,N_5633,N_5927);
and U6204 (N_6204,N_5853,N_5530);
xor U6205 (N_6205,N_5850,N_5732);
and U6206 (N_6206,N_5567,N_5694);
and U6207 (N_6207,N_5989,N_5997);
or U6208 (N_6208,N_5879,N_5805);
xor U6209 (N_6209,N_5897,N_5501);
or U6210 (N_6210,N_5654,N_5792);
or U6211 (N_6211,N_5942,N_5941);
and U6212 (N_6212,N_5641,N_5687);
nand U6213 (N_6213,N_5992,N_5816);
nor U6214 (N_6214,N_5602,N_5952);
and U6215 (N_6215,N_5536,N_5864);
xnor U6216 (N_6216,N_5580,N_5569);
nand U6217 (N_6217,N_5755,N_5570);
and U6218 (N_6218,N_5824,N_5924);
and U6219 (N_6219,N_5638,N_5753);
nor U6220 (N_6220,N_5810,N_5796);
xnor U6221 (N_6221,N_5634,N_5532);
or U6222 (N_6222,N_5878,N_5786);
nand U6223 (N_6223,N_5881,N_5674);
nand U6224 (N_6224,N_5575,N_5685);
nor U6225 (N_6225,N_5937,N_5594);
nand U6226 (N_6226,N_5766,N_5838);
or U6227 (N_6227,N_5690,N_5985);
nand U6228 (N_6228,N_5709,N_5587);
xor U6229 (N_6229,N_5669,N_5919);
xor U6230 (N_6230,N_5652,N_5622);
nand U6231 (N_6231,N_5969,N_5772);
or U6232 (N_6232,N_5675,N_5643);
xor U6233 (N_6233,N_5688,N_5544);
and U6234 (N_6234,N_5899,N_5799);
and U6235 (N_6235,N_5778,N_5925);
xor U6236 (N_6236,N_5507,N_5978);
nand U6237 (N_6237,N_5802,N_5849);
or U6238 (N_6238,N_5597,N_5689);
or U6239 (N_6239,N_5535,N_5913);
and U6240 (N_6240,N_5651,N_5867);
or U6241 (N_6241,N_5696,N_5522);
nand U6242 (N_6242,N_5911,N_5743);
xor U6243 (N_6243,N_5828,N_5851);
and U6244 (N_6244,N_5832,N_5896);
nor U6245 (N_6245,N_5692,N_5944);
nor U6246 (N_6246,N_5959,N_5529);
xnor U6247 (N_6247,N_5784,N_5548);
nand U6248 (N_6248,N_5967,N_5933);
xor U6249 (N_6249,N_5746,N_5647);
nor U6250 (N_6250,N_5604,N_5788);
or U6251 (N_6251,N_5638,N_5884);
xor U6252 (N_6252,N_5846,N_5935);
xnor U6253 (N_6253,N_5707,N_5877);
or U6254 (N_6254,N_5581,N_5852);
or U6255 (N_6255,N_5873,N_5772);
nor U6256 (N_6256,N_5982,N_5566);
nand U6257 (N_6257,N_5977,N_5921);
nand U6258 (N_6258,N_5984,N_5874);
xnor U6259 (N_6259,N_5545,N_5894);
xor U6260 (N_6260,N_5903,N_5893);
or U6261 (N_6261,N_5551,N_5577);
nor U6262 (N_6262,N_5632,N_5815);
and U6263 (N_6263,N_5771,N_5782);
xor U6264 (N_6264,N_5566,N_5668);
and U6265 (N_6265,N_5897,N_5828);
nor U6266 (N_6266,N_5734,N_5799);
and U6267 (N_6267,N_5823,N_5912);
nor U6268 (N_6268,N_5861,N_5782);
or U6269 (N_6269,N_5706,N_5846);
xor U6270 (N_6270,N_5710,N_5990);
nand U6271 (N_6271,N_5917,N_5984);
nor U6272 (N_6272,N_5687,N_5723);
and U6273 (N_6273,N_5702,N_5527);
and U6274 (N_6274,N_5676,N_5541);
nor U6275 (N_6275,N_5983,N_5890);
xnor U6276 (N_6276,N_5566,N_5886);
nand U6277 (N_6277,N_5576,N_5577);
and U6278 (N_6278,N_5579,N_5631);
nor U6279 (N_6279,N_5605,N_5719);
nor U6280 (N_6280,N_5775,N_5974);
xor U6281 (N_6281,N_5972,N_5919);
or U6282 (N_6282,N_5632,N_5568);
nor U6283 (N_6283,N_5640,N_5870);
xor U6284 (N_6284,N_5511,N_5929);
xor U6285 (N_6285,N_5772,N_5638);
and U6286 (N_6286,N_5969,N_5880);
and U6287 (N_6287,N_5920,N_5538);
and U6288 (N_6288,N_5998,N_5651);
and U6289 (N_6289,N_5775,N_5648);
nor U6290 (N_6290,N_5797,N_5843);
nand U6291 (N_6291,N_5556,N_5625);
and U6292 (N_6292,N_5877,N_5789);
nor U6293 (N_6293,N_5748,N_5625);
and U6294 (N_6294,N_5562,N_5840);
nand U6295 (N_6295,N_5867,N_5737);
and U6296 (N_6296,N_5599,N_5587);
xnor U6297 (N_6297,N_5863,N_5579);
xnor U6298 (N_6298,N_5534,N_5913);
nand U6299 (N_6299,N_5575,N_5823);
xnor U6300 (N_6300,N_5696,N_5890);
and U6301 (N_6301,N_5781,N_5523);
and U6302 (N_6302,N_5653,N_5856);
or U6303 (N_6303,N_5743,N_5840);
nor U6304 (N_6304,N_5656,N_5997);
nor U6305 (N_6305,N_5916,N_5680);
nor U6306 (N_6306,N_5761,N_5503);
and U6307 (N_6307,N_5626,N_5649);
or U6308 (N_6308,N_5812,N_5642);
or U6309 (N_6309,N_5749,N_5880);
and U6310 (N_6310,N_5926,N_5722);
nand U6311 (N_6311,N_5655,N_5938);
or U6312 (N_6312,N_5826,N_5561);
and U6313 (N_6313,N_5876,N_5588);
and U6314 (N_6314,N_5753,N_5784);
or U6315 (N_6315,N_5924,N_5703);
xnor U6316 (N_6316,N_5999,N_5917);
nor U6317 (N_6317,N_5677,N_5716);
or U6318 (N_6318,N_5826,N_5539);
or U6319 (N_6319,N_5557,N_5748);
xnor U6320 (N_6320,N_5649,N_5558);
xnor U6321 (N_6321,N_5610,N_5892);
xnor U6322 (N_6322,N_5990,N_5572);
and U6323 (N_6323,N_5682,N_5790);
and U6324 (N_6324,N_5553,N_5933);
and U6325 (N_6325,N_5539,N_5626);
nor U6326 (N_6326,N_5861,N_5898);
or U6327 (N_6327,N_5882,N_5982);
or U6328 (N_6328,N_5851,N_5711);
and U6329 (N_6329,N_5781,N_5902);
nor U6330 (N_6330,N_5545,N_5586);
nor U6331 (N_6331,N_5621,N_5776);
nor U6332 (N_6332,N_5574,N_5563);
nor U6333 (N_6333,N_5522,N_5933);
xnor U6334 (N_6334,N_5758,N_5687);
and U6335 (N_6335,N_5996,N_5758);
nor U6336 (N_6336,N_5960,N_5841);
xnor U6337 (N_6337,N_5816,N_5744);
and U6338 (N_6338,N_5692,N_5865);
or U6339 (N_6339,N_5835,N_5672);
nand U6340 (N_6340,N_5517,N_5793);
or U6341 (N_6341,N_5650,N_5804);
nand U6342 (N_6342,N_5840,N_5581);
and U6343 (N_6343,N_5545,N_5814);
nand U6344 (N_6344,N_5715,N_5813);
nor U6345 (N_6345,N_5517,N_5742);
and U6346 (N_6346,N_5749,N_5595);
xnor U6347 (N_6347,N_5988,N_5878);
or U6348 (N_6348,N_5985,N_5679);
and U6349 (N_6349,N_5748,N_5559);
nand U6350 (N_6350,N_5796,N_5624);
nor U6351 (N_6351,N_5897,N_5968);
nor U6352 (N_6352,N_5731,N_5502);
and U6353 (N_6353,N_5581,N_5637);
or U6354 (N_6354,N_5954,N_5695);
or U6355 (N_6355,N_5685,N_5542);
xor U6356 (N_6356,N_5549,N_5600);
nor U6357 (N_6357,N_5541,N_5850);
nand U6358 (N_6358,N_5704,N_5673);
xnor U6359 (N_6359,N_5852,N_5557);
nand U6360 (N_6360,N_5721,N_5793);
or U6361 (N_6361,N_5774,N_5948);
nand U6362 (N_6362,N_5604,N_5806);
and U6363 (N_6363,N_5924,N_5675);
and U6364 (N_6364,N_5793,N_5887);
xnor U6365 (N_6365,N_5867,N_5682);
nand U6366 (N_6366,N_5944,N_5974);
xor U6367 (N_6367,N_5663,N_5662);
xnor U6368 (N_6368,N_5979,N_5995);
nand U6369 (N_6369,N_5746,N_5598);
nand U6370 (N_6370,N_5845,N_5892);
nor U6371 (N_6371,N_5791,N_5661);
nor U6372 (N_6372,N_5952,N_5961);
nor U6373 (N_6373,N_5790,N_5856);
nand U6374 (N_6374,N_5795,N_5931);
nor U6375 (N_6375,N_5939,N_5828);
xnor U6376 (N_6376,N_5902,N_5835);
nand U6377 (N_6377,N_5818,N_5995);
nand U6378 (N_6378,N_5988,N_5563);
or U6379 (N_6379,N_5921,N_5962);
xnor U6380 (N_6380,N_5552,N_5986);
and U6381 (N_6381,N_5926,N_5607);
nand U6382 (N_6382,N_5724,N_5867);
nand U6383 (N_6383,N_5927,N_5805);
and U6384 (N_6384,N_5970,N_5717);
xnor U6385 (N_6385,N_5901,N_5614);
nor U6386 (N_6386,N_5986,N_5642);
xnor U6387 (N_6387,N_5855,N_5836);
nand U6388 (N_6388,N_5601,N_5854);
xor U6389 (N_6389,N_5873,N_5902);
nor U6390 (N_6390,N_5834,N_5687);
xnor U6391 (N_6391,N_5764,N_5956);
nor U6392 (N_6392,N_5867,N_5904);
xor U6393 (N_6393,N_5977,N_5506);
and U6394 (N_6394,N_5972,N_5895);
or U6395 (N_6395,N_5816,N_5595);
or U6396 (N_6396,N_5755,N_5566);
nand U6397 (N_6397,N_5549,N_5611);
xnor U6398 (N_6398,N_5654,N_5583);
nand U6399 (N_6399,N_5743,N_5752);
nand U6400 (N_6400,N_5885,N_5823);
nor U6401 (N_6401,N_5791,N_5856);
xnor U6402 (N_6402,N_5831,N_5844);
or U6403 (N_6403,N_5942,N_5768);
nand U6404 (N_6404,N_5830,N_5545);
nor U6405 (N_6405,N_5642,N_5989);
or U6406 (N_6406,N_5947,N_5818);
xor U6407 (N_6407,N_5898,N_5996);
and U6408 (N_6408,N_5984,N_5939);
or U6409 (N_6409,N_5799,N_5784);
or U6410 (N_6410,N_5915,N_5669);
and U6411 (N_6411,N_5668,N_5927);
or U6412 (N_6412,N_5784,N_5914);
nand U6413 (N_6413,N_5725,N_5749);
or U6414 (N_6414,N_5646,N_5864);
nor U6415 (N_6415,N_5873,N_5579);
and U6416 (N_6416,N_5683,N_5788);
xnor U6417 (N_6417,N_5964,N_5945);
nand U6418 (N_6418,N_5750,N_5815);
nor U6419 (N_6419,N_5603,N_5899);
or U6420 (N_6420,N_5799,N_5680);
nor U6421 (N_6421,N_5744,N_5575);
or U6422 (N_6422,N_5580,N_5888);
xnor U6423 (N_6423,N_5600,N_5967);
and U6424 (N_6424,N_5793,N_5911);
xor U6425 (N_6425,N_5527,N_5840);
xnor U6426 (N_6426,N_5699,N_5951);
nand U6427 (N_6427,N_5598,N_5959);
nand U6428 (N_6428,N_5798,N_5608);
nand U6429 (N_6429,N_5508,N_5532);
or U6430 (N_6430,N_5760,N_5570);
nor U6431 (N_6431,N_5874,N_5660);
nor U6432 (N_6432,N_5547,N_5608);
nand U6433 (N_6433,N_5903,N_5949);
nand U6434 (N_6434,N_5741,N_5646);
or U6435 (N_6435,N_5864,N_5762);
nor U6436 (N_6436,N_5793,N_5557);
nand U6437 (N_6437,N_5707,N_5770);
nand U6438 (N_6438,N_5693,N_5942);
nand U6439 (N_6439,N_5971,N_5859);
or U6440 (N_6440,N_5608,N_5753);
nor U6441 (N_6441,N_5990,N_5757);
xor U6442 (N_6442,N_5678,N_5596);
nand U6443 (N_6443,N_5771,N_5798);
or U6444 (N_6444,N_5743,N_5861);
and U6445 (N_6445,N_5930,N_5933);
nand U6446 (N_6446,N_5716,N_5525);
xnor U6447 (N_6447,N_5549,N_5578);
and U6448 (N_6448,N_5944,N_5679);
and U6449 (N_6449,N_5648,N_5538);
or U6450 (N_6450,N_5507,N_5599);
xnor U6451 (N_6451,N_5797,N_5575);
xor U6452 (N_6452,N_5746,N_5687);
xnor U6453 (N_6453,N_5601,N_5531);
and U6454 (N_6454,N_5860,N_5913);
nand U6455 (N_6455,N_5821,N_5918);
and U6456 (N_6456,N_5832,N_5796);
nor U6457 (N_6457,N_5852,N_5543);
nor U6458 (N_6458,N_5709,N_5564);
nand U6459 (N_6459,N_5610,N_5989);
xnor U6460 (N_6460,N_5765,N_5541);
nor U6461 (N_6461,N_5537,N_5884);
nand U6462 (N_6462,N_5765,N_5825);
nor U6463 (N_6463,N_5851,N_5656);
nand U6464 (N_6464,N_5529,N_5789);
xor U6465 (N_6465,N_5563,N_5962);
or U6466 (N_6466,N_5877,N_5527);
nor U6467 (N_6467,N_5861,N_5561);
or U6468 (N_6468,N_5866,N_5862);
xnor U6469 (N_6469,N_5921,N_5877);
nand U6470 (N_6470,N_5577,N_5716);
nand U6471 (N_6471,N_5626,N_5762);
or U6472 (N_6472,N_5853,N_5970);
xnor U6473 (N_6473,N_5596,N_5970);
nand U6474 (N_6474,N_5552,N_5818);
xnor U6475 (N_6475,N_5797,N_5742);
nor U6476 (N_6476,N_5869,N_5828);
and U6477 (N_6477,N_5650,N_5677);
or U6478 (N_6478,N_5953,N_5882);
and U6479 (N_6479,N_5630,N_5727);
nand U6480 (N_6480,N_5989,N_5658);
or U6481 (N_6481,N_5857,N_5946);
and U6482 (N_6482,N_5800,N_5950);
or U6483 (N_6483,N_5717,N_5917);
or U6484 (N_6484,N_5940,N_5936);
and U6485 (N_6485,N_5666,N_5965);
or U6486 (N_6486,N_5600,N_5607);
nand U6487 (N_6487,N_5703,N_5689);
xor U6488 (N_6488,N_5860,N_5866);
or U6489 (N_6489,N_5558,N_5797);
nor U6490 (N_6490,N_5859,N_5935);
or U6491 (N_6491,N_5687,N_5913);
nor U6492 (N_6492,N_5857,N_5929);
and U6493 (N_6493,N_5907,N_5645);
or U6494 (N_6494,N_5516,N_5841);
or U6495 (N_6495,N_5708,N_5846);
nand U6496 (N_6496,N_5878,N_5855);
and U6497 (N_6497,N_5620,N_5537);
nor U6498 (N_6498,N_5986,N_5727);
or U6499 (N_6499,N_5570,N_5947);
or U6500 (N_6500,N_6375,N_6278);
nor U6501 (N_6501,N_6388,N_6289);
nand U6502 (N_6502,N_6123,N_6383);
and U6503 (N_6503,N_6168,N_6019);
and U6504 (N_6504,N_6448,N_6055);
and U6505 (N_6505,N_6322,N_6348);
nand U6506 (N_6506,N_6028,N_6265);
nor U6507 (N_6507,N_6136,N_6171);
and U6508 (N_6508,N_6430,N_6426);
xnor U6509 (N_6509,N_6102,N_6064);
or U6510 (N_6510,N_6143,N_6488);
and U6511 (N_6511,N_6090,N_6196);
and U6512 (N_6512,N_6231,N_6207);
and U6513 (N_6513,N_6454,N_6070);
xnor U6514 (N_6514,N_6482,N_6126);
xor U6515 (N_6515,N_6145,N_6398);
xnor U6516 (N_6516,N_6007,N_6342);
or U6517 (N_6517,N_6323,N_6275);
nand U6518 (N_6518,N_6054,N_6310);
and U6519 (N_6519,N_6144,N_6379);
and U6520 (N_6520,N_6023,N_6268);
xnor U6521 (N_6521,N_6436,N_6329);
or U6522 (N_6522,N_6253,N_6072);
and U6523 (N_6523,N_6262,N_6327);
nand U6524 (N_6524,N_6315,N_6319);
or U6525 (N_6525,N_6121,N_6324);
nor U6526 (N_6526,N_6288,N_6490);
or U6527 (N_6527,N_6190,N_6391);
nor U6528 (N_6528,N_6489,N_6321);
and U6529 (N_6529,N_6073,N_6131);
and U6530 (N_6530,N_6456,N_6021);
nor U6531 (N_6531,N_6166,N_6230);
and U6532 (N_6532,N_6420,N_6179);
or U6533 (N_6533,N_6439,N_6014);
nor U6534 (N_6534,N_6421,N_6018);
or U6535 (N_6535,N_6213,N_6229);
or U6536 (N_6536,N_6336,N_6440);
nand U6537 (N_6537,N_6237,N_6115);
nand U6538 (N_6538,N_6099,N_6378);
nand U6539 (N_6539,N_6418,N_6311);
xnor U6540 (N_6540,N_6067,N_6303);
nor U6541 (N_6541,N_6350,N_6113);
and U6542 (N_6542,N_6002,N_6431);
nor U6543 (N_6543,N_6382,N_6432);
nand U6544 (N_6544,N_6088,N_6455);
and U6545 (N_6545,N_6337,N_6453);
xnor U6546 (N_6546,N_6114,N_6024);
or U6547 (N_6547,N_6148,N_6267);
and U6548 (N_6548,N_6218,N_6441);
or U6549 (N_6549,N_6025,N_6367);
nor U6550 (N_6550,N_6380,N_6050);
nor U6551 (N_6551,N_6298,N_6320);
and U6552 (N_6552,N_6347,N_6352);
and U6553 (N_6553,N_6328,N_6344);
and U6554 (N_6554,N_6465,N_6110);
nor U6555 (N_6555,N_6365,N_6239);
xor U6556 (N_6556,N_6437,N_6356);
nor U6557 (N_6557,N_6080,N_6334);
xor U6558 (N_6558,N_6212,N_6447);
or U6559 (N_6559,N_6191,N_6180);
nor U6560 (N_6560,N_6236,N_6247);
nor U6561 (N_6561,N_6009,N_6033);
xor U6562 (N_6562,N_6470,N_6053);
xor U6563 (N_6563,N_6157,N_6097);
nand U6564 (N_6564,N_6345,N_6433);
xnor U6565 (N_6565,N_6079,N_6361);
and U6566 (N_6566,N_6029,N_6473);
and U6567 (N_6567,N_6075,N_6127);
nand U6568 (N_6568,N_6175,N_6165);
nor U6569 (N_6569,N_6346,N_6122);
nand U6570 (N_6570,N_6402,N_6299);
or U6571 (N_6571,N_6373,N_6130);
or U6572 (N_6572,N_6005,N_6251);
or U6573 (N_6573,N_6140,N_6174);
nand U6574 (N_6574,N_6394,N_6246);
xnor U6575 (N_6575,N_6049,N_6086);
nor U6576 (N_6576,N_6249,N_6201);
and U6577 (N_6577,N_6325,N_6296);
or U6578 (N_6578,N_6192,N_6038);
or U6579 (N_6579,N_6227,N_6034);
nand U6580 (N_6580,N_6360,N_6068);
or U6581 (N_6581,N_6195,N_6442);
or U6582 (N_6582,N_6232,N_6458);
or U6583 (N_6583,N_6083,N_6167);
nor U6584 (N_6584,N_6063,N_6184);
xor U6585 (N_6585,N_6294,N_6133);
nor U6586 (N_6586,N_6417,N_6369);
xor U6587 (N_6587,N_6221,N_6381);
nand U6588 (N_6588,N_6235,N_6012);
and U6589 (N_6589,N_6395,N_6491);
nor U6590 (N_6590,N_6318,N_6061);
nand U6591 (N_6591,N_6228,N_6098);
or U6592 (N_6592,N_6284,N_6177);
xor U6593 (N_6593,N_6468,N_6312);
nand U6594 (N_6594,N_6187,N_6031);
nand U6595 (N_6595,N_6172,N_6466);
or U6596 (N_6596,N_6384,N_6156);
nor U6597 (N_6597,N_6343,N_6015);
nand U6598 (N_6598,N_6158,N_6416);
or U6599 (N_6599,N_6052,N_6377);
nor U6600 (N_6600,N_6393,N_6413);
and U6601 (N_6601,N_6139,N_6176);
xor U6602 (N_6602,N_6058,N_6170);
and U6603 (N_6603,N_6095,N_6309);
nand U6604 (N_6604,N_6326,N_6405);
xnor U6605 (N_6605,N_6013,N_6152);
nand U6606 (N_6606,N_6423,N_6254);
nor U6607 (N_6607,N_6459,N_6335);
xnor U6608 (N_6608,N_6464,N_6357);
xor U6609 (N_6609,N_6155,N_6332);
nand U6610 (N_6610,N_6198,N_6186);
nor U6611 (N_6611,N_6477,N_6020);
nand U6612 (N_6612,N_6355,N_6291);
nor U6613 (N_6613,N_6290,N_6486);
nor U6614 (N_6614,N_6371,N_6189);
and U6615 (N_6615,N_6163,N_6017);
xor U6616 (N_6616,N_6208,N_6082);
nand U6617 (N_6617,N_6387,N_6065);
or U6618 (N_6618,N_6103,N_6330);
or U6619 (N_6619,N_6222,N_6415);
xor U6620 (N_6620,N_6406,N_6225);
or U6621 (N_6621,N_6409,N_6480);
or U6622 (N_6622,N_6022,N_6210);
xor U6623 (N_6623,N_6316,N_6071);
or U6624 (N_6624,N_6446,N_6194);
nand U6625 (N_6625,N_6258,N_6435);
nand U6626 (N_6626,N_6162,N_6001);
and U6627 (N_6627,N_6169,N_6016);
and U6628 (N_6628,N_6183,N_6425);
nor U6629 (N_6629,N_6483,N_6153);
or U6630 (N_6630,N_6493,N_6457);
and U6631 (N_6631,N_6469,N_6385);
nand U6632 (N_6632,N_6134,N_6112);
and U6633 (N_6633,N_6363,N_6259);
nor U6634 (N_6634,N_6216,N_6006);
xnor U6635 (N_6635,N_6410,N_6478);
nor U6636 (N_6636,N_6285,N_6217);
or U6637 (N_6637,N_6474,N_6147);
and U6638 (N_6638,N_6339,N_6209);
xor U6639 (N_6639,N_6389,N_6314);
nor U6640 (N_6640,N_6215,N_6399);
nor U6641 (N_6641,N_6331,N_6214);
nand U6642 (N_6642,N_6403,N_6085);
and U6643 (N_6643,N_6250,N_6450);
or U6644 (N_6644,N_6358,N_6317);
or U6645 (N_6645,N_6084,N_6414);
or U6646 (N_6646,N_6044,N_6359);
nor U6647 (N_6647,N_6076,N_6248);
xor U6648 (N_6648,N_6293,N_6269);
nor U6649 (N_6649,N_6492,N_6370);
xnor U6650 (N_6650,N_6241,N_6092);
xor U6651 (N_6651,N_6242,N_6471);
and U6652 (N_6652,N_6264,N_6104);
xor U6653 (N_6653,N_6108,N_6047);
nor U6654 (N_6654,N_6173,N_6100);
or U6655 (N_6655,N_6467,N_6069);
nand U6656 (N_6656,N_6282,N_6074);
nand U6657 (N_6657,N_6392,N_6182);
xor U6658 (N_6658,N_6485,N_6374);
nand U6659 (N_6659,N_6300,N_6164);
xnor U6660 (N_6660,N_6056,N_6185);
nand U6661 (N_6661,N_6461,N_6035);
nand U6662 (N_6662,N_6341,N_6261);
or U6663 (N_6663,N_6245,N_6030);
and U6664 (N_6664,N_6151,N_6041);
nand U6665 (N_6665,N_6449,N_6277);
or U6666 (N_6666,N_6181,N_6066);
or U6667 (N_6667,N_6495,N_6135);
xnor U6668 (N_6668,N_6481,N_6287);
nand U6669 (N_6669,N_6260,N_6101);
or U6670 (N_6670,N_6270,N_6243);
or U6671 (N_6671,N_6256,N_6484);
xnor U6672 (N_6672,N_6472,N_6438);
and U6673 (N_6673,N_6032,N_6271);
and U6674 (N_6674,N_6301,N_6408);
nor U6675 (N_6675,N_6302,N_6105);
xor U6676 (N_6676,N_6349,N_6364);
xor U6677 (N_6677,N_6159,N_6008);
or U6678 (N_6678,N_6116,N_6257);
or U6679 (N_6679,N_6400,N_6305);
and U6680 (N_6680,N_6279,N_6427);
nor U6681 (N_6681,N_6109,N_6091);
nand U6682 (N_6682,N_6202,N_6129);
nand U6683 (N_6683,N_6338,N_6226);
or U6684 (N_6684,N_6276,N_6057);
or U6685 (N_6685,N_6434,N_6146);
nand U6686 (N_6686,N_6238,N_6093);
nand U6687 (N_6687,N_6306,N_6132);
or U6688 (N_6688,N_6204,N_6137);
nand U6689 (N_6689,N_6118,N_6026);
nor U6690 (N_6690,N_6087,N_6263);
nor U6691 (N_6691,N_6460,N_6128);
xnor U6692 (N_6692,N_6004,N_6160);
nand U6693 (N_6693,N_6150,N_6497);
nor U6694 (N_6694,N_6266,N_6106);
or U6695 (N_6695,N_6487,N_6199);
and U6696 (N_6696,N_6233,N_6479);
nand U6697 (N_6697,N_6011,N_6081);
nor U6698 (N_6698,N_6476,N_6295);
or U6699 (N_6699,N_6397,N_6445);
nor U6700 (N_6700,N_6000,N_6366);
or U6701 (N_6701,N_6444,N_6313);
or U6702 (N_6702,N_6205,N_6125);
xnor U6703 (N_6703,N_6178,N_6188);
or U6704 (N_6704,N_6422,N_6039);
xnor U6705 (N_6705,N_6498,N_6094);
xnor U6706 (N_6706,N_6308,N_6220);
nor U6707 (N_6707,N_6224,N_6197);
or U6708 (N_6708,N_6124,N_6048);
xnor U6709 (N_6709,N_6419,N_6424);
nand U6710 (N_6710,N_6412,N_6333);
xor U6711 (N_6711,N_6351,N_6353);
xor U6712 (N_6712,N_6252,N_6244);
nand U6713 (N_6713,N_6060,N_6273);
xnor U6714 (N_6714,N_6119,N_6283);
xnor U6715 (N_6715,N_6281,N_6451);
nor U6716 (N_6716,N_6203,N_6193);
nor U6717 (N_6717,N_6219,N_6045);
or U6718 (N_6718,N_6200,N_6107);
or U6719 (N_6719,N_6206,N_6386);
xor U6720 (N_6720,N_6362,N_6059);
or U6721 (N_6721,N_6274,N_6141);
and U6722 (N_6722,N_6396,N_6111);
and U6723 (N_6723,N_6376,N_6036);
xnor U6724 (N_6724,N_6496,N_6062);
or U6725 (N_6725,N_6161,N_6372);
and U6726 (N_6726,N_6429,N_6077);
and U6727 (N_6727,N_6223,N_6240);
nor U6728 (N_6728,N_6286,N_6407);
xnor U6729 (N_6729,N_6272,N_6089);
xnor U6730 (N_6730,N_6494,N_6401);
nand U6731 (N_6731,N_6304,N_6390);
nor U6732 (N_6732,N_6043,N_6037);
nor U6733 (N_6733,N_6096,N_6463);
or U6734 (N_6734,N_6211,N_6027);
nor U6735 (N_6735,N_6404,N_6051);
nor U6736 (N_6736,N_6120,N_6046);
xor U6737 (N_6737,N_6499,N_6149);
xor U6738 (N_6738,N_6234,N_6307);
or U6739 (N_6739,N_6340,N_6154);
nor U6740 (N_6740,N_6452,N_6042);
xor U6741 (N_6741,N_6428,N_6443);
nor U6742 (N_6742,N_6138,N_6010);
or U6743 (N_6743,N_6280,N_6078);
xnor U6744 (N_6744,N_6255,N_6411);
or U6745 (N_6745,N_6462,N_6003);
xor U6746 (N_6746,N_6354,N_6117);
and U6747 (N_6747,N_6297,N_6475);
xnor U6748 (N_6748,N_6142,N_6292);
and U6749 (N_6749,N_6040,N_6368);
nand U6750 (N_6750,N_6204,N_6150);
nand U6751 (N_6751,N_6227,N_6159);
nor U6752 (N_6752,N_6070,N_6267);
and U6753 (N_6753,N_6458,N_6235);
nor U6754 (N_6754,N_6214,N_6363);
or U6755 (N_6755,N_6345,N_6085);
and U6756 (N_6756,N_6086,N_6246);
nand U6757 (N_6757,N_6031,N_6452);
nor U6758 (N_6758,N_6061,N_6332);
nand U6759 (N_6759,N_6071,N_6285);
xnor U6760 (N_6760,N_6306,N_6240);
nor U6761 (N_6761,N_6348,N_6381);
and U6762 (N_6762,N_6412,N_6414);
xor U6763 (N_6763,N_6495,N_6452);
and U6764 (N_6764,N_6439,N_6402);
xnor U6765 (N_6765,N_6107,N_6318);
xor U6766 (N_6766,N_6015,N_6127);
nand U6767 (N_6767,N_6368,N_6265);
xor U6768 (N_6768,N_6062,N_6392);
xor U6769 (N_6769,N_6478,N_6310);
nand U6770 (N_6770,N_6133,N_6291);
or U6771 (N_6771,N_6128,N_6486);
and U6772 (N_6772,N_6096,N_6413);
nand U6773 (N_6773,N_6307,N_6437);
xor U6774 (N_6774,N_6307,N_6007);
or U6775 (N_6775,N_6273,N_6457);
or U6776 (N_6776,N_6248,N_6196);
xor U6777 (N_6777,N_6479,N_6472);
nor U6778 (N_6778,N_6051,N_6289);
and U6779 (N_6779,N_6252,N_6158);
nand U6780 (N_6780,N_6208,N_6145);
nand U6781 (N_6781,N_6072,N_6388);
and U6782 (N_6782,N_6055,N_6212);
nor U6783 (N_6783,N_6182,N_6163);
nor U6784 (N_6784,N_6328,N_6205);
and U6785 (N_6785,N_6169,N_6301);
xnor U6786 (N_6786,N_6173,N_6122);
and U6787 (N_6787,N_6312,N_6011);
nand U6788 (N_6788,N_6473,N_6233);
xor U6789 (N_6789,N_6291,N_6026);
or U6790 (N_6790,N_6308,N_6019);
xor U6791 (N_6791,N_6408,N_6187);
or U6792 (N_6792,N_6366,N_6395);
xor U6793 (N_6793,N_6361,N_6396);
and U6794 (N_6794,N_6282,N_6235);
nand U6795 (N_6795,N_6024,N_6461);
nand U6796 (N_6796,N_6239,N_6281);
and U6797 (N_6797,N_6439,N_6323);
xnor U6798 (N_6798,N_6286,N_6090);
or U6799 (N_6799,N_6068,N_6281);
and U6800 (N_6800,N_6129,N_6015);
or U6801 (N_6801,N_6381,N_6271);
nor U6802 (N_6802,N_6031,N_6339);
nand U6803 (N_6803,N_6125,N_6430);
nor U6804 (N_6804,N_6235,N_6317);
and U6805 (N_6805,N_6316,N_6008);
xnor U6806 (N_6806,N_6196,N_6161);
nor U6807 (N_6807,N_6189,N_6330);
xnor U6808 (N_6808,N_6091,N_6147);
nand U6809 (N_6809,N_6086,N_6063);
nand U6810 (N_6810,N_6219,N_6200);
and U6811 (N_6811,N_6177,N_6100);
nand U6812 (N_6812,N_6022,N_6139);
xor U6813 (N_6813,N_6304,N_6360);
xnor U6814 (N_6814,N_6184,N_6307);
and U6815 (N_6815,N_6147,N_6319);
or U6816 (N_6816,N_6330,N_6417);
nor U6817 (N_6817,N_6149,N_6268);
nor U6818 (N_6818,N_6248,N_6243);
nand U6819 (N_6819,N_6159,N_6380);
nor U6820 (N_6820,N_6113,N_6314);
nand U6821 (N_6821,N_6125,N_6400);
nor U6822 (N_6822,N_6391,N_6324);
and U6823 (N_6823,N_6209,N_6292);
nand U6824 (N_6824,N_6071,N_6308);
or U6825 (N_6825,N_6008,N_6085);
or U6826 (N_6826,N_6220,N_6057);
nand U6827 (N_6827,N_6318,N_6469);
or U6828 (N_6828,N_6188,N_6319);
nand U6829 (N_6829,N_6019,N_6028);
or U6830 (N_6830,N_6293,N_6202);
xnor U6831 (N_6831,N_6049,N_6424);
nor U6832 (N_6832,N_6435,N_6178);
nand U6833 (N_6833,N_6011,N_6377);
and U6834 (N_6834,N_6109,N_6391);
nand U6835 (N_6835,N_6415,N_6320);
nand U6836 (N_6836,N_6396,N_6416);
or U6837 (N_6837,N_6470,N_6028);
nand U6838 (N_6838,N_6338,N_6227);
nor U6839 (N_6839,N_6322,N_6349);
nor U6840 (N_6840,N_6368,N_6170);
nor U6841 (N_6841,N_6381,N_6302);
and U6842 (N_6842,N_6413,N_6021);
nor U6843 (N_6843,N_6415,N_6423);
nand U6844 (N_6844,N_6128,N_6440);
or U6845 (N_6845,N_6475,N_6353);
and U6846 (N_6846,N_6183,N_6005);
nor U6847 (N_6847,N_6186,N_6437);
xor U6848 (N_6848,N_6288,N_6146);
nand U6849 (N_6849,N_6488,N_6024);
and U6850 (N_6850,N_6406,N_6298);
nand U6851 (N_6851,N_6180,N_6174);
xor U6852 (N_6852,N_6411,N_6454);
nand U6853 (N_6853,N_6096,N_6467);
and U6854 (N_6854,N_6007,N_6069);
or U6855 (N_6855,N_6065,N_6253);
nand U6856 (N_6856,N_6106,N_6462);
nor U6857 (N_6857,N_6013,N_6321);
nor U6858 (N_6858,N_6109,N_6120);
nor U6859 (N_6859,N_6382,N_6353);
and U6860 (N_6860,N_6225,N_6189);
nor U6861 (N_6861,N_6482,N_6164);
xnor U6862 (N_6862,N_6313,N_6375);
nand U6863 (N_6863,N_6006,N_6297);
nor U6864 (N_6864,N_6163,N_6409);
nand U6865 (N_6865,N_6499,N_6461);
nor U6866 (N_6866,N_6327,N_6418);
nand U6867 (N_6867,N_6144,N_6002);
or U6868 (N_6868,N_6257,N_6235);
nand U6869 (N_6869,N_6420,N_6457);
xnor U6870 (N_6870,N_6124,N_6113);
and U6871 (N_6871,N_6092,N_6495);
or U6872 (N_6872,N_6256,N_6492);
nor U6873 (N_6873,N_6280,N_6127);
and U6874 (N_6874,N_6468,N_6268);
or U6875 (N_6875,N_6433,N_6108);
or U6876 (N_6876,N_6127,N_6410);
and U6877 (N_6877,N_6431,N_6368);
xor U6878 (N_6878,N_6009,N_6473);
xor U6879 (N_6879,N_6074,N_6373);
nor U6880 (N_6880,N_6314,N_6017);
xor U6881 (N_6881,N_6439,N_6351);
and U6882 (N_6882,N_6125,N_6204);
nand U6883 (N_6883,N_6206,N_6177);
nor U6884 (N_6884,N_6186,N_6047);
nand U6885 (N_6885,N_6390,N_6182);
nand U6886 (N_6886,N_6034,N_6073);
nor U6887 (N_6887,N_6469,N_6116);
and U6888 (N_6888,N_6051,N_6053);
and U6889 (N_6889,N_6292,N_6016);
xor U6890 (N_6890,N_6008,N_6036);
nor U6891 (N_6891,N_6316,N_6091);
or U6892 (N_6892,N_6053,N_6496);
and U6893 (N_6893,N_6147,N_6330);
xnor U6894 (N_6894,N_6480,N_6050);
and U6895 (N_6895,N_6166,N_6152);
and U6896 (N_6896,N_6305,N_6213);
nor U6897 (N_6897,N_6238,N_6067);
nor U6898 (N_6898,N_6051,N_6133);
xor U6899 (N_6899,N_6489,N_6345);
or U6900 (N_6900,N_6060,N_6152);
or U6901 (N_6901,N_6469,N_6356);
xnor U6902 (N_6902,N_6291,N_6043);
nor U6903 (N_6903,N_6100,N_6081);
nand U6904 (N_6904,N_6368,N_6219);
nand U6905 (N_6905,N_6062,N_6386);
nand U6906 (N_6906,N_6451,N_6133);
or U6907 (N_6907,N_6009,N_6300);
and U6908 (N_6908,N_6487,N_6269);
or U6909 (N_6909,N_6409,N_6283);
xor U6910 (N_6910,N_6372,N_6043);
nor U6911 (N_6911,N_6432,N_6067);
or U6912 (N_6912,N_6044,N_6487);
or U6913 (N_6913,N_6298,N_6015);
nor U6914 (N_6914,N_6145,N_6000);
and U6915 (N_6915,N_6166,N_6318);
xnor U6916 (N_6916,N_6070,N_6324);
nand U6917 (N_6917,N_6448,N_6424);
xnor U6918 (N_6918,N_6420,N_6078);
and U6919 (N_6919,N_6127,N_6293);
or U6920 (N_6920,N_6206,N_6427);
nand U6921 (N_6921,N_6170,N_6006);
xor U6922 (N_6922,N_6022,N_6487);
xor U6923 (N_6923,N_6452,N_6145);
nand U6924 (N_6924,N_6203,N_6101);
and U6925 (N_6925,N_6017,N_6137);
and U6926 (N_6926,N_6322,N_6007);
xnor U6927 (N_6927,N_6323,N_6118);
nor U6928 (N_6928,N_6066,N_6131);
nand U6929 (N_6929,N_6495,N_6072);
or U6930 (N_6930,N_6356,N_6343);
or U6931 (N_6931,N_6406,N_6423);
nand U6932 (N_6932,N_6281,N_6103);
nand U6933 (N_6933,N_6080,N_6239);
nor U6934 (N_6934,N_6289,N_6303);
nor U6935 (N_6935,N_6085,N_6122);
xnor U6936 (N_6936,N_6152,N_6471);
nor U6937 (N_6937,N_6116,N_6404);
and U6938 (N_6938,N_6358,N_6289);
nand U6939 (N_6939,N_6193,N_6117);
or U6940 (N_6940,N_6231,N_6072);
nor U6941 (N_6941,N_6118,N_6066);
or U6942 (N_6942,N_6016,N_6227);
and U6943 (N_6943,N_6363,N_6080);
nand U6944 (N_6944,N_6261,N_6322);
xnor U6945 (N_6945,N_6051,N_6371);
and U6946 (N_6946,N_6229,N_6461);
nor U6947 (N_6947,N_6125,N_6322);
nand U6948 (N_6948,N_6259,N_6430);
xnor U6949 (N_6949,N_6460,N_6408);
xnor U6950 (N_6950,N_6216,N_6482);
xor U6951 (N_6951,N_6126,N_6019);
nand U6952 (N_6952,N_6274,N_6171);
or U6953 (N_6953,N_6344,N_6219);
or U6954 (N_6954,N_6043,N_6144);
or U6955 (N_6955,N_6162,N_6493);
nor U6956 (N_6956,N_6083,N_6061);
or U6957 (N_6957,N_6147,N_6469);
and U6958 (N_6958,N_6495,N_6205);
xor U6959 (N_6959,N_6051,N_6200);
and U6960 (N_6960,N_6053,N_6360);
and U6961 (N_6961,N_6111,N_6018);
or U6962 (N_6962,N_6376,N_6468);
nand U6963 (N_6963,N_6064,N_6082);
nand U6964 (N_6964,N_6277,N_6101);
or U6965 (N_6965,N_6185,N_6139);
xor U6966 (N_6966,N_6036,N_6338);
nor U6967 (N_6967,N_6354,N_6418);
xor U6968 (N_6968,N_6246,N_6045);
and U6969 (N_6969,N_6252,N_6379);
nor U6970 (N_6970,N_6200,N_6379);
nand U6971 (N_6971,N_6181,N_6117);
nor U6972 (N_6972,N_6398,N_6112);
and U6973 (N_6973,N_6289,N_6300);
nor U6974 (N_6974,N_6302,N_6493);
and U6975 (N_6975,N_6363,N_6221);
and U6976 (N_6976,N_6417,N_6128);
and U6977 (N_6977,N_6108,N_6235);
or U6978 (N_6978,N_6050,N_6420);
nand U6979 (N_6979,N_6027,N_6130);
nand U6980 (N_6980,N_6190,N_6029);
xnor U6981 (N_6981,N_6405,N_6409);
xnor U6982 (N_6982,N_6437,N_6204);
or U6983 (N_6983,N_6255,N_6216);
nor U6984 (N_6984,N_6098,N_6217);
nand U6985 (N_6985,N_6301,N_6359);
and U6986 (N_6986,N_6266,N_6075);
nor U6987 (N_6987,N_6412,N_6173);
or U6988 (N_6988,N_6020,N_6459);
xnor U6989 (N_6989,N_6397,N_6349);
nor U6990 (N_6990,N_6015,N_6031);
or U6991 (N_6991,N_6006,N_6233);
and U6992 (N_6992,N_6327,N_6052);
and U6993 (N_6993,N_6380,N_6053);
nand U6994 (N_6994,N_6491,N_6238);
xnor U6995 (N_6995,N_6386,N_6255);
xor U6996 (N_6996,N_6394,N_6319);
or U6997 (N_6997,N_6424,N_6015);
or U6998 (N_6998,N_6136,N_6134);
nand U6999 (N_6999,N_6319,N_6456);
xnor U7000 (N_7000,N_6821,N_6588);
or U7001 (N_7001,N_6632,N_6891);
nor U7002 (N_7002,N_6546,N_6978);
nand U7003 (N_7003,N_6600,N_6793);
xor U7004 (N_7004,N_6753,N_6551);
nor U7005 (N_7005,N_6622,N_6791);
nand U7006 (N_7006,N_6537,N_6956);
nand U7007 (N_7007,N_6807,N_6716);
nand U7008 (N_7008,N_6726,N_6663);
nand U7009 (N_7009,N_6813,N_6902);
xor U7010 (N_7010,N_6987,N_6621);
or U7011 (N_7011,N_6961,N_6779);
nor U7012 (N_7012,N_6989,N_6522);
xor U7013 (N_7013,N_6721,N_6520);
xnor U7014 (N_7014,N_6919,N_6802);
or U7015 (N_7015,N_6921,N_6519);
xor U7016 (N_7016,N_6893,N_6680);
and U7017 (N_7017,N_6831,N_6682);
or U7018 (N_7018,N_6688,N_6900);
and U7019 (N_7019,N_6950,N_6971);
xnor U7020 (N_7020,N_6722,N_6637);
xnor U7021 (N_7021,N_6641,N_6727);
and U7022 (N_7022,N_6604,N_6613);
and U7023 (N_7023,N_6506,N_6589);
xnor U7024 (N_7024,N_6936,N_6881);
or U7025 (N_7025,N_6633,N_6904);
nand U7026 (N_7026,N_6861,N_6804);
xor U7027 (N_7027,N_6918,N_6880);
nor U7028 (N_7028,N_6736,N_6877);
nand U7029 (N_7029,N_6940,N_6835);
or U7030 (N_7030,N_6573,N_6754);
nand U7031 (N_7031,N_6512,N_6781);
nand U7032 (N_7032,N_6647,N_6805);
nor U7033 (N_7033,N_6908,N_6827);
or U7034 (N_7034,N_6640,N_6550);
nor U7035 (N_7035,N_6595,N_6937);
nand U7036 (N_7036,N_6643,N_6742);
nand U7037 (N_7037,N_6645,N_6694);
or U7038 (N_7038,N_6585,N_6664);
xnor U7039 (N_7039,N_6759,N_6549);
nor U7040 (N_7040,N_6684,N_6783);
or U7041 (N_7041,N_6703,N_6543);
xnor U7042 (N_7042,N_6746,N_6887);
nor U7043 (N_7043,N_6623,N_6508);
xor U7044 (N_7044,N_6796,N_6913);
nand U7045 (N_7045,N_6872,N_6922);
and U7046 (N_7046,N_6701,N_6780);
and U7047 (N_7047,N_6614,N_6859);
nor U7048 (N_7048,N_6619,N_6733);
xor U7049 (N_7049,N_6724,N_6625);
or U7050 (N_7050,N_6709,N_6931);
nor U7051 (N_7051,N_6564,N_6725);
and U7052 (N_7052,N_6959,N_6696);
and U7053 (N_7053,N_6552,N_6933);
or U7054 (N_7054,N_6504,N_6609);
or U7055 (N_7055,N_6545,N_6980);
nor U7056 (N_7056,N_6732,N_6958);
xor U7057 (N_7057,N_6533,N_6832);
xnor U7058 (N_7058,N_6756,N_6636);
and U7059 (N_7059,N_6705,N_6639);
and U7060 (N_7060,N_6734,N_6862);
or U7061 (N_7061,N_6955,N_6909);
xnor U7062 (N_7062,N_6778,N_6888);
or U7063 (N_7063,N_6516,N_6882);
xnor U7064 (N_7064,N_6914,N_6523);
nor U7065 (N_7065,N_6953,N_6767);
nor U7066 (N_7066,N_6670,N_6648);
or U7067 (N_7067,N_6984,N_6720);
nor U7068 (N_7068,N_6762,N_6521);
xor U7069 (N_7069,N_6841,N_6842);
nand U7070 (N_7070,N_6917,N_6534);
and U7071 (N_7071,N_6990,N_6879);
and U7072 (N_7072,N_6886,N_6593);
nand U7073 (N_7073,N_6749,N_6566);
and U7074 (N_7074,N_6743,N_6890);
or U7075 (N_7075,N_6706,N_6603);
and U7076 (N_7076,N_6517,N_6991);
or U7077 (N_7077,N_6855,N_6938);
xor U7078 (N_7078,N_6652,N_6620);
or U7079 (N_7079,N_6799,N_6681);
or U7080 (N_7080,N_6849,N_6968);
and U7081 (N_7081,N_6697,N_6826);
and U7082 (N_7082,N_6867,N_6848);
and U7083 (N_7083,N_6577,N_6833);
or U7084 (N_7084,N_6617,N_6760);
nor U7085 (N_7085,N_6692,N_6737);
xnor U7086 (N_7086,N_6998,N_6803);
and U7087 (N_7087,N_6612,N_6624);
nor U7088 (N_7088,N_6592,N_6836);
xnor U7089 (N_7089,N_6634,N_6580);
xor U7090 (N_7090,N_6945,N_6824);
and U7091 (N_7091,N_6771,N_6858);
xor U7092 (N_7092,N_6529,N_6801);
nor U7093 (N_7093,N_6586,N_6815);
nor U7094 (N_7094,N_6571,N_6874);
or U7095 (N_7095,N_6930,N_6626);
xnor U7096 (N_7096,N_6976,N_6773);
and U7097 (N_7097,N_6915,N_6526);
nor U7098 (N_7098,N_6994,N_6739);
or U7099 (N_7099,N_6889,N_6947);
or U7100 (N_7100,N_6563,N_6798);
nor U7101 (N_7101,N_6695,N_6934);
nor U7102 (N_7102,N_6750,N_6986);
or U7103 (N_7103,N_6942,N_6735);
nor U7104 (N_7104,N_6792,N_6656);
nor U7105 (N_7105,N_6729,N_6657);
nand U7106 (N_7106,N_6717,N_6875);
and U7107 (N_7107,N_6618,N_6772);
nand U7108 (N_7108,N_6823,N_6630);
nand U7109 (N_7109,N_6582,N_6608);
nor U7110 (N_7110,N_6977,N_6638);
and U7111 (N_7111,N_6786,N_6704);
and U7112 (N_7112,N_6944,N_6982);
and U7113 (N_7113,N_6857,N_6775);
xor U7114 (N_7114,N_6924,N_6544);
nor U7115 (N_7115,N_6852,N_6527);
nand U7116 (N_7116,N_6751,N_6789);
nand U7117 (N_7117,N_6653,N_6590);
and U7118 (N_7118,N_6960,N_6672);
xnor U7119 (N_7119,N_6776,N_6699);
nor U7120 (N_7120,N_6941,N_6515);
or U7121 (N_7121,N_6927,N_6782);
xnor U7122 (N_7122,N_6501,N_6787);
nor U7123 (N_7123,N_6854,N_6838);
nor U7124 (N_7124,N_6607,N_6669);
xor U7125 (N_7125,N_6627,N_6597);
and U7126 (N_7126,N_6785,N_6605);
or U7127 (N_7127,N_6964,N_6744);
xor U7128 (N_7128,N_6646,N_6567);
and U7129 (N_7129,N_6671,N_6905);
xnor U7130 (N_7130,N_6596,N_6839);
nand U7131 (N_7131,N_6500,N_6999);
nor U7132 (N_7132,N_6675,N_6507);
nor U7133 (N_7133,N_6814,N_6677);
xnor U7134 (N_7134,N_6631,N_6659);
and U7135 (N_7135,N_6578,N_6769);
or U7136 (N_7136,N_6907,N_6660);
nor U7137 (N_7137,N_6558,N_6655);
nand U7138 (N_7138,N_6665,N_6834);
nor U7139 (N_7139,N_6674,N_6518);
and U7140 (N_7140,N_6587,N_6689);
or U7141 (N_7141,N_6768,N_6628);
or U7142 (N_7142,N_6532,N_6707);
or U7143 (N_7143,N_6661,N_6740);
nand U7144 (N_7144,N_6892,N_6540);
xnor U7145 (N_7145,N_6728,N_6822);
nor U7146 (N_7146,N_6810,N_6579);
and U7147 (N_7147,N_6868,N_6837);
and U7148 (N_7148,N_6962,N_6514);
or U7149 (N_7149,N_6531,N_6777);
and U7150 (N_7150,N_6935,N_6951);
nor U7151 (N_7151,N_6993,N_6820);
xnor U7152 (N_7152,N_6911,N_6871);
or U7153 (N_7153,N_6560,N_6687);
or U7154 (N_7154,N_6970,N_6995);
or U7155 (N_7155,N_6635,N_6685);
nor U7156 (N_7156,N_6708,N_6863);
and U7157 (N_7157,N_6554,N_6929);
or U7158 (N_7158,N_6829,N_6758);
nor U7159 (N_7159,N_6594,N_6843);
and U7160 (N_7160,N_6840,N_6869);
nand U7161 (N_7161,N_6992,N_6673);
or U7162 (N_7162,N_6943,N_6818);
nor U7163 (N_7163,N_6745,N_6599);
and U7164 (N_7164,N_6644,N_6860);
and U7165 (N_7165,N_6676,N_6972);
xnor U7166 (N_7166,N_6602,N_6763);
nor U7167 (N_7167,N_6570,N_6748);
xnor U7168 (N_7168,N_6895,N_6666);
xor U7169 (N_7169,N_6581,N_6539);
or U7170 (N_7170,N_6808,N_6731);
nand U7171 (N_7171,N_6654,N_6719);
nor U7172 (N_7172,N_6766,N_6996);
nand U7173 (N_7173,N_6668,N_6809);
xor U7174 (N_7174,N_6513,N_6535);
nor U7175 (N_7175,N_6547,N_6906);
nor U7176 (N_7176,N_6856,N_6606);
and U7177 (N_7177,N_6973,N_6928);
and U7178 (N_7178,N_6981,N_6503);
nand U7179 (N_7179,N_6505,N_6714);
and U7180 (N_7180,N_6642,N_6788);
and U7181 (N_7181,N_6954,N_6693);
xor U7182 (N_7182,N_6713,N_6650);
xnor U7183 (N_7183,N_6797,N_6885);
nor U7184 (N_7184,N_6611,N_6952);
nand U7185 (N_7185,N_6574,N_6565);
nor U7186 (N_7186,N_6530,N_6710);
xor U7187 (N_7187,N_6920,N_6572);
xor U7188 (N_7188,N_6575,N_6884);
or U7189 (N_7189,N_6764,N_6738);
nor U7190 (N_7190,N_6755,N_6932);
nor U7191 (N_7191,N_6903,N_6556);
or U7192 (N_7192,N_6610,N_6747);
or U7193 (N_7193,N_6853,N_6784);
or U7194 (N_7194,N_6538,N_6559);
and U7195 (N_7195,N_6969,N_6730);
xor U7196 (N_7196,N_6555,N_6901);
nor U7197 (N_7197,N_6542,N_6583);
xnor U7198 (N_7198,N_6524,N_6967);
and U7199 (N_7199,N_6741,N_6541);
xnor U7200 (N_7200,N_6790,N_6794);
nand U7201 (N_7201,N_6752,N_6974);
and U7202 (N_7202,N_6761,N_6865);
xor U7203 (N_7203,N_6897,N_6828);
and U7204 (N_7204,N_6916,N_6870);
and U7205 (N_7205,N_6878,N_6667);
nand U7206 (N_7206,N_6569,N_6723);
nand U7207 (N_7207,N_6557,N_6975);
or U7208 (N_7208,N_6819,N_6806);
nand U7209 (N_7209,N_6686,N_6576);
nand U7210 (N_7210,N_6765,N_6502);
or U7211 (N_7211,N_6658,N_6997);
xnor U7212 (N_7212,N_6679,N_6896);
and U7213 (N_7213,N_6651,N_6616);
and U7214 (N_7214,N_6525,N_6844);
xor U7215 (N_7215,N_6774,N_6690);
and U7216 (N_7216,N_6584,N_6946);
nand U7217 (N_7217,N_6715,N_6926);
xnor U7218 (N_7218,N_6988,N_6528);
nand U7219 (N_7219,N_6568,N_6963);
nand U7220 (N_7220,N_6698,N_6830);
xor U7221 (N_7221,N_6811,N_6800);
nor U7222 (N_7222,N_6910,N_6851);
and U7223 (N_7223,N_6949,N_6718);
nand U7224 (N_7224,N_6562,N_6847);
and U7225 (N_7225,N_6817,N_6845);
nor U7226 (N_7226,N_6864,N_6553);
and U7227 (N_7227,N_6691,N_6757);
nand U7228 (N_7228,N_6662,N_6957);
nor U7229 (N_7229,N_6873,N_6700);
nand U7230 (N_7230,N_6678,N_6615);
nand U7231 (N_7231,N_6711,N_6795);
and U7232 (N_7232,N_6509,N_6850);
nand U7233 (N_7233,N_6812,N_6899);
and U7234 (N_7234,N_6939,N_6985);
nand U7235 (N_7235,N_6601,N_6548);
or U7236 (N_7236,N_6898,N_6825);
or U7237 (N_7237,N_6649,N_6912);
nor U7238 (N_7238,N_6536,N_6876);
nand U7239 (N_7239,N_6846,N_6979);
nand U7240 (N_7240,N_6511,N_6816);
nand U7241 (N_7241,N_6702,N_6948);
and U7242 (N_7242,N_6966,N_6598);
or U7243 (N_7243,N_6894,N_6923);
and U7244 (N_7244,N_6925,N_6883);
nand U7245 (N_7245,N_6683,N_6866);
nor U7246 (N_7246,N_6510,N_6770);
xnor U7247 (N_7247,N_6712,N_6591);
nor U7248 (N_7248,N_6965,N_6983);
and U7249 (N_7249,N_6561,N_6629);
and U7250 (N_7250,N_6971,N_6504);
nand U7251 (N_7251,N_6879,N_6820);
and U7252 (N_7252,N_6874,N_6617);
xnor U7253 (N_7253,N_6786,N_6822);
or U7254 (N_7254,N_6925,N_6609);
xnor U7255 (N_7255,N_6609,N_6949);
nand U7256 (N_7256,N_6940,N_6904);
nand U7257 (N_7257,N_6885,N_6990);
or U7258 (N_7258,N_6690,N_6839);
nand U7259 (N_7259,N_6566,N_6578);
xor U7260 (N_7260,N_6578,N_6559);
xor U7261 (N_7261,N_6772,N_6918);
xnor U7262 (N_7262,N_6588,N_6647);
nor U7263 (N_7263,N_6606,N_6540);
and U7264 (N_7264,N_6578,N_6625);
nor U7265 (N_7265,N_6892,N_6914);
or U7266 (N_7266,N_6604,N_6972);
and U7267 (N_7267,N_6563,N_6652);
or U7268 (N_7268,N_6746,N_6971);
nor U7269 (N_7269,N_6649,N_6687);
nor U7270 (N_7270,N_6745,N_6539);
and U7271 (N_7271,N_6899,N_6648);
nor U7272 (N_7272,N_6814,N_6795);
nand U7273 (N_7273,N_6819,N_6691);
nand U7274 (N_7274,N_6836,N_6882);
xor U7275 (N_7275,N_6727,N_6503);
or U7276 (N_7276,N_6857,N_6518);
nor U7277 (N_7277,N_6906,N_6849);
and U7278 (N_7278,N_6899,N_6978);
xor U7279 (N_7279,N_6912,N_6691);
or U7280 (N_7280,N_6702,N_6503);
nand U7281 (N_7281,N_6801,N_6558);
nor U7282 (N_7282,N_6913,N_6576);
nand U7283 (N_7283,N_6671,N_6900);
xor U7284 (N_7284,N_6861,N_6561);
nand U7285 (N_7285,N_6905,N_6513);
and U7286 (N_7286,N_6633,N_6792);
and U7287 (N_7287,N_6548,N_6694);
nand U7288 (N_7288,N_6949,N_6523);
nand U7289 (N_7289,N_6715,N_6923);
or U7290 (N_7290,N_6920,N_6511);
nor U7291 (N_7291,N_6992,N_6568);
or U7292 (N_7292,N_6932,N_6652);
nand U7293 (N_7293,N_6840,N_6606);
and U7294 (N_7294,N_6599,N_6784);
nand U7295 (N_7295,N_6743,N_6604);
nand U7296 (N_7296,N_6718,N_6848);
nor U7297 (N_7297,N_6982,N_6888);
nand U7298 (N_7298,N_6872,N_6902);
nand U7299 (N_7299,N_6704,N_6649);
nand U7300 (N_7300,N_6846,N_6851);
and U7301 (N_7301,N_6938,N_6989);
xor U7302 (N_7302,N_6962,N_6661);
or U7303 (N_7303,N_6613,N_6832);
nand U7304 (N_7304,N_6812,N_6570);
nand U7305 (N_7305,N_6980,N_6967);
xor U7306 (N_7306,N_6886,N_6922);
and U7307 (N_7307,N_6560,N_6816);
nor U7308 (N_7308,N_6789,N_6501);
or U7309 (N_7309,N_6710,N_6620);
and U7310 (N_7310,N_6903,N_6770);
nor U7311 (N_7311,N_6816,N_6630);
nor U7312 (N_7312,N_6905,N_6980);
nor U7313 (N_7313,N_6671,N_6946);
nand U7314 (N_7314,N_6875,N_6649);
and U7315 (N_7315,N_6507,N_6938);
nand U7316 (N_7316,N_6583,N_6930);
xor U7317 (N_7317,N_6501,N_6589);
nand U7318 (N_7318,N_6552,N_6616);
or U7319 (N_7319,N_6915,N_6985);
xnor U7320 (N_7320,N_6577,N_6881);
nor U7321 (N_7321,N_6548,N_6678);
or U7322 (N_7322,N_6521,N_6970);
xor U7323 (N_7323,N_6953,N_6947);
xor U7324 (N_7324,N_6506,N_6742);
xnor U7325 (N_7325,N_6913,N_6927);
xor U7326 (N_7326,N_6977,N_6585);
and U7327 (N_7327,N_6615,N_6913);
nor U7328 (N_7328,N_6629,N_6615);
and U7329 (N_7329,N_6936,N_6545);
and U7330 (N_7330,N_6761,N_6682);
nand U7331 (N_7331,N_6771,N_6643);
nand U7332 (N_7332,N_6581,N_6556);
nor U7333 (N_7333,N_6660,N_6786);
xor U7334 (N_7334,N_6973,N_6888);
nand U7335 (N_7335,N_6556,N_6851);
and U7336 (N_7336,N_6772,N_6508);
xor U7337 (N_7337,N_6696,N_6782);
nand U7338 (N_7338,N_6680,N_6643);
xor U7339 (N_7339,N_6560,N_6954);
nor U7340 (N_7340,N_6861,N_6633);
or U7341 (N_7341,N_6986,N_6692);
xnor U7342 (N_7342,N_6745,N_6834);
or U7343 (N_7343,N_6800,N_6757);
and U7344 (N_7344,N_6598,N_6702);
nand U7345 (N_7345,N_6691,N_6821);
nor U7346 (N_7346,N_6712,N_6988);
and U7347 (N_7347,N_6623,N_6864);
or U7348 (N_7348,N_6658,N_6728);
or U7349 (N_7349,N_6960,N_6512);
xor U7350 (N_7350,N_6686,N_6973);
nor U7351 (N_7351,N_6670,N_6932);
nand U7352 (N_7352,N_6685,N_6990);
nor U7353 (N_7353,N_6983,N_6891);
nor U7354 (N_7354,N_6778,N_6877);
nor U7355 (N_7355,N_6768,N_6547);
xor U7356 (N_7356,N_6546,N_6556);
xnor U7357 (N_7357,N_6922,N_6784);
nor U7358 (N_7358,N_6681,N_6847);
xnor U7359 (N_7359,N_6746,N_6796);
nand U7360 (N_7360,N_6529,N_6882);
or U7361 (N_7361,N_6953,N_6832);
nor U7362 (N_7362,N_6828,N_6532);
xnor U7363 (N_7363,N_6587,N_6512);
and U7364 (N_7364,N_6636,N_6646);
nor U7365 (N_7365,N_6688,N_6750);
nand U7366 (N_7366,N_6946,N_6742);
or U7367 (N_7367,N_6612,N_6844);
or U7368 (N_7368,N_6576,N_6805);
xnor U7369 (N_7369,N_6949,N_6923);
and U7370 (N_7370,N_6718,N_6628);
nor U7371 (N_7371,N_6895,N_6726);
nor U7372 (N_7372,N_6641,N_6683);
and U7373 (N_7373,N_6713,N_6865);
xor U7374 (N_7374,N_6610,N_6837);
xor U7375 (N_7375,N_6966,N_6750);
nor U7376 (N_7376,N_6601,N_6810);
xnor U7377 (N_7377,N_6755,N_6837);
and U7378 (N_7378,N_6595,N_6827);
and U7379 (N_7379,N_6732,N_6640);
and U7380 (N_7380,N_6649,N_6921);
nand U7381 (N_7381,N_6574,N_6857);
or U7382 (N_7382,N_6937,N_6638);
nor U7383 (N_7383,N_6820,N_6754);
nor U7384 (N_7384,N_6940,N_6692);
nor U7385 (N_7385,N_6728,N_6614);
nand U7386 (N_7386,N_6865,N_6773);
and U7387 (N_7387,N_6514,N_6638);
xnor U7388 (N_7388,N_6662,N_6773);
nor U7389 (N_7389,N_6552,N_6979);
nor U7390 (N_7390,N_6611,N_6523);
nand U7391 (N_7391,N_6759,N_6673);
nor U7392 (N_7392,N_6660,N_6628);
nand U7393 (N_7393,N_6830,N_6600);
or U7394 (N_7394,N_6623,N_6924);
nand U7395 (N_7395,N_6608,N_6996);
and U7396 (N_7396,N_6717,N_6804);
xnor U7397 (N_7397,N_6613,N_6798);
nor U7398 (N_7398,N_6981,N_6510);
or U7399 (N_7399,N_6618,N_6919);
nor U7400 (N_7400,N_6746,N_6808);
or U7401 (N_7401,N_6669,N_6589);
nor U7402 (N_7402,N_6577,N_6940);
xnor U7403 (N_7403,N_6636,N_6508);
nor U7404 (N_7404,N_6514,N_6720);
nand U7405 (N_7405,N_6543,N_6510);
nand U7406 (N_7406,N_6522,N_6769);
or U7407 (N_7407,N_6704,N_6511);
nand U7408 (N_7408,N_6779,N_6806);
nand U7409 (N_7409,N_6749,N_6733);
xor U7410 (N_7410,N_6549,N_6895);
and U7411 (N_7411,N_6612,N_6972);
nor U7412 (N_7412,N_6558,N_6860);
nor U7413 (N_7413,N_6659,N_6567);
xor U7414 (N_7414,N_6727,N_6599);
nand U7415 (N_7415,N_6675,N_6641);
xor U7416 (N_7416,N_6549,N_6836);
or U7417 (N_7417,N_6886,N_6937);
nand U7418 (N_7418,N_6686,N_6759);
nor U7419 (N_7419,N_6893,N_6722);
nand U7420 (N_7420,N_6958,N_6692);
and U7421 (N_7421,N_6674,N_6591);
and U7422 (N_7422,N_6710,N_6600);
nand U7423 (N_7423,N_6505,N_6698);
xor U7424 (N_7424,N_6776,N_6879);
nand U7425 (N_7425,N_6500,N_6871);
nand U7426 (N_7426,N_6695,N_6655);
or U7427 (N_7427,N_6648,N_6804);
and U7428 (N_7428,N_6831,N_6575);
nor U7429 (N_7429,N_6770,N_6812);
or U7430 (N_7430,N_6981,N_6674);
or U7431 (N_7431,N_6643,N_6962);
xnor U7432 (N_7432,N_6790,N_6926);
or U7433 (N_7433,N_6795,N_6546);
nand U7434 (N_7434,N_6848,N_6851);
nor U7435 (N_7435,N_6845,N_6999);
nor U7436 (N_7436,N_6975,N_6522);
xor U7437 (N_7437,N_6553,N_6858);
or U7438 (N_7438,N_6772,N_6609);
nor U7439 (N_7439,N_6662,N_6600);
xnor U7440 (N_7440,N_6689,N_6872);
nand U7441 (N_7441,N_6587,N_6615);
nor U7442 (N_7442,N_6812,N_6643);
nand U7443 (N_7443,N_6717,N_6543);
nand U7444 (N_7444,N_6995,N_6961);
or U7445 (N_7445,N_6871,N_6898);
or U7446 (N_7446,N_6782,N_6800);
nor U7447 (N_7447,N_6872,N_6786);
xnor U7448 (N_7448,N_6902,N_6661);
or U7449 (N_7449,N_6606,N_6512);
and U7450 (N_7450,N_6645,N_6903);
nor U7451 (N_7451,N_6688,N_6811);
nand U7452 (N_7452,N_6865,N_6859);
and U7453 (N_7453,N_6842,N_6589);
nand U7454 (N_7454,N_6896,N_6985);
or U7455 (N_7455,N_6681,N_6502);
or U7456 (N_7456,N_6881,N_6830);
xnor U7457 (N_7457,N_6646,N_6684);
and U7458 (N_7458,N_6692,N_6918);
xnor U7459 (N_7459,N_6822,N_6764);
or U7460 (N_7460,N_6816,N_6855);
xor U7461 (N_7461,N_6760,N_6521);
or U7462 (N_7462,N_6841,N_6857);
nor U7463 (N_7463,N_6840,N_6835);
and U7464 (N_7464,N_6811,N_6585);
nand U7465 (N_7465,N_6925,N_6900);
nor U7466 (N_7466,N_6798,N_6600);
xor U7467 (N_7467,N_6819,N_6958);
nor U7468 (N_7468,N_6510,N_6767);
xnor U7469 (N_7469,N_6522,N_6524);
nand U7470 (N_7470,N_6928,N_6689);
and U7471 (N_7471,N_6668,N_6813);
nand U7472 (N_7472,N_6697,N_6646);
xnor U7473 (N_7473,N_6895,N_6863);
and U7474 (N_7474,N_6927,N_6981);
nor U7475 (N_7475,N_6888,N_6612);
nor U7476 (N_7476,N_6696,N_6511);
and U7477 (N_7477,N_6591,N_6850);
or U7478 (N_7478,N_6897,N_6849);
nor U7479 (N_7479,N_6870,N_6707);
xnor U7480 (N_7480,N_6765,N_6609);
nor U7481 (N_7481,N_6666,N_6836);
and U7482 (N_7482,N_6680,N_6935);
and U7483 (N_7483,N_6664,N_6943);
or U7484 (N_7484,N_6667,N_6554);
nor U7485 (N_7485,N_6591,N_6539);
and U7486 (N_7486,N_6986,N_6742);
and U7487 (N_7487,N_6585,N_6966);
xor U7488 (N_7488,N_6666,N_6904);
nor U7489 (N_7489,N_6533,N_6712);
nor U7490 (N_7490,N_6772,N_6532);
xor U7491 (N_7491,N_6713,N_6768);
or U7492 (N_7492,N_6562,N_6733);
xor U7493 (N_7493,N_6896,N_6851);
or U7494 (N_7494,N_6669,N_6920);
and U7495 (N_7495,N_6866,N_6687);
nand U7496 (N_7496,N_6817,N_6901);
nor U7497 (N_7497,N_6926,N_6668);
xnor U7498 (N_7498,N_6610,N_6539);
nor U7499 (N_7499,N_6990,N_6804);
or U7500 (N_7500,N_7117,N_7441);
xnor U7501 (N_7501,N_7359,N_7433);
xor U7502 (N_7502,N_7130,N_7243);
nand U7503 (N_7503,N_7480,N_7279);
and U7504 (N_7504,N_7093,N_7255);
and U7505 (N_7505,N_7059,N_7244);
xnor U7506 (N_7506,N_7140,N_7457);
or U7507 (N_7507,N_7275,N_7110);
or U7508 (N_7508,N_7185,N_7377);
nand U7509 (N_7509,N_7455,N_7091);
or U7510 (N_7510,N_7467,N_7261);
or U7511 (N_7511,N_7021,N_7118);
or U7512 (N_7512,N_7425,N_7241);
nand U7513 (N_7513,N_7295,N_7344);
nand U7514 (N_7514,N_7389,N_7189);
xor U7515 (N_7515,N_7018,N_7342);
or U7516 (N_7516,N_7257,N_7019);
and U7517 (N_7517,N_7099,N_7168);
xor U7518 (N_7518,N_7149,N_7221);
nor U7519 (N_7519,N_7256,N_7408);
xnor U7520 (N_7520,N_7191,N_7379);
xnor U7521 (N_7521,N_7123,N_7006);
nor U7522 (N_7522,N_7495,N_7450);
and U7523 (N_7523,N_7042,N_7274);
nand U7524 (N_7524,N_7171,N_7430);
and U7525 (N_7525,N_7320,N_7054);
or U7526 (N_7526,N_7217,N_7356);
xnor U7527 (N_7527,N_7420,N_7324);
xor U7528 (N_7528,N_7090,N_7158);
xor U7529 (N_7529,N_7399,N_7415);
and U7530 (N_7530,N_7442,N_7025);
or U7531 (N_7531,N_7067,N_7013);
xnor U7532 (N_7532,N_7156,N_7134);
and U7533 (N_7533,N_7368,N_7406);
or U7534 (N_7534,N_7386,N_7499);
xnor U7535 (N_7535,N_7225,N_7174);
nor U7536 (N_7536,N_7456,N_7098);
or U7537 (N_7537,N_7066,N_7285);
xor U7538 (N_7538,N_7064,N_7086);
or U7539 (N_7539,N_7445,N_7082);
nor U7540 (N_7540,N_7112,N_7385);
nor U7541 (N_7541,N_7316,N_7001);
and U7542 (N_7542,N_7265,N_7203);
nor U7543 (N_7543,N_7313,N_7335);
nor U7544 (N_7544,N_7401,N_7372);
nand U7545 (N_7545,N_7052,N_7165);
nand U7546 (N_7546,N_7246,N_7286);
nand U7547 (N_7547,N_7057,N_7443);
and U7548 (N_7548,N_7062,N_7015);
and U7549 (N_7549,N_7383,N_7281);
xor U7550 (N_7550,N_7024,N_7014);
nor U7551 (N_7551,N_7230,N_7362);
and U7552 (N_7552,N_7376,N_7477);
or U7553 (N_7553,N_7249,N_7223);
and U7554 (N_7554,N_7143,N_7296);
and U7555 (N_7555,N_7426,N_7207);
or U7556 (N_7556,N_7459,N_7043);
nand U7557 (N_7557,N_7146,N_7188);
nand U7558 (N_7558,N_7475,N_7330);
or U7559 (N_7559,N_7163,N_7232);
and U7560 (N_7560,N_7229,N_7113);
or U7561 (N_7561,N_7097,N_7439);
nor U7562 (N_7562,N_7023,N_7002);
xnor U7563 (N_7563,N_7305,N_7226);
nor U7564 (N_7564,N_7254,N_7300);
nand U7565 (N_7565,N_7047,N_7291);
nor U7566 (N_7566,N_7150,N_7478);
and U7567 (N_7567,N_7051,N_7298);
and U7568 (N_7568,N_7120,N_7201);
xor U7569 (N_7569,N_7004,N_7186);
nand U7570 (N_7570,N_7107,N_7367);
xor U7571 (N_7571,N_7304,N_7370);
xor U7572 (N_7572,N_7284,N_7077);
or U7573 (N_7573,N_7205,N_7460);
xnor U7574 (N_7574,N_7045,N_7345);
xor U7575 (N_7575,N_7464,N_7483);
or U7576 (N_7576,N_7033,N_7227);
or U7577 (N_7577,N_7224,N_7144);
nand U7578 (N_7578,N_7032,N_7080);
or U7579 (N_7579,N_7177,N_7360);
nor U7580 (N_7580,N_7085,N_7253);
nand U7581 (N_7581,N_7343,N_7010);
xor U7582 (N_7582,N_7154,N_7179);
or U7583 (N_7583,N_7488,N_7105);
xnor U7584 (N_7584,N_7037,N_7103);
or U7585 (N_7585,N_7315,N_7466);
nand U7586 (N_7586,N_7012,N_7096);
or U7587 (N_7587,N_7404,N_7136);
xor U7588 (N_7588,N_7327,N_7041);
and U7589 (N_7589,N_7178,N_7412);
and U7590 (N_7590,N_7382,N_7184);
or U7591 (N_7591,N_7322,N_7166);
or U7592 (N_7592,N_7092,N_7128);
xor U7593 (N_7593,N_7000,N_7473);
nand U7594 (N_7594,N_7282,N_7193);
and U7595 (N_7595,N_7454,N_7378);
and U7596 (N_7596,N_7469,N_7038);
or U7597 (N_7597,N_7381,N_7251);
and U7598 (N_7598,N_7369,N_7252);
and U7599 (N_7599,N_7468,N_7192);
nand U7600 (N_7600,N_7449,N_7338);
nor U7601 (N_7601,N_7310,N_7371);
and U7602 (N_7602,N_7159,N_7048);
xnor U7603 (N_7603,N_7169,N_7049);
xor U7604 (N_7604,N_7198,N_7462);
nand U7605 (N_7605,N_7273,N_7088);
and U7606 (N_7606,N_7352,N_7202);
nor U7607 (N_7607,N_7491,N_7164);
xnor U7608 (N_7608,N_7142,N_7361);
nor U7609 (N_7609,N_7476,N_7287);
xnor U7610 (N_7610,N_7312,N_7437);
xnor U7611 (N_7611,N_7108,N_7407);
and U7612 (N_7612,N_7061,N_7213);
and U7613 (N_7613,N_7470,N_7216);
xnor U7614 (N_7614,N_7109,N_7303);
nor U7615 (N_7615,N_7036,N_7280);
or U7616 (N_7616,N_7029,N_7182);
and U7617 (N_7617,N_7347,N_7497);
or U7618 (N_7618,N_7199,N_7239);
nand U7619 (N_7619,N_7436,N_7181);
nor U7620 (N_7620,N_7121,N_7325);
xnor U7621 (N_7621,N_7063,N_7250);
and U7622 (N_7622,N_7337,N_7214);
nor U7623 (N_7623,N_7209,N_7069);
nand U7624 (N_7624,N_7007,N_7231);
nand U7625 (N_7625,N_7487,N_7271);
nor U7626 (N_7626,N_7290,N_7292);
xor U7627 (N_7627,N_7114,N_7228);
or U7628 (N_7628,N_7272,N_7218);
nor U7629 (N_7629,N_7354,N_7152);
or U7630 (N_7630,N_7332,N_7314);
nor U7631 (N_7631,N_7263,N_7129);
nand U7632 (N_7632,N_7306,N_7486);
nor U7633 (N_7633,N_7268,N_7210);
or U7634 (N_7634,N_7329,N_7100);
nor U7635 (N_7635,N_7039,N_7180);
or U7636 (N_7636,N_7492,N_7339);
and U7637 (N_7637,N_7364,N_7471);
or U7638 (N_7638,N_7076,N_7073);
xor U7639 (N_7639,N_7060,N_7444);
xor U7640 (N_7640,N_7238,N_7390);
nand U7641 (N_7641,N_7133,N_7124);
nor U7642 (N_7642,N_7409,N_7183);
xnor U7643 (N_7643,N_7403,N_7440);
nand U7644 (N_7644,N_7333,N_7009);
xnor U7645 (N_7645,N_7242,N_7479);
xnor U7646 (N_7646,N_7206,N_7294);
and U7647 (N_7647,N_7266,N_7104);
xor U7648 (N_7648,N_7264,N_7490);
nand U7649 (N_7649,N_7204,N_7463);
xor U7650 (N_7650,N_7429,N_7396);
nor U7651 (N_7651,N_7391,N_7481);
or U7652 (N_7652,N_7482,N_7235);
or U7653 (N_7653,N_7167,N_7127);
xnor U7654 (N_7654,N_7299,N_7055);
nor U7655 (N_7655,N_7446,N_7358);
xor U7656 (N_7656,N_7432,N_7387);
nand U7657 (N_7657,N_7153,N_7035);
and U7658 (N_7658,N_7336,N_7340);
xnor U7659 (N_7659,N_7126,N_7119);
xor U7660 (N_7660,N_7289,N_7373);
nand U7661 (N_7661,N_7398,N_7212);
nor U7662 (N_7662,N_7138,N_7309);
and U7663 (N_7663,N_7031,N_7258);
xor U7664 (N_7664,N_7493,N_7068);
or U7665 (N_7665,N_7365,N_7276);
xnor U7666 (N_7666,N_7101,N_7366);
and U7667 (N_7667,N_7453,N_7451);
and U7668 (N_7668,N_7323,N_7245);
or U7669 (N_7669,N_7194,N_7438);
or U7670 (N_7670,N_7374,N_7157);
xnor U7671 (N_7671,N_7046,N_7219);
nor U7672 (N_7672,N_7116,N_7058);
or U7673 (N_7673,N_7106,N_7351);
nor U7674 (N_7674,N_7208,N_7416);
nor U7675 (N_7675,N_7195,N_7040);
xnor U7676 (N_7676,N_7317,N_7353);
nand U7677 (N_7677,N_7414,N_7115);
or U7678 (N_7678,N_7070,N_7075);
and U7679 (N_7679,N_7259,N_7034);
and U7680 (N_7680,N_7418,N_7355);
nor U7681 (N_7681,N_7394,N_7050);
nand U7682 (N_7682,N_7079,N_7461);
xnor U7683 (N_7683,N_7084,N_7111);
xor U7684 (N_7684,N_7301,N_7003);
nor U7685 (N_7685,N_7147,N_7131);
or U7686 (N_7686,N_7222,N_7326);
and U7687 (N_7687,N_7405,N_7422);
and U7688 (N_7688,N_7392,N_7135);
nand U7689 (N_7689,N_7078,N_7465);
nand U7690 (N_7690,N_7005,N_7044);
nor U7691 (N_7691,N_7160,N_7419);
and U7692 (N_7692,N_7411,N_7400);
xnor U7693 (N_7693,N_7237,N_7233);
and U7694 (N_7694,N_7485,N_7056);
and U7695 (N_7695,N_7122,N_7087);
xnor U7696 (N_7696,N_7155,N_7176);
or U7697 (N_7697,N_7262,N_7341);
or U7698 (N_7698,N_7236,N_7065);
nand U7699 (N_7699,N_7270,N_7318);
or U7700 (N_7700,N_7278,N_7145);
nor U7701 (N_7701,N_7071,N_7248);
and U7702 (N_7702,N_7494,N_7072);
and U7703 (N_7703,N_7027,N_7190);
nand U7704 (N_7704,N_7132,N_7346);
nand U7705 (N_7705,N_7020,N_7200);
xor U7706 (N_7706,N_7402,N_7197);
and U7707 (N_7707,N_7348,N_7269);
nor U7708 (N_7708,N_7331,N_7173);
xor U7709 (N_7709,N_7410,N_7074);
nor U7710 (N_7710,N_7447,N_7102);
xnor U7711 (N_7711,N_7267,N_7388);
and U7712 (N_7712,N_7375,N_7139);
xor U7713 (N_7713,N_7452,N_7260);
and U7714 (N_7714,N_7175,N_7008);
nand U7715 (N_7715,N_7125,N_7170);
and U7716 (N_7716,N_7288,N_7094);
nor U7717 (N_7717,N_7431,N_7172);
nor U7718 (N_7718,N_7215,N_7363);
nor U7719 (N_7719,N_7081,N_7384);
and U7720 (N_7720,N_7417,N_7297);
or U7721 (N_7721,N_7283,N_7293);
nor U7722 (N_7722,N_7307,N_7161);
or U7723 (N_7723,N_7141,N_7240);
or U7724 (N_7724,N_7095,N_7395);
or U7725 (N_7725,N_7421,N_7397);
nor U7726 (N_7726,N_7247,N_7427);
nor U7727 (N_7727,N_7137,N_7302);
nand U7728 (N_7728,N_7380,N_7393);
nand U7729 (N_7729,N_7328,N_7349);
and U7730 (N_7730,N_7448,N_7413);
and U7731 (N_7731,N_7308,N_7350);
or U7732 (N_7732,N_7277,N_7089);
nand U7733 (N_7733,N_7162,N_7472);
or U7734 (N_7734,N_7424,N_7498);
or U7735 (N_7735,N_7028,N_7334);
xnor U7736 (N_7736,N_7321,N_7053);
xor U7737 (N_7737,N_7474,N_7428);
and U7738 (N_7738,N_7026,N_7083);
or U7739 (N_7739,N_7211,N_7187);
nor U7740 (N_7740,N_7489,N_7434);
or U7741 (N_7741,N_7220,N_7423);
and U7742 (N_7742,N_7011,N_7458);
nand U7743 (N_7743,N_7435,N_7016);
nor U7744 (N_7744,N_7357,N_7151);
nand U7745 (N_7745,N_7148,N_7496);
xnor U7746 (N_7746,N_7234,N_7030);
and U7747 (N_7747,N_7484,N_7017);
or U7748 (N_7748,N_7196,N_7022);
nor U7749 (N_7749,N_7311,N_7319);
and U7750 (N_7750,N_7132,N_7450);
xnor U7751 (N_7751,N_7472,N_7388);
and U7752 (N_7752,N_7202,N_7260);
or U7753 (N_7753,N_7100,N_7392);
nor U7754 (N_7754,N_7018,N_7095);
nor U7755 (N_7755,N_7457,N_7119);
and U7756 (N_7756,N_7315,N_7121);
nand U7757 (N_7757,N_7113,N_7154);
and U7758 (N_7758,N_7471,N_7045);
xnor U7759 (N_7759,N_7088,N_7390);
xnor U7760 (N_7760,N_7233,N_7117);
and U7761 (N_7761,N_7203,N_7036);
nor U7762 (N_7762,N_7097,N_7356);
or U7763 (N_7763,N_7332,N_7213);
and U7764 (N_7764,N_7111,N_7002);
and U7765 (N_7765,N_7233,N_7122);
nor U7766 (N_7766,N_7388,N_7298);
nand U7767 (N_7767,N_7480,N_7006);
or U7768 (N_7768,N_7085,N_7164);
or U7769 (N_7769,N_7488,N_7370);
or U7770 (N_7770,N_7342,N_7044);
or U7771 (N_7771,N_7496,N_7263);
and U7772 (N_7772,N_7344,N_7260);
and U7773 (N_7773,N_7122,N_7435);
nand U7774 (N_7774,N_7356,N_7464);
or U7775 (N_7775,N_7425,N_7181);
nand U7776 (N_7776,N_7406,N_7001);
nor U7777 (N_7777,N_7125,N_7080);
xnor U7778 (N_7778,N_7069,N_7076);
xnor U7779 (N_7779,N_7238,N_7034);
and U7780 (N_7780,N_7355,N_7277);
xor U7781 (N_7781,N_7429,N_7189);
xnor U7782 (N_7782,N_7081,N_7122);
nand U7783 (N_7783,N_7357,N_7235);
xnor U7784 (N_7784,N_7453,N_7096);
and U7785 (N_7785,N_7073,N_7144);
nor U7786 (N_7786,N_7077,N_7455);
nand U7787 (N_7787,N_7070,N_7419);
xnor U7788 (N_7788,N_7285,N_7345);
or U7789 (N_7789,N_7114,N_7353);
and U7790 (N_7790,N_7070,N_7234);
and U7791 (N_7791,N_7040,N_7395);
nor U7792 (N_7792,N_7480,N_7162);
nand U7793 (N_7793,N_7297,N_7102);
nand U7794 (N_7794,N_7450,N_7086);
xor U7795 (N_7795,N_7022,N_7484);
nor U7796 (N_7796,N_7456,N_7270);
and U7797 (N_7797,N_7311,N_7183);
or U7798 (N_7798,N_7199,N_7036);
nand U7799 (N_7799,N_7001,N_7203);
and U7800 (N_7800,N_7392,N_7276);
nand U7801 (N_7801,N_7160,N_7330);
nand U7802 (N_7802,N_7265,N_7123);
xnor U7803 (N_7803,N_7432,N_7410);
and U7804 (N_7804,N_7190,N_7217);
xor U7805 (N_7805,N_7134,N_7344);
nand U7806 (N_7806,N_7286,N_7150);
xnor U7807 (N_7807,N_7018,N_7308);
xnor U7808 (N_7808,N_7379,N_7133);
and U7809 (N_7809,N_7227,N_7413);
nand U7810 (N_7810,N_7455,N_7368);
and U7811 (N_7811,N_7414,N_7066);
or U7812 (N_7812,N_7058,N_7208);
and U7813 (N_7813,N_7257,N_7127);
xor U7814 (N_7814,N_7201,N_7484);
nand U7815 (N_7815,N_7243,N_7254);
and U7816 (N_7816,N_7096,N_7047);
or U7817 (N_7817,N_7492,N_7029);
nor U7818 (N_7818,N_7260,N_7103);
or U7819 (N_7819,N_7348,N_7171);
and U7820 (N_7820,N_7294,N_7088);
xnor U7821 (N_7821,N_7374,N_7421);
or U7822 (N_7822,N_7341,N_7193);
and U7823 (N_7823,N_7376,N_7452);
and U7824 (N_7824,N_7060,N_7367);
nor U7825 (N_7825,N_7257,N_7252);
and U7826 (N_7826,N_7107,N_7324);
and U7827 (N_7827,N_7190,N_7362);
nor U7828 (N_7828,N_7009,N_7145);
nand U7829 (N_7829,N_7489,N_7080);
or U7830 (N_7830,N_7418,N_7270);
nand U7831 (N_7831,N_7128,N_7174);
nand U7832 (N_7832,N_7449,N_7152);
nor U7833 (N_7833,N_7158,N_7061);
nand U7834 (N_7834,N_7246,N_7005);
nand U7835 (N_7835,N_7174,N_7078);
and U7836 (N_7836,N_7336,N_7459);
nor U7837 (N_7837,N_7000,N_7011);
or U7838 (N_7838,N_7057,N_7051);
nor U7839 (N_7839,N_7110,N_7485);
xor U7840 (N_7840,N_7354,N_7189);
or U7841 (N_7841,N_7434,N_7242);
and U7842 (N_7842,N_7318,N_7174);
and U7843 (N_7843,N_7336,N_7065);
and U7844 (N_7844,N_7405,N_7481);
or U7845 (N_7845,N_7364,N_7367);
xor U7846 (N_7846,N_7073,N_7283);
nand U7847 (N_7847,N_7282,N_7244);
xnor U7848 (N_7848,N_7079,N_7236);
nand U7849 (N_7849,N_7093,N_7261);
nor U7850 (N_7850,N_7190,N_7392);
nor U7851 (N_7851,N_7116,N_7066);
or U7852 (N_7852,N_7005,N_7449);
and U7853 (N_7853,N_7304,N_7383);
xnor U7854 (N_7854,N_7130,N_7027);
or U7855 (N_7855,N_7262,N_7453);
and U7856 (N_7856,N_7065,N_7251);
nor U7857 (N_7857,N_7413,N_7486);
xor U7858 (N_7858,N_7063,N_7326);
and U7859 (N_7859,N_7072,N_7273);
or U7860 (N_7860,N_7320,N_7116);
or U7861 (N_7861,N_7302,N_7366);
or U7862 (N_7862,N_7097,N_7137);
or U7863 (N_7863,N_7070,N_7079);
nand U7864 (N_7864,N_7436,N_7311);
nor U7865 (N_7865,N_7072,N_7081);
nor U7866 (N_7866,N_7183,N_7282);
or U7867 (N_7867,N_7340,N_7212);
nand U7868 (N_7868,N_7308,N_7473);
and U7869 (N_7869,N_7451,N_7318);
nor U7870 (N_7870,N_7126,N_7320);
and U7871 (N_7871,N_7034,N_7393);
nand U7872 (N_7872,N_7273,N_7124);
nor U7873 (N_7873,N_7401,N_7190);
nand U7874 (N_7874,N_7391,N_7420);
or U7875 (N_7875,N_7428,N_7218);
xnor U7876 (N_7876,N_7114,N_7343);
or U7877 (N_7877,N_7073,N_7413);
nor U7878 (N_7878,N_7455,N_7335);
nand U7879 (N_7879,N_7100,N_7328);
or U7880 (N_7880,N_7070,N_7336);
and U7881 (N_7881,N_7031,N_7369);
nor U7882 (N_7882,N_7249,N_7142);
nor U7883 (N_7883,N_7146,N_7294);
nor U7884 (N_7884,N_7415,N_7491);
xnor U7885 (N_7885,N_7446,N_7310);
xor U7886 (N_7886,N_7350,N_7096);
nand U7887 (N_7887,N_7091,N_7316);
xnor U7888 (N_7888,N_7447,N_7481);
and U7889 (N_7889,N_7166,N_7228);
nor U7890 (N_7890,N_7220,N_7164);
nor U7891 (N_7891,N_7231,N_7380);
nand U7892 (N_7892,N_7368,N_7193);
and U7893 (N_7893,N_7460,N_7214);
and U7894 (N_7894,N_7193,N_7034);
and U7895 (N_7895,N_7263,N_7451);
xor U7896 (N_7896,N_7358,N_7420);
or U7897 (N_7897,N_7345,N_7191);
or U7898 (N_7898,N_7225,N_7269);
and U7899 (N_7899,N_7455,N_7089);
xor U7900 (N_7900,N_7277,N_7000);
xnor U7901 (N_7901,N_7036,N_7147);
and U7902 (N_7902,N_7448,N_7376);
xnor U7903 (N_7903,N_7278,N_7259);
nand U7904 (N_7904,N_7109,N_7445);
or U7905 (N_7905,N_7287,N_7471);
and U7906 (N_7906,N_7417,N_7106);
nand U7907 (N_7907,N_7466,N_7006);
or U7908 (N_7908,N_7401,N_7048);
nor U7909 (N_7909,N_7154,N_7047);
or U7910 (N_7910,N_7321,N_7281);
nand U7911 (N_7911,N_7044,N_7443);
or U7912 (N_7912,N_7422,N_7013);
xnor U7913 (N_7913,N_7457,N_7046);
nand U7914 (N_7914,N_7472,N_7068);
nand U7915 (N_7915,N_7280,N_7108);
and U7916 (N_7916,N_7084,N_7298);
and U7917 (N_7917,N_7193,N_7083);
and U7918 (N_7918,N_7213,N_7142);
nand U7919 (N_7919,N_7064,N_7439);
xnor U7920 (N_7920,N_7284,N_7321);
or U7921 (N_7921,N_7273,N_7062);
or U7922 (N_7922,N_7093,N_7410);
or U7923 (N_7923,N_7253,N_7321);
xnor U7924 (N_7924,N_7302,N_7313);
nor U7925 (N_7925,N_7405,N_7289);
nor U7926 (N_7926,N_7355,N_7382);
nand U7927 (N_7927,N_7045,N_7489);
xnor U7928 (N_7928,N_7082,N_7105);
xnor U7929 (N_7929,N_7052,N_7446);
and U7930 (N_7930,N_7027,N_7006);
nor U7931 (N_7931,N_7200,N_7001);
nor U7932 (N_7932,N_7247,N_7354);
xnor U7933 (N_7933,N_7218,N_7424);
and U7934 (N_7934,N_7429,N_7223);
xnor U7935 (N_7935,N_7326,N_7218);
or U7936 (N_7936,N_7417,N_7375);
xnor U7937 (N_7937,N_7305,N_7023);
or U7938 (N_7938,N_7116,N_7063);
nor U7939 (N_7939,N_7453,N_7432);
or U7940 (N_7940,N_7336,N_7305);
or U7941 (N_7941,N_7341,N_7051);
and U7942 (N_7942,N_7115,N_7491);
and U7943 (N_7943,N_7106,N_7038);
nand U7944 (N_7944,N_7488,N_7478);
nor U7945 (N_7945,N_7442,N_7086);
and U7946 (N_7946,N_7284,N_7067);
or U7947 (N_7947,N_7375,N_7278);
or U7948 (N_7948,N_7428,N_7084);
or U7949 (N_7949,N_7203,N_7279);
nand U7950 (N_7950,N_7324,N_7464);
or U7951 (N_7951,N_7279,N_7267);
and U7952 (N_7952,N_7419,N_7115);
nand U7953 (N_7953,N_7047,N_7199);
and U7954 (N_7954,N_7160,N_7071);
and U7955 (N_7955,N_7027,N_7034);
xor U7956 (N_7956,N_7466,N_7340);
nor U7957 (N_7957,N_7486,N_7183);
or U7958 (N_7958,N_7017,N_7364);
xor U7959 (N_7959,N_7261,N_7476);
nor U7960 (N_7960,N_7476,N_7032);
nand U7961 (N_7961,N_7104,N_7365);
or U7962 (N_7962,N_7072,N_7088);
nor U7963 (N_7963,N_7453,N_7031);
and U7964 (N_7964,N_7303,N_7220);
and U7965 (N_7965,N_7060,N_7012);
nor U7966 (N_7966,N_7450,N_7390);
or U7967 (N_7967,N_7076,N_7066);
and U7968 (N_7968,N_7322,N_7068);
xnor U7969 (N_7969,N_7135,N_7260);
or U7970 (N_7970,N_7017,N_7049);
or U7971 (N_7971,N_7269,N_7356);
or U7972 (N_7972,N_7012,N_7179);
nor U7973 (N_7973,N_7073,N_7027);
or U7974 (N_7974,N_7432,N_7279);
and U7975 (N_7975,N_7239,N_7435);
nand U7976 (N_7976,N_7459,N_7231);
xor U7977 (N_7977,N_7028,N_7073);
nand U7978 (N_7978,N_7058,N_7486);
and U7979 (N_7979,N_7318,N_7105);
xor U7980 (N_7980,N_7004,N_7018);
and U7981 (N_7981,N_7378,N_7499);
xnor U7982 (N_7982,N_7313,N_7324);
or U7983 (N_7983,N_7299,N_7051);
and U7984 (N_7984,N_7122,N_7263);
nor U7985 (N_7985,N_7050,N_7324);
nand U7986 (N_7986,N_7491,N_7048);
nor U7987 (N_7987,N_7403,N_7412);
nand U7988 (N_7988,N_7010,N_7270);
nor U7989 (N_7989,N_7098,N_7282);
xor U7990 (N_7990,N_7112,N_7173);
xnor U7991 (N_7991,N_7258,N_7262);
nor U7992 (N_7992,N_7196,N_7444);
or U7993 (N_7993,N_7320,N_7175);
nor U7994 (N_7994,N_7223,N_7268);
or U7995 (N_7995,N_7262,N_7445);
xor U7996 (N_7996,N_7159,N_7282);
and U7997 (N_7997,N_7206,N_7189);
xnor U7998 (N_7998,N_7377,N_7097);
nor U7999 (N_7999,N_7215,N_7200);
and U8000 (N_8000,N_7830,N_7514);
nor U8001 (N_8001,N_7829,N_7803);
or U8002 (N_8002,N_7978,N_7546);
nor U8003 (N_8003,N_7598,N_7763);
and U8004 (N_8004,N_7854,N_7714);
xor U8005 (N_8005,N_7729,N_7739);
xnor U8006 (N_8006,N_7954,N_7879);
and U8007 (N_8007,N_7716,N_7826);
and U8008 (N_8008,N_7755,N_7757);
nor U8009 (N_8009,N_7635,N_7975);
nor U8010 (N_8010,N_7977,N_7562);
nand U8011 (N_8011,N_7528,N_7580);
xor U8012 (N_8012,N_7797,N_7605);
or U8013 (N_8013,N_7929,N_7523);
xnor U8014 (N_8014,N_7502,N_7666);
nor U8015 (N_8015,N_7615,N_7744);
nand U8016 (N_8016,N_7548,N_7821);
nand U8017 (N_8017,N_7708,N_7509);
nor U8018 (N_8018,N_7983,N_7779);
xor U8019 (N_8019,N_7727,N_7815);
xor U8020 (N_8020,N_7599,N_7754);
and U8021 (N_8021,N_7525,N_7658);
or U8022 (N_8022,N_7642,N_7655);
or U8023 (N_8023,N_7623,N_7973);
nand U8024 (N_8024,N_7993,N_7590);
or U8025 (N_8025,N_7967,N_7586);
nor U8026 (N_8026,N_7861,N_7909);
nor U8027 (N_8027,N_7802,N_7697);
xor U8028 (N_8028,N_7640,N_7971);
or U8029 (N_8029,N_7808,N_7933);
nor U8030 (N_8030,N_7520,N_7832);
xor U8031 (N_8031,N_7999,N_7908);
xnor U8032 (N_8032,N_7618,N_7902);
nor U8033 (N_8033,N_7750,N_7718);
or U8034 (N_8034,N_7917,N_7867);
xnor U8035 (N_8035,N_7606,N_7503);
nand U8036 (N_8036,N_7877,N_7787);
and U8037 (N_8037,N_7770,N_7588);
and U8038 (N_8038,N_7863,N_7646);
and U8039 (N_8039,N_7995,N_7573);
nor U8040 (N_8040,N_7532,N_7531);
and U8041 (N_8041,N_7799,N_7907);
and U8042 (N_8042,N_7989,N_7551);
or U8043 (N_8043,N_7912,N_7805);
xnor U8044 (N_8044,N_7741,N_7756);
nand U8045 (N_8045,N_7619,N_7880);
and U8046 (N_8046,N_7698,N_7506);
nor U8047 (N_8047,N_7883,N_7751);
nand U8048 (N_8048,N_7884,N_7679);
and U8049 (N_8049,N_7919,N_7682);
and U8050 (N_8050,N_7876,N_7875);
xor U8051 (N_8051,N_7809,N_7759);
nor U8052 (N_8052,N_7816,N_7602);
xnor U8053 (N_8053,N_7938,N_7935);
or U8054 (N_8054,N_7795,N_7539);
xor U8055 (N_8055,N_7864,N_7671);
nor U8056 (N_8056,N_7604,N_7699);
and U8057 (N_8057,N_7852,N_7637);
nand U8058 (N_8058,N_7540,N_7696);
xnor U8059 (N_8059,N_7676,N_7652);
nand U8060 (N_8060,N_7550,N_7984);
xor U8061 (N_8061,N_7774,N_7762);
and U8062 (N_8062,N_7846,N_7991);
and U8063 (N_8063,N_7567,N_7557);
nor U8064 (N_8064,N_7641,N_7510);
xnor U8065 (N_8065,N_7500,N_7994);
and U8066 (N_8066,N_7643,N_7703);
xnor U8067 (N_8067,N_7969,N_7616);
nor U8068 (N_8068,N_7898,N_7941);
nor U8069 (N_8069,N_7901,N_7847);
nand U8070 (N_8070,N_7656,N_7566);
and U8071 (N_8071,N_7841,N_7626);
and U8072 (N_8072,N_7889,N_7530);
xor U8073 (N_8073,N_7951,N_7725);
nand U8074 (N_8074,N_7860,N_7800);
nand U8075 (N_8075,N_7801,N_7955);
nand U8076 (N_8076,N_7865,N_7845);
nand U8077 (N_8077,N_7786,N_7949);
and U8078 (N_8078,N_7625,N_7707);
nand U8079 (N_8079,N_7892,N_7743);
xor U8080 (N_8080,N_7813,N_7607);
xor U8081 (N_8081,N_7669,N_7900);
nor U8082 (N_8082,N_7851,N_7603);
nand U8083 (N_8083,N_7681,N_7819);
nor U8084 (N_8084,N_7638,N_7549);
nor U8085 (N_8085,N_7953,N_7674);
or U8086 (N_8086,N_7721,N_7897);
nor U8087 (N_8087,N_7715,N_7807);
nand U8088 (N_8088,N_7986,N_7632);
or U8089 (N_8089,N_7569,N_7577);
nor U8090 (N_8090,N_7517,N_7720);
nand U8091 (N_8091,N_7740,N_7584);
nand U8092 (N_8092,N_7613,N_7937);
xor U8093 (N_8093,N_7872,N_7524);
xnor U8094 (N_8094,N_7654,N_7960);
nand U8095 (N_8095,N_7910,N_7563);
xor U8096 (N_8096,N_7657,N_7776);
xor U8097 (N_8097,N_7747,N_7997);
nor U8098 (N_8098,N_7672,N_7559);
or U8099 (N_8099,N_7575,N_7628);
and U8100 (N_8100,N_7663,N_7622);
nand U8101 (N_8101,N_7952,N_7924);
and U8102 (N_8102,N_7527,N_7691);
or U8103 (N_8103,N_7630,N_7874);
and U8104 (N_8104,N_7782,N_7792);
nand U8105 (N_8105,N_7576,N_7677);
or U8106 (N_8106,N_7834,N_7585);
nor U8107 (N_8107,N_7796,N_7579);
xor U8108 (N_8108,N_7600,N_7581);
or U8109 (N_8109,N_7939,N_7695);
or U8110 (N_8110,N_7956,N_7869);
nand U8111 (N_8111,N_7928,N_7966);
nor U8112 (N_8112,N_7724,N_7752);
nand U8113 (N_8113,N_7890,N_7516);
and U8114 (N_8114,N_7634,N_7814);
nand U8115 (N_8115,N_7660,N_7988);
and U8116 (N_8116,N_7916,N_7645);
or U8117 (N_8117,N_7702,N_7649);
and U8118 (N_8118,N_7968,N_7849);
or U8119 (N_8119,N_7667,N_7781);
and U8120 (N_8120,N_7947,N_7513);
and U8121 (N_8121,N_7726,N_7844);
nor U8122 (N_8122,N_7771,N_7694);
nand U8123 (N_8123,N_7507,N_7798);
or U8124 (N_8124,N_7855,N_7943);
and U8125 (N_8125,N_7568,N_7979);
or U8126 (N_8126,N_7537,N_7736);
nand U8127 (N_8127,N_7690,N_7515);
or U8128 (N_8128,N_7959,N_7931);
or U8129 (N_8129,N_7647,N_7878);
nand U8130 (N_8130,N_7817,N_7595);
nand U8131 (N_8131,N_7848,N_7871);
nor U8132 (N_8132,N_7950,N_7593);
nand U8133 (N_8133,N_7717,N_7545);
nor U8134 (N_8134,N_7940,N_7981);
and U8135 (N_8135,N_7620,N_7555);
xnor U8136 (N_8136,N_7859,N_7704);
nand U8137 (N_8137,N_7701,N_7788);
and U8138 (N_8138,N_7582,N_7735);
xor U8139 (N_8139,N_7554,N_7820);
xnor U8140 (N_8140,N_7753,N_7556);
nor U8141 (N_8141,N_7972,N_7894);
and U8142 (N_8142,N_7836,N_7748);
and U8143 (N_8143,N_7790,N_7614);
xor U8144 (N_8144,N_7673,N_7631);
or U8145 (N_8145,N_7730,N_7893);
and U8146 (N_8146,N_7793,N_7964);
and U8147 (N_8147,N_7560,N_7920);
nor U8148 (N_8148,N_7765,N_7824);
and U8149 (N_8149,N_7789,N_7508);
nand U8150 (N_8150,N_7624,N_7772);
xor U8151 (N_8151,N_7742,N_7804);
xor U8152 (N_8152,N_7644,N_7722);
and U8153 (N_8153,N_7737,N_7810);
or U8154 (N_8154,N_7831,N_7621);
nor U8155 (N_8155,N_7843,N_7794);
xor U8156 (N_8156,N_7745,N_7777);
nand U8157 (N_8157,N_7639,N_7965);
nor U8158 (N_8158,N_7544,N_7578);
nand U8159 (N_8159,N_7926,N_7985);
nand U8160 (N_8160,N_7927,N_7574);
xor U8161 (N_8161,N_7827,N_7906);
nor U8162 (N_8162,N_7541,N_7571);
nor U8163 (N_8163,N_7785,N_7963);
nor U8164 (N_8164,N_7932,N_7881);
and U8165 (N_8165,N_7538,N_7749);
and U8166 (N_8166,N_7713,N_7823);
or U8167 (N_8167,N_7957,N_7873);
xor U8168 (N_8168,N_7896,N_7904);
nand U8169 (N_8169,N_7961,N_7930);
and U8170 (N_8170,N_7903,N_7629);
xor U8171 (N_8171,N_7850,N_7685);
or U8172 (N_8172,N_7529,N_7948);
and U8173 (N_8173,N_7633,N_7811);
nor U8174 (N_8174,N_7651,N_7996);
nand U8175 (N_8175,N_7700,N_7840);
nor U8176 (N_8176,N_7731,N_7976);
xor U8177 (N_8177,N_7547,N_7592);
or U8178 (N_8178,N_7526,N_7913);
xnor U8179 (N_8179,N_7990,N_7693);
xor U8180 (N_8180,N_7561,N_7596);
nand U8181 (N_8181,N_7882,N_7710);
and U8182 (N_8182,N_7778,N_7711);
and U8183 (N_8183,N_7936,N_7946);
and U8184 (N_8184,N_7680,N_7839);
nor U8185 (N_8185,N_7870,N_7888);
nor U8186 (N_8186,N_7934,N_7760);
nor U8187 (N_8187,N_7998,N_7914);
xnor U8188 (N_8188,N_7982,N_7818);
nand U8189 (N_8189,N_7536,N_7591);
nand U8190 (N_8190,N_7610,N_7857);
nand U8191 (N_8191,N_7806,N_7992);
nor U8192 (N_8192,N_7609,N_7611);
nor U8193 (N_8193,N_7608,N_7773);
nor U8194 (N_8194,N_7570,N_7670);
xor U8195 (N_8195,N_7709,N_7558);
xnor U8196 (N_8196,N_7712,N_7766);
and U8197 (N_8197,N_7552,N_7733);
or U8198 (N_8198,N_7705,N_7856);
or U8199 (N_8199,N_7895,N_7678);
nor U8200 (N_8200,N_7589,N_7911);
and U8201 (N_8201,N_7518,N_7833);
and U8202 (N_8202,N_7915,N_7533);
nor U8203 (N_8203,N_7706,N_7758);
and U8204 (N_8204,N_7980,N_7668);
xnor U8205 (N_8205,N_7594,N_7858);
nand U8206 (N_8206,N_7812,N_7767);
nand U8207 (N_8207,N_7885,N_7905);
and U8208 (N_8208,N_7945,N_7775);
xor U8209 (N_8209,N_7837,N_7822);
and U8210 (N_8210,N_7769,N_7692);
and U8211 (N_8211,N_7689,N_7887);
nor U8212 (N_8212,N_7987,N_7780);
and U8213 (N_8213,N_7923,N_7583);
nand U8214 (N_8214,N_7825,N_7565);
or U8215 (N_8215,N_7891,N_7791);
or U8216 (N_8216,N_7738,N_7868);
nand U8217 (N_8217,N_7732,N_7962);
or U8218 (N_8218,N_7504,N_7768);
and U8219 (N_8219,N_7866,N_7597);
nand U8220 (N_8220,N_7683,N_7522);
nor U8221 (N_8221,N_7686,N_7521);
xor U8222 (N_8222,N_7659,N_7728);
xnor U8223 (N_8223,N_7835,N_7665);
or U8224 (N_8224,N_7512,N_7601);
nand U8225 (N_8225,N_7675,N_7842);
nand U8226 (N_8226,N_7648,N_7684);
or U8227 (N_8227,N_7746,N_7543);
or U8228 (N_8228,N_7650,N_7783);
and U8229 (N_8229,N_7942,N_7899);
nor U8230 (N_8230,N_7511,N_7587);
nand U8231 (N_8231,N_7572,N_7636);
xnor U8232 (N_8232,N_7958,N_7664);
xor U8233 (N_8233,N_7761,N_7922);
and U8234 (N_8234,N_7688,N_7918);
or U8235 (N_8235,N_7853,N_7535);
nand U8236 (N_8236,N_7505,N_7886);
and U8237 (N_8237,N_7653,N_7925);
xor U8238 (N_8238,N_7553,N_7661);
nor U8239 (N_8239,N_7970,N_7534);
and U8240 (N_8240,N_7838,N_7784);
xnor U8241 (N_8241,N_7734,N_7687);
xnor U8242 (N_8242,N_7764,N_7921);
nor U8243 (N_8243,N_7944,N_7662);
and U8244 (N_8244,N_7719,N_7828);
nor U8245 (N_8245,N_7617,N_7723);
nor U8246 (N_8246,N_7974,N_7627);
nand U8247 (N_8247,N_7862,N_7612);
xnor U8248 (N_8248,N_7542,N_7519);
or U8249 (N_8249,N_7564,N_7501);
nor U8250 (N_8250,N_7852,N_7551);
and U8251 (N_8251,N_7625,N_7538);
nor U8252 (N_8252,N_7880,N_7892);
xor U8253 (N_8253,N_7707,N_7789);
and U8254 (N_8254,N_7901,N_7734);
and U8255 (N_8255,N_7597,N_7854);
or U8256 (N_8256,N_7572,N_7741);
xnor U8257 (N_8257,N_7563,N_7843);
nor U8258 (N_8258,N_7750,N_7734);
nor U8259 (N_8259,N_7665,N_7671);
nand U8260 (N_8260,N_7566,N_7757);
nor U8261 (N_8261,N_7676,N_7578);
and U8262 (N_8262,N_7552,N_7721);
or U8263 (N_8263,N_7734,N_7720);
nand U8264 (N_8264,N_7619,N_7789);
nand U8265 (N_8265,N_7687,N_7988);
or U8266 (N_8266,N_7504,N_7989);
or U8267 (N_8267,N_7642,N_7699);
nand U8268 (N_8268,N_7871,N_7606);
and U8269 (N_8269,N_7575,N_7893);
xor U8270 (N_8270,N_7587,N_7892);
nor U8271 (N_8271,N_7507,N_7629);
nor U8272 (N_8272,N_7963,N_7959);
and U8273 (N_8273,N_7936,N_7665);
xor U8274 (N_8274,N_7543,N_7727);
xnor U8275 (N_8275,N_7619,N_7854);
or U8276 (N_8276,N_7945,N_7604);
or U8277 (N_8277,N_7508,N_7606);
xor U8278 (N_8278,N_7933,N_7622);
or U8279 (N_8279,N_7762,N_7502);
nor U8280 (N_8280,N_7830,N_7964);
nor U8281 (N_8281,N_7726,N_7994);
nand U8282 (N_8282,N_7861,N_7930);
nor U8283 (N_8283,N_7946,N_7541);
nor U8284 (N_8284,N_7501,N_7975);
nand U8285 (N_8285,N_7633,N_7951);
xnor U8286 (N_8286,N_7809,N_7807);
nor U8287 (N_8287,N_7838,N_7668);
nor U8288 (N_8288,N_7699,N_7540);
nor U8289 (N_8289,N_7952,N_7577);
or U8290 (N_8290,N_7980,N_7903);
and U8291 (N_8291,N_7981,N_7985);
xor U8292 (N_8292,N_7992,N_7999);
and U8293 (N_8293,N_7813,N_7597);
and U8294 (N_8294,N_7872,N_7831);
nor U8295 (N_8295,N_7784,N_7909);
xnor U8296 (N_8296,N_7878,N_7651);
or U8297 (N_8297,N_7619,N_7640);
nand U8298 (N_8298,N_7675,N_7831);
nand U8299 (N_8299,N_7652,N_7535);
nor U8300 (N_8300,N_7666,N_7577);
nand U8301 (N_8301,N_7727,N_7834);
nor U8302 (N_8302,N_7929,N_7841);
nand U8303 (N_8303,N_7627,N_7528);
or U8304 (N_8304,N_7723,N_7647);
and U8305 (N_8305,N_7563,N_7878);
nand U8306 (N_8306,N_7912,N_7716);
nor U8307 (N_8307,N_7876,N_7623);
or U8308 (N_8308,N_7569,N_7525);
xnor U8309 (N_8309,N_7556,N_7781);
and U8310 (N_8310,N_7528,N_7929);
nand U8311 (N_8311,N_7541,N_7906);
or U8312 (N_8312,N_7831,N_7695);
and U8313 (N_8313,N_7992,N_7701);
and U8314 (N_8314,N_7642,N_7715);
nand U8315 (N_8315,N_7542,N_7689);
and U8316 (N_8316,N_7804,N_7712);
and U8317 (N_8317,N_7851,N_7709);
or U8318 (N_8318,N_7744,N_7589);
or U8319 (N_8319,N_7519,N_7685);
and U8320 (N_8320,N_7764,N_7600);
nand U8321 (N_8321,N_7596,N_7812);
xnor U8322 (N_8322,N_7925,N_7934);
nor U8323 (N_8323,N_7828,N_7679);
or U8324 (N_8324,N_7629,N_7664);
xor U8325 (N_8325,N_7538,N_7714);
nor U8326 (N_8326,N_7737,N_7595);
xnor U8327 (N_8327,N_7729,N_7914);
or U8328 (N_8328,N_7990,N_7547);
or U8329 (N_8329,N_7627,N_7939);
nor U8330 (N_8330,N_7796,N_7878);
and U8331 (N_8331,N_7751,N_7618);
nand U8332 (N_8332,N_7778,N_7771);
or U8333 (N_8333,N_7528,N_7717);
and U8334 (N_8334,N_7508,N_7528);
nand U8335 (N_8335,N_7663,N_7814);
xnor U8336 (N_8336,N_7882,N_7593);
or U8337 (N_8337,N_7666,N_7806);
or U8338 (N_8338,N_7781,N_7872);
xor U8339 (N_8339,N_7591,N_7801);
or U8340 (N_8340,N_7984,N_7685);
xor U8341 (N_8341,N_7645,N_7706);
and U8342 (N_8342,N_7716,N_7613);
or U8343 (N_8343,N_7698,N_7680);
nand U8344 (N_8344,N_7669,N_7929);
xor U8345 (N_8345,N_7626,N_7747);
xor U8346 (N_8346,N_7748,N_7971);
or U8347 (N_8347,N_7538,N_7629);
nor U8348 (N_8348,N_7522,N_7568);
nand U8349 (N_8349,N_7736,N_7574);
nor U8350 (N_8350,N_7933,N_7773);
and U8351 (N_8351,N_7921,N_7574);
nor U8352 (N_8352,N_7529,N_7577);
nor U8353 (N_8353,N_7838,N_7796);
and U8354 (N_8354,N_7741,N_7778);
xor U8355 (N_8355,N_7950,N_7687);
nand U8356 (N_8356,N_7806,N_7714);
xor U8357 (N_8357,N_7950,N_7518);
or U8358 (N_8358,N_7648,N_7655);
nand U8359 (N_8359,N_7721,N_7689);
and U8360 (N_8360,N_7973,N_7809);
nand U8361 (N_8361,N_7870,N_7855);
nor U8362 (N_8362,N_7834,N_7712);
xnor U8363 (N_8363,N_7821,N_7935);
and U8364 (N_8364,N_7599,N_7901);
or U8365 (N_8365,N_7810,N_7618);
nor U8366 (N_8366,N_7861,N_7710);
or U8367 (N_8367,N_7733,N_7625);
and U8368 (N_8368,N_7669,N_7928);
and U8369 (N_8369,N_7987,N_7722);
and U8370 (N_8370,N_7922,N_7646);
or U8371 (N_8371,N_7504,N_7929);
and U8372 (N_8372,N_7868,N_7869);
and U8373 (N_8373,N_7850,N_7623);
and U8374 (N_8374,N_7697,N_7841);
and U8375 (N_8375,N_7513,N_7913);
nor U8376 (N_8376,N_7699,N_7865);
nand U8377 (N_8377,N_7623,N_7815);
and U8378 (N_8378,N_7831,N_7802);
and U8379 (N_8379,N_7869,N_7739);
or U8380 (N_8380,N_7958,N_7605);
nand U8381 (N_8381,N_7641,N_7841);
nand U8382 (N_8382,N_7510,N_7974);
xnor U8383 (N_8383,N_7613,N_7869);
nand U8384 (N_8384,N_7649,N_7886);
nand U8385 (N_8385,N_7892,N_7723);
nand U8386 (N_8386,N_7891,N_7814);
and U8387 (N_8387,N_7708,N_7960);
nor U8388 (N_8388,N_7761,N_7641);
nand U8389 (N_8389,N_7538,N_7738);
xor U8390 (N_8390,N_7823,N_7981);
nor U8391 (N_8391,N_7946,N_7673);
or U8392 (N_8392,N_7995,N_7790);
nor U8393 (N_8393,N_7679,N_7835);
xor U8394 (N_8394,N_7581,N_7565);
and U8395 (N_8395,N_7585,N_7937);
or U8396 (N_8396,N_7809,N_7872);
nand U8397 (N_8397,N_7666,N_7633);
and U8398 (N_8398,N_7646,N_7558);
xnor U8399 (N_8399,N_7561,N_7533);
nand U8400 (N_8400,N_7905,N_7623);
nand U8401 (N_8401,N_7766,N_7989);
nor U8402 (N_8402,N_7545,N_7548);
nor U8403 (N_8403,N_7981,N_7626);
nor U8404 (N_8404,N_7578,N_7921);
and U8405 (N_8405,N_7523,N_7845);
xnor U8406 (N_8406,N_7743,N_7869);
nand U8407 (N_8407,N_7652,N_7809);
or U8408 (N_8408,N_7831,N_7506);
xor U8409 (N_8409,N_7568,N_7939);
xor U8410 (N_8410,N_7893,N_7642);
nand U8411 (N_8411,N_7518,N_7882);
nor U8412 (N_8412,N_7624,N_7922);
or U8413 (N_8413,N_7587,N_7598);
nor U8414 (N_8414,N_7564,N_7647);
and U8415 (N_8415,N_7856,N_7783);
xor U8416 (N_8416,N_7909,N_7931);
nand U8417 (N_8417,N_7622,N_7869);
and U8418 (N_8418,N_7695,N_7782);
nor U8419 (N_8419,N_7797,N_7650);
nor U8420 (N_8420,N_7890,N_7771);
or U8421 (N_8421,N_7773,N_7786);
or U8422 (N_8422,N_7511,N_7730);
and U8423 (N_8423,N_7559,N_7527);
and U8424 (N_8424,N_7892,N_7574);
xor U8425 (N_8425,N_7603,N_7511);
nand U8426 (N_8426,N_7825,N_7686);
xor U8427 (N_8427,N_7725,N_7743);
xor U8428 (N_8428,N_7997,N_7504);
xnor U8429 (N_8429,N_7964,N_7767);
or U8430 (N_8430,N_7544,N_7700);
nor U8431 (N_8431,N_7977,N_7740);
or U8432 (N_8432,N_7988,N_7565);
or U8433 (N_8433,N_7503,N_7784);
nand U8434 (N_8434,N_7814,N_7678);
nand U8435 (N_8435,N_7764,N_7991);
nor U8436 (N_8436,N_7910,N_7898);
xor U8437 (N_8437,N_7863,N_7640);
and U8438 (N_8438,N_7660,N_7530);
nand U8439 (N_8439,N_7569,N_7552);
and U8440 (N_8440,N_7854,N_7822);
and U8441 (N_8441,N_7682,N_7992);
xnor U8442 (N_8442,N_7887,N_7560);
or U8443 (N_8443,N_7628,N_7675);
nand U8444 (N_8444,N_7734,N_7560);
and U8445 (N_8445,N_7660,N_7797);
or U8446 (N_8446,N_7703,N_7602);
xor U8447 (N_8447,N_7536,N_7539);
xor U8448 (N_8448,N_7811,N_7878);
xor U8449 (N_8449,N_7700,N_7560);
or U8450 (N_8450,N_7882,N_7800);
xor U8451 (N_8451,N_7840,N_7811);
and U8452 (N_8452,N_7920,N_7925);
xnor U8453 (N_8453,N_7650,N_7890);
nor U8454 (N_8454,N_7761,N_7797);
or U8455 (N_8455,N_7811,N_7648);
or U8456 (N_8456,N_7887,N_7555);
nand U8457 (N_8457,N_7923,N_7924);
nand U8458 (N_8458,N_7832,N_7516);
and U8459 (N_8459,N_7809,N_7734);
xor U8460 (N_8460,N_7572,N_7859);
and U8461 (N_8461,N_7657,N_7711);
nor U8462 (N_8462,N_7567,N_7984);
nor U8463 (N_8463,N_7591,N_7876);
nor U8464 (N_8464,N_7663,N_7712);
or U8465 (N_8465,N_7988,N_7561);
nor U8466 (N_8466,N_7722,N_7865);
nand U8467 (N_8467,N_7571,N_7531);
and U8468 (N_8468,N_7935,N_7573);
xnor U8469 (N_8469,N_7872,N_7979);
nor U8470 (N_8470,N_7902,N_7877);
nand U8471 (N_8471,N_7822,N_7951);
nor U8472 (N_8472,N_7736,N_7621);
nor U8473 (N_8473,N_7782,N_7824);
nor U8474 (N_8474,N_7699,N_7515);
nor U8475 (N_8475,N_7620,N_7835);
nand U8476 (N_8476,N_7686,N_7861);
and U8477 (N_8477,N_7934,N_7928);
nand U8478 (N_8478,N_7626,N_7720);
xnor U8479 (N_8479,N_7639,N_7911);
xor U8480 (N_8480,N_7695,N_7937);
nand U8481 (N_8481,N_7530,N_7719);
and U8482 (N_8482,N_7719,N_7604);
xor U8483 (N_8483,N_7846,N_7763);
xor U8484 (N_8484,N_7649,N_7592);
nor U8485 (N_8485,N_7660,N_7970);
nand U8486 (N_8486,N_7888,N_7930);
or U8487 (N_8487,N_7775,N_7550);
and U8488 (N_8488,N_7669,N_7729);
and U8489 (N_8489,N_7764,N_7679);
xor U8490 (N_8490,N_7829,N_7791);
and U8491 (N_8491,N_7985,N_7545);
or U8492 (N_8492,N_7832,N_7694);
nor U8493 (N_8493,N_7915,N_7990);
xnor U8494 (N_8494,N_7889,N_7743);
xnor U8495 (N_8495,N_7920,N_7701);
and U8496 (N_8496,N_7881,N_7622);
or U8497 (N_8497,N_7999,N_7722);
and U8498 (N_8498,N_7657,N_7697);
xor U8499 (N_8499,N_7553,N_7574);
xnor U8500 (N_8500,N_8375,N_8008);
and U8501 (N_8501,N_8183,N_8386);
nand U8502 (N_8502,N_8294,N_8059);
nor U8503 (N_8503,N_8397,N_8248);
or U8504 (N_8504,N_8128,N_8408);
xor U8505 (N_8505,N_8004,N_8211);
and U8506 (N_8506,N_8096,N_8090);
nor U8507 (N_8507,N_8335,N_8066);
or U8508 (N_8508,N_8041,N_8224);
xnor U8509 (N_8509,N_8115,N_8092);
and U8510 (N_8510,N_8409,N_8237);
nand U8511 (N_8511,N_8190,N_8209);
or U8512 (N_8512,N_8444,N_8165);
xor U8513 (N_8513,N_8022,N_8232);
nor U8514 (N_8514,N_8295,N_8137);
nor U8515 (N_8515,N_8253,N_8461);
nand U8516 (N_8516,N_8406,N_8478);
xor U8517 (N_8517,N_8474,N_8158);
xor U8518 (N_8518,N_8496,N_8378);
and U8519 (N_8519,N_8391,N_8364);
nand U8520 (N_8520,N_8304,N_8073);
xnor U8521 (N_8521,N_8194,N_8230);
or U8522 (N_8522,N_8407,N_8291);
or U8523 (N_8523,N_8275,N_8055);
nor U8524 (N_8524,N_8207,N_8220);
or U8525 (N_8525,N_8459,N_8396);
nor U8526 (N_8526,N_8213,N_8104);
or U8527 (N_8527,N_8118,N_8473);
nand U8528 (N_8528,N_8347,N_8219);
or U8529 (N_8529,N_8423,N_8228);
nand U8530 (N_8530,N_8105,N_8257);
nor U8531 (N_8531,N_8164,N_8348);
xor U8532 (N_8532,N_8280,N_8184);
nor U8533 (N_8533,N_8203,N_8465);
or U8534 (N_8534,N_8132,N_8350);
xnor U8535 (N_8535,N_8082,N_8249);
xnor U8536 (N_8536,N_8395,N_8149);
or U8537 (N_8537,N_8269,N_8188);
nand U8538 (N_8538,N_8387,N_8094);
or U8539 (N_8539,N_8307,N_8223);
or U8540 (N_8540,N_8439,N_8365);
or U8541 (N_8541,N_8141,N_8413);
nor U8542 (N_8542,N_8086,N_8298);
and U8543 (N_8543,N_8246,N_8495);
nand U8544 (N_8544,N_8472,N_8101);
xnor U8545 (N_8545,N_8072,N_8468);
nand U8546 (N_8546,N_8368,N_8171);
and U8547 (N_8547,N_8242,N_8259);
and U8548 (N_8548,N_8075,N_8212);
or U8549 (N_8549,N_8060,N_8255);
xor U8550 (N_8550,N_8139,N_8160);
nor U8551 (N_8551,N_8482,N_8310);
nand U8552 (N_8552,N_8093,N_8388);
nand U8553 (N_8553,N_8315,N_8309);
xor U8554 (N_8554,N_8229,N_8360);
or U8555 (N_8555,N_8089,N_8150);
nor U8556 (N_8556,N_8023,N_8447);
xor U8557 (N_8557,N_8061,N_8169);
nand U8558 (N_8558,N_8467,N_8427);
nor U8559 (N_8559,N_8038,N_8369);
nor U8560 (N_8560,N_8216,N_8167);
and U8561 (N_8561,N_8372,N_8177);
xor U8562 (N_8562,N_8120,N_8497);
xor U8563 (N_8563,N_8479,N_8117);
nand U8564 (N_8564,N_8020,N_8130);
or U8565 (N_8565,N_8109,N_8252);
nand U8566 (N_8566,N_8018,N_8341);
xor U8567 (N_8567,N_8499,N_8153);
xnor U8568 (N_8568,N_8371,N_8050);
xor U8569 (N_8569,N_8488,N_8078);
nand U8570 (N_8570,N_8250,N_8454);
nor U8571 (N_8571,N_8178,N_8264);
and U8572 (N_8572,N_8062,N_8057);
nand U8573 (N_8573,N_8483,N_8100);
and U8574 (N_8574,N_8359,N_8056);
or U8575 (N_8575,N_8470,N_8279);
nor U8576 (N_8576,N_8311,N_8452);
xor U8577 (N_8577,N_8205,N_8431);
nor U8578 (N_8578,N_8134,N_8144);
or U8579 (N_8579,N_8035,N_8155);
nand U8580 (N_8580,N_8377,N_8106);
xnor U8581 (N_8581,N_8464,N_8014);
and U8582 (N_8582,N_8374,N_8006);
xnor U8583 (N_8583,N_8111,N_8485);
nor U8584 (N_8584,N_8481,N_8285);
nor U8585 (N_8585,N_8426,N_8446);
xnor U8586 (N_8586,N_8182,N_8438);
nand U8587 (N_8587,N_8079,N_8463);
nand U8588 (N_8588,N_8352,N_8049);
nor U8589 (N_8589,N_8323,N_8052);
nor U8590 (N_8590,N_8270,N_8290);
nand U8591 (N_8591,N_8174,N_8490);
nor U8592 (N_8592,N_8484,N_8027);
xnor U8593 (N_8593,N_8462,N_8168);
xor U8594 (N_8594,N_8487,N_8084);
nand U8595 (N_8595,N_8354,N_8381);
and U8596 (N_8596,N_8260,N_8019);
xor U8597 (N_8597,N_8399,N_8428);
nand U8598 (N_8598,N_8114,N_8091);
xor U8599 (N_8599,N_8015,N_8097);
nand U8600 (N_8600,N_8394,N_8455);
nor U8601 (N_8601,N_8419,N_8453);
nor U8602 (N_8602,N_8021,N_8405);
nand U8603 (N_8603,N_8429,N_8210);
or U8604 (N_8604,N_8276,N_8321);
xnor U8605 (N_8605,N_8493,N_8486);
nor U8606 (N_8606,N_8332,N_8256);
nand U8607 (N_8607,N_8414,N_8028);
xor U8608 (N_8608,N_8379,N_8099);
xor U8609 (N_8609,N_8047,N_8334);
and U8610 (N_8610,N_8245,N_8340);
or U8611 (N_8611,N_8051,N_8425);
and U8612 (N_8612,N_8226,N_8494);
xor U8613 (N_8613,N_8119,N_8272);
nor U8614 (N_8614,N_8342,N_8392);
and U8615 (N_8615,N_8126,N_8054);
and U8616 (N_8616,N_8234,N_8244);
or U8617 (N_8617,N_8030,N_8036);
nor U8618 (N_8618,N_8314,N_8147);
nor U8619 (N_8619,N_8225,N_8287);
nand U8620 (N_8620,N_8327,N_8007);
xnor U8621 (N_8621,N_8476,N_8068);
nor U8622 (N_8622,N_8001,N_8010);
nand U8623 (N_8623,N_8361,N_8357);
nand U8624 (N_8624,N_8284,N_8411);
or U8625 (N_8625,N_8031,N_8238);
and U8626 (N_8626,N_8353,N_8112);
xor U8627 (N_8627,N_8331,N_8319);
nand U8628 (N_8628,N_8159,N_8355);
nor U8629 (N_8629,N_8186,N_8157);
and U8630 (N_8630,N_8013,N_8005);
nor U8631 (N_8631,N_8326,N_8033);
and U8632 (N_8632,N_8161,N_8265);
nand U8633 (N_8633,N_8063,N_8330);
xor U8634 (N_8634,N_8192,N_8067);
and U8635 (N_8635,N_8129,N_8181);
and U8636 (N_8636,N_8324,N_8131);
or U8637 (N_8637,N_8286,N_8201);
and U8638 (N_8638,N_8198,N_8227);
or U8639 (N_8639,N_8443,N_8222);
and U8640 (N_8640,N_8301,N_8363);
or U8641 (N_8641,N_8195,N_8029);
or U8642 (N_8642,N_8123,N_8489);
xor U8643 (N_8643,N_8121,N_8113);
or U8644 (N_8644,N_8384,N_8432);
nand U8645 (N_8645,N_8085,N_8338);
and U8646 (N_8646,N_8045,N_8302);
nor U8647 (N_8647,N_8231,N_8012);
nor U8648 (N_8648,N_8337,N_8058);
xnor U8649 (N_8649,N_8011,N_8032);
nand U8650 (N_8650,N_8122,N_8283);
nor U8651 (N_8651,N_8403,N_8017);
or U8652 (N_8652,N_8125,N_8176);
nor U8653 (N_8653,N_8383,N_8039);
and U8654 (N_8654,N_8268,N_8390);
and U8655 (N_8655,N_8278,N_8448);
xnor U8656 (N_8656,N_8095,N_8366);
and U8657 (N_8657,N_8044,N_8344);
xor U8658 (N_8658,N_8373,N_8345);
nor U8659 (N_8659,N_8197,N_8308);
or U8660 (N_8660,N_8170,N_8136);
xor U8661 (N_8661,N_8305,N_8346);
xor U8662 (N_8662,N_8376,N_8401);
or U8663 (N_8663,N_8235,N_8456);
and U8664 (N_8664,N_8152,N_8313);
or U8665 (N_8665,N_8258,N_8402);
or U8666 (N_8666,N_8214,N_8179);
and U8667 (N_8667,N_8262,N_8065);
xnor U8668 (N_8668,N_8422,N_8303);
nor U8669 (N_8669,N_8243,N_8200);
and U8670 (N_8670,N_8202,N_8292);
or U8671 (N_8671,N_8325,N_8204);
nand U8672 (N_8672,N_8163,N_8440);
nand U8673 (N_8673,N_8077,N_8025);
nand U8674 (N_8674,N_8333,N_8247);
nand U8675 (N_8675,N_8329,N_8288);
nor U8676 (N_8676,N_8215,N_8273);
xnor U8677 (N_8677,N_8380,N_8145);
nor U8678 (N_8678,N_8351,N_8471);
xnor U8679 (N_8679,N_8180,N_8233);
xor U8680 (N_8680,N_8140,N_8138);
and U8681 (N_8681,N_8221,N_8433);
xor U8682 (N_8682,N_8362,N_8103);
or U8683 (N_8683,N_8316,N_8069);
xor U8684 (N_8684,N_8102,N_8124);
and U8685 (N_8685,N_8281,N_8107);
and U8686 (N_8686,N_8175,N_8196);
and U8687 (N_8687,N_8458,N_8274);
and U8688 (N_8688,N_8080,N_8110);
xnor U8689 (N_8689,N_8437,N_8236);
or U8690 (N_8690,N_8451,N_8434);
xor U8691 (N_8691,N_8420,N_8261);
nor U8692 (N_8692,N_8475,N_8173);
or U8693 (N_8693,N_8026,N_8267);
and U8694 (N_8694,N_8339,N_8208);
xor U8695 (N_8695,N_8460,N_8336);
and U8696 (N_8696,N_8081,N_8430);
nor U8697 (N_8697,N_8450,N_8166);
nor U8698 (N_8698,N_8469,N_8436);
nor U8699 (N_8699,N_8083,N_8398);
or U8700 (N_8700,N_8477,N_8410);
xnor U8701 (N_8701,N_8009,N_8116);
nor U8702 (N_8702,N_8343,N_8034);
or U8703 (N_8703,N_8435,N_8441);
or U8704 (N_8704,N_8162,N_8156);
or U8705 (N_8705,N_8254,N_8187);
nor U8706 (N_8706,N_8498,N_8356);
nand U8707 (N_8707,N_8385,N_8206);
or U8708 (N_8708,N_8071,N_8322);
nor U8709 (N_8709,N_8133,N_8393);
nand U8710 (N_8710,N_8306,N_8108);
xnor U8711 (N_8711,N_8400,N_8241);
or U8712 (N_8712,N_8480,N_8142);
or U8713 (N_8713,N_8098,N_8271);
and U8714 (N_8714,N_8240,N_8191);
and U8715 (N_8715,N_8416,N_8076);
or U8716 (N_8716,N_8043,N_8421);
or U8717 (N_8717,N_8299,N_8266);
xnor U8718 (N_8718,N_8296,N_8003);
xnor U8719 (N_8719,N_8087,N_8127);
or U8720 (N_8720,N_8418,N_8037);
or U8721 (N_8721,N_8143,N_8449);
or U8722 (N_8722,N_8088,N_8415);
or U8723 (N_8723,N_8239,N_8492);
nor U8724 (N_8724,N_8466,N_8024);
nor U8725 (N_8725,N_8070,N_8297);
nand U8726 (N_8726,N_8282,N_8000);
and U8727 (N_8727,N_8074,N_8277);
nor U8728 (N_8728,N_8367,N_8317);
and U8729 (N_8729,N_8442,N_8064);
xor U8730 (N_8730,N_8293,N_8358);
or U8731 (N_8731,N_8189,N_8320);
xor U8732 (N_8732,N_8148,N_8193);
or U8733 (N_8733,N_8154,N_8046);
xnor U8734 (N_8734,N_8135,N_8417);
and U8735 (N_8735,N_8042,N_8185);
or U8736 (N_8736,N_8199,N_8445);
or U8737 (N_8737,N_8424,N_8318);
nor U8738 (N_8738,N_8146,N_8016);
or U8739 (N_8739,N_8349,N_8002);
nor U8740 (N_8740,N_8491,N_8412);
xor U8741 (N_8741,N_8382,N_8328);
and U8742 (N_8742,N_8300,N_8053);
and U8743 (N_8743,N_8370,N_8040);
and U8744 (N_8744,N_8389,N_8172);
nor U8745 (N_8745,N_8263,N_8289);
nor U8746 (N_8746,N_8048,N_8151);
xnor U8747 (N_8747,N_8457,N_8312);
and U8748 (N_8748,N_8217,N_8251);
nor U8749 (N_8749,N_8218,N_8404);
nor U8750 (N_8750,N_8341,N_8430);
nand U8751 (N_8751,N_8298,N_8146);
nor U8752 (N_8752,N_8096,N_8225);
nand U8753 (N_8753,N_8405,N_8164);
xnor U8754 (N_8754,N_8261,N_8002);
or U8755 (N_8755,N_8193,N_8171);
and U8756 (N_8756,N_8051,N_8356);
or U8757 (N_8757,N_8445,N_8271);
or U8758 (N_8758,N_8499,N_8381);
nand U8759 (N_8759,N_8266,N_8356);
xnor U8760 (N_8760,N_8449,N_8282);
nor U8761 (N_8761,N_8393,N_8091);
or U8762 (N_8762,N_8320,N_8391);
or U8763 (N_8763,N_8294,N_8296);
nand U8764 (N_8764,N_8051,N_8017);
nand U8765 (N_8765,N_8270,N_8381);
or U8766 (N_8766,N_8185,N_8147);
nand U8767 (N_8767,N_8412,N_8426);
nand U8768 (N_8768,N_8478,N_8111);
nand U8769 (N_8769,N_8096,N_8056);
or U8770 (N_8770,N_8271,N_8494);
and U8771 (N_8771,N_8085,N_8046);
nand U8772 (N_8772,N_8202,N_8472);
xor U8773 (N_8773,N_8310,N_8489);
nand U8774 (N_8774,N_8086,N_8047);
xnor U8775 (N_8775,N_8154,N_8403);
or U8776 (N_8776,N_8305,N_8484);
and U8777 (N_8777,N_8246,N_8296);
or U8778 (N_8778,N_8430,N_8027);
nand U8779 (N_8779,N_8032,N_8368);
xnor U8780 (N_8780,N_8415,N_8336);
nand U8781 (N_8781,N_8371,N_8013);
nor U8782 (N_8782,N_8137,N_8314);
xor U8783 (N_8783,N_8448,N_8330);
xor U8784 (N_8784,N_8224,N_8324);
xnor U8785 (N_8785,N_8037,N_8216);
or U8786 (N_8786,N_8276,N_8443);
and U8787 (N_8787,N_8172,N_8220);
or U8788 (N_8788,N_8460,N_8441);
nand U8789 (N_8789,N_8073,N_8109);
or U8790 (N_8790,N_8005,N_8485);
nor U8791 (N_8791,N_8214,N_8127);
xnor U8792 (N_8792,N_8020,N_8162);
nand U8793 (N_8793,N_8217,N_8270);
nor U8794 (N_8794,N_8431,N_8397);
xnor U8795 (N_8795,N_8490,N_8112);
and U8796 (N_8796,N_8150,N_8404);
nand U8797 (N_8797,N_8473,N_8050);
xnor U8798 (N_8798,N_8438,N_8362);
nand U8799 (N_8799,N_8460,N_8451);
nor U8800 (N_8800,N_8225,N_8312);
nand U8801 (N_8801,N_8281,N_8137);
xor U8802 (N_8802,N_8142,N_8055);
nor U8803 (N_8803,N_8213,N_8146);
nand U8804 (N_8804,N_8005,N_8417);
nand U8805 (N_8805,N_8472,N_8358);
nor U8806 (N_8806,N_8033,N_8259);
and U8807 (N_8807,N_8460,N_8243);
nor U8808 (N_8808,N_8485,N_8253);
and U8809 (N_8809,N_8140,N_8201);
nand U8810 (N_8810,N_8356,N_8399);
and U8811 (N_8811,N_8469,N_8008);
and U8812 (N_8812,N_8034,N_8190);
nand U8813 (N_8813,N_8349,N_8379);
nor U8814 (N_8814,N_8064,N_8278);
xor U8815 (N_8815,N_8245,N_8320);
nor U8816 (N_8816,N_8246,N_8453);
nand U8817 (N_8817,N_8276,N_8195);
and U8818 (N_8818,N_8099,N_8345);
and U8819 (N_8819,N_8341,N_8267);
nand U8820 (N_8820,N_8288,N_8455);
nor U8821 (N_8821,N_8467,N_8370);
nor U8822 (N_8822,N_8452,N_8301);
and U8823 (N_8823,N_8356,N_8014);
xor U8824 (N_8824,N_8317,N_8016);
and U8825 (N_8825,N_8283,N_8130);
and U8826 (N_8826,N_8360,N_8218);
or U8827 (N_8827,N_8147,N_8409);
or U8828 (N_8828,N_8108,N_8488);
xor U8829 (N_8829,N_8101,N_8316);
or U8830 (N_8830,N_8297,N_8159);
xor U8831 (N_8831,N_8311,N_8030);
nor U8832 (N_8832,N_8476,N_8499);
and U8833 (N_8833,N_8068,N_8074);
or U8834 (N_8834,N_8145,N_8118);
or U8835 (N_8835,N_8337,N_8088);
xnor U8836 (N_8836,N_8256,N_8366);
nor U8837 (N_8837,N_8326,N_8488);
xnor U8838 (N_8838,N_8472,N_8249);
nand U8839 (N_8839,N_8449,N_8064);
or U8840 (N_8840,N_8174,N_8227);
and U8841 (N_8841,N_8059,N_8475);
and U8842 (N_8842,N_8044,N_8465);
nor U8843 (N_8843,N_8319,N_8257);
or U8844 (N_8844,N_8345,N_8034);
xor U8845 (N_8845,N_8279,N_8348);
or U8846 (N_8846,N_8016,N_8409);
nand U8847 (N_8847,N_8248,N_8273);
or U8848 (N_8848,N_8251,N_8128);
and U8849 (N_8849,N_8087,N_8149);
and U8850 (N_8850,N_8071,N_8450);
or U8851 (N_8851,N_8184,N_8163);
or U8852 (N_8852,N_8358,N_8160);
and U8853 (N_8853,N_8143,N_8411);
nor U8854 (N_8854,N_8428,N_8161);
nor U8855 (N_8855,N_8412,N_8314);
xnor U8856 (N_8856,N_8276,N_8355);
nor U8857 (N_8857,N_8227,N_8319);
nor U8858 (N_8858,N_8334,N_8245);
and U8859 (N_8859,N_8140,N_8044);
nor U8860 (N_8860,N_8341,N_8182);
nor U8861 (N_8861,N_8246,N_8333);
and U8862 (N_8862,N_8180,N_8131);
nand U8863 (N_8863,N_8185,N_8461);
xor U8864 (N_8864,N_8364,N_8324);
nand U8865 (N_8865,N_8352,N_8253);
xor U8866 (N_8866,N_8429,N_8473);
nand U8867 (N_8867,N_8444,N_8042);
xor U8868 (N_8868,N_8470,N_8012);
and U8869 (N_8869,N_8194,N_8025);
xnor U8870 (N_8870,N_8188,N_8487);
and U8871 (N_8871,N_8138,N_8047);
nand U8872 (N_8872,N_8409,N_8492);
nor U8873 (N_8873,N_8156,N_8010);
and U8874 (N_8874,N_8325,N_8442);
nor U8875 (N_8875,N_8001,N_8330);
and U8876 (N_8876,N_8423,N_8172);
and U8877 (N_8877,N_8141,N_8435);
or U8878 (N_8878,N_8029,N_8154);
nor U8879 (N_8879,N_8221,N_8013);
nor U8880 (N_8880,N_8046,N_8037);
nor U8881 (N_8881,N_8238,N_8456);
or U8882 (N_8882,N_8176,N_8392);
nand U8883 (N_8883,N_8001,N_8309);
nand U8884 (N_8884,N_8451,N_8417);
nand U8885 (N_8885,N_8007,N_8397);
nand U8886 (N_8886,N_8396,N_8208);
or U8887 (N_8887,N_8265,N_8181);
nand U8888 (N_8888,N_8455,N_8184);
or U8889 (N_8889,N_8066,N_8315);
xnor U8890 (N_8890,N_8037,N_8131);
and U8891 (N_8891,N_8152,N_8410);
nand U8892 (N_8892,N_8122,N_8169);
and U8893 (N_8893,N_8489,N_8271);
xnor U8894 (N_8894,N_8007,N_8271);
nor U8895 (N_8895,N_8460,N_8059);
nor U8896 (N_8896,N_8288,N_8204);
or U8897 (N_8897,N_8459,N_8168);
nor U8898 (N_8898,N_8482,N_8152);
or U8899 (N_8899,N_8489,N_8115);
xnor U8900 (N_8900,N_8397,N_8026);
and U8901 (N_8901,N_8176,N_8483);
nor U8902 (N_8902,N_8444,N_8062);
and U8903 (N_8903,N_8010,N_8133);
and U8904 (N_8904,N_8069,N_8323);
nor U8905 (N_8905,N_8447,N_8303);
nor U8906 (N_8906,N_8060,N_8265);
xor U8907 (N_8907,N_8399,N_8121);
and U8908 (N_8908,N_8008,N_8420);
and U8909 (N_8909,N_8208,N_8334);
xnor U8910 (N_8910,N_8160,N_8243);
nand U8911 (N_8911,N_8157,N_8280);
and U8912 (N_8912,N_8471,N_8440);
xnor U8913 (N_8913,N_8464,N_8039);
and U8914 (N_8914,N_8484,N_8105);
nor U8915 (N_8915,N_8441,N_8084);
and U8916 (N_8916,N_8012,N_8097);
nor U8917 (N_8917,N_8051,N_8100);
nand U8918 (N_8918,N_8131,N_8191);
and U8919 (N_8919,N_8238,N_8177);
nand U8920 (N_8920,N_8191,N_8239);
nor U8921 (N_8921,N_8288,N_8008);
nand U8922 (N_8922,N_8207,N_8359);
and U8923 (N_8923,N_8262,N_8105);
nor U8924 (N_8924,N_8449,N_8204);
nand U8925 (N_8925,N_8003,N_8197);
or U8926 (N_8926,N_8050,N_8315);
and U8927 (N_8927,N_8125,N_8002);
nand U8928 (N_8928,N_8186,N_8399);
and U8929 (N_8929,N_8178,N_8009);
xnor U8930 (N_8930,N_8220,N_8043);
nand U8931 (N_8931,N_8071,N_8244);
nand U8932 (N_8932,N_8044,N_8451);
nand U8933 (N_8933,N_8353,N_8179);
nand U8934 (N_8934,N_8390,N_8213);
or U8935 (N_8935,N_8134,N_8397);
xor U8936 (N_8936,N_8167,N_8123);
xnor U8937 (N_8937,N_8069,N_8358);
and U8938 (N_8938,N_8132,N_8044);
or U8939 (N_8939,N_8481,N_8207);
or U8940 (N_8940,N_8488,N_8114);
nor U8941 (N_8941,N_8404,N_8121);
or U8942 (N_8942,N_8025,N_8263);
and U8943 (N_8943,N_8061,N_8074);
nor U8944 (N_8944,N_8342,N_8337);
and U8945 (N_8945,N_8163,N_8106);
or U8946 (N_8946,N_8291,N_8053);
nor U8947 (N_8947,N_8169,N_8456);
or U8948 (N_8948,N_8456,N_8039);
and U8949 (N_8949,N_8133,N_8124);
or U8950 (N_8950,N_8252,N_8279);
and U8951 (N_8951,N_8048,N_8223);
xnor U8952 (N_8952,N_8132,N_8403);
nand U8953 (N_8953,N_8232,N_8471);
and U8954 (N_8954,N_8023,N_8472);
nand U8955 (N_8955,N_8087,N_8383);
nor U8956 (N_8956,N_8015,N_8480);
nor U8957 (N_8957,N_8351,N_8205);
nor U8958 (N_8958,N_8486,N_8380);
or U8959 (N_8959,N_8004,N_8298);
nor U8960 (N_8960,N_8327,N_8063);
nor U8961 (N_8961,N_8183,N_8121);
and U8962 (N_8962,N_8097,N_8474);
nor U8963 (N_8963,N_8053,N_8478);
and U8964 (N_8964,N_8274,N_8281);
or U8965 (N_8965,N_8194,N_8296);
nor U8966 (N_8966,N_8095,N_8425);
nand U8967 (N_8967,N_8076,N_8337);
nor U8968 (N_8968,N_8151,N_8077);
nor U8969 (N_8969,N_8227,N_8256);
nor U8970 (N_8970,N_8434,N_8378);
nor U8971 (N_8971,N_8310,N_8312);
or U8972 (N_8972,N_8034,N_8324);
and U8973 (N_8973,N_8380,N_8088);
nor U8974 (N_8974,N_8061,N_8272);
nand U8975 (N_8975,N_8152,N_8030);
nor U8976 (N_8976,N_8346,N_8421);
nor U8977 (N_8977,N_8493,N_8258);
nor U8978 (N_8978,N_8434,N_8201);
xnor U8979 (N_8979,N_8491,N_8436);
nor U8980 (N_8980,N_8014,N_8313);
nand U8981 (N_8981,N_8085,N_8488);
or U8982 (N_8982,N_8387,N_8323);
xnor U8983 (N_8983,N_8205,N_8433);
nor U8984 (N_8984,N_8341,N_8133);
and U8985 (N_8985,N_8274,N_8295);
and U8986 (N_8986,N_8068,N_8330);
xor U8987 (N_8987,N_8253,N_8136);
nor U8988 (N_8988,N_8295,N_8093);
and U8989 (N_8989,N_8099,N_8341);
nand U8990 (N_8990,N_8330,N_8058);
nor U8991 (N_8991,N_8044,N_8063);
and U8992 (N_8992,N_8302,N_8440);
nor U8993 (N_8993,N_8139,N_8164);
xor U8994 (N_8994,N_8282,N_8065);
or U8995 (N_8995,N_8144,N_8369);
nor U8996 (N_8996,N_8456,N_8150);
nand U8997 (N_8997,N_8169,N_8486);
nand U8998 (N_8998,N_8288,N_8158);
or U8999 (N_8999,N_8081,N_8184);
or U9000 (N_9000,N_8998,N_8829);
xor U9001 (N_9001,N_8686,N_8824);
xnor U9002 (N_9002,N_8999,N_8876);
nor U9003 (N_9003,N_8843,N_8744);
nor U9004 (N_9004,N_8968,N_8530);
nand U9005 (N_9005,N_8882,N_8958);
xor U9006 (N_9006,N_8611,N_8581);
or U9007 (N_9007,N_8650,N_8616);
nand U9008 (N_9008,N_8584,N_8503);
or U9009 (N_9009,N_8796,N_8513);
xnor U9010 (N_9010,N_8870,N_8685);
nand U9011 (N_9011,N_8659,N_8875);
nor U9012 (N_9012,N_8730,N_8733);
xnor U9013 (N_9013,N_8805,N_8562);
and U9014 (N_9014,N_8606,N_8754);
or U9015 (N_9015,N_8945,N_8900);
and U9016 (N_9016,N_8936,N_8745);
nor U9017 (N_9017,N_8831,N_8612);
and U9018 (N_9018,N_8782,N_8897);
or U9019 (N_9019,N_8708,N_8701);
nand U9020 (N_9020,N_8880,N_8813);
nor U9021 (N_9021,N_8605,N_8825);
nand U9022 (N_9022,N_8556,N_8854);
and U9023 (N_9023,N_8535,N_8987);
or U9024 (N_9024,N_8697,N_8981);
or U9025 (N_9025,N_8704,N_8515);
xnor U9026 (N_9026,N_8959,N_8617);
xnor U9027 (N_9027,N_8627,N_8988);
or U9028 (N_9028,N_8523,N_8941);
nor U9029 (N_9029,N_8806,N_8895);
nor U9030 (N_9030,N_8516,N_8888);
nand U9031 (N_9031,N_8613,N_8770);
nand U9032 (N_9032,N_8669,N_8868);
or U9033 (N_9033,N_8544,N_8529);
and U9034 (N_9034,N_8896,N_8756);
nor U9035 (N_9035,N_8543,N_8582);
nand U9036 (N_9036,N_8536,N_8654);
and U9037 (N_9037,N_8852,N_8815);
and U9038 (N_9038,N_8681,N_8711);
or U9039 (N_9039,N_8661,N_8737);
and U9040 (N_9040,N_8548,N_8618);
nor U9041 (N_9041,N_8920,N_8647);
nor U9042 (N_9042,N_8942,N_8952);
nor U9043 (N_9043,N_8692,N_8943);
or U9044 (N_9044,N_8524,N_8632);
or U9045 (N_9045,N_8725,N_8839);
nor U9046 (N_9046,N_8563,N_8828);
xnor U9047 (N_9047,N_8700,N_8629);
xor U9048 (N_9048,N_8694,N_8566);
nand U9049 (N_9049,N_8906,N_8887);
or U9050 (N_9050,N_8560,N_8926);
nand U9051 (N_9051,N_8734,N_8817);
nand U9052 (N_9052,N_8914,N_8757);
xor U9053 (N_9053,N_8575,N_8849);
nand U9054 (N_9054,N_8767,N_8963);
or U9055 (N_9055,N_8539,N_8872);
nor U9056 (N_9056,N_8776,N_8973);
or U9057 (N_9057,N_8643,N_8630);
nand U9058 (N_9058,N_8791,N_8590);
xnor U9059 (N_9059,N_8514,N_8845);
nor U9060 (N_9060,N_8904,N_8889);
nor U9061 (N_9061,N_8979,N_8534);
and U9062 (N_9062,N_8855,N_8785);
nor U9063 (N_9063,N_8804,N_8593);
xor U9064 (N_9064,N_8655,N_8625);
nand U9065 (N_9065,N_8706,N_8878);
and U9066 (N_9066,N_8620,N_8607);
and U9067 (N_9067,N_8518,N_8707);
nand U9068 (N_9068,N_8899,N_8683);
or U9069 (N_9069,N_8937,N_8689);
and U9070 (N_9070,N_8506,N_8760);
and U9071 (N_9071,N_8893,N_8596);
xnor U9072 (N_9072,N_8682,N_8759);
or U9073 (N_9073,N_8568,N_8714);
and U9074 (N_9074,N_8564,N_8832);
xnor U9075 (N_9075,N_8595,N_8634);
and U9076 (N_9076,N_8635,N_8588);
xnor U9077 (N_9077,N_8951,N_8520);
nand U9078 (N_9078,N_8907,N_8751);
nor U9079 (N_9079,N_8820,N_8834);
and U9080 (N_9080,N_8853,N_8980);
and U9081 (N_9081,N_8713,N_8663);
and U9082 (N_9082,N_8724,N_8984);
or U9083 (N_9083,N_8551,N_8719);
and U9084 (N_9084,N_8668,N_8511);
and U9085 (N_9085,N_8765,N_8729);
and U9086 (N_9086,N_8838,N_8718);
xor U9087 (N_9087,N_8690,N_8679);
nand U9088 (N_9088,N_8971,N_8637);
xnor U9089 (N_9089,N_8540,N_8925);
or U9090 (N_9090,N_8976,N_8837);
nor U9091 (N_9091,N_8633,N_8898);
xor U9092 (N_9092,N_8764,N_8809);
nor U9093 (N_9093,N_8991,N_8763);
and U9094 (N_9094,N_8781,N_8555);
nor U9095 (N_9095,N_8772,N_8917);
nand U9096 (N_9096,N_8742,N_8631);
nor U9097 (N_9097,N_8676,N_8665);
or U9098 (N_9098,N_8577,N_8975);
nand U9099 (N_9099,N_8603,N_8609);
nand U9100 (N_9100,N_8996,N_8761);
or U9101 (N_9101,N_8769,N_8646);
nor U9102 (N_9102,N_8934,N_8667);
nor U9103 (N_9103,N_8510,N_8652);
xnor U9104 (N_9104,N_8574,N_8891);
or U9105 (N_9105,N_8940,N_8752);
nor U9106 (N_9106,N_8771,N_8827);
nand U9107 (N_9107,N_8923,N_8519);
nand U9108 (N_9108,N_8826,N_8902);
xor U9109 (N_9109,N_8688,N_8517);
nor U9110 (N_9110,N_8846,N_8867);
xor U9111 (N_9111,N_8915,N_8735);
nor U9112 (N_9112,N_8553,N_8636);
and U9113 (N_9113,N_8787,N_8792);
nand U9114 (N_9114,N_8521,N_8597);
xor U9115 (N_9115,N_8567,N_8600);
xor U9116 (N_9116,N_8547,N_8645);
nor U9117 (N_9117,N_8786,N_8545);
and U9118 (N_9118,N_8788,N_8956);
xnor U9119 (N_9119,N_8779,N_8644);
nand U9120 (N_9120,N_8622,N_8508);
nand U9121 (N_9121,N_8947,N_8978);
nor U9122 (N_9122,N_8598,N_8585);
or U9123 (N_9123,N_8666,N_8847);
or U9124 (N_9124,N_8501,N_8790);
and U9125 (N_9125,N_8935,N_8628);
or U9126 (N_9126,N_8982,N_8569);
nor U9127 (N_9127,N_8842,N_8621);
xor U9128 (N_9128,N_8916,N_8571);
xnor U9129 (N_9129,N_8946,N_8531);
nand U9130 (N_9130,N_8687,N_8933);
or U9131 (N_9131,N_8863,N_8664);
and U9132 (N_9132,N_8589,N_8866);
xnor U9133 (N_9133,N_8723,N_8680);
and U9134 (N_9134,N_8703,N_8758);
nand U9135 (N_9135,N_8901,N_8573);
or U9136 (N_9136,N_8932,N_8848);
xor U9137 (N_9137,N_8747,N_8716);
or U9138 (N_9138,N_8784,N_8881);
and U9139 (N_9139,N_8592,N_8594);
and U9140 (N_9140,N_8921,N_8890);
nand U9141 (N_9141,N_8552,N_8983);
and U9142 (N_9142,N_8823,N_8966);
nor U9143 (N_9143,N_8910,N_8614);
and U9144 (N_9144,N_8957,N_8773);
and U9145 (N_9145,N_8720,N_8850);
xnor U9146 (N_9146,N_8710,N_8526);
and U9147 (N_9147,N_8619,N_8858);
or U9148 (N_9148,N_8794,N_8653);
and U9149 (N_9149,N_8542,N_8918);
nand U9150 (N_9150,N_8836,N_8662);
xor U9151 (N_9151,N_8861,N_8500);
or U9152 (N_9152,N_8702,N_8615);
xor U9153 (N_9153,N_8777,N_8748);
or U9154 (N_9154,N_8572,N_8799);
nand U9155 (N_9155,N_8819,N_8919);
nor U9156 (N_9156,N_8557,N_8985);
or U9157 (N_9157,N_8638,N_8657);
nand U9158 (N_9158,N_8746,N_8728);
xnor U9159 (N_9159,N_8660,N_8648);
nand U9160 (N_9160,N_8783,N_8533);
nand U9161 (N_9161,N_8505,N_8840);
nor U9162 (N_9162,N_8964,N_8801);
and U9163 (N_9163,N_8528,N_8651);
nor U9164 (N_9164,N_8869,N_8579);
and U9165 (N_9165,N_8989,N_8807);
or U9166 (N_9166,N_8802,N_8712);
and U9167 (N_9167,N_8803,N_8905);
nor U9168 (N_9168,N_8955,N_8587);
nand U9169 (N_9169,N_8699,N_8558);
and U9170 (N_9170,N_8623,N_8774);
xor U9171 (N_9171,N_8602,N_8894);
or U9172 (N_9172,N_8693,N_8830);
nor U9173 (N_9173,N_8997,N_8586);
and U9174 (N_9174,N_8775,N_8576);
nor U9175 (N_9175,N_8762,N_8755);
nand U9176 (N_9176,N_8522,N_8580);
nand U9177 (N_9177,N_8865,N_8974);
xor U9178 (N_9178,N_8949,N_8695);
xnor U9179 (N_9179,N_8717,N_8909);
or U9180 (N_9180,N_8559,N_8844);
or U9181 (N_9181,N_8948,N_8859);
xor U9182 (N_9182,N_8884,N_8674);
or U9183 (N_9183,N_8601,N_8738);
xnor U9184 (N_9184,N_8911,N_8986);
or U9185 (N_9185,N_8736,N_8860);
and U9186 (N_9186,N_8578,N_8502);
or U9187 (N_9187,N_8961,N_8509);
nor U9188 (N_9188,N_8504,N_8851);
nor U9189 (N_9189,N_8864,N_8715);
and U9190 (N_9190,N_8903,N_8727);
or U9191 (N_9191,N_8871,N_8570);
nor U9192 (N_9192,N_8722,N_8912);
nand U9193 (N_9193,N_8721,N_8642);
or U9194 (N_9194,N_8750,N_8927);
nand U9195 (N_9195,N_8931,N_8639);
nor U9196 (N_9196,N_8527,N_8798);
or U9197 (N_9197,N_8883,N_8624);
nand U9198 (N_9198,N_8972,N_8554);
nor U9199 (N_9199,N_8822,N_8913);
xnor U9200 (N_9200,N_8684,N_8793);
nand U9201 (N_9201,N_8797,N_8749);
nand U9202 (N_9202,N_8549,N_8892);
and U9203 (N_9203,N_8768,N_8709);
and U9204 (N_9204,N_8641,N_8696);
or U9205 (N_9205,N_8990,N_8583);
nand U9206 (N_9206,N_8670,N_8678);
xnor U9207 (N_9207,N_8739,N_8546);
nand U9208 (N_9208,N_8812,N_8795);
nor U9209 (N_9209,N_8960,N_8732);
nor U9210 (N_9210,N_8950,N_8550);
xor U9211 (N_9211,N_8811,N_8944);
nand U9212 (N_9212,N_8705,N_8640);
or U9213 (N_9213,N_8857,N_8766);
or U9214 (N_9214,N_8879,N_8862);
and U9215 (N_9215,N_8810,N_8789);
nand U9216 (N_9216,N_8877,N_8780);
and U9217 (N_9217,N_8800,N_8541);
xor U9218 (N_9218,N_8953,N_8626);
xnor U9219 (N_9219,N_8929,N_8922);
or U9220 (N_9220,N_8512,N_8928);
nand U9221 (N_9221,N_8726,N_8969);
nand U9222 (N_9222,N_8731,N_8873);
nand U9223 (N_9223,N_8885,N_8954);
nor U9224 (N_9224,N_8992,N_8962);
and U9225 (N_9225,N_8532,N_8608);
or U9226 (N_9226,N_8565,N_8672);
nand U9227 (N_9227,N_8778,N_8677);
nand U9228 (N_9228,N_8835,N_8741);
or U9229 (N_9229,N_8994,N_8930);
nor U9230 (N_9230,N_8938,N_8649);
and U9231 (N_9231,N_8977,N_8841);
or U9232 (N_9232,N_8658,N_8525);
and U9233 (N_9233,N_8993,N_8610);
nand U9234 (N_9234,N_8818,N_8591);
or U9235 (N_9235,N_8856,N_8538);
or U9236 (N_9236,N_8507,N_8816);
nor U9237 (N_9237,N_8908,N_8833);
and U9238 (N_9238,N_8814,N_8874);
or U9239 (N_9239,N_8740,N_8939);
nor U9240 (N_9240,N_8599,N_8965);
nand U9241 (N_9241,N_8561,N_8673);
nor U9242 (N_9242,N_8604,N_8743);
nor U9243 (N_9243,N_8886,N_8675);
or U9244 (N_9244,N_8753,N_8970);
or U9245 (N_9245,N_8698,N_8821);
or U9246 (N_9246,N_8671,N_8691);
nor U9247 (N_9247,N_8808,N_8537);
nand U9248 (N_9248,N_8995,N_8656);
nor U9249 (N_9249,N_8967,N_8924);
nand U9250 (N_9250,N_8536,N_8517);
nand U9251 (N_9251,N_8729,N_8934);
nand U9252 (N_9252,N_8793,N_8716);
and U9253 (N_9253,N_8828,N_8509);
or U9254 (N_9254,N_8653,N_8508);
and U9255 (N_9255,N_8692,N_8781);
nand U9256 (N_9256,N_8781,N_8954);
nand U9257 (N_9257,N_8962,N_8738);
or U9258 (N_9258,N_8765,N_8758);
xor U9259 (N_9259,N_8709,N_8997);
and U9260 (N_9260,N_8809,N_8820);
xor U9261 (N_9261,N_8604,N_8734);
xor U9262 (N_9262,N_8547,N_8960);
xor U9263 (N_9263,N_8533,N_8573);
and U9264 (N_9264,N_8693,N_8869);
and U9265 (N_9265,N_8577,N_8942);
nand U9266 (N_9266,N_8977,N_8531);
nand U9267 (N_9267,N_8586,N_8905);
and U9268 (N_9268,N_8802,N_8644);
xor U9269 (N_9269,N_8997,N_8673);
xor U9270 (N_9270,N_8584,N_8602);
xnor U9271 (N_9271,N_8871,N_8534);
nand U9272 (N_9272,N_8523,N_8565);
nand U9273 (N_9273,N_8912,N_8778);
or U9274 (N_9274,N_8918,N_8968);
nor U9275 (N_9275,N_8601,N_8908);
nand U9276 (N_9276,N_8584,N_8787);
or U9277 (N_9277,N_8991,N_8841);
nor U9278 (N_9278,N_8554,N_8643);
or U9279 (N_9279,N_8754,N_8972);
nand U9280 (N_9280,N_8566,N_8916);
or U9281 (N_9281,N_8700,N_8840);
xnor U9282 (N_9282,N_8926,N_8672);
nor U9283 (N_9283,N_8967,N_8926);
nor U9284 (N_9284,N_8704,N_8812);
nor U9285 (N_9285,N_8874,N_8627);
and U9286 (N_9286,N_8736,N_8799);
and U9287 (N_9287,N_8638,N_8795);
nand U9288 (N_9288,N_8938,N_8508);
nor U9289 (N_9289,N_8814,N_8741);
nand U9290 (N_9290,N_8786,N_8631);
or U9291 (N_9291,N_8743,N_8974);
and U9292 (N_9292,N_8620,N_8940);
nor U9293 (N_9293,N_8781,N_8851);
nand U9294 (N_9294,N_8996,N_8780);
xor U9295 (N_9295,N_8809,N_8742);
or U9296 (N_9296,N_8819,N_8668);
or U9297 (N_9297,N_8926,N_8951);
nand U9298 (N_9298,N_8689,N_8731);
xnor U9299 (N_9299,N_8629,N_8887);
nor U9300 (N_9300,N_8624,N_8686);
nand U9301 (N_9301,N_8561,N_8848);
nand U9302 (N_9302,N_8941,N_8823);
and U9303 (N_9303,N_8577,N_8746);
nand U9304 (N_9304,N_8613,N_8777);
or U9305 (N_9305,N_8978,N_8986);
nand U9306 (N_9306,N_8535,N_8702);
or U9307 (N_9307,N_8575,N_8545);
nor U9308 (N_9308,N_8833,N_8579);
and U9309 (N_9309,N_8627,N_8711);
nand U9310 (N_9310,N_8722,N_8562);
or U9311 (N_9311,N_8979,N_8959);
nand U9312 (N_9312,N_8924,N_8540);
xnor U9313 (N_9313,N_8917,N_8852);
nor U9314 (N_9314,N_8562,N_8581);
nor U9315 (N_9315,N_8937,N_8998);
or U9316 (N_9316,N_8563,N_8800);
and U9317 (N_9317,N_8691,N_8709);
and U9318 (N_9318,N_8879,N_8669);
nand U9319 (N_9319,N_8602,N_8853);
nand U9320 (N_9320,N_8858,N_8552);
or U9321 (N_9321,N_8874,N_8748);
xor U9322 (N_9322,N_8972,N_8979);
or U9323 (N_9323,N_8888,N_8636);
xnor U9324 (N_9324,N_8841,N_8571);
and U9325 (N_9325,N_8661,N_8573);
or U9326 (N_9326,N_8932,N_8736);
xor U9327 (N_9327,N_8595,N_8878);
or U9328 (N_9328,N_8688,N_8511);
nor U9329 (N_9329,N_8568,N_8792);
nor U9330 (N_9330,N_8588,N_8924);
or U9331 (N_9331,N_8984,N_8667);
nand U9332 (N_9332,N_8801,N_8804);
nand U9333 (N_9333,N_8826,N_8727);
xnor U9334 (N_9334,N_8949,N_8901);
or U9335 (N_9335,N_8520,N_8925);
xnor U9336 (N_9336,N_8985,N_8509);
nor U9337 (N_9337,N_8960,N_8715);
nand U9338 (N_9338,N_8969,N_8569);
nor U9339 (N_9339,N_8596,N_8974);
nor U9340 (N_9340,N_8500,N_8953);
and U9341 (N_9341,N_8762,N_8655);
nand U9342 (N_9342,N_8757,N_8617);
nor U9343 (N_9343,N_8603,N_8858);
and U9344 (N_9344,N_8876,N_8725);
and U9345 (N_9345,N_8734,N_8833);
or U9346 (N_9346,N_8708,N_8745);
or U9347 (N_9347,N_8942,N_8905);
nand U9348 (N_9348,N_8909,N_8855);
nand U9349 (N_9349,N_8868,N_8902);
or U9350 (N_9350,N_8674,N_8560);
nor U9351 (N_9351,N_8538,N_8740);
or U9352 (N_9352,N_8852,N_8945);
nand U9353 (N_9353,N_8537,N_8866);
nand U9354 (N_9354,N_8851,N_8538);
and U9355 (N_9355,N_8722,N_8822);
nand U9356 (N_9356,N_8898,N_8913);
and U9357 (N_9357,N_8577,N_8540);
or U9358 (N_9358,N_8682,N_8931);
or U9359 (N_9359,N_8850,N_8537);
or U9360 (N_9360,N_8526,N_8578);
nand U9361 (N_9361,N_8934,N_8662);
xnor U9362 (N_9362,N_8669,N_8766);
nor U9363 (N_9363,N_8882,N_8554);
and U9364 (N_9364,N_8965,N_8624);
nand U9365 (N_9365,N_8903,N_8869);
and U9366 (N_9366,N_8515,N_8688);
xnor U9367 (N_9367,N_8993,N_8830);
nor U9368 (N_9368,N_8993,N_8606);
xor U9369 (N_9369,N_8865,N_8791);
nor U9370 (N_9370,N_8821,N_8581);
and U9371 (N_9371,N_8879,N_8857);
nor U9372 (N_9372,N_8988,N_8603);
xor U9373 (N_9373,N_8539,N_8897);
xnor U9374 (N_9374,N_8929,N_8743);
or U9375 (N_9375,N_8647,N_8912);
and U9376 (N_9376,N_8956,N_8847);
and U9377 (N_9377,N_8870,N_8539);
nor U9378 (N_9378,N_8932,N_8858);
nand U9379 (N_9379,N_8889,N_8756);
or U9380 (N_9380,N_8799,N_8529);
or U9381 (N_9381,N_8778,N_8820);
nor U9382 (N_9382,N_8992,N_8656);
nor U9383 (N_9383,N_8517,N_8716);
nand U9384 (N_9384,N_8719,N_8575);
and U9385 (N_9385,N_8859,N_8839);
nor U9386 (N_9386,N_8993,N_8552);
nor U9387 (N_9387,N_8535,N_8994);
or U9388 (N_9388,N_8924,N_8509);
nand U9389 (N_9389,N_8503,N_8710);
xnor U9390 (N_9390,N_8872,N_8773);
nand U9391 (N_9391,N_8787,N_8865);
nand U9392 (N_9392,N_8800,N_8750);
and U9393 (N_9393,N_8658,N_8641);
nor U9394 (N_9394,N_8629,N_8528);
xor U9395 (N_9395,N_8906,N_8690);
and U9396 (N_9396,N_8812,N_8867);
nand U9397 (N_9397,N_8606,N_8845);
nor U9398 (N_9398,N_8755,N_8923);
xnor U9399 (N_9399,N_8891,N_8860);
nand U9400 (N_9400,N_8613,N_8857);
xor U9401 (N_9401,N_8541,N_8615);
and U9402 (N_9402,N_8784,N_8947);
xor U9403 (N_9403,N_8916,N_8529);
nand U9404 (N_9404,N_8650,N_8950);
nand U9405 (N_9405,N_8632,N_8579);
nor U9406 (N_9406,N_8931,N_8663);
and U9407 (N_9407,N_8728,N_8692);
and U9408 (N_9408,N_8723,N_8942);
xor U9409 (N_9409,N_8933,N_8828);
xnor U9410 (N_9410,N_8783,N_8994);
nand U9411 (N_9411,N_8901,N_8722);
and U9412 (N_9412,N_8998,N_8698);
nor U9413 (N_9413,N_8908,N_8708);
nand U9414 (N_9414,N_8510,N_8981);
or U9415 (N_9415,N_8874,N_8933);
and U9416 (N_9416,N_8885,N_8689);
xnor U9417 (N_9417,N_8777,N_8591);
xnor U9418 (N_9418,N_8989,N_8770);
nand U9419 (N_9419,N_8680,N_8749);
xnor U9420 (N_9420,N_8830,N_8966);
nor U9421 (N_9421,N_8819,N_8776);
and U9422 (N_9422,N_8916,N_8756);
nand U9423 (N_9423,N_8764,N_8666);
or U9424 (N_9424,N_8572,N_8842);
nand U9425 (N_9425,N_8969,N_8735);
or U9426 (N_9426,N_8698,N_8668);
nand U9427 (N_9427,N_8815,N_8753);
nand U9428 (N_9428,N_8537,N_8882);
or U9429 (N_9429,N_8905,N_8679);
nand U9430 (N_9430,N_8987,N_8745);
xor U9431 (N_9431,N_8750,N_8846);
nor U9432 (N_9432,N_8954,N_8552);
xnor U9433 (N_9433,N_8887,N_8771);
or U9434 (N_9434,N_8777,N_8906);
nand U9435 (N_9435,N_8839,N_8797);
xnor U9436 (N_9436,N_8804,N_8631);
or U9437 (N_9437,N_8798,N_8558);
nand U9438 (N_9438,N_8613,N_8737);
xor U9439 (N_9439,N_8604,N_8817);
nor U9440 (N_9440,N_8795,N_8672);
xor U9441 (N_9441,N_8872,N_8881);
or U9442 (N_9442,N_8813,N_8781);
nand U9443 (N_9443,N_8564,N_8517);
or U9444 (N_9444,N_8804,N_8857);
xor U9445 (N_9445,N_8783,N_8885);
nor U9446 (N_9446,N_8926,N_8849);
nand U9447 (N_9447,N_8795,N_8862);
nor U9448 (N_9448,N_8801,N_8596);
nor U9449 (N_9449,N_8936,N_8864);
xnor U9450 (N_9450,N_8957,N_8995);
xnor U9451 (N_9451,N_8530,N_8591);
or U9452 (N_9452,N_8687,N_8639);
nor U9453 (N_9453,N_8864,N_8837);
xor U9454 (N_9454,N_8849,N_8761);
or U9455 (N_9455,N_8712,N_8797);
nand U9456 (N_9456,N_8949,N_8744);
and U9457 (N_9457,N_8512,N_8775);
and U9458 (N_9458,N_8587,N_8691);
and U9459 (N_9459,N_8760,N_8680);
or U9460 (N_9460,N_8828,N_8746);
or U9461 (N_9461,N_8544,N_8530);
nor U9462 (N_9462,N_8759,N_8536);
nor U9463 (N_9463,N_8775,N_8800);
nor U9464 (N_9464,N_8961,N_8867);
xnor U9465 (N_9465,N_8739,N_8772);
xnor U9466 (N_9466,N_8661,N_8675);
xor U9467 (N_9467,N_8941,N_8966);
nand U9468 (N_9468,N_8550,N_8528);
nand U9469 (N_9469,N_8739,N_8673);
nor U9470 (N_9470,N_8985,N_8805);
xor U9471 (N_9471,N_8700,N_8619);
and U9472 (N_9472,N_8733,N_8802);
and U9473 (N_9473,N_8655,N_8574);
or U9474 (N_9474,N_8618,N_8580);
and U9475 (N_9475,N_8985,N_8786);
nor U9476 (N_9476,N_8540,N_8930);
nor U9477 (N_9477,N_8699,N_8507);
and U9478 (N_9478,N_8616,N_8661);
or U9479 (N_9479,N_8534,N_8890);
and U9480 (N_9480,N_8719,N_8664);
xor U9481 (N_9481,N_8573,N_8647);
or U9482 (N_9482,N_8859,N_8891);
or U9483 (N_9483,N_8672,N_8617);
xnor U9484 (N_9484,N_8586,N_8888);
and U9485 (N_9485,N_8855,N_8957);
nand U9486 (N_9486,N_8579,N_8948);
and U9487 (N_9487,N_8962,N_8977);
nor U9488 (N_9488,N_8677,N_8918);
xor U9489 (N_9489,N_8510,N_8630);
nor U9490 (N_9490,N_8728,N_8766);
xnor U9491 (N_9491,N_8613,N_8871);
and U9492 (N_9492,N_8994,N_8551);
or U9493 (N_9493,N_8566,N_8513);
and U9494 (N_9494,N_8825,N_8749);
or U9495 (N_9495,N_8540,N_8884);
nor U9496 (N_9496,N_8894,N_8693);
nand U9497 (N_9497,N_8561,N_8690);
or U9498 (N_9498,N_8836,N_8528);
or U9499 (N_9499,N_8801,N_8832);
or U9500 (N_9500,N_9047,N_9257);
nand U9501 (N_9501,N_9125,N_9219);
nand U9502 (N_9502,N_9068,N_9372);
or U9503 (N_9503,N_9317,N_9324);
xnor U9504 (N_9504,N_9353,N_9398);
nor U9505 (N_9505,N_9164,N_9170);
or U9506 (N_9506,N_9156,N_9109);
nor U9507 (N_9507,N_9344,N_9176);
nor U9508 (N_9508,N_9100,N_9306);
and U9509 (N_9509,N_9333,N_9104);
xnor U9510 (N_9510,N_9387,N_9319);
nor U9511 (N_9511,N_9115,N_9172);
xnor U9512 (N_9512,N_9098,N_9197);
nand U9513 (N_9513,N_9152,N_9392);
and U9514 (N_9514,N_9106,N_9498);
or U9515 (N_9515,N_9182,N_9339);
and U9516 (N_9516,N_9243,N_9013);
nand U9517 (N_9517,N_9433,N_9454);
and U9518 (N_9518,N_9332,N_9383);
or U9519 (N_9519,N_9292,N_9211);
and U9520 (N_9520,N_9058,N_9289);
or U9521 (N_9521,N_9015,N_9034);
xnor U9522 (N_9522,N_9120,N_9088);
xor U9523 (N_9523,N_9030,N_9412);
xnor U9524 (N_9524,N_9010,N_9204);
xor U9525 (N_9525,N_9329,N_9137);
and U9526 (N_9526,N_9143,N_9468);
and U9527 (N_9527,N_9029,N_9420);
nand U9528 (N_9528,N_9441,N_9256);
and U9529 (N_9529,N_9379,N_9128);
and U9530 (N_9530,N_9483,N_9139);
nor U9531 (N_9531,N_9496,N_9476);
nor U9532 (N_9532,N_9192,N_9040);
xor U9533 (N_9533,N_9002,N_9434);
and U9534 (N_9534,N_9178,N_9318);
nand U9535 (N_9535,N_9416,N_9028);
or U9536 (N_9536,N_9325,N_9421);
xor U9537 (N_9537,N_9304,N_9271);
and U9538 (N_9538,N_9432,N_9484);
xor U9539 (N_9539,N_9313,N_9233);
or U9540 (N_9540,N_9050,N_9117);
nand U9541 (N_9541,N_9356,N_9262);
nor U9542 (N_9542,N_9165,N_9019);
nand U9543 (N_9543,N_9275,N_9198);
nand U9544 (N_9544,N_9354,N_9190);
nand U9545 (N_9545,N_9005,N_9186);
nor U9546 (N_9546,N_9393,N_9049);
nand U9547 (N_9547,N_9337,N_9369);
nand U9548 (N_9548,N_9457,N_9250);
nor U9549 (N_9549,N_9495,N_9288);
xnor U9550 (N_9550,N_9024,N_9223);
nand U9551 (N_9551,N_9236,N_9061);
nor U9552 (N_9552,N_9200,N_9373);
or U9553 (N_9553,N_9487,N_9396);
and U9554 (N_9554,N_9453,N_9406);
xnor U9555 (N_9555,N_9048,N_9229);
nor U9556 (N_9556,N_9394,N_9096);
nand U9557 (N_9557,N_9105,N_9064);
and U9558 (N_9558,N_9132,N_9103);
xor U9559 (N_9559,N_9239,N_9153);
and U9560 (N_9560,N_9224,N_9006);
and U9561 (N_9561,N_9264,N_9479);
nand U9562 (N_9562,N_9126,N_9267);
xor U9563 (N_9563,N_9142,N_9003);
and U9564 (N_9564,N_9499,N_9308);
xnor U9565 (N_9565,N_9447,N_9436);
nand U9566 (N_9566,N_9361,N_9080);
xor U9567 (N_9567,N_9382,N_9466);
nor U9568 (N_9568,N_9145,N_9187);
and U9569 (N_9569,N_9340,N_9241);
xor U9570 (N_9570,N_9357,N_9450);
nand U9571 (N_9571,N_9148,N_9222);
nand U9572 (N_9572,N_9491,N_9280);
or U9573 (N_9573,N_9252,N_9465);
nor U9574 (N_9574,N_9168,N_9135);
xnor U9575 (N_9575,N_9166,N_9471);
nand U9576 (N_9576,N_9448,N_9044);
nor U9577 (N_9577,N_9138,N_9221);
nor U9578 (N_9578,N_9431,N_9331);
nor U9579 (N_9579,N_9062,N_9012);
or U9580 (N_9580,N_9458,N_9116);
xor U9581 (N_9581,N_9149,N_9268);
nor U9582 (N_9582,N_9059,N_9171);
xor U9583 (N_9583,N_9445,N_9076);
or U9584 (N_9584,N_9490,N_9060);
or U9585 (N_9585,N_9282,N_9428);
nor U9586 (N_9586,N_9234,N_9402);
xnor U9587 (N_9587,N_9326,N_9123);
nand U9588 (N_9588,N_9131,N_9111);
or U9589 (N_9589,N_9364,N_9460);
or U9590 (N_9590,N_9461,N_9036);
and U9591 (N_9591,N_9492,N_9322);
xor U9592 (N_9592,N_9134,N_9427);
xnor U9593 (N_9593,N_9193,N_9053);
nand U9594 (N_9594,N_9009,N_9199);
nand U9595 (N_9595,N_9079,N_9440);
nand U9596 (N_9596,N_9423,N_9281);
nor U9597 (N_9597,N_9422,N_9063);
and U9598 (N_9598,N_9384,N_9191);
nand U9599 (N_9599,N_9136,N_9194);
nor U9600 (N_9600,N_9147,N_9218);
nand U9601 (N_9601,N_9403,N_9269);
xnor U9602 (N_9602,N_9312,N_9278);
nand U9603 (N_9603,N_9494,N_9022);
xnor U9604 (N_9604,N_9426,N_9266);
nor U9605 (N_9605,N_9245,N_9251);
nor U9606 (N_9606,N_9464,N_9341);
or U9607 (N_9607,N_9263,N_9247);
nand U9608 (N_9608,N_9163,N_9158);
or U9609 (N_9609,N_9021,N_9203);
nand U9610 (N_9610,N_9150,N_9456);
and U9611 (N_9611,N_9375,N_9154);
nand U9612 (N_9612,N_9349,N_9127);
or U9613 (N_9613,N_9213,N_9342);
xnor U9614 (N_9614,N_9184,N_9430);
or U9615 (N_9615,N_9246,N_9347);
nand U9616 (N_9616,N_9374,N_9284);
xor U9617 (N_9617,N_9195,N_9489);
nand U9618 (N_9618,N_9321,N_9473);
xnor U9619 (N_9619,N_9056,N_9214);
xnor U9620 (N_9620,N_9305,N_9386);
xor U9621 (N_9621,N_9451,N_9411);
and U9622 (N_9622,N_9160,N_9260);
xnor U9623 (N_9623,N_9437,N_9419);
and U9624 (N_9624,N_9087,N_9107);
and U9625 (N_9625,N_9385,N_9343);
or U9626 (N_9626,N_9316,N_9455);
or U9627 (N_9627,N_9352,N_9039);
xnor U9628 (N_9628,N_9405,N_9391);
or U9629 (N_9629,N_9378,N_9082);
and U9630 (N_9630,N_9007,N_9418);
nand U9631 (N_9631,N_9114,N_9231);
nor U9632 (N_9632,N_9274,N_9415);
nand U9633 (N_9633,N_9424,N_9095);
xor U9634 (N_9634,N_9046,N_9057);
and U9635 (N_9635,N_9031,N_9181);
and U9636 (N_9636,N_9389,N_9151);
xor U9637 (N_9637,N_9071,N_9279);
nor U9638 (N_9638,N_9066,N_9488);
and U9639 (N_9639,N_9314,N_9225);
and U9640 (N_9640,N_9067,N_9146);
xor U9641 (N_9641,N_9359,N_9025);
nand U9642 (N_9642,N_9452,N_9435);
xnor U9643 (N_9643,N_9085,N_9482);
xnor U9644 (N_9644,N_9065,N_9101);
xnor U9645 (N_9645,N_9303,N_9099);
and U9646 (N_9646,N_9043,N_9237);
or U9647 (N_9647,N_9444,N_9122);
nand U9648 (N_9648,N_9177,N_9409);
nand U9649 (N_9649,N_9390,N_9072);
nand U9650 (N_9650,N_9365,N_9259);
xnor U9651 (N_9651,N_9320,N_9188);
or U9652 (N_9652,N_9074,N_9206);
xor U9653 (N_9653,N_9173,N_9345);
or U9654 (N_9654,N_9472,N_9368);
nor U9655 (N_9655,N_9220,N_9091);
nand U9656 (N_9656,N_9377,N_9285);
xor U9657 (N_9657,N_9293,N_9346);
nand U9658 (N_9658,N_9073,N_9486);
xnor U9659 (N_9659,N_9351,N_9011);
nor U9660 (N_9660,N_9210,N_9118);
nand U9661 (N_9661,N_9032,N_9429);
or U9662 (N_9662,N_9481,N_9283);
or U9663 (N_9663,N_9254,N_9446);
and U9664 (N_9664,N_9045,N_9334);
or U9665 (N_9665,N_9008,N_9407);
nor U9666 (N_9666,N_9227,N_9035);
nor U9667 (N_9667,N_9277,N_9235);
and U9668 (N_9668,N_9242,N_9478);
xor U9669 (N_9669,N_9238,N_9090);
nor U9670 (N_9670,N_9020,N_9215);
xnor U9671 (N_9671,N_9110,N_9205);
and U9672 (N_9672,N_9108,N_9302);
nand U9673 (N_9673,N_9119,N_9404);
nor U9674 (N_9674,N_9474,N_9033);
or U9675 (N_9675,N_9381,N_9323);
nor U9676 (N_9676,N_9093,N_9000);
xor U9677 (N_9677,N_9086,N_9417);
or U9678 (N_9678,N_9443,N_9161);
nor U9679 (N_9679,N_9371,N_9439);
xor U9680 (N_9680,N_9023,N_9477);
nand U9681 (N_9681,N_9270,N_9395);
nand U9682 (N_9682,N_9497,N_9399);
or U9683 (N_9683,N_9244,N_9232);
or U9684 (N_9684,N_9094,N_9300);
nor U9685 (N_9685,N_9363,N_9207);
nor U9686 (N_9686,N_9249,N_9202);
xor U9687 (N_9687,N_9141,N_9258);
and U9688 (N_9688,N_9130,N_9348);
nor U9689 (N_9689,N_9097,N_9027);
xor U9690 (N_9690,N_9366,N_9400);
xnor U9691 (N_9691,N_9248,N_9299);
nand U9692 (N_9692,N_9330,N_9286);
xor U9693 (N_9693,N_9408,N_9273);
or U9694 (N_9694,N_9179,N_9467);
or U9695 (N_9695,N_9480,N_9388);
nand U9696 (N_9696,N_9121,N_9493);
xor U9697 (N_9697,N_9307,N_9016);
xnor U9698 (N_9698,N_9102,N_9189);
and U9699 (N_9699,N_9212,N_9310);
and U9700 (N_9700,N_9078,N_9183);
nor U9701 (N_9701,N_9018,N_9442);
nand U9702 (N_9702,N_9240,N_9077);
and U9703 (N_9703,N_9376,N_9084);
xor U9704 (N_9704,N_9401,N_9296);
or U9705 (N_9705,N_9265,N_9175);
xnor U9706 (N_9706,N_9475,N_9038);
and U9707 (N_9707,N_9004,N_9459);
nor U9708 (N_9708,N_9253,N_9014);
and U9709 (N_9709,N_9124,N_9272);
xnor U9710 (N_9710,N_9276,N_9230);
nand U9711 (N_9711,N_9338,N_9054);
or U9712 (N_9712,N_9350,N_9336);
xnor U9713 (N_9713,N_9162,N_9055);
or U9714 (N_9714,N_9185,N_9140);
nand U9715 (N_9715,N_9089,N_9261);
nand U9716 (N_9716,N_9425,N_9037);
and U9717 (N_9717,N_9169,N_9026);
nor U9718 (N_9718,N_9209,N_9463);
nand U9719 (N_9719,N_9397,N_9414);
or U9720 (N_9720,N_9133,N_9255);
and U9721 (N_9721,N_9410,N_9155);
and U9722 (N_9722,N_9327,N_9129);
or U9723 (N_9723,N_9294,N_9113);
or U9724 (N_9724,N_9070,N_9167);
or U9725 (N_9725,N_9297,N_9355);
xnor U9726 (N_9726,N_9298,N_9083);
nand U9727 (N_9727,N_9069,N_9081);
nor U9728 (N_9728,N_9052,N_9112);
nor U9729 (N_9729,N_9208,N_9217);
nand U9730 (N_9730,N_9075,N_9226);
nand U9731 (N_9731,N_9228,N_9367);
or U9732 (N_9732,N_9201,N_9291);
nand U9733 (N_9733,N_9216,N_9295);
xnor U9734 (N_9734,N_9196,N_9180);
and U9735 (N_9735,N_9485,N_9438);
nor U9736 (N_9736,N_9157,N_9335);
nor U9737 (N_9737,N_9362,N_9360);
and U9738 (N_9738,N_9358,N_9315);
nand U9739 (N_9739,N_9001,N_9413);
nor U9740 (N_9740,N_9301,N_9051);
nor U9741 (N_9741,N_9174,N_9042);
and U9742 (N_9742,N_9092,N_9328);
xor U9743 (N_9743,N_9041,N_9290);
and U9744 (N_9744,N_9159,N_9469);
nand U9745 (N_9745,N_9470,N_9370);
nand U9746 (N_9746,N_9017,N_9287);
or U9747 (N_9747,N_9311,N_9144);
nand U9748 (N_9748,N_9380,N_9309);
nor U9749 (N_9749,N_9462,N_9449);
nor U9750 (N_9750,N_9011,N_9110);
xnor U9751 (N_9751,N_9375,N_9394);
nand U9752 (N_9752,N_9272,N_9156);
and U9753 (N_9753,N_9266,N_9456);
xor U9754 (N_9754,N_9106,N_9227);
and U9755 (N_9755,N_9129,N_9462);
nand U9756 (N_9756,N_9344,N_9189);
or U9757 (N_9757,N_9156,N_9203);
nand U9758 (N_9758,N_9319,N_9075);
or U9759 (N_9759,N_9007,N_9325);
and U9760 (N_9760,N_9299,N_9308);
nand U9761 (N_9761,N_9317,N_9261);
nor U9762 (N_9762,N_9495,N_9341);
nand U9763 (N_9763,N_9073,N_9350);
or U9764 (N_9764,N_9126,N_9145);
xor U9765 (N_9765,N_9148,N_9249);
and U9766 (N_9766,N_9020,N_9260);
xnor U9767 (N_9767,N_9307,N_9157);
or U9768 (N_9768,N_9243,N_9038);
xnor U9769 (N_9769,N_9003,N_9445);
nor U9770 (N_9770,N_9208,N_9231);
xor U9771 (N_9771,N_9359,N_9355);
nand U9772 (N_9772,N_9202,N_9169);
xnor U9773 (N_9773,N_9313,N_9072);
or U9774 (N_9774,N_9041,N_9075);
xor U9775 (N_9775,N_9306,N_9133);
nand U9776 (N_9776,N_9167,N_9297);
nand U9777 (N_9777,N_9133,N_9348);
and U9778 (N_9778,N_9025,N_9135);
nand U9779 (N_9779,N_9394,N_9418);
xor U9780 (N_9780,N_9324,N_9401);
or U9781 (N_9781,N_9306,N_9288);
nor U9782 (N_9782,N_9474,N_9477);
nand U9783 (N_9783,N_9270,N_9330);
xnor U9784 (N_9784,N_9082,N_9200);
and U9785 (N_9785,N_9383,N_9427);
nand U9786 (N_9786,N_9184,N_9010);
xnor U9787 (N_9787,N_9025,N_9174);
xor U9788 (N_9788,N_9339,N_9100);
nand U9789 (N_9789,N_9168,N_9356);
and U9790 (N_9790,N_9055,N_9016);
nand U9791 (N_9791,N_9207,N_9263);
xnor U9792 (N_9792,N_9390,N_9034);
nand U9793 (N_9793,N_9204,N_9187);
nand U9794 (N_9794,N_9169,N_9082);
and U9795 (N_9795,N_9342,N_9476);
and U9796 (N_9796,N_9311,N_9166);
xnor U9797 (N_9797,N_9487,N_9391);
and U9798 (N_9798,N_9485,N_9059);
nand U9799 (N_9799,N_9449,N_9259);
or U9800 (N_9800,N_9308,N_9270);
and U9801 (N_9801,N_9311,N_9401);
nor U9802 (N_9802,N_9221,N_9334);
and U9803 (N_9803,N_9377,N_9491);
nor U9804 (N_9804,N_9122,N_9432);
nand U9805 (N_9805,N_9154,N_9259);
nand U9806 (N_9806,N_9209,N_9405);
xnor U9807 (N_9807,N_9492,N_9254);
and U9808 (N_9808,N_9487,N_9483);
or U9809 (N_9809,N_9444,N_9299);
xnor U9810 (N_9810,N_9428,N_9202);
and U9811 (N_9811,N_9285,N_9186);
xnor U9812 (N_9812,N_9261,N_9161);
and U9813 (N_9813,N_9054,N_9183);
or U9814 (N_9814,N_9000,N_9479);
or U9815 (N_9815,N_9192,N_9376);
or U9816 (N_9816,N_9177,N_9198);
nand U9817 (N_9817,N_9154,N_9036);
nand U9818 (N_9818,N_9080,N_9346);
nand U9819 (N_9819,N_9105,N_9423);
and U9820 (N_9820,N_9445,N_9140);
xor U9821 (N_9821,N_9058,N_9382);
xnor U9822 (N_9822,N_9085,N_9394);
xor U9823 (N_9823,N_9307,N_9441);
nand U9824 (N_9824,N_9060,N_9243);
nand U9825 (N_9825,N_9274,N_9370);
xnor U9826 (N_9826,N_9294,N_9144);
nor U9827 (N_9827,N_9222,N_9073);
nand U9828 (N_9828,N_9102,N_9227);
nand U9829 (N_9829,N_9419,N_9024);
or U9830 (N_9830,N_9353,N_9260);
nor U9831 (N_9831,N_9492,N_9125);
xor U9832 (N_9832,N_9210,N_9086);
xnor U9833 (N_9833,N_9117,N_9377);
nor U9834 (N_9834,N_9257,N_9287);
xor U9835 (N_9835,N_9004,N_9358);
or U9836 (N_9836,N_9107,N_9097);
and U9837 (N_9837,N_9252,N_9277);
nor U9838 (N_9838,N_9272,N_9025);
nor U9839 (N_9839,N_9104,N_9268);
or U9840 (N_9840,N_9210,N_9212);
nand U9841 (N_9841,N_9122,N_9236);
and U9842 (N_9842,N_9343,N_9259);
and U9843 (N_9843,N_9304,N_9119);
nor U9844 (N_9844,N_9192,N_9143);
xor U9845 (N_9845,N_9249,N_9270);
xnor U9846 (N_9846,N_9152,N_9368);
xor U9847 (N_9847,N_9214,N_9226);
and U9848 (N_9848,N_9211,N_9256);
nand U9849 (N_9849,N_9106,N_9172);
nand U9850 (N_9850,N_9405,N_9486);
nand U9851 (N_9851,N_9145,N_9172);
nand U9852 (N_9852,N_9221,N_9390);
or U9853 (N_9853,N_9192,N_9145);
xnor U9854 (N_9854,N_9380,N_9414);
and U9855 (N_9855,N_9055,N_9128);
xor U9856 (N_9856,N_9046,N_9312);
nand U9857 (N_9857,N_9018,N_9150);
or U9858 (N_9858,N_9065,N_9021);
nand U9859 (N_9859,N_9451,N_9125);
nand U9860 (N_9860,N_9499,N_9481);
nand U9861 (N_9861,N_9366,N_9494);
and U9862 (N_9862,N_9457,N_9341);
or U9863 (N_9863,N_9195,N_9184);
nand U9864 (N_9864,N_9069,N_9431);
and U9865 (N_9865,N_9442,N_9195);
nand U9866 (N_9866,N_9197,N_9179);
nand U9867 (N_9867,N_9115,N_9267);
and U9868 (N_9868,N_9278,N_9350);
or U9869 (N_9869,N_9429,N_9241);
xnor U9870 (N_9870,N_9002,N_9360);
and U9871 (N_9871,N_9334,N_9336);
nor U9872 (N_9872,N_9296,N_9048);
xnor U9873 (N_9873,N_9447,N_9167);
and U9874 (N_9874,N_9089,N_9004);
or U9875 (N_9875,N_9316,N_9123);
xor U9876 (N_9876,N_9050,N_9036);
and U9877 (N_9877,N_9189,N_9118);
or U9878 (N_9878,N_9178,N_9224);
or U9879 (N_9879,N_9190,N_9397);
nor U9880 (N_9880,N_9107,N_9292);
or U9881 (N_9881,N_9123,N_9161);
and U9882 (N_9882,N_9109,N_9192);
xnor U9883 (N_9883,N_9024,N_9363);
xor U9884 (N_9884,N_9254,N_9240);
xor U9885 (N_9885,N_9332,N_9359);
xnor U9886 (N_9886,N_9264,N_9343);
and U9887 (N_9887,N_9078,N_9326);
nand U9888 (N_9888,N_9136,N_9148);
and U9889 (N_9889,N_9050,N_9056);
nor U9890 (N_9890,N_9005,N_9355);
and U9891 (N_9891,N_9254,N_9479);
xor U9892 (N_9892,N_9327,N_9402);
and U9893 (N_9893,N_9293,N_9030);
or U9894 (N_9894,N_9368,N_9403);
or U9895 (N_9895,N_9076,N_9436);
or U9896 (N_9896,N_9342,N_9013);
or U9897 (N_9897,N_9164,N_9239);
nand U9898 (N_9898,N_9250,N_9270);
and U9899 (N_9899,N_9438,N_9125);
or U9900 (N_9900,N_9150,N_9428);
xor U9901 (N_9901,N_9312,N_9193);
nor U9902 (N_9902,N_9353,N_9430);
xnor U9903 (N_9903,N_9249,N_9087);
or U9904 (N_9904,N_9132,N_9307);
or U9905 (N_9905,N_9271,N_9150);
nor U9906 (N_9906,N_9090,N_9042);
nor U9907 (N_9907,N_9456,N_9416);
and U9908 (N_9908,N_9433,N_9390);
xor U9909 (N_9909,N_9021,N_9484);
nand U9910 (N_9910,N_9435,N_9298);
nand U9911 (N_9911,N_9459,N_9181);
nor U9912 (N_9912,N_9088,N_9249);
and U9913 (N_9913,N_9421,N_9308);
and U9914 (N_9914,N_9160,N_9333);
or U9915 (N_9915,N_9264,N_9160);
xnor U9916 (N_9916,N_9427,N_9335);
nand U9917 (N_9917,N_9307,N_9139);
nand U9918 (N_9918,N_9379,N_9371);
or U9919 (N_9919,N_9442,N_9345);
xor U9920 (N_9920,N_9438,N_9264);
or U9921 (N_9921,N_9451,N_9431);
and U9922 (N_9922,N_9351,N_9364);
and U9923 (N_9923,N_9157,N_9356);
and U9924 (N_9924,N_9300,N_9170);
or U9925 (N_9925,N_9132,N_9184);
nand U9926 (N_9926,N_9434,N_9372);
nand U9927 (N_9927,N_9442,N_9141);
or U9928 (N_9928,N_9010,N_9488);
or U9929 (N_9929,N_9170,N_9274);
nand U9930 (N_9930,N_9106,N_9280);
nand U9931 (N_9931,N_9266,N_9352);
nand U9932 (N_9932,N_9290,N_9087);
nand U9933 (N_9933,N_9329,N_9150);
nand U9934 (N_9934,N_9011,N_9131);
xor U9935 (N_9935,N_9418,N_9270);
nor U9936 (N_9936,N_9107,N_9460);
and U9937 (N_9937,N_9279,N_9190);
xnor U9938 (N_9938,N_9212,N_9262);
or U9939 (N_9939,N_9372,N_9477);
or U9940 (N_9940,N_9158,N_9064);
or U9941 (N_9941,N_9259,N_9421);
nand U9942 (N_9942,N_9440,N_9180);
or U9943 (N_9943,N_9404,N_9496);
and U9944 (N_9944,N_9463,N_9022);
nor U9945 (N_9945,N_9396,N_9304);
xnor U9946 (N_9946,N_9019,N_9039);
nand U9947 (N_9947,N_9060,N_9372);
nor U9948 (N_9948,N_9451,N_9068);
or U9949 (N_9949,N_9276,N_9024);
nor U9950 (N_9950,N_9037,N_9293);
nor U9951 (N_9951,N_9188,N_9176);
xor U9952 (N_9952,N_9439,N_9096);
and U9953 (N_9953,N_9215,N_9353);
nor U9954 (N_9954,N_9072,N_9114);
nor U9955 (N_9955,N_9434,N_9253);
and U9956 (N_9956,N_9217,N_9193);
nand U9957 (N_9957,N_9154,N_9427);
or U9958 (N_9958,N_9158,N_9182);
or U9959 (N_9959,N_9423,N_9097);
and U9960 (N_9960,N_9394,N_9313);
nand U9961 (N_9961,N_9452,N_9027);
nand U9962 (N_9962,N_9287,N_9364);
nand U9963 (N_9963,N_9036,N_9337);
xnor U9964 (N_9964,N_9090,N_9296);
xor U9965 (N_9965,N_9215,N_9076);
and U9966 (N_9966,N_9172,N_9156);
or U9967 (N_9967,N_9400,N_9185);
and U9968 (N_9968,N_9479,N_9225);
or U9969 (N_9969,N_9320,N_9392);
nand U9970 (N_9970,N_9107,N_9259);
and U9971 (N_9971,N_9194,N_9459);
or U9972 (N_9972,N_9114,N_9432);
nor U9973 (N_9973,N_9324,N_9476);
or U9974 (N_9974,N_9012,N_9441);
or U9975 (N_9975,N_9005,N_9437);
and U9976 (N_9976,N_9456,N_9391);
nand U9977 (N_9977,N_9071,N_9374);
xnor U9978 (N_9978,N_9329,N_9469);
xor U9979 (N_9979,N_9004,N_9290);
or U9980 (N_9980,N_9420,N_9100);
nand U9981 (N_9981,N_9249,N_9081);
and U9982 (N_9982,N_9360,N_9495);
xnor U9983 (N_9983,N_9351,N_9166);
nor U9984 (N_9984,N_9164,N_9025);
xnor U9985 (N_9985,N_9183,N_9298);
nand U9986 (N_9986,N_9428,N_9296);
and U9987 (N_9987,N_9451,N_9134);
and U9988 (N_9988,N_9440,N_9254);
or U9989 (N_9989,N_9119,N_9341);
xor U9990 (N_9990,N_9046,N_9018);
nor U9991 (N_9991,N_9286,N_9400);
or U9992 (N_9992,N_9237,N_9426);
nor U9993 (N_9993,N_9237,N_9301);
and U9994 (N_9994,N_9468,N_9355);
and U9995 (N_9995,N_9297,N_9017);
xor U9996 (N_9996,N_9334,N_9049);
and U9997 (N_9997,N_9469,N_9252);
nand U9998 (N_9998,N_9208,N_9487);
nand U9999 (N_9999,N_9477,N_9035);
or UO_0 (O_0,N_9662,N_9808);
nor UO_1 (O_1,N_9693,N_9544);
nand UO_2 (O_2,N_9568,N_9522);
and UO_3 (O_3,N_9881,N_9961);
nand UO_4 (O_4,N_9997,N_9756);
and UO_5 (O_5,N_9525,N_9669);
or UO_6 (O_6,N_9869,N_9891);
nor UO_7 (O_7,N_9962,N_9939);
nand UO_8 (O_8,N_9797,N_9701);
nand UO_9 (O_9,N_9699,N_9689);
nand UO_10 (O_10,N_9624,N_9806);
or UO_11 (O_11,N_9635,N_9603);
nand UO_12 (O_12,N_9617,N_9802);
xnor UO_13 (O_13,N_9898,N_9695);
nand UO_14 (O_14,N_9683,N_9653);
or UO_15 (O_15,N_9886,N_9675);
nor UO_16 (O_16,N_9668,N_9838);
nand UO_17 (O_17,N_9971,N_9965);
nor UO_18 (O_18,N_9992,N_9505);
nor UO_19 (O_19,N_9696,N_9561);
nand UO_20 (O_20,N_9684,N_9519);
xnor UO_21 (O_21,N_9863,N_9972);
nor UO_22 (O_22,N_9845,N_9550);
or UO_23 (O_23,N_9560,N_9587);
xor UO_24 (O_24,N_9892,N_9822);
xnor UO_25 (O_25,N_9600,N_9993);
xor UO_26 (O_26,N_9620,N_9973);
nor UO_27 (O_27,N_9630,N_9809);
nor UO_28 (O_28,N_9778,N_9958);
nor UO_29 (O_29,N_9588,N_9592);
or UO_30 (O_30,N_9690,N_9807);
and UO_31 (O_31,N_9826,N_9991);
nand UO_32 (O_32,N_9887,N_9558);
or UO_33 (O_33,N_9697,N_9836);
or UO_34 (O_34,N_9864,N_9786);
and UO_35 (O_35,N_9934,N_9880);
or UO_36 (O_36,N_9792,N_9817);
xor UO_37 (O_37,N_9628,N_9677);
nand UO_38 (O_38,N_9619,N_9625);
and UO_39 (O_39,N_9716,N_9754);
nand UO_40 (O_40,N_9974,N_9828);
or UO_41 (O_41,N_9983,N_9614);
xnor UO_42 (O_42,N_9770,N_9937);
nand UO_43 (O_43,N_9657,N_9702);
or UO_44 (O_44,N_9924,N_9918);
or UO_45 (O_45,N_9979,N_9986);
nor UO_46 (O_46,N_9963,N_9503);
and UO_47 (O_47,N_9647,N_9542);
and UO_48 (O_48,N_9582,N_9783);
or UO_49 (O_49,N_9777,N_9506);
nand UO_50 (O_50,N_9938,N_9764);
nor UO_51 (O_51,N_9688,N_9815);
nor UO_52 (O_52,N_9933,N_9910);
or UO_53 (O_53,N_9913,N_9785);
nor UO_54 (O_54,N_9947,N_9780);
or UO_55 (O_55,N_9650,N_9908);
and UO_56 (O_56,N_9906,N_9810);
nand UO_57 (O_57,N_9956,N_9750);
and UO_58 (O_58,N_9897,N_9573);
nand UO_59 (O_59,N_9800,N_9858);
or UO_60 (O_60,N_9884,N_9530);
nand UO_61 (O_61,N_9847,N_9644);
nand UO_62 (O_62,N_9501,N_9841);
nand UO_63 (O_63,N_9586,N_9514);
nand UO_64 (O_64,N_9804,N_9513);
and UO_65 (O_65,N_9745,N_9618);
xnor UO_66 (O_66,N_9541,N_9734);
and UO_67 (O_67,N_9584,N_9609);
nand UO_68 (O_68,N_9873,N_9927);
nor UO_69 (O_69,N_9563,N_9896);
and UO_70 (O_70,N_9596,N_9645);
and UO_71 (O_71,N_9727,N_9984);
xor UO_72 (O_72,N_9949,N_9502);
nor UO_73 (O_73,N_9524,N_9545);
nand UO_74 (O_74,N_9566,N_9957);
xor UO_75 (O_75,N_9945,N_9649);
or UO_76 (O_76,N_9694,N_9827);
and UO_77 (O_77,N_9564,N_9955);
nor UO_78 (O_78,N_9580,N_9682);
nor UO_79 (O_79,N_9776,N_9981);
xnor UO_80 (O_80,N_9814,N_9616);
nor UO_81 (O_81,N_9639,N_9528);
and UO_82 (O_82,N_9929,N_9857);
and UO_83 (O_83,N_9749,N_9865);
and UO_84 (O_84,N_9554,N_9595);
nand UO_85 (O_85,N_9866,N_9549);
or UO_86 (O_86,N_9871,N_9585);
nor UO_87 (O_87,N_9902,N_9591);
or UO_88 (O_88,N_9994,N_9915);
nor UO_89 (O_89,N_9711,N_9976);
or UO_90 (O_90,N_9904,N_9612);
nand UO_91 (O_91,N_9793,N_9951);
xor UO_92 (O_92,N_9607,N_9515);
xor UO_93 (O_93,N_9931,N_9567);
and UO_94 (O_94,N_9579,N_9943);
xnor UO_95 (O_95,N_9537,N_9517);
nor UO_96 (O_96,N_9520,N_9527);
or UO_97 (O_97,N_9922,N_9834);
xnor UO_98 (O_98,N_9593,N_9534);
nor UO_99 (O_99,N_9705,N_9936);
xnor UO_100 (O_100,N_9874,N_9623);
and UO_101 (O_101,N_9876,N_9559);
or UO_102 (O_102,N_9852,N_9708);
xor UO_103 (O_103,N_9736,N_9533);
xor UO_104 (O_104,N_9948,N_9562);
nor UO_105 (O_105,N_9820,N_9899);
nand UO_106 (O_106,N_9538,N_9673);
xnor UO_107 (O_107,N_9854,N_9781);
nand UO_108 (O_108,N_9724,N_9601);
xor UO_109 (O_109,N_9940,N_9547);
xnor UO_110 (O_110,N_9998,N_9622);
nor UO_111 (O_111,N_9977,N_9535);
nand UO_112 (O_112,N_9510,N_9583);
xnor UO_113 (O_113,N_9661,N_9813);
nand UO_114 (O_114,N_9967,N_9680);
xor UO_115 (O_115,N_9659,N_9811);
xor UO_116 (O_116,N_9737,N_9784);
nand UO_117 (O_117,N_9721,N_9531);
or UO_118 (O_118,N_9782,N_9698);
or UO_119 (O_119,N_9674,N_9553);
nand UO_120 (O_120,N_9610,N_9964);
xor UO_121 (O_121,N_9646,N_9921);
xor UO_122 (O_122,N_9599,N_9678);
xor UO_123 (O_123,N_9691,N_9739);
nor UO_124 (O_124,N_9942,N_9521);
and UO_125 (O_125,N_9726,N_9928);
and UO_126 (O_126,N_9594,N_9759);
nand UO_127 (O_127,N_9632,N_9995);
and UO_128 (O_128,N_9769,N_9779);
nor UO_129 (O_129,N_9751,N_9821);
or UO_130 (O_130,N_9926,N_9511);
nand UO_131 (O_131,N_9685,N_9615);
and UO_132 (O_132,N_9757,N_9867);
nand UO_133 (O_133,N_9523,N_9743);
or UO_134 (O_134,N_9752,N_9642);
and UO_135 (O_135,N_9818,N_9885);
nand UO_136 (O_136,N_9732,N_9990);
nand UO_137 (O_137,N_9829,N_9765);
nand UO_138 (O_138,N_9707,N_9848);
and UO_139 (O_139,N_9969,N_9803);
nand UO_140 (O_140,N_9575,N_9551);
or UO_141 (O_141,N_9570,N_9709);
nor UO_142 (O_142,N_9966,N_9733);
xor UO_143 (O_143,N_9722,N_9576);
xor UO_144 (O_144,N_9687,N_9730);
and UO_145 (O_145,N_9577,N_9629);
nand UO_146 (O_146,N_9552,N_9900);
nand UO_147 (O_147,N_9846,N_9982);
or UO_148 (O_148,N_9844,N_9571);
nand UO_149 (O_149,N_9791,N_9970);
or UO_150 (O_150,N_9795,N_9894);
nand UO_151 (O_151,N_9651,N_9911);
nand UO_152 (O_152,N_9602,N_9843);
and UO_153 (O_153,N_9643,N_9508);
nand UO_154 (O_154,N_9888,N_9636);
nand UO_155 (O_155,N_9773,N_9768);
nor UO_156 (O_156,N_9882,N_9837);
xor UO_157 (O_157,N_9988,N_9613);
and UO_158 (O_158,N_9710,N_9812);
nor UO_159 (O_159,N_9671,N_9794);
nand UO_160 (O_160,N_9598,N_9631);
or UO_161 (O_161,N_9923,N_9941);
nor UO_162 (O_162,N_9723,N_9655);
nor UO_163 (O_163,N_9855,N_9539);
nand UO_164 (O_164,N_9789,N_9504);
xor UO_165 (O_165,N_9893,N_9507);
nor UO_166 (O_166,N_9578,N_9608);
xnor UO_167 (O_167,N_9805,N_9851);
and UO_168 (O_168,N_9704,N_9590);
or UO_169 (O_169,N_9832,N_9572);
xnor UO_170 (O_170,N_9824,N_9890);
and UO_171 (O_171,N_9960,N_9676);
or UO_172 (O_172,N_9907,N_9516);
nand UO_173 (O_173,N_9868,N_9889);
nand UO_174 (O_174,N_9664,N_9987);
or UO_175 (O_175,N_9959,N_9703);
nor UO_176 (O_176,N_9731,N_9798);
nand UO_177 (O_177,N_9917,N_9672);
xor UO_178 (O_178,N_9569,N_9746);
xor UO_179 (O_179,N_9509,N_9718);
xnor UO_180 (O_180,N_9903,N_9747);
or UO_181 (O_181,N_9543,N_9762);
and UO_182 (O_182,N_9540,N_9771);
or UO_183 (O_183,N_9728,N_9909);
nor UO_184 (O_184,N_9856,N_9555);
and UO_185 (O_185,N_9996,N_9638);
and UO_186 (O_186,N_9605,N_9760);
nor UO_187 (O_187,N_9611,N_9686);
and UO_188 (O_188,N_9715,N_9912);
or UO_189 (O_189,N_9742,N_9666);
nor UO_190 (O_190,N_9581,N_9692);
nor UO_191 (O_191,N_9859,N_9796);
or UO_192 (O_192,N_9714,N_9860);
nor UO_193 (O_193,N_9774,N_9916);
or UO_194 (O_194,N_9725,N_9665);
or UO_195 (O_195,N_9556,N_9741);
and UO_196 (O_196,N_9788,N_9872);
and UO_197 (O_197,N_9761,N_9557);
and UO_198 (O_198,N_9627,N_9870);
and UO_199 (O_199,N_9713,N_9920);
nand UO_200 (O_200,N_9823,N_9850);
xnor UO_201 (O_201,N_9700,N_9952);
or UO_202 (O_202,N_9621,N_9740);
nor UO_203 (O_203,N_9606,N_9925);
xor UO_204 (O_204,N_9801,N_9830);
nor UO_205 (O_205,N_9633,N_9660);
nand UO_206 (O_206,N_9574,N_9980);
and UO_207 (O_207,N_9862,N_9637);
nor UO_208 (O_208,N_9597,N_9835);
or UO_209 (O_209,N_9681,N_9999);
nand UO_210 (O_210,N_9719,N_9512);
nand UO_211 (O_211,N_9840,N_9626);
nor UO_212 (O_212,N_9720,N_9914);
or UO_213 (O_213,N_9877,N_9875);
and UO_214 (O_214,N_9663,N_9878);
or UO_215 (O_215,N_9775,N_9744);
and UO_216 (O_216,N_9758,N_9946);
nand UO_217 (O_217,N_9831,N_9654);
nand UO_218 (O_218,N_9589,N_9978);
xor UO_219 (O_219,N_9565,N_9895);
xnor UO_220 (O_220,N_9930,N_9932);
nor UO_221 (O_221,N_9748,N_9518);
nand UO_222 (O_222,N_9819,N_9825);
xnor UO_223 (O_223,N_9546,N_9679);
xnor UO_224 (O_224,N_9905,N_9548);
and UO_225 (O_225,N_9879,N_9766);
or UO_226 (O_226,N_9944,N_9640);
xor UO_227 (O_227,N_9529,N_9833);
nor UO_228 (O_228,N_9968,N_9729);
or UO_229 (O_229,N_9634,N_9706);
or UO_230 (O_230,N_9536,N_9861);
and UO_231 (O_231,N_9772,N_9950);
xor UO_232 (O_232,N_9763,N_9738);
or UO_233 (O_233,N_9755,N_9604);
or UO_234 (O_234,N_9849,N_9712);
nor UO_235 (O_235,N_9839,N_9919);
or UO_236 (O_236,N_9790,N_9500);
nor UO_237 (O_237,N_9799,N_9842);
xor UO_238 (O_238,N_9985,N_9717);
and UO_239 (O_239,N_9853,N_9670);
nand UO_240 (O_240,N_9526,N_9641);
and UO_241 (O_241,N_9953,N_9652);
and UO_242 (O_242,N_9767,N_9883);
and UO_243 (O_243,N_9667,N_9735);
xor UO_244 (O_244,N_9658,N_9954);
and UO_245 (O_245,N_9648,N_9816);
xnor UO_246 (O_246,N_9753,N_9532);
nand UO_247 (O_247,N_9901,N_9989);
or UO_248 (O_248,N_9656,N_9935);
xor UO_249 (O_249,N_9975,N_9787);
nand UO_250 (O_250,N_9978,N_9581);
and UO_251 (O_251,N_9679,N_9686);
xnor UO_252 (O_252,N_9742,N_9570);
xnor UO_253 (O_253,N_9740,N_9960);
xnor UO_254 (O_254,N_9647,N_9521);
and UO_255 (O_255,N_9874,N_9964);
nand UO_256 (O_256,N_9876,N_9875);
or UO_257 (O_257,N_9503,N_9648);
and UO_258 (O_258,N_9818,N_9879);
and UO_259 (O_259,N_9593,N_9580);
and UO_260 (O_260,N_9695,N_9920);
xnor UO_261 (O_261,N_9723,N_9934);
xnor UO_262 (O_262,N_9730,N_9803);
nand UO_263 (O_263,N_9977,N_9534);
xor UO_264 (O_264,N_9506,N_9668);
nor UO_265 (O_265,N_9799,N_9742);
and UO_266 (O_266,N_9867,N_9892);
nand UO_267 (O_267,N_9534,N_9786);
or UO_268 (O_268,N_9788,N_9596);
nand UO_269 (O_269,N_9864,N_9665);
or UO_270 (O_270,N_9996,N_9728);
or UO_271 (O_271,N_9806,N_9686);
nand UO_272 (O_272,N_9833,N_9779);
and UO_273 (O_273,N_9798,N_9686);
and UO_274 (O_274,N_9974,N_9742);
or UO_275 (O_275,N_9719,N_9773);
nand UO_276 (O_276,N_9676,N_9832);
nand UO_277 (O_277,N_9847,N_9842);
or UO_278 (O_278,N_9695,N_9796);
nor UO_279 (O_279,N_9543,N_9877);
xnor UO_280 (O_280,N_9948,N_9702);
or UO_281 (O_281,N_9789,N_9637);
and UO_282 (O_282,N_9824,N_9569);
nor UO_283 (O_283,N_9578,N_9567);
and UO_284 (O_284,N_9655,N_9553);
nor UO_285 (O_285,N_9878,N_9918);
nor UO_286 (O_286,N_9964,N_9976);
nor UO_287 (O_287,N_9545,N_9811);
nor UO_288 (O_288,N_9512,N_9662);
xor UO_289 (O_289,N_9927,N_9501);
nor UO_290 (O_290,N_9916,N_9627);
and UO_291 (O_291,N_9530,N_9778);
and UO_292 (O_292,N_9929,N_9738);
nand UO_293 (O_293,N_9885,N_9989);
or UO_294 (O_294,N_9631,N_9547);
or UO_295 (O_295,N_9510,N_9978);
and UO_296 (O_296,N_9608,N_9670);
and UO_297 (O_297,N_9618,N_9548);
xnor UO_298 (O_298,N_9961,N_9678);
and UO_299 (O_299,N_9542,N_9944);
and UO_300 (O_300,N_9971,N_9888);
nand UO_301 (O_301,N_9991,N_9937);
or UO_302 (O_302,N_9747,N_9982);
and UO_303 (O_303,N_9975,N_9671);
nor UO_304 (O_304,N_9833,N_9719);
xnor UO_305 (O_305,N_9611,N_9637);
and UO_306 (O_306,N_9715,N_9691);
xor UO_307 (O_307,N_9965,N_9623);
nor UO_308 (O_308,N_9540,N_9580);
nand UO_309 (O_309,N_9742,N_9783);
xor UO_310 (O_310,N_9626,N_9726);
nor UO_311 (O_311,N_9710,N_9732);
and UO_312 (O_312,N_9844,N_9724);
or UO_313 (O_313,N_9874,N_9911);
nor UO_314 (O_314,N_9871,N_9782);
nand UO_315 (O_315,N_9570,N_9952);
or UO_316 (O_316,N_9892,N_9816);
xnor UO_317 (O_317,N_9998,N_9748);
xor UO_318 (O_318,N_9896,N_9972);
nor UO_319 (O_319,N_9781,N_9657);
nand UO_320 (O_320,N_9969,N_9698);
nand UO_321 (O_321,N_9794,N_9955);
nand UO_322 (O_322,N_9805,N_9853);
or UO_323 (O_323,N_9601,N_9686);
nand UO_324 (O_324,N_9611,N_9840);
xor UO_325 (O_325,N_9595,N_9830);
or UO_326 (O_326,N_9797,N_9970);
nand UO_327 (O_327,N_9605,N_9726);
nor UO_328 (O_328,N_9921,N_9658);
xnor UO_329 (O_329,N_9897,N_9995);
nand UO_330 (O_330,N_9536,N_9693);
nand UO_331 (O_331,N_9555,N_9862);
nand UO_332 (O_332,N_9527,N_9712);
nor UO_333 (O_333,N_9937,N_9561);
and UO_334 (O_334,N_9917,N_9622);
xor UO_335 (O_335,N_9649,N_9741);
or UO_336 (O_336,N_9724,N_9919);
xor UO_337 (O_337,N_9934,N_9758);
nor UO_338 (O_338,N_9615,N_9534);
or UO_339 (O_339,N_9871,N_9643);
nor UO_340 (O_340,N_9506,N_9609);
nor UO_341 (O_341,N_9925,N_9801);
xor UO_342 (O_342,N_9909,N_9619);
nand UO_343 (O_343,N_9521,N_9858);
xor UO_344 (O_344,N_9648,N_9632);
nand UO_345 (O_345,N_9606,N_9538);
nor UO_346 (O_346,N_9600,N_9717);
nand UO_347 (O_347,N_9796,N_9615);
nor UO_348 (O_348,N_9894,N_9815);
nand UO_349 (O_349,N_9836,N_9915);
nor UO_350 (O_350,N_9909,N_9609);
or UO_351 (O_351,N_9809,N_9597);
nand UO_352 (O_352,N_9609,N_9634);
or UO_353 (O_353,N_9635,N_9924);
or UO_354 (O_354,N_9519,N_9541);
and UO_355 (O_355,N_9681,N_9567);
nor UO_356 (O_356,N_9551,N_9946);
xnor UO_357 (O_357,N_9866,N_9697);
nor UO_358 (O_358,N_9653,N_9774);
xor UO_359 (O_359,N_9733,N_9697);
and UO_360 (O_360,N_9949,N_9588);
nand UO_361 (O_361,N_9546,N_9520);
nand UO_362 (O_362,N_9705,N_9760);
nor UO_363 (O_363,N_9893,N_9632);
or UO_364 (O_364,N_9711,N_9864);
xor UO_365 (O_365,N_9922,N_9820);
or UO_366 (O_366,N_9791,N_9767);
nor UO_367 (O_367,N_9930,N_9723);
xnor UO_368 (O_368,N_9542,N_9604);
and UO_369 (O_369,N_9997,N_9785);
or UO_370 (O_370,N_9669,N_9724);
nand UO_371 (O_371,N_9934,N_9515);
or UO_372 (O_372,N_9871,N_9862);
and UO_373 (O_373,N_9816,N_9713);
xnor UO_374 (O_374,N_9809,N_9774);
and UO_375 (O_375,N_9739,N_9867);
xor UO_376 (O_376,N_9919,N_9991);
nor UO_377 (O_377,N_9775,N_9548);
and UO_378 (O_378,N_9984,N_9735);
or UO_379 (O_379,N_9939,N_9920);
and UO_380 (O_380,N_9541,N_9652);
or UO_381 (O_381,N_9891,N_9867);
xor UO_382 (O_382,N_9503,N_9783);
nor UO_383 (O_383,N_9960,N_9695);
and UO_384 (O_384,N_9893,N_9839);
xor UO_385 (O_385,N_9676,N_9576);
and UO_386 (O_386,N_9899,N_9705);
xnor UO_387 (O_387,N_9590,N_9538);
nand UO_388 (O_388,N_9784,N_9954);
and UO_389 (O_389,N_9872,N_9864);
nor UO_390 (O_390,N_9933,N_9973);
and UO_391 (O_391,N_9745,N_9856);
xnor UO_392 (O_392,N_9589,N_9691);
nand UO_393 (O_393,N_9807,N_9540);
nor UO_394 (O_394,N_9767,N_9799);
xnor UO_395 (O_395,N_9882,N_9889);
nor UO_396 (O_396,N_9714,N_9901);
nand UO_397 (O_397,N_9910,N_9801);
or UO_398 (O_398,N_9748,N_9889);
nor UO_399 (O_399,N_9690,N_9716);
and UO_400 (O_400,N_9583,N_9655);
or UO_401 (O_401,N_9723,N_9694);
or UO_402 (O_402,N_9798,N_9891);
nand UO_403 (O_403,N_9913,N_9728);
nor UO_404 (O_404,N_9553,N_9816);
nand UO_405 (O_405,N_9745,N_9572);
and UO_406 (O_406,N_9971,N_9773);
and UO_407 (O_407,N_9799,N_9995);
nor UO_408 (O_408,N_9580,N_9980);
nand UO_409 (O_409,N_9993,N_9591);
and UO_410 (O_410,N_9763,N_9830);
xor UO_411 (O_411,N_9982,N_9945);
nand UO_412 (O_412,N_9900,N_9863);
xor UO_413 (O_413,N_9853,N_9965);
nand UO_414 (O_414,N_9734,N_9986);
nor UO_415 (O_415,N_9877,N_9554);
xor UO_416 (O_416,N_9875,N_9644);
or UO_417 (O_417,N_9687,N_9667);
xnor UO_418 (O_418,N_9881,N_9793);
nand UO_419 (O_419,N_9922,N_9870);
nand UO_420 (O_420,N_9596,N_9821);
nand UO_421 (O_421,N_9530,N_9639);
nor UO_422 (O_422,N_9709,N_9602);
and UO_423 (O_423,N_9661,N_9757);
or UO_424 (O_424,N_9627,N_9853);
nor UO_425 (O_425,N_9731,N_9536);
nor UO_426 (O_426,N_9697,N_9799);
xnor UO_427 (O_427,N_9921,N_9804);
xnor UO_428 (O_428,N_9968,N_9798);
or UO_429 (O_429,N_9870,N_9684);
nand UO_430 (O_430,N_9540,N_9597);
and UO_431 (O_431,N_9723,N_9863);
xor UO_432 (O_432,N_9625,N_9638);
nand UO_433 (O_433,N_9660,N_9598);
nor UO_434 (O_434,N_9801,N_9622);
and UO_435 (O_435,N_9719,N_9920);
or UO_436 (O_436,N_9979,N_9931);
nand UO_437 (O_437,N_9740,N_9622);
and UO_438 (O_438,N_9869,N_9849);
xor UO_439 (O_439,N_9595,N_9633);
and UO_440 (O_440,N_9731,N_9698);
and UO_441 (O_441,N_9902,N_9708);
xor UO_442 (O_442,N_9825,N_9533);
nor UO_443 (O_443,N_9668,N_9917);
nand UO_444 (O_444,N_9861,N_9561);
and UO_445 (O_445,N_9872,N_9687);
nor UO_446 (O_446,N_9506,N_9622);
and UO_447 (O_447,N_9876,N_9913);
xor UO_448 (O_448,N_9646,N_9672);
or UO_449 (O_449,N_9640,N_9869);
and UO_450 (O_450,N_9873,N_9522);
nor UO_451 (O_451,N_9560,N_9512);
xor UO_452 (O_452,N_9747,N_9906);
nand UO_453 (O_453,N_9633,N_9758);
and UO_454 (O_454,N_9838,N_9652);
or UO_455 (O_455,N_9651,N_9628);
nand UO_456 (O_456,N_9876,N_9599);
or UO_457 (O_457,N_9759,N_9581);
xor UO_458 (O_458,N_9679,N_9618);
or UO_459 (O_459,N_9832,N_9936);
nor UO_460 (O_460,N_9621,N_9815);
nor UO_461 (O_461,N_9524,N_9710);
and UO_462 (O_462,N_9543,N_9741);
nand UO_463 (O_463,N_9810,N_9910);
nand UO_464 (O_464,N_9563,N_9880);
or UO_465 (O_465,N_9514,N_9894);
xnor UO_466 (O_466,N_9943,N_9558);
xor UO_467 (O_467,N_9576,N_9601);
and UO_468 (O_468,N_9767,N_9539);
xor UO_469 (O_469,N_9599,N_9583);
nor UO_470 (O_470,N_9890,N_9968);
nand UO_471 (O_471,N_9698,N_9915);
nand UO_472 (O_472,N_9732,N_9897);
and UO_473 (O_473,N_9655,N_9814);
and UO_474 (O_474,N_9646,N_9905);
nor UO_475 (O_475,N_9932,N_9886);
and UO_476 (O_476,N_9874,N_9953);
or UO_477 (O_477,N_9843,N_9787);
nand UO_478 (O_478,N_9728,N_9655);
or UO_479 (O_479,N_9834,N_9914);
or UO_480 (O_480,N_9871,N_9645);
nand UO_481 (O_481,N_9832,N_9893);
nor UO_482 (O_482,N_9639,N_9747);
and UO_483 (O_483,N_9918,N_9895);
and UO_484 (O_484,N_9872,N_9570);
xnor UO_485 (O_485,N_9690,N_9890);
nor UO_486 (O_486,N_9835,N_9547);
nand UO_487 (O_487,N_9680,N_9787);
nand UO_488 (O_488,N_9675,N_9918);
or UO_489 (O_489,N_9843,N_9668);
nand UO_490 (O_490,N_9917,N_9749);
nand UO_491 (O_491,N_9614,N_9626);
or UO_492 (O_492,N_9856,N_9926);
and UO_493 (O_493,N_9880,N_9889);
or UO_494 (O_494,N_9592,N_9694);
xnor UO_495 (O_495,N_9571,N_9612);
nor UO_496 (O_496,N_9636,N_9745);
nor UO_497 (O_497,N_9990,N_9782);
or UO_498 (O_498,N_9594,N_9648);
nor UO_499 (O_499,N_9897,N_9665);
nor UO_500 (O_500,N_9517,N_9561);
or UO_501 (O_501,N_9929,N_9696);
or UO_502 (O_502,N_9772,N_9902);
and UO_503 (O_503,N_9666,N_9522);
xnor UO_504 (O_504,N_9739,N_9925);
nor UO_505 (O_505,N_9716,N_9954);
xor UO_506 (O_506,N_9684,N_9656);
nor UO_507 (O_507,N_9550,N_9940);
or UO_508 (O_508,N_9974,N_9703);
or UO_509 (O_509,N_9743,N_9712);
and UO_510 (O_510,N_9853,N_9847);
nor UO_511 (O_511,N_9587,N_9831);
nand UO_512 (O_512,N_9771,N_9893);
nor UO_513 (O_513,N_9945,N_9628);
xnor UO_514 (O_514,N_9895,N_9732);
nor UO_515 (O_515,N_9587,N_9726);
nand UO_516 (O_516,N_9879,N_9797);
and UO_517 (O_517,N_9580,N_9885);
nand UO_518 (O_518,N_9884,N_9742);
and UO_519 (O_519,N_9735,N_9603);
or UO_520 (O_520,N_9761,N_9652);
xnor UO_521 (O_521,N_9828,N_9543);
and UO_522 (O_522,N_9962,N_9916);
nand UO_523 (O_523,N_9598,N_9828);
nor UO_524 (O_524,N_9637,N_9830);
xor UO_525 (O_525,N_9603,N_9845);
nand UO_526 (O_526,N_9534,N_9839);
nor UO_527 (O_527,N_9757,N_9551);
nor UO_528 (O_528,N_9875,N_9786);
xor UO_529 (O_529,N_9605,N_9563);
xnor UO_530 (O_530,N_9511,N_9565);
xor UO_531 (O_531,N_9614,N_9910);
nor UO_532 (O_532,N_9921,N_9825);
and UO_533 (O_533,N_9755,N_9627);
xor UO_534 (O_534,N_9863,N_9692);
and UO_535 (O_535,N_9685,N_9833);
nor UO_536 (O_536,N_9739,N_9716);
xnor UO_537 (O_537,N_9849,N_9726);
or UO_538 (O_538,N_9588,N_9615);
or UO_539 (O_539,N_9840,N_9868);
nor UO_540 (O_540,N_9675,N_9543);
xnor UO_541 (O_541,N_9586,N_9762);
nor UO_542 (O_542,N_9551,N_9787);
xnor UO_543 (O_543,N_9913,N_9595);
nor UO_544 (O_544,N_9631,N_9868);
xor UO_545 (O_545,N_9653,N_9910);
nor UO_546 (O_546,N_9692,N_9638);
xor UO_547 (O_547,N_9535,N_9773);
or UO_548 (O_548,N_9862,N_9777);
nand UO_549 (O_549,N_9508,N_9575);
nand UO_550 (O_550,N_9899,N_9752);
nor UO_551 (O_551,N_9768,N_9943);
and UO_552 (O_552,N_9695,N_9686);
or UO_553 (O_553,N_9557,N_9571);
and UO_554 (O_554,N_9713,N_9829);
and UO_555 (O_555,N_9636,N_9559);
nor UO_556 (O_556,N_9622,N_9757);
and UO_557 (O_557,N_9829,N_9683);
xor UO_558 (O_558,N_9757,N_9904);
nor UO_559 (O_559,N_9940,N_9564);
nand UO_560 (O_560,N_9618,N_9575);
and UO_561 (O_561,N_9840,N_9939);
xnor UO_562 (O_562,N_9767,N_9741);
xor UO_563 (O_563,N_9568,N_9571);
nand UO_564 (O_564,N_9757,N_9641);
xnor UO_565 (O_565,N_9717,N_9818);
xnor UO_566 (O_566,N_9924,N_9691);
nor UO_567 (O_567,N_9656,N_9816);
xor UO_568 (O_568,N_9768,N_9660);
xor UO_569 (O_569,N_9663,N_9707);
or UO_570 (O_570,N_9556,N_9636);
and UO_571 (O_571,N_9937,N_9501);
and UO_572 (O_572,N_9903,N_9944);
xor UO_573 (O_573,N_9764,N_9838);
and UO_574 (O_574,N_9542,N_9812);
xnor UO_575 (O_575,N_9938,N_9697);
and UO_576 (O_576,N_9708,N_9638);
nand UO_577 (O_577,N_9879,N_9990);
xnor UO_578 (O_578,N_9563,N_9922);
nor UO_579 (O_579,N_9671,N_9521);
xnor UO_580 (O_580,N_9717,N_9719);
or UO_581 (O_581,N_9586,N_9715);
nand UO_582 (O_582,N_9734,N_9531);
nor UO_583 (O_583,N_9908,N_9680);
and UO_584 (O_584,N_9730,N_9760);
and UO_585 (O_585,N_9504,N_9889);
nand UO_586 (O_586,N_9879,N_9596);
nand UO_587 (O_587,N_9863,N_9921);
nor UO_588 (O_588,N_9864,N_9680);
nor UO_589 (O_589,N_9808,N_9898);
and UO_590 (O_590,N_9951,N_9749);
xor UO_591 (O_591,N_9715,N_9732);
nor UO_592 (O_592,N_9924,N_9604);
xnor UO_593 (O_593,N_9891,N_9616);
xor UO_594 (O_594,N_9596,N_9975);
nor UO_595 (O_595,N_9802,N_9578);
xor UO_596 (O_596,N_9611,N_9998);
nor UO_597 (O_597,N_9903,N_9740);
and UO_598 (O_598,N_9847,N_9524);
and UO_599 (O_599,N_9582,N_9607);
xnor UO_600 (O_600,N_9645,N_9721);
nor UO_601 (O_601,N_9766,N_9792);
and UO_602 (O_602,N_9899,N_9877);
nand UO_603 (O_603,N_9603,N_9737);
xnor UO_604 (O_604,N_9519,N_9975);
and UO_605 (O_605,N_9544,N_9817);
nor UO_606 (O_606,N_9541,N_9571);
nor UO_607 (O_607,N_9506,N_9673);
or UO_608 (O_608,N_9790,N_9797);
or UO_609 (O_609,N_9669,N_9790);
xnor UO_610 (O_610,N_9932,N_9865);
or UO_611 (O_611,N_9881,N_9864);
nor UO_612 (O_612,N_9682,N_9997);
xnor UO_613 (O_613,N_9577,N_9500);
nand UO_614 (O_614,N_9722,N_9653);
and UO_615 (O_615,N_9644,N_9673);
nor UO_616 (O_616,N_9544,N_9745);
or UO_617 (O_617,N_9911,N_9902);
nor UO_618 (O_618,N_9920,N_9675);
nand UO_619 (O_619,N_9879,N_9842);
xor UO_620 (O_620,N_9913,N_9842);
nor UO_621 (O_621,N_9511,N_9676);
or UO_622 (O_622,N_9762,N_9748);
or UO_623 (O_623,N_9665,N_9786);
nand UO_624 (O_624,N_9861,N_9825);
nor UO_625 (O_625,N_9934,N_9724);
or UO_626 (O_626,N_9694,N_9769);
nor UO_627 (O_627,N_9858,N_9704);
xor UO_628 (O_628,N_9745,N_9726);
or UO_629 (O_629,N_9765,N_9916);
nor UO_630 (O_630,N_9734,N_9996);
nand UO_631 (O_631,N_9522,N_9940);
and UO_632 (O_632,N_9520,N_9793);
nor UO_633 (O_633,N_9735,N_9810);
nand UO_634 (O_634,N_9568,N_9861);
or UO_635 (O_635,N_9835,N_9896);
and UO_636 (O_636,N_9834,N_9667);
nor UO_637 (O_637,N_9899,N_9715);
and UO_638 (O_638,N_9928,N_9820);
nor UO_639 (O_639,N_9686,N_9851);
nor UO_640 (O_640,N_9632,N_9587);
and UO_641 (O_641,N_9623,N_9797);
nor UO_642 (O_642,N_9818,N_9546);
nand UO_643 (O_643,N_9840,N_9907);
nor UO_644 (O_644,N_9763,N_9652);
xor UO_645 (O_645,N_9915,N_9817);
nand UO_646 (O_646,N_9546,N_9901);
and UO_647 (O_647,N_9733,N_9562);
xnor UO_648 (O_648,N_9901,N_9543);
nor UO_649 (O_649,N_9876,N_9965);
nor UO_650 (O_650,N_9983,N_9535);
xor UO_651 (O_651,N_9639,N_9593);
nor UO_652 (O_652,N_9511,N_9551);
nor UO_653 (O_653,N_9796,N_9827);
nor UO_654 (O_654,N_9929,N_9552);
nor UO_655 (O_655,N_9587,N_9510);
xor UO_656 (O_656,N_9607,N_9728);
or UO_657 (O_657,N_9718,N_9875);
nand UO_658 (O_658,N_9936,N_9814);
or UO_659 (O_659,N_9618,N_9917);
xnor UO_660 (O_660,N_9704,N_9986);
nor UO_661 (O_661,N_9721,N_9551);
nor UO_662 (O_662,N_9912,N_9671);
or UO_663 (O_663,N_9656,N_9688);
nand UO_664 (O_664,N_9996,N_9983);
and UO_665 (O_665,N_9791,N_9633);
nor UO_666 (O_666,N_9601,N_9809);
nand UO_667 (O_667,N_9523,N_9695);
and UO_668 (O_668,N_9777,N_9923);
xor UO_669 (O_669,N_9787,N_9797);
or UO_670 (O_670,N_9648,N_9561);
nor UO_671 (O_671,N_9821,N_9996);
nand UO_672 (O_672,N_9846,N_9590);
nor UO_673 (O_673,N_9794,N_9853);
or UO_674 (O_674,N_9532,N_9738);
or UO_675 (O_675,N_9900,N_9505);
nor UO_676 (O_676,N_9872,N_9629);
and UO_677 (O_677,N_9960,N_9629);
and UO_678 (O_678,N_9815,N_9691);
and UO_679 (O_679,N_9805,N_9762);
or UO_680 (O_680,N_9624,N_9883);
or UO_681 (O_681,N_9784,N_9662);
or UO_682 (O_682,N_9892,N_9679);
or UO_683 (O_683,N_9560,N_9945);
xor UO_684 (O_684,N_9578,N_9544);
nand UO_685 (O_685,N_9805,N_9856);
nand UO_686 (O_686,N_9787,N_9946);
or UO_687 (O_687,N_9944,N_9632);
xor UO_688 (O_688,N_9519,N_9676);
or UO_689 (O_689,N_9664,N_9570);
xnor UO_690 (O_690,N_9643,N_9756);
nor UO_691 (O_691,N_9724,N_9718);
or UO_692 (O_692,N_9664,N_9864);
or UO_693 (O_693,N_9854,N_9595);
nor UO_694 (O_694,N_9797,N_9518);
nand UO_695 (O_695,N_9821,N_9702);
or UO_696 (O_696,N_9754,N_9804);
nand UO_697 (O_697,N_9911,N_9848);
nor UO_698 (O_698,N_9989,N_9605);
or UO_699 (O_699,N_9905,N_9981);
or UO_700 (O_700,N_9623,N_9705);
nor UO_701 (O_701,N_9828,N_9841);
and UO_702 (O_702,N_9943,N_9752);
or UO_703 (O_703,N_9792,N_9771);
xor UO_704 (O_704,N_9960,N_9571);
nand UO_705 (O_705,N_9584,N_9702);
and UO_706 (O_706,N_9543,N_9792);
xnor UO_707 (O_707,N_9645,N_9876);
xnor UO_708 (O_708,N_9966,N_9518);
nand UO_709 (O_709,N_9735,N_9569);
or UO_710 (O_710,N_9889,N_9760);
or UO_711 (O_711,N_9697,N_9648);
xnor UO_712 (O_712,N_9874,N_9620);
xor UO_713 (O_713,N_9870,N_9516);
or UO_714 (O_714,N_9914,N_9943);
and UO_715 (O_715,N_9561,N_9834);
xnor UO_716 (O_716,N_9688,N_9810);
nand UO_717 (O_717,N_9802,N_9798);
nor UO_718 (O_718,N_9780,N_9540);
nor UO_719 (O_719,N_9542,N_9871);
and UO_720 (O_720,N_9607,N_9880);
nor UO_721 (O_721,N_9764,N_9921);
or UO_722 (O_722,N_9544,N_9923);
nor UO_723 (O_723,N_9625,N_9910);
nand UO_724 (O_724,N_9834,N_9659);
nor UO_725 (O_725,N_9748,N_9671);
nor UO_726 (O_726,N_9725,N_9502);
nand UO_727 (O_727,N_9698,N_9724);
nor UO_728 (O_728,N_9895,N_9849);
nor UO_729 (O_729,N_9988,N_9751);
nor UO_730 (O_730,N_9709,N_9909);
nand UO_731 (O_731,N_9547,N_9899);
nor UO_732 (O_732,N_9527,N_9853);
or UO_733 (O_733,N_9608,N_9535);
or UO_734 (O_734,N_9783,N_9516);
or UO_735 (O_735,N_9820,N_9772);
xor UO_736 (O_736,N_9533,N_9507);
nand UO_737 (O_737,N_9958,N_9628);
nor UO_738 (O_738,N_9800,N_9993);
nand UO_739 (O_739,N_9599,N_9864);
nor UO_740 (O_740,N_9819,N_9537);
nor UO_741 (O_741,N_9724,N_9608);
xnor UO_742 (O_742,N_9738,N_9771);
xnor UO_743 (O_743,N_9585,N_9734);
and UO_744 (O_744,N_9734,N_9922);
and UO_745 (O_745,N_9976,N_9762);
and UO_746 (O_746,N_9764,N_9541);
and UO_747 (O_747,N_9545,N_9867);
and UO_748 (O_748,N_9653,N_9712);
nor UO_749 (O_749,N_9711,N_9546);
or UO_750 (O_750,N_9693,N_9756);
nand UO_751 (O_751,N_9536,N_9987);
nand UO_752 (O_752,N_9838,N_9733);
xnor UO_753 (O_753,N_9653,N_9666);
or UO_754 (O_754,N_9534,N_9556);
nor UO_755 (O_755,N_9758,N_9768);
nor UO_756 (O_756,N_9976,N_9614);
nor UO_757 (O_757,N_9637,N_9713);
nand UO_758 (O_758,N_9524,N_9866);
nand UO_759 (O_759,N_9988,N_9562);
or UO_760 (O_760,N_9807,N_9763);
and UO_761 (O_761,N_9829,N_9813);
nand UO_762 (O_762,N_9753,N_9584);
xnor UO_763 (O_763,N_9509,N_9677);
nand UO_764 (O_764,N_9847,N_9952);
nand UO_765 (O_765,N_9987,N_9934);
nor UO_766 (O_766,N_9556,N_9693);
and UO_767 (O_767,N_9771,N_9713);
nand UO_768 (O_768,N_9597,N_9750);
xnor UO_769 (O_769,N_9958,N_9521);
nand UO_770 (O_770,N_9871,N_9830);
or UO_771 (O_771,N_9802,N_9720);
nand UO_772 (O_772,N_9882,N_9542);
nand UO_773 (O_773,N_9664,N_9741);
nor UO_774 (O_774,N_9960,N_9900);
nor UO_775 (O_775,N_9969,N_9745);
xor UO_776 (O_776,N_9712,N_9824);
nor UO_777 (O_777,N_9873,N_9989);
xnor UO_778 (O_778,N_9912,N_9914);
nor UO_779 (O_779,N_9794,N_9625);
nor UO_780 (O_780,N_9872,N_9878);
nand UO_781 (O_781,N_9615,N_9916);
nor UO_782 (O_782,N_9639,N_9759);
nand UO_783 (O_783,N_9558,N_9798);
or UO_784 (O_784,N_9709,N_9596);
and UO_785 (O_785,N_9561,N_9877);
nand UO_786 (O_786,N_9953,N_9914);
and UO_787 (O_787,N_9824,N_9814);
nor UO_788 (O_788,N_9998,N_9686);
nand UO_789 (O_789,N_9985,N_9742);
nand UO_790 (O_790,N_9988,N_9945);
xor UO_791 (O_791,N_9935,N_9926);
xnor UO_792 (O_792,N_9744,N_9508);
or UO_793 (O_793,N_9651,N_9930);
or UO_794 (O_794,N_9824,N_9778);
nor UO_795 (O_795,N_9653,N_9900);
and UO_796 (O_796,N_9648,N_9518);
or UO_797 (O_797,N_9603,N_9851);
xor UO_798 (O_798,N_9695,N_9514);
nand UO_799 (O_799,N_9900,N_9606);
nor UO_800 (O_800,N_9580,N_9901);
xnor UO_801 (O_801,N_9769,N_9919);
nand UO_802 (O_802,N_9763,N_9888);
and UO_803 (O_803,N_9913,N_9592);
and UO_804 (O_804,N_9723,N_9574);
and UO_805 (O_805,N_9609,N_9849);
xnor UO_806 (O_806,N_9578,N_9675);
xor UO_807 (O_807,N_9887,N_9952);
nand UO_808 (O_808,N_9729,N_9545);
nor UO_809 (O_809,N_9613,N_9637);
and UO_810 (O_810,N_9549,N_9985);
and UO_811 (O_811,N_9945,N_9984);
nor UO_812 (O_812,N_9911,N_9900);
nor UO_813 (O_813,N_9509,N_9797);
nand UO_814 (O_814,N_9843,N_9775);
and UO_815 (O_815,N_9684,N_9795);
and UO_816 (O_816,N_9677,N_9933);
nand UO_817 (O_817,N_9676,N_9713);
and UO_818 (O_818,N_9736,N_9686);
or UO_819 (O_819,N_9617,N_9533);
and UO_820 (O_820,N_9598,N_9736);
xor UO_821 (O_821,N_9768,N_9759);
and UO_822 (O_822,N_9638,N_9766);
nor UO_823 (O_823,N_9963,N_9820);
xnor UO_824 (O_824,N_9861,N_9834);
xor UO_825 (O_825,N_9871,N_9597);
or UO_826 (O_826,N_9700,N_9954);
nor UO_827 (O_827,N_9925,N_9782);
and UO_828 (O_828,N_9800,N_9986);
nand UO_829 (O_829,N_9540,N_9785);
nor UO_830 (O_830,N_9647,N_9767);
xor UO_831 (O_831,N_9502,N_9540);
nand UO_832 (O_832,N_9800,N_9895);
or UO_833 (O_833,N_9772,N_9623);
or UO_834 (O_834,N_9885,N_9882);
or UO_835 (O_835,N_9937,N_9940);
nand UO_836 (O_836,N_9648,N_9691);
xor UO_837 (O_837,N_9730,N_9947);
and UO_838 (O_838,N_9590,N_9771);
and UO_839 (O_839,N_9560,N_9810);
or UO_840 (O_840,N_9590,N_9949);
and UO_841 (O_841,N_9519,N_9907);
and UO_842 (O_842,N_9747,N_9678);
and UO_843 (O_843,N_9682,N_9897);
or UO_844 (O_844,N_9568,N_9805);
or UO_845 (O_845,N_9660,N_9925);
or UO_846 (O_846,N_9593,N_9799);
and UO_847 (O_847,N_9653,N_9623);
or UO_848 (O_848,N_9797,N_9654);
or UO_849 (O_849,N_9868,N_9556);
or UO_850 (O_850,N_9977,N_9602);
or UO_851 (O_851,N_9952,N_9575);
or UO_852 (O_852,N_9708,N_9526);
nor UO_853 (O_853,N_9892,N_9776);
xnor UO_854 (O_854,N_9754,N_9519);
nand UO_855 (O_855,N_9786,N_9519);
and UO_856 (O_856,N_9657,N_9753);
nor UO_857 (O_857,N_9720,N_9818);
xnor UO_858 (O_858,N_9533,N_9648);
nand UO_859 (O_859,N_9732,N_9979);
nand UO_860 (O_860,N_9512,N_9629);
nand UO_861 (O_861,N_9523,N_9647);
xor UO_862 (O_862,N_9856,N_9648);
nor UO_863 (O_863,N_9724,N_9754);
or UO_864 (O_864,N_9638,N_9773);
and UO_865 (O_865,N_9782,N_9962);
xnor UO_866 (O_866,N_9500,N_9918);
nor UO_867 (O_867,N_9662,N_9910);
or UO_868 (O_868,N_9891,N_9611);
nand UO_869 (O_869,N_9758,N_9842);
nand UO_870 (O_870,N_9577,N_9801);
nand UO_871 (O_871,N_9914,N_9506);
and UO_872 (O_872,N_9823,N_9583);
nand UO_873 (O_873,N_9834,N_9621);
or UO_874 (O_874,N_9661,N_9586);
and UO_875 (O_875,N_9889,N_9580);
or UO_876 (O_876,N_9844,N_9798);
xor UO_877 (O_877,N_9874,N_9956);
xor UO_878 (O_878,N_9658,N_9834);
xor UO_879 (O_879,N_9593,N_9954);
nor UO_880 (O_880,N_9642,N_9578);
nor UO_881 (O_881,N_9753,N_9574);
or UO_882 (O_882,N_9842,N_9858);
and UO_883 (O_883,N_9506,N_9563);
nand UO_884 (O_884,N_9563,N_9520);
or UO_885 (O_885,N_9526,N_9688);
and UO_886 (O_886,N_9577,N_9848);
nand UO_887 (O_887,N_9909,N_9590);
nand UO_888 (O_888,N_9535,N_9670);
and UO_889 (O_889,N_9957,N_9751);
xor UO_890 (O_890,N_9861,N_9898);
and UO_891 (O_891,N_9952,N_9907);
and UO_892 (O_892,N_9782,N_9697);
and UO_893 (O_893,N_9840,N_9943);
nor UO_894 (O_894,N_9932,N_9660);
or UO_895 (O_895,N_9990,N_9696);
or UO_896 (O_896,N_9812,N_9562);
nand UO_897 (O_897,N_9736,N_9776);
nand UO_898 (O_898,N_9719,N_9687);
or UO_899 (O_899,N_9843,N_9625);
nor UO_900 (O_900,N_9854,N_9664);
or UO_901 (O_901,N_9719,N_9674);
and UO_902 (O_902,N_9637,N_9508);
xnor UO_903 (O_903,N_9692,N_9566);
nor UO_904 (O_904,N_9753,N_9954);
xor UO_905 (O_905,N_9592,N_9875);
nand UO_906 (O_906,N_9920,N_9729);
nand UO_907 (O_907,N_9548,N_9567);
or UO_908 (O_908,N_9636,N_9513);
nor UO_909 (O_909,N_9965,N_9767);
and UO_910 (O_910,N_9678,N_9770);
nand UO_911 (O_911,N_9927,N_9882);
and UO_912 (O_912,N_9596,N_9964);
xnor UO_913 (O_913,N_9868,N_9689);
xor UO_914 (O_914,N_9624,N_9605);
nor UO_915 (O_915,N_9935,N_9908);
nor UO_916 (O_916,N_9920,N_9833);
or UO_917 (O_917,N_9850,N_9902);
nand UO_918 (O_918,N_9811,N_9795);
and UO_919 (O_919,N_9673,N_9554);
nor UO_920 (O_920,N_9654,N_9690);
xor UO_921 (O_921,N_9845,N_9982);
xnor UO_922 (O_922,N_9556,N_9751);
nor UO_923 (O_923,N_9973,N_9814);
nor UO_924 (O_924,N_9601,N_9629);
nor UO_925 (O_925,N_9532,N_9836);
nor UO_926 (O_926,N_9929,N_9762);
nand UO_927 (O_927,N_9985,N_9956);
and UO_928 (O_928,N_9992,N_9964);
nand UO_929 (O_929,N_9758,N_9624);
and UO_930 (O_930,N_9721,N_9801);
nor UO_931 (O_931,N_9948,N_9669);
and UO_932 (O_932,N_9900,N_9516);
nand UO_933 (O_933,N_9576,N_9647);
nand UO_934 (O_934,N_9571,N_9774);
xnor UO_935 (O_935,N_9669,N_9888);
nand UO_936 (O_936,N_9533,N_9565);
xnor UO_937 (O_937,N_9689,N_9632);
or UO_938 (O_938,N_9845,N_9822);
xor UO_939 (O_939,N_9778,N_9820);
or UO_940 (O_940,N_9886,N_9774);
and UO_941 (O_941,N_9876,N_9869);
and UO_942 (O_942,N_9843,N_9821);
nor UO_943 (O_943,N_9505,N_9834);
nand UO_944 (O_944,N_9794,N_9640);
or UO_945 (O_945,N_9509,N_9503);
nor UO_946 (O_946,N_9531,N_9999);
nand UO_947 (O_947,N_9534,N_9871);
xor UO_948 (O_948,N_9583,N_9725);
nand UO_949 (O_949,N_9523,N_9913);
xor UO_950 (O_950,N_9851,N_9788);
xor UO_951 (O_951,N_9842,N_9965);
xnor UO_952 (O_952,N_9995,N_9949);
nand UO_953 (O_953,N_9514,N_9700);
and UO_954 (O_954,N_9834,N_9630);
xnor UO_955 (O_955,N_9612,N_9973);
and UO_956 (O_956,N_9501,N_9944);
or UO_957 (O_957,N_9731,N_9621);
and UO_958 (O_958,N_9586,N_9560);
or UO_959 (O_959,N_9627,N_9532);
nor UO_960 (O_960,N_9933,N_9952);
or UO_961 (O_961,N_9647,N_9682);
and UO_962 (O_962,N_9781,N_9938);
xor UO_963 (O_963,N_9973,N_9745);
nor UO_964 (O_964,N_9754,N_9593);
and UO_965 (O_965,N_9566,N_9555);
nand UO_966 (O_966,N_9660,N_9818);
or UO_967 (O_967,N_9539,N_9711);
or UO_968 (O_968,N_9961,N_9988);
xor UO_969 (O_969,N_9708,N_9671);
nor UO_970 (O_970,N_9963,N_9915);
xnor UO_971 (O_971,N_9657,N_9933);
xnor UO_972 (O_972,N_9855,N_9996);
xnor UO_973 (O_973,N_9947,N_9806);
nand UO_974 (O_974,N_9778,N_9695);
or UO_975 (O_975,N_9588,N_9791);
nor UO_976 (O_976,N_9858,N_9856);
nand UO_977 (O_977,N_9999,N_9553);
nand UO_978 (O_978,N_9935,N_9537);
and UO_979 (O_979,N_9843,N_9535);
and UO_980 (O_980,N_9573,N_9975);
nand UO_981 (O_981,N_9711,N_9558);
nand UO_982 (O_982,N_9613,N_9686);
and UO_983 (O_983,N_9897,N_9691);
or UO_984 (O_984,N_9824,N_9605);
and UO_985 (O_985,N_9595,N_9618);
and UO_986 (O_986,N_9974,N_9706);
nor UO_987 (O_987,N_9788,N_9812);
or UO_988 (O_988,N_9964,N_9817);
xor UO_989 (O_989,N_9550,N_9591);
and UO_990 (O_990,N_9989,N_9986);
and UO_991 (O_991,N_9988,N_9740);
or UO_992 (O_992,N_9785,N_9517);
xor UO_993 (O_993,N_9665,N_9523);
xnor UO_994 (O_994,N_9573,N_9622);
and UO_995 (O_995,N_9621,N_9767);
xnor UO_996 (O_996,N_9721,N_9662);
xnor UO_997 (O_997,N_9805,N_9722);
nand UO_998 (O_998,N_9710,N_9978);
and UO_999 (O_999,N_9851,N_9956);
or UO_1000 (O_1000,N_9680,N_9601);
nand UO_1001 (O_1001,N_9623,N_9786);
and UO_1002 (O_1002,N_9541,N_9506);
xor UO_1003 (O_1003,N_9549,N_9608);
nor UO_1004 (O_1004,N_9588,N_9600);
nor UO_1005 (O_1005,N_9603,N_9642);
xnor UO_1006 (O_1006,N_9503,N_9788);
or UO_1007 (O_1007,N_9645,N_9532);
or UO_1008 (O_1008,N_9864,N_9516);
nor UO_1009 (O_1009,N_9593,N_9543);
nor UO_1010 (O_1010,N_9520,N_9505);
or UO_1011 (O_1011,N_9732,N_9725);
or UO_1012 (O_1012,N_9868,N_9725);
or UO_1013 (O_1013,N_9750,N_9737);
nor UO_1014 (O_1014,N_9862,N_9632);
or UO_1015 (O_1015,N_9984,N_9962);
nand UO_1016 (O_1016,N_9543,N_9597);
or UO_1017 (O_1017,N_9871,N_9969);
or UO_1018 (O_1018,N_9950,N_9869);
or UO_1019 (O_1019,N_9863,N_9597);
nand UO_1020 (O_1020,N_9546,N_9778);
and UO_1021 (O_1021,N_9754,N_9918);
xnor UO_1022 (O_1022,N_9946,N_9667);
and UO_1023 (O_1023,N_9635,N_9814);
nor UO_1024 (O_1024,N_9807,N_9736);
nand UO_1025 (O_1025,N_9530,N_9610);
nor UO_1026 (O_1026,N_9578,N_9893);
xnor UO_1027 (O_1027,N_9951,N_9683);
and UO_1028 (O_1028,N_9860,N_9688);
or UO_1029 (O_1029,N_9838,N_9973);
nor UO_1030 (O_1030,N_9874,N_9650);
xor UO_1031 (O_1031,N_9929,N_9937);
nand UO_1032 (O_1032,N_9972,N_9943);
xor UO_1033 (O_1033,N_9913,N_9513);
nor UO_1034 (O_1034,N_9837,N_9948);
nand UO_1035 (O_1035,N_9923,N_9549);
nor UO_1036 (O_1036,N_9612,N_9772);
xor UO_1037 (O_1037,N_9987,N_9765);
nand UO_1038 (O_1038,N_9914,N_9547);
xor UO_1039 (O_1039,N_9963,N_9512);
xor UO_1040 (O_1040,N_9835,N_9702);
and UO_1041 (O_1041,N_9710,N_9817);
or UO_1042 (O_1042,N_9768,N_9576);
or UO_1043 (O_1043,N_9684,N_9916);
or UO_1044 (O_1044,N_9931,N_9831);
xor UO_1045 (O_1045,N_9938,N_9872);
nand UO_1046 (O_1046,N_9737,N_9709);
or UO_1047 (O_1047,N_9929,N_9560);
nand UO_1048 (O_1048,N_9983,N_9711);
nor UO_1049 (O_1049,N_9621,N_9718);
nor UO_1050 (O_1050,N_9686,N_9592);
nor UO_1051 (O_1051,N_9883,N_9967);
nand UO_1052 (O_1052,N_9690,N_9579);
nor UO_1053 (O_1053,N_9560,N_9588);
nor UO_1054 (O_1054,N_9685,N_9891);
nand UO_1055 (O_1055,N_9601,N_9618);
nor UO_1056 (O_1056,N_9504,N_9562);
xor UO_1057 (O_1057,N_9957,N_9985);
nor UO_1058 (O_1058,N_9814,N_9777);
and UO_1059 (O_1059,N_9510,N_9685);
nand UO_1060 (O_1060,N_9627,N_9528);
and UO_1061 (O_1061,N_9703,N_9630);
nor UO_1062 (O_1062,N_9975,N_9662);
nor UO_1063 (O_1063,N_9990,N_9630);
nor UO_1064 (O_1064,N_9772,N_9511);
xor UO_1065 (O_1065,N_9575,N_9944);
nor UO_1066 (O_1066,N_9884,N_9980);
nand UO_1067 (O_1067,N_9843,N_9571);
and UO_1068 (O_1068,N_9506,N_9544);
and UO_1069 (O_1069,N_9954,N_9989);
xor UO_1070 (O_1070,N_9560,N_9846);
nor UO_1071 (O_1071,N_9727,N_9863);
or UO_1072 (O_1072,N_9615,N_9680);
or UO_1073 (O_1073,N_9531,N_9506);
nand UO_1074 (O_1074,N_9547,N_9644);
nor UO_1075 (O_1075,N_9632,N_9745);
xor UO_1076 (O_1076,N_9806,N_9766);
nor UO_1077 (O_1077,N_9636,N_9542);
nor UO_1078 (O_1078,N_9784,N_9924);
nand UO_1079 (O_1079,N_9557,N_9544);
xnor UO_1080 (O_1080,N_9928,N_9772);
and UO_1081 (O_1081,N_9820,N_9949);
nand UO_1082 (O_1082,N_9749,N_9598);
and UO_1083 (O_1083,N_9675,N_9910);
and UO_1084 (O_1084,N_9902,N_9957);
nor UO_1085 (O_1085,N_9750,N_9724);
and UO_1086 (O_1086,N_9694,N_9829);
nor UO_1087 (O_1087,N_9626,N_9940);
nor UO_1088 (O_1088,N_9502,N_9695);
and UO_1089 (O_1089,N_9509,N_9896);
nor UO_1090 (O_1090,N_9510,N_9589);
nor UO_1091 (O_1091,N_9774,N_9666);
nand UO_1092 (O_1092,N_9628,N_9695);
xor UO_1093 (O_1093,N_9957,N_9885);
nor UO_1094 (O_1094,N_9579,N_9607);
nor UO_1095 (O_1095,N_9982,N_9792);
nand UO_1096 (O_1096,N_9596,N_9854);
or UO_1097 (O_1097,N_9911,N_9789);
nand UO_1098 (O_1098,N_9802,N_9634);
and UO_1099 (O_1099,N_9883,N_9635);
nor UO_1100 (O_1100,N_9933,N_9660);
nand UO_1101 (O_1101,N_9669,N_9503);
or UO_1102 (O_1102,N_9562,N_9798);
nand UO_1103 (O_1103,N_9907,N_9555);
and UO_1104 (O_1104,N_9760,N_9651);
or UO_1105 (O_1105,N_9649,N_9856);
nand UO_1106 (O_1106,N_9742,N_9957);
or UO_1107 (O_1107,N_9893,N_9629);
xor UO_1108 (O_1108,N_9808,N_9625);
xnor UO_1109 (O_1109,N_9816,N_9771);
nand UO_1110 (O_1110,N_9988,N_9793);
or UO_1111 (O_1111,N_9646,N_9609);
or UO_1112 (O_1112,N_9517,N_9694);
and UO_1113 (O_1113,N_9654,N_9596);
or UO_1114 (O_1114,N_9959,N_9517);
nand UO_1115 (O_1115,N_9993,N_9741);
nor UO_1116 (O_1116,N_9723,N_9799);
nand UO_1117 (O_1117,N_9863,N_9821);
nand UO_1118 (O_1118,N_9582,N_9938);
or UO_1119 (O_1119,N_9855,N_9643);
and UO_1120 (O_1120,N_9777,N_9583);
nand UO_1121 (O_1121,N_9649,N_9517);
xor UO_1122 (O_1122,N_9852,N_9602);
xor UO_1123 (O_1123,N_9641,N_9546);
nand UO_1124 (O_1124,N_9614,N_9946);
xor UO_1125 (O_1125,N_9612,N_9657);
xnor UO_1126 (O_1126,N_9623,N_9826);
or UO_1127 (O_1127,N_9686,N_9600);
or UO_1128 (O_1128,N_9934,N_9716);
and UO_1129 (O_1129,N_9599,N_9517);
nand UO_1130 (O_1130,N_9959,N_9738);
nor UO_1131 (O_1131,N_9724,N_9618);
xor UO_1132 (O_1132,N_9705,N_9568);
and UO_1133 (O_1133,N_9530,N_9734);
xor UO_1134 (O_1134,N_9698,N_9946);
nand UO_1135 (O_1135,N_9667,N_9579);
or UO_1136 (O_1136,N_9648,N_9834);
xor UO_1137 (O_1137,N_9572,N_9660);
nand UO_1138 (O_1138,N_9777,N_9686);
nand UO_1139 (O_1139,N_9724,N_9982);
or UO_1140 (O_1140,N_9785,N_9973);
xnor UO_1141 (O_1141,N_9636,N_9574);
or UO_1142 (O_1142,N_9846,N_9870);
or UO_1143 (O_1143,N_9860,N_9573);
nand UO_1144 (O_1144,N_9722,N_9944);
xor UO_1145 (O_1145,N_9693,N_9792);
xor UO_1146 (O_1146,N_9817,N_9591);
or UO_1147 (O_1147,N_9899,N_9510);
xor UO_1148 (O_1148,N_9980,N_9534);
or UO_1149 (O_1149,N_9646,N_9849);
xnor UO_1150 (O_1150,N_9515,N_9805);
xnor UO_1151 (O_1151,N_9645,N_9724);
or UO_1152 (O_1152,N_9676,N_9951);
or UO_1153 (O_1153,N_9894,N_9712);
xor UO_1154 (O_1154,N_9679,N_9947);
nand UO_1155 (O_1155,N_9773,N_9809);
or UO_1156 (O_1156,N_9973,N_9630);
nand UO_1157 (O_1157,N_9664,N_9516);
nor UO_1158 (O_1158,N_9800,N_9956);
or UO_1159 (O_1159,N_9699,N_9953);
nor UO_1160 (O_1160,N_9614,N_9535);
nor UO_1161 (O_1161,N_9863,N_9591);
xor UO_1162 (O_1162,N_9572,N_9922);
nor UO_1163 (O_1163,N_9758,N_9663);
nand UO_1164 (O_1164,N_9952,N_9730);
xnor UO_1165 (O_1165,N_9766,N_9710);
and UO_1166 (O_1166,N_9875,N_9741);
nand UO_1167 (O_1167,N_9872,N_9662);
nand UO_1168 (O_1168,N_9832,N_9764);
and UO_1169 (O_1169,N_9542,N_9914);
xor UO_1170 (O_1170,N_9572,N_9882);
xor UO_1171 (O_1171,N_9510,N_9881);
and UO_1172 (O_1172,N_9743,N_9938);
xor UO_1173 (O_1173,N_9734,N_9664);
nand UO_1174 (O_1174,N_9633,N_9545);
and UO_1175 (O_1175,N_9690,N_9548);
and UO_1176 (O_1176,N_9791,N_9590);
nand UO_1177 (O_1177,N_9691,N_9793);
nor UO_1178 (O_1178,N_9905,N_9950);
xnor UO_1179 (O_1179,N_9873,N_9723);
xnor UO_1180 (O_1180,N_9878,N_9950);
xnor UO_1181 (O_1181,N_9518,N_9728);
and UO_1182 (O_1182,N_9618,N_9637);
nand UO_1183 (O_1183,N_9848,N_9809);
nand UO_1184 (O_1184,N_9734,N_9803);
xor UO_1185 (O_1185,N_9508,N_9832);
and UO_1186 (O_1186,N_9975,N_9841);
and UO_1187 (O_1187,N_9601,N_9648);
xor UO_1188 (O_1188,N_9517,N_9736);
xnor UO_1189 (O_1189,N_9985,N_9526);
xor UO_1190 (O_1190,N_9993,N_9809);
and UO_1191 (O_1191,N_9711,N_9614);
or UO_1192 (O_1192,N_9625,N_9571);
nand UO_1193 (O_1193,N_9524,N_9602);
xnor UO_1194 (O_1194,N_9817,N_9798);
nand UO_1195 (O_1195,N_9672,N_9679);
nor UO_1196 (O_1196,N_9903,N_9875);
nand UO_1197 (O_1197,N_9605,N_9914);
nand UO_1198 (O_1198,N_9974,N_9668);
and UO_1199 (O_1199,N_9946,N_9886);
nand UO_1200 (O_1200,N_9702,N_9955);
nand UO_1201 (O_1201,N_9953,N_9717);
and UO_1202 (O_1202,N_9686,N_9820);
or UO_1203 (O_1203,N_9714,N_9670);
nor UO_1204 (O_1204,N_9570,N_9968);
nor UO_1205 (O_1205,N_9848,N_9612);
nor UO_1206 (O_1206,N_9941,N_9543);
nor UO_1207 (O_1207,N_9824,N_9573);
and UO_1208 (O_1208,N_9957,N_9642);
nor UO_1209 (O_1209,N_9573,N_9781);
nor UO_1210 (O_1210,N_9668,N_9695);
or UO_1211 (O_1211,N_9718,N_9673);
and UO_1212 (O_1212,N_9822,N_9859);
or UO_1213 (O_1213,N_9786,N_9652);
nor UO_1214 (O_1214,N_9867,N_9780);
and UO_1215 (O_1215,N_9671,N_9669);
xnor UO_1216 (O_1216,N_9911,N_9585);
nor UO_1217 (O_1217,N_9906,N_9908);
nand UO_1218 (O_1218,N_9522,N_9893);
xnor UO_1219 (O_1219,N_9612,N_9595);
or UO_1220 (O_1220,N_9828,N_9745);
and UO_1221 (O_1221,N_9665,N_9792);
nand UO_1222 (O_1222,N_9849,N_9806);
or UO_1223 (O_1223,N_9838,N_9675);
or UO_1224 (O_1224,N_9973,N_9673);
or UO_1225 (O_1225,N_9757,N_9695);
nor UO_1226 (O_1226,N_9760,N_9544);
nor UO_1227 (O_1227,N_9775,N_9656);
and UO_1228 (O_1228,N_9854,N_9753);
or UO_1229 (O_1229,N_9889,N_9545);
and UO_1230 (O_1230,N_9815,N_9710);
xnor UO_1231 (O_1231,N_9785,N_9995);
nand UO_1232 (O_1232,N_9716,N_9632);
and UO_1233 (O_1233,N_9610,N_9904);
nand UO_1234 (O_1234,N_9776,N_9860);
xor UO_1235 (O_1235,N_9812,N_9835);
xnor UO_1236 (O_1236,N_9946,N_9956);
or UO_1237 (O_1237,N_9714,N_9838);
or UO_1238 (O_1238,N_9779,N_9655);
or UO_1239 (O_1239,N_9646,N_9781);
or UO_1240 (O_1240,N_9979,N_9533);
xnor UO_1241 (O_1241,N_9745,N_9583);
or UO_1242 (O_1242,N_9651,N_9929);
xor UO_1243 (O_1243,N_9659,N_9910);
nor UO_1244 (O_1244,N_9898,N_9654);
xnor UO_1245 (O_1245,N_9751,N_9896);
nand UO_1246 (O_1246,N_9588,N_9911);
nor UO_1247 (O_1247,N_9834,N_9807);
nor UO_1248 (O_1248,N_9809,N_9502);
and UO_1249 (O_1249,N_9600,N_9769);
nand UO_1250 (O_1250,N_9523,N_9804);
nand UO_1251 (O_1251,N_9591,N_9873);
xor UO_1252 (O_1252,N_9834,N_9515);
nand UO_1253 (O_1253,N_9972,N_9507);
xor UO_1254 (O_1254,N_9948,N_9671);
xnor UO_1255 (O_1255,N_9659,N_9746);
nand UO_1256 (O_1256,N_9533,N_9822);
xor UO_1257 (O_1257,N_9556,N_9794);
nor UO_1258 (O_1258,N_9575,N_9983);
or UO_1259 (O_1259,N_9574,N_9756);
xor UO_1260 (O_1260,N_9672,N_9661);
or UO_1261 (O_1261,N_9707,N_9533);
xnor UO_1262 (O_1262,N_9836,N_9533);
nand UO_1263 (O_1263,N_9891,N_9687);
nor UO_1264 (O_1264,N_9774,N_9600);
nor UO_1265 (O_1265,N_9758,N_9629);
nor UO_1266 (O_1266,N_9672,N_9861);
nand UO_1267 (O_1267,N_9983,N_9777);
or UO_1268 (O_1268,N_9513,N_9991);
or UO_1269 (O_1269,N_9764,N_9778);
and UO_1270 (O_1270,N_9508,N_9796);
and UO_1271 (O_1271,N_9958,N_9534);
or UO_1272 (O_1272,N_9545,N_9963);
nand UO_1273 (O_1273,N_9911,N_9750);
and UO_1274 (O_1274,N_9915,N_9894);
nor UO_1275 (O_1275,N_9817,N_9766);
nor UO_1276 (O_1276,N_9658,N_9635);
nand UO_1277 (O_1277,N_9893,N_9581);
nor UO_1278 (O_1278,N_9969,N_9808);
or UO_1279 (O_1279,N_9579,N_9582);
xor UO_1280 (O_1280,N_9854,N_9956);
nor UO_1281 (O_1281,N_9827,N_9936);
or UO_1282 (O_1282,N_9758,N_9636);
xor UO_1283 (O_1283,N_9746,N_9603);
nor UO_1284 (O_1284,N_9786,N_9914);
nand UO_1285 (O_1285,N_9951,N_9588);
nand UO_1286 (O_1286,N_9674,N_9569);
and UO_1287 (O_1287,N_9573,N_9784);
nand UO_1288 (O_1288,N_9551,N_9653);
nand UO_1289 (O_1289,N_9710,N_9970);
or UO_1290 (O_1290,N_9799,N_9863);
and UO_1291 (O_1291,N_9964,N_9703);
or UO_1292 (O_1292,N_9528,N_9645);
nor UO_1293 (O_1293,N_9576,N_9548);
nor UO_1294 (O_1294,N_9884,N_9998);
xor UO_1295 (O_1295,N_9658,N_9804);
nor UO_1296 (O_1296,N_9868,N_9853);
nor UO_1297 (O_1297,N_9829,N_9729);
nor UO_1298 (O_1298,N_9992,N_9637);
nor UO_1299 (O_1299,N_9875,N_9998);
or UO_1300 (O_1300,N_9662,N_9751);
nor UO_1301 (O_1301,N_9741,N_9903);
xor UO_1302 (O_1302,N_9858,N_9796);
nand UO_1303 (O_1303,N_9765,N_9747);
nor UO_1304 (O_1304,N_9555,N_9654);
xor UO_1305 (O_1305,N_9524,N_9600);
nor UO_1306 (O_1306,N_9706,N_9762);
xor UO_1307 (O_1307,N_9911,N_9653);
and UO_1308 (O_1308,N_9562,N_9588);
xor UO_1309 (O_1309,N_9832,N_9898);
and UO_1310 (O_1310,N_9642,N_9713);
nor UO_1311 (O_1311,N_9858,N_9551);
nand UO_1312 (O_1312,N_9987,N_9535);
or UO_1313 (O_1313,N_9507,N_9851);
or UO_1314 (O_1314,N_9726,N_9776);
and UO_1315 (O_1315,N_9769,N_9642);
or UO_1316 (O_1316,N_9553,N_9572);
nor UO_1317 (O_1317,N_9746,N_9641);
nor UO_1318 (O_1318,N_9605,N_9788);
xnor UO_1319 (O_1319,N_9784,N_9674);
nor UO_1320 (O_1320,N_9864,N_9891);
or UO_1321 (O_1321,N_9527,N_9939);
nor UO_1322 (O_1322,N_9873,N_9890);
xnor UO_1323 (O_1323,N_9559,N_9985);
xor UO_1324 (O_1324,N_9663,N_9575);
nor UO_1325 (O_1325,N_9637,N_9799);
and UO_1326 (O_1326,N_9661,N_9912);
and UO_1327 (O_1327,N_9677,N_9978);
nand UO_1328 (O_1328,N_9990,N_9921);
nand UO_1329 (O_1329,N_9652,N_9843);
or UO_1330 (O_1330,N_9774,N_9648);
nand UO_1331 (O_1331,N_9710,N_9848);
xor UO_1332 (O_1332,N_9526,N_9602);
nand UO_1333 (O_1333,N_9661,N_9518);
nor UO_1334 (O_1334,N_9941,N_9845);
nor UO_1335 (O_1335,N_9720,N_9692);
nor UO_1336 (O_1336,N_9709,N_9780);
and UO_1337 (O_1337,N_9787,N_9601);
or UO_1338 (O_1338,N_9544,N_9681);
nor UO_1339 (O_1339,N_9524,N_9859);
xnor UO_1340 (O_1340,N_9529,N_9509);
and UO_1341 (O_1341,N_9820,N_9880);
nor UO_1342 (O_1342,N_9908,N_9682);
nand UO_1343 (O_1343,N_9932,N_9746);
nand UO_1344 (O_1344,N_9556,N_9993);
and UO_1345 (O_1345,N_9915,N_9970);
and UO_1346 (O_1346,N_9609,N_9547);
nor UO_1347 (O_1347,N_9831,N_9742);
nor UO_1348 (O_1348,N_9866,N_9620);
xor UO_1349 (O_1349,N_9935,N_9897);
and UO_1350 (O_1350,N_9522,N_9654);
nand UO_1351 (O_1351,N_9977,N_9950);
or UO_1352 (O_1352,N_9839,N_9584);
xor UO_1353 (O_1353,N_9731,N_9516);
and UO_1354 (O_1354,N_9817,N_9876);
xnor UO_1355 (O_1355,N_9869,N_9623);
nor UO_1356 (O_1356,N_9728,N_9624);
xor UO_1357 (O_1357,N_9771,N_9600);
xor UO_1358 (O_1358,N_9881,N_9591);
nand UO_1359 (O_1359,N_9932,N_9872);
and UO_1360 (O_1360,N_9898,N_9956);
nor UO_1361 (O_1361,N_9832,N_9700);
nor UO_1362 (O_1362,N_9922,N_9606);
xnor UO_1363 (O_1363,N_9883,N_9724);
nor UO_1364 (O_1364,N_9719,N_9721);
and UO_1365 (O_1365,N_9838,N_9972);
nor UO_1366 (O_1366,N_9877,N_9618);
or UO_1367 (O_1367,N_9504,N_9973);
and UO_1368 (O_1368,N_9569,N_9596);
nor UO_1369 (O_1369,N_9683,N_9953);
or UO_1370 (O_1370,N_9813,N_9741);
nor UO_1371 (O_1371,N_9749,N_9631);
and UO_1372 (O_1372,N_9839,N_9569);
nor UO_1373 (O_1373,N_9633,N_9918);
nor UO_1374 (O_1374,N_9894,N_9636);
nor UO_1375 (O_1375,N_9653,N_9876);
or UO_1376 (O_1376,N_9528,N_9587);
nand UO_1377 (O_1377,N_9866,N_9603);
nor UO_1378 (O_1378,N_9730,N_9980);
and UO_1379 (O_1379,N_9803,N_9756);
nand UO_1380 (O_1380,N_9790,N_9794);
and UO_1381 (O_1381,N_9547,N_9966);
nand UO_1382 (O_1382,N_9636,N_9548);
and UO_1383 (O_1383,N_9527,N_9733);
nor UO_1384 (O_1384,N_9737,N_9782);
nor UO_1385 (O_1385,N_9780,N_9884);
xnor UO_1386 (O_1386,N_9983,N_9952);
xor UO_1387 (O_1387,N_9616,N_9948);
xor UO_1388 (O_1388,N_9968,N_9722);
and UO_1389 (O_1389,N_9996,N_9908);
xnor UO_1390 (O_1390,N_9982,N_9686);
xor UO_1391 (O_1391,N_9653,N_9852);
nor UO_1392 (O_1392,N_9872,N_9865);
and UO_1393 (O_1393,N_9590,N_9765);
nor UO_1394 (O_1394,N_9986,N_9616);
and UO_1395 (O_1395,N_9786,N_9693);
xor UO_1396 (O_1396,N_9661,N_9956);
or UO_1397 (O_1397,N_9895,N_9585);
or UO_1398 (O_1398,N_9767,N_9727);
xor UO_1399 (O_1399,N_9879,N_9917);
or UO_1400 (O_1400,N_9808,N_9740);
nand UO_1401 (O_1401,N_9557,N_9860);
or UO_1402 (O_1402,N_9651,N_9766);
nor UO_1403 (O_1403,N_9545,N_9646);
nor UO_1404 (O_1404,N_9617,N_9663);
and UO_1405 (O_1405,N_9954,N_9544);
or UO_1406 (O_1406,N_9751,N_9678);
nor UO_1407 (O_1407,N_9754,N_9633);
or UO_1408 (O_1408,N_9690,N_9597);
xor UO_1409 (O_1409,N_9970,N_9673);
and UO_1410 (O_1410,N_9736,N_9677);
nand UO_1411 (O_1411,N_9804,N_9860);
nand UO_1412 (O_1412,N_9656,N_9554);
or UO_1413 (O_1413,N_9700,N_9706);
nor UO_1414 (O_1414,N_9649,N_9756);
or UO_1415 (O_1415,N_9745,N_9857);
and UO_1416 (O_1416,N_9505,N_9851);
xor UO_1417 (O_1417,N_9813,N_9653);
and UO_1418 (O_1418,N_9875,N_9951);
or UO_1419 (O_1419,N_9921,N_9826);
and UO_1420 (O_1420,N_9953,N_9657);
or UO_1421 (O_1421,N_9985,N_9619);
xor UO_1422 (O_1422,N_9569,N_9915);
or UO_1423 (O_1423,N_9679,N_9973);
xnor UO_1424 (O_1424,N_9651,N_9893);
xor UO_1425 (O_1425,N_9766,N_9671);
nand UO_1426 (O_1426,N_9728,N_9643);
and UO_1427 (O_1427,N_9713,N_9623);
and UO_1428 (O_1428,N_9648,N_9673);
xnor UO_1429 (O_1429,N_9621,N_9861);
nor UO_1430 (O_1430,N_9731,N_9699);
nor UO_1431 (O_1431,N_9947,N_9789);
or UO_1432 (O_1432,N_9695,N_9748);
or UO_1433 (O_1433,N_9619,N_9531);
xnor UO_1434 (O_1434,N_9777,N_9900);
xnor UO_1435 (O_1435,N_9551,N_9694);
nand UO_1436 (O_1436,N_9629,N_9847);
or UO_1437 (O_1437,N_9913,N_9559);
nand UO_1438 (O_1438,N_9716,N_9784);
and UO_1439 (O_1439,N_9748,N_9699);
and UO_1440 (O_1440,N_9704,N_9522);
nand UO_1441 (O_1441,N_9932,N_9709);
nor UO_1442 (O_1442,N_9997,N_9637);
and UO_1443 (O_1443,N_9565,N_9938);
nand UO_1444 (O_1444,N_9642,N_9958);
nor UO_1445 (O_1445,N_9569,N_9992);
and UO_1446 (O_1446,N_9774,N_9746);
and UO_1447 (O_1447,N_9524,N_9937);
xnor UO_1448 (O_1448,N_9896,N_9638);
nor UO_1449 (O_1449,N_9524,N_9958);
or UO_1450 (O_1450,N_9529,N_9708);
and UO_1451 (O_1451,N_9966,N_9737);
nand UO_1452 (O_1452,N_9607,N_9864);
xnor UO_1453 (O_1453,N_9949,N_9644);
and UO_1454 (O_1454,N_9757,N_9632);
nand UO_1455 (O_1455,N_9715,N_9831);
nand UO_1456 (O_1456,N_9837,N_9823);
xnor UO_1457 (O_1457,N_9839,N_9917);
nand UO_1458 (O_1458,N_9983,N_9809);
or UO_1459 (O_1459,N_9927,N_9801);
or UO_1460 (O_1460,N_9548,N_9522);
nor UO_1461 (O_1461,N_9715,N_9720);
nor UO_1462 (O_1462,N_9697,N_9917);
nand UO_1463 (O_1463,N_9862,N_9963);
xor UO_1464 (O_1464,N_9777,N_9541);
and UO_1465 (O_1465,N_9613,N_9952);
and UO_1466 (O_1466,N_9719,N_9513);
nor UO_1467 (O_1467,N_9744,N_9578);
nand UO_1468 (O_1468,N_9807,N_9890);
and UO_1469 (O_1469,N_9634,N_9667);
and UO_1470 (O_1470,N_9754,N_9890);
nand UO_1471 (O_1471,N_9578,N_9649);
xor UO_1472 (O_1472,N_9645,N_9578);
or UO_1473 (O_1473,N_9845,N_9985);
nor UO_1474 (O_1474,N_9672,N_9932);
and UO_1475 (O_1475,N_9879,N_9978);
nor UO_1476 (O_1476,N_9517,N_9982);
or UO_1477 (O_1477,N_9904,N_9617);
or UO_1478 (O_1478,N_9849,N_9702);
or UO_1479 (O_1479,N_9844,N_9964);
nor UO_1480 (O_1480,N_9806,N_9677);
nor UO_1481 (O_1481,N_9806,N_9736);
xor UO_1482 (O_1482,N_9547,N_9793);
or UO_1483 (O_1483,N_9525,N_9943);
xor UO_1484 (O_1484,N_9761,N_9763);
nand UO_1485 (O_1485,N_9588,N_9726);
xnor UO_1486 (O_1486,N_9594,N_9840);
xor UO_1487 (O_1487,N_9904,N_9866);
nor UO_1488 (O_1488,N_9688,N_9917);
nand UO_1489 (O_1489,N_9911,N_9906);
nor UO_1490 (O_1490,N_9521,N_9765);
nor UO_1491 (O_1491,N_9554,N_9575);
xnor UO_1492 (O_1492,N_9588,N_9904);
and UO_1493 (O_1493,N_9570,N_9727);
or UO_1494 (O_1494,N_9523,N_9708);
nand UO_1495 (O_1495,N_9873,N_9952);
xor UO_1496 (O_1496,N_9640,N_9940);
nand UO_1497 (O_1497,N_9575,N_9814);
nand UO_1498 (O_1498,N_9638,N_9605);
and UO_1499 (O_1499,N_9847,N_9598);
endmodule