module basic_500_3000_500_4_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_307,In_54);
or U1 (N_1,In_427,In_197);
and U2 (N_2,In_315,In_13);
nor U3 (N_3,In_360,In_138);
nor U4 (N_4,In_388,In_278);
or U5 (N_5,In_24,In_372);
nand U6 (N_6,In_120,In_414);
or U7 (N_7,In_119,In_135);
or U8 (N_8,In_469,In_123);
and U9 (N_9,In_96,In_437);
nor U10 (N_10,In_464,In_431);
xnor U11 (N_11,In_29,In_277);
nand U12 (N_12,In_370,In_271);
or U13 (N_13,In_454,In_82);
nand U14 (N_14,In_64,In_199);
or U15 (N_15,In_268,In_171);
or U16 (N_16,In_381,In_185);
or U17 (N_17,In_39,In_352);
nand U18 (N_18,In_239,In_311);
xor U19 (N_19,In_12,In_168);
or U20 (N_20,In_46,In_43);
and U21 (N_21,In_3,In_403);
nand U22 (N_22,In_48,In_457);
and U23 (N_23,In_468,In_139);
or U24 (N_24,In_371,In_72);
and U25 (N_25,In_65,In_250);
nor U26 (N_26,In_182,In_481);
and U27 (N_27,In_1,In_460);
nand U28 (N_28,In_187,In_318);
nand U29 (N_29,In_312,In_261);
nor U30 (N_30,In_462,In_230);
xor U31 (N_31,In_188,In_225);
nand U32 (N_32,In_426,In_68);
nor U33 (N_33,In_452,In_249);
nand U34 (N_34,In_215,In_38);
nand U35 (N_35,In_100,In_145);
nand U36 (N_36,In_206,In_321);
nor U37 (N_37,In_450,In_105);
nand U38 (N_38,In_183,In_297);
or U39 (N_39,In_242,In_156);
and U40 (N_40,In_150,In_329);
nor U41 (N_41,In_298,In_430);
nor U42 (N_42,In_164,In_229);
nand U43 (N_43,In_127,In_303);
and U44 (N_44,In_251,In_418);
nand U45 (N_45,In_219,In_165);
or U46 (N_46,In_198,In_305);
nor U47 (N_47,In_289,In_326);
or U48 (N_48,In_483,In_333);
nor U49 (N_49,In_398,In_196);
nor U50 (N_50,In_233,In_223);
nand U51 (N_51,In_304,In_118);
xor U52 (N_52,In_319,In_189);
nor U53 (N_53,In_415,In_73);
nand U54 (N_54,In_163,In_83);
and U55 (N_55,In_327,In_287);
nor U56 (N_56,In_152,In_461);
and U57 (N_57,In_349,In_9);
nand U58 (N_58,In_47,In_423);
or U59 (N_59,In_476,In_413);
nand U60 (N_60,In_109,In_148);
or U61 (N_61,In_143,In_86);
and U62 (N_62,In_190,In_272);
and U63 (N_63,In_201,In_8);
or U64 (N_64,In_125,In_436);
xnor U65 (N_65,In_320,In_290);
and U66 (N_66,In_309,In_161);
and U67 (N_67,In_107,In_131);
or U68 (N_68,In_15,In_244);
nand U69 (N_69,In_301,In_324);
and U70 (N_70,In_387,In_181);
or U71 (N_71,In_399,In_466);
or U72 (N_72,In_358,In_400);
nor U73 (N_73,In_63,In_367);
nor U74 (N_74,In_151,In_11);
nor U75 (N_75,In_353,In_31);
xor U76 (N_76,In_422,In_276);
nor U77 (N_77,In_255,In_248);
and U78 (N_78,In_232,In_222);
nand U79 (N_79,In_240,In_204);
or U80 (N_80,In_2,In_193);
nand U81 (N_81,In_51,In_459);
and U82 (N_82,In_19,In_499);
nor U83 (N_83,In_97,In_18);
and U84 (N_84,In_32,In_20);
nand U85 (N_85,In_497,In_59);
or U86 (N_86,In_256,In_420);
nand U87 (N_87,In_159,In_465);
nor U88 (N_88,In_378,In_217);
and U89 (N_89,In_75,In_491);
nand U90 (N_90,In_50,In_410);
nor U91 (N_91,In_137,In_402);
nor U92 (N_92,In_220,In_155);
or U93 (N_93,In_392,In_207);
and U94 (N_94,In_254,In_458);
nor U95 (N_95,In_425,In_98);
nand U96 (N_96,In_213,In_103);
nor U97 (N_97,In_373,In_494);
nor U98 (N_98,In_473,In_69);
or U99 (N_99,In_58,In_478);
or U100 (N_100,In_322,In_306);
or U101 (N_101,In_455,In_283);
xnor U102 (N_102,In_179,In_282);
and U103 (N_103,In_295,In_325);
nand U104 (N_104,In_344,In_285);
nor U105 (N_105,In_132,In_88);
or U106 (N_106,In_55,In_406);
nor U107 (N_107,In_379,In_172);
nor U108 (N_108,In_157,In_269);
nor U109 (N_109,In_264,In_258);
and U110 (N_110,In_30,In_112);
nor U111 (N_111,In_361,In_375);
nand U112 (N_112,In_108,In_409);
nand U113 (N_113,In_253,In_210);
nor U114 (N_114,In_343,In_49);
nand U115 (N_115,In_71,In_0);
and U116 (N_116,In_76,In_173);
or U117 (N_117,In_70,In_487);
nand U118 (N_118,In_401,In_167);
and U119 (N_119,In_374,In_121);
and U120 (N_120,In_323,In_60);
xor U121 (N_121,In_84,In_42);
and U122 (N_122,In_192,In_85);
and U123 (N_123,In_36,In_302);
nor U124 (N_124,In_292,In_376);
nor U125 (N_125,In_257,In_140);
or U126 (N_126,In_16,In_262);
nor U127 (N_127,In_175,In_265);
or U128 (N_128,In_448,In_300);
or U129 (N_129,In_133,In_154);
nor U130 (N_130,In_275,In_291);
nand U131 (N_131,In_439,In_432);
and U132 (N_132,In_234,In_160);
nand U133 (N_133,In_61,In_449);
nand U134 (N_134,In_383,In_260);
nand U135 (N_135,In_62,In_359);
xor U136 (N_136,In_332,In_447);
or U137 (N_137,In_328,In_417);
nor U138 (N_138,In_479,In_77);
xor U139 (N_139,In_263,In_40);
nand U140 (N_140,In_453,In_92);
and U141 (N_141,In_52,In_27);
nor U142 (N_142,In_488,In_6);
nand U143 (N_143,In_308,In_365);
nor U144 (N_144,In_480,In_441);
and U145 (N_145,In_477,In_407);
nor U146 (N_146,In_310,In_243);
nand U147 (N_147,In_184,In_110);
xnor U148 (N_148,In_396,In_341);
and U149 (N_149,In_471,In_424);
or U150 (N_150,In_435,In_363);
or U151 (N_151,In_362,In_246);
or U152 (N_152,In_386,In_158);
or U153 (N_153,In_390,In_394);
nand U154 (N_154,In_443,In_470);
nor U155 (N_155,In_177,In_433);
or U156 (N_156,In_115,In_10);
or U157 (N_157,In_66,In_408);
nand U158 (N_158,In_218,In_421);
or U159 (N_159,In_203,In_124);
and U160 (N_160,In_279,In_99);
and U161 (N_161,In_153,In_377);
or U162 (N_162,In_34,In_330);
nor U163 (N_163,In_380,In_147);
and U164 (N_164,In_274,In_366);
nor U165 (N_165,In_128,In_419);
or U166 (N_166,In_126,In_354);
nand U167 (N_167,In_17,In_474);
or U168 (N_168,In_384,In_475);
nor U169 (N_169,In_434,In_369);
nor U170 (N_170,In_364,In_162);
nor U171 (N_171,In_445,In_208);
nor U172 (N_172,In_247,In_80);
or U173 (N_173,In_89,In_116);
nand U174 (N_174,In_486,In_245);
nor U175 (N_175,In_288,In_14);
nand U176 (N_176,In_170,In_5);
nand U177 (N_177,In_94,In_498);
nand U178 (N_178,In_337,In_440);
nor U179 (N_179,In_180,In_281);
nor U180 (N_180,In_382,In_438);
and U181 (N_181,In_467,In_214);
and U182 (N_182,In_385,In_489);
nor U183 (N_183,In_241,In_25);
nand U184 (N_184,In_451,In_259);
xnor U185 (N_185,In_482,In_492);
and U186 (N_186,In_235,In_444);
nor U187 (N_187,In_273,In_356);
nand U188 (N_188,In_228,In_284);
nand U189 (N_189,In_429,In_490);
nor U190 (N_190,In_174,In_91);
or U191 (N_191,In_205,In_238);
and U192 (N_192,In_79,In_212);
xnor U193 (N_193,In_227,In_348);
nand U194 (N_194,In_340,In_87);
nor U195 (N_195,In_130,In_495);
nand U196 (N_196,In_405,In_252);
nand U197 (N_197,In_22,In_221);
nor U198 (N_198,In_339,In_56);
nor U199 (N_199,In_136,In_67);
or U200 (N_200,In_313,In_294);
nor U201 (N_201,In_334,In_114);
and U202 (N_202,In_316,In_21);
nor U203 (N_203,In_57,In_368);
or U204 (N_204,In_37,In_293);
or U205 (N_205,In_496,In_93);
and U206 (N_206,In_347,In_53);
nand U207 (N_207,In_416,In_393);
nor U208 (N_208,In_28,In_141);
nor U209 (N_209,In_270,In_178);
nor U210 (N_210,In_144,In_209);
or U211 (N_211,In_331,In_104);
and U212 (N_212,In_391,In_346);
or U213 (N_213,In_355,In_314);
nor U214 (N_214,In_122,In_299);
or U215 (N_215,In_194,In_351);
and U216 (N_216,In_134,In_412);
nor U217 (N_217,In_428,In_336);
nor U218 (N_218,In_113,In_101);
nand U219 (N_219,In_237,In_166);
nand U220 (N_220,In_146,In_231);
nor U221 (N_221,In_456,In_280);
nand U222 (N_222,In_463,In_266);
or U223 (N_223,In_357,In_397);
nor U224 (N_224,In_395,In_117);
and U225 (N_225,In_44,In_211);
or U226 (N_226,In_267,In_200);
and U227 (N_227,In_191,In_106);
xor U228 (N_228,In_129,In_23);
nand U229 (N_229,In_176,In_286);
or U230 (N_230,In_111,In_26);
and U231 (N_231,In_45,In_102);
and U232 (N_232,In_484,In_317);
or U233 (N_233,In_345,In_335);
nand U234 (N_234,In_169,In_90);
and U235 (N_235,In_224,In_81);
xor U236 (N_236,In_202,In_95);
nor U237 (N_237,In_41,In_404);
xor U238 (N_238,In_389,In_74);
nor U239 (N_239,In_186,In_226);
or U240 (N_240,In_342,In_411);
nor U241 (N_241,In_442,In_350);
xnor U242 (N_242,In_296,In_35);
and U243 (N_243,In_446,In_216);
nor U244 (N_244,In_485,In_33);
and U245 (N_245,In_7,In_78);
or U246 (N_246,In_4,In_338);
or U247 (N_247,In_149,In_493);
nor U248 (N_248,In_195,In_472);
or U249 (N_249,In_142,In_236);
nor U250 (N_250,In_452,In_63);
nand U251 (N_251,In_217,In_411);
and U252 (N_252,In_59,In_18);
or U253 (N_253,In_232,In_241);
nor U254 (N_254,In_74,In_116);
or U255 (N_255,In_95,In_46);
and U256 (N_256,In_160,In_190);
nand U257 (N_257,In_91,In_418);
xor U258 (N_258,In_196,In_25);
nand U259 (N_259,In_97,In_327);
nand U260 (N_260,In_355,In_190);
nand U261 (N_261,In_322,In_128);
nand U262 (N_262,In_464,In_116);
nor U263 (N_263,In_386,In_466);
xnor U264 (N_264,In_219,In_442);
xnor U265 (N_265,In_336,In_474);
and U266 (N_266,In_322,In_113);
nand U267 (N_267,In_323,In_90);
nor U268 (N_268,In_336,In_359);
or U269 (N_269,In_84,In_356);
or U270 (N_270,In_464,In_253);
nor U271 (N_271,In_9,In_10);
nand U272 (N_272,In_129,In_0);
nand U273 (N_273,In_119,In_284);
nand U274 (N_274,In_66,In_120);
or U275 (N_275,In_254,In_188);
xnor U276 (N_276,In_211,In_460);
or U277 (N_277,In_336,In_35);
nand U278 (N_278,In_29,In_332);
nand U279 (N_279,In_309,In_287);
nor U280 (N_280,In_183,In_425);
nand U281 (N_281,In_315,In_341);
or U282 (N_282,In_426,In_360);
nand U283 (N_283,In_226,In_21);
nand U284 (N_284,In_400,In_364);
or U285 (N_285,In_178,In_166);
nand U286 (N_286,In_269,In_391);
nor U287 (N_287,In_152,In_358);
nor U288 (N_288,In_47,In_327);
or U289 (N_289,In_417,In_496);
xor U290 (N_290,In_168,In_45);
nand U291 (N_291,In_468,In_37);
or U292 (N_292,In_32,In_69);
nand U293 (N_293,In_83,In_253);
nand U294 (N_294,In_177,In_431);
nor U295 (N_295,In_209,In_183);
xnor U296 (N_296,In_174,In_119);
or U297 (N_297,In_307,In_110);
or U298 (N_298,In_210,In_289);
nor U299 (N_299,In_99,In_414);
and U300 (N_300,In_190,In_88);
and U301 (N_301,In_442,In_449);
and U302 (N_302,In_380,In_214);
nor U303 (N_303,In_45,In_491);
or U304 (N_304,In_158,In_259);
nand U305 (N_305,In_181,In_157);
nor U306 (N_306,In_279,In_10);
or U307 (N_307,In_422,In_215);
xor U308 (N_308,In_299,In_498);
nand U309 (N_309,In_324,In_363);
nor U310 (N_310,In_131,In_267);
and U311 (N_311,In_132,In_107);
nand U312 (N_312,In_435,In_176);
nor U313 (N_313,In_260,In_406);
nor U314 (N_314,In_316,In_255);
and U315 (N_315,In_122,In_363);
nor U316 (N_316,In_370,In_153);
xnor U317 (N_317,In_48,In_369);
or U318 (N_318,In_173,In_70);
nor U319 (N_319,In_255,In_299);
xnor U320 (N_320,In_420,In_204);
and U321 (N_321,In_72,In_0);
nor U322 (N_322,In_316,In_174);
xnor U323 (N_323,In_202,In_423);
nor U324 (N_324,In_372,In_214);
nor U325 (N_325,In_79,In_168);
and U326 (N_326,In_410,In_180);
nor U327 (N_327,In_210,In_74);
nor U328 (N_328,In_137,In_294);
nor U329 (N_329,In_67,In_361);
nand U330 (N_330,In_268,In_21);
nand U331 (N_331,In_441,In_353);
and U332 (N_332,In_485,In_280);
nor U333 (N_333,In_391,In_499);
or U334 (N_334,In_130,In_488);
or U335 (N_335,In_395,In_201);
nor U336 (N_336,In_397,In_68);
nand U337 (N_337,In_143,In_368);
xor U338 (N_338,In_395,In_409);
xnor U339 (N_339,In_430,In_66);
and U340 (N_340,In_331,In_141);
xnor U341 (N_341,In_467,In_477);
and U342 (N_342,In_333,In_116);
or U343 (N_343,In_339,In_264);
nand U344 (N_344,In_163,In_211);
and U345 (N_345,In_5,In_81);
nor U346 (N_346,In_251,In_398);
and U347 (N_347,In_308,In_42);
or U348 (N_348,In_405,In_254);
nand U349 (N_349,In_82,In_282);
or U350 (N_350,In_52,In_321);
nor U351 (N_351,In_138,In_342);
and U352 (N_352,In_258,In_277);
and U353 (N_353,In_86,In_436);
or U354 (N_354,In_154,In_438);
and U355 (N_355,In_492,In_419);
xor U356 (N_356,In_324,In_328);
nor U357 (N_357,In_232,In_204);
or U358 (N_358,In_153,In_363);
and U359 (N_359,In_6,In_21);
or U360 (N_360,In_100,In_303);
and U361 (N_361,In_12,In_471);
nand U362 (N_362,In_197,In_103);
nor U363 (N_363,In_211,In_72);
or U364 (N_364,In_181,In_277);
and U365 (N_365,In_474,In_186);
and U366 (N_366,In_17,In_382);
nand U367 (N_367,In_403,In_463);
nor U368 (N_368,In_11,In_141);
or U369 (N_369,In_482,In_485);
nor U370 (N_370,In_204,In_469);
nor U371 (N_371,In_205,In_415);
nand U372 (N_372,In_151,In_226);
nand U373 (N_373,In_464,In_157);
and U374 (N_374,In_459,In_101);
or U375 (N_375,In_131,In_163);
nor U376 (N_376,In_477,In_330);
and U377 (N_377,In_115,In_312);
nor U378 (N_378,In_233,In_31);
nand U379 (N_379,In_400,In_195);
nand U380 (N_380,In_293,In_44);
nand U381 (N_381,In_468,In_46);
nor U382 (N_382,In_498,In_54);
nand U383 (N_383,In_433,In_311);
nand U384 (N_384,In_317,In_424);
nor U385 (N_385,In_184,In_120);
or U386 (N_386,In_486,In_283);
nand U387 (N_387,In_13,In_304);
nor U388 (N_388,In_142,In_472);
nand U389 (N_389,In_87,In_368);
nor U390 (N_390,In_441,In_137);
nor U391 (N_391,In_64,In_50);
and U392 (N_392,In_4,In_241);
nand U393 (N_393,In_399,In_52);
or U394 (N_394,In_270,In_192);
nand U395 (N_395,In_281,In_294);
nor U396 (N_396,In_313,In_239);
nor U397 (N_397,In_363,In_28);
xor U398 (N_398,In_371,In_25);
or U399 (N_399,In_32,In_113);
and U400 (N_400,In_273,In_8);
and U401 (N_401,In_233,In_427);
nand U402 (N_402,In_167,In_262);
nand U403 (N_403,In_324,In_177);
nor U404 (N_404,In_183,In_422);
and U405 (N_405,In_481,In_79);
nor U406 (N_406,In_313,In_216);
nand U407 (N_407,In_231,In_265);
and U408 (N_408,In_224,In_79);
nor U409 (N_409,In_95,In_89);
nand U410 (N_410,In_206,In_458);
nand U411 (N_411,In_55,In_124);
nor U412 (N_412,In_301,In_232);
nor U413 (N_413,In_319,In_487);
nor U414 (N_414,In_472,In_229);
and U415 (N_415,In_412,In_484);
nand U416 (N_416,In_371,In_299);
nand U417 (N_417,In_80,In_258);
nor U418 (N_418,In_403,In_68);
nor U419 (N_419,In_350,In_418);
nor U420 (N_420,In_329,In_49);
or U421 (N_421,In_277,In_45);
nor U422 (N_422,In_327,In_89);
nor U423 (N_423,In_281,In_41);
and U424 (N_424,In_241,In_113);
nand U425 (N_425,In_475,In_418);
nand U426 (N_426,In_450,In_357);
and U427 (N_427,In_407,In_351);
and U428 (N_428,In_71,In_221);
xor U429 (N_429,In_23,In_92);
nand U430 (N_430,In_113,In_168);
nor U431 (N_431,In_365,In_264);
nor U432 (N_432,In_307,In_163);
or U433 (N_433,In_405,In_487);
or U434 (N_434,In_282,In_252);
nand U435 (N_435,In_236,In_375);
nor U436 (N_436,In_351,In_390);
and U437 (N_437,In_331,In_376);
nand U438 (N_438,In_267,In_300);
nand U439 (N_439,In_13,In_206);
or U440 (N_440,In_129,In_391);
xnor U441 (N_441,In_333,In_364);
nand U442 (N_442,In_409,In_365);
or U443 (N_443,In_251,In_215);
nor U444 (N_444,In_57,In_116);
nand U445 (N_445,In_47,In_201);
and U446 (N_446,In_28,In_491);
xor U447 (N_447,In_487,In_240);
or U448 (N_448,In_192,In_91);
and U449 (N_449,In_141,In_167);
or U450 (N_450,In_97,In_105);
nor U451 (N_451,In_29,In_283);
xor U452 (N_452,In_351,In_184);
xor U453 (N_453,In_53,In_147);
nor U454 (N_454,In_26,In_48);
or U455 (N_455,In_209,In_179);
nand U456 (N_456,In_389,In_129);
and U457 (N_457,In_213,In_39);
xor U458 (N_458,In_404,In_62);
nand U459 (N_459,In_130,In_364);
or U460 (N_460,In_131,In_134);
and U461 (N_461,In_104,In_34);
nand U462 (N_462,In_248,In_120);
and U463 (N_463,In_197,In_183);
or U464 (N_464,In_130,In_155);
nand U465 (N_465,In_463,In_50);
or U466 (N_466,In_109,In_210);
xor U467 (N_467,In_347,In_247);
nor U468 (N_468,In_343,In_60);
nor U469 (N_469,In_367,In_173);
nor U470 (N_470,In_415,In_346);
nand U471 (N_471,In_5,In_277);
or U472 (N_472,In_78,In_446);
and U473 (N_473,In_136,In_265);
nor U474 (N_474,In_375,In_172);
or U475 (N_475,In_166,In_76);
nor U476 (N_476,In_109,In_427);
and U477 (N_477,In_276,In_40);
nor U478 (N_478,In_32,In_83);
or U479 (N_479,In_118,In_263);
nand U480 (N_480,In_492,In_326);
nor U481 (N_481,In_13,In_169);
nand U482 (N_482,In_413,In_28);
and U483 (N_483,In_303,In_33);
nor U484 (N_484,In_403,In_117);
nor U485 (N_485,In_151,In_409);
xor U486 (N_486,In_153,In_448);
or U487 (N_487,In_248,In_4);
nand U488 (N_488,In_405,In_414);
nand U489 (N_489,In_376,In_347);
nand U490 (N_490,In_108,In_37);
xor U491 (N_491,In_360,In_18);
nand U492 (N_492,In_432,In_79);
nand U493 (N_493,In_78,In_234);
nand U494 (N_494,In_340,In_482);
and U495 (N_495,In_233,In_54);
and U496 (N_496,In_406,In_44);
or U497 (N_497,In_405,In_185);
and U498 (N_498,In_182,In_310);
and U499 (N_499,In_207,In_409);
nor U500 (N_500,In_281,In_340);
nand U501 (N_501,In_30,In_241);
nand U502 (N_502,In_33,In_107);
or U503 (N_503,In_389,In_134);
nor U504 (N_504,In_268,In_26);
nand U505 (N_505,In_405,In_319);
and U506 (N_506,In_367,In_275);
nor U507 (N_507,In_404,In_167);
nor U508 (N_508,In_222,In_223);
nand U509 (N_509,In_301,In_64);
nor U510 (N_510,In_14,In_32);
nand U511 (N_511,In_191,In_445);
and U512 (N_512,In_47,In_250);
or U513 (N_513,In_464,In_190);
or U514 (N_514,In_455,In_121);
or U515 (N_515,In_117,In_294);
nand U516 (N_516,In_199,In_308);
or U517 (N_517,In_229,In_74);
nand U518 (N_518,In_82,In_30);
or U519 (N_519,In_450,In_206);
nor U520 (N_520,In_153,In_256);
or U521 (N_521,In_399,In_421);
xnor U522 (N_522,In_191,In_175);
nand U523 (N_523,In_331,In_233);
nand U524 (N_524,In_190,In_385);
and U525 (N_525,In_96,In_22);
nor U526 (N_526,In_483,In_253);
and U527 (N_527,In_418,In_444);
or U528 (N_528,In_473,In_318);
and U529 (N_529,In_154,In_388);
and U530 (N_530,In_23,In_132);
nand U531 (N_531,In_409,In_211);
nor U532 (N_532,In_232,In_277);
or U533 (N_533,In_172,In_325);
or U534 (N_534,In_12,In_456);
and U535 (N_535,In_296,In_70);
nand U536 (N_536,In_455,In_174);
nand U537 (N_537,In_49,In_492);
nor U538 (N_538,In_18,In_432);
nor U539 (N_539,In_422,In_237);
and U540 (N_540,In_291,In_407);
nor U541 (N_541,In_158,In_122);
nand U542 (N_542,In_342,In_438);
nor U543 (N_543,In_184,In_104);
xnor U544 (N_544,In_161,In_143);
and U545 (N_545,In_116,In_461);
or U546 (N_546,In_155,In_162);
nand U547 (N_547,In_464,In_407);
nand U548 (N_548,In_247,In_488);
nor U549 (N_549,In_349,In_302);
nand U550 (N_550,In_223,In_18);
xor U551 (N_551,In_471,In_392);
xnor U552 (N_552,In_46,In_145);
and U553 (N_553,In_86,In_234);
nor U554 (N_554,In_275,In_234);
or U555 (N_555,In_82,In_289);
nand U556 (N_556,In_243,In_62);
and U557 (N_557,In_448,In_267);
nand U558 (N_558,In_425,In_195);
or U559 (N_559,In_387,In_420);
nand U560 (N_560,In_431,In_427);
xor U561 (N_561,In_209,In_248);
and U562 (N_562,In_112,In_369);
or U563 (N_563,In_408,In_397);
nand U564 (N_564,In_70,In_300);
and U565 (N_565,In_369,In_360);
and U566 (N_566,In_356,In_270);
and U567 (N_567,In_219,In_451);
and U568 (N_568,In_362,In_152);
xnor U569 (N_569,In_251,In_467);
or U570 (N_570,In_332,In_334);
and U571 (N_571,In_298,In_251);
or U572 (N_572,In_231,In_421);
nor U573 (N_573,In_307,In_205);
or U574 (N_574,In_395,In_376);
nor U575 (N_575,In_406,In_136);
and U576 (N_576,In_186,In_257);
nand U577 (N_577,In_309,In_246);
and U578 (N_578,In_495,In_35);
or U579 (N_579,In_418,In_387);
nand U580 (N_580,In_198,In_70);
nor U581 (N_581,In_337,In_416);
and U582 (N_582,In_484,In_448);
xnor U583 (N_583,In_15,In_274);
xor U584 (N_584,In_262,In_379);
nor U585 (N_585,In_394,In_20);
nand U586 (N_586,In_29,In_168);
xor U587 (N_587,In_4,In_280);
or U588 (N_588,In_312,In_267);
or U589 (N_589,In_241,In_342);
nand U590 (N_590,In_135,In_194);
nand U591 (N_591,In_378,In_420);
nand U592 (N_592,In_420,In_474);
nand U593 (N_593,In_301,In_236);
nor U594 (N_594,In_281,In_368);
nand U595 (N_595,In_109,In_54);
and U596 (N_596,In_247,In_75);
nand U597 (N_597,In_320,In_410);
nand U598 (N_598,In_297,In_124);
or U599 (N_599,In_217,In_450);
or U600 (N_600,In_399,In_68);
or U601 (N_601,In_110,In_351);
or U602 (N_602,In_103,In_57);
nand U603 (N_603,In_215,In_302);
nand U604 (N_604,In_148,In_268);
and U605 (N_605,In_184,In_126);
nor U606 (N_606,In_314,In_391);
nand U607 (N_607,In_296,In_438);
xnor U608 (N_608,In_37,In_354);
nor U609 (N_609,In_13,In_238);
nand U610 (N_610,In_27,In_364);
nor U611 (N_611,In_365,In_177);
nand U612 (N_612,In_409,In_304);
nand U613 (N_613,In_423,In_46);
or U614 (N_614,In_202,In_294);
or U615 (N_615,In_494,In_480);
and U616 (N_616,In_232,In_156);
xnor U617 (N_617,In_285,In_318);
and U618 (N_618,In_407,In_340);
or U619 (N_619,In_481,In_298);
and U620 (N_620,In_451,In_39);
xnor U621 (N_621,In_261,In_288);
nor U622 (N_622,In_467,In_232);
or U623 (N_623,In_247,In_159);
and U624 (N_624,In_75,In_415);
xor U625 (N_625,In_445,In_459);
and U626 (N_626,In_378,In_28);
nand U627 (N_627,In_279,In_392);
and U628 (N_628,In_187,In_360);
nand U629 (N_629,In_387,In_350);
and U630 (N_630,In_243,In_18);
or U631 (N_631,In_203,In_47);
and U632 (N_632,In_30,In_376);
and U633 (N_633,In_427,In_443);
or U634 (N_634,In_428,In_499);
xor U635 (N_635,In_110,In_83);
nor U636 (N_636,In_497,In_72);
nand U637 (N_637,In_277,In_367);
and U638 (N_638,In_448,In_428);
nand U639 (N_639,In_109,In_234);
xnor U640 (N_640,In_266,In_229);
and U641 (N_641,In_286,In_473);
or U642 (N_642,In_269,In_397);
nor U643 (N_643,In_364,In_235);
and U644 (N_644,In_471,In_298);
nand U645 (N_645,In_170,In_176);
or U646 (N_646,In_302,In_135);
or U647 (N_647,In_380,In_298);
and U648 (N_648,In_292,In_264);
nand U649 (N_649,In_311,In_72);
nor U650 (N_650,In_458,In_479);
nand U651 (N_651,In_136,In_278);
nand U652 (N_652,In_416,In_292);
and U653 (N_653,In_73,In_270);
nand U654 (N_654,In_89,In_33);
or U655 (N_655,In_455,In_127);
nor U656 (N_656,In_128,In_368);
nor U657 (N_657,In_127,In_226);
and U658 (N_658,In_255,In_31);
xor U659 (N_659,In_469,In_441);
nand U660 (N_660,In_256,In_493);
nand U661 (N_661,In_54,In_460);
xor U662 (N_662,In_221,In_113);
nand U663 (N_663,In_99,In_327);
and U664 (N_664,In_37,In_251);
or U665 (N_665,In_368,In_132);
nor U666 (N_666,In_198,In_59);
nor U667 (N_667,In_186,In_323);
nor U668 (N_668,In_145,In_209);
nand U669 (N_669,In_352,In_85);
or U670 (N_670,In_147,In_167);
nand U671 (N_671,In_437,In_116);
and U672 (N_672,In_28,In_45);
or U673 (N_673,In_21,In_78);
nand U674 (N_674,In_150,In_410);
and U675 (N_675,In_336,In_305);
and U676 (N_676,In_296,In_425);
or U677 (N_677,In_140,In_438);
nor U678 (N_678,In_149,In_404);
nand U679 (N_679,In_248,In_341);
nand U680 (N_680,In_25,In_273);
nand U681 (N_681,In_153,In_75);
or U682 (N_682,In_429,In_259);
nand U683 (N_683,In_406,In_413);
nand U684 (N_684,In_338,In_31);
or U685 (N_685,In_489,In_345);
nand U686 (N_686,In_58,In_3);
and U687 (N_687,In_229,In_277);
xor U688 (N_688,In_153,In_30);
and U689 (N_689,In_303,In_460);
nor U690 (N_690,In_251,In_384);
or U691 (N_691,In_392,In_469);
xor U692 (N_692,In_466,In_420);
nor U693 (N_693,In_273,In_222);
xnor U694 (N_694,In_175,In_444);
nand U695 (N_695,In_420,In_490);
or U696 (N_696,In_175,In_303);
or U697 (N_697,In_372,In_490);
nand U698 (N_698,In_142,In_312);
nand U699 (N_699,In_340,In_477);
and U700 (N_700,In_134,In_317);
xnor U701 (N_701,In_51,In_199);
or U702 (N_702,In_433,In_153);
or U703 (N_703,In_213,In_407);
and U704 (N_704,In_185,In_102);
xnor U705 (N_705,In_435,In_289);
nand U706 (N_706,In_56,In_482);
nor U707 (N_707,In_1,In_298);
or U708 (N_708,In_334,In_107);
nand U709 (N_709,In_106,In_216);
or U710 (N_710,In_312,In_302);
nand U711 (N_711,In_188,In_233);
xor U712 (N_712,In_268,In_152);
nor U713 (N_713,In_93,In_487);
or U714 (N_714,In_449,In_173);
nor U715 (N_715,In_47,In_479);
nor U716 (N_716,In_454,In_149);
or U717 (N_717,In_217,In_231);
and U718 (N_718,In_369,In_295);
nand U719 (N_719,In_81,In_142);
or U720 (N_720,In_91,In_344);
nor U721 (N_721,In_479,In_341);
or U722 (N_722,In_422,In_305);
nand U723 (N_723,In_317,In_403);
or U724 (N_724,In_364,In_489);
nor U725 (N_725,In_115,In_183);
nor U726 (N_726,In_259,In_168);
nor U727 (N_727,In_106,In_396);
and U728 (N_728,In_458,In_193);
or U729 (N_729,In_480,In_146);
and U730 (N_730,In_22,In_68);
and U731 (N_731,In_322,In_169);
xnor U732 (N_732,In_238,In_453);
nor U733 (N_733,In_110,In_485);
nor U734 (N_734,In_212,In_53);
or U735 (N_735,In_251,In_192);
nor U736 (N_736,In_218,In_105);
nand U737 (N_737,In_166,In_455);
nor U738 (N_738,In_281,In_165);
and U739 (N_739,In_366,In_315);
xnor U740 (N_740,In_120,In_6);
and U741 (N_741,In_144,In_152);
or U742 (N_742,In_348,In_163);
and U743 (N_743,In_107,In_86);
and U744 (N_744,In_223,In_298);
or U745 (N_745,In_226,In_389);
xor U746 (N_746,In_226,In_79);
nor U747 (N_747,In_372,In_487);
nand U748 (N_748,In_476,In_282);
nand U749 (N_749,In_50,In_14);
xor U750 (N_750,N_293,N_311);
nor U751 (N_751,N_229,N_384);
xnor U752 (N_752,N_647,N_385);
and U753 (N_753,N_193,N_678);
nand U754 (N_754,N_462,N_590);
or U755 (N_755,N_224,N_412);
nor U756 (N_756,N_52,N_68);
nand U757 (N_757,N_642,N_490);
or U758 (N_758,N_602,N_335);
and U759 (N_759,N_451,N_272);
or U760 (N_760,N_743,N_649);
and U761 (N_761,N_227,N_570);
xnor U762 (N_762,N_664,N_576);
or U763 (N_763,N_436,N_102);
nand U764 (N_764,N_230,N_547);
nor U765 (N_765,N_411,N_13);
nand U766 (N_766,N_500,N_8);
nor U767 (N_767,N_392,N_729);
xor U768 (N_768,N_378,N_679);
and U769 (N_769,N_205,N_103);
or U770 (N_770,N_315,N_34);
and U771 (N_771,N_528,N_79);
nand U772 (N_772,N_17,N_261);
nand U773 (N_773,N_707,N_388);
nor U774 (N_774,N_269,N_353);
and U775 (N_775,N_159,N_208);
xor U776 (N_776,N_23,N_415);
nand U777 (N_777,N_66,N_609);
xnor U778 (N_778,N_288,N_397);
nor U779 (N_779,N_80,N_483);
and U780 (N_780,N_413,N_94);
or U781 (N_781,N_667,N_100);
xnor U782 (N_782,N_135,N_403);
and U783 (N_783,N_401,N_694);
nand U784 (N_784,N_455,N_142);
nor U785 (N_785,N_185,N_457);
or U786 (N_786,N_742,N_471);
nand U787 (N_787,N_111,N_359);
nand U788 (N_788,N_463,N_303);
nor U789 (N_789,N_119,N_190);
nand U790 (N_790,N_705,N_92);
and U791 (N_791,N_43,N_70);
or U792 (N_792,N_644,N_599);
and U793 (N_793,N_48,N_81);
nor U794 (N_794,N_108,N_16);
and U795 (N_795,N_728,N_697);
nor U796 (N_796,N_402,N_452);
xor U797 (N_797,N_726,N_691);
nor U798 (N_798,N_254,N_265);
and U799 (N_799,N_320,N_394);
xor U800 (N_800,N_188,N_178);
nand U801 (N_801,N_489,N_689);
xor U802 (N_802,N_561,N_733);
and U803 (N_803,N_721,N_617);
nor U804 (N_804,N_64,N_423);
xnor U805 (N_805,N_350,N_600);
nor U806 (N_806,N_481,N_550);
or U807 (N_807,N_520,N_136);
or U808 (N_808,N_720,N_372);
or U809 (N_809,N_511,N_274);
nand U810 (N_810,N_255,N_611);
or U811 (N_811,N_184,N_400);
nand U812 (N_812,N_104,N_560);
xor U813 (N_813,N_719,N_492);
nand U814 (N_814,N_321,N_643);
or U815 (N_815,N_316,N_168);
and U816 (N_816,N_331,N_740);
or U817 (N_817,N_165,N_715);
or U818 (N_818,N_630,N_307);
and U819 (N_819,N_131,N_432);
and U820 (N_820,N_129,N_137);
and U821 (N_821,N_695,N_1);
xnor U822 (N_822,N_526,N_292);
nor U823 (N_823,N_552,N_505);
xnor U824 (N_824,N_333,N_238);
nand U825 (N_825,N_579,N_183);
and U826 (N_826,N_544,N_239);
or U827 (N_827,N_660,N_584);
nand U828 (N_828,N_606,N_26);
nor U829 (N_829,N_540,N_515);
nor U830 (N_830,N_109,N_503);
and U831 (N_831,N_712,N_280);
xor U832 (N_832,N_748,N_132);
xnor U833 (N_833,N_460,N_220);
nand U834 (N_834,N_424,N_557);
or U835 (N_835,N_674,N_539);
nor U836 (N_836,N_210,N_594);
and U837 (N_837,N_442,N_198);
or U838 (N_838,N_619,N_203);
nand U839 (N_839,N_266,N_395);
nor U840 (N_840,N_628,N_430);
xnor U841 (N_841,N_744,N_551);
or U842 (N_842,N_655,N_284);
and U843 (N_843,N_398,N_591);
nand U844 (N_844,N_535,N_153);
and U845 (N_845,N_305,N_233);
or U846 (N_846,N_676,N_124);
nor U847 (N_847,N_568,N_745);
nand U848 (N_848,N_449,N_169);
xor U849 (N_849,N_310,N_348);
and U850 (N_850,N_533,N_36);
or U851 (N_851,N_141,N_248);
nor U852 (N_852,N_259,N_240);
and U853 (N_853,N_469,N_126);
xor U854 (N_854,N_672,N_732);
nand U855 (N_855,N_312,N_339);
and U856 (N_856,N_681,N_562);
xor U857 (N_857,N_330,N_597);
nand U858 (N_858,N_456,N_61);
and U859 (N_859,N_308,N_171);
nor U860 (N_860,N_429,N_632);
or U861 (N_861,N_656,N_604);
nor U862 (N_862,N_167,N_29);
or U863 (N_863,N_731,N_680);
nor U864 (N_864,N_166,N_84);
nand U865 (N_865,N_635,N_379);
or U866 (N_866,N_730,N_696);
xor U867 (N_867,N_236,N_358);
nor U868 (N_868,N_298,N_536);
nand U869 (N_869,N_214,N_121);
nand U870 (N_870,N_363,N_377);
xnor U871 (N_871,N_105,N_501);
and U872 (N_872,N_174,N_725);
or U873 (N_873,N_326,N_603);
nand U874 (N_874,N_72,N_18);
nand U875 (N_875,N_309,N_273);
and U876 (N_876,N_291,N_736);
nor U877 (N_877,N_651,N_675);
xor U878 (N_878,N_120,N_625);
nor U879 (N_879,N_313,N_595);
and U880 (N_880,N_427,N_654);
nor U881 (N_881,N_145,N_749);
or U882 (N_882,N_716,N_685);
or U883 (N_883,N_260,N_624);
nand U884 (N_884,N_147,N_74);
and U885 (N_885,N_69,N_148);
nor U886 (N_886,N_56,N_421);
or U887 (N_887,N_30,N_516);
and U888 (N_888,N_256,N_627);
and U889 (N_889,N_473,N_297);
xor U890 (N_890,N_199,N_47);
xnor U891 (N_891,N_612,N_531);
nand U892 (N_892,N_349,N_19);
and U893 (N_893,N_53,N_549);
nor U894 (N_894,N_207,N_62);
nor U895 (N_895,N_294,N_314);
xor U896 (N_896,N_407,N_419);
nor U897 (N_897,N_519,N_268);
or U898 (N_898,N_390,N_14);
nand U899 (N_899,N_328,N_659);
or U900 (N_900,N_182,N_65);
nor U901 (N_901,N_77,N_107);
nor U902 (N_902,N_197,N_671);
nand U903 (N_903,N_614,N_155);
xor U904 (N_904,N_468,N_196);
nor U905 (N_905,N_657,N_698);
or U906 (N_906,N_461,N_202);
nor U907 (N_907,N_342,N_276);
nor U908 (N_908,N_343,N_559);
xor U909 (N_909,N_262,N_152);
nand U910 (N_910,N_445,N_371);
nand U911 (N_911,N_24,N_626);
nor U912 (N_912,N_453,N_33);
or U913 (N_913,N_299,N_82);
nor U914 (N_914,N_409,N_217);
or U915 (N_915,N_682,N_118);
nor U916 (N_916,N_458,N_391);
and U917 (N_917,N_556,N_42);
or U918 (N_918,N_88,N_623);
or U919 (N_919,N_399,N_252);
or U920 (N_920,N_485,N_253);
nand U921 (N_921,N_338,N_63);
or U922 (N_922,N_277,N_502);
and U923 (N_923,N_57,N_668);
or U924 (N_924,N_706,N_573);
nand U925 (N_925,N_480,N_718);
xnor U926 (N_926,N_521,N_582);
or U927 (N_927,N_375,N_574);
and U928 (N_928,N_356,N_156);
nand U929 (N_929,N_631,N_55);
or U930 (N_930,N_571,N_662);
nor U931 (N_931,N_364,N_543);
and U932 (N_932,N_99,N_416);
nor U933 (N_933,N_381,N_361);
nor U934 (N_934,N_714,N_76);
nor U935 (N_935,N_86,N_435);
xnor U936 (N_936,N_404,N_447);
nor U937 (N_937,N_475,N_496);
nor U938 (N_938,N_257,N_440);
xor U939 (N_939,N_620,N_96);
and U940 (N_940,N_189,N_40);
or U941 (N_941,N_666,N_529);
xnor U942 (N_942,N_180,N_243);
nand U943 (N_943,N_739,N_146);
nor U944 (N_944,N_438,N_20);
and U945 (N_945,N_304,N_444);
or U946 (N_946,N_704,N_425);
or U947 (N_947,N_191,N_722);
nand U948 (N_948,N_530,N_78);
or U949 (N_949,N_125,N_652);
or U950 (N_950,N_201,N_665);
or U951 (N_951,N_6,N_162);
nand U952 (N_952,N_368,N_21);
nor U953 (N_953,N_106,N_302);
and U954 (N_954,N_246,N_212);
and U955 (N_955,N_653,N_172);
and U956 (N_956,N_282,N_692);
xnor U957 (N_957,N_441,N_548);
or U958 (N_958,N_270,N_592);
xnor U959 (N_959,N_241,N_279);
and U960 (N_960,N_554,N_645);
xnor U961 (N_961,N_219,N_7);
and U962 (N_962,N_211,N_585);
nor U963 (N_963,N_357,N_488);
nor U964 (N_964,N_746,N_245);
nand U965 (N_965,N_420,N_223);
nor U966 (N_966,N_60,N_232);
and U967 (N_967,N_735,N_130);
and U968 (N_968,N_231,N_487);
nand U969 (N_969,N_408,N_344);
nand U970 (N_970,N_498,N_341);
nand U971 (N_971,N_59,N_115);
nand U972 (N_972,N_90,N_161);
or U973 (N_973,N_360,N_688);
nand U974 (N_974,N_170,N_534);
nor U975 (N_975,N_386,N_366);
or U976 (N_976,N_39,N_417);
or U977 (N_977,N_89,N_354);
and U978 (N_978,N_484,N_323);
nor U979 (N_979,N_608,N_470);
and U980 (N_980,N_177,N_464);
and U981 (N_981,N_509,N_50);
nor U982 (N_982,N_658,N_708);
nor U983 (N_983,N_514,N_143);
or U984 (N_984,N_340,N_127);
or U985 (N_985,N_389,N_482);
nand U986 (N_986,N_45,N_113);
or U987 (N_987,N_151,N_337);
xor U988 (N_988,N_618,N_433);
nand U989 (N_989,N_422,N_640);
and U990 (N_990,N_446,N_286);
xnor U991 (N_991,N_122,N_636);
xor U992 (N_992,N_334,N_163);
nand U993 (N_993,N_186,N_51);
nor U994 (N_994,N_512,N_87);
and U995 (N_995,N_431,N_478);
nor U996 (N_996,N_593,N_44);
nand U997 (N_997,N_418,N_596);
and U998 (N_998,N_493,N_306);
nand U999 (N_999,N_414,N_319);
or U1000 (N_1000,N_9,N_370);
nor U1001 (N_1001,N_459,N_324);
or U1002 (N_1002,N_558,N_247);
or U1003 (N_1003,N_517,N_518);
or U1004 (N_1004,N_641,N_467);
or U1005 (N_1005,N_222,N_234);
nand U1006 (N_1006,N_267,N_513);
nor U1007 (N_1007,N_383,N_607);
and U1008 (N_1008,N_290,N_474);
nand U1009 (N_1009,N_285,N_465);
or U1010 (N_1010,N_322,N_187);
nor U1011 (N_1011,N_154,N_580);
nor U1012 (N_1012,N_225,N_724);
nor U1013 (N_1013,N_633,N_95);
or U1014 (N_1014,N_157,N_541);
or U1015 (N_1015,N_495,N_713);
nand U1016 (N_1016,N_295,N_522);
nand U1017 (N_1017,N_110,N_242);
or U1018 (N_1018,N_701,N_58);
or U1019 (N_1019,N_406,N_387);
nor U1020 (N_1020,N_486,N_615);
nor U1021 (N_1021,N_140,N_439);
nor U1022 (N_1022,N_454,N_537);
nor U1023 (N_1023,N_71,N_637);
nand U1024 (N_1024,N_598,N_737);
nand U1025 (N_1025,N_546,N_215);
nor U1026 (N_1026,N_553,N_97);
nand U1027 (N_1027,N_287,N_160);
nand U1028 (N_1028,N_5,N_67);
nor U1029 (N_1029,N_35,N_49);
or U1030 (N_1030,N_634,N_200);
and U1031 (N_1031,N_437,N_532);
nand U1032 (N_1032,N_525,N_15);
nand U1033 (N_1033,N_426,N_639);
and U1034 (N_1034,N_179,N_382);
and U1035 (N_1035,N_206,N_249);
xor U1036 (N_1036,N_98,N_327);
and U1037 (N_1037,N_101,N_271);
or U1038 (N_1038,N_347,N_376);
nand U1039 (N_1039,N_144,N_527);
nand U1040 (N_1040,N_373,N_158);
nor U1041 (N_1041,N_466,N_613);
nor U1042 (N_1042,N_134,N_648);
nor U1043 (N_1043,N_747,N_351);
and U1044 (N_1044,N_75,N_22);
and U1045 (N_1045,N_283,N_27);
nand U1046 (N_1046,N_683,N_173);
nor U1047 (N_1047,N_710,N_494);
nor U1048 (N_1048,N_116,N_621);
nand U1049 (N_1049,N_128,N_538);
or U1050 (N_1050,N_524,N_684);
or U1051 (N_1051,N_428,N_669);
nor U1052 (N_1052,N_362,N_3);
xnor U1053 (N_1053,N_727,N_703);
xor U1054 (N_1054,N_542,N_507);
or U1055 (N_1055,N_216,N_650);
nor U1056 (N_1056,N_476,N_213);
nand U1057 (N_1057,N_38,N_450);
or U1058 (N_1058,N_393,N_175);
nor U1059 (N_1059,N_587,N_195);
nor U1060 (N_1060,N_563,N_497);
nand U1061 (N_1061,N_616,N_690);
or U1062 (N_1062,N_567,N_629);
nor U1063 (N_1063,N_581,N_263);
xnor U1064 (N_1064,N_702,N_37);
and U1065 (N_1065,N_741,N_583);
or U1066 (N_1066,N_588,N_85);
and U1067 (N_1067,N_4,N_443);
nor U1068 (N_1068,N_499,N_289);
nor U1069 (N_1069,N_296,N_605);
nand U1070 (N_1070,N_192,N_565);
or U1071 (N_1071,N_275,N_10);
nand U1072 (N_1072,N_194,N_380);
and U1073 (N_1073,N_687,N_396);
or U1074 (N_1074,N_138,N_164);
and U1075 (N_1075,N_12,N_93);
and U1076 (N_1076,N_209,N_700);
or U1077 (N_1077,N_638,N_46);
or U1078 (N_1078,N_734,N_278);
nor U1079 (N_1079,N_365,N_575);
nor U1080 (N_1080,N_244,N_300);
or U1081 (N_1081,N_410,N_369);
nand U1082 (N_1082,N_250,N_73);
or U1083 (N_1083,N_610,N_723);
nand U1084 (N_1084,N_235,N_504);
and U1085 (N_1085,N_114,N_83);
and U1086 (N_1086,N_355,N_555);
nand U1087 (N_1087,N_693,N_738);
nand U1088 (N_1088,N_523,N_301);
or U1089 (N_1089,N_545,N_352);
nor U1090 (N_1090,N_264,N_2);
nor U1091 (N_1091,N_601,N_336);
xnor U1092 (N_1092,N_569,N_673);
or U1093 (N_1093,N_345,N_510);
and U1094 (N_1094,N_472,N_677);
nor U1095 (N_1095,N_0,N_41);
nor U1096 (N_1096,N_367,N_228);
or U1097 (N_1097,N_506,N_204);
nand U1098 (N_1098,N_281,N_32);
xnor U1099 (N_1099,N_586,N_572);
nand U1100 (N_1100,N_578,N_717);
and U1101 (N_1101,N_670,N_329);
nor U1102 (N_1102,N_25,N_54);
xor U1103 (N_1103,N_218,N_491);
nor U1104 (N_1104,N_226,N_434);
or U1105 (N_1105,N_133,N_686);
nor U1106 (N_1106,N_150,N_139);
nor U1107 (N_1107,N_28,N_237);
or U1108 (N_1108,N_566,N_91);
nand U1109 (N_1109,N_332,N_589);
nand U1110 (N_1110,N_112,N_508);
and U1111 (N_1111,N_448,N_699);
or U1112 (N_1112,N_149,N_123);
and U1113 (N_1113,N_622,N_318);
or U1114 (N_1114,N_479,N_251);
or U1115 (N_1115,N_374,N_564);
nor U1116 (N_1116,N_317,N_577);
nand U1117 (N_1117,N_181,N_711);
nor U1118 (N_1118,N_11,N_31);
nor U1119 (N_1119,N_176,N_221);
or U1120 (N_1120,N_258,N_405);
and U1121 (N_1121,N_709,N_477);
nand U1122 (N_1122,N_325,N_346);
and U1123 (N_1123,N_663,N_117);
nor U1124 (N_1124,N_661,N_646);
nor U1125 (N_1125,N_90,N_670);
nand U1126 (N_1126,N_316,N_663);
and U1127 (N_1127,N_399,N_262);
and U1128 (N_1128,N_567,N_257);
or U1129 (N_1129,N_99,N_31);
nor U1130 (N_1130,N_396,N_298);
or U1131 (N_1131,N_130,N_414);
or U1132 (N_1132,N_747,N_642);
or U1133 (N_1133,N_731,N_59);
or U1134 (N_1134,N_638,N_271);
and U1135 (N_1135,N_395,N_194);
or U1136 (N_1136,N_642,N_138);
nand U1137 (N_1137,N_176,N_148);
xnor U1138 (N_1138,N_9,N_674);
or U1139 (N_1139,N_656,N_687);
and U1140 (N_1140,N_687,N_464);
nand U1141 (N_1141,N_666,N_114);
nand U1142 (N_1142,N_273,N_140);
or U1143 (N_1143,N_403,N_239);
nor U1144 (N_1144,N_577,N_447);
and U1145 (N_1145,N_217,N_107);
and U1146 (N_1146,N_580,N_337);
and U1147 (N_1147,N_661,N_93);
and U1148 (N_1148,N_650,N_189);
nand U1149 (N_1149,N_118,N_227);
and U1150 (N_1150,N_662,N_504);
and U1151 (N_1151,N_608,N_61);
or U1152 (N_1152,N_710,N_489);
nand U1153 (N_1153,N_278,N_516);
xnor U1154 (N_1154,N_17,N_486);
nand U1155 (N_1155,N_40,N_454);
or U1156 (N_1156,N_170,N_208);
nor U1157 (N_1157,N_343,N_21);
and U1158 (N_1158,N_222,N_718);
and U1159 (N_1159,N_658,N_110);
or U1160 (N_1160,N_708,N_729);
nor U1161 (N_1161,N_62,N_100);
nand U1162 (N_1162,N_582,N_184);
nor U1163 (N_1163,N_373,N_647);
nor U1164 (N_1164,N_17,N_134);
or U1165 (N_1165,N_359,N_477);
and U1166 (N_1166,N_473,N_31);
and U1167 (N_1167,N_614,N_411);
or U1168 (N_1168,N_20,N_362);
and U1169 (N_1169,N_254,N_700);
and U1170 (N_1170,N_558,N_519);
nand U1171 (N_1171,N_40,N_463);
nand U1172 (N_1172,N_694,N_238);
and U1173 (N_1173,N_486,N_205);
nor U1174 (N_1174,N_115,N_310);
or U1175 (N_1175,N_38,N_289);
xnor U1176 (N_1176,N_373,N_438);
and U1177 (N_1177,N_630,N_509);
and U1178 (N_1178,N_45,N_645);
or U1179 (N_1179,N_728,N_66);
and U1180 (N_1180,N_68,N_119);
nor U1181 (N_1181,N_475,N_60);
or U1182 (N_1182,N_478,N_239);
nor U1183 (N_1183,N_419,N_123);
and U1184 (N_1184,N_612,N_445);
or U1185 (N_1185,N_290,N_395);
or U1186 (N_1186,N_429,N_15);
nand U1187 (N_1187,N_652,N_710);
and U1188 (N_1188,N_68,N_490);
and U1189 (N_1189,N_81,N_65);
nor U1190 (N_1190,N_565,N_453);
or U1191 (N_1191,N_41,N_603);
nand U1192 (N_1192,N_376,N_415);
or U1193 (N_1193,N_646,N_113);
nor U1194 (N_1194,N_215,N_237);
nand U1195 (N_1195,N_730,N_390);
nor U1196 (N_1196,N_538,N_508);
nand U1197 (N_1197,N_718,N_299);
xnor U1198 (N_1198,N_154,N_748);
nor U1199 (N_1199,N_525,N_641);
or U1200 (N_1200,N_417,N_403);
nor U1201 (N_1201,N_378,N_137);
nand U1202 (N_1202,N_430,N_515);
or U1203 (N_1203,N_409,N_307);
and U1204 (N_1204,N_293,N_415);
and U1205 (N_1205,N_258,N_328);
or U1206 (N_1206,N_539,N_744);
nand U1207 (N_1207,N_268,N_253);
nand U1208 (N_1208,N_743,N_151);
xnor U1209 (N_1209,N_698,N_230);
and U1210 (N_1210,N_377,N_706);
nor U1211 (N_1211,N_640,N_313);
or U1212 (N_1212,N_340,N_504);
and U1213 (N_1213,N_499,N_18);
or U1214 (N_1214,N_496,N_276);
nor U1215 (N_1215,N_678,N_277);
and U1216 (N_1216,N_584,N_404);
nor U1217 (N_1217,N_407,N_665);
nand U1218 (N_1218,N_306,N_131);
nand U1219 (N_1219,N_499,N_461);
xor U1220 (N_1220,N_725,N_31);
nor U1221 (N_1221,N_229,N_302);
nand U1222 (N_1222,N_96,N_70);
and U1223 (N_1223,N_378,N_406);
and U1224 (N_1224,N_489,N_284);
or U1225 (N_1225,N_707,N_736);
or U1226 (N_1226,N_390,N_217);
nor U1227 (N_1227,N_415,N_380);
nor U1228 (N_1228,N_593,N_728);
nand U1229 (N_1229,N_526,N_713);
nor U1230 (N_1230,N_464,N_457);
or U1231 (N_1231,N_127,N_133);
or U1232 (N_1232,N_438,N_201);
nand U1233 (N_1233,N_320,N_32);
xor U1234 (N_1234,N_241,N_421);
nor U1235 (N_1235,N_397,N_149);
nand U1236 (N_1236,N_690,N_396);
xnor U1237 (N_1237,N_26,N_621);
nand U1238 (N_1238,N_105,N_351);
nor U1239 (N_1239,N_588,N_140);
or U1240 (N_1240,N_630,N_532);
and U1241 (N_1241,N_571,N_315);
and U1242 (N_1242,N_272,N_112);
xor U1243 (N_1243,N_526,N_74);
and U1244 (N_1244,N_205,N_4);
nand U1245 (N_1245,N_332,N_139);
or U1246 (N_1246,N_140,N_584);
and U1247 (N_1247,N_609,N_38);
and U1248 (N_1248,N_331,N_227);
and U1249 (N_1249,N_372,N_156);
or U1250 (N_1250,N_175,N_662);
xor U1251 (N_1251,N_94,N_197);
and U1252 (N_1252,N_211,N_481);
or U1253 (N_1253,N_115,N_261);
nand U1254 (N_1254,N_114,N_180);
and U1255 (N_1255,N_10,N_94);
or U1256 (N_1256,N_556,N_737);
and U1257 (N_1257,N_100,N_181);
and U1258 (N_1258,N_168,N_253);
xor U1259 (N_1259,N_383,N_43);
or U1260 (N_1260,N_215,N_727);
nor U1261 (N_1261,N_742,N_223);
nand U1262 (N_1262,N_379,N_473);
nand U1263 (N_1263,N_1,N_228);
and U1264 (N_1264,N_485,N_341);
nor U1265 (N_1265,N_169,N_106);
or U1266 (N_1266,N_696,N_260);
nor U1267 (N_1267,N_227,N_620);
nor U1268 (N_1268,N_445,N_561);
or U1269 (N_1269,N_617,N_180);
nor U1270 (N_1270,N_119,N_322);
nand U1271 (N_1271,N_4,N_727);
or U1272 (N_1272,N_461,N_407);
or U1273 (N_1273,N_83,N_633);
nand U1274 (N_1274,N_188,N_535);
nor U1275 (N_1275,N_246,N_262);
nand U1276 (N_1276,N_203,N_128);
or U1277 (N_1277,N_681,N_186);
and U1278 (N_1278,N_31,N_50);
or U1279 (N_1279,N_706,N_198);
nand U1280 (N_1280,N_89,N_665);
nor U1281 (N_1281,N_125,N_334);
or U1282 (N_1282,N_526,N_299);
nor U1283 (N_1283,N_107,N_194);
xnor U1284 (N_1284,N_242,N_306);
xnor U1285 (N_1285,N_266,N_333);
xor U1286 (N_1286,N_618,N_276);
nor U1287 (N_1287,N_68,N_279);
and U1288 (N_1288,N_696,N_373);
nand U1289 (N_1289,N_349,N_51);
and U1290 (N_1290,N_630,N_135);
nor U1291 (N_1291,N_115,N_388);
xnor U1292 (N_1292,N_421,N_184);
nand U1293 (N_1293,N_62,N_428);
nor U1294 (N_1294,N_657,N_720);
nor U1295 (N_1295,N_275,N_329);
nand U1296 (N_1296,N_92,N_470);
xnor U1297 (N_1297,N_6,N_513);
or U1298 (N_1298,N_270,N_16);
nor U1299 (N_1299,N_421,N_687);
or U1300 (N_1300,N_579,N_722);
nand U1301 (N_1301,N_408,N_6);
nand U1302 (N_1302,N_738,N_540);
xnor U1303 (N_1303,N_679,N_167);
and U1304 (N_1304,N_665,N_279);
nand U1305 (N_1305,N_130,N_151);
xnor U1306 (N_1306,N_53,N_510);
nor U1307 (N_1307,N_279,N_144);
xnor U1308 (N_1308,N_561,N_222);
or U1309 (N_1309,N_278,N_346);
nor U1310 (N_1310,N_500,N_349);
xor U1311 (N_1311,N_639,N_608);
nor U1312 (N_1312,N_259,N_192);
or U1313 (N_1313,N_143,N_306);
nand U1314 (N_1314,N_424,N_330);
xor U1315 (N_1315,N_509,N_463);
and U1316 (N_1316,N_451,N_20);
and U1317 (N_1317,N_437,N_434);
or U1318 (N_1318,N_160,N_230);
nand U1319 (N_1319,N_267,N_492);
and U1320 (N_1320,N_168,N_38);
or U1321 (N_1321,N_165,N_375);
and U1322 (N_1322,N_247,N_722);
xnor U1323 (N_1323,N_289,N_533);
nor U1324 (N_1324,N_529,N_38);
and U1325 (N_1325,N_63,N_188);
nor U1326 (N_1326,N_103,N_109);
nor U1327 (N_1327,N_262,N_510);
and U1328 (N_1328,N_264,N_702);
and U1329 (N_1329,N_468,N_41);
or U1330 (N_1330,N_710,N_669);
nand U1331 (N_1331,N_669,N_94);
nor U1332 (N_1332,N_91,N_681);
nand U1333 (N_1333,N_679,N_375);
nor U1334 (N_1334,N_612,N_304);
or U1335 (N_1335,N_0,N_189);
xor U1336 (N_1336,N_128,N_652);
nor U1337 (N_1337,N_599,N_371);
nand U1338 (N_1338,N_573,N_616);
or U1339 (N_1339,N_716,N_323);
nand U1340 (N_1340,N_422,N_636);
nand U1341 (N_1341,N_88,N_168);
xnor U1342 (N_1342,N_177,N_62);
or U1343 (N_1343,N_745,N_293);
and U1344 (N_1344,N_706,N_733);
and U1345 (N_1345,N_689,N_165);
xor U1346 (N_1346,N_282,N_44);
and U1347 (N_1347,N_299,N_502);
nand U1348 (N_1348,N_114,N_497);
nor U1349 (N_1349,N_125,N_581);
and U1350 (N_1350,N_534,N_77);
nand U1351 (N_1351,N_359,N_562);
xnor U1352 (N_1352,N_572,N_268);
nor U1353 (N_1353,N_733,N_361);
or U1354 (N_1354,N_238,N_424);
or U1355 (N_1355,N_677,N_483);
nand U1356 (N_1356,N_89,N_449);
xnor U1357 (N_1357,N_96,N_700);
and U1358 (N_1358,N_336,N_352);
xnor U1359 (N_1359,N_26,N_397);
or U1360 (N_1360,N_364,N_456);
or U1361 (N_1361,N_378,N_613);
nor U1362 (N_1362,N_293,N_299);
and U1363 (N_1363,N_482,N_466);
nand U1364 (N_1364,N_292,N_442);
nand U1365 (N_1365,N_257,N_701);
nand U1366 (N_1366,N_707,N_425);
and U1367 (N_1367,N_396,N_619);
xnor U1368 (N_1368,N_749,N_552);
nor U1369 (N_1369,N_337,N_70);
or U1370 (N_1370,N_89,N_339);
and U1371 (N_1371,N_467,N_173);
nand U1372 (N_1372,N_469,N_648);
nand U1373 (N_1373,N_489,N_628);
or U1374 (N_1374,N_415,N_189);
or U1375 (N_1375,N_50,N_325);
and U1376 (N_1376,N_51,N_489);
nand U1377 (N_1377,N_719,N_223);
nand U1378 (N_1378,N_158,N_71);
xor U1379 (N_1379,N_59,N_745);
nor U1380 (N_1380,N_268,N_429);
and U1381 (N_1381,N_21,N_506);
or U1382 (N_1382,N_567,N_643);
or U1383 (N_1383,N_478,N_74);
nand U1384 (N_1384,N_119,N_702);
nor U1385 (N_1385,N_555,N_435);
xor U1386 (N_1386,N_320,N_48);
and U1387 (N_1387,N_247,N_643);
nand U1388 (N_1388,N_576,N_226);
and U1389 (N_1389,N_94,N_618);
xor U1390 (N_1390,N_557,N_170);
nor U1391 (N_1391,N_295,N_239);
nor U1392 (N_1392,N_418,N_622);
and U1393 (N_1393,N_444,N_513);
nand U1394 (N_1394,N_724,N_75);
and U1395 (N_1395,N_348,N_240);
xnor U1396 (N_1396,N_88,N_174);
nand U1397 (N_1397,N_569,N_502);
or U1398 (N_1398,N_352,N_668);
nor U1399 (N_1399,N_196,N_397);
nor U1400 (N_1400,N_484,N_338);
and U1401 (N_1401,N_225,N_20);
and U1402 (N_1402,N_518,N_701);
and U1403 (N_1403,N_520,N_649);
and U1404 (N_1404,N_150,N_73);
and U1405 (N_1405,N_94,N_31);
or U1406 (N_1406,N_453,N_408);
nor U1407 (N_1407,N_194,N_394);
nor U1408 (N_1408,N_288,N_335);
or U1409 (N_1409,N_535,N_696);
nor U1410 (N_1410,N_719,N_100);
nand U1411 (N_1411,N_705,N_553);
and U1412 (N_1412,N_443,N_310);
nor U1413 (N_1413,N_630,N_339);
nor U1414 (N_1414,N_553,N_315);
xnor U1415 (N_1415,N_588,N_340);
or U1416 (N_1416,N_595,N_613);
nor U1417 (N_1417,N_23,N_82);
nand U1418 (N_1418,N_640,N_619);
and U1419 (N_1419,N_743,N_45);
or U1420 (N_1420,N_319,N_651);
and U1421 (N_1421,N_89,N_326);
or U1422 (N_1422,N_536,N_420);
nand U1423 (N_1423,N_664,N_202);
nor U1424 (N_1424,N_356,N_658);
nand U1425 (N_1425,N_643,N_516);
or U1426 (N_1426,N_359,N_141);
and U1427 (N_1427,N_0,N_162);
nor U1428 (N_1428,N_204,N_544);
nor U1429 (N_1429,N_23,N_407);
nor U1430 (N_1430,N_290,N_721);
nand U1431 (N_1431,N_265,N_609);
xor U1432 (N_1432,N_139,N_42);
nor U1433 (N_1433,N_135,N_575);
or U1434 (N_1434,N_290,N_201);
or U1435 (N_1435,N_316,N_343);
nor U1436 (N_1436,N_388,N_9);
nand U1437 (N_1437,N_151,N_196);
nor U1438 (N_1438,N_437,N_94);
or U1439 (N_1439,N_151,N_311);
xnor U1440 (N_1440,N_233,N_604);
nand U1441 (N_1441,N_231,N_97);
or U1442 (N_1442,N_432,N_560);
nand U1443 (N_1443,N_113,N_139);
or U1444 (N_1444,N_278,N_277);
and U1445 (N_1445,N_724,N_169);
nor U1446 (N_1446,N_445,N_58);
and U1447 (N_1447,N_600,N_88);
nand U1448 (N_1448,N_82,N_326);
or U1449 (N_1449,N_167,N_374);
nor U1450 (N_1450,N_390,N_148);
and U1451 (N_1451,N_539,N_701);
nor U1452 (N_1452,N_51,N_749);
xnor U1453 (N_1453,N_381,N_504);
nor U1454 (N_1454,N_575,N_61);
nor U1455 (N_1455,N_84,N_278);
nand U1456 (N_1456,N_17,N_597);
or U1457 (N_1457,N_413,N_523);
and U1458 (N_1458,N_452,N_251);
nand U1459 (N_1459,N_301,N_284);
or U1460 (N_1460,N_749,N_457);
or U1461 (N_1461,N_254,N_546);
or U1462 (N_1462,N_524,N_121);
or U1463 (N_1463,N_206,N_670);
or U1464 (N_1464,N_417,N_152);
xnor U1465 (N_1465,N_327,N_742);
nor U1466 (N_1466,N_466,N_574);
or U1467 (N_1467,N_353,N_404);
or U1468 (N_1468,N_706,N_499);
nand U1469 (N_1469,N_592,N_736);
nand U1470 (N_1470,N_451,N_368);
nand U1471 (N_1471,N_735,N_182);
nor U1472 (N_1472,N_458,N_171);
xnor U1473 (N_1473,N_472,N_31);
xnor U1474 (N_1474,N_582,N_489);
and U1475 (N_1475,N_493,N_298);
nor U1476 (N_1476,N_299,N_542);
nor U1477 (N_1477,N_732,N_440);
nand U1478 (N_1478,N_377,N_178);
nand U1479 (N_1479,N_515,N_391);
and U1480 (N_1480,N_346,N_260);
nor U1481 (N_1481,N_172,N_391);
and U1482 (N_1482,N_676,N_655);
or U1483 (N_1483,N_506,N_731);
and U1484 (N_1484,N_83,N_317);
nor U1485 (N_1485,N_329,N_162);
and U1486 (N_1486,N_389,N_457);
or U1487 (N_1487,N_104,N_131);
nor U1488 (N_1488,N_588,N_103);
nor U1489 (N_1489,N_311,N_17);
nand U1490 (N_1490,N_41,N_324);
nand U1491 (N_1491,N_614,N_149);
xor U1492 (N_1492,N_593,N_173);
nor U1493 (N_1493,N_339,N_561);
or U1494 (N_1494,N_156,N_126);
nor U1495 (N_1495,N_577,N_124);
nand U1496 (N_1496,N_90,N_97);
nand U1497 (N_1497,N_389,N_260);
and U1498 (N_1498,N_320,N_528);
or U1499 (N_1499,N_33,N_158);
or U1500 (N_1500,N_1447,N_886);
nand U1501 (N_1501,N_1271,N_1422);
nand U1502 (N_1502,N_1419,N_888);
and U1503 (N_1503,N_802,N_1106);
or U1504 (N_1504,N_843,N_1269);
nor U1505 (N_1505,N_1311,N_1037);
and U1506 (N_1506,N_1125,N_815);
or U1507 (N_1507,N_1265,N_999);
nor U1508 (N_1508,N_1117,N_924);
nor U1509 (N_1509,N_1052,N_1029);
or U1510 (N_1510,N_1483,N_1245);
nand U1511 (N_1511,N_1266,N_1172);
nand U1512 (N_1512,N_1174,N_1352);
xor U1513 (N_1513,N_1219,N_1489);
nor U1514 (N_1514,N_989,N_1345);
xor U1515 (N_1515,N_1319,N_1458);
and U1516 (N_1516,N_1148,N_1147);
xor U1517 (N_1517,N_1050,N_1010);
nand U1518 (N_1518,N_1003,N_962);
nor U1519 (N_1519,N_1018,N_1334);
nor U1520 (N_1520,N_1014,N_1104);
nor U1521 (N_1521,N_1390,N_1044);
or U1522 (N_1522,N_1385,N_1263);
and U1523 (N_1523,N_1330,N_1142);
and U1524 (N_1524,N_1434,N_852);
nand U1525 (N_1525,N_1120,N_1133);
nor U1526 (N_1526,N_1316,N_1252);
and U1527 (N_1527,N_1471,N_804);
and U1528 (N_1528,N_1135,N_1368);
nor U1529 (N_1529,N_1308,N_1425);
nand U1530 (N_1530,N_1179,N_1303);
or U1531 (N_1531,N_801,N_1166);
and U1532 (N_1532,N_1098,N_1077);
nand U1533 (N_1533,N_903,N_862);
and U1534 (N_1534,N_1378,N_1175);
nand U1535 (N_1535,N_1307,N_1342);
and U1536 (N_1536,N_1242,N_978);
or U1537 (N_1537,N_1047,N_952);
nand U1538 (N_1538,N_1470,N_1468);
nand U1539 (N_1539,N_1270,N_1123);
or U1540 (N_1540,N_1113,N_977);
or U1541 (N_1541,N_775,N_797);
xnor U1542 (N_1542,N_1144,N_1016);
or U1543 (N_1543,N_915,N_1430);
and U1544 (N_1544,N_1177,N_885);
xnor U1545 (N_1545,N_1203,N_1152);
nand U1546 (N_1546,N_1035,N_1296);
xnor U1547 (N_1547,N_943,N_1350);
nor U1548 (N_1548,N_1209,N_773);
nor U1549 (N_1549,N_840,N_803);
or U1550 (N_1550,N_846,N_1153);
or U1551 (N_1551,N_997,N_1409);
nor U1552 (N_1552,N_1401,N_1344);
and U1553 (N_1553,N_941,N_1078);
xnor U1554 (N_1554,N_1085,N_1051);
nand U1555 (N_1555,N_776,N_1402);
nand U1556 (N_1556,N_1143,N_889);
or U1557 (N_1557,N_1075,N_1318);
and U1558 (N_1558,N_1414,N_1107);
and U1559 (N_1559,N_1495,N_1032);
or U1560 (N_1560,N_818,N_875);
nor U1561 (N_1561,N_829,N_764);
and U1562 (N_1562,N_931,N_1155);
and U1563 (N_1563,N_1017,N_851);
and U1564 (N_1564,N_819,N_1176);
and U1565 (N_1565,N_934,N_1235);
nor U1566 (N_1566,N_1217,N_1365);
nor U1567 (N_1567,N_994,N_1432);
or U1568 (N_1568,N_792,N_1025);
and U1569 (N_1569,N_1127,N_1273);
and U1570 (N_1570,N_1171,N_1188);
nand U1571 (N_1571,N_849,N_1317);
or U1572 (N_1572,N_1060,N_778);
xor U1573 (N_1573,N_1313,N_1126);
xnor U1574 (N_1574,N_779,N_1222);
or U1575 (N_1575,N_1041,N_867);
xnor U1576 (N_1576,N_1215,N_905);
or U1577 (N_1577,N_1103,N_1185);
and U1578 (N_1578,N_1040,N_824);
nor U1579 (N_1579,N_900,N_1285);
and U1580 (N_1580,N_1329,N_1099);
and U1581 (N_1581,N_898,N_789);
and U1582 (N_1582,N_1408,N_1165);
nor U1583 (N_1583,N_935,N_1393);
and U1584 (N_1584,N_1225,N_1221);
or U1585 (N_1585,N_766,N_1136);
xnor U1586 (N_1586,N_1472,N_1312);
or U1587 (N_1587,N_1302,N_1255);
nor U1588 (N_1588,N_998,N_1054);
xnor U1589 (N_1589,N_854,N_927);
nor U1590 (N_1590,N_1413,N_970);
and U1591 (N_1591,N_1065,N_1223);
nor U1592 (N_1592,N_1190,N_1068);
and U1593 (N_1593,N_1213,N_884);
or U1594 (N_1594,N_993,N_930);
xnor U1595 (N_1595,N_1056,N_765);
xnor U1596 (N_1596,N_1473,N_908);
or U1597 (N_1597,N_967,N_1005);
nor U1598 (N_1598,N_1100,N_1454);
and U1599 (N_1599,N_1151,N_781);
nand U1600 (N_1600,N_1465,N_842);
nor U1601 (N_1601,N_1397,N_876);
nand U1602 (N_1602,N_1305,N_932);
nand U1603 (N_1603,N_874,N_1241);
or U1604 (N_1604,N_939,N_1064);
nand U1605 (N_1605,N_1469,N_1337);
and U1606 (N_1606,N_853,N_986);
and U1607 (N_1607,N_1247,N_784);
or U1608 (N_1608,N_1448,N_1452);
and U1609 (N_1609,N_957,N_1341);
nor U1610 (N_1610,N_1356,N_1294);
nand U1611 (N_1611,N_928,N_1450);
or U1612 (N_1612,N_1431,N_1343);
nor U1613 (N_1613,N_827,N_968);
or U1614 (N_1614,N_1243,N_1012);
or U1615 (N_1615,N_950,N_1109);
nor U1616 (N_1616,N_793,N_750);
and U1617 (N_1617,N_923,N_1238);
nand U1618 (N_1618,N_1030,N_969);
xor U1619 (N_1619,N_988,N_1083);
nand U1620 (N_1620,N_1272,N_991);
or U1621 (N_1621,N_1295,N_1298);
nand U1622 (N_1622,N_1320,N_1205);
nand U1623 (N_1623,N_1150,N_921);
nor U1624 (N_1624,N_944,N_1115);
or U1625 (N_1625,N_1498,N_1467);
and U1626 (N_1626,N_1421,N_1453);
xor U1627 (N_1627,N_1353,N_1405);
nand U1628 (N_1628,N_1499,N_795);
or U1629 (N_1629,N_1476,N_906);
and U1630 (N_1630,N_878,N_1346);
xor U1631 (N_1631,N_1081,N_963);
nand U1632 (N_1632,N_1191,N_883);
nand U1633 (N_1633,N_831,N_787);
nor U1634 (N_1634,N_1207,N_810);
nand U1635 (N_1635,N_925,N_1493);
nand U1636 (N_1636,N_1158,N_1211);
and U1637 (N_1637,N_1377,N_1360);
nor U1638 (N_1638,N_856,N_806);
xnor U1639 (N_1639,N_1091,N_1310);
nand U1640 (N_1640,N_1057,N_1363);
and U1641 (N_1641,N_1460,N_1210);
nor U1642 (N_1642,N_1290,N_1403);
and U1643 (N_1643,N_951,N_1199);
or U1644 (N_1644,N_1097,N_1333);
nand U1645 (N_1645,N_860,N_893);
or U1646 (N_1646,N_1116,N_1024);
xor U1647 (N_1647,N_913,N_861);
and U1648 (N_1648,N_1328,N_1324);
nand U1649 (N_1649,N_823,N_847);
nand U1650 (N_1650,N_1336,N_850);
or U1651 (N_1651,N_1201,N_942);
or U1652 (N_1652,N_1464,N_1134);
nor U1653 (N_1653,N_1260,N_752);
nor U1654 (N_1654,N_1299,N_1101);
xnor U1655 (N_1655,N_791,N_1229);
nor U1656 (N_1656,N_1224,N_907);
nand U1657 (N_1657,N_899,N_1406);
nand U1658 (N_1658,N_919,N_1218);
and U1659 (N_1659,N_1011,N_839);
and U1660 (N_1660,N_1121,N_1423);
nor U1661 (N_1661,N_1375,N_1236);
or U1662 (N_1662,N_1325,N_1386);
nor U1663 (N_1663,N_917,N_1384);
nor U1664 (N_1664,N_814,N_1293);
nor U1665 (N_1665,N_1045,N_1082);
nand U1666 (N_1666,N_1481,N_1321);
nand U1667 (N_1667,N_1239,N_983);
nand U1668 (N_1668,N_1438,N_774);
or U1669 (N_1669,N_1372,N_794);
nand U1670 (N_1670,N_933,N_1261);
xnor U1671 (N_1671,N_1262,N_961);
and U1672 (N_1672,N_1062,N_835);
or U1673 (N_1673,N_1396,N_868);
and U1674 (N_1674,N_870,N_1132);
nand U1675 (N_1675,N_1327,N_1186);
nand U1676 (N_1676,N_1391,N_1373);
or U1677 (N_1677,N_966,N_1442);
nor U1678 (N_1678,N_1049,N_1366);
nand U1679 (N_1679,N_858,N_1036);
or U1680 (N_1680,N_1072,N_1146);
xnor U1681 (N_1681,N_1208,N_1102);
or U1682 (N_1682,N_965,N_1231);
nand U1683 (N_1683,N_845,N_1335);
and U1684 (N_1684,N_1233,N_882);
nor U1685 (N_1685,N_808,N_1286);
nand U1686 (N_1686,N_947,N_1392);
nand U1687 (N_1687,N_880,N_902);
nor U1688 (N_1688,N_1169,N_1485);
nor U1689 (N_1689,N_1069,N_1444);
or U1690 (N_1690,N_890,N_1292);
nor U1691 (N_1691,N_754,N_1178);
nor U1692 (N_1692,N_822,N_767);
xnor U1693 (N_1693,N_1118,N_976);
or U1694 (N_1694,N_1264,N_1394);
nand U1695 (N_1695,N_1461,N_1008);
or U1696 (N_1696,N_1031,N_959);
or U1697 (N_1697,N_1163,N_1456);
xor U1698 (N_1698,N_1063,N_1309);
and U1699 (N_1699,N_984,N_1487);
nand U1700 (N_1700,N_1331,N_960);
or U1701 (N_1701,N_1415,N_865);
nand U1702 (N_1702,N_937,N_1355);
and U1703 (N_1703,N_1110,N_1258);
or U1704 (N_1704,N_1240,N_830);
nand U1705 (N_1705,N_1080,N_1111);
xnor U1706 (N_1706,N_1256,N_1193);
or U1707 (N_1707,N_914,N_1380);
nor U1708 (N_1708,N_1259,N_1093);
nand U1709 (N_1709,N_1251,N_1043);
nand U1710 (N_1710,N_879,N_1070);
and U1711 (N_1711,N_1197,N_1055);
nor U1712 (N_1712,N_762,N_1283);
nor U1713 (N_1713,N_1234,N_922);
nand U1714 (N_1714,N_1257,N_1092);
and U1715 (N_1715,N_1149,N_1089);
and U1716 (N_1716,N_1039,N_1216);
or U1717 (N_1717,N_866,N_1297);
or U1718 (N_1718,N_1195,N_1323);
nor U1719 (N_1719,N_1347,N_897);
and U1720 (N_1720,N_832,N_751);
or U1721 (N_1721,N_1230,N_1268);
xor U1722 (N_1722,N_864,N_1426);
and U1723 (N_1723,N_756,N_1364);
or U1724 (N_1724,N_1340,N_760);
and U1725 (N_1725,N_758,N_1002);
xor U1726 (N_1726,N_1379,N_1357);
nand U1727 (N_1727,N_1404,N_946);
or U1728 (N_1728,N_1488,N_1486);
and U1729 (N_1729,N_1427,N_974);
and U1730 (N_1730,N_833,N_1276);
and U1731 (N_1731,N_1395,N_1466);
and U1732 (N_1732,N_901,N_1094);
nor U1733 (N_1733,N_958,N_1192);
nor U1734 (N_1734,N_1492,N_1189);
and U1735 (N_1735,N_945,N_1145);
nor U1736 (N_1736,N_1420,N_1028);
nand U1737 (N_1737,N_1059,N_1367);
and U1738 (N_1738,N_1168,N_836);
nor U1739 (N_1739,N_799,N_1315);
or U1740 (N_1740,N_1105,N_848);
xnor U1741 (N_1741,N_1019,N_929);
nor U1742 (N_1742,N_926,N_1141);
nand U1743 (N_1743,N_1226,N_895);
or U1744 (N_1744,N_1455,N_1249);
xor U1745 (N_1745,N_1369,N_1440);
and U1746 (N_1746,N_1084,N_1156);
nand U1747 (N_1747,N_872,N_788);
nor U1748 (N_1748,N_972,N_1314);
nor U1749 (N_1749,N_1370,N_1023);
nor U1750 (N_1750,N_1214,N_837);
or U1751 (N_1751,N_1164,N_785);
or U1752 (N_1752,N_825,N_1009);
or U1753 (N_1753,N_1338,N_1412);
nand U1754 (N_1754,N_1246,N_1277);
or U1755 (N_1755,N_1291,N_1076);
nor U1756 (N_1756,N_777,N_987);
or U1757 (N_1757,N_1306,N_1322);
nand U1758 (N_1758,N_910,N_857);
and U1759 (N_1759,N_1358,N_1300);
nor U1760 (N_1760,N_1048,N_1074);
or U1761 (N_1761,N_1279,N_1387);
or U1762 (N_1762,N_1004,N_783);
nor U1763 (N_1763,N_1228,N_891);
and U1764 (N_1764,N_1253,N_755);
nor U1765 (N_1765,N_1095,N_855);
nand U1766 (N_1766,N_1274,N_1477);
or U1767 (N_1767,N_771,N_800);
nand U1768 (N_1768,N_770,N_757);
nand U1769 (N_1769,N_1326,N_1359);
and U1770 (N_1770,N_1006,N_1496);
and U1771 (N_1771,N_1275,N_1184);
nor U1772 (N_1772,N_816,N_1204);
and U1773 (N_1773,N_1437,N_1167);
xor U1774 (N_1774,N_1162,N_1067);
or U1775 (N_1775,N_1027,N_1200);
or U1776 (N_1776,N_820,N_782);
and U1777 (N_1777,N_1399,N_769);
nor U1778 (N_1778,N_1139,N_918);
xor U1779 (N_1779,N_1436,N_1459);
or U1780 (N_1780,N_1042,N_1157);
and U1781 (N_1781,N_995,N_1022);
nand U1782 (N_1782,N_1173,N_909);
xnor U1783 (N_1783,N_887,N_1119);
and U1784 (N_1784,N_826,N_768);
nand U1785 (N_1785,N_1382,N_1281);
and U1786 (N_1786,N_1278,N_1383);
nand U1787 (N_1787,N_1071,N_949);
nand U1788 (N_1788,N_982,N_1180);
or U1789 (N_1789,N_1348,N_894);
and U1790 (N_1790,N_956,N_1108);
nand U1791 (N_1791,N_912,N_821);
or U1792 (N_1792,N_844,N_841);
and U1793 (N_1793,N_1497,N_955);
or U1794 (N_1794,N_892,N_1474);
or U1795 (N_1795,N_1411,N_1140);
nor U1796 (N_1796,N_1131,N_1090);
nand U1797 (N_1797,N_1087,N_1088);
and U1798 (N_1798,N_1232,N_904);
and U1799 (N_1799,N_1058,N_1374);
and U1800 (N_1800,N_916,N_1398);
or U1801 (N_1801,N_1137,N_1237);
nand U1802 (N_1802,N_1194,N_1202);
and U1803 (N_1803,N_1301,N_1066);
and U1804 (N_1804,N_1288,N_1417);
and U1805 (N_1805,N_1410,N_807);
nor U1806 (N_1806,N_761,N_964);
nor U1807 (N_1807,N_1114,N_975);
or U1808 (N_1808,N_1001,N_1248);
nand U1809 (N_1809,N_1428,N_1122);
nor U1810 (N_1810,N_1013,N_973);
nor U1811 (N_1811,N_1159,N_971);
xnor U1812 (N_1812,N_938,N_1282);
nor U1813 (N_1813,N_786,N_1284);
or U1814 (N_1814,N_1361,N_772);
nand U1815 (N_1815,N_1212,N_1021);
nand U1816 (N_1816,N_1443,N_948);
xnor U1817 (N_1817,N_979,N_1124);
or U1818 (N_1818,N_1441,N_1433);
or U1819 (N_1819,N_985,N_1462);
nand U1820 (N_1820,N_1416,N_1250);
nand U1821 (N_1821,N_811,N_859);
nor U1822 (N_1822,N_1254,N_863);
nand U1823 (N_1823,N_812,N_1244);
nor U1824 (N_1824,N_953,N_1429);
xnor U1825 (N_1825,N_1388,N_1187);
or U1826 (N_1826,N_1160,N_763);
nand U1827 (N_1827,N_1478,N_981);
or U1828 (N_1828,N_1480,N_1073);
nor U1829 (N_1829,N_805,N_834);
or U1830 (N_1830,N_759,N_881);
or U1831 (N_1831,N_1332,N_1439);
nor U1832 (N_1832,N_1445,N_1381);
nor U1833 (N_1833,N_817,N_1015);
xor U1834 (N_1834,N_1007,N_1198);
or U1835 (N_1835,N_1479,N_869);
or U1836 (N_1836,N_1086,N_813);
and U1837 (N_1837,N_1463,N_790);
and U1838 (N_1838,N_798,N_1475);
and U1839 (N_1839,N_1138,N_809);
or U1840 (N_1840,N_1289,N_871);
nor U1841 (N_1841,N_1181,N_1304);
xor U1842 (N_1842,N_1339,N_1457);
or U1843 (N_1843,N_1435,N_1206);
nor U1844 (N_1844,N_1154,N_1183);
nand U1845 (N_1845,N_1096,N_1484);
and U1846 (N_1846,N_1400,N_873);
nand U1847 (N_1847,N_1161,N_828);
nand U1848 (N_1848,N_954,N_1449);
nand U1849 (N_1849,N_936,N_838);
nand U1850 (N_1850,N_1280,N_1128);
and U1851 (N_1851,N_1220,N_1491);
xor U1852 (N_1852,N_1227,N_1407);
or U1853 (N_1853,N_1034,N_1020);
xor U1854 (N_1854,N_877,N_1079);
or U1855 (N_1855,N_1038,N_1362);
nand U1856 (N_1856,N_1196,N_1371);
and U1857 (N_1857,N_1170,N_980);
xor U1858 (N_1858,N_1267,N_990);
nor U1859 (N_1859,N_1354,N_1130);
or U1860 (N_1860,N_940,N_1446);
or U1861 (N_1861,N_1424,N_1026);
nor U1862 (N_1862,N_896,N_911);
or U1863 (N_1863,N_1389,N_753);
or U1864 (N_1864,N_1376,N_1351);
or U1865 (N_1865,N_1112,N_1061);
nor U1866 (N_1866,N_920,N_1482);
nand U1867 (N_1867,N_1490,N_992);
nand U1868 (N_1868,N_1418,N_1046);
nand U1869 (N_1869,N_1053,N_1033);
and U1870 (N_1870,N_1129,N_1349);
nand U1871 (N_1871,N_796,N_996);
nand U1872 (N_1872,N_1287,N_780);
xor U1873 (N_1873,N_1182,N_1451);
nor U1874 (N_1874,N_1494,N_1000);
nor U1875 (N_1875,N_1084,N_1110);
nor U1876 (N_1876,N_1091,N_1064);
or U1877 (N_1877,N_1264,N_1047);
or U1878 (N_1878,N_1475,N_1102);
and U1879 (N_1879,N_1306,N_957);
and U1880 (N_1880,N_1414,N_1317);
nand U1881 (N_1881,N_997,N_896);
and U1882 (N_1882,N_764,N_1167);
xnor U1883 (N_1883,N_1134,N_809);
nand U1884 (N_1884,N_905,N_1332);
nand U1885 (N_1885,N_1361,N_1298);
nand U1886 (N_1886,N_969,N_1241);
xnor U1887 (N_1887,N_1420,N_839);
nand U1888 (N_1888,N_1248,N_980);
nand U1889 (N_1889,N_809,N_1249);
xnor U1890 (N_1890,N_921,N_887);
and U1891 (N_1891,N_1268,N_1260);
xor U1892 (N_1892,N_923,N_1430);
or U1893 (N_1893,N_759,N_1407);
nor U1894 (N_1894,N_1335,N_1214);
xnor U1895 (N_1895,N_849,N_841);
nor U1896 (N_1896,N_838,N_1361);
nor U1897 (N_1897,N_1288,N_1187);
xor U1898 (N_1898,N_1312,N_1476);
nand U1899 (N_1899,N_838,N_1081);
nor U1900 (N_1900,N_909,N_774);
and U1901 (N_1901,N_1079,N_1451);
and U1902 (N_1902,N_1235,N_993);
nor U1903 (N_1903,N_1245,N_774);
or U1904 (N_1904,N_1124,N_1278);
nor U1905 (N_1905,N_1223,N_830);
and U1906 (N_1906,N_846,N_1142);
and U1907 (N_1907,N_1401,N_1172);
nand U1908 (N_1908,N_1159,N_1154);
and U1909 (N_1909,N_964,N_842);
nand U1910 (N_1910,N_1011,N_1484);
nor U1911 (N_1911,N_1051,N_1020);
nor U1912 (N_1912,N_930,N_951);
nor U1913 (N_1913,N_1489,N_1060);
or U1914 (N_1914,N_876,N_1065);
nand U1915 (N_1915,N_1152,N_863);
or U1916 (N_1916,N_780,N_1034);
nor U1917 (N_1917,N_919,N_1089);
nor U1918 (N_1918,N_1272,N_935);
nor U1919 (N_1919,N_815,N_845);
nor U1920 (N_1920,N_1141,N_1398);
xnor U1921 (N_1921,N_1257,N_1182);
nand U1922 (N_1922,N_1009,N_1364);
nor U1923 (N_1923,N_1103,N_1320);
nand U1924 (N_1924,N_775,N_1076);
or U1925 (N_1925,N_816,N_1135);
nor U1926 (N_1926,N_1398,N_1442);
nand U1927 (N_1927,N_1262,N_1421);
nor U1928 (N_1928,N_1075,N_1444);
nor U1929 (N_1929,N_1401,N_1115);
and U1930 (N_1930,N_814,N_1176);
or U1931 (N_1931,N_976,N_1193);
xnor U1932 (N_1932,N_881,N_1441);
nand U1933 (N_1933,N_872,N_938);
or U1934 (N_1934,N_1095,N_1138);
nand U1935 (N_1935,N_1297,N_1131);
nand U1936 (N_1936,N_820,N_1122);
nand U1937 (N_1937,N_872,N_1201);
and U1938 (N_1938,N_1274,N_852);
nor U1939 (N_1939,N_1183,N_1165);
and U1940 (N_1940,N_842,N_1013);
and U1941 (N_1941,N_1142,N_1148);
nor U1942 (N_1942,N_1284,N_1439);
nor U1943 (N_1943,N_955,N_1478);
xor U1944 (N_1944,N_1172,N_1175);
nand U1945 (N_1945,N_922,N_1388);
nand U1946 (N_1946,N_922,N_1387);
and U1947 (N_1947,N_1441,N_1092);
nor U1948 (N_1948,N_1215,N_1018);
nand U1949 (N_1949,N_1435,N_1377);
nand U1950 (N_1950,N_1037,N_1127);
and U1951 (N_1951,N_1381,N_1268);
or U1952 (N_1952,N_1419,N_897);
or U1953 (N_1953,N_796,N_907);
nor U1954 (N_1954,N_1364,N_1422);
nor U1955 (N_1955,N_921,N_1291);
nand U1956 (N_1956,N_1199,N_1102);
or U1957 (N_1957,N_989,N_1065);
nor U1958 (N_1958,N_1086,N_803);
or U1959 (N_1959,N_1064,N_1486);
and U1960 (N_1960,N_1265,N_954);
or U1961 (N_1961,N_755,N_1148);
and U1962 (N_1962,N_958,N_1153);
nand U1963 (N_1963,N_1101,N_1498);
or U1964 (N_1964,N_1318,N_982);
and U1965 (N_1965,N_1373,N_1225);
nand U1966 (N_1966,N_786,N_1152);
xnor U1967 (N_1967,N_786,N_813);
nor U1968 (N_1968,N_783,N_1116);
or U1969 (N_1969,N_1347,N_1193);
xor U1970 (N_1970,N_966,N_1017);
nor U1971 (N_1971,N_1045,N_798);
nor U1972 (N_1972,N_1209,N_1238);
and U1973 (N_1973,N_829,N_982);
xor U1974 (N_1974,N_758,N_1110);
nand U1975 (N_1975,N_1343,N_1467);
or U1976 (N_1976,N_962,N_949);
nor U1977 (N_1977,N_898,N_1131);
xnor U1978 (N_1978,N_1296,N_998);
nor U1979 (N_1979,N_830,N_934);
nor U1980 (N_1980,N_1232,N_1474);
nand U1981 (N_1981,N_1166,N_797);
or U1982 (N_1982,N_1396,N_984);
nor U1983 (N_1983,N_1039,N_1128);
nor U1984 (N_1984,N_914,N_1373);
nand U1985 (N_1985,N_1374,N_1462);
xor U1986 (N_1986,N_865,N_1243);
xor U1987 (N_1987,N_861,N_767);
xor U1988 (N_1988,N_1012,N_1281);
xor U1989 (N_1989,N_1194,N_1106);
xnor U1990 (N_1990,N_805,N_755);
nand U1991 (N_1991,N_1104,N_1452);
nand U1992 (N_1992,N_1210,N_778);
or U1993 (N_1993,N_1227,N_884);
or U1994 (N_1994,N_984,N_1263);
nor U1995 (N_1995,N_922,N_1056);
xnor U1996 (N_1996,N_1391,N_1314);
and U1997 (N_1997,N_1258,N_952);
nand U1998 (N_1998,N_1028,N_1158);
nor U1999 (N_1999,N_812,N_754);
or U2000 (N_2000,N_1314,N_1320);
nand U2001 (N_2001,N_1257,N_1161);
and U2002 (N_2002,N_1101,N_993);
nand U2003 (N_2003,N_982,N_1077);
or U2004 (N_2004,N_1149,N_1175);
or U2005 (N_2005,N_1429,N_1092);
nor U2006 (N_2006,N_998,N_1493);
nand U2007 (N_2007,N_1443,N_799);
nand U2008 (N_2008,N_1128,N_1481);
and U2009 (N_2009,N_1138,N_1026);
nand U2010 (N_2010,N_1023,N_1047);
xor U2011 (N_2011,N_1197,N_1211);
or U2012 (N_2012,N_1141,N_1405);
xnor U2013 (N_2013,N_1040,N_851);
nand U2014 (N_2014,N_1158,N_937);
nor U2015 (N_2015,N_1204,N_781);
or U2016 (N_2016,N_975,N_1475);
or U2017 (N_2017,N_1372,N_1179);
nand U2018 (N_2018,N_860,N_1124);
or U2019 (N_2019,N_1055,N_1313);
nor U2020 (N_2020,N_1437,N_1230);
and U2021 (N_2021,N_1462,N_1311);
and U2022 (N_2022,N_1462,N_1274);
or U2023 (N_2023,N_1104,N_1127);
or U2024 (N_2024,N_846,N_1235);
nand U2025 (N_2025,N_1469,N_1209);
or U2026 (N_2026,N_1018,N_1370);
and U2027 (N_2027,N_1153,N_1430);
nor U2028 (N_2028,N_1072,N_1214);
nor U2029 (N_2029,N_1157,N_1291);
nor U2030 (N_2030,N_1198,N_853);
xnor U2031 (N_2031,N_760,N_1391);
nand U2032 (N_2032,N_1184,N_1085);
and U2033 (N_2033,N_785,N_1233);
nand U2034 (N_2034,N_933,N_1232);
or U2035 (N_2035,N_1452,N_1279);
and U2036 (N_2036,N_978,N_1475);
nor U2037 (N_2037,N_815,N_1472);
nor U2038 (N_2038,N_751,N_835);
nand U2039 (N_2039,N_765,N_816);
xnor U2040 (N_2040,N_1200,N_1398);
nand U2041 (N_2041,N_1248,N_763);
and U2042 (N_2042,N_1032,N_887);
xnor U2043 (N_2043,N_1203,N_1364);
nor U2044 (N_2044,N_1432,N_1079);
and U2045 (N_2045,N_1155,N_841);
and U2046 (N_2046,N_1215,N_1371);
or U2047 (N_2047,N_1491,N_922);
nand U2048 (N_2048,N_1408,N_1292);
nand U2049 (N_2049,N_1257,N_1179);
and U2050 (N_2050,N_1100,N_1469);
and U2051 (N_2051,N_772,N_1153);
and U2052 (N_2052,N_1151,N_1485);
or U2053 (N_2053,N_1280,N_1003);
nand U2054 (N_2054,N_820,N_1325);
and U2055 (N_2055,N_1201,N_1084);
nand U2056 (N_2056,N_1084,N_1285);
nor U2057 (N_2057,N_1223,N_1434);
nor U2058 (N_2058,N_1473,N_1258);
nand U2059 (N_2059,N_819,N_796);
xor U2060 (N_2060,N_1084,N_902);
and U2061 (N_2061,N_1359,N_1170);
and U2062 (N_2062,N_1030,N_978);
and U2063 (N_2063,N_1292,N_988);
nor U2064 (N_2064,N_926,N_899);
nand U2065 (N_2065,N_1044,N_1133);
nand U2066 (N_2066,N_1329,N_994);
nand U2067 (N_2067,N_1177,N_1017);
nand U2068 (N_2068,N_1045,N_1403);
and U2069 (N_2069,N_838,N_862);
and U2070 (N_2070,N_1436,N_1316);
and U2071 (N_2071,N_1465,N_946);
or U2072 (N_2072,N_871,N_1245);
and U2073 (N_2073,N_1083,N_1120);
nor U2074 (N_2074,N_772,N_1379);
and U2075 (N_2075,N_1161,N_1354);
xor U2076 (N_2076,N_1164,N_1156);
or U2077 (N_2077,N_879,N_1382);
or U2078 (N_2078,N_1176,N_1419);
nand U2079 (N_2079,N_945,N_1081);
or U2080 (N_2080,N_1067,N_1420);
nor U2081 (N_2081,N_1496,N_1131);
nand U2082 (N_2082,N_1255,N_1361);
and U2083 (N_2083,N_780,N_1111);
xor U2084 (N_2084,N_884,N_1008);
nor U2085 (N_2085,N_1250,N_1186);
and U2086 (N_2086,N_1096,N_1480);
nand U2087 (N_2087,N_1108,N_927);
xnor U2088 (N_2088,N_1469,N_995);
or U2089 (N_2089,N_1206,N_1337);
nor U2090 (N_2090,N_1223,N_1494);
nor U2091 (N_2091,N_1051,N_1412);
and U2092 (N_2092,N_875,N_1017);
nor U2093 (N_2093,N_837,N_1263);
and U2094 (N_2094,N_1360,N_929);
or U2095 (N_2095,N_1481,N_867);
nand U2096 (N_2096,N_1096,N_1080);
nor U2097 (N_2097,N_1447,N_1084);
and U2098 (N_2098,N_1084,N_858);
or U2099 (N_2099,N_1088,N_1333);
nor U2100 (N_2100,N_1395,N_1187);
or U2101 (N_2101,N_1105,N_796);
xor U2102 (N_2102,N_798,N_1190);
nor U2103 (N_2103,N_1431,N_1488);
or U2104 (N_2104,N_1019,N_852);
nor U2105 (N_2105,N_1273,N_1019);
nand U2106 (N_2106,N_761,N_1124);
nand U2107 (N_2107,N_1347,N_1327);
and U2108 (N_2108,N_1436,N_1245);
and U2109 (N_2109,N_1349,N_957);
and U2110 (N_2110,N_1173,N_1319);
and U2111 (N_2111,N_1372,N_766);
xor U2112 (N_2112,N_1071,N_1110);
nand U2113 (N_2113,N_1204,N_1148);
or U2114 (N_2114,N_990,N_952);
and U2115 (N_2115,N_812,N_1140);
and U2116 (N_2116,N_1056,N_1107);
nand U2117 (N_2117,N_867,N_1369);
and U2118 (N_2118,N_1355,N_1349);
nand U2119 (N_2119,N_1210,N_1461);
nor U2120 (N_2120,N_1033,N_1181);
and U2121 (N_2121,N_1444,N_1479);
xnor U2122 (N_2122,N_808,N_1082);
nor U2123 (N_2123,N_1271,N_1021);
nor U2124 (N_2124,N_1401,N_1236);
nor U2125 (N_2125,N_1249,N_805);
or U2126 (N_2126,N_1468,N_838);
and U2127 (N_2127,N_1331,N_1087);
xnor U2128 (N_2128,N_795,N_763);
or U2129 (N_2129,N_900,N_1139);
nand U2130 (N_2130,N_1031,N_800);
and U2131 (N_2131,N_1419,N_847);
or U2132 (N_2132,N_852,N_1497);
and U2133 (N_2133,N_1408,N_1064);
nor U2134 (N_2134,N_1409,N_1186);
nand U2135 (N_2135,N_1195,N_1032);
nand U2136 (N_2136,N_1350,N_1004);
nand U2137 (N_2137,N_1206,N_1457);
or U2138 (N_2138,N_1411,N_832);
xnor U2139 (N_2139,N_1291,N_1229);
xnor U2140 (N_2140,N_780,N_1123);
and U2141 (N_2141,N_961,N_941);
nor U2142 (N_2142,N_1185,N_970);
or U2143 (N_2143,N_1318,N_918);
nor U2144 (N_2144,N_763,N_1086);
nor U2145 (N_2145,N_1123,N_1260);
nor U2146 (N_2146,N_1059,N_1215);
and U2147 (N_2147,N_1262,N_993);
or U2148 (N_2148,N_791,N_1149);
nand U2149 (N_2149,N_1436,N_1040);
nand U2150 (N_2150,N_1321,N_1221);
xnor U2151 (N_2151,N_1328,N_1496);
xor U2152 (N_2152,N_888,N_1174);
or U2153 (N_2153,N_1280,N_817);
xnor U2154 (N_2154,N_1379,N_962);
or U2155 (N_2155,N_1393,N_1310);
and U2156 (N_2156,N_1224,N_1067);
nor U2157 (N_2157,N_1427,N_1174);
nand U2158 (N_2158,N_1163,N_1110);
and U2159 (N_2159,N_1353,N_818);
or U2160 (N_2160,N_1244,N_905);
nor U2161 (N_2161,N_1085,N_1394);
nor U2162 (N_2162,N_811,N_1463);
nor U2163 (N_2163,N_1349,N_816);
and U2164 (N_2164,N_929,N_1192);
xor U2165 (N_2165,N_1486,N_1179);
or U2166 (N_2166,N_1446,N_1330);
nand U2167 (N_2167,N_765,N_761);
nand U2168 (N_2168,N_1101,N_928);
nor U2169 (N_2169,N_777,N_1355);
nand U2170 (N_2170,N_1471,N_1158);
xor U2171 (N_2171,N_1133,N_835);
and U2172 (N_2172,N_1490,N_1056);
nor U2173 (N_2173,N_890,N_1232);
or U2174 (N_2174,N_1129,N_1242);
or U2175 (N_2175,N_1412,N_1011);
and U2176 (N_2176,N_1393,N_1131);
nor U2177 (N_2177,N_1155,N_1088);
nor U2178 (N_2178,N_802,N_1413);
nor U2179 (N_2179,N_1245,N_1457);
nor U2180 (N_2180,N_953,N_1428);
or U2181 (N_2181,N_1095,N_1387);
and U2182 (N_2182,N_965,N_1450);
nor U2183 (N_2183,N_1130,N_958);
xnor U2184 (N_2184,N_831,N_1401);
nor U2185 (N_2185,N_1214,N_935);
and U2186 (N_2186,N_1049,N_1115);
xor U2187 (N_2187,N_878,N_973);
nor U2188 (N_2188,N_1134,N_1400);
xor U2189 (N_2189,N_946,N_1436);
xor U2190 (N_2190,N_1127,N_759);
nand U2191 (N_2191,N_889,N_1228);
nor U2192 (N_2192,N_1052,N_832);
nand U2193 (N_2193,N_968,N_964);
nand U2194 (N_2194,N_1312,N_1401);
or U2195 (N_2195,N_1185,N_757);
and U2196 (N_2196,N_1282,N_926);
or U2197 (N_2197,N_790,N_1411);
or U2198 (N_2198,N_1175,N_1376);
nand U2199 (N_2199,N_1488,N_1447);
nand U2200 (N_2200,N_1422,N_1295);
nand U2201 (N_2201,N_1393,N_1060);
nand U2202 (N_2202,N_889,N_1023);
nor U2203 (N_2203,N_759,N_1098);
nand U2204 (N_2204,N_879,N_1116);
nor U2205 (N_2205,N_1227,N_1136);
nor U2206 (N_2206,N_1046,N_771);
nor U2207 (N_2207,N_811,N_1440);
nand U2208 (N_2208,N_842,N_951);
nor U2209 (N_2209,N_785,N_1460);
or U2210 (N_2210,N_1009,N_1290);
and U2211 (N_2211,N_916,N_885);
nor U2212 (N_2212,N_1117,N_1197);
nand U2213 (N_2213,N_1135,N_840);
or U2214 (N_2214,N_1155,N_1276);
nand U2215 (N_2215,N_824,N_1287);
nor U2216 (N_2216,N_1304,N_1028);
and U2217 (N_2217,N_1412,N_1395);
nor U2218 (N_2218,N_1363,N_1319);
xor U2219 (N_2219,N_1144,N_870);
nor U2220 (N_2220,N_1219,N_1450);
or U2221 (N_2221,N_1450,N_1222);
nand U2222 (N_2222,N_1199,N_1141);
nor U2223 (N_2223,N_1187,N_798);
nor U2224 (N_2224,N_919,N_1050);
nand U2225 (N_2225,N_857,N_1162);
nor U2226 (N_2226,N_1212,N_1051);
nor U2227 (N_2227,N_1295,N_947);
xor U2228 (N_2228,N_1160,N_1173);
nor U2229 (N_2229,N_1180,N_892);
and U2230 (N_2230,N_969,N_1019);
xnor U2231 (N_2231,N_1177,N_1020);
nor U2232 (N_2232,N_934,N_1399);
nor U2233 (N_2233,N_1426,N_1056);
or U2234 (N_2234,N_950,N_1143);
and U2235 (N_2235,N_835,N_832);
or U2236 (N_2236,N_1295,N_814);
xnor U2237 (N_2237,N_1334,N_1288);
and U2238 (N_2238,N_813,N_1273);
and U2239 (N_2239,N_1378,N_1482);
and U2240 (N_2240,N_1080,N_1013);
and U2241 (N_2241,N_976,N_1122);
nand U2242 (N_2242,N_785,N_1000);
nand U2243 (N_2243,N_1403,N_1035);
or U2244 (N_2244,N_1042,N_904);
nor U2245 (N_2245,N_1389,N_829);
xnor U2246 (N_2246,N_1421,N_1030);
nand U2247 (N_2247,N_1370,N_1134);
nor U2248 (N_2248,N_1405,N_919);
nor U2249 (N_2249,N_1140,N_806);
and U2250 (N_2250,N_1675,N_1903);
nor U2251 (N_2251,N_2089,N_1558);
or U2252 (N_2252,N_1898,N_1798);
or U2253 (N_2253,N_1573,N_2130);
xor U2254 (N_2254,N_1819,N_2221);
nor U2255 (N_2255,N_2132,N_1679);
and U2256 (N_2256,N_1859,N_1935);
nor U2257 (N_2257,N_1923,N_1728);
nand U2258 (N_2258,N_1927,N_2111);
or U2259 (N_2259,N_2035,N_2152);
or U2260 (N_2260,N_2086,N_2137);
xor U2261 (N_2261,N_2147,N_2167);
nand U2262 (N_2262,N_1947,N_2235);
nor U2263 (N_2263,N_1980,N_2170);
and U2264 (N_2264,N_2045,N_1774);
xor U2265 (N_2265,N_2034,N_1534);
and U2266 (N_2266,N_1684,N_1711);
or U2267 (N_2267,N_2107,N_2144);
nand U2268 (N_2268,N_2009,N_2239);
nor U2269 (N_2269,N_1581,N_1755);
xor U2270 (N_2270,N_1960,N_2155);
or U2271 (N_2271,N_1541,N_1674);
or U2272 (N_2272,N_1545,N_1530);
and U2273 (N_2273,N_1589,N_2242);
nand U2274 (N_2274,N_2102,N_1650);
and U2275 (N_2275,N_1669,N_1591);
and U2276 (N_2276,N_1732,N_2098);
nor U2277 (N_2277,N_1824,N_1769);
xor U2278 (N_2278,N_1602,N_1790);
or U2279 (N_2279,N_1951,N_2018);
nor U2280 (N_2280,N_1686,N_1835);
nand U2281 (N_2281,N_1636,N_1954);
nor U2282 (N_2282,N_2210,N_1713);
or U2283 (N_2283,N_2093,N_1531);
and U2284 (N_2284,N_1788,N_1916);
nand U2285 (N_2285,N_1784,N_1995);
or U2286 (N_2286,N_2044,N_2194);
xnor U2287 (N_2287,N_1812,N_2134);
or U2288 (N_2288,N_2218,N_2043);
and U2289 (N_2289,N_1656,N_1629);
nand U2290 (N_2290,N_1685,N_1932);
nor U2291 (N_2291,N_1518,N_1817);
nand U2292 (N_2292,N_1516,N_1867);
nor U2293 (N_2293,N_1642,N_1949);
nand U2294 (N_2294,N_2056,N_1597);
xor U2295 (N_2295,N_1557,N_2165);
or U2296 (N_2296,N_2094,N_1938);
or U2297 (N_2297,N_1576,N_2096);
nand U2298 (N_2298,N_1598,N_2081);
nand U2299 (N_2299,N_1767,N_1751);
nand U2300 (N_2300,N_2225,N_2070);
and U2301 (N_2301,N_1506,N_1512);
and U2302 (N_2302,N_1811,N_2217);
nor U2303 (N_2303,N_1841,N_1918);
nor U2304 (N_2304,N_1894,N_2198);
or U2305 (N_2305,N_1565,N_2157);
and U2306 (N_2306,N_1912,N_1885);
nand U2307 (N_2307,N_1550,N_1974);
or U2308 (N_2308,N_1800,N_1744);
xor U2309 (N_2309,N_1806,N_1723);
or U2310 (N_2310,N_1758,N_1992);
and U2311 (N_2311,N_1846,N_2017);
nor U2312 (N_2312,N_1890,N_1663);
nor U2313 (N_2313,N_1622,N_1771);
nor U2314 (N_2314,N_1941,N_2076);
nor U2315 (N_2315,N_1718,N_1801);
xor U2316 (N_2316,N_2237,N_1639);
nor U2317 (N_2317,N_2050,N_1608);
nor U2318 (N_2318,N_1860,N_1568);
xnor U2319 (N_2319,N_1546,N_1939);
nor U2320 (N_2320,N_1840,N_2088);
xnor U2321 (N_2321,N_1561,N_1925);
xnor U2322 (N_2322,N_1687,N_1627);
nor U2323 (N_2323,N_2247,N_2115);
nand U2324 (N_2324,N_1843,N_2154);
nand U2325 (N_2325,N_1778,N_1962);
nand U2326 (N_2326,N_1535,N_1910);
nor U2327 (N_2327,N_2146,N_2003);
nor U2328 (N_2328,N_1761,N_1854);
and U2329 (N_2329,N_1628,N_2118);
or U2330 (N_2330,N_1651,N_1705);
nor U2331 (N_2331,N_2077,N_1708);
and U2332 (N_2332,N_1845,N_1654);
and U2333 (N_2333,N_2249,N_1507);
or U2334 (N_2334,N_1842,N_2203);
nand U2335 (N_2335,N_1502,N_1552);
xor U2336 (N_2336,N_2151,N_2124);
and U2337 (N_2337,N_2092,N_1961);
and U2338 (N_2338,N_2209,N_1869);
nand U2339 (N_2339,N_1604,N_1830);
nor U2340 (N_2340,N_1765,N_1934);
and U2341 (N_2341,N_2192,N_2214);
nor U2342 (N_2342,N_1839,N_1688);
or U2343 (N_2343,N_1511,N_1500);
nand U2344 (N_2344,N_1795,N_2110);
or U2345 (N_2345,N_1953,N_1920);
xnor U2346 (N_2346,N_1596,N_2238);
and U2347 (N_2347,N_1553,N_1559);
nand U2348 (N_2348,N_2159,N_1979);
or U2349 (N_2349,N_2055,N_1937);
and U2350 (N_2350,N_2000,N_1619);
nand U2351 (N_2351,N_2207,N_1556);
nor U2352 (N_2352,N_1584,N_1532);
and U2353 (N_2353,N_1678,N_2100);
and U2354 (N_2354,N_1831,N_2240);
and U2355 (N_2355,N_1696,N_1536);
nor U2356 (N_2356,N_1641,N_2121);
or U2357 (N_2357,N_1549,N_2069);
or U2358 (N_2358,N_1714,N_2164);
xor U2359 (N_2359,N_2173,N_1733);
and U2360 (N_2360,N_2053,N_1902);
nor U2361 (N_2361,N_1926,N_2143);
or U2362 (N_2362,N_1599,N_1544);
and U2363 (N_2363,N_1689,N_1838);
and U2364 (N_2364,N_1540,N_1870);
nand U2365 (N_2365,N_2227,N_2150);
nand U2366 (N_2366,N_1809,N_1982);
or U2367 (N_2367,N_2156,N_1554);
or U2368 (N_2368,N_2244,N_1970);
nor U2369 (N_2369,N_2114,N_2041);
nor U2370 (N_2370,N_1753,N_2083);
and U2371 (N_2371,N_2188,N_1590);
or U2372 (N_2372,N_1803,N_2185);
nor U2373 (N_2373,N_1924,N_1989);
nor U2374 (N_2374,N_1551,N_1501);
or U2375 (N_2375,N_1818,N_2027);
nor U2376 (N_2376,N_1983,N_1736);
or U2377 (N_2377,N_1853,N_2108);
and U2378 (N_2378,N_1847,N_2020);
nor U2379 (N_2379,N_1682,N_1569);
or U2380 (N_2380,N_2029,N_1702);
nand U2381 (N_2381,N_1746,N_2037);
and U2382 (N_2382,N_1700,N_2106);
xor U2383 (N_2383,N_1644,N_2140);
nand U2384 (N_2384,N_1921,N_2223);
nand U2385 (N_2385,N_1560,N_2176);
and U2386 (N_2386,N_1695,N_1849);
nand U2387 (N_2387,N_1660,N_1704);
or U2388 (N_2388,N_1635,N_1865);
nor U2389 (N_2389,N_1958,N_2048);
or U2390 (N_2390,N_1827,N_2153);
and U2391 (N_2391,N_1889,N_1523);
nand U2392 (N_2392,N_1863,N_1617);
nor U2393 (N_2393,N_1822,N_1878);
or U2394 (N_2394,N_2195,N_1609);
nor U2395 (N_2395,N_2141,N_1738);
nand U2396 (N_2396,N_1647,N_1607);
xor U2397 (N_2397,N_1907,N_1808);
or U2398 (N_2398,N_1826,N_1509);
and U2399 (N_2399,N_1881,N_1710);
or U2400 (N_2400,N_1631,N_1991);
nor U2401 (N_2401,N_1566,N_1524);
or U2402 (N_2402,N_1630,N_2162);
and U2403 (N_2403,N_1868,N_1821);
nand U2404 (N_2404,N_2065,N_1794);
nand U2405 (N_2405,N_1655,N_1836);
or U2406 (N_2406,N_1866,N_2202);
and U2407 (N_2407,N_1929,N_1975);
and U2408 (N_2408,N_1779,N_2233);
and U2409 (N_2409,N_1693,N_2191);
xor U2410 (N_2410,N_2026,N_1786);
and U2411 (N_2411,N_1973,N_2099);
or U2412 (N_2412,N_2113,N_2245);
and U2413 (N_2413,N_2145,N_2142);
and U2414 (N_2414,N_2004,N_1762);
and U2415 (N_2415,N_1747,N_1768);
nand U2416 (N_2416,N_1592,N_1967);
and U2417 (N_2417,N_2193,N_1787);
and U2418 (N_2418,N_1611,N_1580);
nor U2419 (N_2419,N_2011,N_1897);
and U2420 (N_2420,N_1643,N_1943);
nand U2421 (N_2421,N_1579,N_1600);
or U2422 (N_2422,N_1538,N_1972);
nand U2423 (N_2423,N_2126,N_2022);
xor U2424 (N_2424,N_2189,N_1749);
nor U2425 (N_2425,N_1837,N_1857);
nor U2426 (N_2426,N_1701,N_2206);
nor U2427 (N_2427,N_1950,N_2116);
or U2428 (N_2428,N_1883,N_1616);
nor U2429 (N_2429,N_2059,N_1896);
nor U2430 (N_2430,N_1969,N_2030);
and U2431 (N_2431,N_1880,N_1681);
or U2432 (N_2432,N_2234,N_1539);
nor U2433 (N_2433,N_1760,N_2128);
nand U2434 (N_2434,N_1624,N_1677);
or U2435 (N_2435,N_1873,N_1990);
or U2436 (N_2436,N_1529,N_1717);
nand U2437 (N_2437,N_2101,N_1887);
nor U2438 (N_2438,N_1922,N_1882);
nor U2439 (N_2439,N_1993,N_1940);
or U2440 (N_2440,N_2169,N_1913);
nor U2441 (N_2441,N_2119,N_1895);
xor U2442 (N_2442,N_1716,N_1668);
or U2443 (N_2443,N_1741,N_2047);
or U2444 (N_2444,N_1645,N_2248);
or U2445 (N_2445,N_1513,N_2211);
and U2446 (N_2446,N_1740,N_1904);
and U2447 (N_2447,N_2177,N_1931);
and U2448 (N_2448,N_2179,N_1994);
or U2449 (N_2449,N_2212,N_1968);
nand U2450 (N_2450,N_1942,N_1909);
or U2451 (N_2451,N_2133,N_1754);
and U2452 (N_2452,N_1582,N_1661);
or U2453 (N_2453,N_2186,N_1706);
nor U2454 (N_2454,N_1877,N_1725);
or U2455 (N_2455,N_1504,N_2105);
nor U2456 (N_2456,N_1613,N_1875);
nor U2457 (N_2457,N_2057,N_1653);
and U2458 (N_2458,N_1832,N_2138);
and U2459 (N_2459,N_1637,N_1804);
nor U2460 (N_2460,N_2015,N_1911);
and U2461 (N_2461,N_1652,N_1562);
and U2462 (N_2462,N_2163,N_2091);
nor U2463 (N_2463,N_2016,N_1640);
and U2464 (N_2464,N_2012,N_1763);
or U2465 (N_2465,N_2073,N_1595);
nor U2466 (N_2466,N_1662,N_1879);
or U2467 (N_2467,N_1782,N_1621);
and U2468 (N_2468,N_2161,N_1884);
nand U2469 (N_2469,N_1730,N_1720);
xor U2470 (N_2470,N_2236,N_2068);
nor U2471 (N_2471,N_1525,N_1807);
xnor U2472 (N_2472,N_2136,N_2220);
or U2473 (N_2473,N_1690,N_2246);
xor U2474 (N_2474,N_1697,N_1521);
nor U2475 (N_2475,N_1583,N_1930);
xnor U2476 (N_2476,N_1984,N_2122);
nand U2477 (N_2477,N_1862,N_1917);
xnor U2478 (N_2478,N_2120,N_1764);
and U2479 (N_2479,N_1542,N_1585);
nand U2480 (N_2480,N_1721,N_2013);
xor U2481 (N_2481,N_1986,N_1748);
nand U2482 (N_2482,N_1814,N_1646);
nor U2483 (N_2483,N_1892,N_1861);
nor U2484 (N_2484,N_1633,N_1734);
or U2485 (N_2485,N_1743,N_1649);
or U2486 (N_2486,N_1729,N_1900);
or U2487 (N_2487,N_1999,N_1864);
nor U2488 (N_2488,N_1945,N_2184);
or U2489 (N_2489,N_1955,N_2181);
or U2490 (N_2490,N_1978,N_2219);
and U2491 (N_2491,N_1603,N_2149);
and U2492 (N_2492,N_1785,N_1520);
or U2493 (N_2493,N_2172,N_1555);
nor U2494 (N_2494,N_1745,N_1572);
nand U2495 (N_2495,N_1776,N_1810);
nand U2496 (N_2496,N_1850,N_1965);
or U2497 (N_2497,N_2019,N_1606);
nand U2498 (N_2498,N_2006,N_1952);
nand U2499 (N_2499,N_1766,N_1852);
nand U2500 (N_2500,N_1620,N_1618);
nor U2501 (N_2501,N_1671,N_1833);
nand U2502 (N_2502,N_2168,N_2200);
and U2503 (N_2503,N_1759,N_1505);
xnor U2504 (N_2504,N_1739,N_1543);
and U2505 (N_2505,N_1680,N_1672);
nor U2506 (N_2506,N_2052,N_2005);
and U2507 (N_2507,N_1752,N_2040);
nand U2508 (N_2508,N_1998,N_1914);
nand U2509 (N_2509,N_1816,N_2066);
and U2510 (N_2510,N_1574,N_1789);
nand U2511 (N_2511,N_1691,N_1510);
xnor U2512 (N_2512,N_1805,N_1508);
nor U2513 (N_2513,N_1694,N_2085);
nand U2514 (N_2514,N_1527,N_2213);
nor U2515 (N_2515,N_2078,N_2230);
or U2516 (N_2516,N_1515,N_1563);
nor U2517 (N_2517,N_1564,N_2208);
nor U2518 (N_2518,N_1829,N_1692);
and U2519 (N_2519,N_2042,N_1632);
nor U2520 (N_2520,N_2204,N_1594);
and U2521 (N_2521,N_1626,N_2032);
and U2522 (N_2522,N_1673,N_2033);
nor U2523 (N_2523,N_1933,N_1966);
nor U2524 (N_2524,N_1605,N_2104);
and U2525 (N_2525,N_1514,N_2190);
xor U2526 (N_2526,N_2135,N_1855);
nor U2527 (N_2527,N_2166,N_1872);
or U2528 (N_2528,N_1797,N_2231);
or U2529 (N_2529,N_2123,N_1614);
and U2530 (N_2530,N_1737,N_1871);
nand U2531 (N_2531,N_1777,N_1712);
nand U2532 (N_2532,N_2008,N_1570);
nand U2533 (N_2533,N_1683,N_1919);
nor U2534 (N_2534,N_2222,N_2067);
nor U2535 (N_2535,N_1593,N_1815);
nor U2536 (N_2536,N_1665,N_2060);
nand U2537 (N_2537,N_1659,N_2183);
or U2538 (N_2538,N_1775,N_1772);
nor U2539 (N_2539,N_1988,N_1773);
or U2540 (N_2540,N_1844,N_2131);
nor U2541 (N_2541,N_2197,N_2125);
nor U2542 (N_2542,N_2174,N_1780);
xnor U2543 (N_2543,N_1802,N_1963);
or U2544 (N_2544,N_1825,N_2025);
or U2545 (N_2545,N_2087,N_2160);
or U2546 (N_2546,N_1731,N_1715);
or U2547 (N_2547,N_1528,N_1959);
nor U2548 (N_2548,N_2010,N_1670);
and U2549 (N_2549,N_1996,N_2178);
nand U2550 (N_2550,N_2228,N_1699);
or U2551 (N_2551,N_1756,N_2084);
nand U2552 (N_2552,N_1820,N_1526);
nor U2553 (N_2553,N_2054,N_2064);
and U2554 (N_2554,N_2139,N_2051);
nor U2555 (N_2555,N_2196,N_2205);
nand U2556 (N_2556,N_1899,N_1858);
nor U2557 (N_2557,N_2243,N_1948);
nor U2558 (N_2558,N_1905,N_1888);
nor U2559 (N_2559,N_1658,N_1997);
nor U2560 (N_2560,N_2001,N_1908);
xor U2561 (N_2561,N_1735,N_2072);
or U2562 (N_2562,N_1601,N_2180);
or U2563 (N_2563,N_2187,N_2058);
or U2564 (N_2564,N_1577,N_2090);
xnor U2565 (N_2565,N_1987,N_2127);
nand U2566 (N_2566,N_1813,N_1623);
and U2567 (N_2567,N_1727,N_1971);
and U2568 (N_2568,N_1781,N_1547);
xor U2569 (N_2569,N_1928,N_2014);
nor U2570 (N_2570,N_2232,N_1823);
and U2571 (N_2571,N_1783,N_2117);
nor U2572 (N_2572,N_2046,N_1893);
or U2573 (N_2573,N_1664,N_1719);
and U2574 (N_2574,N_1956,N_2074);
nand U2575 (N_2575,N_2201,N_1915);
nand U2576 (N_2576,N_1799,N_1648);
nand U2577 (N_2577,N_1517,N_2002);
nand U2578 (N_2578,N_1634,N_2158);
nor U2579 (N_2579,N_1610,N_1828);
xnor U2580 (N_2580,N_1985,N_2215);
or U2581 (N_2581,N_1703,N_1976);
or U2582 (N_2582,N_1612,N_1944);
xor U2583 (N_2583,N_2049,N_1666);
nor U2584 (N_2584,N_1578,N_2071);
nand U2585 (N_2585,N_2079,N_1901);
or U2586 (N_2586,N_1667,N_1638);
nor U2587 (N_2587,N_2097,N_1792);
nor U2588 (N_2588,N_2109,N_1722);
xor U2589 (N_2589,N_1874,N_2175);
or U2590 (N_2590,N_2216,N_2199);
nand U2591 (N_2591,N_2229,N_1856);
or U2592 (N_2592,N_1709,N_2148);
nand U2593 (N_2593,N_1522,N_1657);
nand U2594 (N_2594,N_1886,N_2023);
nand U2595 (N_2595,N_1977,N_2039);
nor U2596 (N_2596,N_1757,N_2080);
nor U2597 (N_2597,N_1571,N_2038);
nor U2598 (N_2598,N_2031,N_2061);
nor U2599 (N_2599,N_1964,N_2063);
or U2600 (N_2600,N_2062,N_2103);
nor U2601 (N_2601,N_1587,N_1503);
or U2602 (N_2602,N_1698,N_1946);
and U2603 (N_2603,N_1575,N_2007);
nor U2604 (N_2604,N_1876,N_2095);
or U2605 (N_2605,N_2224,N_1533);
xor U2606 (N_2606,N_1957,N_1548);
nand U2607 (N_2607,N_2226,N_1519);
or U2608 (N_2608,N_1936,N_1625);
nand U2609 (N_2609,N_1676,N_1586);
nor U2610 (N_2610,N_2129,N_2075);
and U2611 (N_2611,N_2112,N_2021);
and U2612 (N_2612,N_2028,N_1770);
and U2613 (N_2613,N_1791,N_1537);
and U2614 (N_2614,N_1615,N_1851);
nand U2615 (N_2615,N_2024,N_1726);
nand U2616 (N_2616,N_2171,N_1796);
nor U2617 (N_2617,N_1567,N_1724);
or U2618 (N_2618,N_1891,N_2241);
or U2619 (N_2619,N_1742,N_1588);
or U2620 (N_2620,N_2082,N_1848);
nand U2621 (N_2621,N_1707,N_1793);
xor U2622 (N_2622,N_1981,N_1834);
or U2623 (N_2623,N_2036,N_1750);
or U2624 (N_2624,N_1906,N_2182);
nand U2625 (N_2625,N_1814,N_1889);
and U2626 (N_2626,N_2025,N_2213);
nand U2627 (N_2627,N_1618,N_2044);
nor U2628 (N_2628,N_2186,N_2063);
nor U2629 (N_2629,N_1686,N_2190);
xor U2630 (N_2630,N_1823,N_1581);
nor U2631 (N_2631,N_2176,N_2122);
nand U2632 (N_2632,N_1632,N_2155);
or U2633 (N_2633,N_2138,N_1951);
or U2634 (N_2634,N_1603,N_1644);
nor U2635 (N_2635,N_1571,N_2235);
nor U2636 (N_2636,N_1782,N_1995);
or U2637 (N_2637,N_1543,N_1999);
or U2638 (N_2638,N_2070,N_2186);
or U2639 (N_2639,N_1932,N_1970);
or U2640 (N_2640,N_1736,N_2048);
and U2641 (N_2641,N_1648,N_1691);
and U2642 (N_2642,N_2008,N_1827);
and U2643 (N_2643,N_2154,N_2214);
or U2644 (N_2644,N_2197,N_1734);
nor U2645 (N_2645,N_1937,N_2249);
nor U2646 (N_2646,N_1582,N_2232);
nor U2647 (N_2647,N_2022,N_1609);
or U2648 (N_2648,N_1666,N_1968);
or U2649 (N_2649,N_2090,N_1714);
or U2650 (N_2650,N_1658,N_1899);
nor U2651 (N_2651,N_1896,N_1706);
nor U2652 (N_2652,N_1746,N_1579);
or U2653 (N_2653,N_2164,N_1723);
and U2654 (N_2654,N_2132,N_1629);
or U2655 (N_2655,N_2018,N_1654);
or U2656 (N_2656,N_2104,N_1690);
nor U2657 (N_2657,N_1664,N_2059);
nand U2658 (N_2658,N_1805,N_2180);
nand U2659 (N_2659,N_1928,N_1887);
or U2660 (N_2660,N_2040,N_1542);
and U2661 (N_2661,N_2093,N_2053);
and U2662 (N_2662,N_2138,N_1598);
nand U2663 (N_2663,N_2139,N_1599);
nor U2664 (N_2664,N_1815,N_1819);
and U2665 (N_2665,N_1725,N_1605);
nor U2666 (N_2666,N_2193,N_1930);
nand U2667 (N_2667,N_1725,N_1845);
or U2668 (N_2668,N_1587,N_1919);
nor U2669 (N_2669,N_1665,N_2024);
nor U2670 (N_2670,N_1942,N_1934);
and U2671 (N_2671,N_2090,N_2162);
nand U2672 (N_2672,N_1556,N_1799);
or U2673 (N_2673,N_1854,N_1814);
and U2674 (N_2674,N_2214,N_1911);
and U2675 (N_2675,N_1928,N_1542);
nand U2676 (N_2676,N_1951,N_2125);
and U2677 (N_2677,N_2066,N_1915);
nand U2678 (N_2678,N_1967,N_1712);
nor U2679 (N_2679,N_2237,N_1696);
and U2680 (N_2680,N_1575,N_1719);
and U2681 (N_2681,N_1635,N_1812);
nor U2682 (N_2682,N_1783,N_1949);
or U2683 (N_2683,N_2169,N_1990);
nand U2684 (N_2684,N_1613,N_1842);
nand U2685 (N_2685,N_1534,N_1714);
nor U2686 (N_2686,N_1838,N_1931);
nor U2687 (N_2687,N_1754,N_2212);
nor U2688 (N_2688,N_1631,N_1606);
nand U2689 (N_2689,N_1625,N_1512);
nor U2690 (N_2690,N_2084,N_2160);
nand U2691 (N_2691,N_2023,N_2140);
nand U2692 (N_2692,N_1718,N_2230);
xor U2693 (N_2693,N_1987,N_2129);
and U2694 (N_2694,N_1647,N_2184);
nand U2695 (N_2695,N_2117,N_1807);
and U2696 (N_2696,N_1850,N_1967);
and U2697 (N_2697,N_1733,N_1869);
or U2698 (N_2698,N_2136,N_2189);
xnor U2699 (N_2699,N_2030,N_1904);
nor U2700 (N_2700,N_2199,N_1507);
and U2701 (N_2701,N_1513,N_1561);
and U2702 (N_2702,N_1915,N_2109);
nand U2703 (N_2703,N_1776,N_1891);
nor U2704 (N_2704,N_1990,N_1517);
and U2705 (N_2705,N_1593,N_1967);
nor U2706 (N_2706,N_2185,N_1725);
and U2707 (N_2707,N_1998,N_2205);
or U2708 (N_2708,N_2145,N_1614);
and U2709 (N_2709,N_1692,N_2066);
nor U2710 (N_2710,N_1529,N_2004);
and U2711 (N_2711,N_1859,N_1961);
or U2712 (N_2712,N_2231,N_1981);
nand U2713 (N_2713,N_1941,N_1768);
or U2714 (N_2714,N_1711,N_1633);
xor U2715 (N_2715,N_1651,N_1801);
and U2716 (N_2716,N_2109,N_1751);
or U2717 (N_2717,N_1766,N_2080);
nand U2718 (N_2718,N_2036,N_1881);
nand U2719 (N_2719,N_1818,N_2123);
or U2720 (N_2720,N_2142,N_1559);
or U2721 (N_2721,N_1780,N_1550);
nor U2722 (N_2722,N_2248,N_1903);
nand U2723 (N_2723,N_1939,N_2213);
nand U2724 (N_2724,N_2189,N_1532);
nand U2725 (N_2725,N_1629,N_1601);
xor U2726 (N_2726,N_2230,N_1905);
nand U2727 (N_2727,N_1771,N_1565);
or U2728 (N_2728,N_2026,N_2184);
or U2729 (N_2729,N_1796,N_1892);
or U2730 (N_2730,N_1952,N_1515);
and U2731 (N_2731,N_1805,N_2071);
nand U2732 (N_2732,N_1766,N_1870);
nand U2733 (N_2733,N_1839,N_1617);
nor U2734 (N_2734,N_1639,N_1996);
or U2735 (N_2735,N_1847,N_2113);
and U2736 (N_2736,N_2218,N_2152);
and U2737 (N_2737,N_1811,N_1873);
nand U2738 (N_2738,N_1951,N_1523);
and U2739 (N_2739,N_1968,N_2112);
nor U2740 (N_2740,N_1927,N_2246);
nor U2741 (N_2741,N_1603,N_2025);
nor U2742 (N_2742,N_1726,N_1770);
and U2743 (N_2743,N_2235,N_2212);
nor U2744 (N_2744,N_1962,N_2003);
xnor U2745 (N_2745,N_1845,N_1894);
nand U2746 (N_2746,N_1630,N_2242);
and U2747 (N_2747,N_1720,N_1867);
or U2748 (N_2748,N_2036,N_2040);
nand U2749 (N_2749,N_2191,N_1999);
nor U2750 (N_2750,N_2167,N_1824);
nand U2751 (N_2751,N_1616,N_2094);
nand U2752 (N_2752,N_2157,N_1592);
nor U2753 (N_2753,N_1981,N_1574);
xnor U2754 (N_2754,N_2237,N_2139);
xnor U2755 (N_2755,N_1933,N_1726);
nand U2756 (N_2756,N_1817,N_1709);
nand U2757 (N_2757,N_1682,N_1993);
nor U2758 (N_2758,N_1789,N_1757);
and U2759 (N_2759,N_1791,N_1994);
or U2760 (N_2760,N_1632,N_2244);
nor U2761 (N_2761,N_1959,N_2153);
nor U2762 (N_2762,N_1890,N_1984);
or U2763 (N_2763,N_1893,N_1862);
xnor U2764 (N_2764,N_2188,N_1776);
or U2765 (N_2765,N_2106,N_1651);
nor U2766 (N_2766,N_1562,N_2124);
nand U2767 (N_2767,N_2088,N_1651);
or U2768 (N_2768,N_1752,N_1906);
nand U2769 (N_2769,N_1892,N_1764);
nand U2770 (N_2770,N_1718,N_1826);
or U2771 (N_2771,N_1619,N_2157);
nor U2772 (N_2772,N_1971,N_2198);
nor U2773 (N_2773,N_1698,N_2182);
or U2774 (N_2774,N_2127,N_2202);
nand U2775 (N_2775,N_2169,N_2009);
xor U2776 (N_2776,N_2118,N_2127);
or U2777 (N_2777,N_1785,N_1537);
xor U2778 (N_2778,N_2085,N_1707);
and U2779 (N_2779,N_1936,N_1676);
xor U2780 (N_2780,N_2172,N_1514);
or U2781 (N_2781,N_1900,N_1737);
nor U2782 (N_2782,N_1942,N_1950);
or U2783 (N_2783,N_1709,N_1837);
and U2784 (N_2784,N_1503,N_1514);
nor U2785 (N_2785,N_2012,N_2232);
nor U2786 (N_2786,N_1960,N_1763);
nor U2787 (N_2787,N_1591,N_1541);
or U2788 (N_2788,N_1505,N_1791);
or U2789 (N_2789,N_2086,N_1749);
and U2790 (N_2790,N_1575,N_1807);
nand U2791 (N_2791,N_1538,N_2119);
xnor U2792 (N_2792,N_1750,N_2109);
nand U2793 (N_2793,N_1760,N_1591);
xor U2794 (N_2794,N_1815,N_2103);
nor U2795 (N_2795,N_1901,N_1818);
and U2796 (N_2796,N_1741,N_1658);
or U2797 (N_2797,N_1584,N_1550);
or U2798 (N_2798,N_1842,N_1503);
nand U2799 (N_2799,N_1534,N_1842);
or U2800 (N_2800,N_1616,N_1720);
or U2801 (N_2801,N_1576,N_1725);
and U2802 (N_2802,N_2243,N_1811);
nor U2803 (N_2803,N_1612,N_1524);
or U2804 (N_2804,N_2053,N_2162);
and U2805 (N_2805,N_2221,N_1809);
xnor U2806 (N_2806,N_2070,N_2222);
and U2807 (N_2807,N_2225,N_1774);
nand U2808 (N_2808,N_2019,N_1707);
nor U2809 (N_2809,N_1739,N_1621);
nand U2810 (N_2810,N_1599,N_1618);
xor U2811 (N_2811,N_1924,N_1866);
nor U2812 (N_2812,N_1756,N_2106);
or U2813 (N_2813,N_1833,N_2085);
nand U2814 (N_2814,N_1788,N_1982);
or U2815 (N_2815,N_1960,N_1769);
nand U2816 (N_2816,N_2211,N_2215);
or U2817 (N_2817,N_1875,N_2116);
and U2818 (N_2818,N_1500,N_1917);
and U2819 (N_2819,N_1575,N_2142);
and U2820 (N_2820,N_2171,N_1682);
nand U2821 (N_2821,N_1886,N_2074);
nor U2822 (N_2822,N_2202,N_2206);
nor U2823 (N_2823,N_1691,N_2190);
nor U2824 (N_2824,N_2105,N_2043);
nor U2825 (N_2825,N_1571,N_2197);
or U2826 (N_2826,N_2150,N_1544);
or U2827 (N_2827,N_1740,N_1508);
nand U2828 (N_2828,N_1769,N_2181);
and U2829 (N_2829,N_1584,N_1693);
nor U2830 (N_2830,N_1878,N_1889);
nor U2831 (N_2831,N_2061,N_1554);
nor U2832 (N_2832,N_1527,N_1969);
or U2833 (N_2833,N_2121,N_1771);
and U2834 (N_2834,N_2028,N_2015);
nor U2835 (N_2835,N_1687,N_1942);
nand U2836 (N_2836,N_2149,N_2098);
nand U2837 (N_2837,N_2225,N_1698);
nand U2838 (N_2838,N_2092,N_1766);
and U2839 (N_2839,N_2231,N_1534);
nand U2840 (N_2840,N_1790,N_1859);
nor U2841 (N_2841,N_2197,N_1814);
nand U2842 (N_2842,N_1846,N_1992);
nand U2843 (N_2843,N_2040,N_1957);
nand U2844 (N_2844,N_2115,N_2157);
and U2845 (N_2845,N_1857,N_2198);
nand U2846 (N_2846,N_1806,N_2185);
and U2847 (N_2847,N_1730,N_2244);
nand U2848 (N_2848,N_2089,N_1917);
and U2849 (N_2849,N_1643,N_1565);
nor U2850 (N_2850,N_2153,N_1914);
and U2851 (N_2851,N_1809,N_1622);
and U2852 (N_2852,N_2045,N_1919);
or U2853 (N_2853,N_1906,N_2097);
and U2854 (N_2854,N_1506,N_2248);
and U2855 (N_2855,N_2031,N_1627);
nor U2856 (N_2856,N_1569,N_2244);
nor U2857 (N_2857,N_1974,N_1708);
nand U2858 (N_2858,N_1855,N_2119);
nand U2859 (N_2859,N_1650,N_1685);
and U2860 (N_2860,N_1734,N_1600);
or U2861 (N_2861,N_1660,N_1514);
or U2862 (N_2862,N_2137,N_2075);
nand U2863 (N_2863,N_1731,N_1802);
nand U2864 (N_2864,N_2107,N_1870);
or U2865 (N_2865,N_2077,N_2080);
nand U2866 (N_2866,N_2227,N_1788);
xor U2867 (N_2867,N_1588,N_2005);
nand U2868 (N_2868,N_2227,N_1880);
nand U2869 (N_2869,N_1667,N_1753);
and U2870 (N_2870,N_1855,N_1515);
or U2871 (N_2871,N_2188,N_1892);
nor U2872 (N_2872,N_1829,N_1656);
nor U2873 (N_2873,N_2057,N_1551);
and U2874 (N_2874,N_1921,N_1529);
or U2875 (N_2875,N_1602,N_1830);
or U2876 (N_2876,N_1541,N_1562);
nor U2877 (N_2877,N_1624,N_1630);
xor U2878 (N_2878,N_2108,N_2069);
and U2879 (N_2879,N_1563,N_1867);
and U2880 (N_2880,N_1772,N_2073);
or U2881 (N_2881,N_2230,N_1589);
and U2882 (N_2882,N_1628,N_1709);
nand U2883 (N_2883,N_1701,N_1974);
xor U2884 (N_2884,N_1597,N_1987);
nor U2885 (N_2885,N_1612,N_1753);
nand U2886 (N_2886,N_1677,N_1547);
xor U2887 (N_2887,N_1560,N_2040);
and U2888 (N_2888,N_1724,N_1811);
nor U2889 (N_2889,N_1934,N_1990);
and U2890 (N_2890,N_1751,N_2140);
nor U2891 (N_2891,N_1516,N_1734);
and U2892 (N_2892,N_2012,N_2205);
nor U2893 (N_2893,N_1641,N_2008);
and U2894 (N_2894,N_1747,N_1851);
nor U2895 (N_2895,N_1704,N_2244);
nand U2896 (N_2896,N_1975,N_1650);
nand U2897 (N_2897,N_1797,N_1523);
or U2898 (N_2898,N_1711,N_1502);
and U2899 (N_2899,N_1643,N_2079);
xnor U2900 (N_2900,N_1584,N_1508);
xor U2901 (N_2901,N_1912,N_1961);
and U2902 (N_2902,N_1667,N_2197);
nor U2903 (N_2903,N_1768,N_2089);
and U2904 (N_2904,N_1677,N_1886);
and U2905 (N_2905,N_1686,N_1553);
nand U2906 (N_2906,N_1830,N_2095);
xnor U2907 (N_2907,N_1948,N_1789);
and U2908 (N_2908,N_1911,N_2211);
nand U2909 (N_2909,N_2218,N_1941);
nand U2910 (N_2910,N_2232,N_1654);
and U2911 (N_2911,N_2109,N_1700);
nand U2912 (N_2912,N_1845,N_2137);
nand U2913 (N_2913,N_1702,N_2227);
xor U2914 (N_2914,N_1758,N_2025);
nand U2915 (N_2915,N_1736,N_1640);
nor U2916 (N_2916,N_2097,N_1594);
nand U2917 (N_2917,N_2238,N_1645);
nand U2918 (N_2918,N_2035,N_1913);
xor U2919 (N_2919,N_2220,N_2114);
nor U2920 (N_2920,N_2051,N_1769);
nand U2921 (N_2921,N_2062,N_1855);
or U2922 (N_2922,N_1799,N_1665);
and U2923 (N_2923,N_1929,N_1723);
nand U2924 (N_2924,N_2109,N_1634);
nand U2925 (N_2925,N_1645,N_1804);
nand U2926 (N_2926,N_2137,N_1944);
nor U2927 (N_2927,N_2093,N_1924);
xnor U2928 (N_2928,N_1757,N_1542);
nand U2929 (N_2929,N_1689,N_1546);
nor U2930 (N_2930,N_1766,N_1758);
nand U2931 (N_2931,N_1837,N_1742);
and U2932 (N_2932,N_2119,N_1518);
xnor U2933 (N_2933,N_2208,N_1946);
nand U2934 (N_2934,N_2022,N_1892);
or U2935 (N_2935,N_1810,N_2009);
and U2936 (N_2936,N_1665,N_1577);
xor U2937 (N_2937,N_1998,N_2002);
or U2938 (N_2938,N_2166,N_1851);
nand U2939 (N_2939,N_1689,N_1929);
nor U2940 (N_2940,N_1675,N_1767);
nand U2941 (N_2941,N_1911,N_1835);
nand U2942 (N_2942,N_2167,N_2062);
or U2943 (N_2943,N_1827,N_2100);
nand U2944 (N_2944,N_2227,N_1560);
or U2945 (N_2945,N_1901,N_2092);
or U2946 (N_2946,N_1535,N_1912);
nor U2947 (N_2947,N_1774,N_2013);
or U2948 (N_2948,N_2084,N_1697);
or U2949 (N_2949,N_2222,N_1668);
nand U2950 (N_2950,N_2069,N_1740);
nand U2951 (N_2951,N_1702,N_1583);
nor U2952 (N_2952,N_2019,N_1573);
and U2953 (N_2953,N_1721,N_1591);
nor U2954 (N_2954,N_1892,N_1682);
nand U2955 (N_2955,N_2000,N_1781);
xnor U2956 (N_2956,N_2173,N_1606);
nor U2957 (N_2957,N_1929,N_2004);
or U2958 (N_2958,N_1821,N_1723);
nor U2959 (N_2959,N_1686,N_1874);
or U2960 (N_2960,N_1677,N_2035);
xor U2961 (N_2961,N_2011,N_2240);
xor U2962 (N_2962,N_1508,N_2034);
nand U2963 (N_2963,N_1692,N_1873);
or U2964 (N_2964,N_1994,N_2168);
xor U2965 (N_2965,N_2209,N_1787);
xor U2966 (N_2966,N_1993,N_2207);
nor U2967 (N_2967,N_2032,N_1688);
and U2968 (N_2968,N_1615,N_1712);
or U2969 (N_2969,N_1883,N_1877);
and U2970 (N_2970,N_1634,N_2072);
or U2971 (N_2971,N_1529,N_1969);
nor U2972 (N_2972,N_2043,N_1586);
or U2973 (N_2973,N_1770,N_1730);
and U2974 (N_2974,N_1734,N_1631);
nand U2975 (N_2975,N_1959,N_2225);
xnor U2976 (N_2976,N_1888,N_1967);
nand U2977 (N_2977,N_1572,N_1731);
and U2978 (N_2978,N_2067,N_2198);
nand U2979 (N_2979,N_1886,N_1990);
nand U2980 (N_2980,N_2179,N_1687);
nand U2981 (N_2981,N_2245,N_1901);
xnor U2982 (N_2982,N_2060,N_2249);
and U2983 (N_2983,N_1521,N_1898);
and U2984 (N_2984,N_2214,N_2160);
nor U2985 (N_2985,N_1981,N_2043);
and U2986 (N_2986,N_2119,N_1890);
nand U2987 (N_2987,N_1867,N_1703);
and U2988 (N_2988,N_1603,N_1763);
or U2989 (N_2989,N_1511,N_1834);
and U2990 (N_2990,N_2030,N_1657);
or U2991 (N_2991,N_2190,N_2223);
nand U2992 (N_2992,N_1781,N_1616);
nor U2993 (N_2993,N_1733,N_1915);
nand U2994 (N_2994,N_1766,N_1820);
or U2995 (N_2995,N_1600,N_1878);
nor U2996 (N_2996,N_2049,N_1842);
and U2997 (N_2997,N_1718,N_1613);
and U2998 (N_2998,N_1551,N_2117);
nand U2999 (N_2999,N_1851,N_1977);
and UO_0 (O_0,N_2402,N_2615);
nand UO_1 (O_1,N_2907,N_2604);
or UO_2 (O_2,N_2983,N_2609);
xor UO_3 (O_3,N_2341,N_2773);
and UO_4 (O_4,N_2367,N_2479);
nor UO_5 (O_5,N_2390,N_2380);
and UO_6 (O_6,N_2544,N_2972);
and UO_7 (O_7,N_2499,N_2725);
and UO_8 (O_8,N_2962,N_2373);
nand UO_9 (O_9,N_2484,N_2848);
nand UO_10 (O_10,N_2508,N_2478);
nor UO_11 (O_11,N_2671,N_2502);
nor UO_12 (O_12,N_2886,N_2562);
and UO_13 (O_13,N_2441,N_2446);
nor UO_14 (O_14,N_2767,N_2800);
and UO_15 (O_15,N_2771,N_2985);
and UO_16 (O_16,N_2707,N_2308);
nor UO_17 (O_17,N_2718,N_2444);
and UO_18 (O_18,N_2666,N_2371);
nand UO_19 (O_19,N_2255,N_2860);
or UO_20 (O_20,N_2291,N_2931);
nand UO_21 (O_21,N_2251,N_2625);
nor UO_22 (O_22,N_2558,N_2489);
nor UO_23 (O_23,N_2997,N_2559);
nor UO_24 (O_24,N_2847,N_2525);
nand UO_25 (O_25,N_2394,N_2460);
nor UO_26 (O_26,N_2824,N_2778);
xnor UO_27 (O_27,N_2415,N_2664);
and UO_28 (O_28,N_2293,N_2665);
or UO_29 (O_29,N_2851,N_2328);
nor UO_30 (O_30,N_2651,N_2713);
nor UO_31 (O_31,N_2896,N_2700);
nand UO_32 (O_32,N_2546,N_2762);
nand UO_33 (O_33,N_2335,N_2473);
nand UO_34 (O_34,N_2738,N_2881);
and UO_35 (O_35,N_2463,N_2898);
nand UO_36 (O_36,N_2507,N_2536);
or UO_37 (O_37,N_2472,N_2676);
nor UO_38 (O_38,N_2561,N_2386);
and UO_39 (O_39,N_2693,N_2869);
or UO_40 (O_40,N_2855,N_2864);
nand UO_41 (O_41,N_2570,N_2612);
xor UO_42 (O_42,N_2565,N_2452);
nor UO_43 (O_43,N_2946,N_2978);
or UO_44 (O_44,N_2843,N_2515);
and UO_45 (O_45,N_2289,N_2916);
nor UO_46 (O_46,N_2344,N_2425);
or UO_47 (O_47,N_2370,N_2556);
nand UO_48 (O_48,N_2524,N_2459);
and UO_49 (O_49,N_2528,N_2654);
or UO_50 (O_50,N_2971,N_2863);
and UO_51 (O_51,N_2833,N_2622);
nor UO_52 (O_52,N_2974,N_2590);
or UO_53 (O_53,N_2375,N_2644);
or UO_54 (O_54,N_2492,N_2657);
nor UO_55 (O_55,N_2698,N_2840);
xor UO_56 (O_56,N_2741,N_2831);
nor UO_57 (O_57,N_2826,N_2715);
nand UO_58 (O_58,N_2280,N_2936);
nand UO_59 (O_59,N_2350,N_2769);
nand UO_60 (O_60,N_2277,N_2391);
nor UO_61 (O_61,N_2818,N_2338);
and UO_62 (O_62,N_2469,N_2804);
nor UO_63 (O_63,N_2992,N_2608);
nand UO_64 (O_64,N_2600,N_2772);
nand UO_65 (O_65,N_2828,N_2431);
nor UO_66 (O_66,N_2360,N_2747);
nand UO_67 (O_67,N_2699,N_2634);
and UO_68 (O_68,N_2928,N_2580);
xnor UO_69 (O_69,N_2342,N_2529);
or UO_70 (O_70,N_2926,N_2356);
nor UO_71 (O_71,N_2258,N_2764);
or UO_72 (O_72,N_2626,N_2652);
xnor UO_73 (O_73,N_2279,N_2618);
nor UO_74 (O_74,N_2633,N_2963);
xnor UO_75 (O_75,N_2545,N_2668);
nand UO_76 (O_76,N_2363,N_2254);
nor UO_77 (O_77,N_2690,N_2421);
and UO_78 (O_78,N_2815,N_2811);
or UO_79 (O_79,N_2436,N_2721);
and UO_80 (O_80,N_2880,N_2922);
nand UO_81 (O_81,N_2827,N_2461);
and UO_82 (O_82,N_2788,N_2642);
nor UO_83 (O_83,N_2257,N_2989);
and UO_84 (O_84,N_2494,N_2304);
and UO_85 (O_85,N_2868,N_2495);
nor UO_86 (O_86,N_2361,N_2574);
and UO_87 (O_87,N_2352,N_2532);
or UO_88 (O_88,N_2252,N_2872);
and UO_89 (O_89,N_2903,N_2923);
nor UO_90 (O_90,N_2727,N_2299);
nor UO_91 (O_91,N_2286,N_2599);
nor UO_92 (O_92,N_2712,N_2368);
nand UO_93 (O_93,N_2554,N_2412);
and UO_94 (O_94,N_2566,N_2859);
nand UO_95 (O_95,N_2965,N_2914);
or UO_96 (O_96,N_2591,N_2867);
xnor UO_97 (O_97,N_2913,N_2497);
xor UO_98 (O_98,N_2794,N_2973);
or UO_99 (O_99,N_2862,N_2520);
nor UO_100 (O_100,N_2621,N_2755);
nor UO_101 (O_101,N_2949,N_2732);
xor UO_102 (O_102,N_2284,N_2250);
or UO_103 (O_103,N_2354,N_2387);
nor UO_104 (O_104,N_2806,N_2977);
nor UO_105 (O_105,N_2722,N_2594);
nand UO_106 (O_106,N_2417,N_2758);
nor UO_107 (O_107,N_2841,N_2911);
xnor UO_108 (O_108,N_2742,N_2766);
nand UO_109 (O_109,N_2362,N_2689);
nand UO_110 (O_110,N_2987,N_2939);
or UO_111 (O_111,N_2468,N_2705);
nor UO_112 (O_112,N_2968,N_2466);
or UO_113 (O_113,N_2677,N_2573);
nor UO_114 (O_114,N_2647,N_2364);
or UO_115 (O_115,N_2300,N_2894);
nand UO_116 (O_116,N_2569,N_2694);
nor UO_117 (O_117,N_2887,N_2521);
and UO_118 (O_118,N_2505,N_2260);
or UO_119 (O_119,N_2256,N_2340);
and UO_120 (O_120,N_2948,N_2533);
or UO_121 (O_121,N_2482,N_2799);
and UO_122 (O_122,N_2980,N_2617);
or UO_123 (O_123,N_2940,N_2374);
xnor UO_124 (O_124,N_2288,N_2555);
nand UO_125 (O_125,N_2737,N_2874);
nor UO_126 (O_126,N_2696,N_2435);
nor UO_127 (O_127,N_2263,N_2653);
xnor UO_128 (O_128,N_2637,N_2635);
and UO_129 (O_129,N_2411,N_2623);
nor UO_130 (O_130,N_2519,N_2331);
and UO_131 (O_131,N_2377,N_2480);
nand UO_132 (O_132,N_2746,N_2601);
and UO_133 (O_133,N_2514,N_2661);
or UO_134 (O_134,N_2498,N_2433);
or UO_135 (O_135,N_2271,N_2516);
and UO_136 (O_136,N_2953,N_2541);
or UO_137 (O_137,N_2927,N_2587);
and UO_138 (O_138,N_2547,N_2518);
xor UO_139 (O_139,N_2455,N_2345);
nor UO_140 (O_140,N_2511,N_2849);
and UO_141 (O_141,N_2564,N_2359);
nand UO_142 (O_142,N_2959,N_2982);
nand UO_143 (O_143,N_2274,N_2990);
and UO_144 (O_144,N_2743,N_2768);
nand UO_145 (O_145,N_2845,N_2683);
xor UO_146 (O_146,N_2631,N_2583);
nand UO_147 (O_147,N_2763,N_2606);
or UO_148 (O_148,N_2477,N_2809);
and UO_149 (O_149,N_2383,N_2679);
nand UO_150 (O_150,N_2667,N_2438);
and UO_151 (O_151,N_2607,N_2572);
xnor UO_152 (O_152,N_2724,N_2434);
or UO_153 (O_153,N_2835,N_2920);
or UO_154 (O_154,N_2728,N_2649);
or UO_155 (O_155,N_2884,N_2998);
nand UO_156 (O_156,N_2399,N_2351);
nand UO_157 (O_157,N_2648,N_2616);
nor UO_158 (O_158,N_2389,N_2723);
and UO_159 (O_159,N_2865,N_2403);
xnor UO_160 (O_160,N_2325,N_2673);
xor UO_161 (O_161,N_2357,N_2784);
nand UO_162 (O_162,N_2253,N_2950);
xnor UO_163 (O_163,N_2537,N_2316);
nand UO_164 (O_164,N_2287,N_2264);
or UO_165 (O_165,N_2442,N_2675);
or UO_166 (O_166,N_2330,N_2404);
and UO_167 (O_167,N_2836,N_2629);
and UO_168 (O_168,N_2639,N_2744);
and UO_169 (O_169,N_2292,N_2979);
or UO_170 (O_170,N_2955,N_2850);
nand UO_171 (O_171,N_2889,N_2714);
and UO_172 (O_172,N_2645,N_2686);
and UO_173 (O_173,N_2822,N_2774);
nand UO_174 (O_174,N_2906,N_2932);
and UO_175 (O_175,N_2834,N_2405);
xor UO_176 (O_176,N_2456,N_2589);
nor UO_177 (O_177,N_2921,N_2586);
nand UO_178 (O_178,N_2643,N_2941);
nand UO_179 (O_179,N_2496,N_2853);
nand UO_180 (O_180,N_2901,N_2692);
xnor UO_181 (O_181,N_2994,N_2327);
nor UO_182 (O_182,N_2372,N_2761);
nand UO_183 (O_183,N_2954,N_2646);
or UO_184 (O_184,N_2678,N_2820);
xnor UO_185 (O_185,N_2475,N_2934);
nor UO_186 (O_186,N_2871,N_2797);
nand UO_187 (O_187,N_2995,N_2584);
xnor UO_188 (O_188,N_2603,N_2269);
or UO_189 (O_189,N_2680,N_2311);
or UO_190 (O_190,N_2321,N_2447);
xnor UO_191 (O_191,N_2512,N_2688);
xnor UO_192 (O_192,N_2757,N_2996);
nor UO_193 (O_193,N_2825,N_2481);
and UO_194 (O_194,N_2937,N_2733);
and UO_195 (O_195,N_2796,N_2701);
or UO_196 (O_196,N_2823,N_2709);
nor UO_197 (O_197,N_2333,N_2319);
or UO_198 (O_198,N_2510,N_2613);
and UO_199 (O_199,N_2410,N_2842);
and UO_200 (O_200,N_2343,N_2759);
nor UO_201 (O_201,N_2879,N_2430);
xnor UO_202 (O_202,N_2401,N_2588);
nand UO_203 (O_203,N_2283,N_2483);
or UO_204 (O_204,N_2315,N_2812);
nor UO_205 (O_205,N_2935,N_2720);
or UO_206 (O_206,N_2783,N_2726);
and UO_207 (O_207,N_2813,N_2878);
and UO_208 (O_208,N_2281,N_2294);
nor UO_209 (O_209,N_2407,N_2272);
nor UO_210 (O_210,N_2393,N_2339);
or UO_211 (O_211,N_2844,N_2332);
and UO_212 (O_212,N_2729,N_2422);
and UO_213 (O_213,N_2296,N_2365);
xnor UO_214 (O_214,N_2527,N_2305);
nor UO_215 (O_215,N_2457,N_2307);
and UO_216 (O_216,N_2816,N_2379);
nor UO_217 (O_217,N_2682,N_2999);
and UO_218 (O_218,N_2611,N_2888);
or UO_219 (O_219,N_2875,N_2385);
and UO_220 (O_220,N_2349,N_2355);
nor UO_221 (O_221,N_2890,N_2902);
nor UO_222 (O_222,N_2655,N_2930);
and UO_223 (O_223,N_2899,N_2944);
xnor UO_224 (O_224,N_2802,N_2392);
or UO_225 (O_225,N_2268,N_2553);
and UO_226 (O_226,N_2334,N_2993);
nor UO_227 (O_227,N_2549,N_2961);
nand UO_228 (O_228,N_2567,N_2751);
nor UO_229 (O_229,N_2703,N_2830);
nand UO_230 (O_230,N_2685,N_2706);
and UO_231 (O_231,N_2267,N_2719);
xor UO_232 (O_232,N_2938,N_2531);
and UO_233 (O_233,N_2947,N_2966);
and UO_234 (O_234,N_2777,N_2870);
nor UO_235 (O_235,N_2876,N_2915);
and UO_236 (O_236,N_2449,N_2396);
and UO_237 (O_237,N_2873,N_2620);
or UO_238 (O_238,N_2306,N_2310);
or UO_239 (O_239,N_2577,N_2897);
and UO_240 (O_240,N_2530,N_2917);
nand UO_241 (O_241,N_2418,N_2717);
xor UO_242 (O_242,N_2259,N_2317);
nand UO_243 (O_243,N_2423,N_2563);
or UO_244 (O_244,N_2439,N_2443);
nand UO_245 (O_245,N_2749,N_2658);
nand UO_246 (O_246,N_2925,N_2627);
xor UO_247 (O_247,N_2581,N_2991);
or UO_248 (O_248,N_2585,N_2273);
or UO_249 (O_249,N_2908,N_2793);
or UO_250 (O_250,N_2976,N_2795);
nand UO_251 (O_251,N_2885,N_2988);
or UO_252 (O_252,N_2662,N_2708);
or UO_253 (O_253,N_2323,N_2628);
and UO_254 (O_254,N_2756,N_2697);
nor UO_255 (O_255,N_2597,N_2409);
nor UO_256 (O_256,N_2632,N_2302);
or UO_257 (O_257,N_2951,N_2650);
nand UO_258 (O_258,N_2526,N_2893);
and UO_259 (O_259,N_2910,N_2265);
and UO_260 (O_260,N_2450,N_2610);
nor UO_261 (O_261,N_2501,N_2326);
nor UO_262 (O_262,N_2543,N_2491);
nor UO_263 (O_263,N_2416,N_2490);
nand UO_264 (O_264,N_2942,N_2295);
nand UO_265 (O_265,N_2710,N_2500);
nand UO_266 (O_266,N_2817,N_2413);
nor UO_267 (O_267,N_2382,N_2956);
nand UO_268 (O_268,N_2984,N_2437);
or UO_269 (O_269,N_2301,N_2504);
and UO_270 (O_270,N_2919,N_2659);
or UO_271 (O_271,N_2900,N_2839);
and UO_272 (O_272,N_2905,N_2329);
or UO_273 (O_273,N_2324,N_2388);
or UO_274 (O_274,N_2776,N_2381);
or UO_275 (O_275,N_2909,N_2440);
and UO_276 (O_276,N_2943,N_2560);
and UO_277 (O_277,N_2462,N_2641);
nand UO_278 (O_278,N_2312,N_2453);
nand UO_279 (O_279,N_2303,N_2313);
nand UO_280 (O_280,N_2760,N_2592);
and UO_281 (O_281,N_2964,N_2904);
or UO_282 (O_282,N_2852,N_2857);
nor UO_283 (O_283,N_2471,N_2539);
and UO_284 (O_284,N_2366,N_2467);
or UO_285 (O_285,N_2593,N_2275);
and UO_286 (O_286,N_2320,N_2856);
nand UO_287 (O_287,N_2819,N_2454);
and UO_288 (O_288,N_2270,N_2297);
xnor UO_289 (O_289,N_2426,N_2945);
or UO_290 (O_290,N_2314,N_2493);
nand UO_291 (O_291,N_2786,N_2542);
nand UO_292 (O_292,N_2748,N_2432);
nor UO_293 (O_293,N_2557,N_2266);
or UO_294 (O_294,N_2538,N_2838);
nor UO_295 (O_295,N_2716,N_2798);
and UO_296 (O_296,N_2933,N_2348);
and UO_297 (O_297,N_2261,N_2509);
nor UO_298 (O_298,N_2485,N_2290);
xnor UO_299 (O_299,N_2513,N_2395);
or UO_300 (O_300,N_2282,N_2448);
or UO_301 (O_301,N_2470,N_2740);
nand UO_302 (O_302,N_2318,N_2981);
and UO_303 (O_303,N_2548,N_2384);
and UO_304 (O_304,N_2781,N_2337);
and UO_305 (O_305,N_2735,N_2858);
and UO_306 (O_306,N_2969,N_2877);
nand UO_307 (O_307,N_2420,N_2309);
nor UO_308 (O_308,N_2814,N_2285);
and UO_309 (O_309,N_2619,N_2595);
or UO_310 (O_310,N_2832,N_2821);
and UO_311 (O_311,N_2785,N_2752);
xnor UO_312 (O_312,N_2419,N_2986);
nand UO_313 (O_313,N_2912,N_2458);
nor UO_314 (O_314,N_2967,N_2474);
nand UO_315 (O_315,N_2674,N_2550);
or UO_316 (O_316,N_2779,N_2369);
xor UO_317 (O_317,N_2753,N_2792);
nand UO_318 (O_318,N_2428,N_2801);
or UO_319 (O_319,N_2918,N_2376);
nor UO_320 (O_320,N_2924,N_2670);
nor UO_321 (O_321,N_2672,N_2638);
or UO_322 (O_322,N_2579,N_2540);
or UO_323 (O_323,N_2739,N_2829);
nand UO_324 (O_324,N_2578,N_2517);
nor UO_325 (O_325,N_2782,N_2605);
nand UO_326 (O_326,N_2736,N_2487);
or UO_327 (O_327,N_2681,N_2789);
and UO_328 (O_328,N_2711,N_2803);
and UO_329 (O_329,N_2750,N_2503);
xor UO_330 (O_330,N_2691,N_2575);
nand UO_331 (O_331,N_2775,N_2414);
and UO_332 (O_332,N_2596,N_2745);
and UO_333 (O_333,N_2837,N_2640);
or UO_334 (O_334,N_2624,N_2854);
and UO_335 (O_335,N_2958,N_2765);
and UO_336 (O_336,N_2429,N_2298);
nand UO_337 (O_337,N_2576,N_2656);
and UO_338 (O_338,N_2568,N_2866);
nand UO_339 (O_339,N_2535,N_2861);
and UO_340 (O_340,N_2551,N_2780);
or UO_341 (O_341,N_2695,N_2424);
nor UO_342 (O_342,N_2734,N_2400);
or UO_343 (O_343,N_2262,N_2406);
nand UO_344 (O_344,N_2353,N_2358);
nor UO_345 (O_345,N_2684,N_2397);
or UO_346 (O_346,N_2846,N_2790);
and UO_347 (O_347,N_2810,N_2276);
nand UO_348 (O_348,N_2347,N_2346);
nand UO_349 (O_349,N_2427,N_2704);
nand UO_350 (O_350,N_2929,N_2322);
nor UO_351 (O_351,N_2523,N_2571);
nor UO_352 (O_352,N_2582,N_2808);
nor UO_353 (O_353,N_2770,N_2754);
or UO_354 (O_354,N_2663,N_2464);
nand UO_355 (O_355,N_2731,N_2598);
and UO_356 (O_356,N_2614,N_2882);
nor UO_357 (O_357,N_2660,N_2669);
nor UO_358 (O_358,N_2278,N_2892);
nand UO_359 (O_359,N_2488,N_2975);
nor UO_360 (O_360,N_2636,N_2506);
nor UO_361 (O_361,N_2970,N_2630);
or UO_362 (O_362,N_2378,N_2730);
or UO_363 (O_363,N_2960,N_2534);
and UO_364 (O_364,N_2398,N_2336);
nand UO_365 (O_365,N_2957,N_2883);
nor UO_366 (O_366,N_2807,N_2486);
nand UO_367 (O_367,N_2952,N_2408);
nand UO_368 (O_368,N_2476,N_2805);
nand UO_369 (O_369,N_2787,N_2522);
nand UO_370 (O_370,N_2552,N_2445);
or UO_371 (O_371,N_2602,N_2791);
nor UO_372 (O_372,N_2451,N_2895);
nor UO_373 (O_373,N_2687,N_2465);
and UO_374 (O_374,N_2891,N_2702);
nor UO_375 (O_375,N_2312,N_2908);
and UO_376 (O_376,N_2333,N_2332);
and UO_377 (O_377,N_2417,N_2870);
or UO_378 (O_378,N_2910,N_2447);
or UO_379 (O_379,N_2415,N_2874);
nand UO_380 (O_380,N_2347,N_2647);
and UO_381 (O_381,N_2476,N_2865);
nor UO_382 (O_382,N_2250,N_2807);
nand UO_383 (O_383,N_2473,N_2880);
or UO_384 (O_384,N_2539,N_2727);
or UO_385 (O_385,N_2574,N_2592);
nor UO_386 (O_386,N_2287,N_2796);
or UO_387 (O_387,N_2926,N_2323);
or UO_388 (O_388,N_2297,N_2291);
and UO_389 (O_389,N_2525,N_2609);
nor UO_390 (O_390,N_2894,N_2701);
or UO_391 (O_391,N_2594,N_2546);
or UO_392 (O_392,N_2441,N_2896);
and UO_393 (O_393,N_2353,N_2508);
or UO_394 (O_394,N_2999,N_2496);
nand UO_395 (O_395,N_2780,N_2600);
and UO_396 (O_396,N_2943,N_2453);
nand UO_397 (O_397,N_2424,N_2812);
xnor UO_398 (O_398,N_2369,N_2268);
nor UO_399 (O_399,N_2255,N_2672);
or UO_400 (O_400,N_2422,N_2483);
or UO_401 (O_401,N_2635,N_2395);
nand UO_402 (O_402,N_2279,N_2952);
nand UO_403 (O_403,N_2836,N_2297);
nand UO_404 (O_404,N_2924,N_2392);
nor UO_405 (O_405,N_2511,N_2615);
nor UO_406 (O_406,N_2809,N_2383);
nor UO_407 (O_407,N_2555,N_2753);
or UO_408 (O_408,N_2411,N_2855);
xor UO_409 (O_409,N_2561,N_2952);
xor UO_410 (O_410,N_2761,N_2282);
nand UO_411 (O_411,N_2736,N_2773);
nand UO_412 (O_412,N_2384,N_2852);
nor UO_413 (O_413,N_2788,N_2834);
xnor UO_414 (O_414,N_2411,N_2254);
or UO_415 (O_415,N_2882,N_2768);
nor UO_416 (O_416,N_2950,N_2910);
nand UO_417 (O_417,N_2252,N_2739);
and UO_418 (O_418,N_2439,N_2618);
and UO_419 (O_419,N_2452,N_2692);
nand UO_420 (O_420,N_2998,N_2314);
nand UO_421 (O_421,N_2266,N_2435);
nor UO_422 (O_422,N_2852,N_2880);
nand UO_423 (O_423,N_2837,N_2976);
and UO_424 (O_424,N_2450,N_2804);
nand UO_425 (O_425,N_2991,N_2499);
nand UO_426 (O_426,N_2732,N_2530);
or UO_427 (O_427,N_2937,N_2986);
nor UO_428 (O_428,N_2997,N_2276);
and UO_429 (O_429,N_2948,N_2952);
and UO_430 (O_430,N_2556,N_2389);
or UO_431 (O_431,N_2977,N_2575);
nand UO_432 (O_432,N_2631,N_2653);
nor UO_433 (O_433,N_2978,N_2346);
xnor UO_434 (O_434,N_2711,N_2658);
nor UO_435 (O_435,N_2870,N_2445);
or UO_436 (O_436,N_2562,N_2750);
nor UO_437 (O_437,N_2674,N_2915);
nor UO_438 (O_438,N_2893,N_2262);
and UO_439 (O_439,N_2539,N_2680);
or UO_440 (O_440,N_2748,N_2993);
xor UO_441 (O_441,N_2883,N_2831);
and UO_442 (O_442,N_2788,N_2745);
nor UO_443 (O_443,N_2632,N_2465);
or UO_444 (O_444,N_2757,N_2506);
nand UO_445 (O_445,N_2592,N_2878);
nand UO_446 (O_446,N_2635,N_2469);
or UO_447 (O_447,N_2617,N_2357);
nand UO_448 (O_448,N_2302,N_2999);
or UO_449 (O_449,N_2837,N_2744);
or UO_450 (O_450,N_2307,N_2738);
and UO_451 (O_451,N_2911,N_2720);
or UO_452 (O_452,N_2456,N_2681);
and UO_453 (O_453,N_2960,N_2623);
xnor UO_454 (O_454,N_2413,N_2359);
nand UO_455 (O_455,N_2971,N_2751);
nor UO_456 (O_456,N_2891,N_2779);
nor UO_457 (O_457,N_2293,N_2879);
xnor UO_458 (O_458,N_2813,N_2647);
nand UO_459 (O_459,N_2820,N_2655);
or UO_460 (O_460,N_2884,N_2816);
and UO_461 (O_461,N_2899,N_2251);
xor UO_462 (O_462,N_2870,N_2725);
and UO_463 (O_463,N_2838,N_2444);
nor UO_464 (O_464,N_2745,N_2522);
nor UO_465 (O_465,N_2418,N_2477);
nand UO_466 (O_466,N_2818,N_2273);
and UO_467 (O_467,N_2606,N_2599);
and UO_468 (O_468,N_2438,N_2738);
nand UO_469 (O_469,N_2370,N_2643);
nand UO_470 (O_470,N_2815,N_2904);
nand UO_471 (O_471,N_2616,N_2282);
and UO_472 (O_472,N_2966,N_2990);
and UO_473 (O_473,N_2571,N_2251);
and UO_474 (O_474,N_2461,N_2607);
nor UO_475 (O_475,N_2297,N_2716);
nor UO_476 (O_476,N_2592,N_2555);
or UO_477 (O_477,N_2553,N_2347);
or UO_478 (O_478,N_2829,N_2774);
nor UO_479 (O_479,N_2683,N_2947);
or UO_480 (O_480,N_2892,N_2950);
xor UO_481 (O_481,N_2276,N_2622);
and UO_482 (O_482,N_2593,N_2671);
nor UO_483 (O_483,N_2973,N_2839);
nand UO_484 (O_484,N_2856,N_2884);
xnor UO_485 (O_485,N_2809,N_2393);
nor UO_486 (O_486,N_2490,N_2263);
nor UO_487 (O_487,N_2779,N_2686);
xor UO_488 (O_488,N_2654,N_2581);
or UO_489 (O_489,N_2659,N_2677);
xnor UO_490 (O_490,N_2342,N_2981);
and UO_491 (O_491,N_2794,N_2910);
and UO_492 (O_492,N_2549,N_2735);
nand UO_493 (O_493,N_2638,N_2943);
and UO_494 (O_494,N_2562,N_2748);
xor UO_495 (O_495,N_2545,N_2312);
and UO_496 (O_496,N_2818,N_2375);
nand UO_497 (O_497,N_2436,N_2277);
nand UO_498 (O_498,N_2278,N_2400);
and UO_499 (O_499,N_2311,N_2384);
endmodule