module basic_750_5000_1000_2_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2511,N_2512,N_2515,N_2516,N_2517,N_2519,N_2520,N_2521,N_2522,N_2525,N_2526,N_2527,N_2528,N_2529,N_2531,N_2533,N_2537,N_2538,N_2539,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2580,N_2581,N_2582,N_2583,N_2585,N_2587,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2601,N_2603,N_2604,N_2606,N_2610,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2623,N_2624,N_2625,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2654,N_2655,N_2656,N_2657,N_2660,N_2661,N_2662,N_2663,N_2664,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2688,N_2689,N_2690,N_2692,N_2694,N_2695,N_2696,N_2698,N_2700,N_2701,N_2702,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2711,N_2713,N_2715,N_2716,N_2717,N_2718,N_2720,N_2721,N_2722,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2739,N_2742,N_2744,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2760,N_2762,N_2763,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2784,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2795,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2813,N_2814,N_2815,N_2816,N_2819,N_2820,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2836,N_2837,N_2838,N_2840,N_2841,N_2842,N_2844,N_2845,N_2846,N_2849,N_2851,N_2852,N_2853,N_2854,N_2855,N_2858,N_2859,N_2861,N_2862,N_2863,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2882,N_2883,N_2887,N_2888,N_2890,N_2892,N_2895,N_2897,N_2898,N_2899,N_2900,N_2901,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2915,N_2916,N_2918,N_2919,N_2921,N_2923,N_2925,N_2926,N_2927,N_2928,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2938,N_2939,N_2940,N_2941,N_2943,N_2944,N_2945,N_2946,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2964,N_2965,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2989,N_2991,N_2992,N_2993,N_2995,N_2998,N_3000,N_3001,N_3003,N_3004,N_3005,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3017,N_3018,N_3020,N_3021,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3047,N_3048,N_3050,N_3053,N_3054,N_3055,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3073,N_3074,N_3075,N_3076,N_3078,N_3079,N_3080,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3120,N_3122,N_3123,N_3124,N_3125,N_3126,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3135,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3149,N_3150,N_3152,N_3154,N_3155,N_3156,N_3158,N_3160,N_3161,N_3162,N_3163,N_3165,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3174,N_3175,N_3177,N_3178,N_3179,N_3181,N_3183,N_3185,N_3187,N_3188,N_3191,N_3192,N_3193,N_3195,N_3198,N_3199,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3214,N_3216,N_3219,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3242,N_3243,N_3244,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3258,N_3259,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3289,N_3290,N_3291,N_3292,N_3293,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3304,N_3305,N_3307,N_3309,N_3310,N_3311,N_3314,N_3315,N_3316,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3359,N_3360,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3392,N_3393,N_3394,N_3395,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3431,N_3432,N_3433,N_3434,N_3436,N_3437,N_3439,N_3440,N_3441,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3451,N_3452,N_3453,N_3455,N_3456,N_3458,N_3460,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3490,N_3491,N_3492,N_3493,N_3495,N_3497,N_3499,N_3500,N_3502,N_3503,N_3505,N_3506,N_3507,N_3508,N_3510,N_3511,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3533,N_3534,N_3536,N_3537,N_3538,N_3539,N_3540,N_3542,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3551,N_3552,N_3553,N_3554,N_3556,N_3557,N_3558,N_3559,N_3560,N_3562,N_3563,N_3565,N_3566,N_3567,N_3568,N_3569,N_3571,N_3572,N_3574,N_3576,N_3577,N_3579,N_3582,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3608,N_3610,N_3611,N_3612,N_3615,N_3616,N_3617,N_3620,N_3621,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3636,N_3638,N_3639,N_3641,N_3642,N_3643,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3662,N_3663,N_3664,N_3666,N_3667,N_3670,N_3671,N_3672,N_3673,N_3676,N_3677,N_3678,N_3679,N_3680,N_3682,N_3683,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3712,N_3713,N_3714,N_3716,N_3717,N_3719,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3734,N_3735,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3745,N_3746,N_3748,N_3749,N_3751,N_3752,N_3754,N_3755,N_3756,N_3757,N_3759,N_3760,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3782,N_3785,N_3786,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3796,N_3797,N_3800,N_3801,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3836,N_3837,N_3838,N_3841,N_3842,N_3843,N_3844,N_3845,N_3848,N_3850,N_3851,N_3854,N_3855,N_3856,N_3857,N_3858,N_3862,N_3863,N_3864,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3880,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3889,N_3890,N_3891,N_3892,N_3893,N_3895,N_3896,N_3899,N_3900,N_3901,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3918,N_3919,N_3920,N_3921,N_3922,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3946,N_3947,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3974,N_3975,N_3976,N_3978,N_3980,N_3981,N_3982,N_3984,N_3986,N_3987,N_3988,N_3989,N_3990,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4001,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4013,N_4014,N_4015,N_4016,N_4018,N_4019,N_4021,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4037,N_4039,N_4040,N_4042,N_4044,N_4045,N_4048,N_4049,N_4050,N_4051,N_4052,N_4054,N_4055,N_4056,N_4057,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4067,N_4068,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4086,N_4087,N_4089,N_4090,N_4093,N_4095,N_4096,N_4097,N_4099,N_4102,N_4103,N_4105,N_4106,N_4107,N_4108,N_4109,N_4113,N_4114,N_4115,N_4116,N_4118,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4129,N_4130,N_4131,N_4132,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4141,N_4143,N_4144,N_4145,N_4146,N_4147,N_4149,N_4150,N_4151,N_4154,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4208,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4220,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4231,N_4232,N_4233,N_4234,N_4235,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4249,N_4250,N_4252,N_4253,N_4254,N_4257,N_4258,N_4259,N_4260,N_4262,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4274,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4283,N_4284,N_4285,N_4287,N_4289,N_4290,N_4291,N_4292,N_4293,N_4295,N_4296,N_4297,N_4299,N_4301,N_4302,N_4304,N_4305,N_4306,N_4307,N_4308,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4321,N_4322,N_4323,N_4324,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4361,N_4362,N_4363,N_4364,N_4366,N_4368,N_4369,N_4371,N_4372,N_4373,N_4374,N_4376,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4390,N_4391,N_4392,N_4393,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4414,N_4415,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4426,N_4427,N_4428,N_4430,N_4431,N_4432,N_4433,N_4435,N_4436,N_4437,N_4438,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4491,N_4492,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4503,N_4504,N_4506,N_4508,N_4509,N_4510,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4528,N_4529,N_4531,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4558,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4568,N_4569,N_4570,N_4571,N_4573,N_4576,N_4577,N_4579,N_4581,N_4583,N_4585,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4614,N_4616,N_4617,N_4618,N_4621,N_4622,N_4624,N_4625,N_4626,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4640,N_4641,N_4643,N_4644,N_4646,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4727,N_4728,N_4729,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4771,N_4773,N_4774,N_4776,N_4778,N_4779,N_4781,N_4782,N_4784,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4799,N_4800,N_4801,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4877,N_4878,N_4879,N_4880,N_4882,N_4883,N_4884,N_4885,N_4886,N_4888,N_4889,N_4892,N_4894,N_4895,N_4896,N_4898,N_4899,N_4900,N_4901,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4944,N_4945,N_4947,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4990,N_4991,N_4992,N_4993,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_456,In_80);
or U1 (N_1,In_634,In_184);
nand U2 (N_2,In_330,In_600);
nor U3 (N_3,In_578,In_566);
and U4 (N_4,In_475,In_421);
and U5 (N_5,In_12,In_350);
or U6 (N_6,In_464,In_409);
nand U7 (N_7,In_30,In_270);
and U8 (N_8,In_511,In_316);
nand U9 (N_9,In_549,In_144);
nor U10 (N_10,In_478,In_439);
nand U11 (N_11,In_117,In_177);
and U12 (N_12,In_404,In_325);
nor U13 (N_13,In_708,In_322);
nor U14 (N_14,In_70,In_294);
and U15 (N_15,In_748,In_237);
and U16 (N_16,In_596,In_565);
and U17 (N_17,In_682,In_164);
nand U18 (N_18,In_704,In_429);
or U19 (N_19,In_558,In_283);
and U20 (N_20,In_740,In_631);
or U21 (N_21,In_538,In_366);
or U22 (N_22,In_393,In_696);
and U23 (N_23,In_642,In_155);
and U24 (N_24,In_746,In_373);
nor U25 (N_25,In_611,In_423);
or U26 (N_26,In_305,In_24);
nand U27 (N_27,In_383,In_725);
nor U28 (N_28,In_365,In_715);
and U29 (N_29,In_479,In_238);
or U30 (N_30,In_562,In_138);
and U31 (N_31,In_355,In_34);
nand U32 (N_32,In_13,In_204);
and U33 (N_33,In_339,In_341);
and U34 (N_34,In_85,In_382);
nor U35 (N_35,In_59,In_347);
nor U36 (N_36,In_664,In_326);
and U37 (N_37,In_688,In_160);
nor U38 (N_38,In_180,In_198);
nor U39 (N_39,In_47,In_399);
or U40 (N_40,In_466,In_335);
xnor U41 (N_41,In_497,In_361);
and U42 (N_42,In_287,In_502);
or U43 (N_43,In_581,In_81);
nor U44 (N_44,In_469,In_73);
or U45 (N_45,In_467,In_481);
and U46 (N_46,In_575,In_582);
and U47 (N_47,In_319,In_328);
and U48 (N_48,In_710,In_302);
or U49 (N_49,In_211,In_641);
nand U50 (N_50,In_33,In_541);
or U51 (N_51,In_591,In_156);
or U52 (N_52,In_665,In_118);
nor U53 (N_53,In_52,In_526);
nand U54 (N_54,In_470,In_132);
or U55 (N_55,In_114,In_709);
nand U56 (N_56,In_245,In_711);
nand U57 (N_57,In_419,In_197);
or U58 (N_58,In_308,In_610);
or U59 (N_59,In_430,In_66);
or U60 (N_60,In_327,In_720);
nor U61 (N_61,In_233,In_681);
and U62 (N_62,In_395,In_552);
or U63 (N_63,In_141,In_220);
nand U64 (N_64,In_364,In_391);
nor U65 (N_65,In_62,In_465);
nand U66 (N_66,In_724,In_605);
nand U67 (N_67,In_256,In_97);
and U68 (N_68,In_250,In_677);
nand U69 (N_69,In_309,In_719);
or U70 (N_70,In_252,In_445);
or U71 (N_71,In_574,In_560);
and U72 (N_72,In_263,In_153);
or U73 (N_73,In_448,In_49);
or U74 (N_74,In_647,In_196);
or U75 (N_75,In_277,In_441);
nand U76 (N_76,In_299,In_546);
nand U77 (N_77,In_290,In_1);
and U78 (N_78,In_679,In_346);
and U79 (N_79,In_446,In_616);
and U80 (N_80,In_593,In_95);
and U81 (N_81,In_267,In_480);
or U82 (N_82,In_504,In_225);
nor U83 (N_83,In_45,In_154);
and U84 (N_84,In_743,In_654);
nand U85 (N_85,In_310,In_103);
or U86 (N_86,In_385,In_8);
nor U87 (N_87,In_272,In_730);
nor U88 (N_88,In_337,In_203);
nand U89 (N_89,In_99,In_374);
nand U90 (N_90,In_676,In_656);
nand U91 (N_91,In_78,In_608);
and U92 (N_92,In_63,In_592);
or U93 (N_93,In_249,In_317);
nand U94 (N_94,In_105,In_392);
and U95 (N_95,In_18,In_559);
or U96 (N_96,In_408,In_259);
nor U97 (N_97,In_614,In_500);
or U98 (N_98,In_617,In_300);
nor U99 (N_99,In_274,In_334);
and U100 (N_100,In_597,In_555);
or U101 (N_101,In_210,In_28);
and U102 (N_102,In_484,In_396);
nor U103 (N_103,In_88,In_262);
and U104 (N_104,In_749,In_678);
or U105 (N_105,In_472,In_670);
nand U106 (N_106,In_650,In_590);
nand U107 (N_107,In_255,In_453);
nand U108 (N_108,In_459,In_200);
or U109 (N_109,In_166,In_303);
nor U110 (N_110,In_94,In_436);
nand U111 (N_111,In_454,In_266);
nand U112 (N_112,In_473,In_77);
or U113 (N_113,In_110,In_108);
nand U114 (N_114,In_15,In_633);
and U115 (N_115,In_91,In_359);
or U116 (N_116,In_389,In_496);
nand U117 (N_117,In_662,In_655);
or U118 (N_118,In_702,In_434);
or U119 (N_119,In_675,In_433);
xnor U120 (N_120,In_143,In_607);
nand U121 (N_121,In_168,In_673);
nor U122 (N_122,In_147,In_432);
nand U123 (N_123,In_35,In_488);
and U124 (N_124,In_67,In_304);
nand U125 (N_125,In_625,In_747);
nor U126 (N_126,In_525,In_693);
nand U127 (N_127,In_414,In_39);
nand U128 (N_128,In_426,In_142);
nor U129 (N_129,In_276,In_282);
nand U130 (N_130,In_134,In_74);
nor U131 (N_131,In_222,In_589);
or U132 (N_132,In_553,In_544);
or U133 (N_133,In_570,In_742);
nor U134 (N_134,In_289,In_185);
nand U135 (N_135,In_563,In_627);
or U136 (N_136,In_324,In_653);
and U137 (N_137,In_411,In_232);
and U138 (N_138,In_483,In_745);
and U139 (N_139,In_507,In_60);
or U140 (N_140,In_92,In_295);
and U141 (N_141,In_87,In_636);
nand U142 (N_142,In_437,In_182);
nor U143 (N_143,In_506,In_292);
or U144 (N_144,In_619,In_230);
nand U145 (N_145,In_367,In_726);
and U146 (N_146,In_90,In_206);
or U147 (N_147,In_539,In_615);
and U148 (N_148,In_694,In_424);
nor U149 (N_149,In_447,In_260);
nor U150 (N_150,In_714,In_594);
nor U151 (N_151,In_491,In_509);
nor U152 (N_152,In_638,In_146);
nand U153 (N_153,In_435,In_588);
or U154 (N_154,In_343,In_699);
or U155 (N_155,In_229,In_273);
nand U156 (N_156,In_4,In_712);
xor U157 (N_157,In_19,In_557);
or U158 (N_158,In_519,In_21);
nor U159 (N_159,In_207,In_264);
nor U160 (N_160,In_79,In_666);
and U161 (N_161,In_58,In_318);
nand U162 (N_162,In_425,In_75);
or U163 (N_163,In_518,In_111);
nor U164 (N_164,In_417,In_129);
and U165 (N_165,In_734,In_457);
or U166 (N_166,In_629,In_116);
nor U167 (N_167,In_195,In_162);
or U168 (N_168,In_394,In_126);
nor U169 (N_169,In_234,In_461);
and U170 (N_170,In_668,In_612);
nand U171 (N_171,In_208,In_415);
or U172 (N_172,In_698,In_214);
or U173 (N_173,In_284,In_165);
or U174 (N_174,In_57,In_577);
or U175 (N_175,In_199,In_450);
and U176 (N_176,In_246,In_455);
or U177 (N_177,In_6,In_556);
nand U178 (N_178,In_528,In_191);
nand U179 (N_179,In_201,In_586);
or U180 (N_180,In_43,In_727);
and U181 (N_181,In_223,In_351);
nand U182 (N_182,In_489,In_72);
or U183 (N_183,In_689,In_10);
nor U184 (N_184,In_384,In_651);
and U185 (N_185,In_306,In_236);
or U186 (N_186,In_661,In_713);
nor U187 (N_187,In_427,In_550);
nor U188 (N_188,In_375,In_301);
nand U189 (N_189,In_523,In_127);
and U190 (N_190,In_342,In_368);
and U191 (N_191,In_104,In_603);
nor U192 (N_192,In_169,In_29);
nor U193 (N_193,In_545,In_51);
and U194 (N_194,In_499,In_498);
or U195 (N_195,In_329,In_529);
or U196 (N_196,In_280,In_397);
nor U197 (N_197,In_352,In_44);
or U198 (N_198,In_537,In_171);
or U199 (N_199,In_205,In_505);
nand U200 (N_200,In_403,In_377);
or U201 (N_201,In_468,In_27);
nand U202 (N_202,In_371,In_86);
nor U203 (N_203,In_579,In_84);
nand U204 (N_204,In_400,In_293);
nor U205 (N_205,In_254,In_321);
or U206 (N_206,In_93,In_173);
and U207 (N_207,In_422,In_490);
nand U208 (N_208,In_744,In_46);
or U209 (N_209,In_438,In_644);
or U210 (N_210,In_41,In_444);
and U211 (N_211,In_120,In_569);
nor U212 (N_212,In_109,In_733);
nor U213 (N_213,In_700,In_100);
nand U214 (N_214,In_542,In_248);
nand U215 (N_215,In_189,In_370);
nor U216 (N_216,In_691,In_244);
and U217 (N_217,In_215,In_738);
nor U218 (N_218,In_703,In_40);
and U219 (N_219,In_548,In_50);
nand U220 (N_220,In_261,In_663);
nor U221 (N_221,In_431,In_618);
nor U222 (N_222,In_729,In_452);
and U223 (N_223,In_227,In_463);
or U224 (N_224,In_561,In_279);
or U225 (N_225,In_406,In_163);
and U226 (N_226,In_707,In_64);
nand U227 (N_227,In_551,In_42);
nor U228 (N_228,In_344,In_626);
and U229 (N_229,In_621,In_407);
nor U230 (N_230,In_648,In_536);
nand U231 (N_231,In_428,In_543);
nor U232 (N_232,In_25,In_535);
and U233 (N_233,In_606,In_209);
or U234 (N_234,In_218,In_363);
or U235 (N_235,In_333,In_482);
or U236 (N_236,In_649,In_531);
nor U237 (N_237,In_458,In_674);
and U238 (N_238,In_735,In_130);
and U239 (N_239,In_736,In_721);
or U240 (N_240,In_567,In_336);
nand U241 (N_241,In_686,In_136);
or U242 (N_242,In_486,In_349);
and U243 (N_243,In_96,In_386);
nand U244 (N_244,In_513,In_669);
or U245 (N_245,In_83,In_20);
and U246 (N_246,In_247,In_658);
or U247 (N_247,In_26,In_362);
nand U248 (N_248,In_119,In_172);
nor U249 (N_249,In_583,In_281);
and U250 (N_250,In_253,In_297);
nand U251 (N_251,In_356,In_512);
nand U252 (N_252,In_604,In_573);
or U253 (N_253,In_240,In_106);
nand U254 (N_254,In_527,In_151);
nor U255 (N_255,In_540,In_313);
or U256 (N_256,In_741,In_285);
nand U257 (N_257,In_102,In_474);
or U258 (N_258,In_671,In_471);
or U259 (N_259,In_381,In_599);
nor U260 (N_260,In_320,In_683);
nand U261 (N_261,In_503,In_170);
or U262 (N_262,In_9,In_271);
and U263 (N_263,In_69,In_192);
or U264 (N_264,In_216,In_521);
nand U265 (N_265,In_620,In_652);
or U266 (N_266,In_65,In_379);
nor U267 (N_267,In_728,In_659);
or U268 (N_268,In_167,In_722);
nand U269 (N_269,In_113,In_242);
or U270 (N_270,In_495,In_572);
and U271 (N_271,In_487,In_135);
and U272 (N_272,In_133,In_493);
nor U273 (N_273,In_657,In_98);
or U274 (N_274,In_139,In_646);
and U275 (N_275,In_128,In_291);
and U276 (N_276,In_0,In_585);
or U277 (N_277,In_358,In_32);
and U278 (N_278,In_522,In_315);
nand U279 (N_279,In_732,In_485);
nor U280 (N_280,In_524,In_378);
nor U281 (N_281,In_413,In_462);
or U282 (N_282,In_388,In_137);
xnor U283 (N_283,In_150,In_265);
and U284 (N_284,In_82,In_451);
and U285 (N_285,In_576,In_161);
nand U286 (N_286,In_632,In_178);
nand U287 (N_287,In_348,In_534);
nand U288 (N_288,In_194,In_76);
nor U289 (N_289,In_517,In_251);
nand U290 (N_290,In_739,In_22);
or U291 (N_291,In_390,In_122);
and U292 (N_292,In_323,In_449);
or U293 (N_293,In_17,In_357);
and U294 (N_294,In_213,In_241);
and U295 (N_295,In_623,In_157);
nor U296 (N_296,In_258,In_152);
xnor U297 (N_297,In_376,In_492);
and U298 (N_298,In_602,In_369);
nand U299 (N_299,In_420,In_48);
and U300 (N_300,In_723,In_145);
or U301 (N_301,In_533,In_38);
and U302 (N_302,In_442,In_54);
or U303 (N_303,In_514,In_360);
and U304 (N_304,In_460,In_416);
nor U305 (N_305,In_697,In_212);
nand U306 (N_306,In_554,In_7);
nand U307 (N_307,In_547,In_55);
and U308 (N_308,In_183,In_532);
nor U309 (N_309,In_188,In_598);
and U310 (N_310,In_121,In_68);
and U311 (N_311,In_140,In_3);
nor U312 (N_312,In_193,In_692);
nand U313 (N_313,In_508,In_476);
nand U314 (N_314,In_418,In_5);
nor U315 (N_315,In_338,In_387);
nor U316 (N_316,In_401,In_667);
nand U317 (N_317,In_37,In_187);
nand U318 (N_318,In_53,In_701);
nand U319 (N_319,In_190,In_181);
nand U320 (N_320,In_685,In_690);
or U321 (N_321,In_202,In_645);
nand U322 (N_322,In_717,In_221);
nor U323 (N_323,In_672,In_584);
nand U324 (N_324,In_737,In_515);
or U325 (N_325,In_307,In_695);
or U326 (N_326,In_159,In_115);
and U327 (N_327,In_501,In_345);
nor U328 (N_328,In_71,In_568);
or U329 (N_329,In_36,In_2);
or U330 (N_330,In_148,In_56);
nand U331 (N_331,In_706,In_16);
nor U332 (N_332,In_286,In_175);
nand U333 (N_333,In_372,In_516);
or U334 (N_334,In_530,In_520);
or U335 (N_335,In_298,In_410);
nand U336 (N_336,In_219,In_124);
or U337 (N_337,In_186,In_257);
or U338 (N_338,In_718,In_235);
nor U339 (N_339,In_217,In_331);
or U340 (N_340,In_624,In_23);
nor U341 (N_341,In_680,In_402);
nor U342 (N_342,In_311,In_243);
and U343 (N_343,In_564,In_231);
and U344 (N_344,In_107,In_443);
nand U345 (N_345,In_123,In_226);
and U346 (N_346,In_101,In_622);
nand U347 (N_347,In_609,In_174);
and U348 (N_348,In_510,In_635);
nor U349 (N_349,In_179,In_353);
nand U350 (N_350,In_288,In_314);
nor U351 (N_351,In_660,In_131);
nor U352 (N_352,In_440,In_239);
or U353 (N_353,In_587,In_494);
and U354 (N_354,In_112,In_176);
nand U355 (N_355,In_412,In_716);
and U356 (N_356,In_354,In_89);
or U357 (N_357,In_224,In_61);
and U358 (N_358,In_268,In_684);
and U359 (N_359,In_731,In_639);
and U360 (N_360,In_628,In_613);
or U361 (N_361,In_687,In_14);
nand U362 (N_362,In_571,In_630);
nand U363 (N_363,In_705,In_278);
nand U364 (N_364,In_405,In_31);
nand U365 (N_365,In_477,In_595);
or U366 (N_366,In_340,In_275);
and U367 (N_367,In_312,In_643);
nand U368 (N_368,In_640,In_125);
or U369 (N_369,In_228,In_332);
or U370 (N_370,In_296,In_398);
nand U371 (N_371,In_601,In_149);
nand U372 (N_372,In_637,In_269);
nand U373 (N_373,In_580,In_11);
or U374 (N_374,In_380,In_158);
and U375 (N_375,In_602,In_59);
nand U376 (N_376,In_649,In_302);
and U377 (N_377,In_394,In_204);
or U378 (N_378,In_298,In_424);
nor U379 (N_379,In_734,In_191);
or U380 (N_380,In_637,In_325);
nand U381 (N_381,In_308,In_731);
and U382 (N_382,In_453,In_340);
and U383 (N_383,In_679,In_503);
and U384 (N_384,In_607,In_574);
or U385 (N_385,In_493,In_155);
nand U386 (N_386,In_602,In_225);
nor U387 (N_387,In_571,In_115);
nand U388 (N_388,In_736,In_636);
nand U389 (N_389,In_94,In_87);
nor U390 (N_390,In_160,In_320);
and U391 (N_391,In_243,In_29);
nor U392 (N_392,In_16,In_131);
nand U393 (N_393,In_539,In_162);
or U394 (N_394,In_523,In_697);
and U395 (N_395,In_44,In_563);
nor U396 (N_396,In_332,In_666);
or U397 (N_397,In_107,In_602);
nor U398 (N_398,In_163,In_207);
nand U399 (N_399,In_412,In_2);
nand U400 (N_400,In_72,In_571);
nand U401 (N_401,In_356,In_441);
nor U402 (N_402,In_330,In_719);
and U403 (N_403,In_271,In_627);
nand U404 (N_404,In_363,In_311);
and U405 (N_405,In_191,In_125);
nand U406 (N_406,In_633,In_654);
or U407 (N_407,In_323,In_476);
or U408 (N_408,In_530,In_51);
and U409 (N_409,In_539,In_707);
nor U410 (N_410,In_301,In_140);
nor U411 (N_411,In_417,In_92);
nand U412 (N_412,In_231,In_309);
nor U413 (N_413,In_481,In_411);
or U414 (N_414,In_545,In_14);
nand U415 (N_415,In_352,In_662);
and U416 (N_416,In_78,In_101);
and U417 (N_417,In_333,In_534);
nor U418 (N_418,In_726,In_730);
and U419 (N_419,In_380,In_655);
or U420 (N_420,In_300,In_738);
or U421 (N_421,In_201,In_416);
or U422 (N_422,In_280,In_90);
or U423 (N_423,In_122,In_153);
or U424 (N_424,In_544,In_304);
and U425 (N_425,In_577,In_253);
or U426 (N_426,In_522,In_279);
nor U427 (N_427,In_230,In_515);
or U428 (N_428,In_205,In_663);
nor U429 (N_429,In_404,In_646);
nor U430 (N_430,In_264,In_557);
nand U431 (N_431,In_158,In_143);
nor U432 (N_432,In_96,In_219);
nor U433 (N_433,In_684,In_524);
and U434 (N_434,In_675,In_316);
nor U435 (N_435,In_178,In_551);
or U436 (N_436,In_738,In_686);
nand U437 (N_437,In_297,In_247);
nand U438 (N_438,In_279,In_364);
and U439 (N_439,In_254,In_214);
nand U440 (N_440,In_27,In_301);
nand U441 (N_441,In_246,In_709);
or U442 (N_442,In_468,In_747);
nor U443 (N_443,In_367,In_653);
and U444 (N_444,In_38,In_407);
nand U445 (N_445,In_373,In_285);
and U446 (N_446,In_474,In_112);
nand U447 (N_447,In_438,In_526);
nor U448 (N_448,In_525,In_83);
nand U449 (N_449,In_157,In_292);
nand U450 (N_450,In_326,In_295);
or U451 (N_451,In_557,In_222);
and U452 (N_452,In_507,In_231);
and U453 (N_453,In_743,In_317);
and U454 (N_454,In_726,In_71);
nand U455 (N_455,In_344,In_607);
or U456 (N_456,In_40,In_245);
nand U457 (N_457,In_326,In_633);
nand U458 (N_458,In_533,In_368);
and U459 (N_459,In_94,In_533);
and U460 (N_460,In_554,In_61);
and U461 (N_461,In_520,In_384);
nor U462 (N_462,In_311,In_295);
nand U463 (N_463,In_483,In_145);
nor U464 (N_464,In_635,In_281);
nand U465 (N_465,In_272,In_245);
and U466 (N_466,In_272,In_68);
and U467 (N_467,In_85,In_464);
and U468 (N_468,In_362,In_173);
nand U469 (N_469,In_67,In_26);
nor U470 (N_470,In_748,In_50);
or U471 (N_471,In_288,In_81);
nor U472 (N_472,In_587,In_392);
or U473 (N_473,In_263,In_467);
and U474 (N_474,In_685,In_505);
or U475 (N_475,In_115,In_503);
and U476 (N_476,In_740,In_588);
nand U477 (N_477,In_715,In_597);
or U478 (N_478,In_652,In_605);
and U479 (N_479,In_312,In_219);
nor U480 (N_480,In_600,In_620);
or U481 (N_481,In_733,In_269);
or U482 (N_482,In_443,In_556);
and U483 (N_483,In_636,In_672);
nand U484 (N_484,In_726,In_104);
nor U485 (N_485,In_656,In_736);
and U486 (N_486,In_0,In_569);
and U487 (N_487,In_235,In_232);
and U488 (N_488,In_612,In_715);
nor U489 (N_489,In_99,In_580);
or U490 (N_490,In_382,In_321);
nand U491 (N_491,In_638,In_194);
or U492 (N_492,In_718,In_82);
or U493 (N_493,In_28,In_123);
or U494 (N_494,In_169,In_408);
or U495 (N_495,In_321,In_549);
nand U496 (N_496,In_698,In_89);
nand U497 (N_497,In_429,In_207);
or U498 (N_498,In_587,In_134);
nand U499 (N_499,In_377,In_714);
or U500 (N_500,In_358,In_556);
nand U501 (N_501,In_290,In_244);
or U502 (N_502,In_443,In_199);
nand U503 (N_503,In_45,In_538);
and U504 (N_504,In_591,In_331);
or U505 (N_505,In_93,In_650);
nand U506 (N_506,In_120,In_151);
or U507 (N_507,In_676,In_692);
nand U508 (N_508,In_34,In_253);
nor U509 (N_509,In_135,In_630);
and U510 (N_510,In_96,In_137);
nand U511 (N_511,In_582,In_373);
nor U512 (N_512,In_118,In_129);
nand U513 (N_513,In_175,In_239);
or U514 (N_514,In_321,In_91);
and U515 (N_515,In_567,In_312);
or U516 (N_516,In_400,In_130);
nor U517 (N_517,In_228,In_450);
nand U518 (N_518,In_404,In_584);
and U519 (N_519,In_452,In_263);
and U520 (N_520,In_470,In_599);
nand U521 (N_521,In_262,In_246);
nand U522 (N_522,In_635,In_388);
or U523 (N_523,In_369,In_687);
nor U524 (N_524,In_486,In_298);
nand U525 (N_525,In_329,In_546);
and U526 (N_526,In_105,In_286);
or U527 (N_527,In_159,In_120);
nand U528 (N_528,In_731,In_165);
and U529 (N_529,In_596,In_189);
nand U530 (N_530,In_6,In_637);
nand U531 (N_531,In_629,In_477);
nor U532 (N_532,In_242,In_669);
or U533 (N_533,In_390,In_319);
nand U534 (N_534,In_165,In_453);
nand U535 (N_535,In_619,In_237);
and U536 (N_536,In_538,In_742);
nand U537 (N_537,In_455,In_254);
or U538 (N_538,In_550,In_535);
nor U539 (N_539,In_645,In_592);
nor U540 (N_540,In_355,In_179);
and U541 (N_541,In_196,In_384);
nor U542 (N_542,In_662,In_161);
nand U543 (N_543,In_598,In_594);
nor U544 (N_544,In_366,In_465);
and U545 (N_545,In_626,In_257);
nand U546 (N_546,In_369,In_584);
nor U547 (N_547,In_421,In_554);
or U548 (N_548,In_449,In_480);
or U549 (N_549,In_229,In_668);
or U550 (N_550,In_481,In_103);
nand U551 (N_551,In_118,In_630);
and U552 (N_552,In_16,In_563);
nand U553 (N_553,In_685,In_448);
nor U554 (N_554,In_699,In_29);
nand U555 (N_555,In_438,In_425);
and U556 (N_556,In_472,In_673);
nor U557 (N_557,In_328,In_182);
nand U558 (N_558,In_5,In_420);
nand U559 (N_559,In_392,In_201);
nand U560 (N_560,In_235,In_304);
nand U561 (N_561,In_703,In_374);
nand U562 (N_562,In_2,In_242);
or U563 (N_563,In_417,In_397);
nand U564 (N_564,In_476,In_605);
and U565 (N_565,In_574,In_509);
or U566 (N_566,In_373,In_607);
nand U567 (N_567,In_465,In_585);
or U568 (N_568,In_565,In_587);
or U569 (N_569,In_320,In_624);
or U570 (N_570,In_164,In_702);
and U571 (N_571,In_656,In_212);
and U572 (N_572,In_738,In_651);
nor U573 (N_573,In_1,In_172);
and U574 (N_574,In_570,In_484);
nor U575 (N_575,In_426,In_732);
or U576 (N_576,In_404,In_75);
nor U577 (N_577,In_729,In_119);
nand U578 (N_578,In_274,In_626);
nand U579 (N_579,In_405,In_111);
nor U580 (N_580,In_13,In_513);
nor U581 (N_581,In_586,In_330);
or U582 (N_582,In_402,In_368);
and U583 (N_583,In_255,In_187);
nor U584 (N_584,In_562,In_748);
nor U585 (N_585,In_415,In_682);
or U586 (N_586,In_263,In_115);
nor U587 (N_587,In_9,In_361);
nor U588 (N_588,In_92,In_642);
nand U589 (N_589,In_529,In_202);
nor U590 (N_590,In_174,In_96);
and U591 (N_591,In_521,In_156);
nand U592 (N_592,In_633,In_515);
nor U593 (N_593,In_675,In_175);
nand U594 (N_594,In_34,In_649);
and U595 (N_595,In_488,In_367);
and U596 (N_596,In_492,In_740);
or U597 (N_597,In_712,In_145);
and U598 (N_598,In_338,In_688);
nor U599 (N_599,In_197,In_78);
and U600 (N_600,In_369,In_115);
nand U601 (N_601,In_739,In_392);
and U602 (N_602,In_611,In_229);
nor U603 (N_603,In_727,In_430);
nor U604 (N_604,In_410,In_101);
nand U605 (N_605,In_614,In_31);
and U606 (N_606,In_90,In_472);
nand U607 (N_607,In_252,In_601);
and U608 (N_608,In_202,In_729);
and U609 (N_609,In_425,In_503);
nand U610 (N_610,In_86,In_477);
or U611 (N_611,In_522,In_583);
nor U612 (N_612,In_644,In_380);
nand U613 (N_613,In_348,In_508);
or U614 (N_614,In_480,In_383);
and U615 (N_615,In_396,In_293);
nand U616 (N_616,In_419,In_400);
nor U617 (N_617,In_152,In_621);
or U618 (N_618,In_619,In_148);
nand U619 (N_619,In_720,In_710);
or U620 (N_620,In_524,In_494);
and U621 (N_621,In_44,In_152);
nand U622 (N_622,In_367,In_650);
nor U623 (N_623,In_231,In_236);
and U624 (N_624,In_602,In_455);
nor U625 (N_625,In_3,In_344);
or U626 (N_626,In_649,In_548);
nand U627 (N_627,In_345,In_83);
or U628 (N_628,In_66,In_744);
and U629 (N_629,In_258,In_550);
nand U630 (N_630,In_747,In_195);
or U631 (N_631,In_700,In_380);
and U632 (N_632,In_461,In_697);
nor U633 (N_633,In_67,In_623);
nor U634 (N_634,In_363,In_685);
nand U635 (N_635,In_542,In_479);
nor U636 (N_636,In_692,In_68);
nand U637 (N_637,In_529,In_644);
and U638 (N_638,In_398,In_175);
nand U639 (N_639,In_448,In_263);
or U640 (N_640,In_96,In_621);
or U641 (N_641,In_316,In_486);
nand U642 (N_642,In_234,In_400);
nand U643 (N_643,In_299,In_506);
and U644 (N_644,In_655,In_714);
nor U645 (N_645,In_700,In_140);
and U646 (N_646,In_545,In_42);
or U647 (N_647,In_162,In_428);
and U648 (N_648,In_58,In_338);
or U649 (N_649,In_354,In_269);
and U650 (N_650,In_237,In_712);
nor U651 (N_651,In_628,In_453);
nor U652 (N_652,In_269,In_539);
and U653 (N_653,In_47,In_628);
and U654 (N_654,In_716,In_33);
or U655 (N_655,In_174,In_53);
or U656 (N_656,In_641,In_419);
nor U657 (N_657,In_138,In_281);
and U658 (N_658,In_680,In_255);
and U659 (N_659,In_658,In_692);
or U660 (N_660,In_95,In_85);
and U661 (N_661,In_562,In_445);
nor U662 (N_662,In_590,In_14);
nand U663 (N_663,In_110,In_187);
or U664 (N_664,In_472,In_140);
and U665 (N_665,In_363,In_276);
nor U666 (N_666,In_266,In_497);
nand U667 (N_667,In_141,In_725);
nor U668 (N_668,In_655,In_463);
or U669 (N_669,In_387,In_553);
nor U670 (N_670,In_493,In_302);
or U671 (N_671,In_189,In_290);
nor U672 (N_672,In_161,In_459);
nor U673 (N_673,In_474,In_200);
and U674 (N_674,In_114,In_9);
nor U675 (N_675,In_638,In_136);
or U676 (N_676,In_161,In_615);
or U677 (N_677,In_614,In_298);
and U678 (N_678,In_521,In_71);
nor U679 (N_679,In_596,In_713);
xnor U680 (N_680,In_56,In_469);
and U681 (N_681,In_173,In_290);
nand U682 (N_682,In_316,In_226);
nor U683 (N_683,In_737,In_624);
nor U684 (N_684,In_487,In_26);
and U685 (N_685,In_748,In_391);
nor U686 (N_686,In_179,In_295);
nand U687 (N_687,In_475,In_324);
nor U688 (N_688,In_74,In_340);
nor U689 (N_689,In_534,In_42);
and U690 (N_690,In_318,In_519);
nor U691 (N_691,In_659,In_440);
and U692 (N_692,In_367,In_288);
nor U693 (N_693,In_512,In_43);
or U694 (N_694,In_34,In_310);
nor U695 (N_695,In_167,In_371);
xor U696 (N_696,In_731,In_10);
nand U697 (N_697,In_527,In_349);
nor U698 (N_698,In_632,In_287);
or U699 (N_699,In_623,In_433);
nor U700 (N_700,In_466,In_170);
or U701 (N_701,In_565,In_206);
nor U702 (N_702,In_300,In_440);
nor U703 (N_703,In_116,In_465);
and U704 (N_704,In_397,In_651);
nand U705 (N_705,In_170,In_167);
or U706 (N_706,In_614,In_672);
nand U707 (N_707,In_21,In_284);
and U708 (N_708,In_133,In_673);
nor U709 (N_709,In_531,In_455);
nand U710 (N_710,In_352,In_259);
and U711 (N_711,In_595,In_260);
nand U712 (N_712,In_29,In_216);
nand U713 (N_713,In_138,In_100);
nor U714 (N_714,In_536,In_114);
nand U715 (N_715,In_398,In_724);
and U716 (N_716,In_247,In_468);
or U717 (N_717,In_254,In_88);
or U718 (N_718,In_574,In_438);
or U719 (N_719,In_83,In_188);
nor U720 (N_720,In_247,In_699);
nand U721 (N_721,In_377,In_330);
and U722 (N_722,In_705,In_464);
nand U723 (N_723,In_220,In_676);
and U724 (N_724,In_277,In_32);
and U725 (N_725,In_173,In_673);
and U726 (N_726,In_121,In_568);
or U727 (N_727,In_235,In_295);
nor U728 (N_728,In_319,In_124);
or U729 (N_729,In_37,In_102);
or U730 (N_730,In_154,In_564);
nor U731 (N_731,In_527,In_645);
nand U732 (N_732,In_343,In_605);
nand U733 (N_733,In_184,In_655);
nor U734 (N_734,In_675,In_344);
nand U735 (N_735,In_106,In_335);
nor U736 (N_736,In_207,In_596);
or U737 (N_737,In_631,In_658);
and U738 (N_738,In_329,In_294);
xnor U739 (N_739,In_280,In_309);
and U740 (N_740,In_338,In_7);
or U741 (N_741,In_621,In_743);
nor U742 (N_742,In_614,In_468);
nor U743 (N_743,In_403,In_696);
nand U744 (N_744,In_231,In_407);
nand U745 (N_745,In_219,In_178);
or U746 (N_746,In_352,In_37);
nor U747 (N_747,In_325,In_663);
nand U748 (N_748,In_656,In_520);
and U749 (N_749,In_43,In_403);
nand U750 (N_750,In_302,In_675);
nand U751 (N_751,In_394,In_553);
nor U752 (N_752,In_368,In_300);
and U753 (N_753,In_57,In_237);
and U754 (N_754,In_10,In_246);
nand U755 (N_755,In_335,In_728);
or U756 (N_756,In_284,In_678);
and U757 (N_757,In_156,In_141);
nand U758 (N_758,In_83,In_5);
xnor U759 (N_759,In_67,In_398);
or U760 (N_760,In_175,In_133);
nand U761 (N_761,In_491,In_192);
and U762 (N_762,In_526,In_623);
and U763 (N_763,In_316,In_3);
nor U764 (N_764,In_485,In_96);
nand U765 (N_765,In_673,In_61);
and U766 (N_766,In_215,In_428);
and U767 (N_767,In_707,In_0);
or U768 (N_768,In_367,In_23);
nor U769 (N_769,In_288,In_341);
nor U770 (N_770,In_329,In_264);
and U771 (N_771,In_472,In_634);
nand U772 (N_772,In_202,In_61);
or U773 (N_773,In_355,In_714);
or U774 (N_774,In_377,In_236);
xnor U775 (N_775,In_322,In_390);
and U776 (N_776,In_420,In_217);
and U777 (N_777,In_270,In_408);
nor U778 (N_778,In_493,In_656);
and U779 (N_779,In_548,In_557);
and U780 (N_780,In_125,In_335);
nor U781 (N_781,In_126,In_96);
nand U782 (N_782,In_363,In_737);
nand U783 (N_783,In_356,In_733);
xor U784 (N_784,In_243,In_84);
or U785 (N_785,In_487,In_171);
nor U786 (N_786,In_702,In_245);
and U787 (N_787,In_415,In_154);
nor U788 (N_788,In_377,In_738);
and U789 (N_789,In_559,In_387);
nand U790 (N_790,In_423,In_180);
or U791 (N_791,In_417,In_448);
nand U792 (N_792,In_108,In_280);
or U793 (N_793,In_574,In_403);
nor U794 (N_794,In_151,In_357);
nand U795 (N_795,In_729,In_291);
or U796 (N_796,In_702,In_18);
and U797 (N_797,In_205,In_199);
nor U798 (N_798,In_24,In_221);
and U799 (N_799,In_79,In_698);
nor U800 (N_800,In_270,In_455);
nand U801 (N_801,In_639,In_0);
xnor U802 (N_802,In_27,In_67);
and U803 (N_803,In_21,In_179);
or U804 (N_804,In_586,In_48);
nor U805 (N_805,In_16,In_548);
nor U806 (N_806,In_520,In_500);
or U807 (N_807,In_507,In_89);
and U808 (N_808,In_191,In_548);
nor U809 (N_809,In_451,In_415);
nor U810 (N_810,In_351,In_368);
and U811 (N_811,In_423,In_225);
or U812 (N_812,In_77,In_190);
nand U813 (N_813,In_304,In_299);
nand U814 (N_814,In_246,In_119);
or U815 (N_815,In_491,In_720);
nor U816 (N_816,In_144,In_544);
or U817 (N_817,In_144,In_299);
nor U818 (N_818,In_231,In_184);
nand U819 (N_819,In_591,In_538);
and U820 (N_820,In_477,In_147);
or U821 (N_821,In_285,In_436);
and U822 (N_822,In_180,In_358);
or U823 (N_823,In_638,In_23);
nor U824 (N_824,In_314,In_72);
nor U825 (N_825,In_212,In_489);
nor U826 (N_826,In_180,In_461);
or U827 (N_827,In_695,In_183);
and U828 (N_828,In_609,In_28);
nand U829 (N_829,In_701,In_528);
nand U830 (N_830,In_649,In_255);
nand U831 (N_831,In_121,In_550);
and U832 (N_832,In_103,In_660);
nor U833 (N_833,In_497,In_566);
nand U834 (N_834,In_430,In_636);
and U835 (N_835,In_485,In_729);
and U836 (N_836,In_178,In_563);
or U837 (N_837,In_553,In_529);
or U838 (N_838,In_350,In_80);
nor U839 (N_839,In_630,In_565);
nor U840 (N_840,In_229,In_109);
nor U841 (N_841,In_478,In_350);
or U842 (N_842,In_135,In_155);
nor U843 (N_843,In_344,In_312);
nor U844 (N_844,In_492,In_517);
or U845 (N_845,In_661,In_457);
nor U846 (N_846,In_228,In_535);
and U847 (N_847,In_287,In_276);
nor U848 (N_848,In_673,In_171);
or U849 (N_849,In_249,In_203);
or U850 (N_850,In_684,In_565);
nand U851 (N_851,In_407,In_50);
nand U852 (N_852,In_741,In_697);
or U853 (N_853,In_646,In_602);
or U854 (N_854,In_152,In_354);
and U855 (N_855,In_305,In_282);
and U856 (N_856,In_610,In_618);
and U857 (N_857,In_736,In_385);
and U858 (N_858,In_27,In_510);
or U859 (N_859,In_232,In_58);
nand U860 (N_860,In_740,In_97);
xnor U861 (N_861,In_23,In_307);
nand U862 (N_862,In_517,In_468);
and U863 (N_863,In_433,In_617);
nor U864 (N_864,In_166,In_38);
nor U865 (N_865,In_41,In_686);
and U866 (N_866,In_403,In_607);
xor U867 (N_867,In_598,In_172);
and U868 (N_868,In_204,In_363);
nor U869 (N_869,In_220,In_110);
and U870 (N_870,In_42,In_715);
and U871 (N_871,In_510,In_490);
nand U872 (N_872,In_302,In_102);
nor U873 (N_873,In_563,In_647);
and U874 (N_874,In_363,In_595);
nor U875 (N_875,In_4,In_478);
and U876 (N_876,In_574,In_732);
or U877 (N_877,In_395,In_507);
nand U878 (N_878,In_121,In_79);
nor U879 (N_879,In_55,In_638);
or U880 (N_880,In_669,In_288);
or U881 (N_881,In_118,In_298);
nor U882 (N_882,In_514,In_438);
nand U883 (N_883,In_311,In_672);
or U884 (N_884,In_308,In_168);
or U885 (N_885,In_469,In_139);
and U886 (N_886,In_243,In_392);
or U887 (N_887,In_178,In_489);
nor U888 (N_888,In_291,In_687);
nor U889 (N_889,In_49,In_61);
and U890 (N_890,In_455,In_488);
or U891 (N_891,In_219,In_241);
nand U892 (N_892,In_493,In_373);
nor U893 (N_893,In_126,In_480);
or U894 (N_894,In_317,In_408);
or U895 (N_895,In_363,In_689);
nand U896 (N_896,In_505,In_429);
nand U897 (N_897,In_315,In_717);
nor U898 (N_898,In_560,In_168);
or U899 (N_899,In_689,In_692);
nor U900 (N_900,In_411,In_356);
nor U901 (N_901,In_91,In_250);
or U902 (N_902,In_28,In_57);
and U903 (N_903,In_682,In_683);
nand U904 (N_904,In_288,In_62);
nor U905 (N_905,In_8,In_172);
xor U906 (N_906,In_66,In_189);
nand U907 (N_907,In_267,In_316);
nand U908 (N_908,In_350,In_206);
nor U909 (N_909,In_30,In_156);
nand U910 (N_910,In_402,In_674);
nor U911 (N_911,In_148,In_440);
nand U912 (N_912,In_374,In_457);
nand U913 (N_913,In_26,In_625);
and U914 (N_914,In_72,In_384);
nor U915 (N_915,In_107,In_654);
or U916 (N_916,In_58,In_317);
or U917 (N_917,In_433,In_610);
and U918 (N_918,In_378,In_628);
or U919 (N_919,In_239,In_708);
and U920 (N_920,In_59,In_77);
nand U921 (N_921,In_574,In_323);
and U922 (N_922,In_345,In_551);
or U923 (N_923,In_318,In_483);
nand U924 (N_924,In_657,In_530);
or U925 (N_925,In_483,In_54);
or U926 (N_926,In_737,In_731);
nor U927 (N_927,In_66,In_285);
and U928 (N_928,In_356,In_156);
nor U929 (N_929,In_701,In_256);
nand U930 (N_930,In_293,In_8);
nor U931 (N_931,In_124,In_332);
nand U932 (N_932,In_36,In_744);
or U933 (N_933,In_269,In_644);
or U934 (N_934,In_716,In_638);
nor U935 (N_935,In_546,In_270);
and U936 (N_936,In_333,In_135);
or U937 (N_937,In_736,In_51);
or U938 (N_938,In_252,In_598);
or U939 (N_939,In_303,In_620);
or U940 (N_940,In_346,In_357);
nand U941 (N_941,In_131,In_527);
nor U942 (N_942,In_690,In_56);
or U943 (N_943,In_6,In_314);
nand U944 (N_944,In_39,In_134);
nand U945 (N_945,In_459,In_559);
nand U946 (N_946,In_216,In_509);
and U947 (N_947,In_688,In_198);
nor U948 (N_948,In_725,In_682);
or U949 (N_949,In_554,In_747);
and U950 (N_950,In_589,In_642);
and U951 (N_951,In_391,In_153);
nor U952 (N_952,In_304,In_121);
nor U953 (N_953,In_629,In_705);
nand U954 (N_954,In_119,In_609);
nand U955 (N_955,In_342,In_705);
nor U956 (N_956,In_630,In_126);
nand U957 (N_957,In_457,In_429);
nor U958 (N_958,In_715,In_659);
and U959 (N_959,In_67,In_638);
nand U960 (N_960,In_575,In_563);
nand U961 (N_961,In_425,In_572);
nand U962 (N_962,In_588,In_202);
or U963 (N_963,In_647,In_596);
nand U964 (N_964,In_508,In_182);
and U965 (N_965,In_172,In_614);
nor U966 (N_966,In_608,In_657);
and U967 (N_967,In_371,In_19);
and U968 (N_968,In_529,In_425);
and U969 (N_969,In_18,In_557);
and U970 (N_970,In_233,In_446);
and U971 (N_971,In_541,In_295);
or U972 (N_972,In_674,In_487);
and U973 (N_973,In_146,In_437);
or U974 (N_974,In_537,In_651);
nand U975 (N_975,In_517,In_309);
nand U976 (N_976,In_39,In_357);
or U977 (N_977,In_45,In_532);
xnor U978 (N_978,In_108,In_372);
and U979 (N_979,In_699,In_435);
or U980 (N_980,In_346,In_52);
and U981 (N_981,In_572,In_97);
nor U982 (N_982,In_719,In_431);
nand U983 (N_983,In_290,In_318);
nor U984 (N_984,In_219,In_619);
nand U985 (N_985,In_644,In_351);
and U986 (N_986,In_151,In_58);
and U987 (N_987,In_266,In_273);
or U988 (N_988,In_204,In_749);
nor U989 (N_989,In_164,In_537);
or U990 (N_990,In_306,In_35);
nor U991 (N_991,In_213,In_192);
nand U992 (N_992,In_364,In_363);
or U993 (N_993,In_709,In_732);
nor U994 (N_994,In_278,In_496);
and U995 (N_995,In_588,In_512);
or U996 (N_996,In_698,In_679);
or U997 (N_997,In_367,In_41);
nor U998 (N_998,In_709,In_562);
and U999 (N_999,In_194,In_475);
or U1000 (N_1000,In_734,In_176);
nand U1001 (N_1001,In_477,In_81);
or U1002 (N_1002,In_562,In_85);
and U1003 (N_1003,In_165,In_429);
and U1004 (N_1004,In_310,In_609);
nand U1005 (N_1005,In_580,In_188);
or U1006 (N_1006,In_695,In_614);
and U1007 (N_1007,In_739,In_746);
nor U1008 (N_1008,In_335,In_510);
and U1009 (N_1009,In_169,In_601);
and U1010 (N_1010,In_530,In_153);
nor U1011 (N_1011,In_516,In_189);
nand U1012 (N_1012,In_44,In_476);
nand U1013 (N_1013,In_211,In_275);
and U1014 (N_1014,In_474,In_295);
nor U1015 (N_1015,In_112,In_2);
nor U1016 (N_1016,In_77,In_318);
or U1017 (N_1017,In_684,In_535);
and U1018 (N_1018,In_590,In_496);
or U1019 (N_1019,In_612,In_538);
or U1020 (N_1020,In_698,In_185);
or U1021 (N_1021,In_190,In_371);
nand U1022 (N_1022,In_458,In_76);
or U1023 (N_1023,In_274,In_699);
nor U1024 (N_1024,In_314,In_292);
and U1025 (N_1025,In_317,In_642);
nand U1026 (N_1026,In_163,In_159);
nor U1027 (N_1027,In_218,In_87);
nand U1028 (N_1028,In_408,In_190);
nor U1029 (N_1029,In_193,In_213);
nand U1030 (N_1030,In_141,In_255);
or U1031 (N_1031,In_561,In_362);
nor U1032 (N_1032,In_171,In_305);
and U1033 (N_1033,In_425,In_561);
nand U1034 (N_1034,In_78,In_47);
and U1035 (N_1035,In_694,In_46);
and U1036 (N_1036,In_584,In_492);
nand U1037 (N_1037,In_594,In_562);
or U1038 (N_1038,In_171,In_603);
and U1039 (N_1039,In_646,In_270);
nand U1040 (N_1040,In_22,In_155);
nor U1041 (N_1041,In_53,In_340);
or U1042 (N_1042,In_239,In_561);
and U1043 (N_1043,In_524,In_734);
or U1044 (N_1044,In_209,In_41);
nor U1045 (N_1045,In_508,In_599);
nand U1046 (N_1046,In_702,In_414);
nor U1047 (N_1047,In_590,In_328);
and U1048 (N_1048,In_631,In_347);
nand U1049 (N_1049,In_511,In_16);
nand U1050 (N_1050,In_431,In_589);
nor U1051 (N_1051,In_187,In_98);
or U1052 (N_1052,In_669,In_152);
or U1053 (N_1053,In_685,In_523);
nor U1054 (N_1054,In_739,In_518);
nor U1055 (N_1055,In_468,In_242);
or U1056 (N_1056,In_123,In_510);
and U1057 (N_1057,In_17,In_195);
nand U1058 (N_1058,In_251,In_482);
or U1059 (N_1059,In_366,In_79);
and U1060 (N_1060,In_507,In_170);
nand U1061 (N_1061,In_608,In_317);
nand U1062 (N_1062,In_365,In_739);
nand U1063 (N_1063,In_392,In_347);
nor U1064 (N_1064,In_178,In_74);
and U1065 (N_1065,In_284,In_536);
nor U1066 (N_1066,In_598,In_66);
and U1067 (N_1067,In_703,In_39);
nand U1068 (N_1068,In_706,In_439);
nor U1069 (N_1069,In_202,In_569);
nor U1070 (N_1070,In_149,In_284);
or U1071 (N_1071,In_326,In_24);
or U1072 (N_1072,In_242,In_529);
nand U1073 (N_1073,In_150,In_555);
xor U1074 (N_1074,In_172,In_600);
nor U1075 (N_1075,In_444,In_187);
and U1076 (N_1076,In_507,In_624);
and U1077 (N_1077,In_563,In_295);
or U1078 (N_1078,In_274,In_685);
or U1079 (N_1079,In_567,In_291);
and U1080 (N_1080,In_29,In_250);
and U1081 (N_1081,In_10,In_2);
nor U1082 (N_1082,In_162,In_571);
or U1083 (N_1083,In_446,In_745);
nand U1084 (N_1084,In_712,In_321);
nor U1085 (N_1085,In_722,In_737);
and U1086 (N_1086,In_579,In_327);
nor U1087 (N_1087,In_104,In_506);
nand U1088 (N_1088,In_711,In_207);
nand U1089 (N_1089,In_8,In_233);
or U1090 (N_1090,In_102,In_292);
nand U1091 (N_1091,In_576,In_126);
nor U1092 (N_1092,In_599,In_336);
nand U1093 (N_1093,In_544,In_319);
or U1094 (N_1094,In_355,In_616);
nor U1095 (N_1095,In_120,In_681);
nor U1096 (N_1096,In_587,In_255);
nor U1097 (N_1097,In_707,In_63);
nor U1098 (N_1098,In_247,In_68);
nor U1099 (N_1099,In_434,In_624);
nor U1100 (N_1100,In_356,In_136);
and U1101 (N_1101,In_465,In_343);
nor U1102 (N_1102,In_182,In_118);
and U1103 (N_1103,In_62,In_595);
nand U1104 (N_1104,In_662,In_355);
nand U1105 (N_1105,In_659,In_678);
nand U1106 (N_1106,In_60,In_660);
and U1107 (N_1107,In_234,In_235);
or U1108 (N_1108,In_591,In_418);
nor U1109 (N_1109,In_71,In_648);
and U1110 (N_1110,In_77,In_572);
or U1111 (N_1111,In_175,In_641);
nand U1112 (N_1112,In_340,In_582);
and U1113 (N_1113,In_56,In_2);
nand U1114 (N_1114,In_534,In_359);
or U1115 (N_1115,In_242,In_71);
and U1116 (N_1116,In_508,In_317);
nand U1117 (N_1117,In_665,In_556);
and U1118 (N_1118,In_690,In_453);
or U1119 (N_1119,In_389,In_640);
nand U1120 (N_1120,In_662,In_184);
or U1121 (N_1121,In_513,In_607);
or U1122 (N_1122,In_213,In_426);
nor U1123 (N_1123,In_279,In_216);
and U1124 (N_1124,In_261,In_273);
nand U1125 (N_1125,In_724,In_139);
nor U1126 (N_1126,In_464,In_591);
or U1127 (N_1127,In_519,In_165);
or U1128 (N_1128,In_356,In_665);
or U1129 (N_1129,In_690,In_426);
nor U1130 (N_1130,In_717,In_216);
or U1131 (N_1131,In_173,In_296);
nand U1132 (N_1132,In_265,In_8);
nand U1133 (N_1133,In_441,In_661);
or U1134 (N_1134,In_106,In_181);
nor U1135 (N_1135,In_538,In_235);
and U1136 (N_1136,In_343,In_363);
nand U1137 (N_1137,In_240,In_364);
nor U1138 (N_1138,In_114,In_473);
and U1139 (N_1139,In_555,In_271);
and U1140 (N_1140,In_19,In_511);
and U1141 (N_1141,In_687,In_518);
and U1142 (N_1142,In_85,In_380);
nand U1143 (N_1143,In_122,In_314);
and U1144 (N_1144,In_77,In_167);
or U1145 (N_1145,In_192,In_246);
and U1146 (N_1146,In_655,In_54);
nor U1147 (N_1147,In_401,In_235);
or U1148 (N_1148,In_175,In_528);
and U1149 (N_1149,In_280,In_342);
nand U1150 (N_1150,In_163,In_268);
nor U1151 (N_1151,In_555,In_195);
and U1152 (N_1152,In_500,In_715);
nor U1153 (N_1153,In_439,In_117);
nand U1154 (N_1154,In_637,In_397);
nand U1155 (N_1155,In_2,In_670);
nor U1156 (N_1156,In_310,In_472);
nand U1157 (N_1157,In_165,In_137);
and U1158 (N_1158,In_277,In_619);
and U1159 (N_1159,In_440,In_19);
or U1160 (N_1160,In_262,In_153);
or U1161 (N_1161,In_290,In_463);
nor U1162 (N_1162,In_655,In_713);
nand U1163 (N_1163,In_276,In_717);
and U1164 (N_1164,In_681,In_210);
and U1165 (N_1165,In_599,In_420);
nand U1166 (N_1166,In_147,In_236);
nand U1167 (N_1167,In_640,In_514);
nand U1168 (N_1168,In_359,In_661);
or U1169 (N_1169,In_697,In_213);
nor U1170 (N_1170,In_545,In_301);
nor U1171 (N_1171,In_628,In_413);
or U1172 (N_1172,In_471,In_214);
or U1173 (N_1173,In_334,In_598);
or U1174 (N_1174,In_291,In_566);
nand U1175 (N_1175,In_606,In_271);
nand U1176 (N_1176,In_162,In_608);
and U1177 (N_1177,In_260,In_457);
nand U1178 (N_1178,In_431,In_621);
or U1179 (N_1179,In_549,In_230);
or U1180 (N_1180,In_598,In_569);
nor U1181 (N_1181,In_121,In_514);
nand U1182 (N_1182,In_465,In_533);
and U1183 (N_1183,In_379,In_1);
nor U1184 (N_1184,In_589,In_262);
and U1185 (N_1185,In_288,In_640);
and U1186 (N_1186,In_80,In_56);
nand U1187 (N_1187,In_374,In_174);
or U1188 (N_1188,In_749,In_406);
or U1189 (N_1189,In_362,In_34);
or U1190 (N_1190,In_153,In_126);
nor U1191 (N_1191,In_180,In_81);
and U1192 (N_1192,In_634,In_21);
or U1193 (N_1193,In_335,In_83);
nand U1194 (N_1194,In_612,In_674);
nor U1195 (N_1195,In_534,In_703);
and U1196 (N_1196,In_222,In_536);
nor U1197 (N_1197,In_491,In_482);
nor U1198 (N_1198,In_328,In_159);
nand U1199 (N_1199,In_685,In_504);
or U1200 (N_1200,In_572,In_564);
nand U1201 (N_1201,In_25,In_203);
or U1202 (N_1202,In_7,In_92);
nand U1203 (N_1203,In_462,In_3);
nand U1204 (N_1204,In_542,In_724);
nor U1205 (N_1205,In_412,In_9);
xnor U1206 (N_1206,In_255,In_107);
nand U1207 (N_1207,In_439,In_737);
nand U1208 (N_1208,In_280,In_436);
and U1209 (N_1209,In_197,In_617);
and U1210 (N_1210,In_666,In_302);
and U1211 (N_1211,In_545,In_313);
nor U1212 (N_1212,In_701,In_68);
and U1213 (N_1213,In_516,In_343);
nand U1214 (N_1214,In_81,In_291);
nand U1215 (N_1215,In_376,In_370);
nor U1216 (N_1216,In_447,In_149);
nand U1217 (N_1217,In_258,In_295);
nand U1218 (N_1218,In_23,In_72);
or U1219 (N_1219,In_87,In_251);
or U1220 (N_1220,In_10,In_660);
nor U1221 (N_1221,In_740,In_43);
nand U1222 (N_1222,In_587,In_596);
nand U1223 (N_1223,In_159,In_386);
nor U1224 (N_1224,In_402,In_636);
nor U1225 (N_1225,In_560,In_671);
nand U1226 (N_1226,In_359,In_180);
nor U1227 (N_1227,In_649,In_175);
nand U1228 (N_1228,In_326,In_258);
and U1229 (N_1229,In_322,In_416);
and U1230 (N_1230,In_713,In_194);
nor U1231 (N_1231,In_390,In_545);
nand U1232 (N_1232,In_467,In_610);
and U1233 (N_1233,In_597,In_718);
nand U1234 (N_1234,In_400,In_558);
nand U1235 (N_1235,In_725,In_32);
nand U1236 (N_1236,In_320,In_472);
and U1237 (N_1237,In_585,In_209);
or U1238 (N_1238,In_56,In_189);
and U1239 (N_1239,In_433,In_91);
and U1240 (N_1240,In_359,In_217);
nor U1241 (N_1241,In_207,In_179);
nand U1242 (N_1242,In_356,In_691);
nor U1243 (N_1243,In_728,In_731);
or U1244 (N_1244,In_107,In_82);
and U1245 (N_1245,In_272,In_134);
nor U1246 (N_1246,In_741,In_280);
or U1247 (N_1247,In_73,In_357);
and U1248 (N_1248,In_431,In_635);
or U1249 (N_1249,In_623,In_65);
and U1250 (N_1250,In_229,In_585);
nand U1251 (N_1251,In_563,In_147);
and U1252 (N_1252,In_321,In_209);
and U1253 (N_1253,In_714,In_454);
nor U1254 (N_1254,In_95,In_452);
nand U1255 (N_1255,In_630,In_530);
nand U1256 (N_1256,In_14,In_40);
nand U1257 (N_1257,In_574,In_170);
nor U1258 (N_1258,In_332,In_668);
and U1259 (N_1259,In_620,In_599);
or U1260 (N_1260,In_373,In_670);
and U1261 (N_1261,In_555,In_35);
xor U1262 (N_1262,In_84,In_418);
nand U1263 (N_1263,In_424,In_554);
or U1264 (N_1264,In_111,In_515);
or U1265 (N_1265,In_453,In_614);
nand U1266 (N_1266,In_743,In_472);
nor U1267 (N_1267,In_735,In_102);
nand U1268 (N_1268,In_411,In_252);
or U1269 (N_1269,In_42,In_683);
or U1270 (N_1270,In_88,In_683);
nor U1271 (N_1271,In_452,In_335);
or U1272 (N_1272,In_408,In_431);
or U1273 (N_1273,In_500,In_553);
and U1274 (N_1274,In_177,In_16);
or U1275 (N_1275,In_197,In_610);
or U1276 (N_1276,In_94,In_581);
and U1277 (N_1277,In_517,In_652);
nor U1278 (N_1278,In_608,In_417);
nor U1279 (N_1279,In_406,In_289);
nand U1280 (N_1280,In_725,In_508);
nand U1281 (N_1281,In_407,In_89);
nand U1282 (N_1282,In_473,In_236);
or U1283 (N_1283,In_471,In_357);
or U1284 (N_1284,In_600,In_495);
nand U1285 (N_1285,In_110,In_263);
nor U1286 (N_1286,In_738,In_115);
nor U1287 (N_1287,In_186,In_315);
or U1288 (N_1288,In_217,In_605);
nand U1289 (N_1289,In_80,In_348);
or U1290 (N_1290,In_293,In_592);
or U1291 (N_1291,In_595,In_299);
nand U1292 (N_1292,In_728,In_272);
nor U1293 (N_1293,In_274,In_417);
nor U1294 (N_1294,In_81,In_395);
nand U1295 (N_1295,In_589,In_712);
or U1296 (N_1296,In_295,In_211);
and U1297 (N_1297,In_429,In_40);
nor U1298 (N_1298,In_398,In_418);
and U1299 (N_1299,In_331,In_639);
and U1300 (N_1300,In_690,In_512);
nand U1301 (N_1301,In_194,In_432);
or U1302 (N_1302,In_38,In_534);
and U1303 (N_1303,In_296,In_691);
nand U1304 (N_1304,In_133,In_177);
and U1305 (N_1305,In_402,In_2);
nor U1306 (N_1306,In_332,In_591);
nor U1307 (N_1307,In_293,In_433);
nor U1308 (N_1308,In_717,In_657);
nand U1309 (N_1309,In_166,In_573);
or U1310 (N_1310,In_551,In_153);
nand U1311 (N_1311,In_133,In_620);
nand U1312 (N_1312,In_37,In_92);
nand U1313 (N_1313,In_432,In_115);
nor U1314 (N_1314,In_564,In_686);
nor U1315 (N_1315,In_460,In_517);
nand U1316 (N_1316,In_428,In_398);
nand U1317 (N_1317,In_272,In_158);
nor U1318 (N_1318,In_429,In_348);
and U1319 (N_1319,In_283,In_515);
nor U1320 (N_1320,In_376,In_221);
nor U1321 (N_1321,In_31,In_297);
nor U1322 (N_1322,In_350,In_99);
nand U1323 (N_1323,In_651,In_0);
and U1324 (N_1324,In_368,In_5);
or U1325 (N_1325,In_669,In_391);
nor U1326 (N_1326,In_530,In_165);
nand U1327 (N_1327,In_732,In_324);
nor U1328 (N_1328,In_232,In_606);
and U1329 (N_1329,In_679,In_306);
nand U1330 (N_1330,In_123,In_367);
nor U1331 (N_1331,In_630,In_21);
or U1332 (N_1332,In_158,In_256);
nand U1333 (N_1333,In_668,In_738);
nor U1334 (N_1334,In_425,In_397);
and U1335 (N_1335,In_204,In_693);
nor U1336 (N_1336,In_186,In_279);
and U1337 (N_1337,In_215,In_24);
nor U1338 (N_1338,In_97,In_37);
and U1339 (N_1339,In_703,In_45);
or U1340 (N_1340,In_242,In_741);
and U1341 (N_1341,In_57,In_124);
and U1342 (N_1342,In_346,In_442);
nand U1343 (N_1343,In_616,In_29);
nand U1344 (N_1344,In_358,In_509);
nor U1345 (N_1345,In_136,In_629);
and U1346 (N_1346,In_577,In_140);
or U1347 (N_1347,In_624,In_265);
and U1348 (N_1348,In_687,In_505);
nor U1349 (N_1349,In_40,In_428);
or U1350 (N_1350,In_296,In_564);
or U1351 (N_1351,In_613,In_508);
nand U1352 (N_1352,In_447,In_15);
or U1353 (N_1353,In_110,In_609);
and U1354 (N_1354,In_499,In_544);
or U1355 (N_1355,In_410,In_573);
nand U1356 (N_1356,In_632,In_350);
and U1357 (N_1357,In_77,In_475);
and U1358 (N_1358,In_405,In_227);
or U1359 (N_1359,In_245,In_435);
nand U1360 (N_1360,In_337,In_434);
nand U1361 (N_1361,In_408,In_553);
nand U1362 (N_1362,In_575,In_510);
nand U1363 (N_1363,In_44,In_109);
and U1364 (N_1364,In_470,In_394);
and U1365 (N_1365,In_99,In_231);
nor U1366 (N_1366,In_545,In_123);
and U1367 (N_1367,In_351,In_228);
or U1368 (N_1368,In_388,In_389);
and U1369 (N_1369,In_415,In_519);
nand U1370 (N_1370,In_330,In_75);
and U1371 (N_1371,In_335,In_460);
nand U1372 (N_1372,In_585,In_314);
nand U1373 (N_1373,In_159,In_322);
nand U1374 (N_1374,In_477,In_717);
and U1375 (N_1375,In_247,In_77);
nor U1376 (N_1376,In_26,In_114);
or U1377 (N_1377,In_336,In_275);
nor U1378 (N_1378,In_309,In_701);
nor U1379 (N_1379,In_103,In_88);
and U1380 (N_1380,In_684,In_614);
or U1381 (N_1381,In_41,In_335);
or U1382 (N_1382,In_714,In_722);
or U1383 (N_1383,In_338,In_440);
or U1384 (N_1384,In_425,In_133);
and U1385 (N_1385,In_400,In_449);
nor U1386 (N_1386,In_727,In_579);
nor U1387 (N_1387,In_718,In_320);
or U1388 (N_1388,In_237,In_312);
nand U1389 (N_1389,In_237,In_533);
nor U1390 (N_1390,In_254,In_222);
nor U1391 (N_1391,In_28,In_231);
and U1392 (N_1392,In_158,In_540);
nor U1393 (N_1393,In_475,In_9);
and U1394 (N_1394,In_493,In_291);
and U1395 (N_1395,In_280,In_546);
or U1396 (N_1396,In_544,In_145);
or U1397 (N_1397,In_745,In_341);
and U1398 (N_1398,In_614,In_736);
nor U1399 (N_1399,In_455,In_4);
or U1400 (N_1400,In_376,In_285);
nor U1401 (N_1401,In_21,In_328);
and U1402 (N_1402,In_349,In_555);
nand U1403 (N_1403,In_74,In_467);
nor U1404 (N_1404,In_703,In_657);
nand U1405 (N_1405,In_537,In_388);
and U1406 (N_1406,In_586,In_120);
nor U1407 (N_1407,In_476,In_579);
nor U1408 (N_1408,In_368,In_553);
nand U1409 (N_1409,In_654,In_668);
and U1410 (N_1410,In_455,In_496);
nand U1411 (N_1411,In_413,In_57);
nor U1412 (N_1412,In_103,In_220);
or U1413 (N_1413,In_299,In_501);
or U1414 (N_1414,In_570,In_624);
nand U1415 (N_1415,In_252,In_84);
or U1416 (N_1416,In_68,In_71);
nor U1417 (N_1417,In_406,In_600);
nand U1418 (N_1418,In_234,In_529);
nor U1419 (N_1419,In_242,In_729);
or U1420 (N_1420,In_251,In_316);
and U1421 (N_1421,In_530,In_323);
or U1422 (N_1422,In_289,In_343);
nand U1423 (N_1423,In_340,In_94);
nand U1424 (N_1424,In_319,In_583);
or U1425 (N_1425,In_0,In_709);
nand U1426 (N_1426,In_511,In_218);
nand U1427 (N_1427,In_411,In_118);
and U1428 (N_1428,In_32,In_316);
or U1429 (N_1429,In_441,In_650);
nor U1430 (N_1430,In_381,In_58);
nor U1431 (N_1431,In_138,In_239);
or U1432 (N_1432,In_631,In_171);
nor U1433 (N_1433,In_238,In_619);
nor U1434 (N_1434,In_47,In_70);
or U1435 (N_1435,In_744,In_519);
nand U1436 (N_1436,In_304,In_738);
nor U1437 (N_1437,In_151,In_689);
or U1438 (N_1438,In_295,In_523);
nor U1439 (N_1439,In_609,In_337);
and U1440 (N_1440,In_292,In_391);
nand U1441 (N_1441,In_215,In_744);
nand U1442 (N_1442,In_45,In_301);
nor U1443 (N_1443,In_16,In_151);
or U1444 (N_1444,In_155,In_733);
and U1445 (N_1445,In_320,In_455);
and U1446 (N_1446,In_420,In_285);
and U1447 (N_1447,In_448,In_485);
nand U1448 (N_1448,In_20,In_532);
and U1449 (N_1449,In_413,In_58);
nand U1450 (N_1450,In_693,In_327);
nand U1451 (N_1451,In_100,In_648);
or U1452 (N_1452,In_312,In_496);
and U1453 (N_1453,In_109,In_23);
nor U1454 (N_1454,In_330,In_727);
nand U1455 (N_1455,In_508,In_418);
nand U1456 (N_1456,In_201,In_525);
and U1457 (N_1457,In_206,In_167);
nor U1458 (N_1458,In_471,In_184);
or U1459 (N_1459,In_564,In_405);
xor U1460 (N_1460,In_294,In_629);
nand U1461 (N_1461,In_632,In_142);
nor U1462 (N_1462,In_386,In_167);
or U1463 (N_1463,In_41,In_463);
nand U1464 (N_1464,In_290,In_617);
or U1465 (N_1465,In_610,In_598);
or U1466 (N_1466,In_290,In_483);
nand U1467 (N_1467,In_538,In_167);
nor U1468 (N_1468,In_216,In_696);
xor U1469 (N_1469,In_339,In_287);
nor U1470 (N_1470,In_9,In_252);
and U1471 (N_1471,In_87,In_517);
and U1472 (N_1472,In_571,In_364);
and U1473 (N_1473,In_614,In_742);
nor U1474 (N_1474,In_275,In_680);
nand U1475 (N_1475,In_712,In_188);
and U1476 (N_1476,In_457,In_21);
nor U1477 (N_1477,In_534,In_446);
and U1478 (N_1478,In_594,In_735);
and U1479 (N_1479,In_75,In_261);
or U1480 (N_1480,In_17,In_526);
nand U1481 (N_1481,In_310,In_367);
or U1482 (N_1482,In_184,In_307);
nor U1483 (N_1483,In_216,In_484);
nor U1484 (N_1484,In_549,In_79);
nand U1485 (N_1485,In_38,In_489);
nor U1486 (N_1486,In_21,In_229);
nand U1487 (N_1487,In_202,In_387);
nand U1488 (N_1488,In_566,In_3);
nor U1489 (N_1489,In_301,In_371);
and U1490 (N_1490,In_527,In_467);
and U1491 (N_1491,In_523,In_526);
or U1492 (N_1492,In_645,In_504);
and U1493 (N_1493,In_566,In_118);
and U1494 (N_1494,In_462,In_246);
and U1495 (N_1495,In_175,In_359);
and U1496 (N_1496,In_197,In_620);
and U1497 (N_1497,In_458,In_297);
and U1498 (N_1498,In_446,In_116);
and U1499 (N_1499,In_475,In_247);
nor U1500 (N_1500,In_415,In_277);
nor U1501 (N_1501,In_164,In_539);
and U1502 (N_1502,In_345,In_621);
nor U1503 (N_1503,In_471,In_318);
and U1504 (N_1504,In_325,In_529);
and U1505 (N_1505,In_369,In_612);
or U1506 (N_1506,In_660,In_530);
xor U1507 (N_1507,In_645,In_18);
and U1508 (N_1508,In_630,In_110);
nand U1509 (N_1509,In_39,In_354);
nor U1510 (N_1510,In_206,In_699);
nor U1511 (N_1511,In_368,In_667);
and U1512 (N_1512,In_294,In_188);
nand U1513 (N_1513,In_406,In_677);
nand U1514 (N_1514,In_659,In_367);
nand U1515 (N_1515,In_549,In_588);
or U1516 (N_1516,In_212,In_99);
and U1517 (N_1517,In_700,In_385);
and U1518 (N_1518,In_226,In_614);
nor U1519 (N_1519,In_20,In_326);
nor U1520 (N_1520,In_735,In_699);
and U1521 (N_1521,In_2,In_389);
or U1522 (N_1522,In_382,In_305);
nand U1523 (N_1523,In_641,In_647);
nor U1524 (N_1524,In_390,In_226);
and U1525 (N_1525,In_181,In_313);
nand U1526 (N_1526,In_45,In_713);
nor U1527 (N_1527,In_111,In_175);
nor U1528 (N_1528,In_105,In_169);
nand U1529 (N_1529,In_57,In_557);
nand U1530 (N_1530,In_563,In_316);
nor U1531 (N_1531,In_438,In_688);
nand U1532 (N_1532,In_654,In_384);
or U1533 (N_1533,In_678,In_703);
and U1534 (N_1534,In_692,In_226);
nand U1535 (N_1535,In_216,In_128);
nor U1536 (N_1536,In_741,In_515);
or U1537 (N_1537,In_436,In_527);
and U1538 (N_1538,In_286,In_625);
nor U1539 (N_1539,In_632,In_623);
and U1540 (N_1540,In_251,In_610);
nor U1541 (N_1541,In_71,In_436);
nand U1542 (N_1542,In_396,In_167);
nor U1543 (N_1543,In_399,In_555);
or U1544 (N_1544,In_158,In_1);
or U1545 (N_1545,In_199,In_381);
or U1546 (N_1546,In_20,In_495);
or U1547 (N_1547,In_68,In_378);
nor U1548 (N_1548,In_475,In_393);
nor U1549 (N_1549,In_671,In_266);
nor U1550 (N_1550,In_56,In_288);
and U1551 (N_1551,In_351,In_324);
and U1552 (N_1552,In_636,In_103);
and U1553 (N_1553,In_660,In_30);
nor U1554 (N_1554,In_152,In_443);
or U1555 (N_1555,In_311,In_225);
nor U1556 (N_1556,In_458,In_399);
or U1557 (N_1557,In_357,In_744);
or U1558 (N_1558,In_596,In_372);
nor U1559 (N_1559,In_194,In_261);
or U1560 (N_1560,In_318,In_18);
or U1561 (N_1561,In_405,In_569);
nor U1562 (N_1562,In_90,In_422);
nor U1563 (N_1563,In_358,In_601);
nand U1564 (N_1564,In_405,In_431);
nand U1565 (N_1565,In_665,In_183);
and U1566 (N_1566,In_369,In_670);
nor U1567 (N_1567,In_515,In_395);
nand U1568 (N_1568,In_538,In_671);
nor U1569 (N_1569,In_550,In_38);
and U1570 (N_1570,In_576,In_444);
and U1571 (N_1571,In_581,In_378);
or U1572 (N_1572,In_535,In_8);
nand U1573 (N_1573,In_187,In_357);
nor U1574 (N_1574,In_47,In_397);
or U1575 (N_1575,In_580,In_48);
nand U1576 (N_1576,In_682,In_176);
nor U1577 (N_1577,In_123,In_520);
nand U1578 (N_1578,In_724,In_516);
and U1579 (N_1579,In_368,In_9);
and U1580 (N_1580,In_254,In_689);
nor U1581 (N_1581,In_502,In_81);
nand U1582 (N_1582,In_441,In_147);
and U1583 (N_1583,In_430,In_703);
or U1584 (N_1584,In_747,In_491);
and U1585 (N_1585,In_242,In_362);
or U1586 (N_1586,In_450,In_411);
nand U1587 (N_1587,In_14,In_551);
xor U1588 (N_1588,In_142,In_214);
nand U1589 (N_1589,In_248,In_517);
or U1590 (N_1590,In_45,In_78);
nand U1591 (N_1591,In_484,In_58);
or U1592 (N_1592,In_477,In_604);
and U1593 (N_1593,In_674,In_409);
nand U1594 (N_1594,In_606,In_317);
or U1595 (N_1595,In_712,In_633);
nand U1596 (N_1596,In_263,In_739);
nand U1597 (N_1597,In_713,In_46);
and U1598 (N_1598,In_63,In_410);
nand U1599 (N_1599,In_696,In_286);
and U1600 (N_1600,In_741,In_653);
and U1601 (N_1601,In_569,In_297);
or U1602 (N_1602,In_361,In_684);
or U1603 (N_1603,In_453,In_431);
and U1604 (N_1604,In_603,In_660);
nand U1605 (N_1605,In_500,In_727);
nor U1606 (N_1606,In_713,In_83);
and U1607 (N_1607,In_391,In_271);
nor U1608 (N_1608,In_197,In_424);
xor U1609 (N_1609,In_137,In_469);
nor U1610 (N_1610,In_244,In_714);
nand U1611 (N_1611,In_310,In_449);
nand U1612 (N_1612,In_264,In_293);
nand U1613 (N_1613,In_42,In_140);
and U1614 (N_1614,In_472,In_541);
nor U1615 (N_1615,In_64,In_738);
nor U1616 (N_1616,In_545,In_675);
nor U1617 (N_1617,In_732,In_133);
and U1618 (N_1618,In_644,In_150);
nand U1619 (N_1619,In_351,In_91);
or U1620 (N_1620,In_546,In_11);
nor U1621 (N_1621,In_679,In_317);
nor U1622 (N_1622,In_384,In_328);
nor U1623 (N_1623,In_560,In_392);
and U1624 (N_1624,In_594,In_423);
nand U1625 (N_1625,In_79,In_156);
nand U1626 (N_1626,In_605,In_268);
or U1627 (N_1627,In_107,In_510);
nand U1628 (N_1628,In_33,In_310);
or U1629 (N_1629,In_640,In_701);
or U1630 (N_1630,In_490,In_467);
or U1631 (N_1631,In_423,In_707);
nor U1632 (N_1632,In_503,In_28);
nor U1633 (N_1633,In_239,In_31);
or U1634 (N_1634,In_496,In_231);
and U1635 (N_1635,In_474,In_559);
and U1636 (N_1636,In_0,In_393);
and U1637 (N_1637,In_530,In_358);
or U1638 (N_1638,In_302,In_474);
and U1639 (N_1639,In_674,In_439);
and U1640 (N_1640,In_562,In_446);
or U1641 (N_1641,In_202,In_550);
nor U1642 (N_1642,In_470,In_128);
nor U1643 (N_1643,In_608,In_173);
or U1644 (N_1644,In_548,In_670);
and U1645 (N_1645,In_22,In_105);
and U1646 (N_1646,In_342,In_362);
nand U1647 (N_1647,In_467,In_17);
or U1648 (N_1648,In_344,In_410);
nand U1649 (N_1649,In_249,In_139);
nand U1650 (N_1650,In_591,In_120);
nor U1651 (N_1651,In_168,In_613);
nor U1652 (N_1652,In_13,In_28);
and U1653 (N_1653,In_372,In_476);
or U1654 (N_1654,In_324,In_75);
nor U1655 (N_1655,In_126,In_445);
nand U1656 (N_1656,In_500,In_118);
nor U1657 (N_1657,In_136,In_95);
and U1658 (N_1658,In_363,In_125);
or U1659 (N_1659,In_18,In_254);
nand U1660 (N_1660,In_697,In_749);
or U1661 (N_1661,In_740,In_618);
and U1662 (N_1662,In_420,In_399);
nand U1663 (N_1663,In_433,In_251);
or U1664 (N_1664,In_39,In_55);
nand U1665 (N_1665,In_425,In_284);
and U1666 (N_1666,In_633,In_285);
nor U1667 (N_1667,In_465,In_85);
and U1668 (N_1668,In_735,In_262);
and U1669 (N_1669,In_97,In_422);
nand U1670 (N_1670,In_693,In_271);
and U1671 (N_1671,In_626,In_692);
and U1672 (N_1672,In_32,In_395);
or U1673 (N_1673,In_652,In_475);
nand U1674 (N_1674,In_182,In_150);
nand U1675 (N_1675,In_662,In_493);
nor U1676 (N_1676,In_463,In_190);
nand U1677 (N_1677,In_98,In_93);
and U1678 (N_1678,In_257,In_530);
and U1679 (N_1679,In_347,In_724);
or U1680 (N_1680,In_573,In_111);
nor U1681 (N_1681,In_737,In_605);
or U1682 (N_1682,In_233,In_705);
nand U1683 (N_1683,In_505,In_344);
and U1684 (N_1684,In_102,In_519);
and U1685 (N_1685,In_107,In_606);
or U1686 (N_1686,In_475,In_65);
nand U1687 (N_1687,In_273,In_464);
nand U1688 (N_1688,In_396,In_622);
nand U1689 (N_1689,In_637,In_83);
nor U1690 (N_1690,In_469,In_537);
or U1691 (N_1691,In_272,In_345);
or U1692 (N_1692,In_204,In_225);
nor U1693 (N_1693,In_742,In_233);
nand U1694 (N_1694,In_332,In_46);
nor U1695 (N_1695,In_314,In_286);
nor U1696 (N_1696,In_281,In_74);
nand U1697 (N_1697,In_59,In_420);
nand U1698 (N_1698,In_223,In_610);
or U1699 (N_1699,In_72,In_417);
and U1700 (N_1700,In_145,In_390);
nand U1701 (N_1701,In_154,In_624);
nand U1702 (N_1702,In_387,In_215);
nor U1703 (N_1703,In_686,In_221);
nand U1704 (N_1704,In_94,In_246);
and U1705 (N_1705,In_102,In_272);
nor U1706 (N_1706,In_301,In_173);
and U1707 (N_1707,In_91,In_476);
nand U1708 (N_1708,In_601,In_197);
and U1709 (N_1709,In_466,In_72);
nor U1710 (N_1710,In_30,In_363);
and U1711 (N_1711,In_554,In_234);
and U1712 (N_1712,In_282,In_602);
xor U1713 (N_1713,In_96,In_629);
nand U1714 (N_1714,In_673,In_363);
or U1715 (N_1715,In_317,In_106);
nand U1716 (N_1716,In_444,In_378);
and U1717 (N_1717,In_539,In_485);
nor U1718 (N_1718,In_372,In_423);
or U1719 (N_1719,In_662,In_348);
and U1720 (N_1720,In_84,In_552);
nand U1721 (N_1721,In_540,In_619);
or U1722 (N_1722,In_243,In_510);
nor U1723 (N_1723,In_550,In_478);
nand U1724 (N_1724,In_280,In_22);
nor U1725 (N_1725,In_185,In_60);
and U1726 (N_1726,In_356,In_227);
and U1727 (N_1727,In_670,In_727);
or U1728 (N_1728,In_555,In_371);
and U1729 (N_1729,In_229,In_463);
nor U1730 (N_1730,In_143,In_484);
nor U1731 (N_1731,In_43,In_731);
and U1732 (N_1732,In_453,In_423);
nor U1733 (N_1733,In_58,In_599);
and U1734 (N_1734,In_515,In_476);
and U1735 (N_1735,In_601,In_344);
nor U1736 (N_1736,In_501,In_366);
or U1737 (N_1737,In_209,In_616);
and U1738 (N_1738,In_368,In_551);
and U1739 (N_1739,In_480,In_432);
nand U1740 (N_1740,In_496,In_508);
nor U1741 (N_1741,In_0,In_191);
nor U1742 (N_1742,In_495,In_392);
nor U1743 (N_1743,In_715,In_204);
nor U1744 (N_1744,In_93,In_686);
nor U1745 (N_1745,In_639,In_399);
and U1746 (N_1746,In_724,In_262);
nor U1747 (N_1747,In_330,In_387);
nand U1748 (N_1748,In_45,In_683);
nor U1749 (N_1749,In_268,In_627);
nand U1750 (N_1750,In_9,In_198);
nor U1751 (N_1751,In_573,In_620);
nor U1752 (N_1752,In_405,In_70);
and U1753 (N_1753,In_370,In_198);
nand U1754 (N_1754,In_488,In_467);
and U1755 (N_1755,In_627,In_95);
nand U1756 (N_1756,In_699,In_663);
and U1757 (N_1757,In_16,In_719);
nand U1758 (N_1758,In_248,In_647);
xnor U1759 (N_1759,In_367,In_84);
nor U1760 (N_1760,In_294,In_397);
nor U1761 (N_1761,In_65,In_495);
nor U1762 (N_1762,In_281,In_562);
nor U1763 (N_1763,In_52,In_288);
nand U1764 (N_1764,In_566,In_70);
or U1765 (N_1765,In_146,In_6);
xnor U1766 (N_1766,In_181,In_435);
or U1767 (N_1767,In_560,In_114);
and U1768 (N_1768,In_456,In_511);
nor U1769 (N_1769,In_712,In_578);
or U1770 (N_1770,In_445,In_552);
or U1771 (N_1771,In_413,In_439);
nor U1772 (N_1772,In_116,In_16);
nand U1773 (N_1773,In_214,In_242);
nor U1774 (N_1774,In_333,In_31);
and U1775 (N_1775,In_156,In_539);
and U1776 (N_1776,In_677,In_30);
and U1777 (N_1777,In_502,In_152);
and U1778 (N_1778,In_324,In_459);
or U1779 (N_1779,In_271,In_258);
and U1780 (N_1780,In_572,In_238);
nor U1781 (N_1781,In_475,In_3);
nor U1782 (N_1782,In_723,In_109);
and U1783 (N_1783,In_136,In_427);
nand U1784 (N_1784,In_391,In_254);
nor U1785 (N_1785,In_718,In_238);
or U1786 (N_1786,In_381,In_12);
nand U1787 (N_1787,In_377,In_42);
nor U1788 (N_1788,In_266,In_512);
or U1789 (N_1789,In_363,In_420);
nor U1790 (N_1790,In_553,In_165);
nor U1791 (N_1791,In_48,In_574);
and U1792 (N_1792,In_367,In_674);
nor U1793 (N_1793,In_273,In_298);
or U1794 (N_1794,In_176,In_363);
nor U1795 (N_1795,In_584,In_20);
nor U1796 (N_1796,In_307,In_616);
nand U1797 (N_1797,In_101,In_658);
or U1798 (N_1798,In_452,In_80);
and U1799 (N_1799,In_379,In_572);
or U1800 (N_1800,In_450,In_422);
nand U1801 (N_1801,In_679,In_575);
and U1802 (N_1802,In_296,In_151);
xor U1803 (N_1803,In_555,In_692);
nor U1804 (N_1804,In_705,In_194);
nor U1805 (N_1805,In_317,In_308);
nor U1806 (N_1806,In_500,In_548);
nor U1807 (N_1807,In_525,In_325);
or U1808 (N_1808,In_278,In_516);
or U1809 (N_1809,In_199,In_723);
nand U1810 (N_1810,In_127,In_418);
nand U1811 (N_1811,In_373,In_61);
nor U1812 (N_1812,In_557,In_186);
nand U1813 (N_1813,In_683,In_474);
and U1814 (N_1814,In_353,In_646);
xor U1815 (N_1815,In_463,In_62);
nor U1816 (N_1816,In_272,In_478);
nor U1817 (N_1817,In_566,In_161);
nor U1818 (N_1818,In_596,In_493);
nand U1819 (N_1819,In_420,In_211);
nand U1820 (N_1820,In_304,In_506);
and U1821 (N_1821,In_339,In_584);
and U1822 (N_1822,In_0,In_223);
nand U1823 (N_1823,In_656,In_393);
nor U1824 (N_1824,In_598,In_57);
nor U1825 (N_1825,In_535,In_12);
or U1826 (N_1826,In_357,In_152);
and U1827 (N_1827,In_152,In_283);
and U1828 (N_1828,In_25,In_18);
nand U1829 (N_1829,In_353,In_734);
and U1830 (N_1830,In_390,In_453);
nor U1831 (N_1831,In_662,In_251);
nor U1832 (N_1832,In_322,In_328);
and U1833 (N_1833,In_606,In_575);
and U1834 (N_1834,In_523,In_155);
nor U1835 (N_1835,In_104,In_225);
nand U1836 (N_1836,In_415,In_76);
nor U1837 (N_1837,In_518,In_492);
nor U1838 (N_1838,In_501,In_239);
and U1839 (N_1839,In_677,In_146);
or U1840 (N_1840,In_344,In_140);
nor U1841 (N_1841,In_377,In_396);
nor U1842 (N_1842,In_678,In_322);
and U1843 (N_1843,In_358,In_281);
nand U1844 (N_1844,In_531,In_340);
and U1845 (N_1845,In_661,In_710);
nor U1846 (N_1846,In_22,In_6);
xnor U1847 (N_1847,In_694,In_390);
nor U1848 (N_1848,In_101,In_479);
and U1849 (N_1849,In_658,In_496);
and U1850 (N_1850,In_628,In_573);
and U1851 (N_1851,In_14,In_494);
and U1852 (N_1852,In_136,In_14);
or U1853 (N_1853,In_476,In_667);
nand U1854 (N_1854,In_739,In_322);
or U1855 (N_1855,In_364,In_138);
and U1856 (N_1856,In_724,In_683);
nand U1857 (N_1857,In_729,In_115);
or U1858 (N_1858,In_382,In_366);
or U1859 (N_1859,In_133,In_1);
and U1860 (N_1860,In_178,In_667);
and U1861 (N_1861,In_667,In_52);
nor U1862 (N_1862,In_78,In_505);
nor U1863 (N_1863,In_262,In_592);
and U1864 (N_1864,In_621,In_604);
and U1865 (N_1865,In_441,In_203);
and U1866 (N_1866,In_175,In_448);
nand U1867 (N_1867,In_219,In_218);
nor U1868 (N_1868,In_504,In_340);
nand U1869 (N_1869,In_33,In_513);
or U1870 (N_1870,In_298,In_647);
nand U1871 (N_1871,In_473,In_338);
nor U1872 (N_1872,In_322,In_19);
and U1873 (N_1873,In_613,In_238);
or U1874 (N_1874,In_177,In_578);
and U1875 (N_1875,In_30,In_733);
nor U1876 (N_1876,In_26,In_205);
or U1877 (N_1877,In_141,In_286);
or U1878 (N_1878,In_179,In_201);
nor U1879 (N_1879,In_232,In_274);
and U1880 (N_1880,In_406,In_364);
nand U1881 (N_1881,In_20,In_519);
nand U1882 (N_1882,In_162,In_249);
nand U1883 (N_1883,In_748,In_491);
and U1884 (N_1884,In_183,In_748);
and U1885 (N_1885,In_75,In_353);
nor U1886 (N_1886,In_695,In_290);
nand U1887 (N_1887,In_222,In_458);
or U1888 (N_1888,In_481,In_692);
nand U1889 (N_1889,In_383,In_713);
nor U1890 (N_1890,In_370,In_325);
or U1891 (N_1891,In_526,In_567);
and U1892 (N_1892,In_437,In_519);
nand U1893 (N_1893,In_126,In_627);
nand U1894 (N_1894,In_534,In_72);
and U1895 (N_1895,In_161,In_555);
nor U1896 (N_1896,In_245,In_2);
nor U1897 (N_1897,In_339,In_546);
and U1898 (N_1898,In_507,In_589);
nand U1899 (N_1899,In_440,In_573);
and U1900 (N_1900,In_74,In_705);
or U1901 (N_1901,In_595,In_469);
nand U1902 (N_1902,In_248,In_713);
or U1903 (N_1903,In_599,In_358);
or U1904 (N_1904,In_42,In_588);
nand U1905 (N_1905,In_659,In_120);
and U1906 (N_1906,In_84,In_581);
and U1907 (N_1907,In_518,In_270);
nor U1908 (N_1908,In_593,In_115);
nor U1909 (N_1909,In_488,In_159);
nand U1910 (N_1910,In_393,In_641);
nor U1911 (N_1911,In_448,In_71);
or U1912 (N_1912,In_636,In_476);
and U1913 (N_1913,In_220,In_41);
and U1914 (N_1914,In_20,In_340);
or U1915 (N_1915,In_684,In_87);
nor U1916 (N_1916,In_386,In_130);
and U1917 (N_1917,In_241,In_186);
or U1918 (N_1918,In_562,In_47);
nor U1919 (N_1919,In_642,In_708);
and U1920 (N_1920,In_67,In_429);
and U1921 (N_1921,In_372,In_7);
nand U1922 (N_1922,In_735,In_240);
nor U1923 (N_1923,In_596,In_373);
nand U1924 (N_1924,In_142,In_511);
or U1925 (N_1925,In_240,In_230);
nor U1926 (N_1926,In_648,In_99);
or U1927 (N_1927,In_596,In_690);
and U1928 (N_1928,In_190,In_83);
or U1929 (N_1929,In_45,In_533);
nor U1930 (N_1930,In_454,In_331);
and U1931 (N_1931,In_44,In_570);
nor U1932 (N_1932,In_289,In_535);
nand U1933 (N_1933,In_95,In_360);
nand U1934 (N_1934,In_696,In_356);
nand U1935 (N_1935,In_712,In_678);
or U1936 (N_1936,In_284,In_241);
nor U1937 (N_1937,In_17,In_603);
nand U1938 (N_1938,In_65,In_536);
or U1939 (N_1939,In_572,In_234);
or U1940 (N_1940,In_712,In_422);
nor U1941 (N_1941,In_709,In_742);
and U1942 (N_1942,In_304,In_703);
xnor U1943 (N_1943,In_103,In_320);
nor U1944 (N_1944,In_53,In_590);
or U1945 (N_1945,In_439,In_538);
or U1946 (N_1946,In_572,In_260);
nor U1947 (N_1947,In_308,In_615);
nor U1948 (N_1948,In_290,In_557);
nor U1949 (N_1949,In_472,In_239);
and U1950 (N_1950,In_127,In_298);
and U1951 (N_1951,In_665,In_217);
and U1952 (N_1952,In_217,In_472);
nor U1953 (N_1953,In_115,In_552);
nand U1954 (N_1954,In_137,In_639);
or U1955 (N_1955,In_697,In_131);
nor U1956 (N_1956,In_25,In_285);
or U1957 (N_1957,In_117,In_446);
and U1958 (N_1958,In_528,In_364);
nor U1959 (N_1959,In_257,In_393);
or U1960 (N_1960,In_650,In_515);
xor U1961 (N_1961,In_86,In_609);
and U1962 (N_1962,In_58,In_61);
nor U1963 (N_1963,In_391,In_86);
nor U1964 (N_1964,In_67,In_747);
or U1965 (N_1965,In_703,In_714);
and U1966 (N_1966,In_246,In_599);
nand U1967 (N_1967,In_46,In_88);
nor U1968 (N_1968,In_332,In_102);
and U1969 (N_1969,In_459,In_205);
nand U1970 (N_1970,In_227,In_514);
nor U1971 (N_1971,In_93,In_208);
nor U1972 (N_1972,In_135,In_12);
nand U1973 (N_1973,In_556,In_123);
and U1974 (N_1974,In_379,In_560);
nor U1975 (N_1975,In_680,In_521);
nor U1976 (N_1976,In_204,In_379);
and U1977 (N_1977,In_372,In_74);
or U1978 (N_1978,In_213,In_162);
or U1979 (N_1979,In_348,In_574);
xnor U1980 (N_1980,In_288,In_86);
or U1981 (N_1981,In_460,In_12);
nand U1982 (N_1982,In_118,In_601);
nor U1983 (N_1983,In_697,In_48);
nand U1984 (N_1984,In_607,In_22);
and U1985 (N_1985,In_357,In_604);
nor U1986 (N_1986,In_693,In_471);
nand U1987 (N_1987,In_143,In_542);
or U1988 (N_1988,In_143,In_130);
nor U1989 (N_1989,In_400,In_405);
nand U1990 (N_1990,In_656,In_526);
or U1991 (N_1991,In_612,In_743);
and U1992 (N_1992,In_446,In_693);
nor U1993 (N_1993,In_342,In_143);
or U1994 (N_1994,In_197,In_310);
nand U1995 (N_1995,In_185,In_526);
and U1996 (N_1996,In_546,In_248);
nor U1997 (N_1997,In_361,In_740);
nor U1998 (N_1998,In_479,In_578);
or U1999 (N_1999,In_25,In_499);
nor U2000 (N_2000,In_393,In_100);
nor U2001 (N_2001,In_483,In_179);
xor U2002 (N_2002,In_23,In_70);
or U2003 (N_2003,In_340,In_170);
or U2004 (N_2004,In_519,In_550);
nor U2005 (N_2005,In_582,In_290);
nor U2006 (N_2006,In_536,In_442);
nor U2007 (N_2007,In_318,In_311);
and U2008 (N_2008,In_497,In_269);
nand U2009 (N_2009,In_4,In_421);
and U2010 (N_2010,In_746,In_743);
nor U2011 (N_2011,In_52,In_378);
and U2012 (N_2012,In_478,In_263);
or U2013 (N_2013,In_164,In_449);
nor U2014 (N_2014,In_498,In_333);
nor U2015 (N_2015,In_448,In_604);
nor U2016 (N_2016,In_371,In_354);
or U2017 (N_2017,In_640,In_292);
and U2018 (N_2018,In_18,In_587);
nand U2019 (N_2019,In_377,In_72);
and U2020 (N_2020,In_614,In_556);
or U2021 (N_2021,In_315,In_623);
nor U2022 (N_2022,In_413,In_292);
and U2023 (N_2023,In_517,In_681);
nand U2024 (N_2024,In_239,In_626);
and U2025 (N_2025,In_532,In_708);
or U2026 (N_2026,In_154,In_131);
nand U2027 (N_2027,In_277,In_696);
and U2028 (N_2028,In_647,In_611);
and U2029 (N_2029,In_567,In_420);
nand U2030 (N_2030,In_746,In_227);
or U2031 (N_2031,In_61,In_495);
and U2032 (N_2032,In_603,In_115);
and U2033 (N_2033,In_317,In_636);
and U2034 (N_2034,In_171,In_595);
nor U2035 (N_2035,In_310,In_23);
and U2036 (N_2036,In_586,In_12);
nand U2037 (N_2037,In_157,In_302);
or U2038 (N_2038,In_522,In_348);
or U2039 (N_2039,In_258,In_316);
nor U2040 (N_2040,In_57,In_363);
or U2041 (N_2041,In_296,In_374);
and U2042 (N_2042,In_470,In_431);
and U2043 (N_2043,In_306,In_148);
and U2044 (N_2044,In_233,In_184);
nor U2045 (N_2045,In_420,In_578);
nand U2046 (N_2046,In_445,In_118);
nor U2047 (N_2047,In_562,In_626);
nor U2048 (N_2048,In_167,In_39);
and U2049 (N_2049,In_350,In_582);
nor U2050 (N_2050,In_257,In_616);
and U2051 (N_2051,In_321,In_69);
and U2052 (N_2052,In_390,In_111);
or U2053 (N_2053,In_708,In_5);
or U2054 (N_2054,In_241,In_731);
nor U2055 (N_2055,In_634,In_168);
nor U2056 (N_2056,In_356,In_75);
nor U2057 (N_2057,In_518,In_529);
nor U2058 (N_2058,In_471,In_712);
and U2059 (N_2059,In_108,In_584);
or U2060 (N_2060,In_571,In_736);
or U2061 (N_2061,In_611,In_93);
or U2062 (N_2062,In_540,In_79);
or U2063 (N_2063,In_141,In_355);
or U2064 (N_2064,In_582,In_736);
and U2065 (N_2065,In_260,In_340);
or U2066 (N_2066,In_548,In_398);
xor U2067 (N_2067,In_294,In_345);
nor U2068 (N_2068,In_48,In_328);
nand U2069 (N_2069,In_417,In_17);
nand U2070 (N_2070,In_208,In_128);
nand U2071 (N_2071,In_477,In_315);
nor U2072 (N_2072,In_708,In_292);
nand U2073 (N_2073,In_41,In_153);
and U2074 (N_2074,In_611,In_144);
or U2075 (N_2075,In_474,In_299);
or U2076 (N_2076,In_559,In_69);
and U2077 (N_2077,In_676,In_22);
nor U2078 (N_2078,In_25,In_413);
or U2079 (N_2079,In_589,In_382);
and U2080 (N_2080,In_201,In_299);
nor U2081 (N_2081,In_304,In_500);
nor U2082 (N_2082,In_116,In_415);
or U2083 (N_2083,In_509,In_453);
nor U2084 (N_2084,In_34,In_246);
and U2085 (N_2085,In_662,In_185);
nor U2086 (N_2086,In_363,In_56);
nor U2087 (N_2087,In_263,In_524);
or U2088 (N_2088,In_242,In_22);
or U2089 (N_2089,In_599,In_610);
or U2090 (N_2090,In_462,In_172);
nand U2091 (N_2091,In_69,In_440);
or U2092 (N_2092,In_43,In_684);
or U2093 (N_2093,In_572,In_179);
and U2094 (N_2094,In_266,In_511);
or U2095 (N_2095,In_669,In_633);
or U2096 (N_2096,In_148,In_127);
nand U2097 (N_2097,In_227,In_725);
or U2098 (N_2098,In_160,In_275);
and U2099 (N_2099,In_128,In_608);
nand U2100 (N_2100,In_536,In_41);
nand U2101 (N_2101,In_408,In_351);
nand U2102 (N_2102,In_60,In_607);
nor U2103 (N_2103,In_246,In_370);
or U2104 (N_2104,In_637,In_654);
nand U2105 (N_2105,In_468,In_737);
nand U2106 (N_2106,In_499,In_672);
and U2107 (N_2107,In_392,In_115);
and U2108 (N_2108,In_439,In_470);
or U2109 (N_2109,In_556,In_133);
nand U2110 (N_2110,In_708,In_43);
and U2111 (N_2111,In_535,In_502);
nand U2112 (N_2112,In_439,In_576);
and U2113 (N_2113,In_254,In_4);
nand U2114 (N_2114,In_262,In_491);
and U2115 (N_2115,In_448,In_718);
nand U2116 (N_2116,In_403,In_14);
and U2117 (N_2117,In_370,In_611);
and U2118 (N_2118,In_169,In_719);
nand U2119 (N_2119,In_258,In_241);
nor U2120 (N_2120,In_193,In_95);
nand U2121 (N_2121,In_453,In_224);
nand U2122 (N_2122,In_307,In_380);
nand U2123 (N_2123,In_260,In_309);
or U2124 (N_2124,In_252,In_386);
or U2125 (N_2125,In_309,In_325);
nand U2126 (N_2126,In_155,In_272);
and U2127 (N_2127,In_690,In_678);
or U2128 (N_2128,In_697,In_215);
or U2129 (N_2129,In_482,In_686);
or U2130 (N_2130,In_205,In_73);
nor U2131 (N_2131,In_479,In_360);
nand U2132 (N_2132,In_598,In_114);
and U2133 (N_2133,In_188,In_28);
and U2134 (N_2134,In_298,In_570);
nand U2135 (N_2135,In_408,In_89);
and U2136 (N_2136,In_257,In_621);
and U2137 (N_2137,In_545,In_256);
or U2138 (N_2138,In_154,In_619);
and U2139 (N_2139,In_439,In_558);
nand U2140 (N_2140,In_683,In_595);
nor U2141 (N_2141,In_338,In_496);
nor U2142 (N_2142,In_127,In_449);
xnor U2143 (N_2143,In_720,In_479);
and U2144 (N_2144,In_702,In_75);
nor U2145 (N_2145,In_681,In_219);
nand U2146 (N_2146,In_155,In_468);
nand U2147 (N_2147,In_424,In_87);
nand U2148 (N_2148,In_552,In_359);
nand U2149 (N_2149,In_583,In_329);
nor U2150 (N_2150,In_430,In_385);
and U2151 (N_2151,In_559,In_88);
or U2152 (N_2152,In_54,In_707);
nand U2153 (N_2153,In_667,In_104);
nand U2154 (N_2154,In_473,In_29);
or U2155 (N_2155,In_499,In_106);
or U2156 (N_2156,In_14,In_60);
or U2157 (N_2157,In_568,In_176);
or U2158 (N_2158,In_108,In_69);
or U2159 (N_2159,In_661,In_626);
or U2160 (N_2160,In_618,In_71);
and U2161 (N_2161,In_92,In_563);
and U2162 (N_2162,In_182,In_719);
nand U2163 (N_2163,In_69,In_141);
nand U2164 (N_2164,In_332,In_250);
and U2165 (N_2165,In_397,In_344);
and U2166 (N_2166,In_674,In_585);
nand U2167 (N_2167,In_340,In_720);
and U2168 (N_2168,In_573,In_363);
or U2169 (N_2169,In_54,In_736);
nand U2170 (N_2170,In_519,In_217);
or U2171 (N_2171,In_665,In_210);
nand U2172 (N_2172,In_215,In_275);
nand U2173 (N_2173,In_704,In_179);
nor U2174 (N_2174,In_422,In_8);
nor U2175 (N_2175,In_555,In_107);
and U2176 (N_2176,In_401,In_446);
nand U2177 (N_2177,In_531,In_498);
and U2178 (N_2178,In_576,In_363);
or U2179 (N_2179,In_604,In_394);
or U2180 (N_2180,In_389,In_495);
nor U2181 (N_2181,In_621,In_484);
and U2182 (N_2182,In_165,In_117);
or U2183 (N_2183,In_345,In_111);
or U2184 (N_2184,In_385,In_613);
or U2185 (N_2185,In_715,In_321);
or U2186 (N_2186,In_37,In_25);
nand U2187 (N_2187,In_320,In_143);
or U2188 (N_2188,In_721,In_534);
nand U2189 (N_2189,In_369,In_451);
and U2190 (N_2190,In_64,In_720);
or U2191 (N_2191,In_654,In_78);
nor U2192 (N_2192,In_746,In_526);
and U2193 (N_2193,In_456,In_156);
nor U2194 (N_2194,In_587,In_74);
or U2195 (N_2195,In_375,In_702);
nor U2196 (N_2196,In_42,In_403);
nor U2197 (N_2197,In_647,In_545);
or U2198 (N_2198,In_696,In_655);
nand U2199 (N_2199,In_241,In_462);
nor U2200 (N_2200,In_430,In_96);
and U2201 (N_2201,In_578,In_593);
nor U2202 (N_2202,In_438,In_616);
nor U2203 (N_2203,In_377,In_405);
or U2204 (N_2204,In_325,In_592);
nand U2205 (N_2205,In_507,In_57);
or U2206 (N_2206,In_353,In_167);
nor U2207 (N_2207,In_52,In_304);
or U2208 (N_2208,In_356,In_617);
and U2209 (N_2209,In_327,In_458);
or U2210 (N_2210,In_721,In_394);
or U2211 (N_2211,In_70,In_147);
or U2212 (N_2212,In_139,In_178);
or U2213 (N_2213,In_395,In_208);
and U2214 (N_2214,In_673,In_56);
nand U2215 (N_2215,In_528,In_486);
nand U2216 (N_2216,In_142,In_497);
nor U2217 (N_2217,In_504,In_571);
or U2218 (N_2218,In_433,In_124);
nor U2219 (N_2219,In_257,In_718);
nor U2220 (N_2220,In_471,In_203);
and U2221 (N_2221,In_718,In_539);
and U2222 (N_2222,In_680,In_293);
nor U2223 (N_2223,In_452,In_131);
or U2224 (N_2224,In_320,In_347);
nand U2225 (N_2225,In_133,In_38);
nand U2226 (N_2226,In_280,In_262);
or U2227 (N_2227,In_277,In_547);
nor U2228 (N_2228,In_208,In_245);
or U2229 (N_2229,In_660,In_470);
nor U2230 (N_2230,In_199,In_365);
or U2231 (N_2231,In_563,In_572);
and U2232 (N_2232,In_173,In_73);
and U2233 (N_2233,In_487,In_299);
and U2234 (N_2234,In_114,In_152);
or U2235 (N_2235,In_254,In_490);
nand U2236 (N_2236,In_195,In_503);
nor U2237 (N_2237,In_338,In_54);
nand U2238 (N_2238,In_691,In_557);
or U2239 (N_2239,In_98,In_703);
nand U2240 (N_2240,In_334,In_152);
and U2241 (N_2241,In_570,In_589);
nor U2242 (N_2242,In_407,In_576);
nand U2243 (N_2243,In_705,In_172);
nor U2244 (N_2244,In_81,In_120);
and U2245 (N_2245,In_58,In_503);
nand U2246 (N_2246,In_122,In_400);
and U2247 (N_2247,In_413,In_719);
nor U2248 (N_2248,In_63,In_317);
nor U2249 (N_2249,In_27,In_252);
and U2250 (N_2250,In_40,In_71);
nand U2251 (N_2251,In_205,In_93);
nand U2252 (N_2252,In_212,In_723);
nand U2253 (N_2253,In_584,In_335);
nor U2254 (N_2254,In_650,In_615);
nor U2255 (N_2255,In_325,In_359);
and U2256 (N_2256,In_444,In_122);
or U2257 (N_2257,In_310,In_228);
nor U2258 (N_2258,In_0,In_604);
or U2259 (N_2259,In_483,In_639);
nor U2260 (N_2260,In_193,In_453);
and U2261 (N_2261,In_453,In_330);
xnor U2262 (N_2262,In_474,In_548);
or U2263 (N_2263,In_8,In_524);
nor U2264 (N_2264,In_539,In_104);
nand U2265 (N_2265,In_531,In_141);
nand U2266 (N_2266,In_659,In_531);
or U2267 (N_2267,In_49,In_96);
nand U2268 (N_2268,In_741,In_209);
nand U2269 (N_2269,In_226,In_145);
and U2270 (N_2270,In_37,In_592);
and U2271 (N_2271,In_49,In_105);
or U2272 (N_2272,In_280,In_662);
nor U2273 (N_2273,In_202,In_336);
and U2274 (N_2274,In_349,In_214);
and U2275 (N_2275,In_168,In_497);
and U2276 (N_2276,In_679,In_12);
and U2277 (N_2277,In_251,In_123);
or U2278 (N_2278,In_211,In_69);
and U2279 (N_2279,In_108,In_153);
xor U2280 (N_2280,In_24,In_232);
and U2281 (N_2281,In_437,In_559);
or U2282 (N_2282,In_295,In_610);
and U2283 (N_2283,In_412,In_565);
and U2284 (N_2284,In_64,In_477);
nand U2285 (N_2285,In_62,In_207);
or U2286 (N_2286,In_535,In_496);
and U2287 (N_2287,In_342,In_272);
and U2288 (N_2288,In_322,In_605);
nor U2289 (N_2289,In_553,In_495);
or U2290 (N_2290,In_188,In_445);
nand U2291 (N_2291,In_79,In_633);
nor U2292 (N_2292,In_189,In_225);
or U2293 (N_2293,In_203,In_721);
and U2294 (N_2294,In_383,In_495);
nor U2295 (N_2295,In_568,In_144);
and U2296 (N_2296,In_718,In_592);
and U2297 (N_2297,In_447,In_438);
or U2298 (N_2298,In_105,In_740);
and U2299 (N_2299,In_656,In_568);
nand U2300 (N_2300,In_151,In_289);
nor U2301 (N_2301,In_697,In_111);
or U2302 (N_2302,In_313,In_381);
nand U2303 (N_2303,In_496,In_97);
and U2304 (N_2304,In_242,In_736);
or U2305 (N_2305,In_674,In_263);
nand U2306 (N_2306,In_352,In_536);
nor U2307 (N_2307,In_507,In_198);
nand U2308 (N_2308,In_369,In_278);
nand U2309 (N_2309,In_374,In_367);
nand U2310 (N_2310,In_687,In_615);
nor U2311 (N_2311,In_697,In_138);
or U2312 (N_2312,In_191,In_206);
nor U2313 (N_2313,In_572,In_421);
nor U2314 (N_2314,In_0,In_704);
nor U2315 (N_2315,In_470,In_668);
and U2316 (N_2316,In_267,In_160);
nand U2317 (N_2317,In_270,In_7);
nor U2318 (N_2318,In_632,In_263);
nand U2319 (N_2319,In_499,In_113);
and U2320 (N_2320,In_452,In_633);
or U2321 (N_2321,In_556,In_533);
and U2322 (N_2322,In_399,In_737);
nand U2323 (N_2323,In_14,In_2);
or U2324 (N_2324,In_29,In_551);
nor U2325 (N_2325,In_432,In_496);
and U2326 (N_2326,In_579,In_459);
nand U2327 (N_2327,In_685,In_744);
or U2328 (N_2328,In_306,In_70);
nor U2329 (N_2329,In_513,In_619);
nand U2330 (N_2330,In_414,In_715);
nor U2331 (N_2331,In_246,In_616);
or U2332 (N_2332,In_677,In_495);
and U2333 (N_2333,In_43,In_105);
and U2334 (N_2334,In_665,In_654);
nor U2335 (N_2335,In_471,In_525);
nor U2336 (N_2336,In_56,In_601);
nor U2337 (N_2337,In_365,In_157);
and U2338 (N_2338,In_551,In_276);
or U2339 (N_2339,In_499,In_218);
or U2340 (N_2340,In_16,In_69);
and U2341 (N_2341,In_42,In_476);
or U2342 (N_2342,In_470,In_504);
nor U2343 (N_2343,In_202,In_666);
and U2344 (N_2344,In_138,In_156);
or U2345 (N_2345,In_432,In_124);
and U2346 (N_2346,In_622,In_114);
nand U2347 (N_2347,In_316,In_508);
nand U2348 (N_2348,In_731,In_59);
nand U2349 (N_2349,In_201,In_184);
xor U2350 (N_2350,In_7,In_116);
nand U2351 (N_2351,In_139,In_396);
or U2352 (N_2352,In_220,In_551);
and U2353 (N_2353,In_433,In_647);
or U2354 (N_2354,In_612,In_552);
nor U2355 (N_2355,In_178,In_636);
nand U2356 (N_2356,In_227,In_146);
nand U2357 (N_2357,In_346,In_526);
nand U2358 (N_2358,In_568,In_111);
nor U2359 (N_2359,In_687,In_95);
nor U2360 (N_2360,In_418,In_17);
or U2361 (N_2361,In_131,In_6);
nand U2362 (N_2362,In_572,In_82);
or U2363 (N_2363,In_110,In_495);
xor U2364 (N_2364,In_656,In_238);
nand U2365 (N_2365,In_283,In_271);
and U2366 (N_2366,In_217,In_93);
nand U2367 (N_2367,In_710,In_619);
nand U2368 (N_2368,In_200,In_42);
nor U2369 (N_2369,In_719,In_221);
or U2370 (N_2370,In_595,In_611);
and U2371 (N_2371,In_11,In_177);
and U2372 (N_2372,In_361,In_533);
nand U2373 (N_2373,In_662,In_721);
nand U2374 (N_2374,In_237,In_511);
or U2375 (N_2375,In_364,In_367);
nand U2376 (N_2376,In_305,In_228);
nand U2377 (N_2377,In_18,In_725);
and U2378 (N_2378,In_159,In_616);
nor U2379 (N_2379,In_351,In_289);
nand U2380 (N_2380,In_563,In_601);
nand U2381 (N_2381,In_88,In_146);
or U2382 (N_2382,In_166,In_624);
nor U2383 (N_2383,In_350,In_307);
nor U2384 (N_2384,In_110,In_552);
nand U2385 (N_2385,In_578,In_426);
or U2386 (N_2386,In_359,In_129);
or U2387 (N_2387,In_146,In_56);
or U2388 (N_2388,In_551,In_413);
nor U2389 (N_2389,In_675,In_287);
nand U2390 (N_2390,In_649,In_162);
or U2391 (N_2391,In_452,In_551);
nor U2392 (N_2392,In_198,In_642);
and U2393 (N_2393,In_272,In_671);
and U2394 (N_2394,In_198,In_303);
nand U2395 (N_2395,In_515,In_549);
nand U2396 (N_2396,In_746,In_667);
nand U2397 (N_2397,In_301,In_33);
or U2398 (N_2398,In_104,In_120);
or U2399 (N_2399,In_542,In_457);
nor U2400 (N_2400,In_334,In_632);
nor U2401 (N_2401,In_20,In_618);
nand U2402 (N_2402,In_644,In_275);
or U2403 (N_2403,In_740,In_8);
nand U2404 (N_2404,In_718,In_296);
and U2405 (N_2405,In_427,In_224);
or U2406 (N_2406,In_675,In_406);
or U2407 (N_2407,In_35,In_61);
and U2408 (N_2408,In_494,In_550);
or U2409 (N_2409,In_437,In_18);
and U2410 (N_2410,In_432,In_542);
xnor U2411 (N_2411,In_114,In_292);
or U2412 (N_2412,In_262,In_605);
and U2413 (N_2413,In_197,In_707);
or U2414 (N_2414,In_659,In_67);
and U2415 (N_2415,In_559,In_746);
nand U2416 (N_2416,In_208,In_160);
and U2417 (N_2417,In_676,In_694);
nor U2418 (N_2418,In_259,In_449);
nor U2419 (N_2419,In_461,In_291);
and U2420 (N_2420,In_254,In_470);
nor U2421 (N_2421,In_361,In_479);
or U2422 (N_2422,In_520,In_372);
nand U2423 (N_2423,In_24,In_228);
or U2424 (N_2424,In_183,In_430);
or U2425 (N_2425,In_543,In_144);
or U2426 (N_2426,In_504,In_326);
and U2427 (N_2427,In_420,In_415);
and U2428 (N_2428,In_559,In_693);
or U2429 (N_2429,In_383,In_216);
or U2430 (N_2430,In_306,In_144);
nor U2431 (N_2431,In_309,In_747);
nor U2432 (N_2432,In_203,In_737);
nand U2433 (N_2433,In_90,In_415);
and U2434 (N_2434,In_21,In_459);
or U2435 (N_2435,In_589,In_397);
and U2436 (N_2436,In_123,In_379);
or U2437 (N_2437,In_281,In_100);
nor U2438 (N_2438,In_150,In_541);
nand U2439 (N_2439,In_493,In_114);
and U2440 (N_2440,In_253,In_729);
nor U2441 (N_2441,In_258,In_69);
and U2442 (N_2442,In_509,In_24);
and U2443 (N_2443,In_285,In_360);
and U2444 (N_2444,In_287,In_555);
nand U2445 (N_2445,In_156,In_657);
or U2446 (N_2446,In_464,In_644);
and U2447 (N_2447,In_639,In_364);
and U2448 (N_2448,In_43,In_653);
or U2449 (N_2449,In_46,In_81);
nand U2450 (N_2450,In_297,In_556);
nor U2451 (N_2451,In_475,In_647);
nor U2452 (N_2452,In_306,In_170);
nand U2453 (N_2453,In_385,In_185);
and U2454 (N_2454,In_73,In_159);
and U2455 (N_2455,In_612,In_509);
or U2456 (N_2456,In_102,In_293);
and U2457 (N_2457,In_90,In_365);
and U2458 (N_2458,In_555,In_472);
nor U2459 (N_2459,In_106,In_693);
nand U2460 (N_2460,In_253,In_520);
or U2461 (N_2461,In_112,In_685);
nand U2462 (N_2462,In_155,In_1);
nand U2463 (N_2463,In_514,In_111);
nand U2464 (N_2464,In_671,In_653);
and U2465 (N_2465,In_424,In_120);
nor U2466 (N_2466,In_328,In_475);
nand U2467 (N_2467,In_616,In_524);
nor U2468 (N_2468,In_486,In_589);
or U2469 (N_2469,In_430,In_733);
or U2470 (N_2470,In_233,In_669);
and U2471 (N_2471,In_176,In_267);
nand U2472 (N_2472,In_150,In_519);
and U2473 (N_2473,In_588,In_396);
and U2474 (N_2474,In_479,In_501);
or U2475 (N_2475,In_8,In_110);
and U2476 (N_2476,In_295,In_429);
nand U2477 (N_2477,In_342,In_482);
nand U2478 (N_2478,In_77,In_185);
or U2479 (N_2479,In_517,In_277);
or U2480 (N_2480,In_433,In_129);
nand U2481 (N_2481,In_188,In_310);
nor U2482 (N_2482,In_15,In_413);
xnor U2483 (N_2483,In_82,In_550);
nand U2484 (N_2484,In_352,In_194);
nor U2485 (N_2485,In_358,In_186);
nand U2486 (N_2486,In_406,In_713);
xor U2487 (N_2487,In_288,In_654);
nor U2488 (N_2488,In_237,In_662);
nand U2489 (N_2489,In_165,In_565);
nand U2490 (N_2490,In_505,In_139);
nand U2491 (N_2491,In_225,In_634);
or U2492 (N_2492,In_341,In_391);
nand U2493 (N_2493,In_495,In_241);
nor U2494 (N_2494,In_636,In_181);
nand U2495 (N_2495,In_93,In_693);
and U2496 (N_2496,In_91,In_486);
nor U2497 (N_2497,In_427,In_616);
nand U2498 (N_2498,In_416,In_34);
nand U2499 (N_2499,In_83,In_103);
and U2500 (N_2500,N_604,N_102);
or U2501 (N_2501,N_2488,N_1976);
and U2502 (N_2502,N_1405,N_766);
nor U2503 (N_2503,N_1646,N_28);
and U2504 (N_2504,N_1468,N_630);
nand U2505 (N_2505,N_137,N_30);
and U2506 (N_2506,N_1389,N_1851);
nor U2507 (N_2507,N_552,N_1877);
nand U2508 (N_2508,N_524,N_311);
or U2509 (N_2509,N_962,N_2398);
and U2510 (N_2510,N_1072,N_1221);
and U2511 (N_2511,N_1192,N_2242);
or U2512 (N_2512,N_338,N_675);
and U2513 (N_2513,N_1638,N_833);
and U2514 (N_2514,N_1053,N_1573);
and U2515 (N_2515,N_2463,N_345);
nor U2516 (N_2516,N_2026,N_896);
xor U2517 (N_2517,N_2091,N_360);
nand U2518 (N_2518,N_803,N_2399);
and U2519 (N_2519,N_2316,N_2163);
or U2520 (N_2520,N_1358,N_373);
nor U2521 (N_2521,N_5,N_1472);
and U2522 (N_2522,N_1193,N_1567);
and U2523 (N_2523,N_1157,N_1351);
nand U2524 (N_2524,N_2165,N_1561);
nor U2525 (N_2525,N_1957,N_2396);
xor U2526 (N_2526,N_888,N_405);
nand U2527 (N_2527,N_2111,N_1269);
or U2528 (N_2528,N_1796,N_1060);
or U2529 (N_2529,N_2154,N_2365);
nor U2530 (N_2530,N_1434,N_152);
nand U2531 (N_2531,N_774,N_1922);
nor U2532 (N_2532,N_12,N_238);
nand U2533 (N_2533,N_2344,N_2039);
nand U2534 (N_2534,N_1534,N_1954);
or U2535 (N_2535,N_2182,N_1264);
or U2536 (N_2536,N_1081,N_1489);
nor U2537 (N_2537,N_1572,N_1029);
and U2538 (N_2538,N_1150,N_299);
nor U2539 (N_2539,N_1168,N_1887);
nor U2540 (N_2540,N_1841,N_849);
nand U2541 (N_2541,N_1947,N_2253);
or U2542 (N_2542,N_698,N_1823);
nand U2543 (N_2543,N_595,N_9);
and U2544 (N_2544,N_166,N_747);
nand U2545 (N_2545,N_1844,N_575);
nand U2546 (N_2546,N_1052,N_915);
and U2547 (N_2547,N_1888,N_2128);
nor U2548 (N_2548,N_1104,N_106);
and U2549 (N_2549,N_1963,N_2226);
nand U2550 (N_2550,N_1842,N_2441);
and U2551 (N_2551,N_51,N_1165);
nor U2552 (N_2552,N_2232,N_1680);
nor U2553 (N_2553,N_1798,N_2015);
and U2554 (N_2554,N_2099,N_977);
and U2555 (N_2555,N_2268,N_45);
nand U2556 (N_2556,N_673,N_1375);
or U2557 (N_2557,N_2070,N_113);
nor U2558 (N_2558,N_1691,N_605);
nand U2559 (N_2559,N_2043,N_1525);
and U2560 (N_2560,N_826,N_1202);
nor U2561 (N_2561,N_1324,N_703);
nor U2562 (N_2562,N_1340,N_616);
nor U2563 (N_2563,N_2456,N_475);
or U2564 (N_2564,N_880,N_1142);
nand U2565 (N_2565,N_1817,N_1741);
nor U2566 (N_2566,N_1950,N_2190);
and U2567 (N_2567,N_1800,N_2486);
and U2568 (N_2568,N_1999,N_1587);
or U2569 (N_2569,N_1292,N_449);
nor U2570 (N_2570,N_1768,N_141);
or U2571 (N_2571,N_1827,N_388);
nor U2572 (N_2572,N_1141,N_959);
and U2573 (N_2573,N_417,N_741);
nor U2574 (N_2574,N_573,N_831);
nor U2575 (N_2575,N_1505,N_1021);
or U2576 (N_2576,N_169,N_135);
nor U2577 (N_2577,N_1145,N_505);
nand U2578 (N_2578,N_2093,N_1772);
or U2579 (N_2579,N_83,N_1383);
or U2580 (N_2580,N_2054,N_1644);
nor U2581 (N_2581,N_2181,N_968);
and U2582 (N_2582,N_1542,N_2255);
and U2583 (N_2583,N_1696,N_70);
nand U2584 (N_2584,N_1460,N_1004);
nand U2585 (N_2585,N_2328,N_1735);
or U2586 (N_2586,N_617,N_1738);
and U2587 (N_2587,N_1879,N_2392);
or U2588 (N_2588,N_2056,N_1596);
nor U2589 (N_2589,N_1220,N_300);
and U2590 (N_2590,N_1305,N_986);
nor U2591 (N_2591,N_1514,N_2141);
or U2592 (N_2592,N_853,N_1482);
or U2593 (N_2593,N_291,N_348);
and U2594 (N_2594,N_2312,N_1198);
and U2595 (N_2595,N_121,N_949);
nor U2596 (N_2596,N_466,N_276);
nor U2597 (N_2597,N_1938,N_1439);
and U2598 (N_2598,N_128,N_1752);
and U2599 (N_2599,N_230,N_1391);
nor U2600 (N_2600,N_1604,N_1881);
nor U2601 (N_2601,N_2262,N_1312);
and U2602 (N_2602,N_1589,N_36);
and U2603 (N_2603,N_948,N_767);
nand U2604 (N_2604,N_1027,N_2434);
nor U2605 (N_2605,N_2263,N_1760);
nor U2606 (N_2606,N_512,N_2250);
nor U2607 (N_2607,N_1086,N_2061);
or U2608 (N_2608,N_654,N_1233);
nand U2609 (N_2609,N_491,N_400);
nand U2610 (N_2610,N_782,N_2460);
nand U2611 (N_2611,N_601,N_2103);
nand U2612 (N_2612,N_1899,N_972);
nand U2613 (N_2613,N_1964,N_1012);
and U2614 (N_2614,N_1642,N_1409);
nor U2615 (N_2615,N_2068,N_241);
nand U2616 (N_2616,N_1958,N_85);
and U2617 (N_2617,N_843,N_2083);
nand U2618 (N_2618,N_150,N_2446);
and U2619 (N_2619,N_2325,N_1736);
or U2620 (N_2620,N_1427,N_1921);
and U2621 (N_2621,N_556,N_1766);
and U2622 (N_2622,N_484,N_1013);
or U2623 (N_2623,N_1934,N_2030);
and U2624 (N_2624,N_1240,N_1339);
and U2625 (N_2625,N_1619,N_2310);
nor U2626 (N_2626,N_1538,N_1911);
nor U2627 (N_2627,N_1985,N_1238);
and U2628 (N_2628,N_1727,N_1605);
nand U2629 (N_2629,N_1424,N_794);
and U2630 (N_2630,N_334,N_643);
or U2631 (N_2631,N_738,N_943);
or U2632 (N_2632,N_1419,N_1987);
nand U2633 (N_2633,N_82,N_1906);
nand U2634 (N_2634,N_1762,N_131);
nor U2635 (N_2635,N_69,N_1936);
nor U2636 (N_2636,N_1330,N_515);
and U2637 (N_2637,N_421,N_1040);
nor U2638 (N_2638,N_66,N_1343);
nand U2639 (N_2639,N_2352,N_1792);
nor U2640 (N_2640,N_2331,N_2040);
and U2641 (N_2641,N_932,N_989);
nand U2642 (N_2642,N_2413,N_1133);
nor U2643 (N_2643,N_1437,N_758);
and U2644 (N_2644,N_1321,N_980);
or U2645 (N_2645,N_637,N_1204);
or U2646 (N_2646,N_1010,N_1519);
nor U2647 (N_2647,N_136,N_1668);
nor U2648 (N_2648,N_1652,N_149);
and U2649 (N_2649,N_50,N_1749);
nor U2650 (N_2650,N_236,N_224);
nand U2651 (N_2651,N_1532,N_2300);
nor U2652 (N_2652,N_1663,N_447);
nand U2653 (N_2653,N_946,N_593);
or U2654 (N_2654,N_960,N_2080);
nand U2655 (N_2655,N_1353,N_707);
nor U2656 (N_2656,N_1568,N_2088);
and U2657 (N_2657,N_577,N_1867);
and U2658 (N_2658,N_825,N_728);
nand U2659 (N_2659,N_1135,N_1359);
nor U2660 (N_2660,N_2277,N_2005);
or U2661 (N_2661,N_1059,N_842);
and U2662 (N_2662,N_2069,N_542);
nand U2663 (N_2663,N_756,N_1929);
or U2664 (N_2664,N_2058,N_2495);
nor U2665 (N_2665,N_202,N_581);
nor U2666 (N_2666,N_877,N_39);
nor U2667 (N_2667,N_130,N_270);
nor U2668 (N_2668,N_1694,N_771);
or U2669 (N_2669,N_343,N_1733);
nand U2670 (N_2670,N_391,N_267);
nand U2671 (N_2671,N_438,N_1835);
or U2672 (N_2672,N_1372,N_439);
or U2673 (N_2673,N_839,N_2391);
nor U2674 (N_2674,N_2194,N_2299);
nor U2675 (N_2675,N_1091,N_999);
and U2676 (N_2676,N_440,N_1869);
nor U2677 (N_2677,N_1789,N_194);
or U2678 (N_2678,N_1551,N_2438);
or U2679 (N_2679,N_2454,N_1252);
and U2680 (N_2680,N_1513,N_2119);
or U2681 (N_2681,N_2109,N_1775);
and U2682 (N_2682,N_1674,N_1493);
and U2683 (N_2683,N_1952,N_88);
and U2684 (N_2684,N_1527,N_907);
nand U2685 (N_2685,N_249,N_409);
or U2686 (N_2686,N_614,N_514);
or U2687 (N_2687,N_1748,N_1063);
or U2688 (N_2688,N_536,N_882);
and U2689 (N_2689,N_757,N_1125);
nor U2690 (N_2690,N_1601,N_2304);
and U2691 (N_2691,N_2002,N_1639);
nand U2692 (N_2692,N_1349,N_64);
nor U2693 (N_2693,N_1011,N_1347);
and U2694 (N_2694,N_2335,N_2252);
nor U2695 (N_2695,N_1915,N_2354);
nor U2696 (N_2696,N_1307,N_2306);
and U2697 (N_2697,N_1018,N_1611);
nand U2698 (N_2698,N_1803,N_1352);
nand U2699 (N_2699,N_2195,N_1034);
nand U2700 (N_2700,N_620,N_390);
or U2701 (N_2701,N_2117,N_2322);
nor U2702 (N_2702,N_330,N_1426);
nand U2703 (N_2703,N_1345,N_1476);
nand U2704 (N_2704,N_1089,N_2369);
nor U2705 (N_2705,N_431,N_1032);
and U2706 (N_2706,N_1435,N_679);
or U2707 (N_2707,N_55,N_1837);
and U2708 (N_2708,N_173,N_214);
and U2709 (N_2709,N_2465,N_144);
and U2710 (N_2710,N_27,N_1311);
and U2711 (N_2711,N_171,N_1787);
nand U2712 (N_2712,N_2246,N_1386);
or U2713 (N_2713,N_1284,N_368);
and U2714 (N_2714,N_233,N_1057);
nor U2715 (N_2715,N_2313,N_1315);
nor U2716 (N_2716,N_25,N_711);
xnor U2717 (N_2717,N_2275,N_364);
nor U2718 (N_2718,N_2216,N_2267);
nor U2719 (N_2719,N_1512,N_806);
or U2720 (N_2720,N_786,N_613);
and U2721 (N_2721,N_1515,N_37);
and U2722 (N_2722,N_1385,N_2445);
and U2723 (N_2723,N_687,N_1959);
and U2724 (N_2724,N_1042,N_648);
nor U2725 (N_2725,N_966,N_460);
or U2726 (N_2726,N_1861,N_685);
and U2727 (N_2727,N_294,N_2100);
nand U2728 (N_2728,N_988,N_1393);
or U2729 (N_2729,N_146,N_2453);
nand U2730 (N_2730,N_1747,N_1989);
nand U2731 (N_2731,N_32,N_2143);
nand U2732 (N_2732,N_2382,N_1667);
nand U2733 (N_2733,N_1813,N_809);
and U2734 (N_2734,N_2180,N_1509);
nand U2735 (N_2735,N_2214,N_2390);
xor U2736 (N_2736,N_470,N_48);
nor U2737 (N_2737,N_369,N_418);
or U2738 (N_2738,N_805,N_862);
or U2739 (N_2739,N_2042,N_1797);
or U2740 (N_2740,N_2210,N_20);
and U2741 (N_2741,N_2311,N_2218);
nand U2742 (N_2742,N_1722,N_697);
or U2743 (N_2743,N_1388,N_327);
nand U2744 (N_2744,N_1628,N_1773);
and U2745 (N_2745,N_1606,N_1061);
or U2746 (N_2746,N_2464,N_2025);
or U2747 (N_2747,N_1249,N_925);
nand U2748 (N_2748,N_1382,N_795);
or U2749 (N_2749,N_1428,N_1912);
nor U2750 (N_2750,N_2474,N_2102);
nand U2751 (N_2751,N_1456,N_1648);
nor U2752 (N_2752,N_1276,N_963);
or U2753 (N_2753,N_385,N_1591);
and U2754 (N_2754,N_2108,N_921);
nor U2755 (N_2755,N_1705,N_624);
or U2756 (N_2756,N_2288,N_1054);
or U2757 (N_2757,N_521,N_2321);
and U2758 (N_2758,N_2215,N_2326);
and U2759 (N_2759,N_1173,N_1151);
and U2760 (N_2760,N_186,N_1804);
and U2761 (N_2761,N_2185,N_307);
nand U2762 (N_2762,N_2193,N_635);
and U2763 (N_2763,N_646,N_543);
nand U2764 (N_2764,N_815,N_626);
or U2765 (N_2765,N_2235,N_1784);
nor U2766 (N_2766,N_1718,N_1396);
and U2767 (N_2767,N_340,N_2477);
nor U2768 (N_2768,N_1440,N_991);
and U2769 (N_2769,N_2363,N_1554);
nand U2770 (N_2770,N_112,N_234);
nor U2771 (N_2771,N_970,N_1701);
nand U2772 (N_2772,N_2443,N_1847);
nor U2773 (N_2773,N_269,N_1210);
nor U2774 (N_2774,N_1556,N_1935);
nand U2775 (N_2775,N_535,N_2118);
or U2776 (N_2776,N_665,N_676);
and U2777 (N_2777,N_399,N_1698);
nand U2778 (N_2778,N_90,N_1399);
nand U2779 (N_2779,N_2237,N_1602);
nor U2780 (N_2780,N_325,N_2023);
or U2781 (N_2781,N_664,N_450);
or U2782 (N_2782,N_47,N_906);
nand U2783 (N_2783,N_1671,N_1090);
or U2784 (N_2784,N_2442,N_1660);
nor U2785 (N_2785,N_1043,N_288);
and U2786 (N_2786,N_2082,N_1285);
nand U2787 (N_2787,N_326,N_481);
nor U2788 (N_2788,N_821,N_178);
nand U2789 (N_2789,N_2155,N_1270);
nand U2790 (N_2790,N_663,N_1992);
nor U2791 (N_2791,N_323,N_1214);
or U2792 (N_2792,N_80,N_1932);
and U2793 (N_2793,N_378,N_2047);
nor U2794 (N_2794,N_1387,N_539);
nor U2795 (N_2795,N_702,N_1306);
and U2796 (N_2796,N_253,N_1155);
or U2797 (N_2797,N_336,N_2245);
and U2798 (N_2798,N_2279,N_142);
nand U2799 (N_2799,N_386,N_2254);
or U2800 (N_2800,N_918,N_108);
nand U2801 (N_2801,N_1597,N_1661);
nor U2802 (N_2802,N_1711,N_1451);
and U2803 (N_2803,N_1213,N_2213);
and U2804 (N_2804,N_537,N_1260);
nand U2805 (N_2805,N_791,N_2400);
or U2806 (N_2806,N_212,N_259);
or U2807 (N_2807,N_1469,N_1461);
nor U2808 (N_2808,N_1433,N_1096);
nand U2809 (N_2809,N_1231,N_1949);
and U2810 (N_2810,N_208,N_1993);
and U2811 (N_2811,N_1230,N_7);
nand U2812 (N_2812,N_2243,N_2290);
nor U2813 (N_2813,N_1153,N_122);
nor U2814 (N_2814,N_2222,N_1094);
nor U2815 (N_2815,N_1258,N_84);
nor U2816 (N_2816,N_1250,N_2482);
nand U2817 (N_2817,N_1067,N_525);
nand U2818 (N_2818,N_860,N_863);
and U2819 (N_2819,N_1444,N_1022);
or U2820 (N_2820,N_690,N_352);
and U2821 (N_2821,N_902,N_1531);
nand U2822 (N_2822,N_2285,N_2203);
and U2823 (N_2823,N_2086,N_506);
or U2824 (N_2824,N_2050,N_358);
or U2825 (N_2825,N_1518,N_21);
nand U2826 (N_2826,N_819,N_997);
nor U2827 (N_2827,N_1805,N_519);
and U2828 (N_2828,N_100,N_777);
and U2829 (N_2829,N_101,N_594);
nand U2830 (N_2830,N_2406,N_2449);
nand U2831 (N_2831,N_1009,N_1574);
nor U2832 (N_2832,N_680,N_721);
and U2833 (N_2833,N_723,N_1095);
and U2834 (N_2834,N_2116,N_396);
and U2835 (N_2835,N_1712,N_2319);
and U2836 (N_2836,N_2340,N_2172);
and U2837 (N_2837,N_1986,N_684);
nor U2838 (N_2838,N_255,N_844);
nand U2839 (N_2839,N_172,N_226);
and U2840 (N_2840,N_2457,N_2000);
nand U2841 (N_2841,N_1314,N_1177);
and U2842 (N_2842,N_1970,N_776);
nor U2843 (N_2843,N_205,N_2269);
nor U2844 (N_2844,N_1112,N_1783);
nor U2845 (N_2845,N_2436,N_1066);
and U2846 (N_2846,N_92,N_1833);
nand U2847 (N_2847,N_1281,N_145);
nand U2848 (N_2848,N_1109,N_79);
or U2849 (N_2849,N_1486,N_1273);
nand U2850 (N_2850,N_893,N_1062);
and U2851 (N_2851,N_204,N_2149);
nor U2852 (N_2852,N_1030,N_1008);
and U2853 (N_2853,N_1612,N_744);
nand U2854 (N_2854,N_2168,N_304);
or U2855 (N_2855,N_901,N_554);
and U2856 (N_2856,N_1139,N_1002);
or U2857 (N_2857,N_2271,N_2280);
nor U2858 (N_2858,N_1348,N_1955);
nor U2859 (N_2859,N_1007,N_764);
and U2860 (N_2860,N_2175,N_1689);
nor U2861 (N_2861,N_1378,N_2142);
xor U2862 (N_2862,N_887,N_1684);
nand U2863 (N_2863,N_72,N_847);
and U2864 (N_2864,N_2156,N_1560);
nand U2865 (N_2865,N_770,N_1719);
or U2866 (N_2866,N_179,N_29);
nor U2867 (N_2867,N_1332,N_2355);
and U2868 (N_2868,N_864,N_846);
nand U2869 (N_2869,N_435,N_467);
and U2870 (N_2870,N_1650,N_1319);
nor U2871 (N_2871,N_2414,N_2341);
nor U2872 (N_2872,N_780,N_2238);
nand U2873 (N_2873,N_1170,N_278);
and U2874 (N_2874,N_2053,N_2140);
and U2875 (N_2875,N_1380,N_1453);
or U2876 (N_2876,N_1819,N_800);
nor U2877 (N_2877,N_1761,N_2138);
nor U2878 (N_2878,N_920,N_31);
and U2879 (N_2879,N_58,N_1885);
and U2880 (N_2880,N_2295,N_1076);
or U2881 (N_2881,N_110,N_2492);
and U2882 (N_2882,N_1164,N_2033);
nand U2883 (N_2883,N_2121,N_430);
or U2884 (N_2884,N_1816,N_2158);
nand U2885 (N_2885,N_718,N_1685);
nand U2886 (N_2886,N_2129,N_2373);
nand U2887 (N_2887,N_1501,N_2095);
nand U2888 (N_2888,N_2408,N_1093);
and U2889 (N_2889,N_871,N_1373);
nand U2890 (N_2890,N_1294,N_1140);
or U2891 (N_2891,N_567,N_1156);
nand U2892 (N_2892,N_2303,N_730);
and U2893 (N_2893,N_2127,N_332);
nor U2894 (N_2894,N_810,N_879);
and U2895 (N_2895,N_631,N_1079);
nand U2896 (N_2896,N_1852,N_461);
and U2897 (N_2897,N_1810,N_1529);
nor U2898 (N_2898,N_1209,N_242);
nor U2899 (N_2899,N_2494,N_2051);
and U2900 (N_2900,N_2012,N_1438);
nand U2901 (N_2901,N_1743,N_94);
and U2902 (N_2902,N_404,N_883);
nor U2903 (N_2903,N_2327,N_1739);
and U2904 (N_2904,N_1892,N_1189);
nand U2905 (N_2905,N_1019,N_297);
and U2906 (N_2906,N_1863,N_61);
nand U2907 (N_2907,N_950,N_1997);
nand U2908 (N_2908,N_1297,N_751);
or U2909 (N_2909,N_2298,N_781);
or U2910 (N_2910,N_1483,N_1180);
and U2911 (N_2911,N_432,N_841);
nor U2912 (N_2912,N_517,N_1105);
nor U2913 (N_2913,N_1864,N_1045);
nor U2914 (N_2914,N_649,N_1510);
nor U2915 (N_2915,N_497,N_1854);
nand U2916 (N_2916,N_1295,N_397);
or U2917 (N_2917,N_2130,N_715);
or U2918 (N_2918,N_1248,N_207);
nand U2919 (N_2919,N_588,N_1473);
or U2920 (N_2920,N_1244,N_63);
or U2921 (N_2921,N_1812,N_1676);
or U2922 (N_2922,N_1822,N_2404);
and U2923 (N_2923,N_116,N_1261);
or U2924 (N_2924,N_1025,N_886);
nand U2925 (N_2925,N_722,N_984);
and U2926 (N_2926,N_971,N_2405);
or U2927 (N_2927,N_1508,N_1496);
and U2928 (N_2928,N_2366,N_696);
or U2929 (N_2929,N_219,N_1005);
and U2930 (N_2930,N_1082,N_1099);
or U2931 (N_2931,N_1836,N_1237);
nor U2932 (N_2932,N_884,N_1777);
and U2933 (N_2933,N_1114,N_1313);
or U2934 (N_2934,N_1317,N_1669);
or U2935 (N_2935,N_1651,N_243);
or U2936 (N_2936,N_1037,N_2432);
nor U2937 (N_2937,N_628,N_56);
and U2938 (N_2938,N_2397,N_344);
or U2939 (N_2939,N_2380,N_1415);
nor U2940 (N_2940,N_1298,N_2330);
and U2941 (N_2941,N_1147,N_745);
and U2942 (N_2942,N_1582,N_246);
and U2943 (N_2943,N_35,N_2283);
or U2944 (N_2944,N_2375,N_1750);
nor U2945 (N_2945,N_1790,N_2151);
nand U2946 (N_2946,N_1050,N_1215);
and U2947 (N_2947,N_2,N_444);
and U2948 (N_2948,N_252,N_0);
nand U2949 (N_2949,N_2052,N_739);
nor U2950 (N_2950,N_1251,N_1354);
and U2951 (N_2951,N_1729,N_314);
or U2952 (N_2952,N_1916,N_945);
and U2953 (N_2953,N_1730,N_610);
xor U2954 (N_2954,N_1679,N_1342);
or U2955 (N_2955,N_666,N_454);
or U2956 (N_2956,N_1890,N_1664);
nor U2957 (N_2957,N_2472,N_1579);
nand U2958 (N_2958,N_716,N_2324);
and U2959 (N_2959,N_313,N_2010);
nand U2960 (N_2960,N_2379,N_271);
nand U2961 (N_2961,N_2094,N_2323);
and U2962 (N_2962,N_1896,N_134);
and U2963 (N_2963,N_2276,N_456);
or U2964 (N_2964,N_290,N_489);
and U2965 (N_2965,N_2258,N_1982);
and U2966 (N_2966,N_2125,N_870);
or U2967 (N_2967,N_2435,N_1229);
or U2968 (N_2968,N_892,N_2307);
nor U2969 (N_2969,N_1422,N_1181);
and U2970 (N_2970,N_1595,N_592);
nor U2971 (N_2971,N_4,N_1000);
nand U2972 (N_2972,N_912,N_1759);
xnor U2973 (N_2973,N_1530,N_283);
nand U2974 (N_2974,N_1925,N_42);
or U2975 (N_2975,N_608,N_857);
xnor U2976 (N_2976,N_1980,N_261);
and U2977 (N_2977,N_2332,N_191);
nand U2978 (N_2978,N_2420,N_2192);
and U2979 (N_2979,N_522,N_3);
or U2980 (N_2980,N_1406,N_693);
or U2981 (N_2981,N_425,N_1341);
and U2982 (N_2982,N_900,N_1755);
or U2983 (N_2983,N_155,N_1583);
or U2984 (N_2984,N_670,N_1465);
or U2985 (N_2985,N_1526,N_1316);
nor U2986 (N_2986,N_1367,N_2349);
or U2987 (N_2987,N_762,N_909);
or U2988 (N_2988,N_2187,N_365);
or U2989 (N_2989,N_408,N_2334);
or U2990 (N_2990,N_813,N_811);
or U2991 (N_2991,N_1256,N_899);
or U2992 (N_2992,N_660,N_1878);
or U2993 (N_2993,N_2133,N_2440);
xor U2994 (N_2994,N_1824,N_1889);
nand U2995 (N_2995,N_1268,N_599);
nand U2996 (N_2996,N_732,N_1417);
nand U2997 (N_2997,N_1038,N_941);
and U2998 (N_2998,N_1255,N_1576);
or U2999 (N_2999,N_99,N_2249);
or U3000 (N_3000,N_2459,N_1706);
or U3001 (N_3001,N_1163,N_2476);
and U3002 (N_3002,N_1859,N_196);
nand U3003 (N_3003,N_1570,N_1247);
and U3004 (N_3004,N_1904,N_2320);
nor U3005 (N_3005,N_1566,N_1905);
nand U3006 (N_3006,N_2266,N_2176);
and U3007 (N_3007,N_705,N_392);
and U3008 (N_3008,N_1933,N_737);
nor U3009 (N_3009,N_1121,N_978);
nand U3010 (N_3010,N_414,N_2347);
nand U3011 (N_3011,N_286,N_2428);
and U3012 (N_3012,N_1516,N_1647);
nor U3013 (N_3013,N_2233,N_1106);
nand U3014 (N_3014,N_2227,N_1102);
or U3015 (N_3015,N_1969,N_558);
or U3016 (N_3016,N_2361,N_2171);
nand U3017 (N_3017,N_476,N_623);
nor U3018 (N_3018,N_976,N_324);
nor U3019 (N_3019,N_163,N_1331);
and U3020 (N_3020,N_1463,N_2264);
nand U3021 (N_3021,N_2131,N_1413);
or U3022 (N_3022,N_674,N_1920);
nor U3023 (N_3023,N_894,N_322);
and U3024 (N_3024,N_2212,N_372);
or U3025 (N_3025,N_869,N_861);
nand U3026 (N_3026,N_211,N_985);
nand U3027 (N_3027,N_1400,N_1838);
or U3028 (N_3028,N_49,N_2074);
or U3029 (N_3029,N_1211,N_2106);
or U3030 (N_3030,N_2076,N_1732);
and U3031 (N_3031,N_2225,N_694);
nand U3032 (N_3032,N_2153,N_19);
or U3033 (N_3033,N_2282,N_1471);
and U3034 (N_3034,N_2229,N_1618);
nor U3035 (N_3035,N_1795,N_2006);
or U3036 (N_3036,N_875,N_1290);
nand U3037 (N_3037,N_1449,N_1555);
nand U3038 (N_3038,N_401,N_546);
nor U3039 (N_3039,N_105,N_858);
or U3040 (N_3040,N_1363,N_994);
and U3041 (N_3041,N_889,N_2236);
and U3042 (N_3042,N_223,N_272);
nand U3043 (N_3043,N_1222,N_1682);
nand U3044 (N_3044,N_1965,N_427);
or U3045 (N_3045,N_445,N_2378);
nor U3046 (N_3046,N_2139,N_1876);
and U3047 (N_3047,N_589,N_1080);
nor U3048 (N_3048,N_1418,N_1502);
nand U3049 (N_3049,N_457,N_2113);
or U3050 (N_3050,N_897,N_2090);
nor U3051 (N_3051,N_2305,N_1271);
and U3052 (N_3052,N_1272,N_1267);
nand U3053 (N_3053,N_1159,N_428);
or U3054 (N_3054,N_1624,N_15);
and U3055 (N_3055,N_1423,N_1464);
or U3056 (N_3056,N_1857,N_477);
nand U3057 (N_3057,N_1908,N_133);
nand U3058 (N_3058,N_1455,N_793);
nor U3059 (N_3059,N_2022,N_258);
xor U3060 (N_3060,N_2032,N_1179);
or U3061 (N_3061,N_612,N_1084);
or U3062 (N_3062,N_691,N_905);
nand U3063 (N_3063,N_1742,N_695);
nor U3064 (N_3064,N_2475,N_1448);
nor U3065 (N_3065,N_659,N_420);
nand U3066 (N_3066,N_1636,N_1737);
nand U3067 (N_3067,N_2385,N_509);
or U3068 (N_3068,N_156,N_1829);
or U3069 (N_3069,N_2173,N_499);
nand U3070 (N_3070,N_109,N_2207);
and U3071 (N_3071,N_1128,N_2164);
nor U3072 (N_3072,N_1988,N_655);
and U3073 (N_3073,N_2197,N_2008);
and U3074 (N_3074,N_441,N_1183);
and U3075 (N_3075,N_1765,N_1984);
nor U3076 (N_3076,N_914,N_532);
nor U3077 (N_3077,N_1780,N_1280);
nor U3078 (N_3078,N_328,N_357);
xnor U3079 (N_3079,N_1446,N_538);
and U3080 (N_3080,N_797,N_2407);
xor U3081 (N_3081,N_607,N_1097);
or U3082 (N_3082,N_1443,N_720);
or U3083 (N_3083,N_337,N_2230);
and U3084 (N_3084,N_1543,N_174);
and U3085 (N_3085,N_557,N_295);
and U3086 (N_3086,N_1425,N_1641);
and U3087 (N_3087,N_180,N_1728);
and U3088 (N_3088,N_840,N_2048);
nor U3089 (N_3089,N_1117,N_1633);
or U3090 (N_3090,N_1283,N_2152);
nand U3091 (N_3091,N_2417,N_785);
nand U3092 (N_3092,N_1776,N_2199);
nand U3093 (N_3093,N_1182,N_1707);
nor U3094 (N_3094,N_1416,N_2487);
or U3095 (N_3095,N_474,N_264);
or U3096 (N_3096,N_292,N_768);
and U3097 (N_3097,N_1188,N_500);
nand U3098 (N_3098,N_1174,N_422);
and U3099 (N_3099,N_1462,N_1673);
nand U3100 (N_3100,N_958,N_1654);
or U3101 (N_3101,N_856,N_625);
and U3102 (N_3102,N_1392,N_1593);
and U3103 (N_3103,N_530,N_706);
or U3104 (N_3104,N_579,N_1048);
or U3105 (N_3105,N_2089,N_1724);
nor U3106 (N_3106,N_1630,N_855);
or U3107 (N_3107,N_823,N_1942);
and U3108 (N_3108,N_656,N_1645);
nor U3109 (N_3109,N_2162,N_1242);
nand U3110 (N_3110,N_2433,N_829);
and U3111 (N_3111,N_1715,N_2493);
and U3112 (N_3112,N_1414,N_487);
and U3113 (N_3113,N_1764,N_2274);
nor U3114 (N_3114,N_248,N_2384);
nand U3115 (N_3115,N_1171,N_1323);
or U3116 (N_3116,N_2287,N_1662);
nor U3117 (N_3117,N_1594,N_463);
nor U3118 (N_3118,N_1620,N_2289);
nand U3119 (N_3119,N_265,N_1973);
nor U3120 (N_3120,N_1303,N_2196);
nand U3121 (N_3121,N_570,N_1223);
nand U3122 (N_3122,N_1845,N_1113);
nor U3123 (N_3123,N_1368,N_1404);
and U3124 (N_3124,N_735,N_492);
and U3125 (N_3125,N_341,N_584);
nor U3126 (N_3126,N_792,N_1577);
nor U3127 (N_3127,N_1592,N_1598);
or U3128 (N_3128,N_192,N_2178);
and U3129 (N_3129,N_465,N_1108);
nand U3130 (N_3130,N_1895,N_2293);
and U3131 (N_3131,N_485,N_77);
nand U3132 (N_3132,N_274,N_1293);
nand U3133 (N_3133,N_1394,N_289);
nor U3134 (N_3134,N_602,N_1146);
nor U3135 (N_3135,N_1713,N_2223);
nor U3136 (N_3136,N_2367,N_2483);
xnor U3137 (N_3137,N_1931,N_898);
or U3138 (N_3138,N_154,N_320);
and U3139 (N_3139,N_1480,N_1544);
and U3140 (N_3140,N_2372,N_1700);
nor U3141 (N_3141,N_1866,N_1870);
or U3142 (N_3142,N_1266,N_2296);
nand U3143 (N_3143,N_866,N_2421);
nand U3144 (N_3144,N_1410,N_170);
nor U3145 (N_3145,N_891,N_1055);
nor U3146 (N_3146,N_1226,N_1278);
nor U3147 (N_3147,N_2186,N_1600);
xnor U3148 (N_3148,N_310,N_818);
or U3149 (N_3149,N_634,N_2231);
and U3150 (N_3150,N_1855,N_1994);
or U3151 (N_3151,N_2003,N_2018);
and U3152 (N_3152,N_115,N_2150);
and U3153 (N_3153,N_1882,N_68);
and U3154 (N_3154,N_559,N_1122);
nand U3155 (N_3155,N_1049,N_293);
nor U3156 (N_3156,N_493,N_302);
nor U3157 (N_3157,N_2468,N_583);
nand U3158 (N_3158,N_1550,N_2120);
and U3159 (N_3159,N_2302,N_1088);
nor U3160 (N_3160,N_1160,N_2177);
or U3161 (N_3161,N_571,N_1447);
and U3162 (N_3162,N_854,N_6);
nand U3163 (N_3163,N_2394,N_1186);
or U3164 (N_3164,N_43,N_1672);
nand U3165 (N_3165,N_381,N_382);
nor U3166 (N_3166,N_239,N_1902);
or U3167 (N_3167,N_647,N_1785);
and U3168 (N_3168,N_1763,N_633);
or U3169 (N_3169,N_52,N_2301);
or U3170 (N_3170,N_1035,N_1756);
nor U3171 (N_3171,N_1793,N_2037);
nor U3172 (N_3172,N_2467,N_2470);
nor U3173 (N_3173,N_2358,N_749);
nand U3174 (N_3174,N_1873,N_471);
and U3175 (N_3175,N_1277,N_1001);
nand U3176 (N_3176,N_1167,N_916);
and U3177 (N_3177,N_1071,N_473);
nand U3178 (N_3178,N_2224,N_342);
nor U3179 (N_3179,N_1152,N_1865);
nand U3180 (N_3180,N_423,N_2403);
and U3181 (N_3181,N_177,N_2345);
or U3182 (N_3182,N_2374,N_183);
or U3183 (N_3183,N_416,N_1384);
nor U3184 (N_3184,N_2107,N_1477);
and U3185 (N_3185,N_2067,N_1334);
nand U3186 (N_3186,N_393,N_498);
or U3187 (N_3187,N_1585,N_1176);
nor U3188 (N_3188,N_2122,N_565);
or U3189 (N_3189,N_221,N_362);
nand U3190 (N_3190,N_376,N_2418);
or U3191 (N_3191,N_1395,N_1886);
nand U3192 (N_3192,N_2273,N_1939);
and U3193 (N_3193,N_188,N_746);
and U3194 (N_3194,N_510,N_2239);
or U3195 (N_3195,N_1910,N_1310);
nand U3196 (N_3196,N_931,N_951);
and U3197 (N_3197,N_2166,N_501);
nor U3198 (N_3198,N_200,N_2478);
nand U3199 (N_3199,N_548,N_2059);
nor U3200 (N_3200,N_1903,N_2104);
or U3201 (N_3201,N_553,N_318);
nand U3202 (N_3202,N_979,N_402);
and U3203 (N_3203,N_13,N_692);
nand U3204 (N_3204,N_2339,N_1123);
or U3205 (N_3205,N_1665,N_868);
or U3206 (N_3206,N_713,N_1017);
and U3207 (N_3207,N_1524,N_2427);
nand U3208 (N_3208,N_1617,N_1162);
nor U3209 (N_3209,N_1740,N_263);
or U3210 (N_3210,N_1407,N_719);
nor U3211 (N_3211,N_2201,N_1875);
and U3212 (N_3212,N_1607,N_816);
and U3213 (N_3213,N_1913,N_911);
nor U3214 (N_3214,N_1967,N_2081);
or U3215 (N_3215,N_1690,N_545);
nand U3216 (N_3216,N_835,N_2169);
or U3217 (N_3217,N_2007,N_1432);
or U3218 (N_3218,N_1721,N_2057);
or U3219 (N_3219,N_560,N_644);
and U3220 (N_3220,N_2294,N_653);
and U3221 (N_3221,N_209,N_1521);
and U3222 (N_3222,N_740,N_1127);
nand U3223 (N_3223,N_1143,N_2473);
nor U3224 (N_3224,N_2135,N_1945);
nand U3225 (N_3225,N_572,N_2444);
and U3226 (N_3226,N_1130,N_1033);
or U3227 (N_3227,N_1111,N_1475);
nor U3228 (N_3228,N_247,N_2371);
and U3229 (N_3229,N_1445,N_2217);
nor U3230 (N_3230,N_987,N_1085);
and U3231 (N_3231,N_458,N_1137);
or U3232 (N_3232,N_516,N_2348);
nand U3233 (N_3233,N_1946,N_1734);
or U3234 (N_3234,N_1553,N_1485);
nand U3235 (N_3235,N_672,N_1629);
nor U3236 (N_3236,N_95,N_2448);
nor U3237 (N_3237,N_1028,N_1257);
and U3238 (N_3238,N_1528,N_2309);
and U3239 (N_3239,N_1402,N_1900);
and U3240 (N_3240,N_2211,N_671);
or U3241 (N_3241,N_924,N_836);
or U3242 (N_3242,N_303,N_2362);
nand U3243 (N_3243,N_503,N_14);
and U3244 (N_3244,N_1975,N_919);
nand U3245 (N_3245,N_1241,N_677);
xnor U3246 (N_3246,N_1129,N_1815);
or U3247 (N_3247,N_67,N_1914);
and U3248 (N_3248,N_285,N_1205);
nor U3249 (N_3249,N_2087,N_103);
and U3250 (N_3250,N_2011,N_2046);
nand U3251 (N_3251,N_2179,N_954);
nor U3252 (N_3252,N_359,N_1771);
or U3253 (N_3253,N_927,N_251);
or U3254 (N_3254,N_217,N_2029);
and U3255 (N_3255,N_117,N_411);
nor U3256 (N_3256,N_213,N_2208);
or U3257 (N_3257,N_1814,N_1263);
or U3258 (N_3258,N_1825,N_23);
nand U3259 (N_3259,N_2147,N_240);
nor U3260 (N_3260,N_380,N_339);
or U3261 (N_3261,N_2062,N_2383);
nand U3262 (N_3262,N_1195,N_2401);
or U3263 (N_3263,N_2429,N_22);
and U3264 (N_3264,N_1161,N_2450);
nand U3265 (N_3265,N_1228,N_1458);
nand U3266 (N_3266,N_1523,N_704);
and U3267 (N_3267,N_2049,N_1943);
or U3268 (N_3268,N_1545,N_1782);
nand U3269 (N_3269,N_1723,N_586);
nor U3270 (N_3270,N_689,N_686);
or U3271 (N_3271,N_496,N_1300);
or U3272 (N_3272,N_1930,N_1725);
nand U3273 (N_3273,N_947,N_621);
or U3274 (N_3274,N_446,N_1802);
nor U3275 (N_3275,N_549,N_642);
or U3276 (N_3276,N_890,N_2342);
or U3277 (N_3277,N_1390,N_1041);
and U3278 (N_3278,N_1898,N_1631);
or U3279 (N_3279,N_1794,N_2416);
nor U3280 (N_3280,N_1695,N_308);
nor U3281 (N_3281,N_504,N_563);
nor U3282 (N_3282,N_1610,N_2471);
nor U3283 (N_3283,N_1218,N_353);
and U3284 (N_3284,N_2337,N_775);
and U3285 (N_3285,N_1693,N_1064);
nor U3286 (N_3286,N_830,N_1291);
nor U3287 (N_3287,N_165,N_254);
nand U3288 (N_3288,N_1279,N_1703);
nand U3289 (N_3289,N_2073,N_956);
or U3290 (N_3290,N_1087,N_462);
and U3291 (N_3291,N_773,N_1441);
nor U3292 (N_3292,N_1632,N_215);
or U3293 (N_3293,N_1288,N_2228);
nor U3294 (N_3294,N_284,N_218);
nand U3295 (N_3295,N_1562,N_1184);
and U3296 (N_3296,N_1704,N_1951);
or U3297 (N_3297,N_273,N_1408);
nand U3298 (N_3298,N_658,N_1118);
nor U3299 (N_3299,N_210,N_561);
nand U3300 (N_3300,N_1767,N_1172);
and U3301 (N_3301,N_190,N_316);
or U3302 (N_3302,N_1058,N_784);
or U3303 (N_3303,N_804,N_1232);
and U3304 (N_3304,N_1236,N_1874);
nor U3305 (N_3305,N_928,N_2065);
and U3306 (N_3306,N_1686,N_1016);
nand U3307 (N_3307,N_2458,N_1893);
xnor U3308 (N_3308,N_1586,N_437);
nor U3309 (N_3309,N_2270,N_657);
nand U3310 (N_3310,N_1197,N_2016);
and U3311 (N_3311,N_1274,N_387);
nand U3312 (N_3312,N_2071,N_859);
or U3313 (N_3313,N_1149,N_2044);
and U3314 (N_3314,N_2419,N_2020);
nand U3315 (N_3315,N_451,N_442);
nor U3316 (N_3316,N_930,N_2333);
and U3317 (N_3317,N_1658,N_1046);
or U3318 (N_3318,N_955,N_138);
nor U3319 (N_3319,N_2291,N_1377);
or U3320 (N_3320,N_872,N_367);
nor U3321 (N_3321,N_2336,N_206);
and U3322 (N_3322,N_622,N_1831);
and U3323 (N_3323,N_1745,N_1500);
nor U3324 (N_3324,N_1708,N_750);
nor U3325 (N_3325,N_550,N_725);
nand U3326 (N_3326,N_1075,N_2206);
or U3327 (N_3327,N_1635,N_1467);
nand U3328 (N_3328,N_482,N_938);
and U3329 (N_3329,N_1357,N_2370);
or U3330 (N_3330,N_822,N_1960);
and U3331 (N_3331,N_2314,N_2124);
and U3332 (N_3332,N_1083,N_279);
and U3333 (N_3333,N_40,N_98);
or U3334 (N_3334,N_87,N_1778);
nor U3335 (N_3335,N_335,N_827);
or U3336 (N_3336,N_228,N_34);
and U3337 (N_3337,N_1609,N_355);
or U3338 (N_3338,N_651,N_726);
nor U3339 (N_3339,N_974,N_2105);
nand U3340 (N_3340,N_189,N_1459);
nand U3341 (N_3341,N_123,N_1615);
or U3342 (N_3342,N_407,N_250);
nand U3343 (N_3343,N_1655,N_2160);
nand U3344 (N_3344,N_1981,N_2240);
and U3345 (N_3345,N_1640,N_1622);
or U3346 (N_3346,N_1923,N_1860);
nor U3347 (N_3347,N_662,N_10);
nand U3348 (N_3348,N_2461,N_865);
or U3349 (N_3349,N_2479,N_147);
or U3350 (N_3350,N_488,N_910);
or U3351 (N_3351,N_232,N_1206);
nand U3352 (N_3352,N_2134,N_632);
nor U3353 (N_3353,N_2098,N_1374);
or U3354 (N_3354,N_1811,N_168);
or U3355 (N_3355,N_1666,N_683);
nor U3356 (N_3356,N_2009,N_787);
or U3357 (N_3357,N_526,N_415);
nor U3358 (N_3358,N_2346,N_315);
and U3359 (N_3359,N_867,N_1506);
nor U3360 (N_3360,N_1023,N_580);
nand U3361 (N_3361,N_419,N_2219);
or U3362 (N_3362,N_562,N_1490);
nand U3363 (N_3363,N_216,N_132);
nor U3364 (N_3364,N_1983,N_306);
and U3365 (N_3365,N_1411,N_1203);
nand U3366 (N_3366,N_1036,N_2159);
and U3367 (N_3367,N_1779,N_585);
nor U3368 (N_3368,N_923,N_2481);
and U3369 (N_3369,N_1557,N_983);
nand U3370 (N_3370,N_2447,N_453);
and U3371 (N_3371,N_1474,N_374);
or U3372 (N_3372,N_528,N_383);
nor U3373 (N_3373,N_377,N_1828);
nor U3374 (N_3374,N_114,N_1843);
and U3375 (N_3375,N_2148,N_541);
nand U3376 (N_3376,N_2439,N_1616);
or U3377 (N_3377,N_817,N_1977);
nand U3378 (N_3378,N_2137,N_1070);
nand U3379 (N_3379,N_1626,N_176);
and U3380 (N_3380,N_1287,N_1166);
nand U3381 (N_3381,N_1362,N_1826);
nand U3382 (N_3382,N_596,N_975);
nor U3383 (N_3383,N_1799,N_2045);
or U3384 (N_3384,N_2318,N_1479);
nor U3385 (N_3385,N_1919,N_2188);
and U3386 (N_3386,N_1540,N_917);
nand U3387 (N_3387,N_398,N_1675);
nor U3388 (N_3388,N_603,N_2191);
nor U3389 (N_3389,N_120,N_929);
nor U3390 (N_3390,N_2170,N_1346);
and U3391 (N_3391,N_1239,N_1178);
or U3392 (N_3392,N_2497,N_1692);
and U3393 (N_3393,N_939,N_1962);
nand U3394 (N_3394,N_2491,N_2200);
nand U3395 (N_3395,N_1511,N_1613);
nand U3396 (N_3396,N_2205,N_2350);
and U3397 (N_3397,N_2110,N_41);
nor U3398 (N_3398,N_2357,N_576);
or U3399 (N_3399,N_1442,N_1200);
nand U3400 (N_3400,N_97,N_2343);
or U3401 (N_3401,N_1614,N_1995);
nand U3402 (N_3402,N_157,N_903);
nor U3403 (N_3403,N_2393,N_1716);
or U3404 (N_3404,N_1212,N_1850);
nor U3405 (N_3405,N_1401,N_1883);
or U3406 (N_3406,N_2499,N_185);
or U3407 (N_3407,N_257,N_1891);
and U3408 (N_3408,N_834,N_1403);
nand U3409 (N_3409,N_1308,N_1224);
and U3410 (N_3410,N_564,N_650);
or U3411 (N_3411,N_1430,N_1068);
and U3412 (N_3412,N_1454,N_615);
nor U3413 (N_3413,N_885,N_2256);
or U3414 (N_3414,N_104,N_412);
nand U3415 (N_3415,N_1073,N_375);
nor U3416 (N_3416,N_540,N_235);
and U3417 (N_3417,N_2251,N_1003);
and U3418 (N_3418,N_2027,N_2013);
or U3419 (N_3419,N_523,N_2035);
nand U3420 (N_3420,N_1978,N_2097);
and U3421 (N_3421,N_639,N_1329);
nand U3422 (N_3422,N_2360,N_1296);
nor U3423 (N_3423,N_1971,N_1697);
and U3424 (N_3424,N_2078,N_361);
nand U3425 (N_3425,N_944,N_78);
nand U3426 (N_3426,N_167,N_86);
nand U3427 (N_3427,N_904,N_245);
nor U3428 (N_3428,N_652,N_1834);
nor U3429 (N_3429,N_1699,N_619);
nor U3430 (N_3430,N_371,N_301);
nand U3431 (N_3431,N_1098,N_1687);
and U3432 (N_3432,N_436,N_2484);
nand U3433 (N_3433,N_148,N_837);
and U3434 (N_3434,N_710,N_158);
nand U3435 (N_3435,N_1175,N_2184);
and U3436 (N_3436,N_1194,N_2084);
nand U3437 (N_3437,N_1757,N_2174);
nand U3438 (N_3438,N_1100,N_743);
or U3439 (N_3439,N_2359,N_1974);
or U3440 (N_3440,N_606,N_1136);
nand U3441 (N_3441,N_973,N_661);
nor U3442 (N_3442,N_151,N_57);
nand U3443 (N_3443,N_1216,N_1148);
or U3444 (N_3444,N_2426,N_2490);
nand U3445 (N_3445,N_452,N_824);
and U3446 (N_3446,N_936,N_350);
or U3447 (N_3447,N_2317,N_2248);
or U3448 (N_3448,N_2480,N_1481);
nand U3449 (N_3449,N_2157,N_1356);
nand U3450 (N_3450,N_1412,N_714);
nor U3451 (N_3451,N_480,N_2209);
nand U3452 (N_3452,N_1808,N_349);
nand U3453 (N_3453,N_790,N_16);
nor U3454 (N_3454,N_198,N_1282);
or U3455 (N_3455,N_413,N_1807);
nand U3456 (N_3456,N_2377,N_1436);
nand U3457 (N_3457,N_1235,N_529);
nand U3458 (N_3458,N_1196,N_1365);
or U3459 (N_3459,N_1541,N_2292);
and U3460 (N_3460,N_763,N_1014);
and U3461 (N_3461,N_1450,N_2395);
nand U3462 (N_3462,N_802,N_852);
and U3463 (N_3463,N_89,N_1154);
nand U3464 (N_3464,N_429,N_1517);
nor U3465 (N_3465,N_2411,N_1830);
or U3466 (N_3466,N_2364,N_1956);
nand U3467 (N_3467,N_1116,N_820);
and U3468 (N_3468,N_1208,N_2297);
nor U3469 (N_3469,N_2368,N_998);
and U3470 (N_3470,N_483,N_1520);
nor U3471 (N_3471,N_1948,N_17);
nor U3472 (N_3472,N_518,N_1702);
or U3473 (N_3473,N_1376,N_1926);
nand U3474 (N_3474,N_1039,N_262);
nand U3475 (N_3475,N_2079,N_1092);
nor U3476 (N_3476,N_640,N_1677);
and U3477 (N_3477,N_734,N_609);
nand U3478 (N_3478,N_1966,N_669);
or U3479 (N_3479,N_641,N_1941);
or U3480 (N_3480,N_1535,N_1968);
or U3481 (N_3481,N_568,N_1245);
nand U3482 (N_3482,N_1499,N_1786);
nor U3483 (N_3483,N_2430,N_934);
or U3484 (N_3484,N_363,N_107);
or U3485 (N_3485,N_812,N_1746);
nand U3486 (N_3486,N_1115,N_347);
and U3487 (N_3487,N_1498,N_2004);
or U3488 (N_3488,N_1191,N_1801);
nor U3489 (N_3489,N_44,N_2064);
or U3490 (N_3490,N_2202,N_2241);
nand U3491 (N_3491,N_312,N_2028);
nor U3492 (N_3492,N_256,N_2387);
nor U3493 (N_3493,N_1649,N_490);
or U3494 (N_3494,N_468,N_1588);
nor U3495 (N_3495,N_881,N_1044);
nand U3496 (N_3496,N_351,N_75);
nand U3497 (N_3497,N_2234,N_1169);
nand U3498 (N_3498,N_681,N_65);
nand U3499 (N_3499,N_354,N_1884);
nor U3500 (N_3500,N_590,N_2452);
nand U3501 (N_3501,N_952,N_574);
or U3502 (N_3502,N_712,N_1078);
and U3503 (N_3503,N_701,N_1366);
and U3504 (N_3504,N_331,N_851);
nand U3505 (N_3505,N_8,N_2204);
nor U3506 (N_3506,N_478,N_119);
and U3507 (N_3507,N_1504,N_1187);
nand U3508 (N_3508,N_682,N_908);
nor U3509 (N_3509,N_2261,N_1769);
or U3510 (N_3510,N_1894,N_1643);
nor U3511 (N_3511,N_2498,N_321);
nor U3512 (N_3512,N_161,N_495);
and U3513 (N_3513,N_1907,N_1253);
and U3514 (N_3514,N_287,N_533);
or U3515 (N_3515,N_2001,N_1751);
nor U3516 (N_3516,N_1683,N_788);
and U3517 (N_3517,N_305,N_443);
or U3518 (N_3518,N_511,N_547);
nor U3519 (N_3519,N_922,N_1328);
and U3520 (N_3520,N_878,N_2409);
xnor U3521 (N_3521,N_527,N_1158);
nor U3522 (N_3522,N_1201,N_717);
or U3523 (N_3523,N_2077,N_2308);
or U3524 (N_3524,N_1429,N_667);
and U3525 (N_3525,N_1928,N_1547);
xnor U3526 (N_3526,N_2144,N_753);
or U3527 (N_3527,N_1024,N_333);
nor U3528 (N_3528,N_2422,N_1744);
nand U3529 (N_3529,N_645,N_2247);
nand U3530 (N_3530,N_298,N_60);
nand U3531 (N_3531,N_197,N_1621);
nand U3532 (N_3532,N_1355,N_848);
nand U3533 (N_3533,N_709,N_394);
nand U3534 (N_3534,N_1871,N_587);
nand U3535 (N_3535,N_2353,N_1144);
nand U3536 (N_3536,N_1856,N_1820);
xor U3537 (N_3537,N_379,N_1758);
nor U3538 (N_3538,N_1818,N_1681);
nand U3539 (N_3539,N_736,N_1670);
or U3540 (N_3540,N_2085,N_76);
nor U3541 (N_3541,N_1484,N_678);
or U3542 (N_3542,N_1832,N_1338);
nor U3543 (N_3543,N_143,N_1420);
or U3544 (N_3544,N_384,N_1379);
xnor U3545 (N_3545,N_231,N_965);
nor U3546 (N_3546,N_1026,N_1286);
or U3547 (N_3547,N_508,N_1731);
or U3548 (N_3548,N_2496,N_38);
and U3549 (N_3549,N_1326,N_1492);
and U3550 (N_3550,N_555,N_2451);
or U3551 (N_3551,N_933,N_426);
nor U3552 (N_3552,N_220,N_1656);
or U3553 (N_3553,N_2038,N_1124);
or U3554 (N_3554,N_282,N_2315);
nor U3555 (N_3555,N_942,N_33);
or U3556 (N_3556,N_1503,N_611);
and U3557 (N_3557,N_2265,N_81);
and U3558 (N_3558,N_1625,N_2146);
nand U3559 (N_3559,N_1207,N_1688);
nor U3560 (N_3560,N_2101,N_1849);
and U3561 (N_3561,N_1714,N_798);
and U3562 (N_3562,N_2381,N_2055);
nor U3563 (N_3563,N_1361,N_1103);
or U3564 (N_3564,N_2034,N_129);
nor U3565 (N_3565,N_260,N_2388);
nor U3566 (N_3566,N_434,N_356);
and U3567 (N_3567,N_1259,N_1077);
or U3568 (N_3568,N_1289,N_2183);
nand U3569 (N_3569,N_507,N_627);
and U3570 (N_3570,N_1575,N_1107);
and U3571 (N_3571,N_2161,N_755);
or U3572 (N_3572,N_227,N_578);
nor U3573 (N_3573,N_46,N_1452);
nor U3574 (N_3574,N_222,N_1265);
nor U3575 (N_3575,N_569,N_479);
nor U3576 (N_3576,N_1302,N_1138);
and U3577 (N_3577,N_778,N_1937);
nor U3578 (N_3578,N_1020,N_1132);
or U3579 (N_3579,N_1421,N_940);
or U3580 (N_3580,N_1552,N_772);
and U3581 (N_3581,N_1565,N_1047);
and U3582 (N_3582,N_1564,N_184);
nand U3583 (N_3583,N_992,N_2244);
nand U3584 (N_3584,N_1275,N_455);
nor U3585 (N_3585,N_1497,N_1522);
nand U3586 (N_3586,N_618,N_1327);
and U3587 (N_3587,N_1470,N_1494);
or U3588 (N_3588,N_765,N_1770);
nand U3589 (N_3589,N_1031,N_981);
or U3590 (N_3590,N_1299,N_2145);
or U3591 (N_3591,N_2351,N_1);
nand U3592 (N_3592,N_2424,N_96);
nor U3593 (N_3593,N_1234,N_153);
and U3594 (N_3594,N_926,N_59);
nor U3595 (N_3595,N_2114,N_1006);
nor U3596 (N_3596,N_229,N_1246);
and U3597 (N_3597,N_2123,N_1590);
nor U3598 (N_3598,N_395,N_277);
nand U3599 (N_3599,N_296,N_2024);
nor U3600 (N_3600,N_1397,N_1478);
and U3601 (N_3601,N_139,N_1839);
or U3602 (N_3602,N_464,N_814);
nor U3603 (N_3603,N_1657,N_2466);
nand U3604 (N_3604,N_688,N_1868);
or U3605 (N_3605,N_1563,N_1325);
nor U3606 (N_3606,N_1821,N_1243);
nand U3607 (N_3607,N_91,N_1991);
and U3608 (N_3608,N_62,N_1350);
or U3609 (N_3609,N_329,N_2278);
and U3610 (N_3610,N_175,N_1131);
nor U3611 (N_3611,N_2189,N_1897);
nand U3612 (N_3612,N_201,N_1225);
nor U3613 (N_3613,N_1488,N_1549);
and U3614 (N_3614,N_1872,N_1940);
nor U3615 (N_3615,N_990,N_1333);
and U3616 (N_3616,N_1584,N_2423);
nor U3617 (N_3617,N_193,N_2329);
nor U3618 (N_3618,N_733,N_1431);
or U3619 (N_3619,N_534,N_24);
xor U3620 (N_3620,N_1720,N_597);
and U3621 (N_3621,N_1953,N_1369);
or U3622 (N_3622,N_370,N_159);
and U3623 (N_3623,N_873,N_1840);
and U3624 (N_3624,N_93,N_1781);
nor U3625 (N_3625,N_1344,N_2485);
and U3626 (N_3626,N_1961,N_1487);
nor U3627 (N_3627,N_789,N_2115);
nor U3628 (N_3628,N_1065,N_1809);
xnor U3629 (N_3629,N_638,N_1972);
or U3630 (N_3630,N_225,N_2019);
or U3631 (N_3631,N_520,N_199);
and U3632 (N_3632,N_2017,N_551);
nor U3633 (N_3633,N_1717,N_53);
nor U3634 (N_3634,N_2286,N_1101);
nand U3635 (N_3635,N_2489,N_118);
nor U3636 (N_3636,N_1580,N_127);
and U3637 (N_3637,N_2072,N_1507);
and U3638 (N_3638,N_1074,N_124);
or U3639 (N_3639,N_469,N_486);
nand U3640 (N_3640,N_742,N_2260);
or U3641 (N_3641,N_2092,N_1381);
or U3642 (N_3642,N_748,N_1806);
xor U3643 (N_3643,N_1199,N_2221);
nand U3644 (N_3644,N_913,N_2066);
nand U3645 (N_3645,N_961,N_1110);
nand U3646 (N_3646,N_969,N_2376);
and U3647 (N_3647,N_410,N_1846);
nor U3648 (N_3648,N_2437,N_1320);
or U3649 (N_3649,N_1634,N_1126);
nand U3650 (N_3650,N_2415,N_1301);
and U3651 (N_3651,N_591,N_2075);
or U3652 (N_3652,N_1623,N_727);
or U3653 (N_3653,N_760,N_1337);
xor U3654 (N_3654,N_1653,N_1185);
nor U3655 (N_3655,N_1056,N_2410);
xnor U3656 (N_3656,N_1862,N_203);
nand U3657 (N_3657,N_73,N_403);
nand U3658 (N_3658,N_1217,N_874);
and U3659 (N_3659,N_799,N_268);
and U3660 (N_3660,N_2167,N_1227);
nand U3661 (N_3661,N_1858,N_2014);
and U3662 (N_3662,N_967,N_346);
or U3663 (N_3663,N_1678,N_1996);
and U3664 (N_3664,N_1774,N_1398);
xnor U3665 (N_3665,N_513,N_2469);
and U3666 (N_3666,N_406,N_1571);
nand U3667 (N_3667,N_2060,N_1753);
nand U3668 (N_3668,N_2425,N_876);
nand U3669 (N_3669,N_582,N_832);
and U3670 (N_3670,N_1015,N_1788);
nand U3671 (N_3671,N_2386,N_1710);
nand U3672 (N_3672,N_1909,N_754);
or U3673 (N_3673,N_838,N_18);
nand U3674 (N_3674,N_1578,N_424);
or U3675 (N_3675,N_1546,N_389);
nand U3676 (N_3676,N_1979,N_964);
and U3677 (N_3677,N_1659,N_1309);
nor U3678 (N_3678,N_1603,N_779);
nand U3679 (N_3679,N_472,N_1491);
or U3680 (N_3680,N_1559,N_1917);
and U3681 (N_3681,N_494,N_2112);
and U3682 (N_3682,N_2389,N_126);
or U3683 (N_3683,N_433,N_724);
nor U3684 (N_3684,N_796,N_26);
or U3685 (N_3685,N_769,N_1360);
nor U3686 (N_3686,N_244,N_71);
and U3687 (N_3687,N_1536,N_783);
or U3688 (N_3688,N_11,N_2136);
and U3689 (N_3689,N_1190,N_2220);
nand U3690 (N_3690,N_1726,N_2412);
and U3691 (N_3691,N_1709,N_1533);
nand U3692 (N_3692,N_182,N_2259);
and U3693 (N_3693,N_957,N_1853);
and U3694 (N_3694,N_111,N_2462);
and U3695 (N_3695,N_731,N_2036);
and U3696 (N_3696,N_1924,N_531);
nor U3697 (N_3697,N_2356,N_668);
and U3698 (N_3698,N_2402,N_54);
nand U3699 (N_3699,N_1998,N_160);
or U3700 (N_3700,N_2281,N_1119);
and U3701 (N_3701,N_1548,N_1120);
nor U3702 (N_3702,N_1336,N_1927);
and U3703 (N_3703,N_319,N_708);
or U3704 (N_3704,N_808,N_2284);
nand U3705 (N_3705,N_982,N_1539);
nand U3706 (N_3706,N_140,N_729);
nor U3707 (N_3707,N_996,N_2198);
nor U3708 (N_3708,N_1457,N_275);
and U3709 (N_3709,N_74,N_1364);
and U3710 (N_3710,N_2257,N_566);
and U3711 (N_3711,N_280,N_850);
or U3712 (N_3712,N_1537,N_1880);
or U3713 (N_3713,N_1370,N_187);
nand U3714 (N_3714,N_1627,N_636);
or U3715 (N_3715,N_162,N_448);
nor U3716 (N_3716,N_1051,N_1581);
nand U3717 (N_3717,N_1599,N_1069);
nor U3718 (N_3718,N_309,N_281);
or U3719 (N_3719,N_752,N_807);
and U3720 (N_3720,N_544,N_2132);
or U3721 (N_3721,N_600,N_125);
and U3722 (N_3722,N_1848,N_828);
or U3723 (N_3723,N_366,N_993);
or U3724 (N_3724,N_1495,N_1254);
nor U3725 (N_3725,N_164,N_1791);
nand U3726 (N_3726,N_845,N_629);
nand U3727 (N_3727,N_2021,N_2031);
nand U3728 (N_3728,N_1371,N_2431);
nor U3729 (N_3729,N_1558,N_1901);
and U3730 (N_3730,N_195,N_1134);
nor U3731 (N_3731,N_700,N_2096);
or U3732 (N_3732,N_459,N_801);
or U3733 (N_3733,N_1754,N_1944);
nand U3734 (N_3734,N_1262,N_317);
and U3735 (N_3735,N_237,N_502);
or U3736 (N_3736,N_761,N_2063);
or U3737 (N_3737,N_2041,N_598);
nor U3738 (N_3738,N_1918,N_1569);
nand U3739 (N_3739,N_2338,N_2272);
nor U3740 (N_3740,N_181,N_953);
and U3741 (N_3741,N_1318,N_1608);
nand U3742 (N_3742,N_1637,N_266);
and U3743 (N_3743,N_895,N_1219);
nand U3744 (N_3744,N_1322,N_759);
nand U3745 (N_3745,N_2455,N_2126);
nand U3746 (N_3746,N_699,N_1466);
and U3747 (N_3747,N_935,N_995);
nand U3748 (N_3748,N_1304,N_1335);
nand U3749 (N_3749,N_937,N_1990);
nor U3750 (N_3750,N_470,N_715);
or U3751 (N_3751,N_1217,N_1503);
nor U3752 (N_3752,N_1007,N_2462);
or U3753 (N_3753,N_1341,N_1253);
nand U3754 (N_3754,N_1070,N_1748);
and U3755 (N_3755,N_246,N_206);
and U3756 (N_3756,N_698,N_1554);
nand U3757 (N_3757,N_537,N_2305);
nand U3758 (N_3758,N_28,N_373);
or U3759 (N_3759,N_1916,N_403);
and U3760 (N_3760,N_1260,N_2360);
nand U3761 (N_3761,N_2010,N_570);
nor U3762 (N_3762,N_2098,N_1893);
nor U3763 (N_3763,N_1459,N_2319);
or U3764 (N_3764,N_89,N_2165);
nand U3765 (N_3765,N_2257,N_343);
or U3766 (N_3766,N_684,N_773);
nand U3767 (N_3767,N_996,N_1466);
and U3768 (N_3768,N_434,N_1322);
and U3769 (N_3769,N_2058,N_830);
or U3770 (N_3770,N_931,N_452);
nand U3771 (N_3771,N_925,N_222);
xnor U3772 (N_3772,N_295,N_1623);
xor U3773 (N_3773,N_2450,N_537);
and U3774 (N_3774,N_871,N_934);
nor U3775 (N_3775,N_1998,N_403);
nand U3776 (N_3776,N_390,N_2255);
nor U3777 (N_3777,N_2226,N_1950);
nand U3778 (N_3778,N_2307,N_938);
or U3779 (N_3779,N_890,N_911);
or U3780 (N_3780,N_394,N_2066);
nand U3781 (N_3781,N_2328,N_2383);
nor U3782 (N_3782,N_1977,N_303);
or U3783 (N_3783,N_2413,N_2406);
or U3784 (N_3784,N_1678,N_1526);
or U3785 (N_3785,N_257,N_997);
and U3786 (N_3786,N_1570,N_506);
nor U3787 (N_3787,N_1278,N_159);
xnor U3788 (N_3788,N_16,N_499);
or U3789 (N_3789,N_1989,N_2105);
nor U3790 (N_3790,N_1777,N_1682);
nand U3791 (N_3791,N_1291,N_1769);
nand U3792 (N_3792,N_1853,N_2155);
or U3793 (N_3793,N_727,N_564);
and U3794 (N_3794,N_447,N_2141);
nor U3795 (N_3795,N_2161,N_1078);
and U3796 (N_3796,N_1211,N_792);
nand U3797 (N_3797,N_1617,N_1458);
xor U3798 (N_3798,N_537,N_683);
nand U3799 (N_3799,N_1757,N_381);
or U3800 (N_3800,N_2130,N_61);
nor U3801 (N_3801,N_757,N_1748);
nor U3802 (N_3802,N_192,N_1237);
and U3803 (N_3803,N_1681,N_1366);
nand U3804 (N_3804,N_1030,N_655);
or U3805 (N_3805,N_1968,N_1031);
or U3806 (N_3806,N_1850,N_1295);
or U3807 (N_3807,N_2030,N_1636);
or U3808 (N_3808,N_1146,N_520);
nor U3809 (N_3809,N_182,N_1704);
or U3810 (N_3810,N_1230,N_1895);
or U3811 (N_3811,N_355,N_556);
or U3812 (N_3812,N_2283,N_267);
or U3813 (N_3813,N_2356,N_2011);
or U3814 (N_3814,N_1919,N_2130);
nand U3815 (N_3815,N_316,N_281);
nor U3816 (N_3816,N_1997,N_918);
and U3817 (N_3817,N_1914,N_1809);
or U3818 (N_3818,N_2092,N_478);
nor U3819 (N_3819,N_1208,N_1139);
and U3820 (N_3820,N_635,N_2318);
or U3821 (N_3821,N_2,N_792);
or U3822 (N_3822,N_716,N_1892);
or U3823 (N_3823,N_735,N_1073);
and U3824 (N_3824,N_2344,N_98);
nor U3825 (N_3825,N_739,N_957);
nor U3826 (N_3826,N_244,N_689);
or U3827 (N_3827,N_588,N_741);
or U3828 (N_3828,N_1997,N_2390);
and U3829 (N_3829,N_428,N_1760);
or U3830 (N_3830,N_751,N_1106);
nand U3831 (N_3831,N_1,N_483);
nor U3832 (N_3832,N_362,N_1501);
nor U3833 (N_3833,N_2076,N_2066);
nor U3834 (N_3834,N_1380,N_1749);
nand U3835 (N_3835,N_330,N_169);
or U3836 (N_3836,N_1374,N_1395);
nand U3837 (N_3837,N_2131,N_32);
and U3838 (N_3838,N_650,N_1722);
nand U3839 (N_3839,N_1252,N_4);
and U3840 (N_3840,N_1962,N_838);
nor U3841 (N_3841,N_11,N_963);
or U3842 (N_3842,N_791,N_1307);
and U3843 (N_3843,N_582,N_1823);
or U3844 (N_3844,N_819,N_1679);
and U3845 (N_3845,N_2119,N_157);
nor U3846 (N_3846,N_776,N_595);
or U3847 (N_3847,N_748,N_698);
and U3848 (N_3848,N_2233,N_176);
nand U3849 (N_3849,N_1118,N_2046);
nor U3850 (N_3850,N_976,N_255);
and U3851 (N_3851,N_1070,N_1006);
nand U3852 (N_3852,N_453,N_2302);
or U3853 (N_3853,N_1459,N_940);
nand U3854 (N_3854,N_685,N_733);
nand U3855 (N_3855,N_240,N_1432);
nor U3856 (N_3856,N_1965,N_407);
or U3857 (N_3857,N_152,N_2095);
or U3858 (N_3858,N_1530,N_613);
nand U3859 (N_3859,N_1821,N_2235);
and U3860 (N_3860,N_257,N_887);
and U3861 (N_3861,N_2213,N_845);
or U3862 (N_3862,N_556,N_2155);
and U3863 (N_3863,N_2301,N_1555);
nor U3864 (N_3864,N_529,N_1395);
nand U3865 (N_3865,N_1676,N_1430);
or U3866 (N_3866,N_2110,N_1408);
nand U3867 (N_3867,N_1980,N_2061);
or U3868 (N_3868,N_405,N_1953);
or U3869 (N_3869,N_58,N_1775);
or U3870 (N_3870,N_115,N_413);
or U3871 (N_3871,N_1352,N_2212);
nor U3872 (N_3872,N_86,N_837);
and U3873 (N_3873,N_247,N_320);
and U3874 (N_3874,N_139,N_288);
or U3875 (N_3875,N_2405,N_1069);
nor U3876 (N_3876,N_2362,N_413);
nand U3877 (N_3877,N_1320,N_795);
nor U3878 (N_3878,N_155,N_2459);
nor U3879 (N_3879,N_1472,N_1398);
or U3880 (N_3880,N_1379,N_1365);
or U3881 (N_3881,N_29,N_1748);
and U3882 (N_3882,N_1936,N_1081);
or U3883 (N_3883,N_1343,N_1103);
nand U3884 (N_3884,N_1194,N_2029);
or U3885 (N_3885,N_2160,N_648);
and U3886 (N_3886,N_376,N_1682);
nor U3887 (N_3887,N_543,N_257);
and U3888 (N_3888,N_1238,N_2022);
nor U3889 (N_3889,N_1285,N_346);
and U3890 (N_3890,N_1738,N_1159);
and U3891 (N_3891,N_994,N_843);
nor U3892 (N_3892,N_1228,N_997);
and U3893 (N_3893,N_1890,N_250);
or U3894 (N_3894,N_568,N_22);
nor U3895 (N_3895,N_464,N_1067);
nand U3896 (N_3896,N_1350,N_1290);
nor U3897 (N_3897,N_2078,N_951);
and U3898 (N_3898,N_13,N_847);
nor U3899 (N_3899,N_2258,N_960);
or U3900 (N_3900,N_2415,N_1809);
nor U3901 (N_3901,N_710,N_108);
nand U3902 (N_3902,N_1701,N_16);
or U3903 (N_3903,N_1393,N_1582);
nor U3904 (N_3904,N_1891,N_497);
nor U3905 (N_3905,N_1739,N_1422);
nor U3906 (N_3906,N_70,N_164);
and U3907 (N_3907,N_468,N_973);
or U3908 (N_3908,N_757,N_1320);
or U3909 (N_3909,N_150,N_2413);
nor U3910 (N_3910,N_59,N_1943);
and U3911 (N_3911,N_1015,N_522);
nor U3912 (N_3912,N_1449,N_1989);
and U3913 (N_3913,N_1043,N_2249);
nor U3914 (N_3914,N_570,N_520);
or U3915 (N_3915,N_1653,N_680);
or U3916 (N_3916,N_962,N_2184);
nor U3917 (N_3917,N_1125,N_1728);
nand U3918 (N_3918,N_1393,N_2204);
nor U3919 (N_3919,N_714,N_1113);
nor U3920 (N_3920,N_1146,N_1836);
and U3921 (N_3921,N_1758,N_1357);
or U3922 (N_3922,N_1109,N_396);
nor U3923 (N_3923,N_2496,N_760);
nand U3924 (N_3924,N_1316,N_1955);
nand U3925 (N_3925,N_2467,N_730);
or U3926 (N_3926,N_365,N_881);
nand U3927 (N_3927,N_2360,N_2127);
nor U3928 (N_3928,N_2485,N_1182);
nor U3929 (N_3929,N_1774,N_160);
and U3930 (N_3930,N_1302,N_996);
nor U3931 (N_3931,N_2173,N_981);
and U3932 (N_3932,N_1216,N_1054);
or U3933 (N_3933,N_1180,N_1233);
or U3934 (N_3934,N_1766,N_1509);
nand U3935 (N_3935,N_719,N_2218);
nor U3936 (N_3936,N_618,N_525);
nor U3937 (N_3937,N_877,N_1078);
nand U3938 (N_3938,N_2418,N_2016);
nor U3939 (N_3939,N_374,N_1132);
nand U3940 (N_3940,N_2277,N_2477);
nor U3941 (N_3941,N_978,N_1401);
nand U3942 (N_3942,N_2361,N_1583);
and U3943 (N_3943,N_1946,N_2266);
nor U3944 (N_3944,N_1858,N_1834);
or U3945 (N_3945,N_53,N_1543);
nor U3946 (N_3946,N_1471,N_592);
nor U3947 (N_3947,N_491,N_950);
nor U3948 (N_3948,N_860,N_95);
nor U3949 (N_3949,N_2180,N_2425);
nor U3950 (N_3950,N_366,N_1726);
nand U3951 (N_3951,N_617,N_1744);
nor U3952 (N_3952,N_701,N_1060);
and U3953 (N_3953,N_1711,N_1599);
and U3954 (N_3954,N_1406,N_912);
or U3955 (N_3955,N_1366,N_2275);
nand U3956 (N_3956,N_1805,N_2332);
and U3957 (N_3957,N_2116,N_173);
and U3958 (N_3958,N_2256,N_1709);
or U3959 (N_3959,N_755,N_2306);
nand U3960 (N_3960,N_838,N_1032);
and U3961 (N_3961,N_1645,N_1731);
and U3962 (N_3962,N_776,N_1013);
and U3963 (N_3963,N_267,N_2420);
and U3964 (N_3964,N_259,N_541);
or U3965 (N_3965,N_1674,N_1200);
nor U3966 (N_3966,N_50,N_1514);
nor U3967 (N_3967,N_1279,N_2185);
nand U3968 (N_3968,N_509,N_448);
xnor U3969 (N_3969,N_1571,N_749);
and U3970 (N_3970,N_2035,N_1152);
or U3971 (N_3971,N_1726,N_1926);
or U3972 (N_3972,N_1096,N_130);
nor U3973 (N_3973,N_1014,N_675);
and U3974 (N_3974,N_673,N_1953);
or U3975 (N_3975,N_1004,N_2413);
and U3976 (N_3976,N_22,N_1299);
nor U3977 (N_3977,N_2326,N_1347);
and U3978 (N_3978,N_1569,N_1033);
and U3979 (N_3979,N_600,N_1465);
or U3980 (N_3980,N_1560,N_1314);
and U3981 (N_3981,N_1046,N_2241);
nor U3982 (N_3982,N_2411,N_2207);
and U3983 (N_3983,N_373,N_53);
and U3984 (N_3984,N_2127,N_1407);
or U3985 (N_3985,N_126,N_730);
nor U3986 (N_3986,N_1135,N_1442);
nand U3987 (N_3987,N_608,N_1361);
nor U3988 (N_3988,N_919,N_2070);
xor U3989 (N_3989,N_1155,N_544);
and U3990 (N_3990,N_1030,N_1867);
xnor U3991 (N_3991,N_1316,N_896);
nand U3992 (N_3992,N_2209,N_1391);
nand U3993 (N_3993,N_1548,N_2128);
nand U3994 (N_3994,N_2103,N_722);
and U3995 (N_3995,N_914,N_2498);
nand U3996 (N_3996,N_1653,N_1200);
nand U3997 (N_3997,N_1215,N_855);
or U3998 (N_3998,N_2463,N_771);
nand U3999 (N_3999,N_1458,N_1031);
and U4000 (N_4000,N_1511,N_235);
nor U4001 (N_4001,N_1988,N_2489);
nand U4002 (N_4002,N_124,N_9);
nor U4003 (N_4003,N_1751,N_1580);
and U4004 (N_4004,N_1589,N_2275);
nor U4005 (N_4005,N_1794,N_2342);
or U4006 (N_4006,N_2161,N_455);
nor U4007 (N_4007,N_788,N_993);
nand U4008 (N_4008,N_477,N_2010);
nand U4009 (N_4009,N_1766,N_1976);
or U4010 (N_4010,N_4,N_641);
and U4011 (N_4011,N_2311,N_572);
and U4012 (N_4012,N_975,N_747);
or U4013 (N_4013,N_1971,N_1876);
nand U4014 (N_4014,N_564,N_2020);
nand U4015 (N_4015,N_957,N_1168);
nand U4016 (N_4016,N_1340,N_2114);
xor U4017 (N_4017,N_2038,N_2332);
or U4018 (N_4018,N_1534,N_1323);
or U4019 (N_4019,N_1458,N_2238);
and U4020 (N_4020,N_1710,N_1143);
and U4021 (N_4021,N_2345,N_2337);
and U4022 (N_4022,N_2457,N_1241);
nor U4023 (N_4023,N_2315,N_1323);
nor U4024 (N_4024,N_1952,N_1512);
and U4025 (N_4025,N_367,N_1623);
nand U4026 (N_4026,N_2079,N_1417);
nand U4027 (N_4027,N_1279,N_1701);
nand U4028 (N_4028,N_196,N_738);
and U4029 (N_4029,N_656,N_884);
or U4030 (N_4030,N_1881,N_680);
and U4031 (N_4031,N_2463,N_1001);
and U4032 (N_4032,N_120,N_604);
and U4033 (N_4033,N_83,N_1273);
and U4034 (N_4034,N_1190,N_337);
or U4035 (N_4035,N_81,N_2499);
or U4036 (N_4036,N_1514,N_2355);
or U4037 (N_4037,N_2133,N_266);
or U4038 (N_4038,N_1731,N_2129);
and U4039 (N_4039,N_1885,N_179);
or U4040 (N_4040,N_2384,N_1319);
and U4041 (N_4041,N_1254,N_2497);
and U4042 (N_4042,N_1961,N_1533);
nor U4043 (N_4043,N_1941,N_2454);
nor U4044 (N_4044,N_852,N_2333);
nand U4045 (N_4045,N_1031,N_694);
nand U4046 (N_4046,N_170,N_1442);
nor U4047 (N_4047,N_1505,N_2049);
or U4048 (N_4048,N_1049,N_1633);
or U4049 (N_4049,N_1082,N_645);
nand U4050 (N_4050,N_2420,N_175);
and U4051 (N_4051,N_747,N_1780);
or U4052 (N_4052,N_412,N_2470);
and U4053 (N_4053,N_2065,N_1311);
or U4054 (N_4054,N_2347,N_239);
or U4055 (N_4055,N_1638,N_1799);
and U4056 (N_4056,N_1871,N_262);
nor U4057 (N_4057,N_2057,N_622);
nor U4058 (N_4058,N_53,N_959);
nand U4059 (N_4059,N_1558,N_2057);
or U4060 (N_4060,N_1379,N_1226);
nand U4061 (N_4061,N_1702,N_1283);
nor U4062 (N_4062,N_2328,N_1249);
and U4063 (N_4063,N_1877,N_1258);
and U4064 (N_4064,N_620,N_806);
nor U4065 (N_4065,N_2305,N_1836);
or U4066 (N_4066,N_1131,N_491);
and U4067 (N_4067,N_1008,N_10);
nand U4068 (N_4068,N_40,N_1263);
nand U4069 (N_4069,N_382,N_2140);
nand U4070 (N_4070,N_1165,N_1135);
and U4071 (N_4071,N_697,N_539);
nand U4072 (N_4072,N_1360,N_1384);
nor U4073 (N_4073,N_875,N_541);
and U4074 (N_4074,N_1415,N_1617);
and U4075 (N_4075,N_2107,N_334);
nand U4076 (N_4076,N_1891,N_1204);
nand U4077 (N_4077,N_617,N_1547);
nor U4078 (N_4078,N_680,N_902);
nor U4079 (N_4079,N_1409,N_1871);
and U4080 (N_4080,N_1830,N_1548);
or U4081 (N_4081,N_2345,N_2313);
or U4082 (N_4082,N_2266,N_2076);
nand U4083 (N_4083,N_1873,N_1400);
nor U4084 (N_4084,N_2090,N_2099);
nor U4085 (N_4085,N_51,N_1545);
and U4086 (N_4086,N_1010,N_1258);
and U4087 (N_4087,N_1470,N_1793);
or U4088 (N_4088,N_32,N_2184);
nor U4089 (N_4089,N_1445,N_264);
or U4090 (N_4090,N_1632,N_1782);
nand U4091 (N_4091,N_1879,N_1995);
nand U4092 (N_4092,N_342,N_587);
and U4093 (N_4093,N_1182,N_2128);
nand U4094 (N_4094,N_1467,N_1915);
and U4095 (N_4095,N_1866,N_710);
or U4096 (N_4096,N_1841,N_2021);
and U4097 (N_4097,N_1894,N_1688);
or U4098 (N_4098,N_2318,N_1190);
and U4099 (N_4099,N_263,N_11);
or U4100 (N_4100,N_764,N_1503);
nand U4101 (N_4101,N_2291,N_1853);
or U4102 (N_4102,N_804,N_2063);
or U4103 (N_4103,N_112,N_2046);
or U4104 (N_4104,N_2415,N_857);
and U4105 (N_4105,N_446,N_1966);
and U4106 (N_4106,N_263,N_2382);
nor U4107 (N_4107,N_2049,N_1105);
and U4108 (N_4108,N_163,N_1744);
or U4109 (N_4109,N_1960,N_580);
nand U4110 (N_4110,N_2103,N_2305);
nor U4111 (N_4111,N_574,N_1076);
nor U4112 (N_4112,N_899,N_2052);
nor U4113 (N_4113,N_373,N_2449);
nand U4114 (N_4114,N_1631,N_1294);
or U4115 (N_4115,N_1405,N_2186);
nand U4116 (N_4116,N_86,N_379);
nand U4117 (N_4117,N_206,N_81);
nor U4118 (N_4118,N_1783,N_2439);
nand U4119 (N_4119,N_653,N_305);
nand U4120 (N_4120,N_2486,N_377);
and U4121 (N_4121,N_1013,N_1712);
nor U4122 (N_4122,N_1226,N_601);
and U4123 (N_4123,N_256,N_146);
nand U4124 (N_4124,N_648,N_1684);
and U4125 (N_4125,N_957,N_2364);
and U4126 (N_4126,N_678,N_1598);
and U4127 (N_4127,N_2498,N_305);
nand U4128 (N_4128,N_1223,N_1885);
xnor U4129 (N_4129,N_1560,N_1987);
or U4130 (N_4130,N_1621,N_2054);
or U4131 (N_4131,N_763,N_1593);
or U4132 (N_4132,N_226,N_904);
and U4133 (N_4133,N_1793,N_49);
nor U4134 (N_4134,N_1489,N_736);
nor U4135 (N_4135,N_2252,N_469);
nor U4136 (N_4136,N_1056,N_1136);
and U4137 (N_4137,N_817,N_1579);
and U4138 (N_4138,N_12,N_463);
nor U4139 (N_4139,N_1422,N_891);
and U4140 (N_4140,N_21,N_1362);
or U4141 (N_4141,N_2021,N_1971);
nor U4142 (N_4142,N_1065,N_2254);
or U4143 (N_4143,N_69,N_1783);
nor U4144 (N_4144,N_1418,N_2181);
nor U4145 (N_4145,N_2450,N_1701);
nor U4146 (N_4146,N_1737,N_349);
nor U4147 (N_4147,N_2488,N_772);
and U4148 (N_4148,N_647,N_2453);
or U4149 (N_4149,N_2204,N_1033);
nand U4150 (N_4150,N_377,N_286);
nand U4151 (N_4151,N_657,N_832);
or U4152 (N_4152,N_2467,N_1336);
or U4153 (N_4153,N_1007,N_2471);
nor U4154 (N_4154,N_793,N_2446);
or U4155 (N_4155,N_757,N_1596);
nand U4156 (N_4156,N_684,N_1507);
nand U4157 (N_4157,N_588,N_1049);
or U4158 (N_4158,N_203,N_1036);
or U4159 (N_4159,N_1933,N_1200);
nor U4160 (N_4160,N_11,N_1098);
and U4161 (N_4161,N_1867,N_1157);
nand U4162 (N_4162,N_2238,N_1695);
nand U4163 (N_4163,N_740,N_796);
nand U4164 (N_4164,N_2121,N_2309);
or U4165 (N_4165,N_2047,N_2093);
or U4166 (N_4166,N_21,N_2280);
or U4167 (N_4167,N_23,N_1599);
nor U4168 (N_4168,N_905,N_569);
and U4169 (N_4169,N_609,N_1148);
xnor U4170 (N_4170,N_1003,N_485);
and U4171 (N_4171,N_1038,N_118);
or U4172 (N_4172,N_2280,N_1510);
nor U4173 (N_4173,N_1787,N_929);
or U4174 (N_4174,N_2492,N_1938);
and U4175 (N_4175,N_246,N_1407);
or U4176 (N_4176,N_559,N_2047);
or U4177 (N_4177,N_1761,N_1953);
nand U4178 (N_4178,N_1739,N_2075);
and U4179 (N_4179,N_2363,N_2310);
nand U4180 (N_4180,N_2141,N_293);
or U4181 (N_4181,N_2355,N_505);
or U4182 (N_4182,N_1846,N_1091);
nor U4183 (N_4183,N_137,N_112);
or U4184 (N_4184,N_968,N_563);
or U4185 (N_4185,N_370,N_1932);
nand U4186 (N_4186,N_2238,N_1482);
or U4187 (N_4187,N_885,N_1978);
xnor U4188 (N_4188,N_2270,N_960);
nor U4189 (N_4189,N_1060,N_559);
nand U4190 (N_4190,N_2248,N_356);
and U4191 (N_4191,N_1927,N_1857);
or U4192 (N_4192,N_2166,N_2469);
nor U4193 (N_4193,N_1071,N_1894);
nand U4194 (N_4194,N_1963,N_789);
or U4195 (N_4195,N_1080,N_2063);
or U4196 (N_4196,N_521,N_870);
nor U4197 (N_4197,N_1003,N_883);
or U4198 (N_4198,N_713,N_1542);
nor U4199 (N_4199,N_1598,N_1467);
and U4200 (N_4200,N_171,N_2080);
nand U4201 (N_4201,N_100,N_577);
nand U4202 (N_4202,N_2293,N_1321);
or U4203 (N_4203,N_239,N_1356);
nand U4204 (N_4204,N_1003,N_1976);
nand U4205 (N_4205,N_972,N_1187);
or U4206 (N_4206,N_414,N_2330);
or U4207 (N_4207,N_1775,N_1803);
or U4208 (N_4208,N_173,N_1418);
and U4209 (N_4209,N_1038,N_1186);
and U4210 (N_4210,N_920,N_1659);
nor U4211 (N_4211,N_1888,N_624);
nor U4212 (N_4212,N_1394,N_840);
and U4213 (N_4213,N_1852,N_501);
nand U4214 (N_4214,N_1185,N_1711);
or U4215 (N_4215,N_2293,N_2173);
nand U4216 (N_4216,N_7,N_2295);
and U4217 (N_4217,N_77,N_1782);
or U4218 (N_4218,N_1798,N_1551);
and U4219 (N_4219,N_740,N_1828);
or U4220 (N_4220,N_1261,N_1490);
and U4221 (N_4221,N_1777,N_2439);
or U4222 (N_4222,N_2027,N_212);
nand U4223 (N_4223,N_2470,N_2084);
nor U4224 (N_4224,N_1285,N_33);
nor U4225 (N_4225,N_2267,N_2185);
or U4226 (N_4226,N_1749,N_1647);
nor U4227 (N_4227,N_881,N_1213);
and U4228 (N_4228,N_559,N_229);
nand U4229 (N_4229,N_717,N_488);
nor U4230 (N_4230,N_1572,N_182);
nand U4231 (N_4231,N_1906,N_2319);
or U4232 (N_4232,N_759,N_1439);
and U4233 (N_4233,N_1633,N_1610);
or U4234 (N_4234,N_179,N_838);
or U4235 (N_4235,N_1579,N_2042);
nor U4236 (N_4236,N_694,N_850);
and U4237 (N_4237,N_382,N_1639);
or U4238 (N_4238,N_1880,N_966);
nor U4239 (N_4239,N_630,N_366);
and U4240 (N_4240,N_100,N_2142);
nand U4241 (N_4241,N_925,N_1456);
nor U4242 (N_4242,N_2069,N_2282);
and U4243 (N_4243,N_1784,N_550);
nand U4244 (N_4244,N_678,N_2030);
nand U4245 (N_4245,N_883,N_2335);
and U4246 (N_4246,N_719,N_2476);
nor U4247 (N_4247,N_209,N_1181);
nand U4248 (N_4248,N_2128,N_2401);
nand U4249 (N_4249,N_1218,N_617);
nor U4250 (N_4250,N_511,N_611);
nor U4251 (N_4251,N_125,N_2328);
and U4252 (N_4252,N_1543,N_689);
and U4253 (N_4253,N_2382,N_1212);
nand U4254 (N_4254,N_1529,N_1192);
and U4255 (N_4255,N_1009,N_1367);
and U4256 (N_4256,N_1573,N_269);
nor U4257 (N_4257,N_1511,N_2364);
or U4258 (N_4258,N_705,N_1605);
nand U4259 (N_4259,N_84,N_1714);
and U4260 (N_4260,N_362,N_1439);
nor U4261 (N_4261,N_783,N_1521);
nand U4262 (N_4262,N_2149,N_1764);
or U4263 (N_4263,N_1248,N_878);
and U4264 (N_4264,N_1036,N_762);
and U4265 (N_4265,N_1022,N_2214);
nand U4266 (N_4266,N_2461,N_1519);
nor U4267 (N_4267,N_1002,N_1393);
and U4268 (N_4268,N_443,N_855);
nand U4269 (N_4269,N_572,N_615);
nand U4270 (N_4270,N_965,N_1999);
xor U4271 (N_4271,N_2468,N_611);
or U4272 (N_4272,N_151,N_378);
or U4273 (N_4273,N_823,N_1734);
nor U4274 (N_4274,N_995,N_1699);
or U4275 (N_4275,N_2191,N_1041);
or U4276 (N_4276,N_907,N_1493);
or U4277 (N_4277,N_1951,N_279);
and U4278 (N_4278,N_1693,N_2065);
and U4279 (N_4279,N_19,N_440);
or U4280 (N_4280,N_753,N_2120);
and U4281 (N_4281,N_2018,N_1208);
and U4282 (N_4282,N_1830,N_580);
and U4283 (N_4283,N_975,N_1218);
or U4284 (N_4284,N_257,N_542);
or U4285 (N_4285,N_1807,N_1117);
and U4286 (N_4286,N_2082,N_1267);
and U4287 (N_4287,N_2218,N_1911);
and U4288 (N_4288,N_806,N_1302);
or U4289 (N_4289,N_1766,N_1333);
or U4290 (N_4290,N_159,N_2482);
and U4291 (N_4291,N_2173,N_142);
nor U4292 (N_4292,N_2400,N_70);
or U4293 (N_4293,N_953,N_1857);
nor U4294 (N_4294,N_2244,N_2110);
nand U4295 (N_4295,N_1401,N_506);
nand U4296 (N_4296,N_2250,N_1091);
or U4297 (N_4297,N_1200,N_325);
and U4298 (N_4298,N_48,N_685);
or U4299 (N_4299,N_2013,N_678);
and U4300 (N_4300,N_790,N_881);
nand U4301 (N_4301,N_777,N_468);
nand U4302 (N_4302,N_291,N_68);
and U4303 (N_4303,N_1561,N_1088);
or U4304 (N_4304,N_2073,N_2484);
and U4305 (N_4305,N_1270,N_357);
or U4306 (N_4306,N_630,N_324);
or U4307 (N_4307,N_1216,N_228);
or U4308 (N_4308,N_467,N_1131);
nor U4309 (N_4309,N_842,N_964);
and U4310 (N_4310,N_1630,N_1277);
nor U4311 (N_4311,N_775,N_733);
or U4312 (N_4312,N_574,N_1343);
nor U4313 (N_4313,N_1333,N_827);
nor U4314 (N_4314,N_458,N_1150);
and U4315 (N_4315,N_1781,N_470);
nor U4316 (N_4316,N_2112,N_1772);
nand U4317 (N_4317,N_450,N_1014);
nor U4318 (N_4318,N_2409,N_1176);
nand U4319 (N_4319,N_511,N_723);
or U4320 (N_4320,N_386,N_855);
nand U4321 (N_4321,N_202,N_1896);
and U4322 (N_4322,N_568,N_1570);
nand U4323 (N_4323,N_1907,N_171);
nor U4324 (N_4324,N_282,N_534);
nor U4325 (N_4325,N_475,N_1330);
and U4326 (N_4326,N_1485,N_1371);
nor U4327 (N_4327,N_1508,N_2255);
or U4328 (N_4328,N_2470,N_355);
or U4329 (N_4329,N_1542,N_2080);
or U4330 (N_4330,N_1415,N_289);
nor U4331 (N_4331,N_1331,N_2089);
or U4332 (N_4332,N_1702,N_511);
and U4333 (N_4333,N_942,N_2116);
and U4334 (N_4334,N_271,N_1547);
and U4335 (N_4335,N_598,N_1566);
nor U4336 (N_4336,N_5,N_736);
nand U4337 (N_4337,N_395,N_2190);
nor U4338 (N_4338,N_77,N_1156);
or U4339 (N_4339,N_1495,N_1566);
or U4340 (N_4340,N_1763,N_2197);
and U4341 (N_4341,N_2498,N_1953);
or U4342 (N_4342,N_474,N_71);
and U4343 (N_4343,N_29,N_648);
or U4344 (N_4344,N_1066,N_1413);
nand U4345 (N_4345,N_2259,N_1758);
or U4346 (N_4346,N_1754,N_1530);
and U4347 (N_4347,N_1321,N_2488);
nand U4348 (N_4348,N_281,N_1953);
nor U4349 (N_4349,N_2066,N_2455);
and U4350 (N_4350,N_1524,N_563);
and U4351 (N_4351,N_415,N_660);
nand U4352 (N_4352,N_1339,N_1870);
nor U4353 (N_4353,N_1062,N_2078);
nor U4354 (N_4354,N_1378,N_695);
and U4355 (N_4355,N_1689,N_2465);
nor U4356 (N_4356,N_237,N_1605);
nand U4357 (N_4357,N_2059,N_604);
and U4358 (N_4358,N_287,N_458);
or U4359 (N_4359,N_1973,N_2199);
and U4360 (N_4360,N_1868,N_965);
nor U4361 (N_4361,N_135,N_1877);
or U4362 (N_4362,N_1696,N_2351);
nor U4363 (N_4363,N_2139,N_1899);
and U4364 (N_4364,N_424,N_1469);
and U4365 (N_4365,N_2103,N_795);
nand U4366 (N_4366,N_2134,N_2047);
and U4367 (N_4367,N_1717,N_2374);
nand U4368 (N_4368,N_894,N_792);
and U4369 (N_4369,N_2388,N_1770);
nand U4370 (N_4370,N_134,N_22);
nor U4371 (N_4371,N_1718,N_407);
nor U4372 (N_4372,N_1443,N_1790);
and U4373 (N_4373,N_371,N_2043);
nor U4374 (N_4374,N_1323,N_1199);
nor U4375 (N_4375,N_2006,N_947);
nor U4376 (N_4376,N_2463,N_2420);
and U4377 (N_4377,N_1510,N_148);
or U4378 (N_4378,N_1631,N_78);
and U4379 (N_4379,N_1369,N_1756);
nand U4380 (N_4380,N_1095,N_843);
and U4381 (N_4381,N_1920,N_477);
and U4382 (N_4382,N_1967,N_547);
or U4383 (N_4383,N_748,N_1639);
and U4384 (N_4384,N_1423,N_1477);
nor U4385 (N_4385,N_626,N_1373);
or U4386 (N_4386,N_2377,N_954);
and U4387 (N_4387,N_490,N_515);
nand U4388 (N_4388,N_1584,N_1734);
or U4389 (N_4389,N_2280,N_1101);
and U4390 (N_4390,N_1047,N_650);
or U4391 (N_4391,N_1228,N_2297);
and U4392 (N_4392,N_2409,N_2492);
nor U4393 (N_4393,N_495,N_1243);
or U4394 (N_4394,N_1574,N_2181);
nand U4395 (N_4395,N_1721,N_1745);
nand U4396 (N_4396,N_1331,N_440);
or U4397 (N_4397,N_1937,N_611);
nor U4398 (N_4398,N_1612,N_1289);
nand U4399 (N_4399,N_2051,N_2163);
nor U4400 (N_4400,N_2067,N_560);
and U4401 (N_4401,N_1947,N_1065);
or U4402 (N_4402,N_1736,N_5);
nor U4403 (N_4403,N_431,N_561);
nor U4404 (N_4404,N_2277,N_949);
and U4405 (N_4405,N_878,N_1296);
or U4406 (N_4406,N_1144,N_558);
xor U4407 (N_4407,N_1509,N_2000);
xor U4408 (N_4408,N_876,N_289);
and U4409 (N_4409,N_1290,N_2330);
and U4410 (N_4410,N_75,N_1689);
and U4411 (N_4411,N_1198,N_261);
nand U4412 (N_4412,N_1584,N_787);
or U4413 (N_4413,N_918,N_2233);
and U4414 (N_4414,N_608,N_874);
or U4415 (N_4415,N_354,N_143);
nor U4416 (N_4416,N_1917,N_1350);
or U4417 (N_4417,N_55,N_364);
nand U4418 (N_4418,N_676,N_426);
nand U4419 (N_4419,N_1543,N_541);
nand U4420 (N_4420,N_1348,N_249);
and U4421 (N_4421,N_801,N_772);
nand U4422 (N_4422,N_1474,N_493);
nand U4423 (N_4423,N_1315,N_297);
nand U4424 (N_4424,N_996,N_903);
and U4425 (N_4425,N_92,N_1172);
and U4426 (N_4426,N_934,N_478);
or U4427 (N_4427,N_2085,N_1738);
nand U4428 (N_4428,N_459,N_1455);
nor U4429 (N_4429,N_638,N_1382);
and U4430 (N_4430,N_391,N_2076);
nor U4431 (N_4431,N_1952,N_725);
or U4432 (N_4432,N_1592,N_1647);
nand U4433 (N_4433,N_727,N_2287);
or U4434 (N_4434,N_1169,N_2277);
and U4435 (N_4435,N_1428,N_2172);
and U4436 (N_4436,N_224,N_1389);
nor U4437 (N_4437,N_308,N_1538);
or U4438 (N_4438,N_1739,N_1367);
and U4439 (N_4439,N_973,N_696);
nor U4440 (N_4440,N_809,N_2044);
or U4441 (N_4441,N_464,N_375);
nand U4442 (N_4442,N_461,N_2249);
nand U4443 (N_4443,N_1700,N_1011);
nor U4444 (N_4444,N_789,N_99);
nor U4445 (N_4445,N_18,N_1613);
nor U4446 (N_4446,N_1998,N_2033);
nand U4447 (N_4447,N_971,N_2162);
nor U4448 (N_4448,N_1084,N_298);
or U4449 (N_4449,N_1355,N_1122);
nor U4450 (N_4450,N_2361,N_482);
nor U4451 (N_4451,N_2472,N_777);
nand U4452 (N_4452,N_593,N_2321);
nand U4453 (N_4453,N_1401,N_1730);
and U4454 (N_4454,N_1820,N_119);
nand U4455 (N_4455,N_2018,N_915);
nor U4456 (N_4456,N_2271,N_1850);
and U4457 (N_4457,N_1681,N_1407);
nor U4458 (N_4458,N_1728,N_1454);
or U4459 (N_4459,N_734,N_67);
or U4460 (N_4460,N_263,N_2152);
and U4461 (N_4461,N_18,N_1324);
nand U4462 (N_4462,N_2399,N_0);
or U4463 (N_4463,N_1422,N_1600);
nor U4464 (N_4464,N_866,N_1684);
or U4465 (N_4465,N_1262,N_2359);
nand U4466 (N_4466,N_1719,N_98);
nor U4467 (N_4467,N_228,N_14);
nor U4468 (N_4468,N_1427,N_1838);
nand U4469 (N_4469,N_1659,N_2449);
and U4470 (N_4470,N_332,N_51);
or U4471 (N_4471,N_1068,N_1907);
nand U4472 (N_4472,N_2064,N_1446);
or U4473 (N_4473,N_2261,N_207);
nand U4474 (N_4474,N_281,N_235);
and U4475 (N_4475,N_2036,N_1855);
nand U4476 (N_4476,N_1478,N_1917);
and U4477 (N_4477,N_244,N_77);
nor U4478 (N_4478,N_2093,N_791);
nand U4479 (N_4479,N_1708,N_170);
nand U4480 (N_4480,N_1911,N_2224);
nor U4481 (N_4481,N_1430,N_2310);
nand U4482 (N_4482,N_2396,N_463);
or U4483 (N_4483,N_871,N_2245);
or U4484 (N_4484,N_714,N_2260);
or U4485 (N_4485,N_259,N_141);
or U4486 (N_4486,N_1767,N_1488);
and U4487 (N_4487,N_997,N_579);
nand U4488 (N_4488,N_60,N_279);
nor U4489 (N_4489,N_419,N_1759);
nand U4490 (N_4490,N_665,N_142);
or U4491 (N_4491,N_332,N_2250);
and U4492 (N_4492,N_484,N_744);
or U4493 (N_4493,N_2361,N_1559);
and U4494 (N_4494,N_148,N_1969);
or U4495 (N_4495,N_830,N_430);
or U4496 (N_4496,N_1168,N_1284);
and U4497 (N_4497,N_1108,N_1284);
and U4498 (N_4498,N_1033,N_2354);
nor U4499 (N_4499,N_612,N_945);
or U4500 (N_4500,N_631,N_753);
or U4501 (N_4501,N_1968,N_2178);
nand U4502 (N_4502,N_1840,N_1077);
nand U4503 (N_4503,N_247,N_1226);
nand U4504 (N_4504,N_1288,N_650);
nand U4505 (N_4505,N_2019,N_55);
nor U4506 (N_4506,N_1561,N_1029);
and U4507 (N_4507,N_939,N_187);
nand U4508 (N_4508,N_357,N_298);
and U4509 (N_4509,N_554,N_1698);
or U4510 (N_4510,N_1913,N_194);
or U4511 (N_4511,N_2448,N_712);
and U4512 (N_4512,N_2340,N_1844);
or U4513 (N_4513,N_193,N_1547);
nor U4514 (N_4514,N_1221,N_1060);
and U4515 (N_4515,N_2273,N_43);
nand U4516 (N_4516,N_929,N_320);
nor U4517 (N_4517,N_1577,N_1289);
nor U4518 (N_4518,N_2263,N_1148);
nand U4519 (N_4519,N_1019,N_2112);
and U4520 (N_4520,N_838,N_2205);
nand U4521 (N_4521,N_1072,N_1573);
nand U4522 (N_4522,N_2324,N_157);
nor U4523 (N_4523,N_990,N_514);
and U4524 (N_4524,N_108,N_411);
and U4525 (N_4525,N_2332,N_401);
or U4526 (N_4526,N_1766,N_1245);
nand U4527 (N_4527,N_20,N_1384);
or U4528 (N_4528,N_2467,N_1354);
nand U4529 (N_4529,N_1584,N_2448);
nor U4530 (N_4530,N_1253,N_26);
and U4531 (N_4531,N_495,N_837);
nand U4532 (N_4532,N_2185,N_308);
or U4533 (N_4533,N_270,N_906);
nor U4534 (N_4534,N_378,N_1911);
xor U4535 (N_4535,N_1203,N_2432);
nor U4536 (N_4536,N_2027,N_840);
nand U4537 (N_4537,N_1826,N_1018);
nor U4538 (N_4538,N_269,N_293);
and U4539 (N_4539,N_837,N_876);
nand U4540 (N_4540,N_1891,N_1916);
and U4541 (N_4541,N_630,N_660);
nor U4542 (N_4542,N_99,N_2107);
and U4543 (N_4543,N_1713,N_2415);
xor U4544 (N_4544,N_2480,N_2261);
nand U4545 (N_4545,N_1375,N_2409);
and U4546 (N_4546,N_1537,N_1947);
and U4547 (N_4547,N_114,N_864);
nand U4548 (N_4548,N_172,N_358);
or U4549 (N_4549,N_659,N_522);
or U4550 (N_4550,N_1088,N_688);
nor U4551 (N_4551,N_1415,N_967);
nor U4552 (N_4552,N_1056,N_1519);
and U4553 (N_4553,N_1081,N_2343);
nor U4554 (N_4554,N_2134,N_29);
or U4555 (N_4555,N_1560,N_1501);
and U4556 (N_4556,N_46,N_2275);
nor U4557 (N_4557,N_325,N_7);
or U4558 (N_4558,N_770,N_1620);
and U4559 (N_4559,N_1417,N_1041);
or U4560 (N_4560,N_1619,N_1857);
nand U4561 (N_4561,N_1,N_1120);
nor U4562 (N_4562,N_537,N_2221);
and U4563 (N_4563,N_670,N_1616);
nand U4564 (N_4564,N_2173,N_12);
and U4565 (N_4565,N_1058,N_172);
nand U4566 (N_4566,N_298,N_512);
and U4567 (N_4567,N_383,N_630);
and U4568 (N_4568,N_420,N_1557);
and U4569 (N_4569,N_1741,N_1714);
nor U4570 (N_4570,N_2047,N_1671);
nor U4571 (N_4571,N_17,N_1426);
nor U4572 (N_4572,N_1765,N_779);
and U4573 (N_4573,N_852,N_1496);
and U4574 (N_4574,N_10,N_383);
nor U4575 (N_4575,N_1477,N_2375);
and U4576 (N_4576,N_526,N_151);
nand U4577 (N_4577,N_946,N_825);
nand U4578 (N_4578,N_1116,N_2031);
nor U4579 (N_4579,N_713,N_2419);
nor U4580 (N_4580,N_543,N_274);
nor U4581 (N_4581,N_1592,N_1737);
or U4582 (N_4582,N_2433,N_1875);
or U4583 (N_4583,N_1876,N_2160);
nand U4584 (N_4584,N_981,N_2192);
and U4585 (N_4585,N_1328,N_1626);
or U4586 (N_4586,N_901,N_2484);
or U4587 (N_4587,N_124,N_520);
nor U4588 (N_4588,N_1725,N_675);
or U4589 (N_4589,N_4,N_1775);
and U4590 (N_4590,N_1762,N_940);
and U4591 (N_4591,N_842,N_1387);
and U4592 (N_4592,N_957,N_1090);
and U4593 (N_4593,N_20,N_1208);
nand U4594 (N_4594,N_1110,N_2085);
nand U4595 (N_4595,N_280,N_368);
nand U4596 (N_4596,N_1284,N_1446);
nor U4597 (N_4597,N_138,N_1885);
nor U4598 (N_4598,N_1324,N_1606);
and U4599 (N_4599,N_1299,N_2085);
nand U4600 (N_4600,N_1322,N_2057);
or U4601 (N_4601,N_180,N_196);
nor U4602 (N_4602,N_1747,N_1926);
nand U4603 (N_4603,N_2482,N_443);
and U4604 (N_4604,N_1912,N_255);
or U4605 (N_4605,N_1252,N_1702);
and U4606 (N_4606,N_1198,N_932);
and U4607 (N_4607,N_377,N_800);
nor U4608 (N_4608,N_2281,N_2000);
xor U4609 (N_4609,N_1831,N_971);
nand U4610 (N_4610,N_2422,N_228);
nor U4611 (N_4611,N_1115,N_74);
nand U4612 (N_4612,N_786,N_268);
or U4613 (N_4613,N_583,N_896);
or U4614 (N_4614,N_493,N_2412);
xor U4615 (N_4615,N_1502,N_2299);
or U4616 (N_4616,N_1877,N_2469);
or U4617 (N_4617,N_1576,N_382);
or U4618 (N_4618,N_1510,N_1419);
nor U4619 (N_4619,N_884,N_1391);
or U4620 (N_4620,N_1387,N_21);
or U4621 (N_4621,N_415,N_2382);
or U4622 (N_4622,N_1862,N_726);
nand U4623 (N_4623,N_455,N_2114);
nor U4624 (N_4624,N_197,N_2259);
and U4625 (N_4625,N_1790,N_2174);
nand U4626 (N_4626,N_368,N_893);
nor U4627 (N_4627,N_2238,N_2105);
and U4628 (N_4628,N_2337,N_1396);
nor U4629 (N_4629,N_78,N_1769);
and U4630 (N_4630,N_2270,N_692);
or U4631 (N_4631,N_1642,N_1619);
and U4632 (N_4632,N_1969,N_1123);
nand U4633 (N_4633,N_1280,N_976);
or U4634 (N_4634,N_309,N_889);
nand U4635 (N_4635,N_86,N_599);
nor U4636 (N_4636,N_2253,N_2299);
or U4637 (N_4637,N_1830,N_2313);
nand U4638 (N_4638,N_1774,N_1432);
or U4639 (N_4639,N_564,N_773);
nor U4640 (N_4640,N_1947,N_1423);
or U4641 (N_4641,N_524,N_992);
nand U4642 (N_4642,N_115,N_2184);
nand U4643 (N_4643,N_90,N_140);
nor U4644 (N_4644,N_938,N_318);
or U4645 (N_4645,N_1961,N_646);
nand U4646 (N_4646,N_640,N_733);
nor U4647 (N_4647,N_2335,N_1190);
and U4648 (N_4648,N_1154,N_879);
and U4649 (N_4649,N_1695,N_1347);
and U4650 (N_4650,N_705,N_1256);
or U4651 (N_4651,N_1852,N_1228);
or U4652 (N_4652,N_28,N_1112);
or U4653 (N_4653,N_428,N_1359);
and U4654 (N_4654,N_2012,N_1378);
or U4655 (N_4655,N_2279,N_2009);
nand U4656 (N_4656,N_2304,N_1060);
and U4657 (N_4657,N_1845,N_883);
nor U4658 (N_4658,N_1742,N_1852);
or U4659 (N_4659,N_2079,N_243);
nand U4660 (N_4660,N_2289,N_2235);
nand U4661 (N_4661,N_46,N_2342);
nand U4662 (N_4662,N_1304,N_982);
or U4663 (N_4663,N_468,N_49);
and U4664 (N_4664,N_421,N_792);
nand U4665 (N_4665,N_1246,N_469);
nand U4666 (N_4666,N_282,N_394);
nor U4667 (N_4667,N_691,N_340);
nand U4668 (N_4668,N_1566,N_984);
and U4669 (N_4669,N_859,N_1935);
nand U4670 (N_4670,N_1560,N_131);
nor U4671 (N_4671,N_1150,N_1207);
nand U4672 (N_4672,N_1023,N_73);
and U4673 (N_4673,N_155,N_767);
nor U4674 (N_4674,N_2483,N_328);
and U4675 (N_4675,N_2293,N_222);
nor U4676 (N_4676,N_1298,N_1170);
nand U4677 (N_4677,N_2223,N_2158);
nand U4678 (N_4678,N_93,N_325);
nor U4679 (N_4679,N_2239,N_471);
or U4680 (N_4680,N_1103,N_2100);
and U4681 (N_4681,N_549,N_1716);
nand U4682 (N_4682,N_2272,N_1244);
or U4683 (N_4683,N_1712,N_738);
nand U4684 (N_4684,N_2374,N_436);
nand U4685 (N_4685,N_178,N_1959);
nand U4686 (N_4686,N_1752,N_633);
nand U4687 (N_4687,N_1418,N_2349);
and U4688 (N_4688,N_893,N_1160);
and U4689 (N_4689,N_2039,N_961);
nand U4690 (N_4690,N_1004,N_2089);
and U4691 (N_4691,N_49,N_1975);
nand U4692 (N_4692,N_1140,N_294);
nand U4693 (N_4693,N_1206,N_2237);
and U4694 (N_4694,N_257,N_1451);
nor U4695 (N_4695,N_405,N_133);
and U4696 (N_4696,N_1017,N_1753);
nand U4697 (N_4697,N_67,N_2091);
and U4698 (N_4698,N_326,N_1811);
nand U4699 (N_4699,N_801,N_1923);
nor U4700 (N_4700,N_1994,N_1335);
nand U4701 (N_4701,N_1624,N_1333);
nor U4702 (N_4702,N_908,N_929);
and U4703 (N_4703,N_212,N_1378);
or U4704 (N_4704,N_686,N_2285);
nor U4705 (N_4705,N_441,N_299);
nand U4706 (N_4706,N_468,N_952);
and U4707 (N_4707,N_77,N_1624);
and U4708 (N_4708,N_94,N_2370);
nor U4709 (N_4709,N_2489,N_492);
nor U4710 (N_4710,N_2466,N_1606);
or U4711 (N_4711,N_2065,N_1932);
and U4712 (N_4712,N_2065,N_983);
and U4713 (N_4713,N_366,N_1850);
nor U4714 (N_4714,N_1965,N_54);
nor U4715 (N_4715,N_651,N_1728);
nor U4716 (N_4716,N_965,N_355);
or U4717 (N_4717,N_1473,N_1621);
nand U4718 (N_4718,N_2193,N_2081);
or U4719 (N_4719,N_2108,N_211);
nor U4720 (N_4720,N_1487,N_1952);
or U4721 (N_4721,N_1258,N_398);
nor U4722 (N_4722,N_585,N_1074);
nand U4723 (N_4723,N_750,N_1658);
nand U4724 (N_4724,N_376,N_2231);
nor U4725 (N_4725,N_1321,N_2189);
or U4726 (N_4726,N_639,N_396);
or U4727 (N_4727,N_479,N_1525);
or U4728 (N_4728,N_968,N_714);
and U4729 (N_4729,N_250,N_1015);
and U4730 (N_4730,N_2330,N_212);
xor U4731 (N_4731,N_1196,N_1990);
and U4732 (N_4732,N_1930,N_2492);
and U4733 (N_4733,N_1188,N_607);
nor U4734 (N_4734,N_1711,N_1477);
nor U4735 (N_4735,N_435,N_2195);
or U4736 (N_4736,N_454,N_1695);
nand U4737 (N_4737,N_2189,N_1822);
nor U4738 (N_4738,N_1258,N_1861);
or U4739 (N_4739,N_1656,N_1676);
and U4740 (N_4740,N_1594,N_1201);
nor U4741 (N_4741,N_1532,N_1993);
nand U4742 (N_4742,N_945,N_1798);
nand U4743 (N_4743,N_1822,N_1438);
xor U4744 (N_4744,N_1596,N_915);
nor U4745 (N_4745,N_196,N_2446);
and U4746 (N_4746,N_983,N_2098);
and U4747 (N_4747,N_1964,N_433);
nand U4748 (N_4748,N_1541,N_413);
nand U4749 (N_4749,N_728,N_1326);
xnor U4750 (N_4750,N_1767,N_1324);
and U4751 (N_4751,N_1858,N_2231);
nor U4752 (N_4752,N_11,N_762);
nor U4753 (N_4753,N_2184,N_955);
or U4754 (N_4754,N_1954,N_2336);
nand U4755 (N_4755,N_2240,N_772);
nand U4756 (N_4756,N_344,N_458);
or U4757 (N_4757,N_2499,N_263);
or U4758 (N_4758,N_1343,N_2483);
or U4759 (N_4759,N_773,N_1236);
and U4760 (N_4760,N_338,N_1635);
nand U4761 (N_4761,N_1518,N_2176);
or U4762 (N_4762,N_141,N_1665);
or U4763 (N_4763,N_2229,N_2034);
and U4764 (N_4764,N_2095,N_1444);
and U4765 (N_4765,N_250,N_303);
nand U4766 (N_4766,N_2361,N_2216);
nand U4767 (N_4767,N_1339,N_1473);
nor U4768 (N_4768,N_2063,N_1925);
nor U4769 (N_4769,N_2118,N_2164);
and U4770 (N_4770,N_517,N_1591);
nand U4771 (N_4771,N_1597,N_1188);
nand U4772 (N_4772,N_385,N_891);
and U4773 (N_4773,N_2404,N_1384);
or U4774 (N_4774,N_397,N_1309);
nand U4775 (N_4775,N_649,N_2337);
nor U4776 (N_4776,N_727,N_1249);
and U4777 (N_4777,N_923,N_1811);
or U4778 (N_4778,N_1115,N_1575);
and U4779 (N_4779,N_1241,N_153);
or U4780 (N_4780,N_885,N_530);
nor U4781 (N_4781,N_668,N_2438);
nor U4782 (N_4782,N_866,N_1833);
or U4783 (N_4783,N_1450,N_1540);
xor U4784 (N_4784,N_2110,N_2235);
or U4785 (N_4785,N_116,N_1175);
and U4786 (N_4786,N_1239,N_2233);
and U4787 (N_4787,N_2477,N_1225);
xor U4788 (N_4788,N_627,N_2094);
nand U4789 (N_4789,N_1713,N_1935);
nor U4790 (N_4790,N_1226,N_1941);
xnor U4791 (N_4791,N_2421,N_617);
and U4792 (N_4792,N_432,N_402);
nor U4793 (N_4793,N_146,N_1352);
nor U4794 (N_4794,N_315,N_763);
nand U4795 (N_4795,N_63,N_981);
and U4796 (N_4796,N_1096,N_1637);
nor U4797 (N_4797,N_1006,N_898);
nor U4798 (N_4798,N_425,N_7);
or U4799 (N_4799,N_560,N_2077);
nor U4800 (N_4800,N_175,N_2006);
and U4801 (N_4801,N_328,N_128);
nor U4802 (N_4802,N_136,N_1821);
nor U4803 (N_4803,N_1723,N_554);
and U4804 (N_4804,N_1538,N_2140);
nor U4805 (N_4805,N_1597,N_657);
or U4806 (N_4806,N_172,N_1146);
nand U4807 (N_4807,N_875,N_879);
nand U4808 (N_4808,N_1460,N_1696);
nor U4809 (N_4809,N_1162,N_1163);
or U4810 (N_4810,N_1221,N_2322);
nor U4811 (N_4811,N_1216,N_881);
or U4812 (N_4812,N_1356,N_1407);
nor U4813 (N_4813,N_278,N_815);
or U4814 (N_4814,N_1696,N_192);
or U4815 (N_4815,N_2213,N_1818);
and U4816 (N_4816,N_2323,N_2350);
and U4817 (N_4817,N_2013,N_579);
or U4818 (N_4818,N_631,N_2335);
nor U4819 (N_4819,N_2043,N_293);
and U4820 (N_4820,N_494,N_735);
or U4821 (N_4821,N_601,N_204);
and U4822 (N_4822,N_1945,N_934);
or U4823 (N_4823,N_2046,N_86);
or U4824 (N_4824,N_1879,N_1562);
nor U4825 (N_4825,N_2479,N_263);
and U4826 (N_4826,N_463,N_61);
nor U4827 (N_4827,N_1884,N_1454);
or U4828 (N_4828,N_1684,N_20);
and U4829 (N_4829,N_1051,N_1363);
nand U4830 (N_4830,N_670,N_2207);
nand U4831 (N_4831,N_2190,N_1864);
and U4832 (N_4832,N_1599,N_1977);
and U4833 (N_4833,N_311,N_2357);
and U4834 (N_4834,N_1004,N_2347);
or U4835 (N_4835,N_2280,N_2433);
and U4836 (N_4836,N_925,N_2266);
nor U4837 (N_4837,N_460,N_248);
nor U4838 (N_4838,N_1541,N_1092);
nor U4839 (N_4839,N_331,N_2432);
nor U4840 (N_4840,N_1863,N_1025);
and U4841 (N_4841,N_539,N_2449);
nand U4842 (N_4842,N_496,N_1252);
or U4843 (N_4843,N_863,N_2389);
or U4844 (N_4844,N_1572,N_1923);
nor U4845 (N_4845,N_1352,N_247);
nand U4846 (N_4846,N_1311,N_1063);
nor U4847 (N_4847,N_1590,N_274);
nor U4848 (N_4848,N_2229,N_1530);
or U4849 (N_4849,N_261,N_1169);
nand U4850 (N_4850,N_289,N_1839);
and U4851 (N_4851,N_1406,N_1382);
nand U4852 (N_4852,N_1144,N_193);
nand U4853 (N_4853,N_2073,N_10);
nor U4854 (N_4854,N_677,N_357);
nand U4855 (N_4855,N_678,N_91);
nand U4856 (N_4856,N_186,N_2381);
or U4857 (N_4857,N_868,N_1662);
nor U4858 (N_4858,N_1701,N_520);
and U4859 (N_4859,N_1570,N_1771);
and U4860 (N_4860,N_1995,N_486);
and U4861 (N_4861,N_2058,N_2432);
nand U4862 (N_4862,N_2236,N_2144);
and U4863 (N_4863,N_317,N_2042);
nand U4864 (N_4864,N_1294,N_1488);
nor U4865 (N_4865,N_2182,N_1709);
nor U4866 (N_4866,N_1906,N_1244);
nor U4867 (N_4867,N_309,N_677);
nand U4868 (N_4868,N_518,N_1673);
nand U4869 (N_4869,N_2228,N_252);
and U4870 (N_4870,N_1561,N_99);
or U4871 (N_4871,N_1497,N_694);
nand U4872 (N_4872,N_2321,N_92);
and U4873 (N_4873,N_1539,N_2310);
nor U4874 (N_4874,N_290,N_2329);
and U4875 (N_4875,N_2454,N_314);
nand U4876 (N_4876,N_579,N_1563);
and U4877 (N_4877,N_362,N_1883);
nor U4878 (N_4878,N_2257,N_2459);
or U4879 (N_4879,N_1170,N_1491);
or U4880 (N_4880,N_165,N_961);
nand U4881 (N_4881,N_1817,N_1926);
or U4882 (N_4882,N_2234,N_2146);
and U4883 (N_4883,N_70,N_582);
or U4884 (N_4884,N_1145,N_2144);
nand U4885 (N_4885,N_759,N_181);
nand U4886 (N_4886,N_1317,N_1274);
nand U4887 (N_4887,N_892,N_2077);
and U4888 (N_4888,N_266,N_96);
or U4889 (N_4889,N_1240,N_242);
nand U4890 (N_4890,N_963,N_1200);
or U4891 (N_4891,N_200,N_874);
nand U4892 (N_4892,N_1378,N_729);
and U4893 (N_4893,N_2474,N_1038);
nand U4894 (N_4894,N_2449,N_919);
nor U4895 (N_4895,N_1351,N_1946);
and U4896 (N_4896,N_336,N_410);
and U4897 (N_4897,N_1809,N_1245);
and U4898 (N_4898,N_2127,N_1889);
and U4899 (N_4899,N_1508,N_199);
and U4900 (N_4900,N_2456,N_1200);
nor U4901 (N_4901,N_1782,N_1512);
or U4902 (N_4902,N_1386,N_310);
nor U4903 (N_4903,N_755,N_873);
nor U4904 (N_4904,N_1467,N_451);
or U4905 (N_4905,N_1053,N_2336);
and U4906 (N_4906,N_345,N_1100);
and U4907 (N_4907,N_213,N_1605);
or U4908 (N_4908,N_1999,N_1931);
or U4909 (N_4909,N_405,N_750);
nand U4910 (N_4910,N_664,N_1997);
or U4911 (N_4911,N_1141,N_1497);
nand U4912 (N_4912,N_2197,N_519);
and U4913 (N_4913,N_1944,N_1965);
or U4914 (N_4914,N_996,N_262);
nor U4915 (N_4915,N_1828,N_165);
nor U4916 (N_4916,N_1316,N_724);
nand U4917 (N_4917,N_496,N_90);
or U4918 (N_4918,N_1105,N_599);
nor U4919 (N_4919,N_1636,N_1145);
and U4920 (N_4920,N_339,N_452);
nand U4921 (N_4921,N_770,N_945);
and U4922 (N_4922,N_606,N_227);
and U4923 (N_4923,N_493,N_1555);
and U4924 (N_4924,N_1711,N_230);
and U4925 (N_4925,N_1724,N_1843);
nand U4926 (N_4926,N_1944,N_1127);
and U4927 (N_4927,N_2411,N_1019);
nor U4928 (N_4928,N_996,N_832);
nand U4929 (N_4929,N_2258,N_1835);
nand U4930 (N_4930,N_81,N_1715);
nor U4931 (N_4931,N_1713,N_178);
nand U4932 (N_4932,N_748,N_531);
and U4933 (N_4933,N_2486,N_2188);
nor U4934 (N_4934,N_1753,N_2484);
or U4935 (N_4935,N_2246,N_475);
or U4936 (N_4936,N_859,N_1635);
nand U4937 (N_4937,N_2463,N_2416);
nand U4938 (N_4938,N_1989,N_1797);
nor U4939 (N_4939,N_1251,N_567);
nand U4940 (N_4940,N_999,N_1475);
and U4941 (N_4941,N_1770,N_1688);
or U4942 (N_4942,N_1971,N_533);
nor U4943 (N_4943,N_1534,N_1667);
nor U4944 (N_4944,N_363,N_1601);
nor U4945 (N_4945,N_1792,N_7);
or U4946 (N_4946,N_1554,N_464);
and U4947 (N_4947,N_1719,N_2394);
nor U4948 (N_4948,N_116,N_1780);
nand U4949 (N_4949,N_2048,N_2337);
nand U4950 (N_4950,N_447,N_1616);
nor U4951 (N_4951,N_387,N_1784);
and U4952 (N_4952,N_814,N_673);
nand U4953 (N_4953,N_248,N_867);
or U4954 (N_4954,N_1310,N_1187);
or U4955 (N_4955,N_2016,N_2463);
nor U4956 (N_4956,N_1307,N_1881);
or U4957 (N_4957,N_34,N_2360);
or U4958 (N_4958,N_626,N_372);
and U4959 (N_4959,N_562,N_2451);
or U4960 (N_4960,N_1659,N_551);
or U4961 (N_4961,N_1417,N_1569);
and U4962 (N_4962,N_630,N_726);
and U4963 (N_4963,N_2480,N_1849);
nand U4964 (N_4964,N_144,N_1659);
nand U4965 (N_4965,N_1459,N_211);
nor U4966 (N_4966,N_1559,N_606);
nor U4967 (N_4967,N_1308,N_1747);
or U4968 (N_4968,N_347,N_780);
and U4969 (N_4969,N_684,N_1070);
and U4970 (N_4970,N_73,N_1234);
and U4971 (N_4971,N_2050,N_708);
and U4972 (N_4972,N_308,N_1996);
or U4973 (N_4973,N_1465,N_2354);
or U4974 (N_4974,N_1691,N_1742);
nand U4975 (N_4975,N_373,N_469);
or U4976 (N_4976,N_2193,N_707);
or U4977 (N_4977,N_1071,N_2043);
nor U4978 (N_4978,N_724,N_713);
nor U4979 (N_4979,N_1854,N_2057);
nand U4980 (N_4980,N_447,N_117);
or U4981 (N_4981,N_277,N_635);
or U4982 (N_4982,N_2114,N_2442);
and U4983 (N_4983,N_1027,N_1062);
or U4984 (N_4984,N_1396,N_688);
and U4985 (N_4985,N_2490,N_230);
and U4986 (N_4986,N_1464,N_264);
nand U4987 (N_4987,N_1762,N_224);
nand U4988 (N_4988,N_851,N_1382);
and U4989 (N_4989,N_499,N_189);
nor U4990 (N_4990,N_913,N_282);
nand U4991 (N_4991,N_1501,N_1698);
or U4992 (N_4992,N_2181,N_1486);
and U4993 (N_4993,N_1297,N_557);
nor U4994 (N_4994,N_853,N_81);
nand U4995 (N_4995,N_267,N_185);
nand U4996 (N_4996,N_1123,N_2464);
and U4997 (N_4997,N_455,N_691);
nor U4998 (N_4998,N_427,N_43);
nor U4999 (N_4999,N_2296,N_2351);
and UO_0 (O_0,N_3207,N_3971);
nor UO_1 (O_1,N_3782,N_2507);
nand UO_2 (O_2,N_2502,N_4083);
or UO_3 (O_3,N_2668,N_4537);
nor UO_4 (O_4,N_3058,N_3988);
nand UO_5 (O_5,N_3658,N_4061);
or UO_6 (O_6,N_2938,N_2914);
or UO_7 (O_7,N_3955,N_4165);
nand UO_8 (O_8,N_2721,N_3612);
nand UO_9 (O_9,N_3476,N_4596);
nor UO_10 (O_10,N_4179,N_3602);
and UO_11 (O_11,N_3960,N_3814);
nand UO_12 (O_12,N_3150,N_3628);
or UO_13 (O_13,N_2982,N_3407);
or UO_14 (O_14,N_3209,N_3082);
nor UO_15 (O_15,N_4079,N_2822);
nand UO_16 (O_16,N_4976,N_4706);
nand UO_17 (O_17,N_3416,N_3226);
and UO_18 (O_18,N_2688,N_2819);
or UO_19 (O_19,N_4378,N_4199);
or UO_20 (O_20,N_3141,N_3086);
or UO_21 (O_21,N_3275,N_4406);
nand UO_22 (O_22,N_4759,N_3378);
nor UO_23 (O_23,N_4355,N_3497);
or UO_24 (O_24,N_4628,N_3484);
nand UO_25 (O_25,N_4488,N_3170);
nor UO_26 (O_26,N_3043,N_3625);
or UO_27 (O_27,N_4287,N_2978);
and UO_28 (O_28,N_4042,N_2797);
nor UO_29 (O_29,N_3469,N_4196);
or UO_30 (O_30,N_2807,N_3970);
nand UO_31 (O_31,N_3806,N_3601);
nand UO_32 (O_32,N_3269,N_4238);
or UO_33 (O_33,N_3600,N_4605);
and UO_34 (O_34,N_2790,N_4215);
nor UO_35 (O_35,N_3107,N_3690);
and UO_36 (O_36,N_2707,N_4169);
and UO_37 (O_37,N_2760,N_3506);
and UO_38 (O_38,N_3376,N_4591);
nand UO_39 (O_39,N_3899,N_3334);
nor UO_40 (O_40,N_4340,N_3291);
and UO_41 (O_41,N_3090,N_3490);
nand UO_42 (O_42,N_2521,N_4329);
and UO_43 (O_43,N_3280,N_3488);
nand UO_44 (O_44,N_4222,N_3403);
nor UO_45 (O_45,N_2630,N_4712);
or UO_46 (O_46,N_4508,N_4352);
nand UO_47 (O_47,N_4782,N_4858);
nor UO_48 (O_48,N_2952,N_2934);
and UO_49 (O_49,N_3460,N_3367);
nor UO_50 (O_50,N_4996,N_2508);
nor UO_51 (O_51,N_3801,N_4460);
nand UO_52 (O_52,N_4109,N_4433);
nor UO_53 (O_53,N_3168,N_3520);
nand UO_54 (O_54,N_4609,N_3500);
and UO_55 (O_55,N_4515,N_3202);
and UO_56 (O_56,N_4161,N_4411);
and UO_57 (O_57,N_3105,N_3697);
and UO_58 (O_58,N_4725,N_2643);
or UO_59 (O_59,N_2636,N_4321);
nand UO_60 (O_60,N_3229,N_4728);
nand UO_61 (O_61,N_3359,N_4846);
nand UO_62 (O_62,N_2960,N_2970);
and UO_63 (O_63,N_3446,N_2851);
nand UO_64 (O_64,N_4495,N_4980);
nand UO_65 (O_65,N_4936,N_2951);
or UO_66 (O_66,N_3253,N_2977);
nand UO_67 (O_67,N_3708,N_3379);
nor UO_68 (O_68,N_4990,N_3604);
or UO_69 (O_69,N_3638,N_4060);
nand UO_70 (O_70,N_2766,N_4805);
or UO_71 (O_71,N_4594,N_4844);
or UO_72 (O_72,N_4652,N_3223);
nand UO_73 (O_73,N_3178,N_4659);
nand UO_74 (O_74,N_3187,N_3112);
nor UO_75 (O_75,N_3211,N_4836);
nor UO_76 (O_76,N_3206,N_3616);
nand UO_77 (O_77,N_4931,N_3522);
and UO_78 (O_78,N_3032,N_4347);
nor UO_79 (O_79,N_4264,N_3123);
or UO_80 (O_80,N_4517,N_3406);
or UO_81 (O_81,N_3426,N_4539);
or UO_82 (O_82,N_3585,N_4632);
or UO_83 (O_83,N_4981,N_2834);
nor UO_84 (O_84,N_4545,N_4952);
nand UO_85 (O_85,N_2620,N_2702);
nand UO_86 (O_86,N_3485,N_3339);
nand UO_87 (O_87,N_4731,N_3576);
and UO_88 (O_88,N_3836,N_4840);
nand UO_89 (O_89,N_3528,N_3608);
nor UO_90 (O_90,N_3336,N_3871);
nor UO_91 (O_91,N_2555,N_3422);
nor UO_92 (O_92,N_4558,N_3691);
or UO_93 (O_93,N_4441,N_3412);
nand UO_94 (O_94,N_3870,N_4570);
or UO_95 (O_95,N_4392,N_3741);
or UO_96 (O_96,N_2713,N_2823);
nand UO_97 (O_97,N_3617,N_4114);
or UO_98 (O_98,N_2672,N_3261);
and UO_99 (O_99,N_4721,N_3863);
or UO_100 (O_100,N_2955,N_3290);
and UO_101 (O_101,N_4895,N_4281);
nand UO_102 (O_102,N_4830,N_2648);
or UO_103 (O_103,N_3595,N_2671);
or UO_104 (O_104,N_3360,N_3586);
and UO_105 (O_105,N_3243,N_2769);
nor UO_106 (O_106,N_2910,N_3154);
or UO_107 (O_107,N_4040,N_3950);
nor UO_108 (O_108,N_4939,N_2776);
nand UO_109 (O_109,N_3083,N_3231);
nor UO_110 (O_110,N_2733,N_2979);
nor UO_111 (O_111,N_3688,N_3309);
nand UO_112 (O_112,N_3716,N_3965);
and UO_113 (O_113,N_2520,N_3366);
and UO_114 (O_114,N_4143,N_3319);
and UO_115 (O_115,N_3259,N_3848);
and UO_116 (O_116,N_3343,N_4229);
nor UO_117 (O_117,N_3751,N_4898);
and UO_118 (O_118,N_4239,N_4851);
or UO_119 (O_119,N_3167,N_4194);
nor UO_120 (O_120,N_3800,N_2698);
nor UO_121 (O_121,N_3008,N_3893);
nor UO_122 (O_122,N_3943,N_4681);
nand UO_123 (O_123,N_3192,N_3962);
or UO_124 (O_124,N_3000,N_2731);
xnor UO_125 (O_125,N_3792,N_4214);
nand UO_126 (O_126,N_4972,N_3872);
or UO_127 (O_127,N_2925,N_2644);
nand UO_128 (O_128,N_4003,N_2916);
and UO_129 (O_129,N_2569,N_3938);
or UO_130 (O_130,N_3627,N_4538);
or UO_131 (O_131,N_3824,N_2618);
or UO_132 (O_132,N_4404,N_2768);
and UO_133 (O_133,N_3745,N_4465);
and UO_134 (O_134,N_3817,N_4501);
nor UO_135 (O_135,N_3920,N_4059);
nor UO_136 (O_136,N_2711,N_3993);
or UO_137 (O_137,N_2641,N_4354);
and UO_138 (O_138,N_3513,N_4476);
nand UO_139 (O_139,N_3656,N_4644);
or UO_140 (O_140,N_3858,N_3208);
and UO_141 (O_141,N_3514,N_3268);
nand UO_142 (O_142,N_4984,N_2597);
or UO_143 (O_143,N_2828,N_3951);
and UO_144 (O_144,N_2545,N_3624);
and UO_145 (O_145,N_4136,N_2541);
or UO_146 (O_146,N_3278,N_4751);
nor UO_147 (O_147,N_3250,N_4453);
and UO_148 (O_148,N_3694,N_4250);
nor UO_149 (O_149,N_3717,N_3040);
and UO_150 (O_150,N_3689,N_4107);
nand UO_151 (O_151,N_3020,N_2767);
and UO_152 (O_152,N_4603,N_3124);
and UO_153 (O_153,N_4801,N_4915);
xnor UO_154 (O_154,N_4074,N_4758);
nand UO_155 (O_155,N_4492,N_4927);
nor UO_156 (O_156,N_4600,N_3735);
nor UO_157 (O_157,N_4084,N_2676);
and UO_158 (O_158,N_4479,N_3837);
nand UO_159 (O_159,N_2558,N_2747);
nand UO_160 (O_160,N_3465,N_2853);
or UO_161 (O_161,N_4171,N_3411);
nor UO_162 (O_162,N_3557,N_4919);
nand UO_163 (O_163,N_3244,N_3232);
or UO_164 (O_164,N_3597,N_4422);
nor UO_165 (O_165,N_3193,N_4982);
and UO_166 (O_166,N_4975,N_3059);
nand UO_167 (O_167,N_3932,N_2739);
nor UO_168 (O_168,N_2517,N_3797);
or UO_169 (O_169,N_4693,N_2538);
nor UO_170 (O_170,N_3701,N_4708);
nor UO_171 (O_171,N_3757,N_3031);
and UO_172 (O_172,N_3286,N_2593);
or UO_173 (O_173,N_3982,N_4743);
nand UO_174 (O_174,N_2813,N_4299);
nand UO_175 (O_175,N_3175,N_2946);
and UO_176 (O_176,N_2515,N_4856);
and UO_177 (O_177,N_3368,N_3472);
and UO_178 (O_178,N_4497,N_3523);
or UO_179 (O_179,N_3821,N_4124);
and UO_180 (O_180,N_4588,N_4374);
nor UO_181 (O_181,N_4121,N_4247);
and UO_182 (O_182,N_4684,N_4173);
and UO_183 (O_183,N_2932,N_2619);
and UO_184 (O_184,N_4740,N_2948);
nand UO_185 (O_185,N_2919,N_4713);
or UO_186 (O_186,N_3001,N_3048);
and UO_187 (O_187,N_4963,N_4737);
and UO_188 (O_188,N_3544,N_4616);
nor UO_189 (O_189,N_4401,N_3096);
nand UO_190 (O_190,N_4694,N_4097);
or UO_191 (O_191,N_3205,N_2971);
or UO_192 (O_192,N_3163,N_2887);
nand UO_193 (O_193,N_4138,N_3120);
and UO_194 (O_194,N_3762,N_4385);
nand UO_195 (O_195,N_3569,N_4387);
and UO_196 (O_196,N_3764,N_3867);
nand UO_197 (O_197,N_3789,N_2685);
and UO_198 (O_198,N_2678,N_4486);
nand UO_199 (O_199,N_4296,N_2832);
and UO_200 (O_200,N_4923,N_3816);
nand UO_201 (O_201,N_4978,N_3387);
nor UO_202 (O_202,N_2679,N_3714);
nor UO_203 (O_203,N_3603,N_4704);
or UO_204 (O_204,N_2991,N_3418);
nand UO_205 (O_205,N_4668,N_4823);
nor UO_206 (O_206,N_4529,N_4016);
and UO_207 (O_207,N_2717,N_3969);
nand UO_208 (O_208,N_3554,N_4292);
and UO_209 (O_209,N_3341,N_4436);
nor UO_210 (O_210,N_4951,N_2567);
nand UO_211 (O_211,N_4509,N_3521);
and UO_212 (O_212,N_3843,N_3394);
or UO_213 (O_213,N_3165,N_3834);
nor UO_214 (O_214,N_3479,N_3855);
and UO_215 (O_215,N_3350,N_4957);
nor UO_216 (O_216,N_3300,N_3940);
or UO_217 (O_217,N_3731,N_4774);
xnor UO_218 (O_218,N_4498,N_2616);
nor UO_219 (O_219,N_3203,N_3256);
and UO_220 (O_220,N_3692,N_4983);
or UO_221 (O_221,N_3307,N_4614);
or UO_222 (O_222,N_2604,N_3636);
nand UO_223 (O_223,N_4253,N_3335);
nor UO_224 (O_224,N_4457,N_4156);
or UO_225 (O_225,N_3537,N_4064);
and UO_226 (O_226,N_4940,N_4870);
or UO_227 (O_227,N_3649,N_4223);
nand UO_228 (O_228,N_3062,N_2728);
nand UO_229 (O_229,N_4680,N_4129);
nand UO_230 (O_230,N_3380,N_4986);
nand UO_231 (O_231,N_2556,N_4849);
and UO_232 (O_232,N_3087,N_4637);
nor UO_233 (O_233,N_3067,N_4466);
nand UO_234 (O_234,N_4028,N_3161);
and UO_235 (O_235,N_4626,N_3505);
and UO_236 (O_236,N_3743,N_3089);
or UO_237 (O_237,N_3633,N_3265);
nor UO_238 (O_238,N_4450,N_3491);
and UO_239 (O_239,N_2692,N_4262);
nor UO_240 (O_240,N_3986,N_4362);
and UO_241 (O_241,N_3769,N_2596);
nor UO_242 (O_242,N_2664,N_4912);
and UO_243 (O_243,N_4388,N_3420);
and UO_244 (O_244,N_4125,N_4874);
nor UO_245 (O_245,N_4944,N_4225);
or UO_246 (O_246,N_2729,N_3483);
nor UO_247 (O_247,N_3776,N_3949);
nand UO_248 (O_248,N_3473,N_3910);
nand UO_249 (O_249,N_2594,N_4033);
or UO_250 (O_250,N_4013,N_3279);
or UO_251 (O_251,N_2795,N_4688);
or UO_252 (O_252,N_4617,N_4689);
nand UO_253 (O_253,N_4270,N_4930);
and UO_254 (O_254,N_3941,N_4315);
xnor UO_255 (O_255,N_2561,N_2646);
nor UO_256 (O_256,N_4932,N_3937);
nand UO_257 (O_257,N_2592,N_3662);
nor UO_258 (O_258,N_3158,N_4023);
nor UO_259 (O_259,N_3314,N_4833);
nand UO_260 (O_260,N_4857,N_4555);
nor UO_261 (O_261,N_4654,N_4190);
or UO_262 (O_262,N_3091,N_3695);
nor UO_263 (O_263,N_4108,N_4993);
nor UO_264 (O_264,N_4418,N_3615);
and UO_265 (O_265,N_3593,N_4606);
nor UO_266 (O_266,N_4968,N_3475);
and UO_267 (O_267,N_4564,N_4232);
nor UO_268 (O_268,N_3864,N_3053);
and UO_269 (O_269,N_3103,N_4788);
nand UO_270 (O_270,N_2708,N_3034);
nor UO_271 (O_271,N_2599,N_4373);
and UO_272 (O_272,N_3549,N_2566);
nand UO_273 (O_273,N_3444,N_4301);
or UO_274 (O_274,N_4044,N_3880);
nor UO_275 (O_275,N_4757,N_3092);
or UO_276 (O_276,N_4648,N_4322);
and UO_277 (O_277,N_2875,N_4487);
or UO_278 (O_278,N_3423,N_4428);
nor UO_279 (O_279,N_3997,N_4878);
nor UO_280 (O_280,N_3079,N_3921);
nand UO_281 (O_281,N_4750,N_3263);
nor UO_282 (O_282,N_3791,N_4141);
and UO_283 (O_283,N_2831,N_4516);
and UO_284 (O_284,N_2950,N_2897);
and UO_285 (O_285,N_3143,N_2613);
nand UO_286 (O_286,N_4739,N_2751);
nand UO_287 (O_287,N_3954,N_2696);
and UO_288 (O_288,N_3642,N_4078);
or UO_289 (O_289,N_4472,N_2589);
or UO_290 (O_290,N_4482,N_4180);
nor UO_291 (O_291,N_3807,N_4293);
and UO_292 (O_292,N_2968,N_3742);
or UO_293 (O_293,N_4563,N_4150);
nor UO_294 (O_294,N_3754,N_4916);
nor UO_295 (O_295,N_4473,N_3630);
and UO_296 (O_296,N_3272,N_4650);
nand UO_297 (O_297,N_3156,N_3122);
nand UO_298 (O_298,N_4348,N_4571);
nand UO_299 (O_299,N_2898,N_3183);
nand UO_300 (O_300,N_3347,N_4234);
and UO_301 (O_301,N_2716,N_2762);
nand UO_302 (O_302,N_2778,N_3672);
nand UO_303 (O_303,N_2976,N_3527);
and UO_304 (O_304,N_3013,N_3942);
or UO_305 (O_305,N_2557,N_3765);
nor UO_306 (O_306,N_4202,N_4019);
and UO_307 (O_307,N_4716,N_2798);
or UO_308 (O_308,N_4252,N_4781);
and UO_309 (O_309,N_4618,N_2912);
or UO_310 (O_310,N_3676,N_4847);
or UO_311 (O_311,N_2974,N_3644);
nor UO_312 (O_312,N_2526,N_2940);
and UO_313 (O_313,N_4099,N_3240);
and UO_314 (O_314,N_4127,N_2773);
nor UO_315 (O_315,N_4267,N_3351);
or UO_316 (O_316,N_4368,N_4451);
and UO_317 (O_317,N_4191,N_3667);
nor UO_318 (O_318,N_4550,N_2837);
or UO_319 (O_319,N_3889,N_4396);
and UO_320 (O_320,N_2512,N_3978);
or UO_321 (O_321,N_4711,N_2927);
or UO_322 (O_322,N_4888,N_4703);
nand UO_323 (O_323,N_3666,N_4590);
and UO_324 (O_324,N_3248,N_3448);
nand UO_325 (O_325,N_4842,N_3646);
nor UO_326 (O_326,N_3856,N_3337);
or UO_327 (O_327,N_3866,N_3829);
and UO_328 (O_328,N_4926,N_3310);
or UO_329 (O_329,N_2758,N_3365);
and UO_330 (O_330,N_4192,N_4860);
or UO_331 (O_331,N_2872,N_4423);
nor UO_332 (O_332,N_3639,N_4050);
or UO_333 (O_333,N_2628,N_4146);
and UO_334 (O_334,N_2706,N_4656);
or UO_335 (O_335,N_3388,N_3101);
and UO_336 (O_336,N_3093,N_4265);
and UO_337 (O_337,N_4351,N_3673);
nand UO_338 (O_338,N_3219,N_2718);
nor UO_339 (O_339,N_2606,N_3548);
nand UO_340 (O_340,N_3029,N_4581);
nand UO_341 (O_341,N_3149,N_2661);
nand UO_342 (O_342,N_3320,N_4542);
nand UO_343 (O_343,N_2820,N_2695);
or UO_344 (O_344,N_3233,N_3740);
and UO_345 (O_345,N_3927,N_2585);
or UO_346 (O_346,N_4268,N_3957);
or UO_347 (O_347,N_2560,N_3873);
xnor UO_348 (O_348,N_3326,N_4062);
nor UO_349 (O_349,N_4499,N_2673);
nor UO_350 (O_350,N_4973,N_4102);
or UO_351 (O_351,N_3539,N_3384);
nand UO_352 (O_352,N_4105,N_4187);
or UO_353 (O_353,N_2944,N_3778);
nand UO_354 (O_354,N_4841,N_3629);
nand UO_355 (O_355,N_4589,N_3671);
nor UO_356 (O_356,N_4510,N_4646);
xor UO_357 (O_357,N_2892,N_4868);
nand UO_358 (O_358,N_4257,N_3728);
or UO_359 (O_359,N_4157,N_4792);
or UO_360 (O_360,N_4935,N_3216);
nand UO_361 (O_361,N_2542,N_4200);
and UO_362 (O_362,N_3657,N_3913);
nor UO_363 (O_363,N_4707,N_3382);
nand UO_364 (O_364,N_4599,N_4987);
nor UO_365 (O_365,N_4496,N_3826);
and UO_366 (O_366,N_4896,N_3037);
nor UO_367 (O_367,N_3221,N_4467);
nand UO_368 (O_368,N_3068,N_4621);
or UO_369 (O_369,N_4778,N_3162);
and UO_370 (O_370,N_4188,N_2638);
nand UO_371 (O_371,N_3390,N_4475);
nand UO_372 (O_372,N_3463,N_4369);
and UO_373 (O_373,N_3998,N_3352);
or UO_374 (O_374,N_3721,N_2953);
nor UO_375 (O_375,N_4649,N_3785);
nand UO_376 (O_376,N_4795,N_2655);
nand UO_377 (O_377,N_3678,N_4683);
or UO_378 (O_378,N_2651,N_2575);
and UO_379 (O_379,N_2601,N_4285);
or UO_380 (O_380,N_4607,N_2615);
or UO_381 (O_381,N_3383,N_2531);
xor UO_382 (O_382,N_4602,N_3254);
or UO_383 (O_383,N_2610,N_3237);
and UO_384 (O_384,N_4067,N_4380);
nor UO_385 (O_385,N_2799,N_4960);
and UO_386 (O_386,N_3805,N_3650);
nand UO_387 (O_387,N_4638,N_3631);
nand UO_388 (O_388,N_3886,N_3562);
nand UO_389 (O_389,N_3204,N_4345);
and UO_390 (O_390,N_4723,N_4624);
or UO_391 (O_391,N_3953,N_3409);
nor UO_392 (O_392,N_3443,N_2801);
or UO_393 (O_393,N_3315,N_4254);
nor UO_394 (O_394,N_2949,N_2539);
nor UO_395 (O_395,N_2746,N_2867);
or UO_396 (O_396,N_3551,N_4906);
nand UO_397 (O_397,N_3987,N_4346);
nor UO_398 (O_398,N_3930,N_4364);
nor UO_399 (O_399,N_4027,N_2844);
nor UO_400 (O_400,N_3752,N_4154);
nor UO_401 (O_401,N_2882,N_2683);
or UO_402 (O_402,N_4715,N_3693);
nor UO_403 (O_403,N_4997,N_4123);
nor UO_404 (O_404,N_2883,N_3047);
and UO_405 (O_405,N_4697,N_3517);
or UO_406 (O_406,N_4544,N_3131);
nand UO_407 (O_407,N_4167,N_3340);
nor UO_408 (O_408,N_3097,N_2701);
nor UO_409 (O_409,N_2734,N_2926);
nor UO_410 (O_410,N_4535,N_3605);
nor UO_411 (O_411,N_4536,N_3984);
or UO_412 (O_412,N_3588,N_4827);
nor UO_413 (O_413,N_3516,N_2553);
or UO_414 (O_414,N_3191,N_3830);
nor UO_415 (O_415,N_3247,N_2623);
nand UO_416 (O_416,N_3236,N_4848);
nand UO_417 (O_417,N_3819,N_4025);
and UO_418 (O_418,N_3854,N_3025);
and UO_419 (O_419,N_4316,N_2780);
nand UO_420 (O_420,N_3138,N_4259);
and UO_421 (O_421,N_3098,N_3251);
nor UO_422 (O_422,N_4096,N_4660);
nor UO_423 (O_423,N_4709,N_4920);
or UO_424 (O_424,N_2901,N_4813);
and UO_425 (O_425,N_3292,N_3892);
nand UO_426 (O_426,N_4569,N_2995);
nand UO_427 (O_427,N_4068,N_4579);
or UO_428 (O_428,N_3952,N_2727);
and UO_429 (O_429,N_3428,N_4667);
nand UO_430 (O_430,N_4390,N_4736);
and UO_431 (O_431,N_4344,N_4181);
or UO_432 (O_432,N_4633,N_2529);
nand UO_433 (O_433,N_4818,N_3338);
or UO_434 (O_434,N_3467,N_4203);
nor UO_435 (O_435,N_3106,N_2935);
and UO_436 (O_436,N_3293,N_4790);
nor UO_437 (O_437,N_3883,N_4039);
or UO_438 (O_438,N_3558,N_2983);
and UO_439 (O_439,N_3530,N_4937);
nand UO_440 (O_440,N_3809,N_4326);
nand UO_441 (O_441,N_3453,N_4699);
nor UO_442 (O_442,N_3385,N_3568);
and UO_443 (O_443,N_3571,N_2931);
nand UO_444 (O_444,N_4686,N_4357);
or UO_445 (O_445,N_2939,N_2564);
or UO_446 (O_446,N_3371,N_4386);
and UO_447 (O_447,N_2656,N_4561);
and UO_448 (O_448,N_4086,N_3142);
nor UO_449 (O_449,N_3130,N_4722);
nand UO_450 (O_450,N_3975,N_4045);
and UO_451 (O_451,N_4228,N_2715);
nor UO_452 (O_452,N_4622,N_4941);
nor UO_453 (O_453,N_4822,N_3399);
nor UO_454 (O_454,N_3822,N_2617);
or UO_455 (O_455,N_4440,N_4953);
and UO_456 (O_456,N_4377,N_4961);
nand UO_457 (O_457,N_4410,N_4231);
and UO_458 (O_458,N_4875,N_3685);
or UO_459 (O_459,N_4032,N_2732);
and UO_460 (O_460,N_3304,N_4449);
or UO_461 (O_461,N_3036,N_2533);
and UO_462 (O_462,N_3926,N_2631);
and UO_463 (O_463,N_4010,N_2573);
nand UO_464 (O_464,N_4009,N_4008);
and UO_465 (O_465,N_4796,N_3828);
nor UO_466 (O_466,N_4217,N_4809);
nor UO_467 (O_467,N_2865,N_2905);
nor UO_468 (O_468,N_3749,N_4323);
nand UO_469 (O_469,N_2505,N_4658);
or UO_470 (O_470,N_4057,N_2954);
nor UO_471 (O_471,N_4933,N_3851);
or UO_472 (O_472,N_4184,N_4882);
or UO_473 (O_473,N_4048,N_3281);
and UO_474 (O_474,N_3198,N_4037);
and UO_475 (O_475,N_4330,N_3510);
nor UO_476 (O_476,N_3174,N_3125);
nor UO_477 (O_477,N_2836,N_4799);
and UO_478 (O_478,N_2677,N_2725);
and UO_479 (O_479,N_4208,N_2918);
nor UO_480 (O_480,N_4004,N_3277);
and UO_481 (O_481,N_2765,N_4991);
nor UO_482 (O_482,N_4444,N_4745);
or UO_483 (O_483,N_4076,N_3579);
nor UO_484 (O_484,N_3372,N_2700);
nor UO_485 (O_485,N_3386,N_3768);
and UO_486 (O_486,N_3818,N_4103);
nor UO_487 (O_487,N_3311,N_3129);
and UO_488 (O_488,N_4954,N_3298);
or UO_489 (O_489,N_3239,N_4260);
nand UO_490 (O_490,N_4359,N_3328);
and UO_491 (O_491,N_3003,N_2958);
and UO_492 (O_492,N_3999,N_3349);
nor UO_493 (O_493,N_4026,N_4835);
and UO_494 (O_494,N_3427,N_2595);
or UO_495 (O_495,N_3890,N_4071);
nand UO_496 (O_496,N_3024,N_3038);
and UO_497 (O_497,N_4391,N_4929);
nor UO_498 (O_498,N_2933,N_2544);
and UO_499 (O_499,N_3009,N_3698);
nand UO_500 (O_500,N_2967,N_2972);
nand UO_501 (O_501,N_2635,N_3811);
nand UO_502 (O_502,N_2985,N_4714);
and UO_503 (O_503,N_3084,N_3102);
nand UO_504 (O_504,N_3647,N_3850);
nor UO_505 (O_505,N_3255,N_3995);
or UO_506 (O_506,N_3794,N_3111);
or UO_507 (O_507,N_3302,N_4029);
nand UO_508 (O_508,N_2543,N_3429);
or UO_509 (O_509,N_3730,N_4024);
xor UO_510 (O_510,N_3786,N_4803);
nor UO_511 (O_511,N_3393,N_2645);
nand UO_512 (O_512,N_4903,N_3972);
nor UO_513 (O_513,N_4913,N_3862);
nor UO_514 (O_514,N_3110,N_4904);
nand UO_515 (O_515,N_4147,N_4754);
or UO_516 (O_516,N_2824,N_4817);
nor UO_517 (O_517,N_4283,N_4284);
or UO_518 (O_518,N_2878,N_3566);
and UO_519 (O_519,N_4295,N_4717);
and UO_520 (O_520,N_3181,N_3147);
and UO_521 (O_521,N_3369,N_4177);
and UO_522 (O_522,N_4106,N_3529);
nand UO_523 (O_523,N_2845,N_4548);
nand UO_524 (O_524,N_3214,N_2858);
nand UO_525 (O_525,N_3230,N_3980);
or UO_526 (O_526,N_3525,N_3994);
and UO_527 (O_527,N_2789,N_3790);
nand UO_528 (O_528,N_3918,N_3456);
and UO_529 (O_529,N_2782,N_3777);
or UO_530 (O_530,N_3374,N_4332);
nor UO_531 (O_531,N_4565,N_4861);
xor UO_532 (O_532,N_3078,N_2921);
and UO_533 (O_533,N_3276,N_4269);
and UO_534 (O_534,N_3511,N_4018);
nand UO_535 (O_535,N_2726,N_4072);
nor UO_536 (O_536,N_4877,N_4164);
and UO_537 (O_537,N_4312,N_3912);
or UO_538 (O_538,N_4966,N_4985);
and UO_539 (O_539,N_4562,N_4118);
nor UO_540 (O_540,N_3515,N_4641);
or UO_541 (O_541,N_3780,N_4304);
nor UO_542 (O_542,N_4546,N_4741);
and UO_543 (O_543,N_4291,N_4137);
xor UO_544 (O_544,N_4333,N_4520);
nor UO_545 (O_545,N_3026,N_4484);
nand UO_546 (O_546,N_2753,N_4806);
or UO_547 (O_547,N_4892,N_4307);
nor UO_548 (O_548,N_3774,N_4185);
or UO_549 (O_549,N_3563,N_4075);
nor UO_550 (O_550,N_2504,N_3400);
nand UO_551 (O_551,N_3827,N_4674);
and UO_552 (O_552,N_3356,N_4393);
nand UO_553 (O_553,N_3075,N_4629);
and UO_554 (O_554,N_4854,N_3723);
nand UO_555 (O_555,N_4767,N_2913);
or UO_556 (O_556,N_4399,N_3775);
or UO_557 (O_557,N_2800,N_2899);
or UO_558 (O_558,N_3264,N_3874);
or UO_559 (O_559,N_4998,N_2888);
and UO_560 (O_560,N_3305,N_3707);
nor UO_561 (O_561,N_4372,N_3763);
nand UO_562 (O_562,N_3055,N_4964);
nand UO_563 (O_563,N_2509,N_3589);
nor UO_564 (O_564,N_4720,N_2657);
nor UO_565 (O_565,N_4006,N_2637);
or UO_566 (O_566,N_3914,N_3594);
nor UO_567 (O_567,N_3793,N_3424);
and UO_568 (O_568,N_3452,N_3030);
and UO_569 (O_569,N_4816,N_2749);
nor UO_570 (O_570,N_2600,N_3133);
or UO_571 (O_571,N_3042,N_3242);
nand UO_572 (O_572,N_3907,N_4524);
or UO_573 (O_573,N_4839,N_4866);
or UO_574 (O_574,N_4363,N_2748);
nand UO_575 (O_575,N_2784,N_4763);
and UO_576 (O_576,N_4829,N_4685);
nand UO_577 (O_577,N_4598,N_3503);
nand UO_578 (O_578,N_2772,N_3238);
nor UO_579 (O_579,N_4526,N_3480);
or UO_580 (O_580,N_4063,N_4014);
or UO_581 (O_581,N_3432,N_4865);
nor UO_582 (O_582,N_4768,N_3389);
and UO_583 (O_583,N_4400,N_3808);
xnor UO_584 (O_584,N_3100,N_3076);
nand UO_585 (O_585,N_3683,N_2842);
or UO_586 (O_586,N_3234,N_3679);
or UO_587 (O_587,N_3331,N_2866);
and UO_588 (O_588,N_4883,N_4459);
nand UO_589 (O_589,N_4631,N_3823);
or UO_590 (O_590,N_3996,N_3282);
nand UO_591 (O_591,N_4872,N_2957);
nand UO_592 (O_592,N_4577,N_2742);
nand UO_593 (O_593,N_4464,N_4162);
and UO_594 (O_594,N_3116,N_2900);
or UO_595 (O_595,N_4115,N_3477);
xor UO_596 (O_596,N_4356,N_4093);
and UO_597 (O_597,N_4894,N_2694);
nor UO_598 (O_598,N_4489,N_4403);
xor UO_599 (O_599,N_3065,N_3017);
nand UO_600 (O_600,N_2674,N_3486);
nand UO_601 (O_601,N_3611,N_2750);
nand UO_602 (O_602,N_4139,N_3773);
or UO_603 (O_603,N_3825,N_4015);
or UO_604 (O_604,N_2511,N_4021);
xor UO_605 (O_605,N_4341,N_4431);
nor UO_606 (O_606,N_3682,N_2690);
or UO_607 (O_607,N_4863,N_4764);
nor UO_608 (O_608,N_3546,N_3070);
nor UO_609 (O_609,N_4477,N_2829);
nor UO_610 (O_610,N_3018,N_3115);
nor UO_611 (O_611,N_4224,N_4458);
nand UO_612 (O_612,N_3401,N_2973);
nand UO_613 (O_613,N_2624,N_3050);
nand UO_614 (O_614,N_2670,N_4211);
nor UO_615 (O_615,N_4478,N_3857);
xor UO_616 (O_616,N_4820,N_2827);
nand UO_617 (O_617,N_3464,N_3591);
nand UO_618 (O_618,N_4342,N_3922);
nand UO_619 (O_619,N_3064,N_4186);
and UO_620 (O_620,N_3274,N_2863);
nand UO_621 (O_621,N_4744,N_4807);
nor UO_622 (O_622,N_2647,N_2633);
nand UO_623 (O_623,N_4131,N_3540);
nor UO_624 (O_624,N_4879,N_3188);
nor UO_625 (O_625,N_4427,N_2590);
or UO_626 (O_626,N_2786,N_4787);
and UO_627 (O_627,N_4899,N_4967);
or UO_628 (O_628,N_4773,N_3283);
and UO_629 (O_629,N_4468,N_4938);
and UO_630 (O_630,N_3946,N_3246);
or UO_631 (O_631,N_3756,N_3526);
or UO_632 (O_632,N_4445,N_3552);
nor UO_633 (O_633,N_2554,N_3670);
and UO_634 (O_634,N_4553,N_4794);
nor UO_635 (O_635,N_3474,N_4205);
and UO_636 (O_636,N_4669,N_3363);
and UO_637 (O_637,N_4337,N_4958);
or UO_638 (O_638,N_3478,N_4665);
or UO_639 (O_639,N_2632,N_2528);
nor UO_640 (O_640,N_3258,N_4463);
and UO_641 (O_641,N_3322,N_4672);
and UO_642 (O_642,N_3329,N_3833);
nor UO_643 (O_643,N_4756,N_3455);
or UO_644 (O_644,N_2930,N_4506);
or UO_645 (O_645,N_2868,N_4521);
and UO_646 (O_646,N_4197,N_3906);
and UO_647 (O_647,N_2907,N_3405);
and UO_648 (O_648,N_3332,N_3702);
and UO_649 (O_649,N_4210,N_3916);
nor UO_650 (O_650,N_4666,N_3536);
nor UO_651 (O_651,N_4608,N_2838);
or UO_652 (O_652,N_4049,N_2877);
or UO_653 (O_653,N_4718,N_3487);
and UO_654 (O_654,N_4007,N_3439);
or UO_655 (O_655,N_4503,N_4971);
nor UO_656 (O_656,N_3653,N_4272);
nor UO_657 (O_657,N_3706,N_3434);
nand UO_658 (O_658,N_4158,N_4528);
and UO_659 (O_659,N_4358,N_4625);
nor UO_660 (O_660,N_2565,N_2603);
nor UO_661 (O_661,N_3655,N_4974);
nor UO_662 (O_662,N_4760,N_3876);
or UO_663 (O_663,N_4907,N_2840);
nor UO_664 (O_664,N_3080,N_3441);
or UO_665 (O_665,N_2870,N_3507);
nand UO_666 (O_666,N_3903,N_4749);
or UO_667 (O_667,N_4001,N_2909);
nand UO_668 (O_668,N_4193,N_2787);
nor UO_669 (O_669,N_2522,N_4183);
and UO_670 (O_670,N_2506,N_3534);
nor UO_671 (O_671,N_3722,N_4349);
and UO_672 (O_672,N_3508,N_4811);
nor UO_673 (O_673,N_2830,N_2779);
and UO_674 (O_674,N_4766,N_3128);
nand UO_675 (O_675,N_4519,N_3071);
nor UO_676 (O_676,N_4336,N_4080);
nor UO_677 (O_677,N_4266,N_3687);
nor UO_678 (O_678,N_3144,N_3703);
and UO_679 (O_679,N_3132,N_4381);
nand UO_680 (O_680,N_4448,N_4552);
or UO_681 (O_681,N_3844,N_4178);
nor UO_682 (O_682,N_4918,N_4962);
and UO_683 (O_683,N_4677,N_3074);
or UO_684 (O_684,N_3567,N_2775);
and UO_685 (O_685,N_3895,N_3599);
or UO_686 (O_686,N_3992,N_3968);
or UO_687 (O_687,N_2568,N_4945);
or UO_688 (O_688,N_4421,N_3734);
nor UO_689 (O_689,N_4512,N_3632);
or UO_690 (O_690,N_4864,N_4166);
nand UO_691 (O_691,N_4695,N_4549);
and UO_692 (O_692,N_3324,N_4126);
nor UO_693 (O_693,N_3495,N_4784);
nor UO_694 (O_694,N_3299,N_4145);
nor UO_695 (O_695,N_4729,N_4485);
and UO_696 (O_696,N_4583,N_2503);
and UO_697 (O_697,N_2781,N_4361);
or UO_698 (O_698,N_3289,N_4052);
and UO_699 (O_699,N_3598,N_4800);
and UO_700 (O_700,N_2964,N_4825);
nor UO_701 (O_701,N_3553,N_4604);
and UO_702 (O_702,N_3559,N_4651);
nor UO_703 (O_703,N_4640,N_3414);
and UO_704 (O_704,N_2704,N_2965);
nand UO_705 (O_705,N_2639,N_2559);
and UO_706 (O_706,N_4999,N_4701);
nor UO_707 (O_707,N_4314,N_2998);
or UO_708 (O_708,N_4245,N_3011);
and UO_709 (O_709,N_3346,N_3719);
nand UO_710 (O_710,N_3841,N_4908);
nor UO_711 (O_711,N_2587,N_4438);
nand UO_712 (O_712,N_4437,N_2755);
or UO_713 (O_713,N_4910,N_3010);
and UO_714 (O_714,N_3610,N_4852);
or UO_715 (O_715,N_2989,N_3779);
and UO_716 (O_716,N_4732,N_2689);
nor UO_717 (O_717,N_4350,N_3445);
or UO_718 (O_718,N_4543,N_4174);
nand UO_719 (O_719,N_2722,N_3095);
or UO_720 (O_720,N_3590,N_3210);
or UO_721 (O_721,N_4843,N_4241);
nand UO_722 (O_722,N_3148,N_2525);
and UO_723 (O_723,N_2763,N_3974);
or UO_724 (O_724,N_4405,N_4924);
and UO_725 (O_725,N_3989,N_3724);
and UO_726 (O_726,N_3931,N_2984);
nand UO_727 (O_727,N_3869,N_2757);
nand UO_728 (O_728,N_3911,N_2852);
nor UO_729 (O_729,N_4661,N_4914);
nor UO_730 (O_730,N_3437,N_3704);
or UO_731 (O_731,N_3832,N_4327);
or UO_732 (O_732,N_4371,N_4522);
nand UO_733 (O_733,N_3061,N_4585);
and UO_734 (O_734,N_2825,N_4696);
and UO_735 (O_735,N_2709,N_3152);
and UO_736 (O_736,N_4134,N_3582);
and UO_737 (O_737,N_4905,N_4748);
nand UO_738 (O_738,N_2756,N_2552);
and UO_739 (O_739,N_4213,N_4313);
and UO_740 (O_740,N_3353,N_3963);
and UO_741 (O_741,N_3759,N_4765);
nor UO_742 (O_742,N_3705,N_4554);
and UO_743 (O_743,N_3641,N_3905);
nand UO_744 (O_744,N_2915,N_3054);
and UO_745 (O_745,N_4735,N_4855);
nand UO_746 (O_746,N_3748,N_3297);
and UO_747 (O_747,N_2969,N_3831);
nand UO_748 (O_748,N_3330,N_3760);
nand UO_749 (O_749,N_4965,N_3357);
and UO_750 (O_750,N_3410,N_2945);
nand UO_751 (O_751,N_4456,N_4738);
nor UO_752 (O_752,N_3212,N_4867);
and UO_753 (O_753,N_4442,N_3738);
and UO_754 (O_754,N_3440,N_3739);
nor UO_755 (O_755,N_3468,N_3066);
or UO_756 (O_756,N_4791,N_3033);
nand UO_757 (O_757,N_2992,N_4249);
or UO_758 (O_758,N_3135,N_4643);
nand UO_759 (O_759,N_4832,N_4432);
nor UO_760 (O_760,N_4310,N_2986);
nor UO_761 (O_761,N_4383,N_4885);
nand UO_762 (O_762,N_4664,N_4087);
and UO_763 (O_763,N_3395,N_4311);
or UO_764 (O_764,N_4452,N_4481);
nand UO_765 (O_765,N_4338,N_3225);
or UO_766 (O_766,N_3755,N_3421);
nor UO_767 (O_767,N_4277,N_4901);
nor UO_768 (O_768,N_4601,N_4279);
or UO_769 (O_769,N_4705,N_4135);
or UO_770 (O_770,N_3686,N_4671);
nor UO_771 (O_771,N_3285,N_4455);
nand UO_772 (O_772,N_4679,N_4779);
or UO_773 (O_773,N_3224,N_4318);
nand UO_774 (O_774,N_3201,N_3364);
nand UO_775 (O_775,N_2629,N_3574);
and UO_776 (O_776,N_3547,N_4149);
and UO_777 (O_777,N_4850,N_2663);
nor UO_778 (O_778,N_4682,N_3545);
nor UO_779 (O_779,N_4663,N_2500);
nand UO_780 (O_780,N_2771,N_4747);
and UO_781 (O_781,N_3947,N_3502);
nor UO_782 (O_782,N_2879,N_3531);
and UO_783 (O_783,N_3958,N_3935);
nand UO_784 (O_784,N_3252,N_2537);
nand UO_785 (O_785,N_3060,N_2980);
and UO_786 (O_786,N_2682,N_4474);
nand UO_787 (O_787,N_3104,N_2571);
and UO_788 (O_788,N_2814,N_3939);
or UO_789 (O_789,N_2849,N_4130);
nor UO_790 (O_790,N_3419,N_3542);
and UO_791 (O_791,N_3085,N_4838);
or UO_792 (O_792,N_2580,N_3560);
nor UO_793 (O_793,N_4576,N_4159);
nor UO_794 (O_794,N_3185,N_4630);
nor UO_795 (O_795,N_3392,N_4308);
or UO_796 (O_796,N_4216,N_4302);
or UO_797 (O_797,N_4376,N_4170);
nand UO_798 (O_798,N_3099,N_4491);
nand UO_799 (O_799,N_4243,N_2654);
nor UO_800 (O_800,N_4673,N_4873);
or UO_801 (O_801,N_2861,N_2546);
nand UO_802 (O_802,N_2547,N_4834);
nor UO_803 (O_803,N_4917,N_3041);
nand UO_804 (O_804,N_3449,N_4030);
xnor UO_805 (O_805,N_3884,N_3323);
and UO_806 (O_806,N_2816,N_3373);
or UO_807 (O_807,N_3887,N_3284);
or UO_808 (O_808,N_3966,N_3458);
nor UO_809 (O_809,N_4531,N_4398);
or UO_810 (O_810,N_2791,N_3842);
and UO_811 (O_811,N_4762,N_4676);
nor UO_812 (O_812,N_3325,N_2730);
and UO_813 (O_813,N_2582,N_3727);
and UO_814 (O_814,N_4402,N_2846);
and UO_815 (O_815,N_3967,N_4235);
or UO_816 (O_816,N_3928,N_3524);
nand UO_817 (O_817,N_3039,N_2777);
or UO_818 (O_818,N_3094,N_3915);
and UO_819 (O_819,N_4568,N_4733);
nor UO_820 (O_820,N_3925,N_3408);
nor UO_821 (O_821,N_3235,N_2943);
and UO_822 (O_822,N_4734,N_3327);
nand UO_823 (O_823,N_3169,N_3088);
and UO_824 (O_824,N_2859,N_3725);
or UO_825 (O_825,N_4073,N_3634);
and UO_826 (O_826,N_4415,N_4595);
and UO_827 (O_827,N_4500,N_4828);
or UO_828 (O_828,N_2669,N_3901);
xnor UO_829 (O_829,N_3160,N_3354);
nor UO_830 (O_830,N_4339,N_4306);
and UO_831 (O_831,N_4116,N_4692);
nor UO_832 (O_832,N_2612,N_2548);
and UO_833 (O_833,N_4297,N_4274);
nor UO_834 (O_834,N_4808,N_4242);
nor UO_835 (O_835,N_4771,N_4420);
and UO_836 (O_836,N_4690,N_2961);
nor UO_837 (O_837,N_4382,N_2563);
nor UO_838 (O_838,N_3956,N_2841);
nor UO_839 (O_839,N_2735,N_3262);
nand UO_840 (O_840,N_3659,N_2652);
or UO_841 (O_841,N_4698,N_2802);
nand UO_842 (O_842,N_3810,N_4233);
nor UO_843 (O_843,N_4082,N_3709);
nor UO_844 (O_844,N_4949,N_3924);
nand UO_845 (O_845,N_4513,N_3402);
and UO_846 (O_846,N_4278,N_3381);
or UO_847 (O_847,N_4461,N_3199);
and UO_848 (O_848,N_4246,N_2650);
nand UO_849 (O_849,N_3267,N_4525);
nor UO_850 (O_850,N_4810,N_4407);
and UO_851 (O_851,N_2826,N_3028);
or UO_852 (O_852,N_4826,N_4397);
nand UO_853 (O_853,N_4691,N_3417);
or UO_854 (O_854,N_4160,N_4435);
and UO_855 (O_855,N_4483,N_2803);
nor UO_856 (O_856,N_2975,N_4454);
and UO_857 (O_857,N_4776,N_4653);
or UO_858 (O_858,N_3146,N_3415);
nor UO_859 (O_859,N_3348,N_4724);
or UO_860 (O_860,N_3451,N_4541);
and UO_861 (O_861,N_3713,N_3398);
or UO_862 (O_862,N_4560,N_3177);
nor UO_863 (O_863,N_2642,N_4244);
nor UO_864 (O_864,N_2519,N_4353);
and UO_865 (O_865,N_4176,N_2640);
or UO_866 (O_866,N_3342,N_3990);
or UO_867 (O_867,N_4005,N_4480);
and UO_868 (O_868,N_2928,N_4955);
or UO_869 (O_869,N_3273,N_3316);
nand UO_870 (O_870,N_3228,N_3266);
and UO_871 (O_871,N_3014,N_4670);
nand UO_872 (O_872,N_4789,N_3620);
nor UO_873 (O_873,N_3964,N_3868);
nor UO_874 (O_874,N_2869,N_3431);
and UO_875 (O_875,N_4122,N_4551);
nor UO_876 (O_876,N_3838,N_2574);
and UO_877 (O_877,N_3919,N_3249);
and UO_878 (O_878,N_4727,N_4220);
or UO_879 (O_879,N_2959,N_3005);
nand UO_880 (O_880,N_3664,N_2614);
and UO_881 (O_881,N_2987,N_2591);
or UO_882 (O_882,N_2680,N_2724);
nand UO_883 (O_883,N_3767,N_3114);
and UO_884 (O_884,N_3587,N_2770);
nand UO_885 (O_885,N_4540,N_3195);
nand UO_886 (O_886,N_2621,N_3877);
nand UO_887 (O_887,N_4054,N_4120);
nand UO_888 (O_888,N_3900,N_2923);
nor UO_889 (O_889,N_4884,N_3108);
nand UO_890 (O_890,N_4462,N_2720);
nor UO_891 (O_891,N_4331,N_3904);
nand UO_892 (O_892,N_4409,N_4056);
nand UO_893 (O_893,N_3572,N_2993);
or UO_894 (O_894,N_2862,N_4430);
or UO_895 (O_895,N_3885,N_3556);
or UO_896 (O_896,N_4769,N_4859);
and UO_897 (O_897,N_4227,N_3027);
or UO_898 (O_898,N_3413,N_2660);
nand UO_899 (O_899,N_3976,N_3462);
nand UO_900 (O_900,N_3896,N_4151);
or UO_901 (O_901,N_3651,N_3680);
and UO_902 (O_902,N_4922,N_4636);
nand UO_903 (O_903,N_2792,N_2906);
and UO_904 (O_904,N_4328,N_4655);
and UO_905 (O_905,N_4469,N_3929);
and UO_906 (O_906,N_4819,N_3404);
nand UO_907 (O_907,N_3012,N_3804);
or UO_908 (O_908,N_2675,N_4611);
nand UO_909 (O_909,N_4909,N_3355);
or UO_910 (O_910,N_4831,N_4317);
nor UO_911 (O_911,N_4206,N_2815);
nor UO_912 (O_912,N_2551,N_4212);
nand UO_913 (O_913,N_2705,N_4366);
and UO_914 (O_914,N_4742,N_3345);
or UO_915 (O_915,N_4290,N_3677);
nor UO_916 (O_916,N_3815,N_3626);
nor UO_917 (O_917,N_4886,N_4900);
nand UO_918 (O_918,N_3648,N_3934);
and UO_919 (O_919,N_2854,N_3113);
and UO_920 (O_920,N_4514,N_3222);
or UO_921 (O_921,N_4928,N_3004);
nand UO_922 (O_922,N_2806,N_3981);
and UO_923 (O_923,N_3908,N_4419);
nor UO_924 (O_924,N_4168,N_4095);
and UO_925 (O_925,N_2549,N_4950);
nand UO_926 (O_926,N_3820,N_3875);
nor UO_927 (O_927,N_2572,N_3172);
or UO_928 (O_928,N_3584,N_4956);
and UO_929 (O_929,N_4815,N_3447);
and UO_930 (O_930,N_2681,N_4979);
nand UO_931 (O_931,N_3592,N_2649);
nand UO_932 (O_932,N_2570,N_4424);
nand UO_933 (O_933,N_4889,N_4113);
nand UO_934 (O_934,N_2662,N_3533);
nor UO_935 (O_935,N_4065,N_3021);
or UO_936 (O_936,N_3936,N_3538);
or UO_937 (O_937,N_2754,N_4824);
or UO_938 (O_938,N_3466,N_3139);
nand UO_939 (O_939,N_3577,N_4195);
nor UO_940 (O_940,N_4090,N_2908);
or UO_941 (O_941,N_4793,N_2890);
or UO_942 (O_942,N_4755,N_2516);
nor UO_943 (O_943,N_4523,N_4504);
or UO_944 (O_944,N_2855,N_2962);
nand UO_945 (O_945,N_3499,N_3063);
and UO_946 (O_946,N_4880,N_2788);
and UO_947 (O_947,N_4408,N_3660);
nor UO_948 (O_948,N_3729,N_3726);
nor UO_949 (O_949,N_3518,N_3436);
and UO_950 (O_950,N_3845,N_3301);
or UO_951 (O_951,N_4280,N_4240);
nor UO_952 (O_952,N_4219,N_4189);
or UO_953 (O_953,N_4276,N_2876);
nand UO_954 (O_954,N_3643,N_4786);
and UO_955 (O_955,N_4324,N_3370);
nor UO_956 (O_956,N_4443,N_4871);
and UO_957 (O_957,N_3377,N_4055);
nand UO_958 (O_958,N_4031,N_3803);
nor UO_959 (O_959,N_4702,N_4426);
or UO_960 (O_960,N_3179,N_2527);
or UO_961 (O_961,N_4258,N_3891);
nor UO_962 (O_962,N_4593,N_3696);
nor UO_963 (O_963,N_4635,N_3796);
nand UO_964 (O_964,N_4657,N_3663);
nor UO_965 (O_965,N_3126,N_4271);
or UO_966 (O_966,N_3712,N_3425);
or UO_967 (O_967,N_2625,N_4592);
and UO_968 (O_968,N_4556,N_3746);
nand UO_969 (O_969,N_3375,N_4610);
or UO_970 (O_970,N_2744,N_4812);
and UO_971 (O_971,N_2581,N_2904);
or UO_972 (O_972,N_4089,N_4804);
and UO_973 (O_973,N_4289,N_3321);
or UO_974 (O_974,N_3171,N_4678);
nand UO_975 (O_975,N_2833,N_4612);
nand UO_976 (O_976,N_4947,N_2684);
or UO_977 (O_977,N_2627,N_4051);
and UO_978 (O_978,N_2736,N_4746);
nor UO_979 (O_979,N_4414,N_2873);
and UO_980 (O_980,N_3433,N_3878);
and UO_981 (O_981,N_2956,N_2880);
nand UO_982 (O_982,N_2583,N_2895);
or UO_983 (O_983,N_2941,N_3812);
nand UO_984 (O_984,N_4995,N_4144);
nand UO_985 (O_985,N_2805,N_4305);
xor UO_986 (O_986,N_4132,N_4573);
or UO_987 (O_987,N_3493,N_4081);
nand UO_988 (O_988,N_3362,N_2981);
nor UO_989 (O_989,N_3565,N_4925);
nand UO_990 (O_990,N_4969,N_3492);
and UO_991 (O_991,N_3155,N_2874);
and UO_992 (O_992,N_3772,N_4204);
nor UO_993 (O_993,N_3140,N_4992);
nor UO_994 (O_994,N_3882,N_3621);
or UO_995 (O_995,N_3069,N_4845);
nor UO_996 (O_996,N_4201,N_2804);
nand UO_997 (O_997,N_4853,N_4182);
and UO_998 (O_998,N_3073,N_4412);
nand UO_999 (O_999,N_4384,N_4634);
endmodule