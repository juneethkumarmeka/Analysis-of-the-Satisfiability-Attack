module basic_1500_15000_2000_3_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10002,N_10004,N_10005,N_10006,N_10007,N_10008,N_10010,N_10011,N_10012,N_10014,N_10015,N_10016,N_10017,N_10019,N_10020,N_10021,N_10022,N_10024,N_10026,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10062,N_10063,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10074,N_10076,N_10078,N_10080,N_10082,N_10084,N_10085,N_10086,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10095,N_10096,N_10097,N_10098,N_10099,N_10101,N_10103,N_10107,N_10108,N_10109,N_10110,N_10111,N_10113,N_10116,N_10117,N_10118,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10129,N_10131,N_10132,N_10133,N_10134,N_10136,N_10137,N_10138,N_10139,N_10140,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10152,N_10153,N_10154,N_10155,N_10157,N_10159,N_10160,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10199,N_10200,N_10202,N_10203,N_10205,N_10208,N_10209,N_10210,N_10211,N_10212,N_10214,N_10215,N_10217,N_10218,N_10219,N_10220,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10243,N_10244,N_10248,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10279,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10308,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10319,N_10320,N_10321,N_10322,N_10324,N_10326,N_10327,N_10328,N_10330,N_10331,N_10332,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10354,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10365,N_10367,N_10368,N_10369,N_10370,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10416,N_10417,N_10418,N_10419,N_10420,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10446,N_10447,N_10448,N_10449,N_10450,N_10452,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10480,N_10482,N_10483,N_10485,N_10488,N_10490,N_10491,N_10492,N_10493,N_10494,N_10496,N_10498,N_10499,N_10500,N_10501,N_10503,N_10504,N_10505,N_10507,N_10508,N_10509,N_10510,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10523,N_10524,N_10526,N_10527,N_10528,N_10529,N_10531,N_10532,N_10533,N_10535,N_10536,N_10537,N_10538,N_10540,N_10541,N_10543,N_10546,N_10547,N_10548,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10563,N_10564,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10578,N_10579,N_10580,N_10581,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10625,N_10626,N_10627,N_10629,N_10630,N_10631,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10649,N_10651,N_10652,N_10653,N_10654,N_10655,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10670,N_10671,N_10672,N_10674,N_10675,N_10677,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10698,N_10699,N_10700,N_10701,N_10702,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10721,N_10722,N_10723,N_10724,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10750,N_10751,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10760,N_10761,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10771,N_10772,N_10773,N_10777,N_10778,N_10780,N_10781,N_10782,N_10783,N_10785,N_10786,N_10787,N_10788,N_10789,N_10791,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10800,N_10801,N_10802,N_10803,N_10804,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10826,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10838,N_10839,N_10841,N_10842,N_10844,N_10846,N_10848,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10875,N_10876,N_10877,N_10878,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10891,N_10892,N_10893,N_10894,N_10895,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10925,N_10927,N_10928,N_10930,N_10932,N_10934,N_10935,N_10936,N_10938,N_10939,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10952,N_10953,N_10954,N_10955,N_10956,N_10958,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10969,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10985,N_10986,N_10987,N_10988,N_10989,N_10991,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_11000,N_11001,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11012,N_11015,N_11016,N_11017,N_11018,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11032,N_11033,N_11034,N_11036,N_11037,N_11038,N_11039,N_11040,N_11042,N_11043,N_11044,N_11045,N_11047,N_11049,N_11050,N_11051,N_11052,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11061,N_11062,N_11064,N_11065,N_11066,N_11067,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11077,N_11078,N_11079,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11095,N_11096,N_11097,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11112,N_11113,N_11114,N_11115,N_11116,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11150,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11164,N_11165,N_11167,N_11168,N_11170,N_11171,N_11172,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11186,N_11188,N_11189,N_11190,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11210,N_11211,N_11213,N_11214,N_11215,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11228,N_11229,N_11230,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11247,N_11248,N_11249,N_11250,N_11251,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11266,N_11268,N_11269,N_11270,N_11273,N_11275,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11302,N_11303,N_11304,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11318,N_11319,N_11320,N_11321,N_11323,N_11324,N_11325,N_11326,N_11328,N_11329,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11380,N_11381,N_11382,N_11384,N_11385,N_11386,N_11387,N_11388,N_11392,N_11393,N_11394,N_11395,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11405,N_11406,N_11408,N_11410,N_11412,N_11415,N_11416,N_11417,N_11418,N_11419,N_11421,N_11422,N_11425,N_11426,N_11427,N_11428,N_11430,N_11431,N_11432,N_11433,N_11434,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11469,N_11472,N_11473,N_11474,N_11475,N_11476,N_11479,N_11480,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11492,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11502,N_11503,N_11504,N_11505,N_11506,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11542,N_11543,N_11544,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11573,N_11574,N_11576,N_11577,N_11578,N_11581,N_11582,N_11584,N_11586,N_11587,N_11588,N_11589,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11600,N_11601,N_11602,N_11604,N_11606,N_11607,N_11608,N_11609,N_11610,N_11612,N_11613,N_11614,N_11615,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11633,N_11634,N_11635,N_11636,N_11637,N_11640,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11662,N_11663,N_11665,N_11666,N_11667,N_11669,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11692,N_11694,N_11697,N_11698,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11713,N_11714,N_11715,N_11716,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11725,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11734,N_11735,N_11736,N_11737,N_11738,N_11741,N_11742,N_11743,N_11745,N_11746,N_11748,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11759,N_11761,N_11763,N_11764,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11776,N_11777,N_11780,N_11782,N_11783,N_11784,N_11785,N_11787,N_11788,N_11790,N_11791,N_11793,N_11794,N_11796,N_11798,N_11799,N_11800,N_11801,N_11803,N_11804,N_11805,N_11807,N_11808,N_11810,N_11811,N_11812,N_11814,N_11815,N_11817,N_11818,N_11819,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11829,N_11830,N_11831,N_11833,N_11834,N_11835,N_11836,N_11837,N_11839,N_11841,N_11844,N_11845,N_11846,N_11849,N_11850,N_11851,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11873,N_11874,N_11875,N_11877,N_11880,N_11882,N_11883,N_11884,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11895,N_11896,N_11898,N_11899,N_11900,N_11902,N_11903,N_11904,N_11906,N_11908,N_11909,N_11910,N_11911,N_11912,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11951,N_11952,N_11953,N_11955,N_11956,N_11958,N_11960,N_11961,N_11962,N_11963,N_11965,N_11967,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11984,N_11985,N_11986,N_11987,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12010,N_12011,N_12013,N_12014,N_12015,N_12017,N_12018,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12046,N_12048,N_12049,N_12050,N_12051,N_12052,N_12054,N_12056,N_12058,N_12059,N_12060,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12077,N_12078,N_12079,N_12080,N_12082,N_12083,N_12085,N_12087,N_12088,N_12089,N_12090,N_12092,N_12093,N_12094,N_12096,N_12097,N_12099,N_12100,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12110,N_12112,N_12114,N_12115,N_12116,N_12118,N_12119,N_12121,N_12123,N_12125,N_12126,N_12128,N_12130,N_12132,N_12133,N_12134,N_12135,N_12137,N_12138,N_12139,N_12140,N_12141,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12154,N_12155,N_12156,N_12157,N_12158,N_12160,N_12161,N_12163,N_12164,N_12165,N_12166,N_12167,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12183,N_12184,N_12186,N_12187,N_12188,N_12189,N_12191,N_12192,N_12193,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12203,N_12204,N_12205,N_12207,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12218,N_12219,N_12220,N_12221,N_12223,N_12225,N_12227,N_12228,N_12229,N_12230,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12246,N_12247,N_12248,N_12249,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12264,N_12265,N_12267,N_12269,N_12270,N_12271,N_12272,N_12274,N_12275,N_12276,N_12278,N_12279,N_12280,N_12281,N_12285,N_12286,N_12287,N_12288,N_12289,N_12291,N_12292,N_12293,N_12294,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12303,N_12304,N_12305,N_12306,N_12308,N_12309,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12321,N_12322,N_12323,N_12324,N_12325,N_12327,N_12328,N_12329,N_12330,N_12332,N_12333,N_12334,N_12335,N_12336,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12372,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12382,N_12385,N_12386,N_12389,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12412,N_12413,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12432,N_12433,N_12434,N_12435,N_12436,N_12440,N_12441,N_12442,N_12443,N_12444,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12464,N_12465,N_12467,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12479,N_12480,N_12481,N_12482,N_12483,N_12485,N_12486,N_12487,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12548,N_12549,N_12550,N_12552,N_12553,N_12554,N_12555,N_12556,N_12558,N_12560,N_12561,N_12562,N_12564,N_12565,N_12566,N_12567,N_12569,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12593,N_12594,N_12595,N_12596,N_12597,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12626,N_12627,N_12632,N_12634,N_12635,N_12638,N_12639,N_12640,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12650,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12660,N_12661,N_12662,N_12663,N_12664,N_12667,N_12669,N_12670,N_12671,N_12673,N_12674,N_12676,N_12679,N_12680,N_12681,N_12683,N_12684,N_12685,N_12686,N_12687,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12716,N_12717,N_12718,N_12719,N_12721,N_12722,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12740,N_12741,N_12742,N_12743,N_12744,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12760,N_12761,N_12762,N_12764,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12779,N_12780,N_12781,N_12782,N_12784,N_12785,N_12787,N_12788,N_12790,N_12793,N_12794,N_12795,N_12796,N_12797,N_12799,N_12800,N_12801,N_12804,N_12805,N_12806,N_12807,N_12809,N_12810,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12823,N_12824,N_12826,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12865,N_12866,N_12867,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12885,N_12886,N_12887,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12907,N_12909,N_12910,N_12912,N_12913,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12928,N_12929,N_12930,N_12932,N_12933,N_12934,N_12935,N_12936,N_12938,N_12939,N_12940,N_12941,N_12943,N_12944,N_12945,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12962,N_12963,N_12964,N_12965,N_12967,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12981,N_12983,N_12984,N_12985,N_12986,N_12987,N_12989,N_12990,N_12991,N_12994,N_12995,N_12996,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13027,N_13028,N_13030,N_13032,N_13034,N_13035,N_13036,N_13038,N_13040,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13065,N_13066,N_13067,N_13069,N_13070,N_13072,N_13073,N_13075,N_13076,N_13077,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13092,N_13094,N_13095,N_13096,N_13097,N_13099,N_13101,N_13102,N_13104,N_13105,N_13106,N_13108,N_13109,N_13111,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13137,N_13138,N_13140,N_13141,N_13142,N_13143,N_13145,N_13146,N_13147,N_13148,N_13150,N_13151,N_13152,N_13153,N_13155,N_13156,N_13158,N_13160,N_13161,N_13162,N_13164,N_13165,N_13167,N_13168,N_13169,N_13170,N_13171,N_13175,N_13176,N_13177,N_13179,N_13181,N_13182,N_13183,N_13184,N_13186,N_13187,N_13188,N_13189,N_13190,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13227,N_13228,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13237,N_13238,N_13240,N_13241,N_13243,N_13245,N_13246,N_13248,N_13250,N_13251,N_13252,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13262,N_13264,N_13265,N_13266,N_13267,N_13268,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13310,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13319,N_13320,N_13321,N_13322,N_13323,N_13325,N_13326,N_13327,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13339,N_13340,N_13344,N_13345,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13358,N_13359,N_13361,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13374,N_13377,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13390,N_13392,N_13394,N_13395,N_13396,N_13397,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13418,N_13419,N_13420,N_13421,N_13422,N_13424,N_13425,N_13426,N_13429,N_13430,N_13432,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13453,N_13455,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13475,N_13476,N_13477,N_13478,N_13480,N_13481,N_13483,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13512,N_13514,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13538,N_13539,N_13540,N_13541,N_13542,N_13544,N_13545,N_13546,N_13548,N_13549,N_13550,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13560,N_13564,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13577,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13588,N_13589,N_13590,N_13591,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13613,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13634,N_13635,N_13636,N_13637,N_13638,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13647,N_13648,N_13649,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13665,N_13667,N_13668,N_13670,N_13671,N_13672,N_13673,N_13675,N_13676,N_13677,N_13679,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13700,N_13701,N_13702,N_13703,N_13704,N_13706,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13716,N_13717,N_13718,N_13719,N_13720,N_13722,N_13725,N_13726,N_13727,N_13728,N_13730,N_13734,N_13735,N_13736,N_13737,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13768,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13780,N_13781,N_13782,N_13783,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13803,N_13804,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13852,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13888,N_13889,N_13890,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13919,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13951,N_13954,N_13955,N_13956,N_13958,N_13960,N_13962,N_13963,N_13964,N_13965,N_13966,N_13969,N_13971,N_13972,N_13973,N_13974,N_13975,N_13977,N_13978,N_13979,N_13980,N_13981,N_13983,N_13985,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14007,N_14008,N_14009,N_14010,N_14013,N_14014,N_14016,N_14017,N_14018,N_14020,N_14021,N_14022,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14034,N_14035,N_14036,N_14037,N_14038,N_14040,N_14042,N_14043,N_14044,N_14045,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14054,N_14055,N_14057,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14075,N_14076,N_14078,N_14079,N_14080,N_14082,N_14083,N_14085,N_14087,N_14089,N_14090,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14107,N_14109,N_14110,N_14111,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14127,N_14128,N_14129,N_14130,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14145,N_14146,N_14147,N_14148,N_14150,N_14151,N_14152,N_14153,N_14155,N_14156,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14171,N_14173,N_14176,N_14177,N_14178,N_14179,N_14180,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14236,N_14238,N_14239,N_14240,N_14241,N_14243,N_14244,N_14245,N_14247,N_14250,N_14251,N_14253,N_14254,N_14255,N_14256,N_14257,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14289,N_14290,N_14291,N_14292,N_14294,N_14295,N_14297,N_14299,N_14300,N_14301,N_14302,N_14303,N_14305,N_14306,N_14307,N_14309,N_14310,N_14311,N_14313,N_14315,N_14317,N_14318,N_14320,N_14322,N_14323,N_14324,N_14325,N_14326,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14338,N_14339,N_14341,N_14342,N_14343,N_14344,N_14345,N_14347,N_14348,N_14349,N_14350,N_14351,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14393,N_14394,N_14395,N_14398,N_14399,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14412,N_14413,N_14414,N_14415,N_14417,N_14418,N_14420,N_14421,N_14422,N_14423,N_14425,N_14426,N_14427,N_14428,N_14429,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14445,N_14448,N_14450,N_14451,N_14453,N_14454,N_14455,N_14457,N_14458,N_14460,N_14461,N_14462,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14473,N_14474,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14486,N_14487,N_14489,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14512,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14529,N_14530,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14544,N_14545,N_14546,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14566,N_14567,N_14569,N_14570,N_14571,N_14572,N_14573,N_14577,N_14578,N_14579,N_14580,N_14581,N_14583,N_14584,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14598,N_14600,N_14602,N_14603,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14617,N_14618,N_14619,N_14620,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14630,N_14631,N_14632,N_14634,N_14635,N_14636,N_14637,N_14638,N_14640,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14653,N_14654,N_14655,N_14657,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14667,N_14668,N_14672,N_14673,N_14674,N_14675,N_14676,N_14679,N_14680,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14715,N_14716,N_14717,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14734,N_14737,N_14739,N_14740,N_14741,N_14742,N_14743,N_14745,N_14746,N_14747,N_14748,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14761,N_14762,N_14764,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14787,N_14789,N_14790,N_14791,N_14792,N_14793,N_14795,N_14796,N_14797,N_14799,N_14800,N_14801,N_14802,N_14803,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14833,N_14834,N_14835,N_14836,N_14838,N_14839,N_14840,N_14841,N_14842,N_14844,N_14845,N_14846,N_14847,N_14850,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14886,N_14888,N_14891,N_14892,N_14893,N_14894,N_14895,N_14897,N_14898,N_14899,N_14902,N_14904,N_14906,N_14908,N_14909,N_14911,N_14912,N_14913,N_14916,N_14918,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14936,N_14937,N_14938,N_14939,N_14940,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14981,N_14982,N_14985,N_14990,N_14991,N_14993,N_14994,N_14995,N_14998,N_14999;
nor U0 (N_0,In_319,In_235);
xnor U1 (N_1,In_70,In_1267);
nor U2 (N_2,In_173,In_21);
xor U3 (N_3,In_1088,In_841);
or U4 (N_4,In_1085,In_400);
xor U5 (N_5,In_674,In_473);
nand U6 (N_6,In_968,In_1303);
nand U7 (N_7,In_974,In_1290);
xnor U8 (N_8,In_518,In_1104);
xor U9 (N_9,In_859,In_588);
nand U10 (N_10,In_528,In_347);
xnor U11 (N_11,In_356,In_754);
and U12 (N_12,In_1406,In_48);
and U13 (N_13,In_230,In_1336);
nor U14 (N_14,In_836,In_545);
xor U15 (N_15,In_679,In_677);
nor U16 (N_16,In_708,In_1471);
and U17 (N_17,In_690,In_1201);
nand U18 (N_18,In_863,In_165);
and U19 (N_19,In_989,In_307);
nand U20 (N_20,In_902,In_131);
nor U21 (N_21,In_176,In_1443);
and U22 (N_22,In_595,In_412);
and U23 (N_23,In_1316,In_200);
nor U24 (N_24,In_261,In_313);
and U25 (N_25,In_1340,In_1282);
nand U26 (N_26,In_757,In_1241);
xnor U27 (N_27,In_1126,In_1036);
or U28 (N_28,In_954,In_1479);
xor U29 (N_29,In_377,In_629);
xor U30 (N_30,In_1151,In_369);
or U31 (N_31,In_969,In_193);
nor U32 (N_32,In_1347,In_281);
or U33 (N_33,In_431,In_1299);
or U34 (N_34,In_1141,In_189);
xor U35 (N_35,In_1477,In_581);
and U36 (N_36,In_1293,In_882);
xor U37 (N_37,In_361,In_546);
nand U38 (N_38,In_1215,In_920);
xor U39 (N_39,In_0,In_124);
xor U40 (N_40,In_1363,In_496);
nand U41 (N_41,In_117,In_827);
and U42 (N_42,In_1450,In_1481);
nand U43 (N_43,In_443,In_330);
nand U44 (N_44,In_94,In_401);
nor U45 (N_45,In_306,In_1433);
xnor U46 (N_46,In_977,In_320);
xnor U47 (N_47,In_442,In_490);
nand U48 (N_48,In_828,In_459);
nand U49 (N_49,In_271,In_565);
or U50 (N_50,In_272,In_1484);
and U51 (N_51,In_553,In_1352);
nand U52 (N_52,In_354,In_78);
nor U53 (N_53,In_1073,In_418);
nand U54 (N_54,In_1279,In_1135);
and U55 (N_55,In_1378,In_839);
nand U56 (N_56,In_1380,In_1192);
nand U57 (N_57,In_205,In_1211);
xor U58 (N_58,In_793,In_843);
and U59 (N_59,In_423,In_955);
nand U60 (N_60,In_1338,In_4);
nor U61 (N_61,In_577,In_460);
nor U62 (N_62,In_1187,In_917);
or U63 (N_63,In_907,In_915);
and U64 (N_64,In_519,In_684);
nor U65 (N_65,In_860,In_248);
nor U66 (N_66,In_402,In_829);
nor U67 (N_67,In_567,In_975);
or U68 (N_68,In_227,In_709);
nand U69 (N_69,In_1254,In_1233);
xor U70 (N_70,In_409,In_19);
xor U71 (N_71,In_1002,In_339);
xor U72 (N_72,In_1062,In_991);
nand U73 (N_73,In_962,In_1238);
xnor U74 (N_74,In_341,In_717);
nand U75 (N_75,In_1493,In_91);
xor U76 (N_76,In_665,In_300);
xnor U77 (N_77,In_380,In_1425);
and U78 (N_78,In_801,In_1043);
nor U79 (N_79,In_1269,In_864);
nor U80 (N_80,In_374,In_245);
xnor U81 (N_81,In_299,In_1328);
nor U82 (N_82,In_1418,In_468);
and U83 (N_83,In_876,In_1193);
nand U84 (N_84,In_1499,In_1277);
nand U85 (N_85,In_1053,In_18);
nor U86 (N_86,In_635,In_1237);
or U87 (N_87,In_982,In_928);
nor U88 (N_88,In_1167,In_922);
nand U89 (N_89,In_1125,In_1345);
xnor U90 (N_90,In_1495,In_1230);
or U91 (N_91,In_1,In_521);
and U92 (N_92,In_1438,In_384);
and U93 (N_93,In_225,In_119);
xnor U94 (N_94,In_174,In_1330);
nor U95 (N_95,In_956,In_23);
or U96 (N_96,In_47,In_981);
or U97 (N_97,In_650,In_233);
and U98 (N_98,In_1497,In_448);
or U99 (N_99,In_137,In_729);
nand U100 (N_100,In_638,In_344);
nor U101 (N_101,In_666,In_331);
nor U102 (N_102,In_256,In_334);
nor U103 (N_103,In_392,In_396);
nor U104 (N_104,In_772,In_391);
and U105 (N_105,In_501,In_857);
nand U106 (N_106,In_76,In_593);
or U107 (N_107,In_1412,In_549);
and U108 (N_108,In_651,In_1055);
nand U109 (N_109,In_1353,In_1391);
nor U110 (N_110,In_1030,In_868);
xor U111 (N_111,In_726,In_1173);
or U112 (N_112,In_1225,In_206);
and U113 (N_113,In_1474,In_95);
xnor U114 (N_114,In_622,In_1307);
or U115 (N_115,In_1009,In_1091);
and U116 (N_116,In_24,In_122);
nor U117 (N_117,In_965,In_492);
xnor U118 (N_118,In_1323,In_606);
xnor U119 (N_119,In_1019,In_1152);
and U120 (N_120,In_1035,In_121);
or U121 (N_121,In_1457,In_696);
xor U122 (N_122,In_455,In_1161);
nand U123 (N_123,In_536,In_181);
xnor U124 (N_124,In_763,In_1178);
nor U125 (N_125,In_452,In_202);
xnor U126 (N_126,In_834,In_1068);
nor U127 (N_127,In_185,In_1414);
nand U128 (N_128,In_865,In_10);
or U129 (N_129,In_610,In_3);
nand U130 (N_130,In_967,In_364);
nor U131 (N_131,In_215,In_1332);
xnor U132 (N_132,In_1143,In_984);
and U133 (N_133,In_83,In_1075);
and U134 (N_134,In_197,In_1295);
and U135 (N_135,In_596,In_668);
or U136 (N_136,In_1081,In_619);
xnor U137 (N_137,In_736,In_54);
or U138 (N_138,In_279,In_1301);
nor U139 (N_139,In_949,In_1115);
nand U140 (N_140,In_385,In_444);
or U141 (N_141,In_1171,In_680);
or U142 (N_142,In_351,In_25);
nor U143 (N_143,In_923,In_766);
xnor U144 (N_144,In_513,In_109);
nand U145 (N_145,In_632,In_1439);
or U146 (N_146,In_438,In_1118);
or U147 (N_147,In_1024,In_617);
xnor U148 (N_148,In_778,In_760);
or U149 (N_149,In_932,In_951);
or U150 (N_150,In_771,In_976);
xnor U151 (N_151,In_1224,In_601);
and U152 (N_152,In_1058,In_723);
or U153 (N_153,In_647,In_777);
or U154 (N_154,In_735,In_1228);
and U155 (N_155,In_274,In_1221);
or U156 (N_156,In_1177,In_463);
or U157 (N_157,In_1403,In_101);
nor U158 (N_158,In_1146,In_1098);
or U159 (N_159,In_1417,In_850);
nor U160 (N_160,In_81,In_1138);
nor U161 (N_161,In_1287,In_219);
nor U162 (N_162,In_37,In_1016);
nor U163 (N_163,In_1475,In_375);
xor U164 (N_164,In_1008,In_789);
and U165 (N_165,In_184,In_591);
nor U166 (N_166,In_837,In_732);
or U167 (N_167,In_699,In_1342);
nor U168 (N_168,In_942,In_508);
or U169 (N_169,In_335,In_776);
or U170 (N_170,In_1396,In_290);
nor U171 (N_171,In_832,In_1382);
xnor U172 (N_172,In_616,In_345);
nand U173 (N_173,In_1208,In_1090);
xnor U174 (N_174,In_733,In_1061);
xor U175 (N_175,In_929,In_825);
and U176 (N_176,In_390,In_901);
xnor U177 (N_177,In_1229,In_75);
nand U178 (N_178,In_1154,In_426);
nor U179 (N_179,In_544,In_1272);
xnor U180 (N_180,In_627,In_820);
xor U181 (N_181,In_180,In_1358);
nor U182 (N_182,In_1478,In_1446);
or U183 (N_183,In_212,In_770);
or U184 (N_184,In_583,In_569);
and U185 (N_185,In_49,In_887);
or U186 (N_186,In_1262,In_940);
xor U187 (N_187,In_257,In_156);
nand U188 (N_188,In_739,In_166);
nor U189 (N_189,In_744,In_561);
and U190 (N_190,In_1223,In_873);
and U191 (N_191,In_1464,In_1087);
nor U192 (N_192,In_695,In_1372);
or U193 (N_193,In_39,In_31);
nor U194 (N_194,In_346,In_379);
nand U195 (N_195,In_1028,In_1416);
nor U196 (N_196,In_1047,In_861);
nor U197 (N_197,In_862,In_422);
nor U198 (N_198,In_1011,In_767);
nand U199 (N_199,In_782,In_1180);
nor U200 (N_200,In_986,In_1374);
and U201 (N_201,In_148,In_909);
or U202 (N_202,In_1089,In_216);
nand U203 (N_203,In_142,In_1069);
nor U204 (N_204,In_29,In_67);
xor U205 (N_205,In_1367,In_897);
nor U206 (N_206,In_849,In_813);
and U207 (N_207,In_1181,In_1407);
nor U208 (N_208,In_608,In_660);
or U209 (N_209,In_1082,In_872);
or U210 (N_210,In_786,In_764);
xnor U211 (N_211,In_648,In_636);
xnor U212 (N_212,In_1064,In_106);
nand U213 (N_213,In_605,In_1294);
and U214 (N_214,In_11,In_477);
nand U215 (N_215,In_275,In_218);
or U216 (N_216,In_611,In_552);
and U217 (N_217,In_563,In_669);
nand U218 (N_218,In_223,In_160);
nand U219 (N_219,In_103,In_742);
and U220 (N_220,In_1271,In_846);
xnor U221 (N_221,In_139,In_482);
and U222 (N_222,In_558,In_1315);
nand U223 (N_223,In_231,In_727);
xnor U224 (N_224,In_946,In_1071);
nor U225 (N_225,In_875,In_509);
or U226 (N_226,In_1333,In_710);
or U227 (N_227,In_481,In_870);
and U228 (N_228,In_61,In_779);
and U229 (N_229,In_434,In_931);
nand U230 (N_230,In_1067,In_286);
and U231 (N_231,In_102,In_311);
nor U232 (N_232,In_1429,In_111);
nand U233 (N_233,In_971,In_51);
nor U234 (N_234,In_1127,In_298);
or U235 (N_235,In_745,In_582);
or U236 (N_236,In_112,In_430);
or U237 (N_237,In_898,In_46);
xnor U238 (N_238,In_1437,In_99);
nand U239 (N_239,In_945,In_885);
or U240 (N_240,In_1095,In_1051);
nand U241 (N_241,In_1496,In_476);
or U242 (N_242,In_1139,In_1434);
nor U243 (N_243,In_440,In_1106);
nand U244 (N_244,In_291,In_220);
and U245 (N_245,In_1013,In_663);
nand U246 (N_246,In_791,In_1157);
nand U247 (N_247,In_807,In_357);
xor U248 (N_248,In_675,In_654);
nand U249 (N_249,In_310,In_906);
nor U250 (N_250,In_376,In_13);
nor U251 (N_251,In_598,In_316);
or U252 (N_252,In_1029,In_1451);
nor U253 (N_253,In_1317,In_338);
nand U254 (N_254,In_1166,In_108);
or U255 (N_255,In_1476,In_520);
and U256 (N_256,In_485,In_1296);
xor U257 (N_257,In_277,In_82);
and U258 (N_258,In_1054,In_822);
nand U259 (N_259,In_1387,In_524);
or U260 (N_260,In_45,In_217);
nand U261 (N_261,In_833,In_1252);
nor U262 (N_262,In_1298,In_72);
or U263 (N_263,In_891,In_785);
or U264 (N_264,In_851,In_600);
and U265 (N_265,In_979,In_645);
and U266 (N_266,In_73,In_603);
and U267 (N_267,In_312,In_87);
or U268 (N_268,In_28,In_348);
and U269 (N_269,In_1218,In_1274);
xnor U270 (N_270,In_858,In_1093);
and U271 (N_271,In_664,In_493);
or U272 (N_272,In_343,In_1465);
or U273 (N_273,In_133,In_1116);
nor U274 (N_274,In_762,In_1148);
nor U275 (N_275,In_1306,In_1189);
and U276 (N_276,In_394,In_250);
and U277 (N_277,In_360,In_1226);
and U278 (N_278,In_315,In_242);
and U279 (N_279,In_644,In_883);
and U280 (N_280,In_580,In_1400);
and U281 (N_281,In_692,In_98);
xor U282 (N_282,In_1174,In_479);
and U283 (N_283,In_506,In_743);
or U284 (N_284,In_568,In_855);
nand U285 (N_285,In_224,In_251);
xnor U286 (N_286,In_625,In_1292);
nor U287 (N_287,In_751,In_450);
and U288 (N_288,In_824,In_912);
xnor U289 (N_289,In_734,In_1168);
nor U290 (N_290,In_652,In_208);
nand U291 (N_291,In_1351,In_691);
nor U292 (N_292,In_869,In_1249);
nand U293 (N_293,In_337,In_1145);
and U294 (N_294,In_17,In_389);
or U295 (N_295,In_34,In_147);
nor U296 (N_296,In_1248,In_326);
xnor U297 (N_297,In_584,In_781);
nand U298 (N_298,In_1227,In_399);
nand U299 (N_299,In_113,In_1099);
nor U300 (N_300,In_135,In_682);
xor U301 (N_301,In_936,In_1205);
nor U302 (N_302,In_555,In_363);
xnor U303 (N_303,In_226,In_1040);
and U304 (N_304,In_171,In_1096);
xor U305 (N_305,In_1033,In_276);
or U306 (N_306,In_814,In_1172);
nand U307 (N_307,In_643,In_1355);
and U308 (N_308,In_515,In_159);
xor U309 (N_309,In_1409,In_1384);
nor U310 (N_310,In_457,In_480);
or U311 (N_311,In_318,In_1411);
and U312 (N_312,In_908,In_1423);
nand U313 (N_313,In_966,In_1203);
nor U314 (N_314,In_768,In_721);
nand U315 (N_315,In_1128,In_784);
and U316 (N_316,In_1335,In_58);
nor U317 (N_317,In_362,In_615);
and U318 (N_318,In_1430,In_921);
and U319 (N_319,In_323,In_530);
or U320 (N_320,In_1026,In_285);
xnor U321 (N_321,In_325,In_1357);
xor U322 (N_322,In_383,In_308);
nand U323 (N_323,In_985,In_1456);
nand U324 (N_324,In_1462,In_1066);
and U325 (N_325,In_1113,In_1350);
or U326 (N_326,In_201,In_1006);
xnor U327 (N_327,In_1014,In_1398);
or U328 (N_328,In_512,In_1236);
nor U329 (N_329,In_856,In_1265);
xor U330 (N_330,In_158,In_1150);
nand U331 (N_331,In_572,In_994);
or U332 (N_332,In_186,In_871);
xnor U333 (N_333,In_136,In_1428);
xnor U334 (N_334,In_794,In_826);
nor U335 (N_335,In_324,In_952);
nor U336 (N_336,In_810,In_84);
or U337 (N_337,In_609,In_191);
or U338 (N_338,In_529,In_1001);
nor U339 (N_339,In_1235,In_1385);
xor U340 (N_340,In_462,In_190);
and U341 (N_341,In_57,In_228);
xor U342 (N_342,In_1212,In_775);
xor U343 (N_343,In_1204,In_720);
and U344 (N_344,In_747,In_342);
and U345 (N_345,In_210,In_322);
nor U346 (N_346,In_237,In_491);
or U347 (N_347,In_150,In_421);
and U348 (N_348,In_557,In_238);
or U349 (N_349,In_1232,In_1182);
xnor U350 (N_350,In_12,In_1305);
and U351 (N_351,In_523,In_1140);
and U352 (N_352,In_1320,In_607);
and U353 (N_353,In_1100,In_1377);
nor U354 (N_354,In_1313,In_1183);
xnor U355 (N_355,In_1371,In_1243);
and U356 (N_356,In_303,In_472);
nand U357 (N_357,In_406,In_1222);
nand U358 (N_358,In_1124,In_1190);
or U359 (N_359,In_464,In_461);
and U360 (N_360,In_1449,In_1155);
nor U361 (N_361,In_446,In_145);
or U362 (N_362,In_573,In_712);
or U363 (N_363,In_808,In_818);
xnor U364 (N_364,In_953,In_1220);
xnor U365 (N_365,In_8,In_1133);
and U366 (N_366,In_1217,In_1112);
nor U367 (N_367,In_484,In_854);
nor U368 (N_368,In_498,In_1413);
nand U369 (N_369,In_105,In_213);
and U370 (N_370,In_157,In_559);
and U371 (N_371,In_260,In_129);
nand U372 (N_372,In_681,In_146);
and U373 (N_373,In_259,In_1000);
xnor U374 (N_374,In_1120,In_532);
xnor U375 (N_375,In_1264,In_1408);
xor U376 (N_376,In_1179,In_478);
xnor U377 (N_377,In_713,In_415);
nand U378 (N_378,In_33,In_1199);
and U379 (N_379,In_1390,In_340);
nand U380 (N_380,In_806,In_1078);
and U381 (N_381,In_52,In_270);
nand U382 (N_382,In_43,In_787);
nor U383 (N_383,In_239,In_1072);
or U384 (N_384,In_420,In_1034);
xor U385 (N_385,In_130,In_823);
nor U386 (N_386,In_1197,In_1334);
xnor U387 (N_387,In_957,In_1454);
xor U388 (N_388,In_1468,In_143);
or U389 (N_389,In_60,In_56);
or U390 (N_390,In_1444,In_809);
xnor U391 (N_391,In_642,In_1261);
nand U392 (N_392,In_404,In_1038);
or U393 (N_393,In_798,In_811);
nand U394 (N_394,In_366,In_1480);
or U395 (N_395,In_1063,In_686);
xnor U396 (N_396,In_995,In_847);
and U397 (N_397,In_718,In_1119);
or U398 (N_398,In_86,In_69);
xnor U399 (N_399,In_1132,In_983);
xnor U400 (N_400,In_53,In_941);
or U401 (N_401,In_845,In_1300);
and U402 (N_402,In_378,In_26);
nand U403 (N_403,In_1388,In_1275);
and U404 (N_404,In_511,In_192);
or U405 (N_405,In_737,In_63);
nand U406 (N_406,In_1492,In_999);
nor U407 (N_407,In_353,In_1131);
xor U408 (N_408,In_1448,In_1086);
nor U409 (N_409,In_203,In_141);
nor U410 (N_410,In_1319,In_687);
xor U411 (N_411,In_1121,In_698);
xnor U412 (N_412,In_589,In_1327);
or U413 (N_413,In_1037,In_333);
and U414 (N_414,In_89,In_543);
and U415 (N_415,In_640,In_1498);
nand U416 (N_416,In_819,In_1239);
or U417 (N_417,In_658,In_1389);
nor U418 (N_418,In_571,In_435);
xnor U419 (N_419,In_355,In_1253);
nor U420 (N_420,In_38,In_269);
nand U421 (N_421,In_204,In_1266);
xor U422 (N_422,In_656,In_110);
nand U423 (N_423,In_1165,In_1200);
xor U424 (N_424,In_1399,In_916);
nor U425 (N_425,In_128,In_1289);
nor U426 (N_426,In_1458,In_800);
or U427 (N_427,In_1210,In_125);
or U428 (N_428,In_407,In_93);
and U429 (N_429,In_1280,In_783);
xor U430 (N_430,In_542,In_881);
xnor U431 (N_431,In_314,In_840);
xnor U432 (N_432,In_264,In_1103);
nor U433 (N_433,In_1010,In_55);
nor U434 (N_434,In_1012,In_474);
and U435 (N_435,In_358,In_884);
and U436 (N_436,In_978,In_738);
xor U437 (N_437,In_458,In_649);
nor U438 (N_438,In_1185,In_893);
xor U439 (N_439,In_716,In_741);
nand U440 (N_440,In_79,In_927);
and U441 (N_441,In_288,In_66);
nor U442 (N_442,In_755,In_1130);
nor U443 (N_443,In_525,In_247);
nor U444 (N_444,In_1356,In_1170);
xor U445 (N_445,In_370,In_151);
nor U446 (N_446,In_1278,In_1346);
nand U447 (N_447,In_365,In_410);
nor U448 (N_448,In_503,In_1270);
nor U449 (N_449,In_517,In_469);
nor U450 (N_450,In_514,In_678);
nor U451 (N_451,In_258,In_294);
nand U452 (N_452,In_540,In_537);
xnor U453 (N_453,In_877,In_1324);
nor U454 (N_454,In_905,In_620);
xnor U455 (N_455,In_398,In_797);
nand U456 (N_456,In_1025,In_1488);
and U457 (N_457,In_867,In_278);
nand U458 (N_458,In_948,In_758);
or U459 (N_459,In_1404,In_107);
nand U460 (N_460,In_924,In_1017);
and U461 (N_461,In_328,In_541);
nand U462 (N_462,In_602,In_790);
or U463 (N_463,In_722,In_1045);
and U464 (N_464,In_222,In_1196);
nor U465 (N_465,In_821,In_414);
or U466 (N_466,In_22,In_662);
and U467 (N_467,In_1111,In_1459);
or U468 (N_468,In_911,In_1304);
xor U469 (N_469,In_938,In_980);
xnor U470 (N_470,In_350,In_305);
and U471 (N_471,In_296,In_1326);
nand U472 (N_472,In_970,In_531);
or U473 (N_473,In_118,In_1392);
nor U474 (N_474,In_1046,In_504);
or U475 (N_475,In_749,In_534);
nor U476 (N_476,In_1312,In_85);
nand U477 (N_477,In_104,In_1259);
nor U478 (N_478,In_64,In_633);
xor U479 (N_479,In_466,In_1003);
and U480 (N_480,In_178,In_714);
nand U481 (N_481,In_1245,In_154);
xnor U482 (N_482,In_706,In_670);
xnor U483 (N_483,In_1129,In_866);
xor U484 (N_484,In_548,In_1422);
nor U485 (N_485,In_397,In_774);
nor U486 (N_486,In_641,In_284);
or U487 (N_487,In_179,In_594);
or U488 (N_488,In_1005,In_1369);
nor U489 (N_489,In_7,In_1216);
or U490 (N_490,In_240,In_676);
or U491 (N_491,In_1436,In_163);
or U492 (N_492,In_510,In_1318);
xnor U493 (N_493,In_5,In_254);
xor U494 (N_494,In_560,In_30);
or U495 (N_495,In_1021,In_746);
or U496 (N_496,In_899,In_973);
xor U497 (N_497,In_1349,In_232);
nand U498 (N_498,In_1122,In_688);
nor U499 (N_499,In_427,In_62);
xor U500 (N_500,In_367,In_694);
nor U501 (N_501,In_329,In_667);
xor U502 (N_502,In_1049,In_878);
or U503 (N_503,In_1395,In_387);
and U504 (N_504,In_1027,In_1370);
xor U505 (N_505,In_1206,In_910);
xnor U506 (N_506,In_1302,In_556);
nor U507 (N_507,In_429,In_41);
nand U508 (N_508,In_1453,In_1373);
nand U509 (N_509,In_255,In_65);
nand U510 (N_510,In_892,In_283);
and U511 (N_511,In_1137,In_702);
nor U512 (N_512,In_138,In_701);
nor U513 (N_513,In_1114,In_1447);
and U514 (N_514,In_395,In_1344);
xnor U515 (N_515,In_689,In_1393);
xnor U516 (N_516,In_249,In_262);
nor U517 (N_517,In_454,In_317);
and U518 (N_518,In_1214,In_425);
xor U519 (N_519,In_578,In_1470);
xnor U520 (N_520,In_467,In_1314);
xnor U521 (N_521,In_1041,In_495);
nand U522 (N_522,In_1421,In_1405);
nand U523 (N_523,In_1065,In_996);
nand U524 (N_524,In_471,In_817);
nor U525 (N_525,In_1386,In_715);
and U526 (N_526,In_6,In_812);
xnor U527 (N_527,In_424,In_252);
nand U528 (N_528,In_624,In_780);
nand U529 (N_529,In_198,In_570);
nand U530 (N_530,In_792,In_287);
or U531 (N_531,In_16,In_1048);
and U532 (N_532,In_214,In_586);
nand U533 (N_533,In_74,In_1186);
or U534 (N_534,In_655,In_268);
or U535 (N_535,In_1117,In_321);
nand U536 (N_536,In_1360,In_1195);
nor U537 (N_537,In_961,In_1452);
xnor U538 (N_538,In_765,In_693);
nand U539 (N_539,In_1427,In_1213);
nand U540 (N_540,In_579,In_388);
xnor U541 (N_541,In_1286,In_1175);
and U542 (N_542,In_445,In_120);
and U543 (N_543,In_1079,In_175);
and U544 (N_544,In_116,In_672);
and U545 (N_545,In_1341,In_700);
nand U546 (N_546,In_796,In_590);
nor U547 (N_547,In_295,In_273);
nand U548 (N_548,In_1250,In_172);
and U549 (N_549,In_896,In_1348);
xnor U550 (N_550,In_1198,In_1426);
or U551 (N_551,In_1039,In_1321);
or U552 (N_552,In_1325,In_1020);
and U553 (N_553,In_913,In_950);
or U554 (N_554,In_1365,In_740);
nor U555 (N_555,In_1092,In_1149);
nand U556 (N_556,In_432,In_1018);
nand U557 (N_557,In_815,In_169);
xnor U558 (N_558,In_1147,In_539);
nor U559 (N_559,In_36,In_1440);
and U560 (N_560,In_576,In_1361);
nand U561 (N_561,In_35,In_1331);
and U562 (N_562,In_439,In_874);
or U563 (N_563,In_1163,In_1176);
xor U564 (N_564,In_1489,In_1052);
or U565 (N_565,In_1310,In_1397);
and U566 (N_566,In_1184,In_1160);
nand U567 (N_567,In_161,In_756);
xnor U568 (N_568,In_1379,In_831);
and U569 (N_569,In_748,In_1297);
nor U570 (N_570,In_1256,In_88);
xor U571 (N_571,In_960,In_1076);
nand U572 (N_572,In_411,In_149);
nand U573 (N_573,In_1077,In_403);
and U574 (N_574,In_44,In_550);
nand U575 (N_575,In_890,In_947);
nand U576 (N_576,In_1366,In_368);
nor U577 (N_577,In_1472,In_816);
and U578 (N_578,In_705,In_724);
nor U579 (N_579,In_1284,In_1159);
xnor U580 (N_580,In_453,In_1234);
xnor U581 (N_581,In_263,In_1074);
nand U582 (N_582,In_998,In_997);
nor U583 (N_583,In_436,In_123);
nand U584 (N_584,In_711,In_132);
nor U585 (N_585,In_1247,In_1107);
and U586 (N_586,In_114,In_944);
or U587 (N_587,In_332,In_750);
nand U588 (N_588,In_90,In_575);
xor U589 (N_589,In_433,In_853);
nand U590 (N_590,In_731,In_304);
nand U591 (N_591,In_993,In_155);
xor U592 (N_592,In_562,In_1309);
nand U593 (N_593,In_1031,In_683);
nor U594 (N_594,In_1219,In_487);
xor U595 (N_595,In_634,In_1490);
xor U596 (N_596,In_1268,In_50);
nor U597 (N_597,In_1022,In_183);
nand U598 (N_598,In_904,In_804);
and U599 (N_599,In_386,In_1101);
and U600 (N_600,In_253,In_32);
or U601 (N_601,In_1402,In_144);
or U602 (N_602,In_1015,In_488);
nand U603 (N_603,In_80,In_1463);
and U604 (N_604,In_621,In_1097);
nor U605 (N_605,In_1431,In_470);
xnor U606 (N_606,In_1004,In_1281);
and U607 (N_607,In_1194,In_1467);
xnor U608 (N_608,In_1381,In_1109);
xor U609 (N_609,In_1110,In_162);
nand U610 (N_610,In_1102,In_194);
or U611 (N_611,In_1162,In_547);
nand U612 (N_612,In_393,In_526);
or U613 (N_613,In_1359,In_788);
or U614 (N_614,In_685,In_1466);
xor U615 (N_615,In_1415,In_894);
or U616 (N_616,In_1368,In_1376);
and U617 (N_617,In_1244,In_1083);
and U618 (N_618,In_167,In_838);
xnor U619 (N_619,In_933,In_1251);
or U620 (N_620,In_1246,In_9);
and U621 (N_621,In_241,In_551);
and U622 (N_622,In_1142,In_1276);
nand U623 (N_623,In_659,In_1445);
nand U624 (N_624,In_1240,In_505);
and U625 (N_625,In_243,In_209);
xor U626 (N_626,In_538,In_14);
xnor U627 (N_627,In_359,In_919);
nand U628 (N_628,In_168,In_623);
xor U629 (N_629,In_68,In_992);
nand U630 (N_630,In_1383,In_1435);
nor U631 (N_631,In_1060,In_914);
or U632 (N_632,In_221,In_990);
xor U633 (N_633,In_1136,In_1257);
nor U634 (N_634,In_483,In_1419);
xor U635 (N_635,In_943,In_127);
nand U636 (N_636,In_1337,In_1231);
xor U637 (N_637,In_140,In_888);
xnor U638 (N_638,In_1375,In_1134);
xnor U639 (N_639,In_852,In_637);
xnor U640 (N_640,In_799,In_631);
nor U641 (N_641,In_959,In_381);
nor U642 (N_642,In_371,In_42);
nor U643 (N_643,In_1242,In_1487);
and U644 (N_644,In_1260,In_266);
and U645 (N_645,In_97,In_152);
or U646 (N_646,In_1032,In_437);
and U647 (N_647,In_958,In_1486);
xor U648 (N_648,In_895,In_207);
nand U649 (N_649,In_1473,In_972);
nor U650 (N_650,In_1153,In_587);
xnor U651 (N_651,In_1258,In_417);
or U652 (N_652,In_1108,In_848);
or U653 (N_653,In_449,In_1255);
and U654 (N_654,In_416,In_934);
nand U655 (N_655,In_1207,In_177);
nand U656 (N_656,In_626,In_1050);
xor U657 (N_657,In_1044,In_280);
and U658 (N_658,In_1007,In_126);
or U659 (N_659,In_327,In_653);
xor U660 (N_660,In_1059,In_153);
xor U661 (N_661,In_842,In_199);
or U662 (N_662,In_759,In_830);
or U663 (N_663,In_592,In_302);
nor U664 (N_664,In_1042,In_925);
or U665 (N_665,In_336,In_92);
nand U666 (N_666,In_889,In_1123);
xor U667 (N_667,In_289,In_497);
xor U668 (N_668,In_657,In_673);
or U669 (N_669,In_599,In_502);
or U670 (N_670,In_1288,In_188);
nor U671 (N_671,In_752,In_1401);
xor U672 (N_672,In_428,In_234);
nor U673 (N_673,In_671,In_1322);
nand U674 (N_674,In_494,In_1329);
nand U675 (N_675,In_1056,In_77);
xnor U676 (N_676,In_1343,In_773);
nor U677 (N_677,In_533,In_292);
nand U678 (N_678,In_1482,In_844);
and U679 (N_679,In_1424,In_293);
and U680 (N_680,In_1442,In_803);
nor U681 (N_681,In_486,In_1483);
xor U682 (N_682,In_1188,In_535);
and U683 (N_683,In_282,In_301);
nand U684 (N_684,In_182,In_1420);
or U685 (N_685,In_40,In_1156);
nor U686 (N_686,In_507,In_935);
xor U687 (N_687,In_988,In_164);
nand U688 (N_688,In_769,In_1283);
and U689 (N_689,In_1164,In_1202);
or U690 (N_690,In_447,In_1469);
xnor U691 (N_691,In_1364,In_1191);
nand U692 (N_692,In_697,In_1461);
nand U693 (N_693,In_566,In_522);
xor U694 (N_694,In_918,In_879);
nand U695 (N_695,In_1441,In_1410);
nand U696 (N_696,In_1273,In_297);
and U697 (N_697,In_229,In_1080);
or U698 (N_698,In_1491,In_1339);
or U699 (N_699,In_1144,In_630);
nor U700 (N_700,In_880,In_725);
nor U701 (N_701,In_196,In_703);
nand U702 (N_702,In_1158,In_499);
or U703 (N_703,In_930,In_903);
nor U704 (N_704,In_574,In_639);
nand U705 (N_705,In_516,In_96);
or U706 (N_706,In_1394,In_115);
nor U707 (N_707,In_187,In_20);
xnor U708 (N_708,In_382,In_100);
and U709 (N_709,In_15,In_500);
or U710 (N_710,In_900,In_456);
or U711 (N_711,In_1023,In_728);
xor U712 (N_712,In_475,In_604);
and U713 (N_713,In_59,In_597);
xnor U714 (N_714,In_1460,In_1455);
nand U715 (N_715,In_661,In_1285);
or U716 (N_716,In_170,In_835);
nand U717 (N_717,In_1094,In_373);
nand U718 (N_718,In_753,In_618);
nor U719 (N_719,In_408,In_964);
nor U720 (N_720,In_963,In_1432);
xnor U721 (N_721,In_413,In_1362);
xnor U722 (N_722,In_564,In_405);
xnor U723 (N_723,In_795,In_646);
xor U724 (N_724,In_27,In_244);
nor U725 (N_725,In_372,In_441);
nor U726 (N_726,In_1209,In_585);
xor U727 (N_727,In_246,In_1057);
or U728 (N_728,In_805,In_2);
or U729 (N_729,In_612,In_1354);
xnor U730 (N_730,In_309,In_614);
and U731 (N_731,In_1084,In_352);
or U732 (N_732,In_802,In_761);
xnor U733 (N_733,In_1485,In_1070);
nor U734 (N_734,In_1169,In_451);
nor U735 (N_735,In_236,In_704);
and U736 (N_736,In_628,In_71);
xnor U737 (N_737,In_1311,In_730);
or U738 (N_738,In_265,In_554);
and U739 (N_739,In_987,In_939);
nand U740 (N_740,In_926,In_465);
nand U741 (N_741,In_707,In_1291);
nor U742 (N_742,In_886,In_211);
xnor U743 (N_743,In_419,In_613);
nor U744 (N_744,In_1263,In_1105);
nand U745 (N_745,In_134,In_349);
nor U746 (N_746,In_527,In_719);
xor U747 (N_747,In_195,In_937);
nor U748 (N_748,In_1308,In_489);
and U749 (N_749,In_267,In_1494);
xnor U750 (N_750,In_1439,In_67);
nor U751 (N_751,In_779,In_411);
and U752 (N_752,In_848,In_1191);
or U753 (N_753,In_1278,In_1190);
nand U754 (N_754,In_944,In_1335);
and U755 (N_755,In_338,In_1194);
nand U756 (N_756,In_765,In_631);
and U757 (N_757,In_1002,In_225);
and U758 (N_758,In_1198,In_1376);
nor U759 (N_759,In_251,In_1359);
or U760 (N_760,In_1075,In_597);
and U761 (N_761,In_1282,In_4);
nor U762 (N_762,In_16,In_748);
nor U763 (N_763,In_617,In_1225);
or U764 (N_764,In_1125,In_1169);
or U765 (N_765,In_565,In_1289);
nor U766 (N_766,In_567,In_206);
and U767 (N_767,In_201,In_393);
or U768 (N_768,In_772,In_830);
xnor U769 (N_769,In_732,In_1023);
xnor U770 (N_770,In_201,In_114);
or U771 (N_771,In_943,In_1341);
xnor U772 (N_772,In_1138,In_405);
or U773 (N_773,In_990,In_1219);
or U774 (N_774,In_1110,In_1185);
nor U775 (N_775,In_901,In_1294);
or U776 (N_776,In_1222,In_187);
xor U777 (N_777,In_1372,In_1066);
xor U778 (N_778,In_13,In_1113);
and U779 (N_779,In_1240,In_768);
nor U780 (N_780,In_294,In_234);
or U781 (N_781,In_1119,In_60);
nor U782 (N_782,In_842,In_611);
and U783 (N_783,In_1210,In_907);
xor U784 (N_784,In_63,In_242);
or U785 (N_785,In_720,In_840);
and U786 (N_786,In_171,In_980);
nor U787 (N_787,In_764,In_19);
nor U788 (N_788,In_1184,In_865);
xnor U789 (N_789,In_1363,In_526);
nor U790 (N_790,In_1186,In_757);
nor U791 (N_791,In_1096,In_76);
xor U792 (N_792,In_988,In_981);
nor U793 (N_793,In_1286,In_1);
nand U794 (N_794,In_1020,In_690);
or U795 (N_795,In_1025,In_1475);
xor U796 (N_796,In_1345,In_1098);
and U797 (N_797,In_734,In_1354);
or U798 (N_798,In_490,In_95);
nor U799 (N_799,In_422,In_289);
or U800 (N_800,In_1004,In_859);
nor U801 (N_801,In_197,In_1036);
or U802 (N_802,In_303,In_53);
nor U803 (N_803,In_1372,In_1404);
xor U804 (N_804,In_594,In_172);
or U805 (N_805,In_1159,In_158);
or U806 (N_806,In_655,In_546);
or U807 (N_807,In_782,In_1140);
and U808 (N_808,In_105,In_1018);
or U809 (N_809,In_1294,In_6);
nor U810 (N_810,In_292,In_118);
and U811 (N_811,In_517,In_473);
and U812 (N_812,In_1055,In_622);
nor U813 (N_813,In_419,In_754);
xor U814 (N_814,In_633,In_321);
or U815 (N_815,In_1270,In_889);
and U816 (N_816,In_1173,In_249);
or U817 (N_817,In_849,In_438);
nor U818 (N_818,In_802,In_1359);
nand U819 (N_819,In_1333,In_1214);
nand U820 (N_820,In_430,In_766);
or U821 (N_821,In_329,In_360);
and U822 (N_822,In_281,In_288);
xor U823 (N_823,In_575,In_739);
or U824 (N_824,In_758,In_887);
xnor U825 (N_825,In_981,In_1426);
nand U826 (N_826,In_988,In_663);
nor U827 (N_827,In_924,In_340);
and U828 (N_828,In_482,In_415);
or U829 (N_829,In_456,In_1421);
nand U830 (N_830,In_228,In_1029);
or U831 (N_831,In_1470,In_372);
or U832 (N_832,In_84,In_95);
xnor U833 (N_833,In_122,In_372);
nand U834 (N_834,In_44,In_1379);
or U835 (N_835,In_766,In_1180);
nor U836 (N_836,In_149,In_799);
or U837 (N_837,In_1122,In_467);
xor U838 (N_838,In_870,In_1091);
and U839 (N_839,In_1077,In_196);
nand U840 (N_840,In_463,In_32);
or U841 (N_841,In_941,In_1043);
or U842 (N_842,In_982,In_410);
nor U843 (N_843,In_621,In_578);
or U844 (N_844,In_138,In_344);
xor U845 (N_845,In_622,In_196);
xor U846 (N_846,In_20,In_592);
or U847 (N_847,In_386,In_407);
nor U848 (N_848,In_147,In_116);
and U849 (N_849,In_788,In_1065);
and U850 (N_850,In_1468,In_869);
or U851 (N_851,In_1495,In_201);
and U852 (N_852,In_85,In_599);
or U853 (N_853,In_1363,In_326);
nor U854 (N_854,In_463,In_775);
nor U855 (N_855,In_182,In_897);
and U856 (N_856,In_1190,In_698);
or U857 (N_857,In_1281,In_229);
and U858 (N_858,In_567,In_534);
xnor U859 (N_859,In_1037,In_182);
and U860 (N_860,In_777,In_1106);
or U861 (N_861,In_1422,In_841);
xor U862 (N_862,In_799,In_1092);
xnor U863 (N_863,In_123,In_852);
and U864 (N_864,In_663,In_1200);
and U865 (N_865,In_17,In_148);
xor U866 (N_866,In_806,In_1150);
nand U867 (N_867,In_16,In_1332);
xor U868 (N_868,In_110,In_920);
or U869 (N_869,In_666,In_670);
nor U870 (N_870,In_356,In_0);
nand U871 (N_871,In_565,In_232);
nor U872 (N_872,In_992,In_765);
xor U873 (N_873,In_77,In_551);
and U874 (N_874,In_880,In_1469);
or U875 (N_875,In_956,In_693);
nand U876 (N_876,In_886,In_1258);
xor U877 (N_877,In_431,In_1238);
nand U878 (N_878,In_280,In_463);
nor U879 (N_879,In_644,In_1391);
nand U880 (N_880,In_574,In_275);
xnor U881 (N_881,In_898,In_420);
or U882 (N_882,In_914,In_144);
or U883 (N_883,In_1198,In_1026);
nor U884 (N_884,In_966,In_756);
nand U885 (N_885,In_845,In_469);
nand U886 (N_886,In_474,In_766);
nor U887 (N_887,In_1422,In_1299);
or U888 (N_888,In_33,In_752);
xor U889 (N_889,In_1320,In_883);
xnor U890 (N_890,In_1217,In_170);
xnor U891 (N_891,In_141,In_378);
xor U892 (N_892,In_427,In_1460);
xnor U893 (N_893,In_1007,In_990);
nor U894 (N_894,In_460,In_822);
xnor U895 (N_895,In_1106,In_1294);
xnor U896 (N_896,In_1227,In_1422);
and U897 (N_897,In_682,In_727);
and U898 (N_898,In_240,In_1134);
or U899 (N_899,In_974,In_30);
nand U900 (N_900,In_929,In_1405);
xnor U901 (N_901,In_14,In_1430);
xnor U902 (N_902,In_1040,In_1192);
nand U903 (N_903,In_1281,In_962);
nor U904 (N_904,In_581,In_591);
xnor U905 (N_905,In_1280,In_255);
nor U906 (N_906,In_1172,In_1212);
nor U907 (N_907,In_1458,In_531);
nand U908 (N_908,In_1420,In_1481);
nor U909 (N_909,In_484,In_487);
nand U910 (N_910,In_851,In_698);
nand U911 (N_911,In_1014,In_61);
nor U912 (N_912,In_241,In_733);
nor U913 (N_913,In_989,In_332);
and U914 (N_914,In_1437,In_602);
and U915 (N_915,In_1292,In_16);
and U916 (N_916,In_1377,In_1301);
xor U917 (N_917,In_1006,In_120);
or U918 (N_918,In_352,In_135);
or U919 (N_919,In_414,In_1438);
nor U920 (N_920,In_98,In_879);
and U921 (N_921,In_729,In_364);
and U922 (N_922,In_736,In_867);
and U923 (N_923,In_1477,In_1201);
nand U924 (N_924,In_607,In_1235);
and U925 (N_925,In_1242,In_940);
nor U926 (N_926,In_1167,In_1329);
nand U927 (N_927,In_1253,In_1209);
nand U928 (N_928,In_599,In_842);
xor U929 (N_929,In_1032,In_1491);
or U930 (N_930,In_254,In_902);
xor U931 (N_931,In_18,In_300);
or U932 (N_932,In_383,In_809);
nand U933 (N_933,In_1444,In_69);
nand U934 (N_934,In_1099,In_1076);
and U935 (N_935,In_1225,In_506);
nor U936 (N_936,In_744,In_1035);
nand U937 (N_937,In_789,In_570);
or U938 (N_938,In_1442,In_1130);
and U939 (N_939,In_988,In_1447);
and U940 (N_940,In_646,In_757);
nand U941 (N_941,In_1199,In_575);
nand U942 (N_942,In_1181,In_1134);
nand U943 (N_943,In_452,In_1344);
nor U944 (N_944,In_843,In_895);
nor U945 (N_945,In_975,In_1234);
or U946 (N_946,In_920,In_964);
xor U947 (N_947,In_953,In_1159);
xor U948 (N_948,In_619,In_1179);
xor U949 (N_949,In_495,In_9);
or U950 (N_950,In_792,In_911);
nor U951 (N_951,In_485,In_114);
or U952 (N_952,In_707,In_32);
xor U953 (N_953,In_609,In_1387);
nor U954 (N_954,In_977,In_1386);
or U955 (N_955,In_32,In_1099);
nand U956 (N_956,In_254,In_1089);
and U957 (N_957,In_1275,In_193);
nor U958 (N_958,In_717,In_501);
or U959 (N_959,In_1043,In_507);
or U960 (N_960,In_672,In_1399);
and U961 (N_961,In_245,In_850);
xor U962 (N_962,In_1099,In_78);
nor U963 (N_963,In_527,In_304);
and U964 (N_964,In_274,In_1010);
nor U965 (N_965,In_158,In_202);
xor U966 (N_966,In_688,In_559);
or U967 (N_967,In_1203,In_747);
or U968 (N_968,In_1271,In_1100);
nand U969 (N_969,In_50,In_586);
or U970 (N_970,In_232,In_1169);
xnor U971 (N_971,In_754,In_1058);
xor U972 (N_972,In_1451,In_441);
nand U973 (N_973,In_453,In_1208);
nand U974 (N_974,In_920,In_614);
and U975 (N_975,In_846,In_607);
nand U976 (N_976,In_1257,In_1460);
or U977 (N_977,In_331,In_1008);
nor U978 (N_978,In_201,In_601);
nand U979 (N_979,In_1492,In_156);
or U980 (N_980,In_1196,In_102);
nand U981 (N_981,In_642,In_1354);
and U982 (N_982,In_1454,In_1270);
xnor U983 (N_983,In_1138,In_1251);
and U984 (N_984,In_479,In_701);
or U985 (N_985,In_228,In_1392);
nand U986 (N_986,In_1141,In_684);
nand U987 (N_987,In_1037,In_0);
xnor U988 (N_988,In_995,In_856);
xnor U989 (N_989,In_911,In_527);
xnor U990 (N_990,In_773,In_1125);
nor U991 (N_991,In_1396,In_613);
nor U992 (N_992,In_881,In_554);
and U993 (N_993,In_1185,In_557);
nand U994 (N_994,In_784,In_1225);
and U995 (N_995,In_1077,In_1267);
or U996 (N_996,In_40,In_1270);
xor U997 (N_997,In_660,In_938);
nand U998 (N_998,In_325,In_1407);
xnor U999 (N_999,In_1182,In_108);
and U1000 (N_1000,In_256,In_429);
xnor U1001 (N_1001,In_217,In_256);
and U1002 (N_1002,In_348,In_372);
or U1003 (N_1003,In_968,In_1425);
or U1004 (N_1004,In_561,In_1277);
or U1005 (N_1005,In_966,In_787);
nor U1006 (N_1006,In_661,In_44);
nand U1007 (N_1007,In_804,In_1413);
xnor U1008 (N_1008,In_1461,In_431);
nor U1009 (N_1009,In_842,In_850);
xor U1010 (N_1010,In_927,In_263);
xor U1011 (N_1011,In_995,In_164);
or U1012 (N_1012,In_172,In_444);
and U1013 (N_1013,In_481,In_365);
xor U1014 (N_1014,In_1257,In_734);
xnor U1015 (N_1015,In_1466,In_850);
nor U1016 (N_1016,In_761,In_1435);
nor U1017 (N_1017,In_1037,In_200);
nand U1018 (N_1018,In_815,In_324);
and U1019 (N_1019,In_1171,In_1457);
nand U1020 (N_1020,In_602,In_651);
nand U1021 (N_1021,In_1135,In_631);
and U1022 (N_1022,In_728,In_1393);
and U1023 (N_1023,In_625,In_1253);
xor U1024 (N_1024,In_1480,In_865);
or U1025 (N_1025,In_321,In_925);
nor U1026 (N_1026,In_1001,In_107);
xnor U1027 (N_1027,In_282,In_631);
xor U1028 (N_1028,In_775,In_801);
xnor U1029 (N_1029,In_1000,In_375);
nor U1030 (N_1030,In_1345,In_540);
and U1031 (N_1031,In_1353,In_697);
xnor U1032 (N_1032,In_1404,In_584);
xor U1033 (N_1033,In_972,In_704);
or U1034 (N_1034,In_1138,In_89);
nand U1035 (N_1035,In_1297,In_332);
nor U1036 (N_1036,In_1348,In_1017);
or U1037 (N_1037,In_84,In_795);
or U1038 (N_1038,In_1188,In_745);
xnor U1039 (N_1039,In_195,In_236);
or U1040 (N_1040,In_1367,In_561);
nand U1041 (N_1041,In_438,In_475);
nand U1042 (N_1042,In_483,In_762);
and U1043 (N_1043,In_1268,In_1032);
nor U1044 (N_1044,In_1259,In_1282);
nand U1045 (N_1045,In_1065,In_626);
nand U1046 (N_1046,In_543,In_1426);
nor U1047 (N_1047,In_369,In_264);
and U1048 (N_1048,In_885,In_131);
xor U1049 (N_1049,In_382,In_1282);
and U1050 (N_1050,In_680,In_1377);
and U1051 (N_1051,In_21,In_25);
nand U1052 (N_1052,In_1133,In_629);
or U1053 (N_1053,In_1221,In_131);
xnor U1054 (N_1054,In_832,In_537);
or U1055 (N_1055,In_1228,In_292);
nand U1056 (N_1056,In_1102,In_171);
xor U1057 (N_1057,In_1091,In_901);
nand U1058 (N_1058,In_760,In_112);
and U1059 (N_1059,In_990,In_1193);
nor U1060 (N_1060,In_389,In_58);
and U1061 (N_1061,In_510,In_652);
xnor U1062 (N_1062,In_611,In_249);
nand U1063 (N_1063,In_1346,In_499);
and U1064 (N_1064,In_1234,In_1050);
xor U1065 (N_1065,In_258,In_727);
or U1066 (N_1066,In_502,In_1300);
or U1067 (N_1067,In_764,In_610);
and U1068 (N_1068,In_1199,In_876);
nor U1069 (N_1069,In_774,In_98);
and U1070 (N_1070,In_1397,In_255);
and U1071 (N_1071,In_573,In_230);
nand U1072 (N_1072,In_1347,In_1093);
xor U1073 (N_1073,In_450,In_544);
and U1074 (N_1074,In_1294,In_1398);
xor U1075 (N_1075,In_287,In_1478);
nand U1076 (N_1076,In_988,In_103);
nor U1077 (N_1077,In_12,In_237);
and U1078 (N_1078,In_404,In_367);
xnor U1079 (N_1079,In_161,In_872);
and U1080 (N_1080,In_477,In_435);
xnor U1081 (N_1081,In_1332,In_1353);
nor U1082 (N_1082,In_1232,In_458);
or U1083 (N_1083,In_1481,In_291);
nand U1084 (N_1084,In_144,In_1249);
xnor U1085 (N_1085,In_497,In_914);
nand U1086 (N_1086,In_504,In_91);
nor U1087 (N_1087,In_216,In_373);
or U1088 (N_1088,In_339,In_1043);
nand U1089 (N_1089,In_293,In_1314);
or U1090 (N_1090,In_851,In_758);
nor U1091 (N_1091,In_190,In_250);
and U1092 (N_1092,In_419,In_1350);
xnor U1093 (N_1093,In_1404,In_28);
and U1094 (N_1094,In_1194,In_1061);
nor U1095 (N_1095,In_959,In_52);
nor U1096 (N_1096,In_1484,In_740);
nor U1097 (N_1097,In_1068,In_770);
xnor U1098 (N_1098,In_633,In_957);
xor U1099 (N_1099,In_754,In_979);
or U1100 (N_1100,In_756,In_805);
xor U1101 (N_1101,In_1419,In_1334);
nor U1102 (N_1102,In_908,In_1477);
and U1103 (N_1103,In_873,In_329);
and U1104 (N_1104,In_694,In_40);
and U1105 (N_1105,In_229,In_697);
nor U1106 (N_1106,In_568,In_188);
xnor U1107 (N_1107,In_623,In_1213);
and U1108 (N_1108,In_608,In_1345);
xnor U1109 (N_1109,In_1270,In_394);
nor U1110 (N_1110,In_493,In_1008);
or U1111 (N_1111,In_499,In_210);
and U1112 (N_1112,In_328,In_1264);
xor U1113 (N_1113,In_635,In_658);
or U1114 (N_1114,In_1277,In_1075);
nor U1115 (N_1115,In_889,In_975);
xnor U1116 (N_1116,In_431,In_1322);
nand U1117 (N_1117,In_1387,In_260);
nor U1118 (N_1118,In_1333,In_436);
and U1119 (N_1119,In_529,In_849);
nand U1120 (N_1120,In_847,In_424);
nor U1121 (N_1121,In_284,In_368);
or U1122 (N_1122,In_429,In_440);
xor U1123 (N_1123,In_62,In_735);
xor U1124 (N_1124,In_1477,In_302);
or U1125 (N_1125,In_299,In_950);
xor U1126 (N_1126,In_228,In_95);
nor U1127 (N_1127,In_215,In_945);
nor U1128 (N_1128,In_388,In_1142);
nor U1129 (N_1129,In_257,In_1134);
and U1130 (N_1130,In_1430,In_880);
or U1131 (N_1131,In_359,In_416);
nor U1132 (N_1132,In_1493,In_1237);
nand U1133 (N_1133,In_478,In_266);
xor U1134 (N_1134,In_784,In_78);
and U1135 (N_1135,In_389,In_486);
or U1136 (N_1136,In_481,In_374);
or U1137 (N_1137,In_0,In_296);
and U1138 (N_1138,In_778,In_569);
nor U1139 (N_1139,In_1229,In_1455);
nor U1140 (N_1140,In_603,In_743);
and U1141 (N_1141,In_889,In_354);
and U1142 (N_1142,In_1379,In_825);
xor U1143 (N_1143,In_463,In_1307);
or U1144 (N_1144,In_444,In_794);
nor U1145 (N_1145,In_340,In_1395);
and U1146 (N_1146,In_459,In_284);
xor U1147 (N_1147,In_51,In_603);
nand U1148 (N_1148,In_421,In_521);
xnor U1149 (N_1149,In_1412,In_1442);
xor U1150 (N_1150,In_369,In_969);
and U1151 (N_1151,In_933,In_609);
and U1152 (N_1152,In_876,In_197);
xor U1153 (N_1153,In_667,In_361);
nor U1154 (N_1154,In_263,In_1436);
nand U1155 (N_1155,In_1283,In_1392);
nor U1156 (N_1156,In_1287,In_1495);
nor U1157 (N_1157,In_1383,In_1094);
nand U1158 (N_1158,In_798,In_385);
nand U1159 (N_1159,In_1063,In_98);
nor U1160 (N_1160,In_384,In_371);
and U1161 (N_1161,In_557,In_7);
xnor U1162 (N_1162,In_499,In_184);
nand U1163 (N_1163,In_1137,In_1418);
nor U1164 (N_1164,In_316,In_39);
nor U1165 (N_1165,In_1233,In_412);
xor U1166 (N_1166,In_821,In_255);
nor U1167 (N_1167,In_870,In_939);
and U1168 (N_1168,In_707,In_190);
xor U1169 (N_1169,In_826,In_681);
xnor U1170 (N_1170,In_366,In_965);
xnor U1171 (N_1171,In_1199,In_370);
xnor U1172 (N_1172,In_442,In_98);
and U1173 (N_1173,In_1410,In_237);
and U1174 (N_1174,In_194,In_804);
nor U1175 (N_1175,In_671,In_60);
nand U1176 (N_1176,In_1421,In_597);
nor U1177 (N_1177,In_23,In_1084);
and U1178 (N_1178,In_447,In_1112);
and U1179 (N_1179,In_1335,In_1099);
nor U1180 (N_1180,In_186,In_1228);
or U1181 (N_1181,In_1045,In_244);
nand U1182 (N_1182,In_442,In_108);
nor U1183 (N_1183,In_167,In_1454);
nor U1184 (N_1184,In_1210,In_1163);
nor U1185 (N_1185,In_1014,In_362);
nor U1186 (N_1186,In_511,In_63);
and U1187 (N_1187,In_313,In_1314);
xnor U1188 (N_1188,In_182,In_808);
and U1189 (N_1189,In_36,In_423);
and U1190 (N_1190,In_1238,In_1163);
nor U1191 (N_1191,In_1274,In_203);
and U1192 (N_1192,In_498,In_1290);
xor U1193 (N_1193,In_452,In_573);
nor U1194 (N_1194,In_336,In_271);
xnor U1195 (N_1195,In_819,In_470);
nor U1196 (N_1196,In_1231,In_1475);
nand U1197 (N_1197,In_1359,In_654);
nor U1198 (N_1198,In_1484,In_979);
and U1199 (N_1199,In_1287,In_1083);
nand U1200 (N_1200,In_920,In_721);
xor U1201 (N_1201,In_67,In_789);
and U1202 (N_1202,In_38,In_877);
nand U1203 (N_1203,In_1195,In_312);
and U1204 (N_1204,In_1332,In_1174);
xnor U1205 (N_1205,In_1260,In_397);
xnor U1206 (N_1206,In_1371,In_191);
and U1207 (N_1207,In_827,In_945);
nor U1208 (N_1208,In_988,In_493);
nor U1209 (N_1209,In_427,In_771);
nand U1210 (N_1210,In_267,In_1212);
or U1211 (N_1211,In_811,In_202);
or U1212 (N_1212,In_1200,In_76);
nor U1213 (N_1213,In_952,In_26);
or U1214 (N_1214,In_775,In_635);
and U1215 (N_1215,In_828,In_688);
nor U1216 (N_1216,In_911,In_542);
and U1217 (N_1217,In_592,In_626);
nor U1218 (N_1218,In_86,In_960);
nor U1219 (N_1219,In_1117,In_1284);
nand U1220 (N_1220,In_887,In_729);
nor U1221 (N_1221,In_919,In_963);
nor U1222 (N_1222,In_334,In_360);
or U1223 (N_1223,In_75,In_548);
nand U1224 (N_1224,In_510,In_1252);
and U1225 (N_1225,In_548,In_61);
nor U1226 (N_1226,In_72,In_1077);
nand U1227 (N_1227,In_14,In_920);
xnor U1228 (N_1228,In_1019,In_1146);
xor U1229 (N_1229,In_389,In_626);
nand U1230 (N_1230,In_1460,In_460);
xnor U1231 (N_1231,In_1356,In_398);
nor U1232 (N_1232,In_748,In_919);
nand U1233 (N_1233,In_1335,In_727);
or U1234 (N_1234,In_25,In_994);
and U1235 (N_1235,In_282,In_1158);
nand U1236 (N_1236,In_1070,In_1381);
xor U1237 (N_1237,In_653,In_797);
or U1238 (N_1238,In_1072,In_492);
nand U1239 (N_1239,In_1064,In_596);
or U1240 (N_1240,In_161,In_1358);
or U1241 (N_1241,In_550,In_538);
nor U1242 (N_1242,In_781,In_1217);
nor U1243 (N_1243,In_1419,In_307);
nand U1244 (N_1244,In_249,In_1135);
nand U1245 (N_1245,In_493,In_1480);
nand U1246 (N_1246,In_1354,In_1305);
nand U1247 (N_1247,In_729,In_1467);
nand U1248 (N_1248,In_97,In_1001);
nand U1249 (N_1249,In_1326,In_319);
nor U1250 (N_1250,In_1135,In_1119);
nor U1251 (N_1251,In_1216,In_1268);
and U1252 (N_1252,In_294,In_178);
and U1253 (N_1253,In_1164,In_782);
or U1254 (N_1254,In_1182,In_1357);
and U1255 (N_1255,In_1378,In_874);
nand U1256 (N_1256,In_487,In_536);
xnor U1257 (N_1257,In_63,In_1453);
or U1258 (N_1258,In_584,In_664);
nand U1259 (N_1259,In_94,In_1313);
xnor U1260 (N_1260,In_505,In_76);
or U1261 (N_1261,In_702,In_199);
nand U1262 (N_1262,In_1168,In_794);
and U1263 (N_1263,In_1134,In_26);
or U1264 (N_1264,In_1359,In_17);
or U1265 (N_1265,In_1147,In_1011);
or U1266 (N_1266,In_92,In_22);
xnor U1267 (N_1267,In_1482,In_1123);
nand U1268 (N_1268,In_637,In_1461);
and U1269 (N_1269,In_1153,In_690);
nand U1270 (N_1270,In_819,In_336);
xor U1271 (N_1271,In_539,In_376);
or U1272 (N_1272,In_1240,In_359);
and U1273 (N_1273,In_66,In_1120);
nor U1274 (N_1274,In_767,In_461);
xnor U1275 (N_1275,In_234,In_304);
nor U1276 (N_1276,In_855,In_359);
or U1277 (N_1277,In_1184,In_310);
nand U1278 (N_1278,In_1149,In_1414);
xnor U1279 (N_1279,In_663,In_1276);
or U1280 (N_1280,In_514,In_94);
nor U1281 (N_1281,In_412,In_1195);
nand U1282 (N_1282,In_649,In_229);
nor U1283 (N_1283,In_114,In_85);
and U1284 (N_1284,In_371,In_805);
or U1285 (N_1285,In_1409,In_1310);
and U1286 (N_1286,In_772,In_11);
nand U1287 (N_1287,In_918,In_886);
or U1288 (N_1288,In_1048,In_825);
or U1289 (N_1289,In_27,In_1439);
nor U1290 (N_1290,In_1415,In_747);
nor U1291 (N_1291,In_1379,In_412);
or U1292 (N_1292,In_714,In_100);
nor U1293 (N_1293,In_238,In_19);
nand U1294 (N_1294,In_1217,In_1065);
nor U1295 (N_1295,In_349,In_1403);
xor U1296 (N_1296,In_185,In_869);
nor U1297 (N_1297,In_1205,In_979);
xnor U1298 (N_1298,In_1260,In_1095);
or U1299 (N_1299,In_723,In_1425);
xnor U1300 (N_1300,In_455,In_813);
xnor U1301 (N_1301,In_675,In_787);
nand U1302 (N_1302,In_966,In_49);
or U1303 (N_1303,In_215,In_824);
nand U1304 (N_1304,In_236,In_959);
or U1305 (N_1305,In_983,In_336);
and U1306 (N_1306,In_252,In_872);
and U1307 (N_1307,In_570,In_1022);
or U1308 (N_1308,In_1458,In_766);
or U1309 (N_1309,In_616,In_824);
or U1310 (N_1310,In_436,In_953);
nand U1311 (N_1311,In_675,In_380);
nor U1312 (N_1312,In_201,In_260);
xor U1313 (N_1313,In_455,In_711);
or U1314 (N_1314,In_1492,In_1072);
and U1315 (N_1315,In_1238,In_928);
and U1316 (N_1316,In_162,In_718);
or U1317 (N_1317,In_398,In_1319);
nand U1318 (N_1318,In_352,In_1296);
nor U1319 (N_1319,In_756,In_1280);
or U1320 (N_1320,In_1178,In_589);
nor U1321 (N_1321,In_1173,In_100);
and U1322 (N_1322,In_930,In_896);
or U1323 (N_1323,In_297,In_71);
and U1324 (N_1324,In_5,In_21);
xnor U1325 (N_1325,In_865,In_376);
nand U1326 (N_1326,In_478,In_915);
xor U1327 (N_1327,In_704,In_1114);
and U1328 (N_1328,In_554,In_1353);
and U1329 (N_1329,In_1298,In_1027);
and U1330 (N_1330,In_46,In_82);
or U1331 (N_1331,In_427,In_806);
nand U1332 (N_1332,In_872,In_322);
and U1333 (N_1333,In_782,In_855);
nor U1334 (N_1334,In_1223,In_802);
xor U1335 (N_1335,In_1472,In_1259);
nor U1336 (N_1336,In_823,In_471);
nor U1337 (N_1337,In_424,In_71);
xnor U1338 (N_1338,In_1136,In_1476);
and U1339 (N_1339,In_1337,In_215);
nor U1340 (N_1340,In_1008,In_555);
xnor U1341 (N_1341,In_852,In_754);
nor U1342 (N_1342,In_398,In_1145);
nor U1343 (N_1343,In_385,In_70);
xor U1344 (N_1344,In_1445,In_410);
nor U1345 (N_1345,In_215,In_582);
nand U1346 (N_1346,In_1268,In_1102);
nor U1347 (N_1347,In_707,In_221);
nor U1348 (N_1348,In_602,In_1020);
nor U1349 (N_1349,In_1082,In_633);
and U1350 (N_1350,In_1473,In_854);
and U1351 (N_1351,In_879,In_703);
or U1352 (N_1352,In_410,In_1376);
or U1353 (N_1353,In_99,In_251);
and U1354 (N_1354,In_648,In_0);
or U1355 (N_1355,In_833,In_480);
nor U1356 (N_1356,In_1012,In_145);
nand U1357 (N_1357,In_433,In_809);
nor U1358 (N_1358,In_18,In_221);
and U1359 (N_1359,In_1286,In_872);
nor U1360 (N_1360,In_1189,In_1014);
xnor U1361 (N_1361,In_585,In_1240);
and U1362 (N_1362,In_1109,In_1282);
nor U1363 (N_1363,In_816,In_139);
nor U1364 (N_1364,In_547,In_1494);
and U1365 (N_1365,In_556,In_126);
or U1366 (N_1366,In_1374,In_541);
nand U1367 (N_1367,In_290,In_788);
or U1368 (N_1368,In_444,In_235);
nand U1369 (N_1369,In_779,In_1099);
and U1370 (N_1370,In_1167,In_930);
xnor U1371 (N_1371,In_1192,In_1230);
or U1372 (N_1372,In_461,In_981);
and U1373 (N_1373,In_1491,In_624);
xnor U1374 (N_1374,In_644,In_462);
nor U1375 (N_1375,In_1119,In_1049);
xor U1376 (N_1376,In_506,In_51);
and U1377 (N_1377,In_1243,In_923);
nand U1378 (N_1378,In_1046,In_500);
xnor U1379 (N_1379,In_1048,In_136);
xor U1380 (N_1380,In_322,In_951);
or U1381 (N_1381,In_1305,In_847);
nor U1382 (N_1382,In_528,In_542);
xor U1383 (N_1383,In_768,In_1142);
or U1384 (N_1384,In_869,In_8);
nor U1385 (N_1385,In_641,In_1050);
xor U1386 (N_1386,In_758,In_1491);
or U1387 (N_1387,In_1021,In_1091);
xnor U1388 (N_1388,In_451,In_879);
xor U1389 (N_1389,In_582,In_894);
nand U1390 (N_1390,In_740,In_602);
or U1391 (N_1391,In_60,In_97);
or U1392 (N_1392,In_1067,In_69);
and U1393 (N_1393,In_971,In_50);
nor U1394 (N_1394,In_1417,In_837);
nand U1395 (N_1395,In_460,In_39);
and U1396 (N_1396,In_114,In_1394);
xor U1397 (N_1397,In_544,In_1340);
nor U1398 (N_1398,In_418,In_162);
xor U1399 (N_1399,In_940,In_577);
or U1400 (N_1400,In_1237,In_392);
and U1401 (N_1401,In_237,In_437);
or U1402 (N_1402,In_1408,In_399);
nand U1403 (N_1403,In_21,In_814);
or U1404 (N_1404,In_874,In_1001);
nand U1405 (N_1405,In_315,In_128);
nor U1406 (N_1406,In_1350,In_935);
nand U1407 (N_1407,In_663,In_1460);
nor U1408 (N_1408,In_935,In_743);
and U1409 (N_1409,In_281,In_294);
xor U1410 (N_1410,In_838,In_1232);
xnor U1411 (N_1411,In_1126,In_508);
xor U1412 (N_1412,In_215,In_688);
or U1413 (N_1413,In_1370,In_1001);
nor U1414 (N_1414,In_541,In_772);
or U1415 (N_1415,In_1263,In_643);
nand U1416 (N_1416,In_452,In_1434);
or U1417 (N_1417,In_1218,In_381);
or U1418 (N_1418,In_876,In_476);
xnor U1419 (N_1419,In_510,In_70);
or U1420 (N_1420,In_508,In_577);
xnor U1421 (N_1421,In_1315,In_42);
nand U1422 (N_1422,In_449,In_1153);
or U1423 (N_1423,In_142,In_24);
or U1424 (N_1424,In_997,In_291);
and U1425 (N_1425,In_394,In_1108);
xnor U1426 (N_1426,In_1283,In_569);
xor U1427 (N_1427,In_1242,In_377);
nor U1428 (N_1428,In_1052,In_274);
nand U1429 (N_1429,In_789,In_1079);
or U1430 (N_1430,In_187,In_870);
nand U1431 (N_1431,In_688,In_472);
xor U1432 (N_1432,In_1461,In_119);
nand U1433 (N_1433,In_1246,In_33);
nand U1434 (N_1434,In_508,In_1317);
and U1435 (N_1435,In_978,In_79);
xnor U1436 (N_1436,In_989,In_423);
or U1437 (N_1437,In_531,In_616);
nand U1438 (N_1438,In_372,In_281);
nor U1439 (N_1439,In_162,In_360);
xnor U1440 (N_1440,In_1447,In_1087);
or U1441 (N_1441,In_800,In_604);
nand U1442 (N_1442,In_961,In_1485);
xor U1443 (N_1443,In_196,In_728);
nor U1444 (N_1444,In_839,In_585);
nor U1445 (N_1445,In_169,In_1182);
and U1446 (N_1446,In_1251,In_257);
or U1447 (N_1447,In_297,In_1494);
and U1448 (N_1448,In_180,In_511);
nor U1449 (N_1449,In_637,In_259);
nor U1450 (N_1450,In_567,In_19);
and U1451 (N_1451,In_625,In_146);
and U1452 (N_1452,In_840,In_332);
nand U1453 (N_1453,In_1428,In_744);
and U1454 (N_1454,In_772,In_406);
nand U1455 (N_1455,In_658,In_212);
nor U1456 (N_1456,In_156,In_518);
or U1457 (N_1457,In_1268,In_923);
or U1458 (N_1458,In_1088,In_399);
and U1459 (N_1459,In_363,In_1187);
nand U1460 (N_1460,In_1202,In_903);
or U1461 (N_1461,In_284,In_213);
nor U1462 (N_1462,In_951,In_1270);
or U1463 (N_1463,In_732,In_81);
and U1464 (N_1464,In_1258,In_1108);
nand U1465 (N_1465,In_862,In_1137);
or U1466 (N_1466,In_643,In_296);
nand U1467 (N_1467,In_414,In_458);
xnor U1468 (N_1468,In_874,In_181);
and U1469 (N_1469,In_1079,In_44);
and U1470 (N_1470,In_629,In_728);
nand U1471 (N_1471,In_949,In_1413);
or U1472 (N_1472,In_1233,In_1245);
nor U1473 (N_1473,In_1050,In_320);
xnor U1474 (N_1474,In_756,In_473);
and U1475 (N_1475,In_1322,In_17);
nor U1476 (N_1476,In_668,In_766);
nand U1477 (N_1477,In_728,In_1057);
nor U1478 (N_1478,In_808,In_1268);
nor U1479 (N_1479,In_682,In_27);
xor U1480 (N_1480,In_1483,In_922);
or U1481 (N_1481,In_539,In_419);
or U1482 (N_1482,In_1146,In_481);
xor U1483 (N_1483,In_1151,In_967);
nor U1484 (N_1484,In_529,In_633);
or U1485 (N_1485,In_151,In_593);
nand U1486 (N_1486,In_324,In_444);
xor U1487 (N_1487,In_524,In_508);
xnor U1488 (N_1488,In_228,In_859);
xnor U1489 (N_1489,In_1213,In_462);
and U1490 (N_1490,In_432,In_771);
nor U1491 (N_1491,In_1243,In_246);
or U1492 (N_1492,In_750,In_1034);
and U1493 (N_1493,In_1381,In_1420);
nand U1494 (N_1494,In_141,In_148);
or U1495 (N_1495,In_1179,In_200);
xnor U1496 (N_1496,In_890,In_413);
or U1497 (N_1497,In_1276,In_1188);
xnor U1498 (N_1498,In_1466,In_1002);
nor U1499 (N_1499,In_1345,In_146);
nand U1500 (N_1500,In_1367,In_1166);
xnor U1501 (N_1501,In_471,In_132);
xor U1502 (N_1502,In_800,In_284);
and U1503 (N_1503,In_729,In_1300);
or U1504 (N_1504,In_969,In_740);
nand U1505 (N_1505,In_229,In_606);
and U1506 (N_1506,In_707,In_1484);
xnor U1507 (N_1507,In_379,In_1310);
and U1508 (N_1508,In_1102,In_1283);
or U1509 (N_1509,In_7,In_529);
or U1510 (N_1510,In_987,In_792);
or U1511 (N_1511,In_140,In_1252);
nor U1512 (N_1512,In_1098,In_787);
nand U1513 (N_1513,In_1387,In_1020);
and U1514 (N_1514,In_1376,In_547);
xor U1515 (N_1515,In_1234,In_149);
nor U1516 (N_1516,In_1182,In_699);
and U1517 (N_1517,In_657,In_38);
nand U1518 (N_1518,In_260,In_41);
or U1519 (N_1519,In_656,In_857);
nand U1520 (N_1520,In_1049,In_1272);
nor U1521 (N_1521,In_796,In_1444);
or U1522 (N_1522,In_1465,In_355);
xnor U1523 (N_1523,In_1186,In_58);
or U1524 (N_1524,In_563,In_1139);
or U1525 (N_1525,In_565,In_1119);
or U1526 (N_1526,In_1240,In_968);
xor U1527 (N_1527,In_180,In_1030);
xnor U1528 (N_1528,In_390,In_341);
or U1529 (N_1529,In_61,In_1141);
xnor U1530 (N_1530,In_766,In_578);
nor U1531 (N_1531,In_1085,In_223);
xor U1532 (N_1532,In_1357,In_174);
or U1533 (N_1533,In_1231,In_1246);
xnor U1534 (N_1534,In_234,In_279);
nor U1535 (N_1535,In_1073,In_19);
nand U1536 (N_1536,In_183,In_493);
xor U1537 (N_1537,In_1294,In_502);
nor U1538 (N_1538,In_866,In_1477);
or U1539 (N_1539,In_1291,In_650);
nand U1540 (N_1540,In_573,In_818);
nand U1541 (N_1541,In_706,In_1342);
and U1542 (N_1542,In_638,In_1253);
xnor U1543 (N_1543,In_900,In_876);
and U1544 (N_1544,In_1384,In_265);
nand U1545 (N_1545,In_1186,In_1171);
or U1546 (N_1546,In_991,In_277);
nand U1547 (N_1547,In_15,In_1085);
nor U1548 (N_1548,In_129,In_12);
and U1549 (N_1549,In_364,In_112);
or U1550 (N_1550,In_1355,In_1362);
or U1551 (N_1551,In_408,In_618);
and U1552 (N_1552,In_748,In_1282);
xnor U1553 (N_1553,In_450,In_728);
or U1554 (N_1554,In_1000,In_625);
or U1555 (N_1555,In_970,In_1018);
nand U1556 (N_1556,In_1,In_1351);
nand U1557 (N_1557,In_488,In_1371);
or U1558 (N_1558,In_564,In_454);
nor U1559 (N_1559,In_730,In_1369);
nor U1560 (N_1560,In_870,In_910);
and U1561 (N_1561,In_989,In_1176);
nor U1562 (N_1562,In_1027,In_861);
or U1563 (N_1563,In_447,In_586);
nor U1564 (N_1564,In_958,In_397);
or U1565 (N_1565,In_1398,In_950);
xnor U1566 (N_1566,In_1044,In_1161);
xor U1567 (N_1567,In_586,In_1368);
nand U1568 (N_1568,In_1255,In_1164);
nor U1569 (N_1569,In_1358,In_893);
nor U1570 (N_1570,In_715,In_414);
xnor U1571 (N_1571,In_169,In_660);
nand U1572 (N_1572,In_1293,In_500);
nor U1573 (N_1573,In_145,In_377);
and U1574 (N_1574,In_375,In_643);
xor U1575 (N_1575,In_268,In_1272);
xnor U1576 (N_1576,In_844,In_1192);
xnor U1577 (N_1577,In_717,In_260);
xor U1578 (N_1578,In_1125,In_1262);
xnor U1579 (N_1579,In_48,In_86);
and U1580 (N_1580,In_438,In_419);
xnor U1581 (N_1581,In_954,In_856);
nand U1582 (N_1582,In_744,In_29);
nor U1583 (N_1583,In_324,In_1216);
or U1584 (N_1584,In_936,In_103);
xnor U1585 (N_1585,In_1485,In_165);
and U1586 (N_1586,In_183,In_1394);
and U1587 (N_1587,In_1044,In_798);
xnor U1588 (N_1588,In_633,In_280);
nor U1589 (N_1589,In_193,In_730);
xnor U1590 (N_1590,In_755,In_1440);
nand U1591 (N_1591,In_91,In_1378);
xor U1592 (N_1592,In_1144,In_390);
nand U1593 (N_1593,In_683,In_1091);
or U1594 (N_1594,In_922,In_677);
nor U1595 (N_1595,In_302,In_1217);
or U1596 (N_1596,In_1011,In_326);
xor U1597 (N_1597,In_253,In_321);
or U1598 (N_1598,In_1279,In_337);
xor U1599 (N_1599,In_493,In_992);
and U1600 (N_1600,In_1222,In_314);
and U1601 (N_1601,In_1387,In_1458);
xor U1602 (N_1602,In_162,In_860);
nand U1603 (N_1603,In_437,In_347);
nor U1604 (N_1604,In_1160,In_927);
and U1605 (N_1605,In_625,In_606);
or U1606 (N_1606,In_1406,In_628);
nand U1607 (N_1607,In_422,In_1057);
and U1608 (N_1608,In_620,In_501);
nand U1609 (N_1609,In_982,In_1116);
or U1610 (N_1610,In_1110,In_815);
and U1611 (N_1611,In_228,In_1394);
nand U1612 (N_1612,In_1190,In_852);
xnor U1613 (N_1613,In_1007,In_276);
and U1614 (N_1614,In_1300,In_836);
nand U1615 (N_1615,In_298,In_516);
and U1616 (N_1616,In_775,In_1122);
or U1617 (N_1617,In_101,In_420);
nand U1618 (N_1618,In_1476,In_605);
or U1619 (N_1619,In_595,In_1493);
or U1620 (N_1620,In_131,In_1179);
nand U1621 (N_1621,In_1185,In_82);
nor U1622 (N_1622,In_408,In_916);
nand U1623 (N_1623,In_1076,In_1495);
nand U1624 (N_1624,In_913,In_1371);
nor U1625 (N_1625,In_573,In_400);
nand U1626 (N_1626,In_340,In_377);
nor U1627 (N_1627,In_664,In_596);
nor U1628 (N_1628,In_250,In_983);
xor U1629 (N_1629,In_378,In_582);
nor U1630 (N_1630,In_349,In_506);
nor U1631 (N_1631,In_1363,In_865);
or U1632 (N_1632,In_1131,In_147);
nand U1633 (N_1633,In_1402,In_733);
xor U1634 (N_1634,In_1034,In_850);
and U1635 (N_1635,In_1067,In_1188);
nand U1636 (N_1636,In_228,In_927);
nor U1637 (N_1637,In_1057,In_1426);
and U1638 (N_1638,In_990,In_41);
and U1639 (N_1639,In_1120,In_1305);
nand U1640 (N_1640,In_1482,In_971);
nand U1641 (N_1641,In_1040,In_864);
or U1642 (N_1642,In_259,In_419);
or U1643 (N_1643,In_581,In_247);
nor U1644 (N_1644,In_448,In_505);
xor U1645 (N_1645,In_356,In_1018);
nor U1646 (N_1646,In_666,In_1483);
xnor U1647 (N_1647,In_979,In_1347);
and U1648 (N_1648,In_893,In_1472);
or U1649 (N_1649,In_836,In_1232);
xor U1650 (N_1650,In_10,In_1272);
nand U1651 (N_1651,In_400,In_186);
nand U1652 (N_1652,In_808,In_1096);
nand U1653 (N_1653,In_496,In_1441);
nand U1654 (N_1654,In_860,In_897);
and U1655 (N_1655,In_815,In_441);
nand U1656 (N_1656,In_692,In_565);
nand U1657 (N_1657,In_672,In_25);
nand U1658 (N_1658,In_466,In_128);
nor U1659 (N_1659,In_1123,In_826);
nand U1660 (N_1660,In_493,In_1155);
xor U1661 (N_1661,In_1208,In_31);
nand U1662 (N_1662,In_819,In_167);
nand U1663 (N_1663,In_1411,In_1003);
nor U1664 (N_1664,In_1370,In_883);
nor U1665 (N_1665,In_1043,In_628);
xnor U1666 (N_1666,In_1425,In_1372);
xor U1667 (N_1667,In_819,In_307);
and U1668 (N_1668,In_205,In_120);
or U1669 (N_1669,In_137,In_942);
xor U1670 (N_1670,In_166,In_820);
nor U1671 (N_1671,In_657,In_41);
or U1672 (N_1672,In_517,In_1360);
and U1673 (N_1673,In_276,In_1427);
and U1674 (N_1674,In_19,In_137);
nand U1675 (N_1675,In_1380,In_287);
nand U1676 (N_1676,In_448,In_1235);
and U1677 (N_1677,In_1279,In_966);
or U1678 (N_1678,In_1110,In_1306);
and U1679 (N_1679,In_734,In_64);
nor U1680 (N_1680,In_719,In_1330);
nor U1681 (N_1681,In_1385,In_1295);
or U1682 (N_1682,In_157,In_1067);
or U1683 (N_1683,In_1118,In_300);
xor U1684 (N_1684,In_617,In_544);
xor U1685 (N_1685,In_814,In_541);
and U1686 (N_1686,In_1236,In_1165);
nand U1687 (N_1687,In_561,In_875);
xnor U1688 (N_1688,In_145,In_739);
or U1689 (N_1689,In_514,In_776);
nor U1690 (N_1690,In_852,In_742);
or U1691 (N_1691,In_806,In_1334);
nand U1692 (N_1692,In_288,In_644);
xor U1693 (N_1693,In_937,In_370);
nor U1694 (N_1694,In_1316,In_1128);
nand U1695 (N_1695,In_1062,In_526);
nand U1696 (N_1696,In_1016,In_514);
and U1697 (N_1697,In_845,In_735);
or U1698 (N_1698,In_218,In_729);
xor U1699 (N_1699,In_1018,In_979);
and U1700 (N_1700,In_670,In_308);
and U1701 (N_1701,In_1305,In_1048);
and U1702 (N_1702,In_1061,In_485);
and U1703 (N_1703,In_1198,In_239);
xor U1704 (N_1704,In_1090,In_615);
or U1705 (N_1705,In_541,In_1441);
and U1706 (N_1706,In_85,In_151);
nand U1707 (N_1707,In_1029,In_129);
and U1708 (N_1708,In_215,In_700);
nand U1709 (N_1709,In_649,In_353);
nor U1710 (N_1710,In_1366,In_100);
nand U1711 (N_1711,In_779,In_1137);
and U1712 (N_1712,In_1465,In_1472);
and U1713 (N_1713,In_225,In_729);
nor U1714 (N_1714,In_922,In_949);
or U1715 (N_1715,In_1218,In_904);
nor U1716 (N_1716,In_100,In_134);
nand U1717 (N_1717,In_737,In_328);
or U1718 (N_1718,In_899,In_44);
nor U1719 (N_1719,In_1262,In_226);
xor U1720 (N_1720,In_978,In_85);
nand U1721 (N_1721,In_390,In_1401);
nand U1722 (N_1722,In_1250,In_1384);
nand U1723 (N_1723,In_455,In_1242);
and U1724 (N_1724,In_1494,In_816);
nor U1725 (N_1725,In_515,In_524);
xnor U1726 (N_1726,In_169,In_529);
and U1727 (N_1727,In_710,In_53);
nor U1728 (N_1728,In_1438,In_731);
nand U1729 (N_1729,In_255,In_667);
nor U1730 (N_1730,In_1123,In_360);
nor U1731 (N_1731,In_1093,In_1171);
nand U1732 (N_1732,In_1324,In_1022);
nand U1733 (N_1733,In_585,In_1499);
or U1734 (N_1734,In_492,In_1317);
or U1735 (N_1735,In_530,In_763);
or U1736 (N_1736,In_662,In_754);
and U1737 (N_1737,In_431,In_298);
or U1738 (N_1738,In_856,In_1122);
nand U1739 (N_1739,In_199,In_301);
nand U1740 (N_1740,In_330,In_171);
nor U1741 (N_1741,In_840,In_846);
nor U1742 (N_1742,In_559,In_1380);
or U1743 (N_1743,In_1229,In_570);
and U1744 (N_1744,In_294,In_595);
nand U1745 (N_1745,In_1228,In_1483);
nor U1746 (N_1746,In_1123,In_857);
nor U1747 (N_1747,In_409,In_2);
and U1748 (N_1748,In_829,In_990);
or U1749 (N_1749,In_1044,In_823);
xnor U1750 (N_1750,In_1228,In_14);
and U1751 (N_1751,In_1493,In_1155);
nand U1752 (N_1752,In_1123,In_1109);
nor U1753 (N_1753,In_451,In_994);
or U1754 (N_1754,In_1279,In_148);
nand U1755 (N_1755,In_389,In_992);
xnor U1756 (N_1756,In_821,In_999);
or U1757 (N_1757,In_1449,In_793);
nor U1758 (N_1758,In_881,In_1212);
or U1759 (N_1759,In_566,In_585);
xnor U1760 (N_1760,In_74,In_1411);
xor U1761 (N_1761,In_744,In_295);
nand U1762 (N_1762,In_126,In_802);
and U1763 (N_1763,In_125,In_1077);
or U1764 (N_1764,In_626,In_607);
or U1765 (N_1765,In_1475,In_797);
nand U1766 (N_1766,In_733,In_624);
xor U1767 (N_1767,In_786,In_511);
nand U1768 (N_1768,In_1305,In_231);
or U1769 (N_1769,In_868,In_701);
nand U1770 (N_1770,In_184,In_19);
nand U1771 (N_1771,In_487,In_192);
or U1772 (N_1772,In_1314,In_56);
nor U1773 (N_1773,In_180,In_525);
or U1774 (N_1774,In_1364,In_671);
xor U1775 (N_1775,In_1173,In_474);
and U1776 (N_1776,In_1286,In_166);
nor U1777 (N_1777,In_1366,In_509);
xor U1778 (N_1778,In_372,In_889);
xor U1779 (N_1779,In_820,In_1262);
nand U1780 (N_1780,In_1216,In_436);
nand U1781 (N_1781,In_527,In_1241);
xnor U1782 (N_1782,In_1300,In_1262);
and U1783 (N_1783,In_509,In_1098);
xnor U1784 (N_1784,In_681,In_1244);
xnor U1785 (N_1785,In_110,In_500);
nor U1786 (N_1786,In_585,In_1484);
xnor U1787 (N_1787,In_1353,In_1073);
xor U1788 (N_1788,In_1010,In_1108);
and U1789 (N_1789,In_1224,In_1447);
and U1790 (N_1790,In_1225,In_403);
nand U1791 (N_1791,In_639,In_505);
and U1792 (N_1792,In_1491,In_769);
nand U1793 (N_1793,In_214,In_188);
nand U1794 (N_1794,In_1451,In_1079);
xnor U1795 (N_1795,In_1126,In_1250);
and U1796 (N_1796,In_365,In_828);
or U1797 (N_1797,In_895,In_1086);
nor U1798 (N_1798,In_1064,In_1499);
xnor U1799 (N_1799,In_354,In_1103);
xnor U1800 (N_1800,In_328,In_80);
or U1801 (N_1801,In_28,In_793);
and U1802 (N_1802,In_1395,In_129);
nand U1803 (N_1803,In_945,In_863);
nand U1804 (N_1804,In_664,In_987);
nand U1805 (N_1805,In_997,In_1096);
and U1806 (N_1806,In_1331,In_581);
or U1807 (N_1807,In_67,In_445);
nand U1808 (N_1808,In_1477,In_625);
nand U1809 (N_1809,In_958,In_622);
nor U1810 (N_1810,In_931,In_78);
and U1811 (N_1811,In_977,In_442);
nand U1812 (N_1812,In_216,In_1090);
nor U1813 (N_1813,In_94,In_46);
and U1814 (N_1814,In_491,In_1254);
nor U1815 (N_1815,In_427,In_1368);
nor U1816 (N_1816,In_1356,In_1055);
nor U1817 (N_1817,In_940,In_1056);
nand U1818 (N_1818,In_504,In_58);
nor U1819 (N_1819,In_420,In_975);
or U1820 (N_1820,In_752,In_377);
or U1821 (N_1821,In_1016,In_242);
and U1822 (N_1822,In_1173,In_1067);
and U1823 (N_1823,In_906,In_421);
and U1824 (N_1824,In_432,In_1255);
nor U1825 (N_1825,In_164,In_695);
and U1826 (N_1826,In_508,In_549);
nor U1827 (N_1827,In_881,In_1194);
and U1828 (N_1828,In_303,In_1059);
and U1829 (N_1829,In_856,In_549);
xor U1830 (N_1830,In_193,In_508);
nor U1831 (N_1831,In_1225,In_665);
nand U1832 (N_1832,In_673,In_1106);
or U1833 (N_1833,In_1424,In_1263);
or U1834 (N_1834,In_145,In_271);
nand U1835 (N_1835,In_1041,In_428);
nand U1836 (N_1836,In_679,In_1067);
or U1837 (N_1837,In_890,In_21);
or U1838 (N_1838,In_634,In_1086);
nor U1839 (N_1839,In_506,In_1367);
xor U1840 (N_1840,In_460,In_831);
or U1841 (N_1841,In_736,In_1328);
or U1842 (N_1842,In_1139,In_1371);
xnor U1843 (N_1843,In_1293,In_596);
xnor U1844 (N_1844,In_1100,In_391);
or U1845 (N_1845,In_1154,In_1130);
nand U1846 (N_1846,In_83,In_1231);
and U1847 (N_1847,In_495,In_134);
nor U1848 (N_1848,In_955,In_1419);
nand U1849 (N_1849,In_1208,In_1245);
nand U1850 (N_1850,In_1028,In_1049);
nand U1851 (N_1851,In_1140,In_1440);
and U1852 (N_1852,In_711,In_208);
nand U1853 (N_1853,In_1065,In_1005);
xnor U1854 (N_1854,In_459,In_201);
xor U1855 (N_1855,In_147,In_607);
nor U1856 (N_1856,In_337,In_85);
nor U1857 (N_1857,In_284,In_1371);
or U1858 (N_1858,In_821,In_896);
and U1859 (N_1859,In_993,In_1008);
or U1860 (N_1860,In_837,In_623);
nor U1861 (N_1861,In_377,In_1420);
nor U1862 (N_1862,In_151,In_1196);
xnor U1863 (N_1863,In_470,In_144);
nand U1864 (N_1864,In_280,In_345);
and U1865 (N_1865,In_499,In_1179);
xor U1866 (N_1866,In_118,In_192);
or U1867 (N_1867,In_449,In_197);
nand U1868 (N_1868,In_584,In_83);
xnor U1869 (N_1869,In_1344,In_1138);
or U1870 (N_1870,In_1139,In_364);
xor U1871 (N_1871,In_524,In_1479);
nor U1872 (N_1872,In_1320,In_1327);
xnor U1873 (N_1873,In_223,In_1479);
or U1874 (N_1874,In_385,In_628);
xnor U1875 (N_1875,In_988,In_1100);
or U1876 (N_1876,In_371,In_1123);
xor U1877 (N_1877,In_1212,In_407);
or U1878 (N_1878,In_1294,In_1028);
and U1879 (N_1879,In_961,In_272);
xnor U1880 (N_1880,In_275,In_1354);
and U1881 (N_1881,In_360,In_958);
and U1882 (N_1882,In_1347,In_333);
nand U1883 (N_1883,In_1011,In_793);
and U1884 (N_1884,In_1326,In_985);
xnor U1885 (N_1885,In_1463,In_1329);
nor U1886 (N_1886,In_13,In_1148);
or U1887 (N_1887,In_605,In_55);
or U1888 (N_1888,In_1277,In_818);
xor U1889 (N_1889,In_827,In_1249);
or U1890 (N_1890,In_107,In_490);
xnor U1891 (N_1891,In_619,In_150);
or U1892 (N_1892,In_1282,In_1299);
or U1893 (N_1893,In_46,In_1019);
and U1894 (N_1894,In_1298,In_1067);
and U1895 (N_1895,In_1154,In_6);
nor U1896 (N_1896,In_292,In_350);
nor U1897 (N_1897,In_482,In_1385);
xor U1898 (N_1898,In_120,In_73);
and U1899 (N_1899,In_1115,In_734);
nand U1900 (N_1900,In_1144,In_657);
or U1901 (N_1901,In_1297,In_321);
and U1902 (N_1902,In_204,In_512);
nand U1903 (N_1903,In_1335,In_1076);
xor U1904 (N_1904,In_307,In_1003);
or U1905 (N_1905,In_887,In_862);
nand U1906 (N_1906,In_1360,In_925);
nand U1907 (N_1907,In_266,In_286);
nand U1908 (N_1908,In_303,In_1155);
nor U1909 (N_1909,In_1431,In_548);
or U1910 (N_1910,In_219,In_664);
and U1911 (N_1911,In_1271,In_440);
nand U1912 (N_1912,In_503,In_729);
xnor U1913 (N_1913,In_960,In_1);
nand U1914 (N_1914,In_1313,In_116);
nand U1915 (N_1915,In_621,In_904);
nor U1916 (N_1916,In_1070,In_213);
nor U1917 (N_1917,In_1006,In_1240);
nor U1918 (N_1918,In_1372,In_1225);
and U1919 (N_1919,In_936,In_1137);
xor U1920 (N_1920,In_170,In_109);
and U1921 (N_1921,In_691,In_283);
nor U1922 (N_1922,In_677,In_866);
nand U1923 (N_1923,In_708,In_1441);
nor U1924 (N_1924,In_888,In_1485);
xnor U1925 (N_1925,In_957,In_880);
and U1926 (N_1926,In_1116,In_363);
and U1927 (N_1927,In_123,In_742);
xnor U1928 (N_1928,In_96,In_171);
and U1929 (N_1929,In_1355,In_111);
and U1930 (N_1930,In_229,In_800);
nor U1931 (N_1931,In_1271,In_99);
and U1932 (N_1932,In_496,In_105);
or U1933 (N_1933,In_1030,In_119);
or U1934 (N_1934,In_288,In_932);
or U1935 (N_1935,In_784,In_102);
and U1936 (N_1936,In_195,In_176);
or U1937 (N_1937,In_239,In_105);
and U1938 (N_1938,In_379,In_285);
and U1939 (N_1939,In_1404,In_1142);
nor U1940 (N_1940,In_97,In_695);
nor U1941 (N_1941,In_1091,In_219);
nand U1942 (N_1942,In_428,In_661);
nand U1943 (N_1943,In_195,In_529);
or U1944 (N_1944,In_487,In_1420);
or U1945 (N_1945,In_492,In_810);
xor U1946 (N_1946,In_1420,In_662);
or U1947 (N_1947,In_273,In_692);
and U1948 (N_1948,In_944,In_995);
xor U1949 (N_1949,In_522,In_1229);
or U1950 (N_1950,In_522,In_302);
and U1951 (N_1951,In_867,In_987);
nand U1952 (N_1952,In_274,In_345);
nor U1953 (N_1953,In_880,In_113);
nand U1954 (N_1954,In_421,In_1487);
or U1955 (N_1955,In_196,In_319);
or U1956 (N_1956,In_540,In_776);
xor U1957 (N_1957,In_1011,In_299);
or U1958 (N_1958,In_1022,In_1002);
or U1959 (N_1959,In_240,In_334);
xnor U1960 (N_1960,In_802,In_1313);
nand U1961 (N_1961,In_1019,In_611);
or U1962 (N_1962,In_688,In_15);
and U1963 (N_1963,In_428,In_681);
and U1964 (N_1964,In_1136,In_906);
xor U1965 (N_1965,In_102,In_320);
or U1966 (N_1966,In_133,In_1029);
nand U1967 (N_1967,In_1095,In_139);
nand U1968 (N_1968,In_555,In_937);
nor U1969 (N_1969,In_1066,In_728);
nor U1970 (N_1970,In_759,In_971);
and U1971 (N_1971,In_266,In_892);
nand U1972 (N_1972,In_1040,In_590);
nand U1973 (N_1973,In_515,In_574);
or U1974 (N_1974,In_120,In_192);
nand U1975 (N_1975,In_1296,In_119);
nor U1976 (N_1976,In_1390,In_803);
nor U1977 (N_1977,In_1032,In_317);
xnor U1978 (N_1978,In_1025,In_689);
nand U1979 (N_1979,In_1191,In_878);
or U1980 (N_1980,In_307,In_899);
nor U1981 (N_1981,In_1314,In_741);
xnor U1982 (N_1982,In_995,In_1155);
and U1983 (N_1983,In_1366,In_538);
xor U1984 (N_1984,In_1040,In_1385);
xor U1985 (N_1985,In_1413,In_1161);
nand U1986 (N_1986,In_183,In_1379);
xor U1987 (N_1987,In_402,In_3);
nor U1988 (N_1988,In_637,In_243);
xnor U1989 (N_1989,In_1398,In_81);
nor U1990 (N_1990,In_1286,In_983);
xor U1991 (N_1991,In_818,In_1274);
nand U1992 (N_1992,In_1370,In_659);
nand U1993 (N_1993,In_1342,In_210);
or U1994 (N_1994,In_819,In_1295);
and U1995 (N_1995,In_1405,In_622);
nand U1996 (N_1996,In_1204,In_565);
xor U1997 (N_1997,In_92,In_978);
nand U1998 (N_1998,In_1046,In_1134);
or U1999 (N_1999,In_1437,In_667);
nand U2000 (N_2000,In_1475,In_834);
or U2001 (N_2001,In_662,In_460);
and U2002 (N_2002,In_1100,In_1487);
nor U2003 (N_2003,In_623,In_1377);
or U2004 (N_2004,In_396,In_516);
or U2005 (N_2005,In_1191,In_706);
nand U2006 (N_2006,In_1336,In_340);
nand U2007 (N_2007,In_1239,In_289);
nor U2008 (N_2008,In_1301,In_1391);
xnor U2009 (N_2009,In_622,In_909);
and U2010 (N_2010,In_1190,In_1428);
nor U2011 (N_2011,In_1116,In_546);
or U2012 (N_2012,In_705,In_943);
nand U2013 (N_2013,In_129,In_1223);
xor U2014 (N_2014,In_1234,In_187);
and U2015 (N_2015,In_72,In_1288);
nand U2016 (N_2016,In_151,In_953);
and U2017 (N_2017,In_713,In_977);
and U2018 (N_2018,In_1326,In_815);
nand U2019 (N_2019,In_288,In_161);
xnor U2020 (N_2020,In_615,In_415);
xor U2021 (N_2021,In_1027,In_13);
xnor U2022 (N_2022,In_712,In_1331);
xnor U2023 (N_2023,In_1313,In_196);
nand U2024 (N_2024,In_762,In_872);
nor U2025 (N_2025,In_500,In_860);
nor U2026 (N_2026,In_461,In_677);
or U2027 (N_2027,In_1272,In_1150);
xor U2028 (N_2028,In_93,In_537);
or U2029 (N_2029,In_1,In_180);
nand U2030 (N_2030,In_1100,In_473);
or U2031 (N_2031,In_845,In_758);
or U2032 (N_2032,In_836,In_864);
xnor U2033 (N_2033,In_285,In_1059);
xnor U2034 (N_2034,In_878,In_199);
nand U2035 (N_2035,In_310,In_17);
nor U2036 (N_2036,In_643,In_676);
nor U2037 (N_2037,In_992,In_964);
nand U2038 (N_2038,In_448,In_1103);
nor U2039 (N_2039,In_1337,In_806);
nor U2040 (N_2040,In_554,In_626);
nand U2041 (N_2041,In_333,In_655);
nand U2042 (N_2042,In_235,In_639);
or U2043 (N_2043,In_291,In_686);
or U2044 (N_2044,In_302,In_97);
nor U2045 (N_2045,In_972,In_298);
or U2046 (N_2046,In_271,In_897);
nand U2047 (N_2047,In_1352,In_353);
nor U2048 (N_2048,In_124,In_1350);
and U2049 (N_2049,In_33,In_1391);
xnor U2050 (N_2050,In_50,In_1338);
or U2051 (N_2051,In_1090,In_725);
nand U2052 (N_2052,In_902,In_1424);
nand U2053 (N_2053,In_88,In_237);
and U2054 (N_2054,In_293,In_760);
and U2055 (N_2055,In_184,In_1136);
nand U2056 (N_2056,In_1424,In_176);
nor U2057 (N_2057,In_473,In_515);
and U2058 (N_2058,In_1490,In_1209);
xor U2059 (N_2059,In_344,In_524);
nand U2060 (N_2060,In_813,In_978);
or U2061 (N_2061,In_31,In_475);
nor U2062 (N_2062,In_736,In_880);
xor U2063 (N_2063,In_1309,In_504);
or U2064 (N_2064,In_990,In_858);
or U2065 (N_2065,In_1359,In_738);
nor U2066 (N_2066,In_1103,In_1434);
xor U2067 (N_2067,In_1473,In_255);
nor U2068 (N_2068,In_1228,In_908);
nor U2069 (N_2069,In_364,In_194);
nor U2070 (N_2070,In_144,In_773);
and U2071 (N_2071,In_263,In_941);
xor U2072 (N_2072,In_1456,In_1054);
nor U2073 (N_2073,In_508,In_726);
xnor U2074 (N_2074,In_112,In_666);
and U2075 (N_2075,In_863,In_718);
and U2076 (N_2076,In_1073,In_325);
nand U2077 (N_2077,In_190,In_175);
nor U2078 (N_2078,In_684,In_1269);
nand U2079 (N_2079,In_739,In_284);
xnor U2080 (N_2080,In_572,In_921);
nand U2081 (N_2081,In_936,In_320);
and U2082 (N_2082,In_31,In_1345);
and U2083 (N_2083,In_767,In_1418);
nor U2084 (N_2084,In_1020,In_715);
xor U2085 (N_2085,In_733,In_589);
xor U2086 (N_2086,In_1190,In_1167);
xnor U2087 (N_2087,In_569,In_1050);
nor U2088 (N_2088,In_925,In_937);
or U2089 (N_2089,In_921,In_873);
nand U2090 (N_2090,In_46,In_752);
xnor U2091 (N_2091,In_220,In_1375);
xor U2092 (N_2092,In_1368,In_976);
and U2093 (N_2093,In_678,In_1206);
xor U2094 (N_2094,In_128,In_291);
nand U2095 (N_2095,In_1434,In_688);
and U2096 (N_2096,In_380,In_510);
xnor U2097 (N_2097,In_263,In_314);
or U2098 (N_2098,In_1356,In_963);
xor U2099 (N_2099,In_483,In_489);
nor U2100 (N_2100,In_582,In_1061);
nand U2101 (N_2101,In_1425,In_1410);
xnor U2102 (N_2102,In_1150,In_611);
or U2103 (N_2103,In_26,In_724);
and U2104 (N_2104,In_87,In_616);
and U2105 (N_2105,In_788,In_1267);
or U2106 (N_2106,In_208,In_966);
nor U2107 (N_2107,In_330,In_853);
and U2108 (N_2108,In_467,In_713);
xnor U2109 (N_2109,In_57,In_896);
or U2110 (N_2110,In_899,In_191);
xnor U2111 (N_2111,In_1372,In_1298);
nor U2112 (N_2112,In_1019,In_955);
xnor U2113 (N_2113,In_314,In_134);
nor U2114 (N_2114,In_1019,In_427);
or U2115 (N_2115,In_1199,In_1337);
xnor U2116 (N_2116,In_1243,In_1034);
xor U2117 (N_2117,In_448,In_938);
nand U2118 (N_2118,In_1018,In_478);
nor U2119 (N_2119,In_65,In_210);
nand U2120 (N_2120,In_196,In_23);
or U2121 (N_2121,In_1406,In_1244);
nand U2122 (N_2122,In_368,In_344);
and U2123 (N_2123,In_449,In_1444);
xor U2124 (N_2124,In_292,In_710);
nor U2125 (N_2125,In_792,In_731);
nor U2126 (N_2126,In_1189,In_474);
nor U2127 (N_2127,In_1035,In_1450);
and U2128 (N_2128,In_608,In_1024);
nand U2129 (N_2129,In_819,In_968);
xor U2130 (N_2130,In_1295,In_172);
xnor U2131 (N_2131,In_261,In_288);
and U2132 (N_2132,In_809,In_535);
or U2133 (N_2133,In_102,In_394);
and U2134 (N_2134,In_77,In_1058);
and U2135 (N_2135,In_107,In_709);
xor U2136 (N_2136,In_377,In_48);
nor U2137 (N_2137,In_255,In_412);
or U2138 (N_2138,In_587,In_913);
nand U2139 (N_2139,In_1465,In_813);
xor U2140 (N_2140,In_258,In_1226);
or U2141 (N_2141,In_1340,In_1387);
nor U2142 (N_2142,In_902,In_1364);
nor U2143 (N_2143,In_546,In_1308);
nor U2144 (N_2144,In_1341,In_311);
nor U2145 (N_2145,In_293,In_257);
or U2146 (N_2146,In_1386,In_1069);
and U2147 (N_2147,In_391,In_1057);
nand U2148 (N_2148,In_42,In_623);
or U2149 (N_2149,In_1482,In_1078);
and U2150 (N_2150,In_1019,In_1098);
nor U2151 (N_2151,In_995,In_467);
and U2152 (N_2152,In_809,In_1393);
and U2153 (N_2153,In_1020,In_909);
nand U2154 (N_2154,In_706,In_657);
nor U2155 (N_2155,In_364,In_805);
or U2156 (N_2156,In_670,In_100);
nand U2157 (N_2157,In_730,In_708);
and U2158 (N_2158,In_531,In_743);
xnor U2159 (N_2159,In_459,In_1229);
nor U2160 (N_2160,In_132,In_1497);
nor U2161 (N_2161,In_25,In_330);
xor U2162 (N_2162,In_876,In_1144);
nand U2163 (N_2163,In_303,In_468);
xnor U2164 (N_2164,In_1011,In_697);
nand U2165 (N_2165,In_710,In_901);
nand U2166 (N_2166,In_1361,In_585);
and U2167 (N_2167,In_311,In_14);
nand U2168 (N_2168,In_267,In_364);
xor U2169 (N_2169,In_830,In_124);
nand U2170 (N_2170,In_296,In_1418);
nor U2171 (N_2171,In_53,In_1487);
nand U2172 (N_2172,In_1164,In_1331);
or U2173 (N_2173,In_751,In_733);
xnor U2174 (N_2174,In_1342,In_336);
nand U2175 (N_2175,In_977,In_1170);
or U2176 (N_2176,In_223,In_1207);
nor U2177 (N_2177,In_374,In_1295);
or U2178 (N_2178,In_959,In_1356);
xor U2179 (N_2179,In_939,In_1212);
or U2180 (N_2180,In_737,In_644);
or U2181 (N_2181,In_387,In_1123);
and U2182 (N_2182,In_257,In_146);
and U2183 (N_2183,In_1253,In_1221);
or U2184 (N_2184,In_337,In_404);
and U2185 (N_2185,In_888,In_636);
xnor U2186 (N_2186,In_1294,In_1322);
nor U2187 (N_2187,In_807,In_677);
or U2188 (N_2188,In_1130,In_118);
nand U2189 (N_2189,In_1401,In_1287);
nor U2190 (N_2190,In_415,In_490);
nor U2191 (N_2191,In_150,In_1048);
nor U2192 (N_2192,In_833,In_693);
xor U2193 (N_2193,In_686,In_23);
nand U2194 (N_2194,In_1257,In_711);
or U2195 (N_2195,In_1054,In_1180);
nor U2196 (N_2196,In_603,In_659);
or U2197 (N_2197,In_971,In_186);
nor U2198 (N_2198,In_674,In_1282);
nor U2199 (N_2199,In_916,In_1496);
nor U2200 (N_2200,In_414,In_1363);
and U2201 (N_2201,In_1450,In_1447);
nor U2202 (N_2202,In_615,In_291);
nand U2203 (N_2203,In_912,In_1067);
and U2204 (N_2204,In_1080,In_1180);
nor U2205 (N_2205,In_1420,In_613);
or U2206 (N_2206,In_1362,In_1160);
nand U2207 (N_2207,In_1055,In_517);
and U2208 (N_2208,In_1092,In_943);
and U2209 (N_2209,In_1036,In_1065);
nand U2210 (N_2210,In_153,In_149);
xnor U2211 (N_2211,In_1049,In_1282);
xor U2212 (N_2212,In_538,In_740);
nand U2213 (N_2213,In_1372,In_302);
nand U2214 (N_2214,In_1400,In_107);
nand U2215 (N_2215,In_1165,In_143);
or U2216 (N_2216,In_1455,In_933);
xnor U2217 (N_2217,In_414,In_599);
nor U2218 (N_2218,In_454,In_1279);
and U2219 (N_2219,In_241,In_1100);
xor U2220 (N_2220,In_62,In_1013);
nor U2221 (N_2221,In_839,In_333);
and U2222 (N_2222,In_34,In_235);
nor U2223 (N_2223,In_311,In_572);
or U2224 (N_2224,In_583,In_265);
and U2225 (N_2225,In_880,In_589);
and U2226 (N_2226,In_559,In_360);
nand U2227 (N_2227,In_1231,In_1309);
nor U2228 (N_2228,In_1215,In_130);
and U2229 (N_2229,In_1137,In_810);
and U2230 (N_2230,In_1166,In_8);
nand U2231 (N_2231,In_1182,In_379);
nand U2232 (N_2232,In_1407,In_759);
and U2233 (N_2233,In_544,In_349);
or U2234 (N_2234,In_1314,In_79);
nand U2235 (N_2235,In_1436,In_72);
nor U2236 (N_2236,In_593,In_1083);
xor U2237 (N_2237,In_1008,In_72);
and U2238 (N_2238,In_1330,In_1111);
and U2239 (N_2239,In_171,In_1186);
or U2240 (N_2240,In_1476,In_567);
xnor U2241 (N_2241,In_550,In_372);
xnor U2242 (N_2242,In_894,In_906);
nor U2243 (N_2243,In_1429,In_898);
and U2244 (N_2244,In_105,In_615);
xor U2245 (N_2245,In_447,In_1306);
nand U2246 (N_2246,In_1341,In_330);
nand U2247 (N_2247,In_1089,In_969);
and U2248 (N_2248,In_987,In_167);
xnor U2249 (N_2249,In_757,In_1419);
xor U2250 (N_2250,In_965,In_1055);
xor U2251 (N_2251,In_1101,In_852);
nand U2252 (N_2252,In_1220,In_673);
nand U2253 (N_2253,In_1424,In_763);
or U2254 (N_2254,In_1479,In_69);
nand U2255 (N_2255,In_1004,In_192);
nor U2256 (N_2256,In_341,In_510);
and U2257 (N_2257,In_318,In_939);
or U2258 (N_2258,In_417,In_844);
nor U2259 (N_2259,In_1411,In_751);
or U2260 (N_2260,In_1344,In_103);
and U2261 (N_2261,In_419,In_1384);
or U2262 (N_2262,In_131,In_739);
xnor U2263 (N_2263,In_164,In_174);
or U2264 (N_2264,In_1157,In_63);
nor U2265 (N_2265,In_1178,In_493);
nand U2266 (N_2266,In_1498,In_1249);
and U2267 (N_2267,In_860,In_636);
nor U2268 (N_2268,In_1256,In_55);
nor U2269 (N_2269,In_1451,In_10);
xor U2270 (N_2270,In_951,In_1408);
or U2271 (N_2271,In_500,In_31);
nor U2272 (N_2272,In_117,In_153);
and U2273 (N_2273,In_1156,In_1377);
nor U2274 (N_2274,In_959,In_676);
nand U2275 (N_2275,In_384,In_1093);
or U2276 (N_2276,In_846,In_304);
nor U2277 (N_2277,In_270,In_419);
nor U2278 (N_2278,In_990,In_868);
or U2279 (N_2279,In_213,In_49);
and U2280 (N_2280,In_1037,In_890);
or U2281 (N_2281,In_1437,In_440);
or U2282 (N_2282,In_772,In_266);
nand U2283 (N_2283,In_1013,In_1441);
xor U2284 (N_2284,In_1374,In_1455);
nor U2285 (N_2285,In_1387,In_867);
xnor U2286 (N_2286,In_466,In_1103);
xnor U2287 (N_2287,In_1496,In_958);
xor U2288 (N_2288,In_883,In_704);
or U2289 (N_2289,In_1304,In_893);
xor U2290 (N_2290,In_101,In_1183);
nand U2291 (N_2291,In_690,In_266);
nor U2292 (N_2292,In_809,In_1425);
and U2293 (N_2293,In_1423,In_1408);
and U2294 (N_2294,In_998,In_676);
xnor U2295 (N_2295,In_207,In_276);
or U2296 (N_2296,In_1248,In_144);
and U2297 (N_2297,In_956,In_1336);
nor U2298 (N_2298,In_664,In_25);
xnor U2299 (N_2299,In_80,In_1435);
nor U2300 (N_2300,In_106,In_870);
nand U2301 (N_2301,In_1077,In_1424);
and U2302 (N_2302,In_591,In_1149);
or U2303 (N_2303,In_901,In_1022);
xnor U2304 (N_2304,In_786,In_866);
nand U2305 (N_2305,In_636,In_844);
xnor U2306 (N_2306,In_1133,In_528);
and U2307 (N_2307,In_89,In_674);
or U2308 (N_2308,In_627,In_1168);
or U2309 (N_2309,In_970,In_812);
and U2310 (N_2310,In_503,In_1086);
xor U2311 (N_2311,In_1093,In_1064);
and U2312 (N_2312,In_1312,In_1313);
nand U2313 (N_2313,In_389,In_426);
nor U2314 (N_2314,In_244,In_988);
xnor U2315 (N_2315,In_980,In_431);
xnor U2316 (N_2316,In_680,In_378);
and U2317 (N_2317,In_963,In_946);
nand U2318 (N_2318,In_467,In_1007);
nand U2319 (N_2319,In_1381,In_1468);
or U2320 (N_2320,In_835,In_1000);
nand U2321 (N_2321,In_1416,In_401);
and U2322 (N_2322,In_1126,In_147);
nor U2323 (N_2323,In_896,In_1309);
nand U2324 (N_2324,In_446,In_560);
and U2325 (N_2325,In_1139,In_167);
nand U2326 (N_2326,In_29,In_72);
or U2327 (N_2327,In_335,In_110);
nor U2328 (N_2328,In_123,In_785);
xor U2329 (N_2329,In_1041,In_1147);
xor U2330 (N_2330,In_1399,In_1372);
nand U2331 (N_2331,In_497,In_826);
nor U2332 (N_2332,In_483,In_1126);
xor U2333 (N_2333,In_362,In_791);
nand U2334 (N_2334,In_772,In_305);
or U2335 (N_2335,In_1246,In_680);
and U2336 (N_2336,In_1130,In_710);
xnor U2337 (N_2337,In_386,In_72);
nor U2338 (N_2338,In_244,In_424);
or U2339 (N_2339,In_1452,In_1403);
nor U2340 (N_2340,In_1254,In_1237);
or U2341 (N_2341,In_1168,In_665);
nand U2342 (N_2342,In_908,In_30);
nor U2343 (N_2343,In_231,In_1067);
and U2344 (N_2344,In_772,In_320);
and U2345 (N_2345,In_402,In_712);
and U2346 (N_2346,In_359,In_291);
and U2347 (N_2347,In_1365,In_1304);
nor U2348 (N_2348,In_235,In_1471);
xor U2349 (N_2349,In_1184,In_1193);
xnor U2350 (N_2350,In_1239,In_1379);
nor U2351 (N_2351,In_951,In_97);
and U2352 (N_2352,In_1040,In_370);
xor U2353 (N_2353,In_1214,In_670);
and U2354 (N_2354,In_878,In_494);
xnor U2355 (N_2355,In_574,In_572);
nand U2356 (N_2356,In_592,In_809);
nand U2357 (N_2357,In_927,In_1421);
nor U2358 (N_2358,In_18,In_922);
or U2359 (N_2359,In_286,In_1039);
xnor U2360 (N_2360,In_120,In_1344);
nand U2361 (N_2361,In_1162,In_398);
nand U2362 (N_2362,In_488,In_188);
nor U2363 (N_2363,In_955,In_238);
nand U2364 (N_2364,In_1496,In_169);
nand U2365 (N_2365,In_302,In_1399);
nor U2366 (N_2366,In_311,In_67);
or U2367 (N_2367,In_685,In_791);
xnor U2368 (N_2368,In_1464,In_234);
xor U2369 (N_2369,In_453,In_1382);
nor U2370 (N_2370,In_695,In_1115);
xor U2371 (N_2371,In_163,In_1168);
or U2372 (N_2372,In_118,In_339);
nand U2373 (N_2373,In_153,In_407);
nor U2374 (N_2374,In_747,In_468);
nand U2375 (N_2375,In_353,In_233);
or U2376 (N_2376,In_524,In_1170);
nor U2377 (N_2377,In_568,In_422);
xor U2378 (N_2378,In_431,In_54);
or U2379 (N_2379,In_932,In_696);
and U2380 (N_2380,In_324,In_140);
or U2381 (N_2381,In_603,In_485);
and U2382 (N_2382,In_8,In_827);
nor U2383 (N_2383,In_613,In_1126);
and U2384 (N_2384,In_638,In_1132);
or U2385 (N_2385,In_1106,In_1273);
xor U2386 (N_2386,In_680,In_694);
or U2387 (N_2387,In_426,In_1014);
xor U2388 (N_2388,In_1034,In_848);
nor U2389 (N_2389,In_1445,In_916);
xor U2390 (N_2390,In_19,In_781);
and U2391 (N_2391,In_574,In_698);
or U2392 (N_2392,In_791,In_754);
nand U2393 (N_2393,In_401,In_780);
or U2394 (N_2394,In_398,In_1015);
nor U2395 (N_2395,In_1479,In_1358);
and U2396 (N_2396,In_1318,In_128);
xnor U2397 (N_2397,In_738,In_1251);
xor U2398 (N_2398,In_42,In_450);
and U2399 (N_2399,In_1025,In_419);
xor U2400 (N_2400,In_1023,In_677);
xor U2401 (N_2401,In_227,In_239);
xor U2402 (N_2402,In_592,In_898);
nand U2403 (N_2403,In_169,In_651);
and U2404 (N_2404,In_89,In_711);
and U2405 (N_2405,In_189,In_906);
and U2406 (N_2406,In_1153,In_815);
nor U2407 (N_2407,In_967,In_980);
nand U2408 (N_2408,In_1459,In_296);
nand U2409 (N_2409,In_1056,In_644);
xnor U2410 (N_2410,In_223,In_110);
xor U2411 (N_2411,In_166,In_444);
or U2412 (N_2412,In_324,In_1078);
nand U2413 (N_2413,In_1148,In_112);
or U2414 (N_2414,In_1326,In_76);
nor U2415 (N_2415,In_1408,In_284);
and U2416 (N_2416,In_874,In_1416);
and U2417 (N_2417,In_1212,In_202);
nand U2418 (N_2418,In_1228,In_353);
and U2419 (N_2419,In_1016,In_414);
xnor U2420 (N_2420,In_37,In_67);
and U2421 (N_2421,In_1437,In_1187);
nor U2422 (N_2422,In_268,In_1354);
nor U2423 (N_2423,In_13,In_331);
and U2424 (N_2424,In_656,In_1431);
nor U2425 (N_2425,In_878,In_261);
xor U2426 (N_2426,In_392,In_876);
or U2427 (N_2427,In_729,In_846);
nand U2428 (N_2428,In_3,In_795);
nor U2429 (N_2429,In_412,In_584);
xnor U2430 (N_2430,In_1213,In_1180);
xnor U2431 (N_2431,In_310,In_470);
nand U2432 (N_2432,In_1079,In_867);
nor U2433 (N_2433,In_1248,In_125);
nand U2434 (N_2434,In_1320,In_586);
or U2435 (N_2435,In_823,In_939);
and U2436 (N_2436,In_147,In_1274);
or U2437 (N_2437,In_344,In_790);
or U2438 (N_2438,In_457,In_207);
and U2439 (N_2439,In_1230,In_153);
nor U2440 (N_2440,In_1068,In_184);
and U2441 (N_2441,In_637,In_855);
and U2442 (N_2442,In_1035,In_82);
nand U2443 (N_2443,In_887,In_226);
xnor U2444 (N_2444,In_356,In_1042);
xor U2445 (N_2445,In_977,In_1138);
and U2446 (N_2446,In_1069,In_790);
xor U2447 (N_2447,In_375,In_339);
xnor U2448 (N_2448,In_762,In_730);
nand U2449 (N_2449,In_1183,In_469);
or U2450 (N_2450,In_1071,In_57);
or U2451 (N_2451,In_126,In_1283);
xnor U2452 (N_2452,In_632,In_62);
nand U2453 (N_2453,In_700,In_810);
xnor U2454 (N_2454,In_38,In_534);
and U2455 (N_2455,In_927,In_1325);
and U2456 (N_2456,In_1022,In_1156);
and U2457 (N_2457,In_865,In_1188);
xnor U2458 (N_2458,In_956,In_391);
nor U2459 (N_2459,In_1276,In_1369);
xnor U2460 (N_2460,In_623,In_863);
nor U2461 (N_2461,In_727,In_166);
nand U2462 (N_2462,In_837,In_562);
nor U2463 (N_2463,In_351,In_1171);
and U2464 (N_2464,In_1185,In_16);
nand U2465 (N_2465,In_275,In_278);
xnor U2466 (N_2466,In_1002,In_1292);
nor U2467 (N_2467,In_597,In_252);
nor U2468 (N_2468,In_398,In_1462);
nand U2469 (N_2469,In_607,In_15);
and U2470 (N_2470,In_654,In_1228);
and U2471 (N_2471,In_1444,In_490);
xnor U2472 (N_2472,In_172,In_437);
xnor U2473 (N_2473,In_598,In_690);
or U2474 (N_2474,In_892,In_577);
xnor U2475 (N_2475,In_1145,In_729);
nand U2476 (N_2476,In_1486,In_243);
nor U2477 (N_2477,In_375,In_854);
nor U2478 (N_2478,In_151,In_1218);
nor U2479 (N_2479,In_1328,In_1331);
nor U2480 (N_2480,In_61,In_1412);
or U2481 (N_2481,In_1419,In_1212);
nor U2482 (N_2482,In_1306,In_526);
and U2483 (N_2483,In_1091,In_1317);
or U2484 (N_2484,In_314,In_1465);
xor U2485 (N_2485,In_1372,In_857);
or U2486 (N_2486,In_915,In_942);
xnor U2487 (N_2487,In_891,In_440);
and U2488 (N_2488,In_1393,In_653);
nand U2489 (N_2489,In_609,In_567);
xnor U2490 (N_2490,In_1451,In_1222);
xnor U2491 (N_2491,In_1359,In_1163);
nand U2492 (N_2492,In_1375,In_817);
xor U2493 (N_2493,In_29,In_20);
and U2494 (N_2494,In_1088,In_386);
nor U2495 (N_2495,In_1189,In_1125);
nand U2496 (N_2496,In_292,In_968);
nand U2497 (N_2497,In_97,In_962);
or U2498 (N_2498,In_755,In_485);
nand U2499 (N_2499,In_314,In_955);
xnor U2500 (N_2500,In_211,In_702);
and U2501 (N_2501,In_1117,In_197);
and U2502 (N_2502,In_1392,In_773);
nor U2503 (N_2503,In_119,In_284);
nor U2504 (N_2504,In_166,In_1274);
and U2505 (N_2505,In_1404,In_997);
nor U2506 (N_2506,In_912,In_883);
and U2507 (N_2507,In_1388,In_179);
nor U2508 (N_2508,In_1451,In_1204);
nand U2509 (N_2509,In_1259,In_118);
and U2510 (N_2510,In_1181,In_661);
or U2511 (N_2511,In_466,In_1341);
xor U2512 (N_2512,In_778,In_1383);
and U2513 (N_2513,In_367,In_41);
or U2514 (N_2514,In_1310,In_1070);
nand U2515 (N_2515,In_1354,In_1313);
xor U2516 (N_2516,In_534,In_720);
and U2517 (N_2517,In_1311,In_482);
nand U2518 (N_2518,In_103,In_6);
or U2519 (N_2519,In_325,In_301);
nor U2520 (N_2520,In_947,In_109);
nor U2521 (N_2521,In_488,In_570);
nand U2522 (N_2522,In_534,In_1388);
xor U2523 (N_2523,In_1081,In_1305);
and U2524 (N_2524,In_881,In_190);
or U2525 (N_2525,In_582,In_1210);
and U2526 (N_2526,In_255,In_908);
xnor U2527 (N_2527,In_248,In_802);
xnor U2528 (N_2528,In_101,In_207);
nor U2529 (N_2529,In_829,In_410);
or U2530 (N_2530,In_161,In_27);
or U2531 (N_2531,In_1197,In_794);
nor U2532 (N_2532,In_1128,In_194);
or U2533 (N_2533,In_1293,In_768);
xnor U2534 (N_2534,In_434,In_457);
xor U2535 (N_2535,In_1406,In_543);
xnor U2536 (N_2536,In_520,In_1295);
nand U2537 (N_2537,In_1324,In_508);
and U2538 (N_2538,In_504,In_486);
or U2539 (N_2539,In_1063,In_111);
or U2540 (N_2540,In_975,In_373);
nand U2541 (N_2541,In_736,In_472);
and U2542 (N_2542,In_1325,In_1141);
xnor U2543 (N_2543,In_988,In_25);
and U2544 (N_2544,In_961,In_225);
nand U2545 (N_2545,In_1151,In_1427);
nor U2546 (N_2546,In_1307,In_1379);
and U2547 (N_2547,In_477,In_1227);
and U2548 (N_2548,In_709,In_352);
or U2549 (N_2549,In_369,In_505);
xor U2550 (N_2550,In_22,In_935);
or U2551 (N_2551,In_1415,In_343);
or U2552 (N_2552,In_806,In_397);
nor U2553 (N_2553,In_1409,In_231);
xnor U2554 (N_2554,In_326,In_285);
and U2555 (N_2555,In_825,In_1268);
nand U2556 (N_2556,In_1428,In_752);
or U2557 (N_2557,In_746,In_741);
or U2558 (N_2558,In_973,In_298);
or U2559 (N_2559,In_1042,In_1321);
or U2560 (N_2560,In_37,In_1095);
nor U2561 (N_2561,In_1454,In_919);
and U2562 (N_2562,In_1150,In_0);
nand U2563 (N_2563,In_485,In_1222);
or U2564 (N_2564,In_1291,In_155);
nor U2565 (N_2565,In_1128,In_54);
nor U2566 (N_2566,In_521,In_426);
and U2567 (N_2567,In_1233,In_1163);
nor U2568 (N_2568,In_749,In_958);
and U2569 (N_2569,In_910,In_623);
or U2570 (N_2570,In_79,In_562);
xnor U2571 (N_2571,In_653,In_950);
nor U2572 (N_2572,In_328,In_770);
and U2573 (N_2573,In_655,In_447);
and U2574 (N_2574,In_610,In_237);
nand U2575 (N_2575,In_1144,In_62);
xnor U2576 (N_2576,In_656,In_719);
or U2577 (N_2577,In_1496,In_1004);
xnor U2578 (N_2578,In_932,In_1128);
nand U2579 (N_2579,In_746,In_1351);
and U2580 (N_2580,In_720,In_1471);
xnor U2581 (N_2581,In_209,In_901);
nor U2582 (N_2582,In_390,In_681);
xnor U2583 (N_2583,In_327,In_107);
nand U2584 (N_2584,In_667,In_303);
nor U2585 (N_2585,In_848,In_302);
or U2586 (N_2586,In_1488,In_801);
nand U2587 (N_2587,In_370,In_611);
or U2588 (N_2588,In_676,In_552);
nand U2589 (N_2589,In_73,In_421);
or U2590 (N_2590,In_518,In_620);
nor U2591 (N_2591,In_1407,In_827);
xnor U2592 (N_2592,In_950,In_53);
nand U2593 (N_2593,In_210,In_872);
nor U2594 (N_2594,In_801,In_732);
nand U2595 (N_2595,In_857,In_151);
xnor U2596 (N_2596,In_1087,In_497);
or U2597 (N_2597,In_176,In_753);
or U2598 (N_2598,In_1495,In_446);
nand U2599 (N_2599,In_1036,In_574);
or U2600 (N_2600,In_950,In_1044);
nor U2601 (N_2601,In_338,In_886);
and U2602 (N_2602,In_394,In_627);
nand U2603 (N_2603,In_1335,In_218);
xnor U2604 (N_2604,In_927,In_847);
or U2605 (N_2605,In_605,In_377);
and U2606 (N_2606,In_23,In_276);
nand U2607 (N_2607,In_671,In_182);
and U2608 (N_2608,In_966,In_523);
and U2609 (N_2609,In_395,In_1260);
xor U2610 (N_2610,In_87,In_294);
and U2611 (N_2611,In_23,In_1478);
and U2612 (N_2612,In_1267,In_1036);
nand U2613 (N_2613,In_646,In_1001);
nor U2614 (N_2614,In_1403,In_462);
xnor U2615 (N_2615,In_839,In_1258);
nand U2616 (N_2616,In_781,In_469);
nand U2617 (N_2617,In_1293,In_561);
or U2618 (N_2618,In_599,In_786);
xor U2619 (N_2619,In_99,In_744);
and U2620 (N_2620,In_1249,In_747);
or U2621 (N_2621,In_1058,In_200);
or U2622 (N_2622,In_1186,In_1052);
nor U2623 (N_2623,In_1113,In_398);
xnor U2624 (N_2624,In_986,In_1084);
or U2625 (N_2625,In_787,In_425);
xnor U2626 (N_2626,In_327,In_859);
nand U2627 (N_2627,In_284,In_421);
xnor U2628 (N_2628,In_241,In_97);
nand U2629 (N_2629,In_1169,In_925);
nand U2630 (N_2630,In_170,In_249);
nand U2631 (N_2631,In_250,In_163);
nand U2632 (N_2632,In_999,In_673);
nor U2633 (N_2633,In_533,In_1321);
nand U2634 (N_2634,In_589,In_1092);
nand U2635 (N_2635,In_936,In_895);
or U2636 (N_2636,In_359,In_906);
and U2637 (N_2637,In_632,In_1170);
or U2638 (N_2638,In_7,In_563);
nor U2639 (N_2639,In_1056,In_822);
and U2640 (N_2640,In_1370,In_1228);
or U2641 (N_2641,In_346,In_1053);
nor U2642 (N_2642,In_739,In_1108);
and U2643 (N_2643,In_1314,In_761);
nor U2644 (N_2644,In_1470,In_0);
nand U2645 (N_2645,In_277,In_858);
or U2646 (N_2646,In_1450,In_65);
nand U2647 (N_2647,In_913,In_1144);
and U2648 (N_2648,In_1350,In_356);
nor U2649 (N_2649,In_1001,In_1253);
nor U2650 (N_2650,In_526,In_355);
nand U2651 (N_2651,In_1379,In_1390);
xnor U2652 (N_2652,In_1339,In_1487);
xor U2653 (N_2653,In_1080,In_609);
nor U2654 (N_2654,In_891,In_1055);
xor U2655 (N_2655,In_35,In_630);
and U2656 (N_2656,In_1107,In_1212);
nand U2657 (N_2657,In_994,In_360);
or U2658 (N_2658,In_600,In_420);
nor U2659 (N_2659,In_467,In_619);
and U2660 (N_2660,In_1146,In_1163);
or U2661 (N_2661,In_1190,In_1419);
or U2662 (N_2662,In_876,In_501);
xor U2663 (N_2663,In_691,In_68);
nor U2664 (N_2664,In_1436,In_390);
nand U2665 (N_2665,In_131,In_77);
nand U2666 (N_2666,In_28,In_700);
nor U2667 (N_2667,In_790,In_438);
xor U2668 (N_2668,In_158,In_1080);
or U2669 (N_2669,In_532,In_1350);
nor U2670 (N_2670,In_286,In_824);
nand U2671 (N_2671,In_1016,In_416);
xnor U2672 (N_2672,In_258,In_242);
or U2673 (N_2673,In_1078,In_1026);
xnor U2674 (N_2674,In_1280,In_883);
nand U2675 (N_2675,In_1008,In_1005);
nand U2676 (N_2676,In_1190,In_349);
or U2677 (N_2677,In_968,In_670);
nand U2678 (N_2678,In_410,In_290);
nand U2679 (N_2679,In_79,In_716);
and U2680 (N_2680,In_1233,In_207);
or U2681 (N_2681,In_356,In_802);
and U2682 (N_2682,In_410,In_601);
nor U2683 (N_2683,In_1089,In_866);
nor U2684 (N_2684,In_1141,In_803);
and U2685 (N_2685,In_783,In_185);
nor U2686 (N_2686,In_1220,In_34);
nor U2687 (N_2687,In_36,In_709);
or U2688 (N_2688,In_370,In_542);
xor U2689 (N_2689,In_252,In_147);
and U2690 (N_2690,In_1449,In_882);
or U2691 (N_2691,In_1247,In_1175);
or U2692 (N_2692,In_539,In_1092);
xnor U2693 (N_2693,In_489,In_1203);
and U2694 (N_2694,In_186,In_84);
and U2695 (N_2695,In_754,In_605);
xnor U2696 (N_2696,In_807,In_436);
and U2697 (N_2697,In_324,In_119);
and U2698 (N_2698,In_674,In_1021);
nor U2699 (N_2699,In_694,In_1318);
and U2700 (N_2700,In_676,In_32);
nor U2701 (N_2701,In_761,In_661);
nor U2702 (N_2702,In_460,In_713);
nand U2703 (N_2703,In_687,In_1169);
xor U2704 (N_2704,In_1258,In_421);
nor U2705 (N_2705,In_1229,In_1290);
nand U2706 (N_2706,In_1410,In_1477);
nor U2707 (N_2707,In_480,In_519);
and U2708 (N_2708,In_123,In_319);
nand U2709 (N_2709,In_908,In_536);
or U2710 (N_2710,In_658,In_251);
or U2711 (N_2711,In_1265,In_1405);
and U2712 (N_2712,In_769,In_1167);
xnor U2713 (N_2713,In_308,In_1258);
and U2714 (N_2714,In_799,In_334);
nor U2715 (N_2715,In_1208,In_276);
or U2716 (N_2716,In_724,In_7);
xor U2717 (N_2717,In_67,In_1207);
xnor U2718 (N_2718,In_1316,In_843);
nand U2719 (N_2719,In_340,In_809);
nand U2720 (N_2720,In_1280,In_1484);
nand U2721 (N_2721,In_781,In_845);
xor U2722 (N_2722,In_942,In_141);
nor U2723 (N_2723,In_519,In_412);
and U2724 (N_2724,In_378,In_778);
and U2725 (N_2725,In_413,In_711);
nand U2726 (N_2726,In_46,In_1107);
and U2727 (N_2727,In_12,In_770);
and U2728 (N_2728,In_1227,In_1258);
and U2729 (N_2729,In_650,In_677);
or U2730 (N_2730,In_143,In_650);
and U2731 (N_2731,In_1244,In_608);
nor U2732 (N_2732,In_1275,In_397);
or U2733 (N_2733,In_908,In_387);
nor U2734 (N_2734,In_698,In_897);
nor U2735 (N_2735,In_572,In_926);
xor U2736 (N_2736,In_446,In_710);
nor U2737 (N_2737,In_933,In_1156);
and U2738 (N_2738,In_701,In_655);
or U2739 (N_2739,In_1316,In_1326);
xor U2740 (N_2740,In_1045,In_751);
nor U2741 (N_2741,In_936,In_1258);
nand U2742 (N_2742,In_383,In_418);
or U2743 (N_2743,In_732,In_598);
nand U2744 (N_2744,In_61,In_1394);
and U2745 (N_2745,In_1457,In_960);
xor U2746 (N_2746,In_1064,In_937);
and U2747 (N_2747,In_963,In_214);
nor U2748 (N_2748,In_1470,In_847);
xor U2749 (N_2749,In_890,In_75);
xor U2750 (N_2750,In_1182,In_936);
and U2751 (N_2751,In_591,In_1474);
xnor U2752 (N_2752,In_1252,In_1262);
and U2753 (N_2753,In_321,In_847);
and U2754 (N_2754,In_585,In_842);
nor U2755 (N_2755,In_156,In_1376);
and U2756 (N_2756,In_268,In_147);
xnor U2757 (N_2757,In_486,In_1109);
and U2758 (N_2758,In_1100,In_299);
and U2759 (N_2759,In_1188,In_619);
xor U2760 (N_2760,In_471,In_394);
xor U2761 (N_2761,In_500,In_915);
or U2762 (N_2762,In_344,In_432);
xnor U2763 (N_2763,In_1055,In_1492);
or U2764 (N_2764,In_958,In_280);
or U2765 (N_2765,In_1228,In_1218);
xor U2766 (N_2766,In_1093,In_970);
and U2767 (N_2767,In_948,In_826);
and U2768 (N_2768,In_1192,In_73);
and U2769 (N_2769,In_1250,In_730);
and U2770 (N_2770,In_533,In_1419);
nand U2771 (N_2771,In_270,In_636);
xnor U2772 (N_2772,In_944,In_618);
and U2773 (N_2773,In_326,In_771);
nand U2774 (N_2774,In_432,In_1285);
and U2775 (N_2775,In_293,In_982);
or U2776 (N_2776,In_331,In_852);
nor U2777 (N_2777,In_667,In_1174);
xor U2778 (N_2778,In_1184,In_252);
or U2779 (N_2779,In_13,In_1278);
xnor U2780 (N_2780,In_371,In_610);
or U2781 (N_2781,In_586,In_1131);
nand U2782 (N_2782,In_1315,In_539);
or U2783 (N_2783,In_1109,In_805);
and U2784 (N_2784,In_90,In_993);
or U2785 (N_2785,In_786,In_1010);
and U2786 (N_2786,In_683,In_10);
or U2787 (N_2787,In_419,In_913);
xnor U2788 (N_2788,In_1013,In_299);
or U2789 (N_2789,In_340,In_1496);
xor U2790 (N_2790,In_1085,In_927);
nor U2791 (N_2791,In_1287,In_1048);
and U2792 (N_2792,In_196,In_347);
nand U2793 (N_2793,In_1313,In_56);
or U2794 (N_2794,In_1434,In_980);
nand U2795 (N_2795,In_1289,In_1310);
xnor U2796 (N_2796,In_771,In_1056);
nand U2797 (N_2797,In_389,In_516);
nor U2798 (N_2798,In_332,In_1038);
xor U2799 (N_2799,In_622,In_320);
xnor U2800 (N_2800,In_702,In_289);
xnor U2801 (N_2801,In_1271,In_881);
nor U2802 (N_2802,In_1127,In_383);
or U2803 (N_2803,In_1147,In_607);
nor U2804 (N_2804,In_1088,In_1410);
xor U2805 (N_2805,In_378,In_1289);
nand U2806 (N_2806,In_884,In_977);
and U2807 (N_2807,In_276,In_434);
xor U2808 (N_2808,In_1457,In_1388);
nand U2809 (N_2809,In_253,In_1452);
nand U2810 (N_2810,In_943,In_483);
nor U2811 (N_2811,In_392,In_994);
or U2812 (N_2812,In_1078,In_457);
nor U2813 (N_2813,In_383,In_751);
nand U2814 (N_2814,In_210,In_1339);
or U2815 (N_2815,In_1408,In_863);
or U2816 (N_2816,In_1220,In_560);
or U2817 (N_2817,In_52,In_1114);
and U2818 (N_2818,In_703,In_1371);
nand U2819 (N_2819,In_1455,In_1021);
and U2820 (N_2820,In_261,In_1242);
nand U2821 (N_2821,In_239,In_78);
xnor U2822 (N_2822,In_312,In_1453);
or U2823 (N_2823,In_844,In_168);
nand U2824 (N_2824,In_947,In_585);
and U2825 (N_2825,In_544,In_386);
or U2826 (N_2826,In_757,In_1381);
nand U2827 (N_2827,In_995,In_918);
nor U2828 (N_2828,In_880,In_101);
and U2829 (N_2829,In_1343,In_1404);
nor U2830 (N_2830,In_459,In_1053);
and U2831 (N_2831,In_1446,In_594);
nand U2832 (N_2832,In_1223,In_415);
or U2833 (N_2833,In_72,In_177);
nand U2834 (N_2834,In_1279,In_581);
nand U2835 (N_2835,In_1417,In_502);
and U2836 (N_2836,In_213,In_542);
and U2837 (N_2837,In_624,In_373);
or U2838 (N_2838,In_1315,In_680);
nand U2839 (N_2839,In_481,In_839);
xor U2840 (N_2840,In_1223,In_352);
and U2841 (N_2841,In_1481,In_3);
or U2842 (N_2842,In_1,In_1091);
nor U2843 (N_2843,In_52,In_1004);
nand U2844 (N_2844,In_1428,In_596);
and U2845 (N_2845,In_599,In_122);
nor U2846 (N_2846,In_204,In_89);
nand U2847 (N_2847,In_1337,In_936);
nand U2848 (N_2848,In_1248,In_863);
or U2849 (N_2849,In_932,In_101);
nand U2850 (N_2850,In_151,In_435);
nand U2851 (N_2851,In_869,In_1433);
xor U2852 (N_2852,In_825,In_918);
xnor U2853 (N_2853,In_1072,In_510);
and U2854 (N_2854,In_253,In_1092);
nand U2855 (N_2855,In_404,In_1341);
or U2856 (N_2856,In_213,In_459);
xor U2857 (N_2857,In_1167,In_1296);
xor U2858 (N_2858,In_1369,In_1097);
nor U2859 (N_2859,In_841,In_130);
nor U2860 (N_2860,In_919,In_561);
nor U2861 (N_2861,In_59,In_521);
or U2862 (N_2862,In_205,In_924);
or U2863 (N_2863,In_596,In_929);
or U2864 (N_2864,In_1213,In_168);
xor U2865 (N_2865,In_432,In_196);
or U2866 (N_2866,In_1092,In_1442);
nand U2867 (N_2867,In_513,In_384);
nor U2868 (N_2868,In_275,In_1454);
and U2869 (N_2869,In_50,In_188);
or U2870 (N_2870,In_45,In_638);
nor U2871 (N_2871,In_1447,In_633);
nand U2872 (N_2872,In_116,In_1151);
nor U2873 (N_2873,In_482,In_330);
nand U2874 (N_2874,In_841,In_1165);
and U2875 (N_2875,In_1274,In_1057);
or U2876 (N_2876,In_1275,In_1280);
nand U2877 (N_2877,In_1239,In_334);
and U2878 (N_2878,In_165,In_479);
and U2879 (N_2879,In_291,In_1458);
xor U2880 (N_2880,In_489,In_966);
nand U2881 (N_2881,In_262,In_1387);
and U2882 (N_2882,In_262,In_1446);
or U2883 (N_2883,In_24,In_1226);
and U2884 (N_2884,In_622,In_388);
and U2885 (N_2885,In_563,In_515);
xnor U2886 (N_2886,In_1421,In_528);
nor U2887 (N_2887,In_1433,In_479);
xnor U2888 (N_2888,In_130,In_42);
nor U2889 (N_2889,In_553,In_843);
or U2890 (N_2890,In_1384,In_616);
xnor U2891 (N_2891,In_65,In_1145);
xnor U2892 (N_2892,In_1207,In_182);
and U2893 (N_2893,In_525,In_248);
nor U2894 (N_2894,In_209,In_889);
or U2895 (N_2895,In_292,In_263);
and U2896 (N_2896,In_879,In_1021);
nor U2897 (N_2897,In_87,In_1078);
nor U2898 (N_2898,In_703,In_1111);
xor U2899 (N_2899,In_971,In_405);
nor U2900 (N_2900,In_1112,In_315);
or U2901 (N_2901,In_571,In_979);
nor U2902 (N_2902,In_1419,In_1182);
nor U2903 (N_2903,In_774,In_1439);
or U2904 (N_2904,In_1129,In_869);
and U2905 (N_2905,In_567,In_761);
nand U2906 (N_2906,In_912,In_1459);
and U2907 (N_2907,In_913,In_1498);
xnor U2908 (N_2908,In_757,In_177);
nor U2909 (N_2909,In_863,In_117);
or U2910 (N_2910,In_934,In_809);
and U2911 (N_2911,In_844,In_552);
nor U2912 (N_2912,In_193,In_421);
xnor U2913 (N_2913,In_898,In_1366);
or U2914 (N_2914,In_1259,In_706);
nor U2915 (N_2915,In_1136,In_628);
nor U2916 (N_2916,In_1135,In_1484);
or U2917 (N_2917,In_1147,In_535);
nor U2918 (N_2918,In_1174,In_387);
or U2919 (N_2919,In_516,In_468);
nor U2920 (N_2920,In_866,In_966);
nor U2921 (N_2921,In_637,In_1086);
or U2922 (N_2922,In_792,In_941);
and U2923 (N_2923,In_1458,In_368);
xnor U2924 (N_2924,In_1315,In_34);
xnor U2925 (N_2925,In_299,In_542);
xnor U2926 (N_2926,In_748,In_545);
nand U2927 (N_2927,In_621,In_161);
nor U2928 (N_2928,In_531,In_527);
or U2929 (N_2929,In_720,In_767);
or U2930 (N_2930,In_961,In_1350);
and U2931 (N_2931,In_1376,In_133);
xor U2932 (N_2932,In_934,In_4);
or U2933 (N_2933,In_706,In_1438);
or U2934 (N_2934,In_679,In_1343);
or U2935 (N_2935,In_775,In_1431);
and U2936 (N_2936,In_991,In_643);
and U2937 (N_2937,In_1473,In_1059);
xnor U2938 (N_2938,In_583,In_826);
nand U2939 (N_2939,In_936,In_695);
xor U2940 (N_2940,In_310,In_514);
nand U2941 (N_2941,In_525,In_939);
nor U2942 (N_2942,In_853,In_22);
xor U2943 (N_2943,In_285,In_691);
xnor U2944 (N_2944,In_686,In_918);
or U2945 (N_2945,In_169,In_988);
nor U2946 (N_2946,In_491,In_35);
xnor U2947 (N_2947,In_63,In_35);
xor U2948 (N_2948,In_328,In_799);
xnor U2949 (N_2949,In_899,In_960);
nand U2950 (N_2950,In_128,In_190);
or U2951 (N_2951,In_1238,In_1374);
and U2952 (N_2952,In_647,In_938);
and U2953 (N_2953,In_442,In_205);
xor U2954 (N_2954,In_94,In_464);
or U2955 (N_2955,In_233,In_1377);
nor U2956 (N_2956,In_1455,In_305);
and U2957 (N_2957,In_1317,In_1188);
xor U2958 (N_2958,In_567,In_1355);
nor U2959 (N_2959,In_583,In_1380);
nor U2960 (N_2960,In_709,In_1221);
nor U2961 (N_2961,In_1344,In_973);
nor U2962 (N_2962,In_754,In_521);
xor U2963 (N_2963,In_456,In_1248);
xnor U2964 (N_2964,In_764,In_794);
or U2965 (N_2965,In_906,In_1122);
nand U2966 (N_2966,In_387,In_391);
xnor U2967 (N_2967,In_1303,In_1227);
xor U2968 (N_2968,In_1164,In_1167);
nand U2969 (N_2969,In_621,In_1156);
or U2970 (N_2970,In_285,In_869);
nand U2971 (N_2971,In_514,In_501);
and U2972 (N_2972,In_248,In_152);
nand U2973 (N_2973,In_570,In_62);
xnor U2974 (N_2974,In_951,In_905);
or U2975 (N_2975,In_857,In_392);
xor U2976 (N_2976,In_527,In_1268);
or U2977 (N_2977,In_473,In_1423);
nand U2978 (N_2978,In_369,In_938);
xor U2979 (N_2979,In_1109,In_861);
nor U2980 (N_2980,In_181,In_174);
or U2981 (N_2981,In_824,In_513);
or U2982 (N_2982,In_604,In_751);
nand U2983 (N_2983,In_611,In_319);
nand U2984 (N_2984,In_886,In_832);
and U2985 (N_2985,In_3,In_26);
or U2986 (N_2986,In_128,In_1086);
nand U2987 (N_2987,In_940,In_614);
nor U2988 (N_2988,In_718,In_196);
or U2989 (N_2989,In_459,In_1304);
or U2990 (N_2990,In_393,In_745);
nand U2991 (N_2991,In_362,In_1025);
xor U2992 (N_2992,In_120,In_1268);
or U2993 (N_2993,In_697,In_33);
nand U2994 (N_2994,In_1196,In_1363);
nor U2995 (N_2995,In_730,In_20);
or U2996 (N_2996,In_1151,In_1048);
nor U2997 (N_2997,In_424,In_1318);
xor U2998 (N_2998,In_1474,In_1088);
or U2999 (N_2999,In_1246,In_746);
and U3000 (N_3000,In_770,In_1468);
and U3001 (N_3001,In_115,In_662);
or U3002 (N_3002,In_1042,In_556);
xnor U3003 (N_3003,In_789,In_882);
or U3004 (N_3004,In_407,In_429);
xor U3005 (N_3005,In_414,In_527);
and U3006 (N_3006,In_921,In_1031);
or U3007 (N_3007,In_240,In_885);
nand U3008 (N_3008,In_1420,In_348);
xnor U3009 (N_3009,In_0,In_1162);
or U3010 (N_3010,In_400,In_1312);
or U3011 (N_3011,In_1252,In_1203);
or U3012 (N_3012,In_30,In_455);
xnor U3013 (N_3013,In_820,In_300);
nor U3014 (N_3014,In_1065,In_1089);
nor U3015 (N_3015,In_943,In_490);
and U3016 (N_3016,In_595,In_235);
nand U3017 (N_3017,In_593,In_1219);
or U3018 (N_3018,In_109,In_353);
xor U3019 (N_3019,In_1464,In_1039);
and U3020 (N_3020,In_1483,In_736);
nor U3021 (N_3021,In_760,In_239);
or U3022 (N_3022,In_336,In_355);
nand U3023 (N_3023,In_251,In_268);
or U3024 (N_3024,In_900,In_35);
nand U3025 (N_3025,In_1165,In_1407);
and U3026 (N_3026,In_399,In_1320);
or U3027 (N_3027,In_403,In_839);
and U3028 (N_3028,In_402,In_386);
nand U3029 (N_3029,In_1046,In_959);
and U3030 (N_3030,In_955,In_1267);
nor U3031 (N_3031,In_1251,In_1460);
and U3032 (N_3032,In_63,In_30);
and U3033 (N_3033,In_318,In_147);
nor U3034 (N_3034,In_868,In_369);
or U3035 (N_3035,In_1206,In_1393);
nor U3036 (N_3036,In_1254,In_1452);
or U3037 (N_3037,In_957,In_373);
and U3038 (N_3038,In_1091,In_1365);
nor U3039 (N_3039,In_755,In_1131);
nand U3040 (N_3040,In_504,In_906);
and U3041 (N_3041,In_769,In_1180);
nor U3042 (N_3042,In_1200,In_1393);
and U3043 (N_3043,In_626,In_730);
nor U3044 (N_3044,In_638,In_1101);
or U3045 (N_3045,In_1151,In_1261);
nand U3046 (N_3046,In_813,In_118);
or U3047 (N_3047,In_3,In_203);
nor U3048 (N_3048,In_70,In_454);
xnor U3049 (N_3049,In_87,In_1458);
xor U3050 (N_3050,In_1396,In_1237);
nor U3051 (N_3051,In_1090,In_1479);
and U3052 (N_3052,In_875,In_715);
nand U3053 (N_3053,In_1442,In_551);
nor U3054 (N_3054,In_659,In_58);
nor U3055 (N_3055,In_398,In_374);
xnor U3056 (N_3056,In_1305,In_315);
nor U3057 (N_3057,In_168,In_783);
nor U3058 (N_3058,In_580,In_843);
and U3059 (N_3059,In_1203,In_3);
nand U3060 (N_3060,In_554,In_108);
or U3061 (N_3061,In_1152,In_1144);
or U3062 (N_3062,In_781,In_1441);
xnor U3063 (N_3063,In_20,In_452);
or U3064 (N_3064,In_678,In_970);
xor U3065 (N_3065,In_1081,In_1394);
xor U3066 (N_3066,In_485,In_496);
xnor U3067 (N_3067,In_568,In_820);
nand U3068 (N_3068,In_469,In_624);
xor U3069 (N_3069,In_608,In_213);
xor U3070 (N_3070,In_604,In_72);
nor U3071 (N_3071,In_698,In_786);
and U3072 (N_3072,In_954,In_845);
nor U3073 (N_3073,In_1448,In_976);
and U3074 (N_3074,In_1421,In_794);
xor U3075 (N_3075,In_415,In_569);
nand U3076 (N_3076,In_1439,In_40);
nor U3077 (N_3077,In_1242,In_1048);
nand U3078 (N_3078,In_503,In_1142);
and U3079 (N_3079,In_1295,In_866);
or U3080 (N_3080,In_395,In_764);
nand U3081 (N_3081,In_1075,In_1425);
nor U3082 (N_3082,In_114,In_541);
xnor U3083 (N_3083,In_1271,In_497);
nand U3084 (N_3084,In_379,In_198);
and U3085 (N_3085,In_743,In_361);
xor U3086 (N_3086,In_219,In_1223);
nor U3087 (N_3087,In_697,In_377);
or U3088 (N_3088,In_57,In_1415);
nor U3089 (N_3089,In_904,In_816);
nand U3090 (N_3090,In_937,In_970);
nor U3091 (N_3091,In_1251,In_637);
nand U3092 (N_3092,In_1245,In_826);
nand U3093 (N_3093,In_737,In_1000);
or U3094 (N_3094,In_702,In_75);
or U3095 (N_3095,In_1201,In_319);
nand U3096 (N_3096,In_512,In_842);
nand U3097 (N_3097,In_1230,In_924);
and U3098 (N_3098,In_520,In_326);
nor U3099 (N_3099,In_487,In_339);
nand U3100 (N_3100,In_1376,In_918);
nor U3101 (N_3101,In_1492,In_171);
nand U3102 (N_3102,In_654,In_657);
and U3103 (N_3103,In_1398,In_893);
xnor U3104 (N_3104,In_474,In_298);
nand U3105 (N_3105,In_1009,In_775);
nand U3106 (N_3106,In_1259,In_1454);
nand U3107 (N_3107,In_500,In_62);
xor U3108 (N_3108,In_1132,In_202);
nand U3109 (N_3109,In_84,In_1326);
or U3110 (N_3110,In_1283,In_485);
or U3111 (N_3111,In_1470,In_287);
and U3112 (N_3112,In_888,In_782);
nand U3113 (N_3113,In_1326,In_547);
or U3114 (N_3114,In_560,In_9);
nor U3115 (N_3115,In_173,In_363);
or U3116 (N_3116,In_1119,In_1162);
nor U3117 (N_3117,In_442,In_946);
and U3118 (N_3118,In_128,In_1346);
xor U3119 (N_3119,In_986,In_1347);
nand U3120 (N_3120,In_7,In_467);
xnor U3121 (N_3121,In_1138,In_1434);
nand U3122 (N_3122,In_713,In_106);
nor U3123 (N_3123,In_1085,In_555);
nor U3124 (N_3124,In_149,In_320);
nand U3125 (N_3125,In_1309,In_463);
or U3126 (N_3126,In_1103,In_584);
nor U3127 (N_3127,In_285,In_306);
and U3128 (N_3128,In_285,In_1474);
nand U3129 (N_3129,In_1317,In_1478);
xor U3130 (N_3130,In_1267,In_790);
and U3131 (N_3131,In_913,In_184);
and U3132 (N_3132,In_561,In_509);
or U3133 (N_3133,In_323,In_1446);
and U3134 (N_3134,In_1150,In_1129);
and U3135 (N_3135,In_299,In_717);
xor U3136 (N_3136,In_145,In_1034);
and U3137 (N_3137,In_943,In_361);
nand U3138 (N_3138,In_1002,In_1124);
and U3139 (N_3139,In_975,In_1155);
xnor U3140 (N_3140,In_109,In_184);
xor U3141 (N_3141,In_39,In_1440);
nand U3142 (N_3142,In_346,In_44);
and U3143 (N_3143,In_425,In_311);
or U3144 (N_3144,In_1016,In_1196);
xnor U3145 (N_3145,In_1153,In_233);
or U3146 (N_3146,In_940,In_941);
nor U3147 (N_3147,In_1028,In_186);
or U3148 (N_3148,In_943,In_990);
or U3149 (N_3149,In_1096,In_781);
nor U3150 (N_3150,In_338,In_1170);
nand U3151 (N_3151,In_545,In_1356);
and U3152 (N_3152,In_317,In_491);
nand U3153 (N_3153,In_965,In_1425);
nand U3154 (N_3154,In_752,In_134);
or U3155 (N_3155,In_57,In_418);
nor U3156 (N_3156,In_1325,In_613);
and U3157 (N_3157,In_893,In_290);
or U3158 (N_3158,In_526,In_79);
nor U3159 (N_3159,In_240,In_471);
xnor U3160 (N_3160,In_312,In_251);
nor U3161 (N_3161,In_172,In_649);
xnor U3162 (N_3162,In_1074,In_1277);
xor U3163 (N_3163,In_1227,In_1327);
xnor U3164 (N_3164,In_1215,In_1094);
xor U3165 (N_3165,In_1480,In_1053);
nand U3166 (N_3166,In_391,In_768);
nor U3167 (N_3167,In_110,In_451);
or U3168 (N_3168,In_505,In_1047);
nand U3169 (N_3169,In_651,In_274);
or U3170 (N_3170,In_298,In_1080);
nand U3171 (N_3171,In_308,In_639);
and U3172 (N_3172,In_270,In_1022);
and U3173 (N_3173,In_1051,In_1385);
xor U3174 (N_3174,In_246,In_969);
nor U3175 (N_3175,In_313,In_95);
xnor U3176 (N_3176,In_153,In_392);
nand U3177 (N_3177,In_427,In_646);
xor U3178 (N_3178,In_25,In_137);
xnor U3179 (N_3179,In_338,In_53);
xnor U3180 (N_3180,In_91,In_1394);
nor U3181 (N_3181,In_462,In_467);
and U3182 (N_3182,In_566,In_1279);
nand U3183 (N_3183,In_1226,In_1447);
or U3184 (N_3184,In_1073,In_523);
or U3185 (N_3185,In_774,In_1083);
and U3186 (N_3186,In_1250,In_940);
nand U3187 (N_3187,In_483,In_275);
nand U3188 (N_3188,In_244,In_1220);
xnor U3189 (N_3189,In_722,In_665);
nand U3190 (N_3190,In_569,In_344);
xor U3191 (N_3191,In_961,In_1402);
nand U3192 (N_3192,In_596,In_1430);
nor U3193 (N_3193,In_62,In_449);
or U3194 (N_3194,In_1416,In_654);
nand U3195 (N_3195,In_1281,In_387);
nand U3196 (N_3196,In_1239,In_282);
nand U3197 (N_3197,In_510,In_548);
and U3198 (N_3198,In_17,In_1097);
nor U3199 (N_3199,In_693,In_548);
or U3200 (N_3200,In_547,In_490);
nand U3201 (N_3201,In_1488,In_791);
and U3202 (N_3202,In_563,In_2);
xnor U3203 (N_3203,In_1043,In_723);
xor U3204 (N_3204,In_1268,In_1326);
nor U3205 (N_3205,In_824,In_1244);
xor U3206 (N_3206,In_1089,In_84);
nor U3207 (N_3207,In_1193,In_587);
and U3208 (N_3208,In_1127,In_766);
xor U3209 (N_3209,In_1307,In_794);
and U3210 (N_3210,In_216,In_629);
nand U3211 (N_3211,In_304,In_821);
xnor U3212 (N_3212,In_577,In_853);
nand U3213 (N_3213,In_590,In_420);
or U3214 (N_3214,In_945,In_1157);
nand U3215 (N_3215,In_1017,In_1212);
xnor U3216 (N_3216,In_686,In_820);
or U3217 (N_3217,In_503,In_1207);
and U3218 (N_3218,In_829,In_568);
nand U3219 (N_3219,In_1049,In_6);
and U3220 (N_3220,In_1327,In_273);
nand U3221 (N_3221,In_41,In_596);
and U3222 (N_3222,In_713,In_78);
nor U3223 (N_3223,In_998,In_59);
nand U3224 (N_3224,In_1233,In_258);
or U3225 (N_3225,In_1142,In_1012);
nor U3226 (N_3226,In_400,In_1107);
or U3227 (N_3227,In_425,In_270);
or U3228 (N_3228,In_392,In_1138);
and U3229 (N_3229,In_590,In_330);
xor U3230 (N_3230,In_1315,In_664);
nand U3231 (N_3231,In_959,In_1373);
nor U3232 (N_3232,In_877,In_76);
nor U3233 (N_3233,In_1290,In_1212);
and U3234 (N_3234,In_40,In_142);
xor U3235 (N_3235,In_1218,In_114);
nand U3236 (N_3236,In_196,In_1246);
nand U3237 (N_3237,In_246,In_572);
xor U3238 (N_3238,In_1431,In_827);
xor U3239 (N_3239,In_954,In_1048);
or U3240 (N_3240,In_777,In_659);
nor U3241 (N_3241,In_1310,In_598);
or U3242 (N_3242,In_1406,In_1274);
nor U3243 (N_3243,In_199,In_372);
and U3244 (N_3244,In_847,In_513);
nand U3245 (N_3245,In_501,In_854);
or U3246 (N_3246,In_51,In_7);
or U3247 (N_3247,In_1420,In_532);
nor U3248 (N_3248,In_906,In_482);
xnor U3249 (N_3249,In_713,In_116);
nor U3250 (N_3250,In_945,In_1338);
or U3251 (N_3251,In_75,In_804);
nand U3252 (N_3252,In_573,In_310);
nand U3253 (N_3253,In_1350,In_1210);
or U3254 (N_3254,In_1253,In_249);
nor U3255 (N_3255,In_368,In_860);
nor U3256 (N_3256,In_658,In_804);
xnor U3257 (N_3257,In_172,In_652);
nor U3258 (N_3258,In_640,In_664);
xor U3259 (N_3259,In_280,In_43);
nor U3260 (N_3260,In_943,In_443);
or U3261 (N_3261,In_463,In_1337);
xor U3262 (N_3262,In_1443,In_1447);
nand U3263 (N_3263,In_328,In_222);
or U3264 (N_3264,In_1140,In_848);
nor U3265 (N_3265,In_752,In_1227);
or U3266 (N_3266,In_21,In_18);
or U3267 (N_3267,In_663,In_495);
nand U3268 (N_3268,In_477,In_413);
nor U3269 (N_3269,In_127,In_314);
and U3270 (N_3270,In_875,In_451);
xnor U3271 (N_3271,In_468,In_1158);
nor U3272 (N_3272,In_119,In_746);
or U3273 (N_3273,In_1138,In_780);
and U3274 (N_3274,In_466,In_16);
or U3275 (N_3275,In_387,In_1310);
nand U3276 (N_3276,In_1268,In_609);
nor U3277 (N_3277,In_1160,In_48);
nand U3278 (N_3278,In_512,In_495);
nor U3279 (N_3279,In_261,In_1143);
and U3280 (N_3280,In_404,In_82);
and U3281 (N_3281,In_1356,In_241);
xnor U3282 (N_3282,In_425,In_1370);
nand U3283 (N_3283,In_1035,In_1360);
xor U3284 (N_3284,In_1136,In_305);
nand U3285 (N_3285,In_1358,In_285);
or U3286 (N_3286,In_1118,In_885);
nand U3287 (N_3287,In_1444,In_1243);
nor U3288 (N_3288,In_24,In_311);
and U3289 (N_3289,In_442,In_341);
nor U3290 (N_3290,In_621,In_99);
xor U3291 (N_3291,In_1407,In_1246);
and U3292 (N_3292,In_306,In_301);
xor U3293 (N_3293,In_445,In_854);
nor U3294 (N_3294,In_438,In_597);
or U3295 (N_3295,In_826,In_516);
and U3296 (N_3296,In_689,In_870);
nor U3297 (N_3297,In_1460,In_1377);
or U3298 (N_3298,In_810,In_583);
nand U3299 (N_3299,In_1148,In_249);
xnor U3300 (N_3300,In_446,In_534);
xnor U3301 (N_3301,In_83,In_393);
nor U3302 (N_3302,In_335,In_992);
nand U3303 (N_3303,In_908,In_712);
nor U3304 (N_3304,In_453,In_363);
xnor U3305 (N_3305,In_260,In_786);
nand U3306 (N_3306,In_20,In_87);
xnor U3307 (N_3307,In_409,In_1116);
nor U3308 (N_3308,In_550,In_589);
xnor U3309 (N_3309,In_780,In_798);
and U3310 (N_3310,In_1371,In_325);
and U3311 (N_3311,In_210,In_88);
and U3312 (N_3312,In_1360,In_943);
nor U3313 (N_3313,In_809,In_1132);
or U3314 (N_3314,In_1369,In_1048);
xnor U3315 (N_3315,In_752,In_414);
nand U3316 (N_3316,In_1113,In_1110);
and U3317 (N_3317,In_969,In_708);
xor U3318 (N_3318,In_379,In_1185);
nor U3319 (N_3319,In_940,In_1021);
nand U3320 (N_3320,In_742,In_1478);
or U3321 (N_3321,In_988,In_1381);
nor U3322 (N_3322,In_919,In_786);
and U3323 (N_3323,In_285,In_1290);
xnor U3324 (N_3324,In_1329,In_1445);
and U3325 (N_3325,In_35,In_210);
xor U3326 (N_3326,In_411,In_739);
or U3327 (N_3327,In_519,In_1088);
xnor U3328 (N_3328,In_361,In_660);
xor U3329 (N_3329,In_709,In_622);
or U3330 (N_3330,In_967,In_1394);
xor U3331 (N_3331,In_774,In_1328);
nand U3332 (N_3332,In_538,In_504);
nand U3333 (N_3333,In_1261,In_63);
and U3334 (N_3334,In_715,In_317);
nor U3335 (N_3335,In_1399,In_171);
and U3336 (N_3336,In_371,In_123);
or U3337 (N_3337,In_57,In_1437);
nand U3338 (N_3338,In_1385,In_1418);
nand U3339 (N_3339,In_968,In_1145);
nand U3340 (N_3340,In_1237,In_250);
and U3341 (N_3341,In_1420,In_1493);
nand U3342 (N_3342,In_70,In_446);
or U3343 (N_3343,In_58,In_609);
or U3344 (N_3344,In_1421,In_65);
nand U3345 (N_3345,In_336,In_793);
xor U3346 (N_3346,In_1092,In_287);
and U3347 (N_3347,In_1026,In_1121);
nand U3348 (N_3348,In_1171,In_926);
nand U3349 (N_3349,In_144,In_1139);
or U3350 (N_3350,In_469,In_1223);
xnor U3351 (N_3351,In_1408,In_503);
nor U3352 (N_3352,In_644,In_948);
and U3353 (N_3353,In_89,In_497);
xor U3354 (N_3354,In_1455,In_515);
and U3355 (N_3355,In_323,In_1272);
xnor U3356 (N_3356,In_73,In_439);
or U3357 (N_3357,In_834,In_1440);
xor U3358 (N_3358,In_297,In_755);
nor U3359 (N_3359,In_1209,In_74);
or U3360 (N_3360,In_962,In_255);
nor U3361 (N_3361,In_890,In_1063);
nor U3362 (N_3362,In_209,In_775);
or U3363 (N_3363,In_621,In_469);
nor U3364 (N_3364,In_1344,In_756);
and U3365 (N_3365,In_633,In_1246);
xor U3366 (N_3366,In_1417,In_738);
nand U3367 (N_3367,In_1394,In_908);
and U3368 (N_3368,In_290,In_76);
or U3369 (N_3369,In_894,In_1123);
nand U3370 (N_3370,In_39,In_1181);
and U3371 (N_3371,In_449,In_1218);
and U3372 (N_3372,In_363,In_287);
nand U3373 (N_3373,In_0,In_1243);
and U3374 (N_3374,In_1321,In_1194);
xnor U3375 (N_3375,In_1063,In_1218);
nand U3376 (N_3376,In_1094,In_116);
xor U3377 (N_3377,In_122,In_492);
xor U3378 (N_3378,In_865,In_122);
and U3379 (N_3379,In_1051,In_825);
nand U3380 (N_3380,In_520,In_118);
xor U3381 (N_3381,In_580,In_825);
nand U3382 (N_3382,In_264,In_690);
nor U3383 (N_3383,In_1177,In_487);
nor U3384 (N_3384,In_978,In_850);
nor U3385 (N_3385,In_630,In_377);
nand U3386 (N_3386,In_56,In_1332);
nor U3387 (N_3387,In_1400,In_405);
xor U3388 (N_3388,In_1315,In_252);
nor U3389 (N_3389,In_947,In_1330);
nand U3390 (N_3390,In_703,In_620);
or U3391 (N_3391,In_1429,In_254);
and U3392 (N_3392,In_365,In_901);
and U3393 (N_3393,In_244,In_537);
xnor U3394 (N_3394,In_563,In_1254);
xnor U3395 (N_3395,In_65,In_702);
nor U3396 (N_3396,In_266,In_816);
and U3397 (N_3397,In_1162,In_349);
and U3398 (N_3398,In_566,In_982);
nor U3399 (N_3399,In_388,In_243);
nor U3400 (N_3400,In_424,In_1422);
nor U3401 (N_3401,In_1380,In_58);
xor U3402 (N_3402,In_1147,In_768);
and U3403 (N_3403,In_105,In_430);
xor U3404 (N_3404,In_897,In_416);
nand U3405 (N_3405,In_1010,In_20);
or U3406 (N_3406,In_823,In_1322);
xor U3407 (N_3407,In_596,In_217);
nand U3408 (N_3408,In_1360,In_1437);
xnor U3409 (N_3409,In_889,In_793);
or U3410 (N_3410,In_118,In_1308);
xor U3411 (N_3411,In_351,In_771);
xor U3412 (N_3412,In_1136,In_1144);
or U3413 (N_3413,In_189,In_464);
and U3414 (N_3414,In_379,In_676);
nand U3415 (N_3415,In_1027,In_1256);
nor U3416 (N_3416,In_465,In_217);
nand U3417 (N_3417,In_847,In_1209);
and U3418 (N_3418,In_269,In_863);
nor U3419 (N_3419,In_1047,In_900);
xor U3420 (N_3420,In_1444,In_92);
nor U3421 (N_3421,In_858,In_535);
and U3422 (N_3422,In_632,In_1002);
or U3423 (N_3423,In_1485,In_192);
or U3424 (N_3424,In_936,In_1271);
or U3425 (N_3425,In_389,In_1);
nor U3426 (N_3426,In_998,In_198);
nor U3427 (N_3427,In_1407,In_124);
nand U3428 (N_3428,In_1481,In_906);
nor U3429 (N_3429,In_158,In_514);
xnor U3430 (N_3430,In_103,In_608);
and U3431 (N_3431,In_1484,In_1009);
and U3432 (N_3432,In_740,In_165);
xor U3433 (N_3433,In_946,In_1418);
nor U3434 (N_3434,In_70,In_220);
xnor U3435 (N_3435,In_409,In_176);
nand U3436 (N_3436,In_1129,In_535);
xor U3437 (N_3437,In_974,In_1417);
nand U3438 (N_3438,In_1195,In_61);
xnor U3439 (N_3439,In_1249,In_541);
nand U3440 (N_3440,In_189,In_1025);
xnor U3441 (N_3441,In_376,In_895);
xnor U3442 (N_3442,In_1418,In_729);
nand U3443 (N_3443,In_3,In_437);
nor U3444 (N_3444,In_1423,In_37);
nand U3445 (N_3445,In_220,In_855);
nand U3446 (N_3446,In_1456,In_557);
nor U3447 (N_3447,In_1425,In_388);
nand U3448 (N_3448,In_264,In_377);
nand U3449 (N_3449,In_27,In_509);
and U3450 (N_3450,In_322,In_1441);
or U3451 (N_3451,In_360,In_851);
or U3452 (N_3452,In_315,In_506);
and U3453 (N_3453,In_1195,In_1068);
and U3454 (N_3454,In_737,In_1313);
xor U3455 (N_3455,In_768,In_1400);
nor U3456 (N_3456,In_1112,In_588);
or U3457 (N_3457,In_256,In_1213);
nor U3458 (N_3458,In_1219,In_87);
nor U3459 (N_3459,In_485,In_1403);
nor U3460 (N_3460,In_131,In_394);
nor U3461 (N_3461,In_24,In_469);
or U3462 (N_3462,In_1068,In_1305);
nor U3463 (N_3463,In_1392,In_1356);
nand U3464 (N_3464,In_1482,In_527);
xor U3465 (N_3465,In_652,In_368);
or U3466 (N_3466,In_246,In_1115);
or U3467 (N_3467,In_210,In_750);
nand U3468 (N_3468,In_20,In_190);
or U3469 (N_3469,In_650,In_86);
or U3470 (N_3470,In_850,In_113);
or U3471 (N_3471,In_678,In_182);
xnor U3472 (N_3472,In_829,In_1079);
nand U3473 (N_3473,In_100,In_553);
or U3474 (N_3474,In_1342,In_456);
nand U3475 (N_3475,In_1031,In_218);
nand U3476 (N_3476,In_1142,In_1437);
nor U3477 (N_3477,In_275,In_228);
or U3478 (N_3478,In_218,In_1238);
nor U3479 (N_3479,In_948,In_235);
nor U3480 (N_3480,In_228,In_1118);
nand U3481 (N_3481,In_1227,In_253);
nand U3482 (N_3482,In_742,In_872);
or U3483 (N_3483,In_32,In_1399);
or U3484 (N_3484,In_1158,In_522);
or U3485 (N_3485,In_1001,In_955);
nand U3486 (N_3486,In_1308,In_1120);
nand U3487 (N_3487,In_748,In_161);
xor U3488 (N_3488,In_994,In_13);
and U3489 (N_3489,In_125,In_1131);
xnor U3490 (N_3490,In_1355,In_350);
nor U3491 (N_3491,In_107,In_789);
and U3492 (N_3492,In_1009,In_577);
and U3493 (N_3493,In_664,In_1339);
xor U3494 (N_3494,In_837,In_653);
and U3495 (N_3495,In_467,In_612);
nor U3496 (N_3496,In_211,In_691);
nor U3497 (N_3497,In_201,In_582);
xnor U3498 (N_3498,In_153,In_794);
nand U3499 (N_3499,In_557,In_611);
nor U3500 (N_3500,In_1019,In_1086);
nor U3501 (N_3501,In_692,In_874);
xnor U3502 (N_3502,In_438,In_476);
nand U3503 (N_3503,In_858,In_999);
nor U3504 (N_3504,In_8,In_444);
and U3505 (N_3505,In_904,In_526);
xnor U3506 (N_3506,In_1308,In_165);
xnor U3507 (N_3507,In_1388,In_1031);
and U3508 (N_3508,In_877,In_1312);
and U3509 (N_3509,In_84,In_222);
and U3510 (N_3510,In_142,In_1257);
or U3511 (N_3511,In_1230,In_1409);
xnor U3512 (N_3512,In_1483,In_809);
or U3513 (N_3513,In_1161,In_1303);
xnor U3514 (N_3514,In_1090,In_574);
nand U3515 (N_3515,In_1420,In_228);
nor U3516 (N_3516,In_1401,In_832);
xor U3517 (N_3517,In_1403,In_184);
and U3518 (N_3518,In_1194,In_1167);
xnor U3519 (N_3519,In_5,In_1478);
xor U3520 (N_3520,In_373,In_344);
nand U3521 (N_3521,In_1257,In_500);
or U3522 (N_3522,In_1102,In_760);
nand U3523 (N_3523,In_785,In_770);
xnor U3524 (N_3524,In_351,In_967);
xnor U3525 (N_3525,In_15,In_956);
nand U3526 (N_3526,In_85,In_1193);
xor U3527 (N_3527,In_721,In_102);
and U3528 (N_3528,In_698,In_199);
nor U3529 (N_3529,In_444,In_345);
nand U3530 (N_3530,In_912,In_1007);
and U3531 (N_3531,In_202,In_398);
nor U3532 (N_3532,In_504,In_794);
nand U3533 (N_3533,In_1152,In_327);
or U3534 (N_3534,In_1367,In_986);
xnor U3535 (N_3535,In_933,In_444);
or U3536 (N_3536,In_330,In_960);
and U3537 (N_3537,In_331,In_1315);
xnor U3538 (N_3538,In_814,In_1479);
nor U3539 (N_3539,In_1166,In_796);
nor U3540 (N_3540,In_662,In_1303);
or U3541 (N_3541,In_1146,In_162);
and U3542 (N_3542,In_710,In_815);
and U3543 (N_3543,In_852,In_764);
nor U3544 (N_3544,In_392,In_1298);
xor U3545 (N_3545,In_670,In_1345);
nand U3546 (N_3546,In_350,In_809);
or U3547 (N_3547,In_250,In_735);
nor U3548 (N_3548,In_288,In_593);
nor U3549 (N_3549,In_821,In_1450);
or U3550 (N_3550,In_1021,In_282);
or U3551 (N_3551,In_262,In_344);
nand U3552 (N_3552,In_2,In_1289);
xnor U3553 (N_3553,In_1323,In_1484);
or U3554 (N_3554,In_881,In_905);
xnor U3555 (N_3555,In_582,In_438);
nor U3556 (N_3556,In_1479,In_535);
or U3557 (N_3557,In_198,In_1266);
nor U3558 (N_3558,In_459,In_862);
or U3559 (N_3559,In_1274,In_1017);
and U3560 (N_3560,In_1278,In_1050);
nor U3561 (N_3561,In_515,In_672);
or U3562 (N_3562,In_482,In_665);
or U3563 (N_3563,In_920,In_198);
and U3564 (N_3564,In_226,In_540);
nand U3565 (N_3565,In_1373,In_152);
nand U3566 (N_3566,In_1209,In_279);
or U3567 (N_3567,In_332,In_170);
nor U3568 (N_3568,In_1120,In_1156);
or U3569 (N_3569,In_246,In_123);
xor U3570 (N_3570,In_426,In_1231);
xnor U3571 (N_3571,In_1161,In_1061);
and U3572 (N_3572,In_906,In_1313);
nor U3573 (N_3573,In_1119,In_1381);
nor U3574 (N_3574,In_557,In_115);
or U3575 (N_3575,In_19,In_1130);
or U3576 (N_3576,In_1381,In_439);
xor U3577 (N_3577,In_1289,In_982);
or U3578 (N_3578,In_617,In_300);
and U3579 (N_3579,In_216,In_424);
nor U3580 (N_3580,In_772,In_174);
nor U3581 (N_3581,In_807,In_1137);
or U3582 (N_3582,In_147,In_408);
and U3583 (N_3583,In_780,In_133);
nand U3584 (N_3584,In_351,In_1346);
or U3585 (N_3585,In_1206,In_858);
or U3586 (N_3586,In_417,In_943);
nand U3587 (N_3587,In_340,In_269);
nor U3588 (N_3588,In_603,In_1278);
or U3589 (N_3589,In_482,In_858);
or U3590 (N_3590,In_1409,In_1211);
nor U3591 (N_3591,In_449,In_263);
nor U3592 (N_3592,In_544,In_183);
xnor U3593 (N_3593,In_512,In_1133);
nand U3594 (N_3594,In_344,In_1429);
nand U3595 (N_3595,In_1071,In_1275);
xor U3596 (N_3596,In_20,In_575);
xnor U3597 (N_3597,In_201,In_1367);
nor U3598 (N_3598,In_320,In_336);
or U3599 (N_3599,In_787,In_855);
xnor U3600 (N_3600,In_1465,In_1428);
nand U3601 (N_3601,In_1116,In_653);
nand U3602 (N_3602,In_865,In_1106);
nand U3603 (N_3603,In_276,In_101);
and U3604 (N_3604,In_1001,In_636);
nor U3605 (N_3605,In_1157,In_846);
nor U3606 (N_3606,In_1152,In_275);
xnor U3607 (N_3607,In_1015,In_1469);
xor U3608 (N_3608,In_1071,In_643);
and U3609 (N_3609,In_563,In_631);
nand U3610 (N_3610,In_1477,In_1487);
or U3611 (N_3611,In_1236,In_1006);
nor U3612 (N_3612,In_634,In_287);
and U3613 (N_3613,In_1323,In_891);
xor U3614 (N_3614,In_855,In_1306);
nor U3615 (N_3615,In_85,In_1021);
nand U3616 (N_3616,In_1223,In_1303);
nand U3617 (N_3617,In_294,In_775);
nand U3618 (N_3618,In_439,In_1489);
and U3619 (N_3619,In_344,In_961);
and U3620 (N_3620,In_298,In_784);
nor U3621 (N_3621,In_1463,In_1071);
and U3622 (N_3622,In_1334,In_1389);
nor U3623 (N_3623,In_14,In_1495);
nor U3624 (N_3624,In_859,In_244);
xnor U3625 (N_3625,In_1042,In_7);
or U3626 (N_3626,In_563,In_738);
nor U3627 (N_3627,In_16,In_246);
and U3628 (N_3628,In_504,In_1045);
or U3629 (N_3629,In_1032,In_1358);
and U3630 (N_3630,In_455,In_54);
nand U3631 (N_3631,In_1140,In_439);
and U3632 (N_3632,In_183,In_1071);
nand U3633 (N_3633,In_676,In_185);
and U3634 (N_3634,In_1232,In_224);
nand U3635 (N_3635,In_775,In_943);
xor U3636 (N_3636,In_1274,In_597);
and U3637 (N_3637,In_569,In_730);
nand U3638 (N_3638,In_65,In_1278);
and U3639 (N_3639,In_1461,In_1207);
or U3640 (N_3640,In_686,In_782);
xor U3641 (N_3641,In_779,In_1216);
xnor U3642 (N_3642,In_1458,In_1008);
xor U3643 (N_3643,In_1223,In_484);
nor U3644 (N_3644,In_511,In_1222);
nand U3645 (N_3645,In_1209,In_405);
nor U3646 (N_3646,In_51,In_340);
or U3647 (N_3647,In_158,In_836);
xor U3648 (N_3648,In_414,In_1089);
nand U3649 (N_3649,In_403,In_1028);
or U3650 (N_3650,In_95,In_191);
nand U3651 (N_3651,In_1035,In_1123);
nand U3652 (N_3652,In_1313,In_1327);
and U3653 (N_3653,In_1103,In_603);
nor U3654 (N_3654,In_1376,In_193);
nor U3655 (N_3655,In_1013,In_296);
and U3656 (N_3656,In_1336,In_321);
nor U3657 (N_3657,In_1119,In_14);
xnor U3658 (N_3658,In_803,In_24);
xnor U3659 (N_3659,In_947,In_1185);
or U3660 (N_3660,In_224,In_110);
and U3661 (N_3661,In_241,In_757);
or U3662 (N_3662,In_1299,In_49);
xnor U3663 (N_3663,In_1117,In_1123);
xor U3664 (N_3664,In_1460,In_1005);
nand U3665 (N_3665,In_1389,In_19);
and U3666 (N_3666,In_716,In_793);
or U3667 (N_3667,In_181,In_879);
xnor U3668 (N_3668,In_353,In_577);
nor U3669 (N_3669,In_1067,In_3);
nor U3670 (N_3670,In_121,In_793);
nor U3671 (N_3671,In_1475,In_232);
or U3672 (N_3672,In_1174,In_847);
xor U3673 (N_3673,In_1013,In_1077);
nor U3674 (N_3674,In_46,In_62);
xor U3675 (N_3675,In_1269,In_95);
nor U3676 (N_3676,In_1253,In_1175);
or U3677 (N_3677,In_911,In_153);
nand U3678 (N_3678,In_209,In_9);
nand U3679 (N_3679,In_236,In_1043);
and U3680 (N_3680,In_787,In_1255);
nor U3681 (N_3681,In_76,In_1232);
nor U3682 (N_3682,In_777,In_1018);
xnor U3683 (N_3683,In_979,In_1187);
nand U3684 (N_3684,In_1272,In_469);
nor U3685 (N_3685,In_1464,In_490);
xnor U3686 (N_3686,In_712,In_255);
nor U3687 (N_3687,In_126,In_4);
or U3688 (N_3688,In_1499,In_1323);
and U3689 (N_3689,In_968,In_576);
xnor U3690 (N_3690,In_1146,In_1479);
xor U3691 (N_3691,In_878,In_214);
and U3692 (N_3692,In_613,In_421);
nor U3693 (N_3693,In_1094,In_948);
nand U3694 (N_3694,In_1264,In_508);
nor U3695 (N_3695,In_87,In_560);
nor U3696 (N_3696,In_643,In_1205);
xor U3697 (N_3697,In_942,In_923);
and U3698 (N_3698,In_1124,In_918);
xnor U3699 (N_3699,In_768,In_1158);
nand U3700 (N_3700,In_387,In_616);
xor U3701 (N_3701,In_176,In_187);
nor U3702 (N_3702,In_872,In_521);
xnor U3703 (N_3703,In_605,In_751);
xnor U3704 (N_3704,In_773,In_475);
and U3705 (N_3705,In_527,In_896);
or U3706 (N_3706,In_737,In_475);
nand U3707 (N_3707,In_1268,In_981);
or U3708 (N_3708,In_218,In_1111);
nand U3709 (N_3709,In_1259,In_1381);
and U3710 (N_3710,In_891,In_34);
nand U3711 (N_3711,In_557,In_285);
xor U3712 (N_3712,In_498,In_1149);
and U3713 (N_3713,In_1426,In_1317);
nor U3714 (N_3714,In_1325,In_705);
nand U3715 (N_3715,In_194,In_1394);
and U3716 (N_3716,In_1340,In_822);
or U3717 (N_3717,In_886,In_1212);
nand U3718 (N_3718,In_1194,In_488);
and U3719 (N_3719,In_464,In_1387);
nand U3720 (N_3720,In_1165,In_369);
xnor U3721 (N_3721,In_822,In_1404);
xor U3722 (N_3722,In_731,In_1419);
or U3723 (N_3723,In_89,In_1193);
xor U3724 (N_3724,In_719,In_345);
xnor U3725 (N_3725,In_1116,In_1377);
xnor U3726 (N_3726,In_538,In_555);
and U3727 (N_3727,In_182,In_209);
xor U3728 (N_3728,In_865,In_1467);
nor U3729 (N_3729,In_1397,In_248);
nand U3730 (N_3730,In_1278,In_172);
and U3731 (N_3731,In_1225,In_706);
or U3732 (N_3732,In_1002,In_264);
xor U3733 (N_3733,In_601,In_445);
or U3734 (N_3734,In_1193,In_915);
and U3735 (N_3735,In_592,In_1141);
xor U3736 (N_3736,In_837,In_898);
nand U3737 (N_3737,In_624,In_550);
nor U3738 (N_3738,In_594,In_1031);
xor U3739 (N_3739,In_218,In_1038);
xor U3740 (N_3740,In_1388,In_1126);
xor U3741 (N_3741,In_819,In_161);
and U3742 (N_3742,In_432,In_567);
or U3743 (N_3743,In_241,In_1200);
or U3744 (N_3744,In_784,In_1348);
nand U3745 (N_3745,In_47,In_1164);
nor U3746 (N_3746,In_1145,In_10);
nand U3747 (N_3747,In_56,In_143);
nor U3748 (N_3748,In_1269,In_14);
or U3749 (N_3749,In_1195,In_82);
nor U3750 (N_3750,In_655,In_1274);
and U3751 (N_3751,In_661,In_1289);
or U3752 (N_3752,In_876,In_316);
or U3753 (N_3753,In_1021,In_1479);
nand U3754 (N_3754,In_334,In_1399);
nand U3755 (N_3755,In_220,In_351);
nor U3756 (N_3756,In_895,In_480);
or U3757 (N_3757,In_1010,In_562);
nand U3758 (N_3758,In_497,In_357);
or U3759 (N_3759,In_1006,In_1303);
and U3760 (N_3760,In_1121,In_881);
or U3761 (N_3761,In_425,In_645);
xor U3762 (N_3762,In_690,In_15);
and U3763 (N_3763,In_1175,In_576);
or U3764 (N_3764,In_1316,In_378);
and U3765 (N_3765,In_239,In_298);
nor U3766 (N_3766,In_1316,In_1084);
nor U3767 (N_3767,In_665,In_1059);
or U3768 (N_3768,In_631,In_1063);
nor U3769 (N_3769,In_782,In_991);
nor U3770 (N_3770,In_466,In_582);
nand U3771 (N_3771,In_1163,In_1115);
or U3772 (N_3772,In_603,In_1085);
and U3773 (N_3773,In_774,In_922);
and U3774 (N_3774,In_15,In_1384);
and U3775 (N_3775,In_1453,In_586);
or U3776 (N_3776,In_15,In_179);
or U3777 (N_3777,In_991,In_506);
nand U3778 (N_3778,In_1411,In_181);
nand U3779 (N_3779,In_1490,In_554);
and U3780 (N_3780,In_1454,In_1287);
xnor U3781 (N_3781,In_496,In_330);
nor U3782 (N_3782,In_664,In_888);
and U3783 (N_3783,In_511,In_1118);
nor U3784 (N_3784,In_1481,In_554);
nor U3785 (N_3785,In_667,In_556);
nand U3786 (N_3786,In_1390,In_786);
or U3787 (N_3787,In_899,In_406);
xnor U3788 (N_3788,In_198,In_383);
xnor U3789 (N_3789,In_116,In_1483);
xor U3790 (N_3790,In_1238,In_12);
nor U3791 (N_3791,In_257,In_458);
nor U3792 (N_3792,In_1343,In_149);
xor U3793 (N_3793,In_223,In_396);
or U3794 (N_3794,In_1147,In_1368);
nor U3795 (N_3795,In_144,In_1085);
and U3796 (N_3796,In_1042,In_305);
or U3797 (N_3797,In_355,In_1141);
or U3798 (N_3798,In_218,In_641);
xor U3799 (N_3799,In_739,In_567);
nand U3800 (N_3800,In_1136,In_1343);
or U3801 (N_3801,In_1419,In_999);
nand U3802 (N_3802,In_986,In_164);
and U3803 (N_3803,In_541,In_606);
or U3804 (N_3804,In_1105,In_452);
nor U3805 (N_3805,In_535,In_610);
xor U3806 (N_3806,In_801,In_977);
and U3807 (N_3807,In_1266,In_856);
xnor U3808 (N_3808,In_1228,In_546);
and U3809 (N_3809,In_322,In_1293);
or U3810 (N_3810,In_1364,In_1457);
or U3811 (N_3811,In_1276,In_1401);
nand U3812 (N_3812,In_781,In_227);
nor U3813 (N_3813,In_331,In_1415);
nor U3814 (N_3814,In_382,In_439);
xor U3815 (N_3815,In_1069,In_967);
or U3816 (N_3816,In_458,In_881);
or U3817 (N_3817,In_349,In_250);
nor U3818 (N_3818,In_1228,In_94);
or U3819 (N_3819,In_408,In_619);
nor U3820 (N_3820,In_1456,In_1414);
nor U3821 (N_3821,In_1052,In_949);
nand U3822 (N_3822,In_15,In_456);
nor U3823 (N_3823,In_378,In_622);
and U3824 (N_3824,In_1235,In_1018);
nor U3825 (N_3825,In_1145,In_169);
xor U3826 (N_3826,In_946,In_287);
or U3827 (N_3827,In_1032,In_1248);
xor U3828 (N_3828,In_271,In_286);
and U3829 (N_3829,In_199,In_87);
nor U3830 (N_3830,In_248,In_1186);
or U3831 (N_3831,In_304,In_68);
nor U3832 (N_3832,In_615,In_798);
nor U3833 (N_3833,In_625,In_148);
or U3834 (N_3834,In_572,In_761);
or U3835 (N_3835,In_80,In_1449);
and U3836 (N_3836,In_1456,In_1191);
or U3837 (N_3837,In_201,In_161);
or U3838 (N_3838,In_4,In_1343);
xnor U3839 (N_3839,In_831,In_1163);
nor U3840 (N_3840,In_1424,In_94);
nor U3841 (N_3841,In_365,In_803);
and U3842 (N_3842,In_318,In_57);
nor U3843 (N_3843,In_11,In_793);
or U3844 (N_3844,In_521,In_389);
xnor U3845 (N_3845,In_342,In_59);
and U3846 (N_3846,In_500,In_1188);
or U3847 (N_3847,In_1418,In_866);
or U3848 (N_3848,In_1395,In_1045);
and U3849 (N_3849,In_266,In_140);
and U3850 (N_3850,In_235,In_943);
nor U3851 (N_3851,In_360,In_551);
xor U3852 (N_3852,In_152,In_939);
or U3853 (N_3853,In_1230,In_30);
nand U3854 (N_3854,In_19,In_813);
nor U3855 (N_3855,In_110,In_1231);
xor U3856 (N_3856,In_886,In_627);
and U3857 (N_3857,In_437,In_200);
xnor U3858 (N_3858,In_761,In_1307);
or U3859 (N_3859,In_1237,In_30);
and U3860 (N_3860,In_1434,In_649);
nand U3861 (N_3861,In_808,In_1192);
nand U3862 (N_3862,In_178,In_1328);
or U3863 (N_3863,In_684,In_406);
nor U3864 (N_3864,In_278,In_783);
or U3865 (N_3865,In_524,In_550);
nor U3866 (N_3866,In_869,In_71);
nor U3867 (N_3867,In_185,In_900);
nand U3868 (N_3868,In_249,In_448);
nor U3869 (N_3869,In_779,In_449);
or U3870 (N_3870,In_1271,In_1065);
xnor U3871 (N_3871,In_43,In_506);
xor U3872 (N_3872,In_1221,In_146);
or U3873 (N_3873,In_717,In_832);
nor U3874 (N_3874,In_1241,In_279);
and U3875 (N_3875,In_717,In_380);
nand U3876 (N_3876,In_1085,In_1025);
or U3877 (N_3877,In_491,In_1210);
nor U3878 (N_3878,In_888,In_576);
or U3879 (N_3879,In_818,In_727);
nand U3880 (N_3880,In_1037,In_1345);
nand U3881 (N_3881,In_767,In_1382);
xor U3882 (N_3882,In_778,In_1334);
nor U3883 (N_3883,In_1045,In_670);
or U3884 (N_3884,In_998,In_853);
nor U3885 (N_3885,In_399,In_570);
nor U3886 (N_3886,In_680,In_1429);
xnor U3887 (N_3887,In_777,In_834);
nand U3888 (N_3888,In_696,In_140);
nor U3889 (N_3889,In_5,In_1228);
xor U3890 (N_3890,In_955,In_746);
nor U3891 (N_3891,In_508,In_263);
nand U3892 (N_3892,In_940,In_1497);
and U3893 (N_3893,In_778,In_432);
nor U3894 (N_3894,In_230,In_586);
and U3895 (N_3895,In_1091,In_70);
nand U3896 (N_3896,In_997,In_1278);
nand U3897 (N_3897,In_363,In_1354);
xnor U3898 (N_3898,In_864,In_43);
xnor U3899 (N_3899,In_1454,In_746);
xnor U3900 (N_3900,In_448,In_220);
nand U3901 (N_3901,In_335,In_283);
and U3902 (N_3902,In_397,In_1005);
nand U3903 (N_3903,In_707,In_942);
xor U3904 (N_3904,In_162,In_1489);
nor U3905 (N_3905,In_705,In_315);
nor U3906 (N_3906,In_761,In_104);
or U3907 (N_3907,In_1079,In_1406);
xor U3908 (N_3908,In_737,In_1367);
xor U3909 (N_3909,In_738,In_1058);
nor U3910 (N_3910,In_738,In_557);
nand U3911 (N_3911,In_103,In_943);
nand U3912 (N_3912,In_4,In_952);
and U3913 (N_3913,In_78,In_1038);
or U3914 (N_3914,In_1130,In_159);
or U3915 (N_3915,In_402,In_647);
or U3916 (N_3916,In_577,In_422);
nor U3917 (N_3917,In_831,In_807);
or U3918 (N_3918,In_318,In_752);
nor U3919 (N_3919,In_854,In_305);
nand U3920 (N_3920,In_1229,In_303);
nand U3921 (N_3921,In_598,In_309);
xnor U3922 (N_3922,In_1032,In_615);
nor U3923 (N_3923,In_439,In_150);
and U3924 (N_3924,In_894,In_785);
nor U3925 (N_3925,In_1205,In_1034);
nand U3926 (N_3926,In_163,In_432);
nor U3927 (N_3927,In_439,In_43);
nand U3928 (N_3928,In_155,In_1475);
xor U3929 (N_3929,In_1197,In_554);
xnor U3930 (N_3930,In_146,In_418);
nor U3931 (N_3931,In_318,In_153);
or U3932 (N_3932,In_328,In_173);
nor U3933 (N_3933,In_996,In_591);
and U3934 (N_3934,In_1206,In_68);
nor U3935 (N_3935,In_433,In_122);
nor U3936 (N_3936,In_187,In_1379);
nor U3937 (N_3937,In_124,In_687);
or U3938 (N_3938,In_1278,In_486);
and U3939 (N_3939,In_1241,In_129);
xor U3940 (N_3940,In_882,In_553);
or U3941 (N_3941,In_440,In_1154);
nand U3942 (N_3942,In_669,In_997);
nor U3943 (N_3943,In_582,In_285);
nand U3944 (N_3944,In_818,In_770);
nand U3945 (N_3945,In_182,In_282);
and U3946 (N_3946,In_466,In_1018);
nand U3947 (N_3947,In_578,In_1343);
and U3948 (N_3948,In_132,In_1486);
and U3949 (N_3949,In_246,In_974);
and U3950 (N_3950,In_803,In_1251);
and U3951 (N_3951,In_402,In_650);
xnor U3952 (N_3952,In_769,In_617);
nand U3953 (N_3953,In_867,In_190);
or U3954 (N_3954,In_377,In_456);
xnor U3955 (N_3955,In_1079,In_619);
xor U3956 (N_3956,In_449,In_195);
nand U3957 (N_3957,In_1414,In_1478);
nand U3958 (N_3958,In_1138,In_87);
nor U3959 (N_3959,In_1352,In_1420);
nor U3960 (N_3960,In_1463,In_299);
nand U3961 (N_3961,In_482,In_1021);
or U3962 (N_3962,In_1155,In_1237);
xnor U3963 (N_3963,In_907,In_1234);
nand U3964 (N_3964,In_1003,In_1017);
nand U3965 (N_3965,In_1360,In_162);
or U3966 (N_3966,In_1175,In_1448);
nor U3967 (N_3967,In_1172,In_1255);
nor U3968 (N_3968,In_644,In_278);
and U3969 (N_3969,In_170,In_1074);
and U3970 (N_3970,In_1192,In_1275);
and U3971 (N_3971,In_734,In_752);
or U3972 (N_3972,In_1051,In_994);
nand U3973 (N_3973,In_946,In_527);
nand U3974 (N_3974,In_1348,In_746);
nand U3975 (N_3975,In_359,In_526);
or U3976 (N_3976,In_735,In_453);
or U3977 (N_3977,In_897,In_719);
xor U3978 (N_3978,In_483,In_1107);
and U3979 (N_3979,In_1148,In_767);
nand U3980 (N_3980,In_252,In_1442);
nand U3981 (N_3981,In_136,In_412);
nand U3982 (N_3982,In_247,In_1159);
or U3983 (N_3983,In_60,In_391);
nor U3984 (N_3984,In_1396,In_683);
or U3985 (N_3985,In_126,In_605);
nor U3986 (N_3986,In_768,In_648);
nand U3987 (N_3987,In_268,In_675);
nor U3988 (N_3988,In_731,In_92);
and U3989 (N_3989,In_1429,In_992);
or U3990 (N_3990,In_1375,In_552);
and U3991 (N_3991,In_1335,In_129);
and U3992 (N_3992,In_782,In_832);
xor U3993 (N_3993,In_428,In_1021);
xor U3994 (N_3994,In_912,In_1269);
nor U3995 (N_3995,In_1309,In_286);
and U3996 (N_3996,In_1035,In_1057);
xnor U3997 (N_3997,In_1212,In_861);
or U3998 (N_3998,In_247,In_968);
and U3999 (N_3999,In_1107,In_36);
nor U4000 (N_4000,In_966,In_449);
or U4001 (N_4001,In_1239,In_1345);
nand U4002 (N_4002,In_1191,In_834);
nor U4003 (N_4003,In_1242,In_1376);
nor U4004 (N_4004,In_317,In_347);
xnor U4005 (N_4005,In_1183,In_306);
nor U4006 (N_4006,In_782,In_977);
xor U4007 (N_4007,In_309,In_1444);
or U4008 (N_4008,In_192,In_1492);
xnor U4009 (N_4009,In_1486,In_399);
xor U4010 (N_4010,In_1105,In_128);
and U4011 (N_4011,In_599,In_873);
xnor U4012 (N_4012,In_1085,In_1402);
or U4013 (N_4013,In_317,In_567);
and U4014 (N_4014,In_487,In_758);
or U4015 (N_4015,In_1470,In_1404);
and U4016 (N_4016,In_178,In_629);
or U4017 (N_4017,In_647,In_1056);
and U4018 (N_4018,In_921,In_707);
or U4019 (N_4019,In_699,In_690);
xor U4020 (N_4020,In_1492,In_424);
nor U4021 (N_4021,In_1329,In_327);
and U4022 (N_4022,In_1120,In_65);
or U4023 (N_4023,In_999,In_1312);
nand U4024 (N_4024,In_1448,In_410);
nor U4025 (N_4025,In_768,In_106);
nand U4026 (N_4026,In_667,In_5);
nand U4027 (N_4027,In_1366,In_175);
nor U4028 (N_4028,In_1327,In_341);
nor U4029 (N_4029,In_1158,In_693);
and U4030 (N_4030,In_17,In_641);
nor U4031 (N_4031,In_744,In_1153);
nor U4032 (N_4032,In_633,In_500);
and U4033 (N_4033,In_1310,In_1128);
or U4034 (N_4034,In_1328,In_230);
or U4035 (N_4035,In_968,In_113);
nor U4036 (N_4036,In_468,In_136);
or U4037 (N_4037,In_1051,In_449);
xor U4038 (N_4038,In_146,In_855);
nor U4039 (N_4039,In_843,In_630);
or U4040 (N_4040,In_79,In_368);
nand U4041 (N_4041,In_1029,In_1062);
nand U4042 (N_4042,In_747,In_559);
xor U4043 (N_4043,In_1191,In_465);
and U4044 (N_4044,In_1067,In_1010);
and U4045 (N_4045,In_835,In_1315);
xor U4046 (N_4046,In_949,In_711);
or U4047 (N_4047,In_1440,In_738);
xor U4048 (N_4048,In_165,In_1339);
nand U4049 (N_4049,In_1490,In_688);
nand U4050 (N_4050,In_1034,In_459);
or U4051 (N_4051,In_984,In_1092);
nor U4052 (N_4052,In_799,In_560);
or U4053 (N_4053,In_1171,In_79);
nand U4054 (N_4054,In_694,In_872);
and U4055 (N_4055,In_946,In_1103);
xor U4056 (N_4056,In_1313,In_1404);
or U4057 (N_4057,In_800,In_81);
nor U4058 (N_4058,In_1250,In_988);
and U4059 (N_4059,In_717,In_528);
xnor U4060 (N_4060,In_666,In_1433);
or U4061 (N_4061,In_449,In_541);
nor U4062 (N_4062,In_1016,In_1450);
xnor U4063 (N_4063,In_520,In_497);
and U4064 (N_4064,In_1074,In_1406);
nand U4065 (N_4065,In_24,In_557);
nand U4066 (N_4066,In_154,In_1207);
and U4067 (N_4067,In_1160,In_615);
and U4068 (N_4068,In_1232,In_216);
nand U4069 (N_4069,In_592,In_70);
xor U4070 (N_4070,In_63,In_878);
nand U4071 (N_4071,In_590,In_426);
or U4072 (N_4072,In_126,In_682);
and U4073 (N_4073,In_365,In_1416);
nand U4074 (N_4074,In_238,In_717);
nand U4075 (N_4075,In_705,In_707);
nor U4076 (N_4076,In_817,In_1201);
xor U4077 (N_4077,In_791,In_971);
nor U4078 (N_4078,In_136,In_1213);
or U4079 (N_4079,In_211,In_27);
nand U4080 (N_4080,In_1443,In_1047);
or U4081 (N_4081,In_290,In_566);
or U4082 (N_4082,In_914,In_370);
or U4083 (N_4083,In_1080,In_183);
nand U4084 (N_4084,In_337,In_149);
nand U4085 (N_4085,In_105,In_131);
nand U4086 (N_4086,In_909,In_1414);
nand U4087 (N_4087,In_487,In_811);
or U4088 (N_4088,In_883,In_87);
nand U4089 (N_4089,In_1360,In_249);
or U4090 (N_4090,In_1480,In_1141);
nor U4091 (N_4091,In_992,In_642);
or U4092 (N_4092,In_1212,In_1032);
xor U4093 (N_4093,In_1491,In_1244);
xor U4094 (N_4094,In_327,In_1181);
and U4095 (N_4095,In_409,In_1);
and U4096 (N_4096,In_782,In_956);
or U4097 (N_4097,In_765,In_947);
nand U4098 (N_4098,In_866,In_224);
xor U4099 (N_4099,In_803,In_210);
nor U4100 (N_4100,In_1436,In_408);
xor U4101 (N_4101,In_537,In_844);
and U4102 (N_4102,In_570,In_98);
xor U4103 (N_4103,In_711,In_653);
or U4104 (N_4104,In_113,In_339);
or U4105 (N_4105,In_1485,In_491);
nand U4106 (N_4106,In_1125,In_545);
or U4107 (N_4107,In_91,In_1165);
or U4108 (N_4108,In_541,In_1433);
and U4109 (N_4109,In_1234,In_50);
nor U4110 (N_4110,In_871,In_125);
nand U4111 (N_4111,In_1193,In_395);
and U4112 (N_4112,In_403,In_334);
or U4113 (N_4113,In_604,In_1261);
nand U4114 (N_4114,In_1001,In_501);
xor U4115 (N_4115,In_1124,In_831);
xnor U4116 (N_4116,In_84,In_802);
nand U4117 (N_4117,In_104,In_887);
or U4118 (N_4118,In_41,In_1276);
xor U4119 (N_4119,In_57,In_1032);
nor U4120 (N_4120,In_1096,In_269);
and U4121 (N_4121,In_1261,In_326);
nand U4122 (N_4122,In_269,In_223);
nor U4123 (N_4123,In_1339,In_1084);
nor U4124 (N_4124,In_676,In_1189);
nand U4125 (N_4125,In_588,In_127);
xor U4126 (N_4126,In_182,In_1276);
and U4127 (N_4127,In_1155,In_227);
xor U4128 (N_4128,In_287,In_575);
or U4129 (N_4129,In_406,In_1408);
and U4130 (N_4130,In_420,In_179);
xor U4131 (N_4131,In_887,In_1063);
and U4132 (N_4132,In_410,In_1312);
nand U4133 (N_4133,In_317,In_750);
or U4134 (N_4134,In_843,In_691);
nor U4135 (N_4135,In_1064,In_1287);
and U4136 (N_4136,In_1412,In_1348);
nand U4137 (N_4137,In_699,In_1073);
xor U4138 (N_4138,In_326,In_621);
and U4139 (N_4139,In_679,In_172);
nor U4140 (N_4140,In_1116,In_1388);
xnor U4141 (N_4141,In_615,In_1377);
xor U4142 (N_4142,In_550,In_677);
or U4143 (N_4143,In_1025,In_428);
nand U4144 (N_4144,In_444,In_264);
and U4145 (N_4145,In_1435,In_1228);
and U4146 (N_4146,In_207,In_271);
nand U4147 (N_4147,In_1162,In_776);
nor U4148 (N_4148,In_97,In_930);
xor U4149 (N_4149,In_839,In_1171);
or U4150 (N_4150,In_1367,In_702);
nand U4151 (N_4151,In_426,In_112);
xor U4152 (N_4152,In_687,In_838);
xnor U4153 (N_4153,In_661,In_342);
xnor U4154 (N_4154,In_58,In_858);
or U4155 (N_4155,In_171,In_637);
or U4156 (N_4156,In_421,In_499);
nand U4157 (N_4157,In_1050,In_1123);
and U4158 (N_4158,In_1234,In_204);
and U4159 (N_4159,In_713,In_1184);
xor U4160 (N_4160,In_293,In_1408);
xnor U4161 (N_4161,In_208,In_41);
or U4162 (N_4162,In_194,In_368);
nand U4163 (N_4163,In_284,In_261);
xor U4164 (N_4164,In_413,In_1151);
or U4165 (N_4165,In_427,In_287);
or U4166 (N_4166,In_720,In_52);
xnor U4167 (N_4167,In_81,In_366);
and U4168 (N_4168,In_832,In_939);
nand U4169 (N_4169,In_1323,In_1449);
and U4170 (N_4170,In_462,In_1271);
or U4171 (N_4171,In_627,In_823);
xor U4172 (N_4172,In_831,In_1423);
and U4173 (N_4173,In_518,In_645);
nor U4174 (N_4174,In_1492,In_893);
nor U4175 (N_4175,In_1351,In_1031);
nor U4176 (N_4176,In_311,In_534);
nor U4177 (N_4177,In_682,In_1335);
or U4178 (N_4178,In_426,In_296);
or U4179 (N_4179,In_138,In_50);
or U4180 (N_4180,In_1030,In_608);
nand U4181 (N_4181,In_791,In_1175);
and U4182 (N_4182,In_321,In_1257);
and U4183 (N_4183,In_1363,In_317);
nand U4184 (N_4184,In_1486,In_1065);
nand U4185 (N_4185,In_986,In_558);
or U4186 (N_4186,In_522,In_1362);
and U4187 (N_4187,In_558,In_818);
xnor U4188 (N_4188,In_772,In_390);
xor U4189 (N_4189,In_1464,In_927);
or U4190 (N_4190,In_150,In_1006);
nor U4191 (N_4191,In_1211,In_1166);
and U4192 (N_4192,In_576,In_799);
xor U4193 (N_4193,In_42,In_1371);
nand U4194 (N_4194,In_803,In_281);
nand U4195 (N_4195,In_34,In_1358);
or U4196 (N_4196,In_1092,In_323);
nand U4197 (N_4197,In_1371,In_1153);
nor U4198 (N_4198,In_1444,In_815);
xor U4199 (N_4199,In_69,In_445);
nor U4200 (N_4200,In_133,In_898);
nand U4201 (N_4201,In_190,In_384);
and U4202 (N_4202,In_645,In_835);
or U4203 (N_4203,In_901,In_810);
and U4204 (N_4204,In_458,In_388);
nand U4205 (N_4205,In_675,In_1035);
and U4206 (N_4206,In_1265,In_552);
or U4207 (N_4207,In_570,In_444);
or U4208 (N_4208,In_626,In_1199);
xor U4209 (N_4209,In_1382,In_919);
nand U4210 (N_4210,In_1454,In_506);
and U4211 (N_4211,In_1272,In_914);
or U4212 (N_4212,In_349,In_1005);
xnor U4213 (N_4213,In_951,In_1013);
nand U4214 (N_4214,In_301,In_443);
nand U4215 (N_4215,In_1492,In_1345);
nand U4216 (N_4216,In_1197,In_421);
nand U4217 (N_4217,In_389,In_608);
nor U4218 (N_4218,In_1341,In_364);
or U4219 (N_4219,In_374,In_565);
nand U4220 (N_4220,In_813,In_77);
nand U4221 (N_4221,In_1287,In_902);
or U4222 (N_4222,In_128,In_924);
and U4223 (N_4223,In_365,In_471);
and U4224 (N_4224,In_1307,In_979);
xor U4225 (N_4225,In_247,In_627);
nor U4226 (N_4226,In_725,In_643);
nand U4227 (N_4227,In_771,In_960);
xor U4228 (N_4228,In_931,In_854);
or U4229 (N_4229,In_310,In_1436);
or U4230 (N_4230,In_855,In_646);
xor U4231 (N_4231,In_90,In_1084);
or U4232 (N_4232,In_520,In_1252);
and U4233 (N_4233,In_1022,In_516);
or U4234 (N_4234,In_37,In_1263);
xnor U4235 (N_4235,In_343,In_548);
and U4236 (N_4236,In_158,In_242);
and U4237 (N_4237,In_1265,In_868);
or U4238 (N_4238,In_69,In_14);
nor U4239 (N_4239,In_465,In_962);
and U4240 (N_4240,In_1400,In_1011);
or U4241 (N_4241,In_904,In_1125);
xnor U4242 (N_4242,In_1477,In_918);
nor U4243 (N_4243,In_1090,In_222);
or U4244 (N_4244,In_792,In_214);
and U4245 (N_4245,In_446,In_151);
nor U4246 (N_4246,In_190,In_780);
xor U4247 (N_4247,In_1382,In_1496);
nor U4248 (N_4248,In_189,In_1247);
nor U4249 (N_4249,In_784,In_966);
xnor U4250 (N_4250,In_935,In_272);
nand U4251 (N_4251,In_520,In_1406);
nand U4252 (N_4252,In_629,In_852);
nor U4253 (N_4253,In_967,In_253);
nand U4254 (N_4254,In_746,In_1384);
and U4255 (N_4255,In_1490,In_557);
and U4256 (N_4256,In_1171,In_296);
or U4257 (N_4257,In_727,In_1294);
and U4258 (N_4258,In_390,In_1161);
nand U4259 (N_4259,In_1018,In_117);
nor U4260 (N_4260,In_106,In_208);
and U4261 (N_4261,In_273,In_675);
or U4262 (N_4262,In_39,In_937);
xnor U4263 (N_4263,In_774,In_255);
and U4264 (N_4264,In_1157,In_798);
nor U4265 (N_4265,In_985,In_427);
nand U4266 (N_4266,In_282,In_669);
or U4267 (N_4267,In_665,In_1037);
nand U4268 (N_4268,In_844,In_594);
nand U4269 (N_4269,In_702,In_552);
or U4270 (N_4270,In_101,In_591);
nand U4271 (N_4271,In_173,In_64);
nor U4272 (N_4272,In_773,In_1082);
xnor U4273 (N_4273,In_51,In_1002);
xnor U4274 (N_4274,In_575,In_1128);
and U4275 (N_4275,In_1441,In_839);
nor U4276 (N_4276,In_260,In_426);
nand U4277 (N_4277,In_472,In_1170);
or U4278 (N_4278,In_957,In_1347);
nor U4279 (N_4279,In_1429,In_510);
and U4280 (N_4280,In_1495,In_862);
or U4281 (N_4281,In_879,In_1439);
nand U4282 (N_4282,In_642,In_568);
nor U4283 (N_4283,In_167,In_1497);
nand U4284 (N_4284,In_1366,In_126);
and U4285 (N_4285,In_1004,In_619);
nor U4286 (N_4286,In_1283,In_1197);
or U4287 (N_4287,In_1379,In_202);
xnor U4288 (N_4288,In_1233,In_1176);
and U4289 (N_4289,In_1257,In_713);
or U4290 (N_4290,In_68,In_1063);
or U4291 (N_4291,In_325,In_792);
nand U4292 (N_4292,In_959,In_317);
xor U4293 (N_4293,In_829,In_240);
and U4294 (N_4294,In_626,In_16);
nand U4295 (N_4295,In_1013,In_653);
nor U4296 (N_4296,In_1216,In_564);
or U4297 (N_4297,In_1084,In_656);
and U4298 (N_4298,In_991,In_311);
nand U4299 (N_4299,In_1408,In_414);
xor U4300 (N_4300,In_210,In_835);
or U4301 (N_4301,In_1239,In_854);
nor U4302 (N_4302,In_1046,In_1380);
nand U4303 (N_4303,In_856,In_759);
and U4304 (N_4304,In_1096,In_602);
nor U4305 (N_4305,In_1236,In_31);
xnor U4306 (N_4306,In_1175,In_187);
nand U4307 (N_4307,In_1330,In_1011);
or U4308 (N_4308,In_644,In_732);
nor U4309 (N_4309,In_69,In_588);
xnor U4310 (N_4310,In_648,In_857);
xnor U4311 (N_4311,In_960,In_433);
nor U4312 (N_4312,In_1380,In_395);
or U4313 (N_4313,In_441,In_163);
and U4314 (N_4314,In_310,In_1159);
xor U4315 (N_4315,In_1374,In_231);
nand U4316 (N_4316,In_1478,In_705);
or U4317 (N_4317,In_453,In_90);
or U4318 (N_4318,In_352,In_636);
nor U4319 (N_4319,In_692,In_179);
or U4320 (N_4320,In_1136,In_521);
and U4321 (N_4321,In_945,In_385);
or U4322 (N_4322,In_1096,In_425);
nand U4323 (N_4323,In_1032,In_111);
xor U4324 (N_4324,In_49,In_660);
or U4325 (N_4325,In_253,In_672);
xor U4326 (N_4326,In_123,In_977);
nor U4327 (N_4327,In_1116,In_782);
or U4328 (N_4328,In_46,In_813);
nand U4329 (N_4329,In_159,In_699);
and U4330 (N_4330,In_586,In_1354);
xor U4331 (N_4331,In_1432,In_565);
nand U4332 (N_4332,In_699,In_820);
and U4333 (N_4333,In_513,In_1137);
and U4334 (N_4334,In_329,In_286);
and U4335 (N_4335,In_1103,In_314);
nor U4336 (N_4336,In_892,In_1194);
xor U4337 (N_4337,In_437,In_372);
xor U4338 (N_4338,In_1139,In_1491);
nor U4339 (N_4339,In_1079,In_1044);
xor U4340 (N_4340,In_50,In_859);
xnor U4341 (N_4341,In_1248,In_873);
nor U4342 (N_4342,In_1086,In_1071);
xnor U4343 (N_4343,In_460,In_1440);
or U4344 (N_4344,In_531,In_85);
or U4345 (N_4345,In_594,In_586);
and U4346 (N_4346,In_1075,In_562);
nand U4347 (N_4347,In_1459,In_826);
nor U4348 (N_4348,In_1389,In_97);
and U4349 (N_4349,In_1139,In_1269);
xnor U4350 (N_4350,In_423,In_1325);
nor U4351 (N_4351,In_132,In_682);
xor U4352 (N_4352,In_467,In_842);
nand U4353 (N_4353,In_1232,In_205);
xor U4354 (N_4354,In_1429,In_1316);
nand U4355 (N_4355,In_1476,In_659);
or U4356 (N_4356,In_352,In_1281);
xnor U4357 (N_4357,In_480,In_162);
xnor U4358 (N_4358,In_142,In_433);
xnor U4359 (N_4359,In_830,In_625);
nand U4360 (N_4360,In_508,In_682);
and U4361 (N_4361,In_1134,In_64);
nand U4362 (N_4362,In_965,In_623);
or U4363 (N_4363,In_744,In_150);
xor U4364 (N_4364,In_864,In_298);
nor U4365 (N_4365,In_453,In_517);
or U4366 (N_4366,In_1251,In_449);
or U4367 (N_4367,In_1087,In_605);
or U4368 (N_4368,In_1391,In_407);
and U4369 (N_4369,In_113,In_1026);
and U4370 (N_4370,In_1479,In_569);
nor U4371 (N_4371,In_861,In_1009);
nor U4372 (N_4372,In_1475,In_450);
nor U4373 (N_4373,In_1378,In_1436);
nand U4374 (N_4374,In_859,In_1334);
nand U4375 (N_4375,In_1042,In_790);
and U4376 (N_4376,In_892,In_237);
xor U4377 (N_4377,In_952,In_1486);
nor U4378 (N_4378,In_1230,In_1235);
or U4379 (N_4379,In_1089,In_1221);
nor U4380 (N_4380,In_228,In_824);
and U4381 (N_4381,In_780,In_888);
nand U4382 (N_4382,In_258,In_640);
or U4383 (N_4383,In_767,In_170);
or U4384 (N_4384,In_1239,In_349);
or U4385 (N_4385,In_1060,In_1394);
xor U4386 (N_4386,In_1179,In_15);
or U4387 (N_4387,In_1322,In_504);
nor U4388 (N_4388,In_1009,In_78);
and U4389 (N_4389,In_1144,In_857);
or U4390 (N_4390,In_574,In_1020);
xnor U4391 (N_4391,In_809,In_810);
nor U4392 (N_4392,In_468,In_508);
and U4393 (N_4393,In_879,In_150);
and U4394 (N_4394,In_1338,In_698);
xor U4395 (N_4395,In_1156,In_1320);
or U4396 (N_4396,In_1025,In_248);
nand U4397 (N_4397,In_1213,In_877);
and U4398 (N_4398,In_296,In_1049);
and U4399 (N_4399,In_1001,In_650);
nand U4400 (N_4400,In_1139,In_1040);
or U4401 (N_4401,In_1457,In_795);
or U4402 (N_4402,In_427,In_239);
nand U4403 (N_4403,In_1065,In_287);
and U4404 (N_4404,In_1225,In_741);
or U4405 (N_4405,In_75,In_76);
nand U4406 (N_4406,In_771,In_515);
and U4407 (N_4407,In_824,In_125);
nor U4408 (N_4408,In_937,In_87);
nand U4409 (N_4409,In_1412,In_647);
nand U4410 (N_4410,In_585,In_203);
or U4411 (N_4411,In_1359,In_1383);
and U4412 (N_4412,In_1251,In_1196);
xnor U4413 (N_4413,In_25,In_488);
and U4414 (N_4414,In_60,In_932);
and U4415 (N_4415,In_1027,In_144);
nand U4416 (N_4416,In_1311,In_920);
nand U4417 (N_4417,In_842,In_487);
nor U4418 (N_4418,In_883,In_1379);
nand U4419 (N_4419,In_424,In_1103);
nand U4420 (N_4420,In_330,In_1387);
or U4421 (N_4421,In_185,In_248);
and U4422 (N_4422,In_353,In_1496);
nand U4423 (N_4423,In_829,In_861);
and U4424 (N_4424,In_1177,In_353);
nor U4425 (N_4425,In_1393,In_1467);
or U4426 (N_4426,In_758,In_204);
or U4427 (N_4427,In_808,In_890);
and U4428 (N_4428,In_981,In_994);
nand U4429 (N_4429,In_1148,In_1047);
xor U4430 (N_4430,In_714,In_1074);
and U4431 (N_4431,In_248,In_732);
nand U4432 (N_4432,In_739,In_1434);
xor U4433 (N_4433,In_268,In_1217);
or U4434 (N_4434,In_412,In_283);
nor U4435 (N_4435,In_173,In_763);
nor U4436 (N_4436,In_1106,In_159);
and U4437 (N_4437,In_57,In_445);
or U4438 (N_4438,In_981,In_222);
and U4439 (N_4439,In_454,In_418);
nand U4440 (N_4440,In_15,In_1184);
nor U4441 (N_4441,In_1216,In_1085);
or U4442 (N_4442,In_716,In_788);
xnor U4443 (N_4443,In_954,In_553);
nand U4444 (N_4444,In_990,In_713);
nor U4445 (N_4445,In_462,In_729);
or U4446 (N_4446,In_893,In_709);
nor U4447 (N_4447,In_510,In_729);
and U4448 (N_4448,In_1161,In_1488);
xnor U4449 (N_4449,In_501,In_149);
or U4450 (N_4450,In_292,In_47);
nor U4451 (N_4451,In_654,In_338);
and U4452 (N_4452,In_1221,In_58);
or U4453 (N_4453,In_417,In_460);
nand U4454 (N_4454,In_309,In_1178);
nor U4455 (N_4455,In_464,In_474);
and U4456 (N_4456,In_874,In_87);
or U4457 (N_4457,In_1316,In_1234);
and U4458 (N_4458,In_552,In_169);
and U4459 (N_4459,In_727,In_986);
nor U4460 (N_4460,In_604,In_1359);
xor U4461 (N_4461,In_97,In_958);
and U4462 (N_4462,In_1368,In_1148);
or U4463 (N_4463,In_1487,In_933);
nor U4464 (N_4464,In_818,In_1055);
xnor U4465 (N_4465,In_103,In_319);
and U4466 (N_4466,In_1020,In_1045);
xor U4467 (N_4467,In_101,In_1459);
nor U4468 (N_4468,In_154,In_440);
xnor U4469 (N_4469,In_536,In_144);
and U4470 (N_4470,In_449,In_1145);
or U4471 (N_4471,In_1283,In_412);
or U4472 (N_4472,In_321,In_222);
xor U4473 (N_4473,In_482,In_889);
and U4474 (N_4474,In_303,In_845);
or U4475 (N_4475,In_1086,In_1281);
nand U4476 (N_4476,In_1042,In_1195);
and U4477 (N_4477,In_1074,In_584);
or U4478 (N_4478,In_1330,In_362);
nor U4479 (N_4479,In_424,In_752);
xor U4480 (N_4480,In_519,In_1416);
or U4481 (N_4481,In_599,In_469);
xnor U4482 (N_4482,In_422,In_761);
nand U4483 (N_4483,In_1495,In_1259);
or U4484 (N_4484,In_1338,In_329);
nor U4485 (N_4485,In_195,In_991);
nand U4486 (N_4486,In_1495,In_90);
nor U4487 (N_4487,In_1157,In_1431);
nand U4488 (N_4488,In_411,In_1283);
or U4489 (N_4489,In_1102,In_759);
and U4490 (N_4490,In_869,In_1006);
nand U4491 (N_4491,In_783,In_1090);
or U4492 (N_4492,In_412,In_1466);
nor U4493 (N_4493,In_1312,In_1311);
or U4494 (N_4494,In_1161,In_187);
nor U4495 (N_4495,In_234,In_1108);
nor U4496 (N_4496,In_645,In_988);
xor U4497 (N_4497,In_679,In_174);
or U4498 (N_4498,In_1356,In_1235);
nand U4499 (N_4499,In_1348,In_1036);
xor U4500 (N_4500,In_19,In_187);
and U4501 (N_4501,In_127,In_31);
nand U4502 (N_4502,In_1380,In_275);
or U4503 (N_4503,In_370,In_113);
nor U4504 (N_4504,In_181,In_1455);
xnor U4505 (N_4505,In_1008,In_736);
xnor U4506 (N_4506,In_851,In_83);
nor U4507 (N_4507,In_393,In_604);
nor U4508 (N_4508,In_1238,In_775);
nor U4509 (N_4509,In_1072,In_1403);
and U4510 (N_4510,In_877,In_403);
nor U4511 (N_4511,In_762,In_1176);
nand U4512 (N_4512,In_5,In_1211);
or U4513 (N_4513,In_1493,In_271);
or U4514 (N_4514,In_1049,In_1072);
and U4515 (N_4515,In_434,In_350);
nand U4516 (N_4516,In_783,In_842);
or U4517 (N_4517,In_871,In_495);
nand U4518 (N_4518,In_1276,In_1317);
nand U4519 (N_4519,In_1368,In_1119);
and U4520 (N_4520,In_574,In_109);
and U4521 (N_4521,In_883,In_468);
nor U4522 (N_4522,In_576,In_1105);
nor U4523 (N_4523,In_1307,In_1136);
or U4524 (N_4524,In_20,In_365);
or U4525 (N_4525,In_637,In_60);
and U4526 (N_4526,In_40,In_160);
xor U4527 (N_4527,In_1070,In_1040);
or U4528 (N_4528,In_865,In_286);
nor U4529 (N_4529,In_1310,In_824);
nor U4530 (N_4530,In_359,In_977);
nand U4531 (N_4531,In_166,In_878);
and U4532 (N_4532,In_870,In_992);
xor U4533 (N_4533,In_167,In_719);
nand U4534 (N_4534,In_378,In_957);
and U4535 (N_4535,In_562,In_1308);
and U4536 (N_4536,In_983,In_500);
xor U4537 (N_4537,In_903,In_289);
nor U4538 (N_4538,In_841,In_685);
and U4539 (N_4539,In_206,In_610);
and U4540 (N_4540,In_825,In_1332);
xnor U4541 (N_4541,In_239,In_682);
nand U4542 (N_4542,In_1380,In_741);
xnor U4543 (N_4543,In_609,In_448);
nor U4544 (N_4544,In_630,In_502);
or U4545 (N_4545,In_232,In_6);
xnor U4546 (N_4546,In_25,In_1085);
or U4547 (N_4547,In_1002,In_324);
or U4548 (N_4548,In_373,In_1447);
and U4549 (N_4549,In_139,In_764);
xor U4550 (N_4550,In_1274,In_563);
nor U4551 (N_4551,In_728,In_1434);
nor U4552 (N_4552,In_239,In_440);
xor U4553 (N_4553,In_1062,In_407);
xnor U4554 (N_4554,In_273,In_1353);
or U4555 (N_4555,In_195,In_209);
nor U4556 (N_4556,In_540,In_534);
nand U4557 (N_4557,In_996,In_318);
nor U4558 (N_4558,In_916,In_842);
nor U4559 (N_4559,In_977,In_1290);
nor U4560 (N_4560,In_526,In_1043);
xnor U4561 (N_4561,In_1189,In_555);
xor U4562 (N_4562,In_838,In_968);
and U4563 (N_4563,In_743,In_247);
and U4564 (N_4564,In_676,In_1074);
or U4565 (N_4565,In_754,In_211);
or U4566 (N_4566,In_1214,In_571);
or U4567 (N_4567,In_798,In_497);
or U4568 (N_4568,In_286,In_1127);
nand U4569 (N_4569,In_989,In_1138);
nor U4570 (N_4570,In_1083,In_1061);
nor U4571 (N_4571,In_992,In_362);
nor U4572 (N_4572,In_369,In_437);
or U4573 (N_4573,In_675,In_139);
and U4574 (N_4574,In_514,In_746);
xnor U4575 (N_4575,In_201,In_269);
or U4576 (N_4576,In_149,In_1131);
nor U4577 (N_4577,In_807,In_1185);
xor U4578 (N_4578,In_731,In_839);
or U4579 (N_4579,In_931,In_938);
xor U4580 (N_4580,In_528,In_1072);
and U4581 (N_4581,In_1173,In_1240);
nand U4582 (N_4582,In_1111,In_735);
nand U4583 (N_4583,In_313,In_1042);
xnor U4584 (N_4584,In_1075,In_1041);
nor U4585 (N_4585,In_204,In_49);
and U4586 (N_4586,In_252,In_1385);
nand U4587 (N_4587,In_1362,In_1368);
and U4588 (N_4588,In_238,In_587);
nand U4589 (N_4589,In_531,In_1339);
and U4590 (N_4590,In_354,In_1434);
xnor U4591 (N_4591,In_76,In_733);
nor U4592 (N_4592,In_1407,In_418);
nor U4593 (N_4593,In_795,In_456);
xnor U4594 (N_4594,In_999,In_690);
nand U4595 (N_4595,In_696,In_953);
or U4596 (N_4596,In_605,In_1438);
nand U4597 (N_4597,In_355,In_1307);
nand U4598 (N_4598,In_310,In_1433);
and U4599 (N_4599,In_668,In_1440);
and U4600 (N_4600,In_691,In_605);
nor U4601 (N_4601,In_1407,In_571);
nand U4602 (N_4602,In_665,In_245);
xnor U4603 (N_4603,In_480,In_1027);
nor U4604 (N_4604,In_1420,In_946);
nor U4605 (N_4605,In_1151,In_382);
nand U4606 (N_4606,In_45,In_406);
or U4607 (N_4607,In_1196,In_1068);
and U4608 (N_4608,In_489,In_820);
or U4609 (N_4609,In_221,In_1480);
or U4610 (N_4610,In_813,In_1137);
or U4611 (N_4611,In_273,In_1056);
and U4612 (N_4612,In_580,In_1237);
or U4613 (N_4613,In_354,In_38);
nor U4614 (N_4614,In_296,In_793);
or U4615 (N_4615,In_877,In_97);
or U4616 (N_4616,In_298,In_1239);
nand U4617 (N_4617,In_1287,In_1316);
xor U4618 (N_4618,In_55,In_1129);
nor U4619 (N_4619,In_564,In_609);
or U4620 (N_4620,In_1350,In_1062);
and U4621 (N_4621,In_244,In_238);
nand U4622 (N_4622,In_433,In_510);
nand U4623 (N_4623,In_906,In_833);
nand U4624 (N_4624,In_666,In_187);
nor U4625 (N_4625,In_1379,In_552);
xnor U4626 (N_4626,In_1007,In_488);
xor U4627 (N_4627,In_182,In_615);
nand U4628 (N_4628,In_1324,In_449);
and U4629 (N_4629,In_1287,In_727);
nor U4630 (N_4630,In_500,In_1198);
nand U4631 (N_4631,In_1487,In_360);
nor U4632 (N_4632,In_768,In_630);
and U4633 (N_4633,In_1490,In_944);
or U4634 (N_4634,In_536,In_1439);
or U4635 (N_4635,In_584,In_1350);
or U4636 (N_4636,In_527,In_293);
xnor U4637 (N_4637,In_327,In_541);
nor U4638 (N_4638,In_495,In_551);
nor U4639 (N_4639,In_1170,In_130);
xnor U4640 (N_4640,In_418,In_667);
or U4641 (N_4641,In_27,In_461);
xnor U4642 (N_4642,In_1026,In_1331);
nand U4643 (N_4643,In_270,In_1000);
nor U4644 (N_4644,In_1277,In_872);
and U4645 (N_4645,In_605,In_834);
xor U4646 (N_4646,In_699,In_413);
and U4647 (N_4647,In_1357,In_661);
and U4648 (N_4648,In_745,In_918);
nand U4649 (N_4649,In_1283,In_1140);
or U4650 (N_4650,In_1187,In_219);
xnor U4651 (N_4651,In_362,In_876);
or U4652 (N_4652,In_895,In_1401);
nand U4653 (N_4653,In_38,In_559);
or U4654 (N_4654,In_117,In_1165);
or U4655 (N_4655,In_499,In_1188);
nor U4656 (N_4656,In_541,In_1375);
xor U4657 (N_4657,In_387,In_864);
xnor U4658 (N_4658,In_1424,In_498);
and U4659 (N_4659,In_23,In_1341);
and U4660 (N_4660,In_919,In_912);
or U4661 (N_4661,In_437,In_1151);
and U4662 (N_4662,In_1139,In_312);
xnor U4663 (N_4663,In_698,In_1144);
xor U4664 (N_4664,In_185,In_888);
nand U4665 (N_4665,In_379,In_1350);
or U4666 (N_4666,In_925,In_1031);
or U4667 (N_4667,In_982,In_775);
nor U4668 (N_4668,In_835,In_844);
xor U4669 (N_4669,In_1199,In_1445);
and U4670 (N_4670,In_500,In_1018);
or U4671 (N_4671,In_41,In_1190);
xnor U4672 (N_4672,In_738,In_1077);
nor U4673 (N_4673,In_1327,In_1256);
nor U4674 (N_4674,In_987,In_979);
or U4675 (N_4675,In_553,In_1154);
or U4676 (N_4676,In_1151,In_1416);
xor U4677 (N_4677,In_315,In_462);
xnor U4678 (N_4678,In_542,In_709);
and U4679 (N_4679,In_229,In_732);
xor U4680 (N_4680,In_1218,In_1183);
or U4681 (N_4681,In_1335,In_1381);
xnor U4682 (N_4682,In_174,In_705);
xnor U4683 (N_4683,In_5,In_859);
nand U4684 (N_4684,In_1268,In_623);
or U4685 (N_4685,In_175,In_1193);
or U4686 (N_4686,In_906,In_153);
nor U4687 (N_4687,In_1247,In_1430);
nor U4688 (N_4688,In_1356,In_1398);
and U4689 (N_4689,In_107,In_1264);
and U4690 (N_4690,In_1467,In_1456);
nor U4691 (N_4691,In_676,In_36);
nor U4692 (N_4692,In_1300,In_1243);
nor U4693 (N_4693,In_530,In_20);
nor U4694 (N_4694,In_415,In_307);
nand U4695 (N_4695,In_1140,In_78);
and U4696 (N_4696,In_403,In_210);
and U4697 (N_4697,In_795,In_568);
or U4698 (N_4698,In_1411,In_443);
xor U4699 (N_4699,In_677,In_418);
and U4700 (N_4700,In_320,In_324);
xor U4701 (N_4701,In_300,In_1207);
xor U4702 (N_4702,In_340,In_925);
or U4703 (N_4703,In_933,In_1252);
nand U4704 (N_4704,In_760,In_5);
xor U4705 (N_4705,In_735,In_1012);
nor U4706 (N_4706,In_452,In_1338);
xnor U4707 (N_4707,In_505,In_159);
nor U4708 (N_4708,In_1254,In_185);
or U4709 (N_4709,In_225,In_690);
nand U4710 (N_4710,In_1259,In_1167);
xor U4711 (N_4711,In_1168,In_1064);
or U4712 (N_4712,In_311,In_1086);
or U4713 (N_4713,In_727,In_1175);
nand U4714 (N_4714,In_893,In_1406);
or U4715 (N_4715,In_1159,In_79);
nor U4716 (N_4716,In_774,In_390);
xnor U4717 (N_4717,In_415,In_82);
and U4718 (N_4718,In_472,In_573);
and U4719 (N_4719,In_1047,In_908);
and U4720 (N_4720,In_975,In_1207);
or U4721 (N_4721,In_746,In_943);
nand U4722 (N_4722,In_1039,In_1032);
nor U4723 (N_4723,In_109,In_972);
or U4724 (N_4724,In_1313,In_1385);
or U4725 (N_4725,In_1009,In_22);
nand U4726 (N_4726,In_274,In_760);
or U4727 (N_4727,In_1414,In_211);
nor U4728 (N_4728,In_218,In_763);
xor U4729 (N_4729,In_1283,In_778);
nand U4730 (N_4730,In_339,In_1054);
and U4731 (N_4731,In_541,In_908);
nor U4732 (N_4732,In_354,In_747);
or U4733 (N_4733,In_372,In_506);
xor U4734 (N_4734,In_276,In_204);
xnor U4735 (N_4735,In_451,In_322);
nor U4736 (N_4736,In_1198,In_466);
nand U4737 (N_4737,In_482,In_74);
and U4738 (N_4738,In_296,In_336);
nand U4739 (N_4739,In_137,In_705);
and U4740 (N_4740,In_1209,In_1040);
and U4741 (N_4741,In_1057,In_1442);
and U4742 (N_4742,In_469,In_336);
nand U4743 (N_4743,In_7,In_1211);
xor U4744 (N_4744,In_5,In_1456);
nor U4745 (N_4745,In_1429,In_1418);
nor U4746 (N_4746,In_845,In_1306);
xnor U4747 (N_4747,In_520,In_338);
nor U4748 (N_4748,In_1078,In_784);
nor U4749 (N_4749,In_597,In_612);
xor U4750 (N_4750,In_698,In_1195);
or U4751 (N_4751,In_1186,In_1445);
nor U4752 (N_4752,In_616,In_1036);
nor U4753 (N_4753,In_567,In_157);
nand U4754 (N_4754,In_224,In_654);
nand U4755 (N_4755,In_1054,In_1372);
nand U4756 (N_4756,In_1088,In_760);
xor U4757 (N_4757,In_689,In_149);
nor U4758 (N_4758,In_757,In_495);
or U4759 (N_4759,In_1226,In_616);
xnor U4760 (N_4760,In_600,In_185);
xor U4761 (N_4761,In_1205,In_14);
or U4762 (N_4762,In_826,In_789);
xor U4763 (N_4763,In_336,In_574);
nand U4764 (N_4764,In_165,In_1231);
and U4765 (N_4765,In_1040,In_420);
and U4766 (N_4766,In_1420,In_819);
and U4767 (N_4767,In_235,In_935);
or U4768 (N_4768,In_234,In_416);
or U4769 (N_4769,In_944,In_1421);
and U4770 (N_4770,In_551,In_521);
nand U4771 (N_4771,In_1130,In_171);
and U4772 (N_4772,In_1172,In_71);
or U4773 (N_4773,In_295,In_1320);
nand U4774 (N_4774,In_347,In_856);
and U4775 (N_4775,In_1327,In_1078);
nand U4776 (N_4776,In_991,In_1094);
nor U4777 (N_4777,In_688,In_110);
xor U4778 (N_4778,In_160,In_120);
nor U4779 (N_4779,In_1390,In_143);
nor U4780 (N_4780,In_871,In_367);
nor U4781 (N_4781,In_1445,In_473);
nor U4782 (N_4782,In_1104,In_356);
xnor U4783 (N_4783,In_815,In_712);
nor U4784 (N_4784,In_1151,In_1250);
and U4785 (N_4785,In_1077,In_544);
nor U4786 (N_4786,In_1180,In_26);
or U4787 (N_4787,In_1399,In_482);
and U4788 (N_4788,In_568,In_1153);
nor U4789 (N_4789,In_908,In_1113);
or U4790 (N_4790,In_1054,In_1276);
xnor U4791 (N_4791,In_374,In_1132);
xnor U4792 (N_4792,In_582,In_648);
nor U4793 (N_4793,In_878,In_106);
and U4794 (N_4794,In_1431,In_181);
nor U4795 (N_4795,In_434,In_1350);
nand U4796 (N_4796,In_813,In_208);
nand U4797 (N_4797,In_914,In_1490);
nor U4798 (N_4798,In_150,In_272);
nand U4799 (N_4799,In_85,In_970);
nor U4800 (N_4800,In_1363,In_523);
nor U4801 (N_4801,In_223,In_853);
nand U4802 (N_4802,In_1497,In_83);
nor U4803 (N_4803,In_1427,In_625);
and U4804 (N_4804,In_499,In_150);
or U4805 (N_4805,In_388,In_1227);
and U4806 (N_4806,In_927,In_72);
or U4807 (N_4807,In_686,In_892);
or U4808 (N_4808,In_1346,In_1331);
nand U4809 (N_4809,In_336,In_243);
xor U4810 (N_4810,In_322,In_1142);
xnor U4811 (N_4811,In_1176,In_1445);
nor U4812 (N_4812,In_513,In_64);
xor U4813 (N_4813,In_1171,In_550);
nor U4814 (N_4814,In_541,In_40);
xor U4815 (N_4815,In_163,In_1323);
or U4816 (N_4816,In_493,In_896);
and U4817 (N_4817,In_1026,In_729);
nand U4818 (N_4818,In_744,In_360);
and U4819 (N_4819,In_988,In_673);
nor U4820 (N_4820,In_1480,In_919);
xnor U4821 (N_4821,In_1342,In_150);
nor U4822 (N_4822,In_258,In_1347);
xor U4823 (N_4823,In_962,In_938);
xor U4824 (N_4824,In_1487,In_497);
and U4825 (N_4825,In_1020,In_827);
nand U4826 (N_4826,In_1218,In_833);
or U4827 (N_4827,In_1047,In_681);
or U4828 (N_4828,In_300,In_1329);
and U4829 (N_4829,In_1038,In_1301);
xor U4830 (N_4830,In_900,In_1229);
nand U4831 (N_4831,In_1384,In_864);
nand U4832 (N_4832,In_1200,In_918);
nand U4833 (N_4833,In_352,In_659);
xnor U4834 (N_4834,In_907,In_1155);
xor U4835 (N_4835,In_199,In_486);
and U4836 (N_4836,In_327,In_873);
and U4837 (N_4837,In_558,In_78);
or U4838 (N_4838,In_762,In_577);
nor U4839 (N_4839,In_324,In_884);
nand U4840 (N_4840,In_669,In_570);
nand U4841 (N_4841,In_306,In_1243);
nor U4842 (N_4842,In_198,In_171);
nand U4843 (N_4843,In_5,In_969);
xor U4844 (N_4844,In_1143,In_557);
or U4845 (N_4845,In_843,In_1221);
and U4846 (N_4846,In_957,In_895);
nor U4847 (N_4847,In_401,In_112);
or U4848 (N_4848,In_631,In_132);
xor U4849 (N_4849,In_492,In_108);
nand U4850 (N_4850,In_1191,In_774);
nor U4851 (N_4851,In_198,In_80);
nor U4852 (N_4852,In_602,In_490);
xnor U4853 (N_4853,In_305,In_1346);
nor U4854 (N_4854,In_1369,In_551);
or U4855 (N_4855,In_280,In_1425);
and U4856 (N_4856,In_917,In_397);
or U4857 (N_4857,In_941,In_649);
or U4858 (N_4858,In_645,In_815);
nand U4859 (N_4859,In_116,In_213);
nor U4860 (N_4860,In_578,In_1071);
and U4861 (N_4861,In_493,In_859);
nor U4862 (N_4862,In_14,In_815);
and U4863 (N_4863,In_876,In_49);
xnor U4864 (N_4864,In_81,In_1308);
xor U4865 (N_4865,In_789,In_931);
xnor U4866 (N_4866,In_1376,In_259);
or U4867 (N_4867,In_413,In_1200);
and U4868 (N_4868,In_840,In_146);
or U4869 (N_4869,In_336,In_1071);
nand U4870 (N_4870,In_594,In_1440);
and U4871 (N_4871,In_425,In_1234);
or U4872 (N_4872,In_1211,In_431);
xor U4873 (N_4873,In_1227,In_1446);
or U4874 (N_4874,In_18,In_794);
xor U4875 (N_4875,In_802,In_1292);
nor U4876 (N_4876,In_737,In_1341);
xnor U4877 (N_4877,In_923,In_951);
xor U4878 (N_4878,In_79,In_307);
and U4879 (N_4879,In_409,In_413);
and U4880 (N_4880,In_365,In_1448);
nor U4881 (N_4881,In_836,In_1119);
xnor U4882 (N_4882,In_1475,In_452);
nand U4883 (N_4883,In_1348,In_541);
or U4884 (N_4884,In_57,In_100);
nand U4885 (N_4885,In_1274,In_256);
nand U4886 (N_4886,In_1049,In_743);
and U4887 (N_4887,In_1406,In_1295);
xor U4888 (N_4888,In_1255,In_1045);
or U4889 (N_4889,In_1345,In_26);
xnor U4890 (N_4890,In_808,In_537);
and U4891 (N_4891,In_743,In_1265);
or U4892 (N_4892,In_1185,In_1172);
nand U4893 (N_4893,In_1368,In_1422);
and U4894 (N_4894,In_1316,In_993);
or U4895 (N_4895,In_1208,In_1046);
or U4896 (N_4896,In_22,In_915);
nor U4897 (N_4897,In_1057,In_967);
xor U4898 (N_4898,In_1253,In_117);
and U4899 (N_4899,In_447,In_374);
xor U4900 (N_4900,In_1207,In_574);
nand U4901 (N_4901,In_419,In_1338);
or U4902 (N_4902,In_1178,In_1101);
nand U4903 (N_4903,In_1181,In_917);
or U4904 (N_4904,In_922,In_720);
and U4905 (N_4905,In_543,In_221);
nand U4906 (N_4906,In_764,In_648);
and U4907 (N_4907,In_652,In_291);
nor U4908 (N_4908,In_672,In_103);
nand U4909 (N_4909,In_780,In_1316);
xor U4910 (N_4910,In_62,In_351);
or U4911 (N_4911,In_10,In_285);
xor U4912 (N_4912,In_1399,In_859);
nand U4913 (N_4913,In_427,In_581);
and U4914 (N_4914,In_214,In_1316);
and U4915 (N_4915,In_403,In_57);
or U4916 (N_4916,In_784,In_1392);
xnor U4917 (N_4917,In_1021,In_655);
and U4918 (N_4918,In_239,In_1405);
and U4919 (N_4919,In_358,In_1182);
or U4920 (N_4920,In_711,In_21);
nand U4921 (N_4921,In_1330,In_1171);
nor U4922 (N_4922,In_1129,In_897);
and U4923 (N_4923,In_1373,In_1405);
or U4924 (N_4924,In_1168,In_292);
xor U4925 (N_4925,In_363,In_848);
xnor U4926 (N_4926,In_349,In_874);
nand U4927 (N_4927,In_1214,In_1159);
and U4928 (N_4928,In_157,In_356);
nor U4929 (N_4929,In_283,In_1155);
and U4930 (N_4930,In_521,In_906);
or U4931 (N_4931,In_1176,In_916);
or U4932 (N_4932,In_40,In_1138);
xor U4933 (N_4933,In_961,In_988);
or U4934 (N_4934,In_1230,In_1481);
nor U4935 (N_4935,In_321,In_216);
and U4936 (N_4936,In_373,In_1317);
or U4937 (N_4937,In_870,In_1311);
nor U4938 (N_4938,In_1020,In_40);
or U4939 (N_4939,In_203,In_446);
xor U4940 (N_4940,In_63,In_227);
and U4941 (N_4941,In_1390,In_1096);
nor U4942 (N_4942,In_1115,In_1300);
and U4943 (N_4943,In_96,In_924);
nor U4944 (N_4944,In_521,In_1034);
or U4945 (N_4945,In_243,In_203);
xor U4946 (N_4946,In_543,In_1469);
and U4947 (N_4947,In_625,In_1380);
and U4948 (N_4948,In_812,In_673);
xnor U4949 (N_4949,In_736,In_1498);
xor U4950 (N_4950,In_255,In_1372);
nor U4951 (N_4951,In_1070,In_1009);
and U4952 (N_4952,In_541,In_206);
and U4953 (N_4953,In_608,In_1348);
and U4954 (N_4954,In_1364,In_1154);
nor U4955 (N_4955,In_1029,In_633);
nand U4956 (N_4956,In_892,In_59);
nor U4957 (N_4957,In_1341,In_887);
nand U4958 (N_4958,In_1048,In_290);
xnor U4959 (N_4959,In_1331,In_345);
nor U4960 (N_4960,In_656,In_883);
and U4961 (N_4961,In_490,In_892);
and U4962 (N_4962,In_1009,In_763);
and U4963 (N_4963,In_600,In_258);
or U4964 (N_4964,In_385,In_1249);
and U4965 (N_4965,In_2,In_445);
or U4966 (N_4966,In_505,In_139);
nand U4967 (N_4967,In_1231,In_190);
xnor U4968 (N_4968,In_346,In_1105);
nor U4969 (N_4969,In_1389,In_285);
and U4970 (N_4970,In_920,In_1379);
or U4971 (N_4971,In_730,In_1299);
and U4972 (N_4972,In_969,In_1463);
or U4973 (N_4973,In_1449,In_1462);
or U4974 (N_4974,In_188,In_533);
xor U4975 (N_4975,In_705,In_306);
and U4976 (N_4976,In_1253,In_1422);
xnor U4977 (N_4977,In_1271,In_477);
or U4978 (N_4978,In_232,In_1103);
or U4979 (N_4979,In_83,In_561);
nand U4980 (N_4980,In_528,In_27);
xnor U4981 (N_4981,In_559,In_709);
and U4982 (N_4982,In_212,In_1446);
xor U4983 (N_4983,In_342,In_1110);
nor U4984 (N_4984,In_878,In_460);
and U4985 (N_4985,In_1330,In_1262);
xnor U4986 (N_4986,In_1083,In_1306);
and U4987 (N_4987,In_474,In_1360);
xnor U4988 (N_4988,In_1000,In_576);
and U4989 (N_4989,In_1015,In_397);
nand U4990 (N_4990,In_553,In_431);
xnor U4991 (N_4991,In_42,In_364);
and U4992 (N_4992,In_419,In_1119);
or U4993 (N_4993,In_747,In_1278);
xnor U4994 (N_4994,In_929,In_717);
nand U4995 (N_4995,In_921,In_575);
nand U4996 (N_4996,In_183,In_354);
nand U4997 (N_4997,In_287,In_10);
and U4998 (N_4998,In_1224,In_128);
and U4999 (N_4999,In_1480,In_834);
and U5000 (N_5000,N_773,N_4515);
xor U5001 (N_5001,N_4590,N_3734);
nor U5002 (N_5002,N_4588,N_3880);
or U5003 (N_5003,N_442,N_3365);
xor U5004 (N_5004,N_4034,N_2525);
or U5005 (N_5005,N_4978,N_1546);
or U5006 (N_5006,N_2392,N_1206);
nor U5007 (N_5007,N_345,N_1766);
xnor U5008 (N_5008,N_3908,N_1405);
xnor U5009 (N_5009,N_241,N_1392);
xnor U5010 (N_5010,N_3104,N_1502);
nor U5011 (N_5011,N_2207,N_1114);
nand U5012 (N_5012,N_4691,N_4662);
xor U5013 (N_5013,N_1493,N_3299);
and U5014 (N_5014,N_313,N_3242);
nand U5015 (N_5015,N_4521,N_2945);
and U5016 (N_5016,N_1371,N_272);
xor U5017 (N_5017,N_1861,N_1927);
and U5018 (N_5018,N_2236,N_1803);
or U5019 (N_5019,N_505,N_3685);
nand U5020 (N_5020,N_1485,N_3395);
nor U5021 (N_5021,N_1393,N_4591);
xnor U5022 (N_5022,N_3222,N_1433);
and U5023 (N_5023,N_2531,N_2056);
or U5024 (N_5024,N_1092,N_1491);
or U5025 (N_5025,N_1951,N_741);
nand U5026 (N_5026,N_4747,N_1020);
or U5027 (N_5027,N_2860,N_2017);
xnor U5028 (N_5028,N_4121,N_3260);
and U5029 (N_5029,N_909,N_3695);
xor U5030 (N_5030,N_3739,N_2808);
and U5031 (N_5031,N_420,N_2031);
or U5032 (N_5032,N_2584,N_3214);
nor U5033 (N_5033,N_114,N_1014);
and U5034 (N_5034,N_1361,N_2633);
nand U5035 (N_5035,N_4518,N_4060);
or U5036 (N_5036,N_4697,N_4058);
nand U5037 (N_5037,N_1057,N_447);
nand U5038 (N_5038,N_4057,N_2163);
nor U5039 (N_5039,N_2904,N_4346);
nand U5040 (N_5040,N_191,N_1532);
nor U5041 (N_5041,N_3752,N_2907);
xor U5042 (N_5042,N_1196,N_3029);
nor U5043 (N_5043,N_854,N_3736);
nor U5044 (N_5044,N_223,N_729);
xor U5045 (N_5045,N_101,N_474);
nor U5046 (N_5046,N_4274,N_2006);
xor U5047 (N_5047,N_1709,N_4499);
and U5048 (N_5048,N_4157,N_1427);
nor U5049 (N_5049,N_1655,N_1016);
or U5050 (N_5050,N_3667,N_283);
and U5051 (N_5051,N_1091,N_1323);
or U5052 (N_5052,N_4433,N_4541);
or U5053 (N_5053,N_163,N_328);
and U5054 (N_5054,N_2179,N_2129);
nand U5055 (N_5055,N_2449,N_944);
or U5056 (N_5056,N_831,N_4266);
nand U5057 (N_5057,N_2204,N_4907);
nor U5058 (N_5058,N_4733,N_641);
and U5059 (N_5059,N_4509,N_4218);
nand U5060 (N_5060,N_870,N_4592);
nand U5061 (N_5061,N_2354,N_4349);
xor U5062 (N_5062,N_4307,N_3781);
or U5063 (N_5063,N_2950,N_993);
or U5064 (N_5064,N_3162,N_4746);
or U5065 (N_5065,N_4155,N_1854);
and U5066 (N_5066,N_3692,N_3709);
xor U5067 (N_5067,N_4717,N_2721);
xnor U5068 (N_5068,N_295,N_3426);
xor U5069 (N_5069,N_1037,N_2308);
and U5070 (N_5070,N_2772,N_4508);
xnor U5071 (N_5071,N_4839,N_23);
or U5072 (N_5072,N_2867,N_406);
nor U5073 (N_5073,N_4769,N_1339);
nor U5074 (N_5074,N_2057,N_3553);
xor U5075 (N_5075,N_2238,N_3530);
xnor U5076 (N_5076,N_1116,N_4589);
or U5077 (N_5077,N_1970,N_3241);
nand U5078 (N_5078,N_3337,N_1475);
or U5079 (N_5079,N_4069,N_1700);
and U5080 (N_5080,N_168,N_337);
or U5081 (N_5081,N_457,N_2981);
nand U5082 (N_5082,N_2460,N_4781);
or U5083 (N_5083,N_2258,N_3179);
xor U5084 (N_5084,N_1516,N_1638);
xnor U5085 (N_5085,N_3506,N_4262);
nor U5086 (N_5086,N_2751,N_2281);
nor U5087 (N_5087,N_1722,N_467);
or U5088 (N_5088,N_4072,N_2288);
and U5089 (N_5089,N_3678,N_737);
xor U5090 (N_5090,N_4438,N_2612);
or U5091 (N_5091,N_2949,N_4260);
and U5092 (N_5092,N_2796,N_3262);
nand U5093 (N_5093,N_2989,N_419);
nor U5094 (N_5094,N_1859,N_2505);
xnor U5095 (N_5095,N_4621,N_318);
and U5096 (N_5096,N_2254,N_3433);
nand U5097 (N_5097,N_49,N_2091);
or U5098 (N_5098,N_3082,N_3634);
and U5099 (N_5099,N_4551,N_2978);
or U5100 (N_5100,N_2788,N_1935);
or U5101 (N_5101,N_4224,N_1451);
nor U5102 (N_5102,N_973,N_4986);
or U5103 (N_5103,N_2383,N_2208);
and U5104 (N_5104,N_4889,N_4390);
nand U5105 (N_5105,N_1587,N_455);
xnor U5106 (N_5106,N_3289,N_3891);
or U5107 (N_5107,N_3170,N_386);
nand U5108 (N_5108,N_4884,N_1787);
or U5109 (N_5109,N_1496,N_3534);
and U5110 (N_5110,N_2757,N_463);
xnor U5111 (N_5111,N_4685,N_952);
and U5112 (N_5112,N_824,N_255);
nor U5113 (N_5113,N_3507,N_2622);
xnor U5114 (N_5114,N_4998,N_2188);
nor U5115 (N_5115,N_4983,N_1942);
nor U5116 (N_5116,N_2866,N_4392);
and U5117 (N_5117,N_2851,N_704);
xor U5118 (N_5118,N_2465,N_826);
xnor U5119 (N_5119,N_1737,N_3776);
nand U5120 (N_5120,N_1173,N_820);
or U5121 (N_5121,N_2873,N_1620);
nor U5122 (N_5122,N_4113,N_1593);
xnor U5123 (N_5123,N_494,N_3556);
nand U5124 (N_5124,N_960,N_3652);
nor U5125 (N_5125,N_2371,N_3959);
and U5126 (N_5126,N_2070,N_2361);
nor U5127 (N_5127,N_362,N_2976);
nand U5128 (N_5128,N_2260,N_2852);
or U5129 (N_5129,N_1424,N_3157);
nand U5130 (N_5130,N_3915,N_4004);
or U5131 (N_5131,N_12,N_1224);
xor U5132 (N_5132,N_2464,N_1997);
nand U5133 (N_5133,N_4759,N_2169);
or U5134 (N_5134,N_2799,N_1431);
or U5135 (N_5135,N_2014,N_1675);
xor U5136 (N_5136,N_2473,N_4073);
and U5137 (N_5137,N_2559,N_2754);
xor U5138 (N_5138,N_2709,N_649);
and U5139 (N_5139,N_3073,N_4795);
nand U5140 (N_5140,N_2128,N_4596);
or U5141 (N_5141,N_2364,N_1623);
or U5142 (N_5142,N_4263,N_3503);
or U5143 (N_5143,N_3822,N_2651);
and U5144 (N_5144,N_3898,N_3620);
xnor U5145 (N_5145,N_2266,N_1536);
nand U5146 (N_5146,N_2979,N_2840);
nand U5147 (N_5147,N_268,N_2146);
nand U5148 (N_5148,N_1876,N_2043);
nor U5149 (N_5149,N_1106,N_4139);
and U5150 (N_5150,N_2016,N_4114);
and U5151 (N_5151,N_1466,N_3995);
xnor U5152 (N_5152,N_1313,N_4253);
or U5153 (N_5153,N_2075,N_4820);
nor U5154 (N_5154,N_290,N_3630);
nor U5155 (N_5155,N_2412,N_4186);
or U5156 (N_5156,N_4085,N_4446);
nor U5157 (N_5157,N_771,N_3571);
or U5158 (N_5158,N_4873,N_1017);
nand U5159 (N_5159,N_4491,N_4627);
nand U5160 (N_5160,N_1525,N_666);
xnor U5161 (N_5161,N_3255,N_3129);
and U5162 (N_5162,N_2180,N_4129);
or U5163 (N_5163,N_3797,N_1239);
or U5164 (N_5164,N_4549,N_2565);
nand U5165 (N_5165,N_4776,N_4294);
nor U5166 (N_5166,N_1778,N_2804);
xor U5167 (N_5167,N_4394,N_3462);
or U5168 (N_5168,N_3862,N_3669);
nand U5169 (N_5169,N_4844,N_2269);
xor U5170 (N_5170,N_558,N_3471);
xnor U5171 (N_5171,N_2320,N_3075);
and U5172 (N_5172,N_2630,N_84);
or U5173 (N_5173,N_2246,N_5);
or U5174 (N_5174,N_1812,N_2481);
and U5175 (N_5175,N_3294,N_2454);
nand U5176 (N_5176,N_2629,N_786);
nand U5177 (N_5177,N_722,N_4232);
nand U5178 (N_5178,N_1893,N_4900);
nand U5179 (N_5179,N_2106,N_1726);
and U5180 (N_5180,N_1899,N_144);
nor U5181 (N_5181,N_3084,N_1376);
and U5182 (N_5182,N_2265,N_1053);
nand U5183 (N_5183,N_2870,N_2899);
nor U5184 (N_5184,N_2319,N_1968);
or U5185 (N_5185,N_2199,N_932);
or U5186 (N_5186,N_4205,N_1343);
and U5187 (N_5187,N_4337,N_3671);
xor U5188 (N_5188,N_2488,N_3682);
or U5189 (N_5189,N_1497,N_2432);
and U5190 (N_5190,N_4951,N_143);
nor U5191 (N_5191,N_2170,N_1896);
nor U5192 (N_5192,N_1465,N_3836);
xor U5193 (N_5193,N_425,N_2386);
nand U5194 (N_5194,N_1608,N_3410);
nand U5195 (N_5195,N_2385,N_343);
xor U5196 (N_5196,N_39,N_2774);
xnor U5197 (N_5197,N_1971,N_1048);
nand U5198 (N_5198,N_3713,N_2399);
and U5199 (N_5199,N_4152,N_2741);
nand U5200 (N_5200,N_3960,N_465);
nor U5201 (N_5201,N_545,N_2752);
xnor U5202 (N_5202,N_2409,N_4361);
xor U5203 (N_5203,N_2289,N_2092);
nor U5204 (N_5204,N_3013,N_4929);
and U5205 (N_5205,N_231,N_2303);
nor U5206 (N_5206,N_4049,N_1674);
xnor U5207 (N_5207,N_11,N_2506);
or U5208 (N_5208,N_4582,N_4030);
xor U5209 (N_5209,N_2839,N_1295);
nor U5210 (N_5210,N_2099,N_3352);
nand U5211 (N_5211,N_617,N_1093);
nor U5212 (N_5212,N_3581,N_2939);
xor U5213 (N_5213,N_154,N_4966);
or U5214 (N_5214,N_4031,N_1571);
xor U5215 (N_5215,N_2275,N_506);
and U5216 (N_5216,N_2843,N_2942);
and U5217 (N_5217,N_1097,N_2060);
nor U5218 (N_5218,N_1658,N_1187);
nand U5219 (N_5219,N_939,N_2183);
or U5220 (N_5220,N_1462,N_1013);
and U5221 (N_5221,N_1203,N_3541);
or U5222 (N_5222,N_3422,N_3258);
xor U5223 (N_5223,N_730,N_3805);
and U5224 (N_5224,N_3917,N_1910);
nand U5225 (N_5225,N_1642,N_2102);
nand U5226 (N_5226,N_1622,N_2532);
nand U5227 (N_5227,N_172,N_596);
xnor U5228 (N_5228,N_1260,N_203);
or U5229 (N_5229,N_4869,N_4735);
or U5230 (N_5230,N_2470,N_597);
xnor U5231 (N_5231,N_949,N_4243);
and U5232 (N_5232,N_2592,N_1380);
nand U5233 (N_5233,N_3557,N_4829);
or U5234 (N_5234,N_685,N_2143);
xor U5235 (N_5235,N_1128,N_1998);
nor U5236 (N_5236,N_3193,N_1448);
and U5237 (N_5237,N_1567,N_1625);
xor U5238 (N_5238,N_2457,N_3924);
and U5239 (N_5239,N_4938,N_2677);
nor U5240 (N_5240,N_4504,N_1241);
and U5241 (N_5241,N_3527,N_4649);
xnor U5242 (N_5242,N_3487,N_1936);
and U5243 (N_5243,N_91,N_4953);
and U5244 (N_5244,N_211,N_2570);
nand U5245 (N_5245,N_3957,N_1221);
nor U5246 (N_5246,N_4854,N_3024);
xor U5247 (N_5247,N_2517,N_4311);
nand U5248 (N_5248,N_401,N_2039);
or U5249 (N_5249,N_2007,N_276);
nand U5250 (N_5250,N_443,N_1247);
and U5251 (N_5251,N_4424,N_716);
and U5252 (N_5252,N_3755,N_3972);
and U5253 (N_5253,N_1394,N_3857);
and U5254 (N_5254,N_3148,N_2462);
nor U5255 (N_5255,N_1989,N_2737);
and U5256 (N_5256,N_3470,N_621);
xnor U5257 (N_5257,N_3818,N_4342);
xor U5258 (N_5258,N_4377,N_1118);
and U5259 (N_5259,N_2656,N_3386);
nor U5260 (N_5260,N_4089,N_4503);
or U5261 (N_5261,N_3187,N_4773);
nor U5262 (N_5262,N_553,N_2356);
and U5263 (N_5263,N_1333,N_3374);
nand U5264 (N_5264,N_1663,N_2909);
and U5265 (N_5265,N_2218,N_2975);
or U5266 (N_5266,N_4163,N_1719);
or U5267 (N_5267,N_1902,N_1165);
nor U5268 (N_5268,N_431,N_721);
or U5269 (N_5269,N_1850,N_4895);
nand U5270 (N_5270,N_1975,N_3207);
nor U5271 (N_5271,N_429,N_2539);
nor U5272 (N_5272,N_2398,N_703);
or U5273 (N_5273,N_1569,N_2337);
or U5274 (N_5274,N_1024,N_1157);
and U5275 (N_5275,N_1319,N_81);
and U5276 (N_5276,N_4798,N_1820);
nor U5277 (N_5277,N_68,N_4940);
xor U5278 (N_5278,N_1487,N_978);
nor U5279 (N_5279,N_857,N_3770);
xnor U5280 (N_5280,N_3688,N_4899);
xnor U5281 (N_5281,N_2453,N_3497);
xnor U5282 (N_5282,N_1327,N_2413);
nor U5283 (N_5283,N_2263,N_540);
nand U5284 (N_5284,N_265,N_2684);
xnor U5285 (N_5285,N_4570,N_2815);
or U5286 (N_5286,N_70,N_2881);
nor U5287 (N_5287,N_2639,N_2631);
nor U5288 (N_5288,N_53,N_4604);
nor U5289 (N_5289,N_2307,N_3074);
and U5290 (N_5290,N_4693,N_2913);
and U5291 (N_5291,N_3225,N_1320);
nand U5292 (N_5292,N_2704,N_1796);
or U5293 (N_5293,N_3684,N_4749);
and U5294 (N_5294,N_492,N_2540);
and U5295 (N_5295,N_2609,N_4875);
or U5296 (N_5296,N_118,N_747);
xor U5297 (N_5297,N_1214,N_1129);
or U5298 (N_5298,N_2159,N_1692);
and U5299 (N_5299,N_1768,N_3201);
or U5300 (N_5300,N_853,N_4456);
and U5301 (N_5301,N_3650,N_1089);
nand U5302 (N_5302,N_4314,N_934);
nand U5303 (N_5303,N_3830,N_2348);
nor U5304 (N_5304,N_3033,N_3708);
nor U5305 (N_5305,N_4335,N_2195);
nor U5306 (N_5306,N_513,N_3921);
or U5307 (N_5307,N_622,N_3820);
and U5308 (N_5308,N_3551,N_1305);
and U5309 (N_5309,N_387,N_2551);
or U5310 (N_5310,N_1712,N_1202);
xor U5311 (N_5311,N_1384,N_3637);
and U5312 (N_5312,N_1182,N_3293);
xnor U5313 (N_5313,N_3078,N_1857);
xor U5314 (N_5314,N_4906,N_1685);
and U5315 (N_5315,N_294,N_3764);
xor U5316 (N_5316,N_3699,N_720);
nand U5317 (N_5317,N_4511,N_862);
or U5318 (N_5318,N_1261,N_2894);
nand U5319 (N_5319,N_2345,N_1784);
or U5320 (N_5320,N_2703,N_4422);
nor U5321 (N_5321,N_2344,N_4930);
nand U5322 (N_5322,N_1590,N_3922);
nand U5323 (N_5323,N_3228,N_798);
xnor U5324 (N_5324,N_2330,N_4320);
nor U5325 (N_5325,N_483,N_1527);
and U5326 (N_5326,N_4531,N_2952);
nor U5327 (N_5327,N_1518,N_4387);
nand U5328 (N_5328,N_2668,N_2632);
nor U5329 (N_5329,N_2053,N_503);
nor U5330 (N_5330,N_2705,N_3850);
nand U5331 (N_5331,N_1417,N_335);
xor U5332 (N_5332,N_4370,N_607);
nand U5333 (N_5333,N_1031,N_466);
xor U5334 (N_5334,N_3611,N_692);
or U5335 (N_5335,N_3377,N_1336);
and U5336 (N_5336,N_2244,N_4528);
nor U5337 (N_5337,N_3500,N_3756);
or U5338 (N_5338,N_2917,N_3322);
or U5339 (N_5339,N_998,N_1085);
xor U5340 (N_5340,N_1793,N_4386);
xor U5341 (N_5341,N_3750,N_1707);
nand U5342 (N_5342,N_670,N_2022);
and U5343 (N_5343,N_3769,N_1956);
or U5344 (N_5344,N_3184,N_3054);
xor U5345 (N_5345,N_4671,N_4497);
nand U5346 (N_5346,N_719,N_1508);
or U5347 (N_5347,N_3544,N_2301);
xor U5348 (N_5348,N_4360,N_3070);
xor U5349 (N_5349,N_4296,N_970);
or U5350 (N_5350,N_1826,N_3409);
nor U5351 (N_5351,N_60,N_3169);
and U5352 (N_5352,N_602,N_4395);
nor U5353 (N_5353,N_2058,N_3430);
nor U5354 (N_5354,N_239,N_4577);
xnor U5355 (N_5355,N_2864,N_4571);
nor U5356 (N_5356,N_1180,N_1283);
and U5357 (N_5357,N_4874,N_3119);
xor U5358 (N_5358,N_4202,N_2436);
nor U5359 (N_5359,N_637,N_2463);
nor U5360 (N_5360,N_1457,N_2906);
nor U5361 (N_5361,N_2770,N_41);
xnor U5362 (N_5362,N_985,N_1695);
and U5363 (N_5363,N_863,N_3702);
xnor U5364 (N_5364,N_1222,N_2189);
or U5365 (N_5365,N_1410,N_2977);
or U5366 (N_5366,N_1352,N_1363);
nor U5367 (N_5367,N_825,N_1795);
nor U5368 (N_5368,N_4306,N_2544);
xnor U5369 (N_5369,N_3899,N_3389);
xnor U5370 (N_5370,N_1422,N_4505);
or U5371 (N_5371,N_3363,N_384);
nand U5372 (N_5372,N_2523,N_103);
and U5373 (N_5373,N_1467,N_181);
xor U5374 (N_5374,N_1842,N_3944);
or U5375 (N_5375,N_2599,N_1752);
nor U5376 (N_5376,N_2963,N_4280);
nand U5377 (N_5377,N_4475,N_2600);
and U5378 (N_5378,N_3384,N_2489);
nand U5379 (N_5379,N_2594,N_4179);
nand U5380 (N_5380,N_4648,N_4097);
xnor U5381 (N_5381,N_1120,N_4134);
or U5382 (N_5382,N_4706,N_4680);
and U5383 (N_5383,N_1537,N_2495);
or U5384 (N_5384,N_2181,N_125);
or U5385 (N_5385,N_1055,N_4107);
nor U5386 (N_5386,N_2325,N_864);
nor U5387 (N_5387,N_2965,N_4087);
nand U5388 (N_5388,N_2928,N_4240);
or U5389 (N_5389,N_1140,N_1176);
nand U5390 (N_5390,N_808,N_681);
nand U5391 (N_5391,N_2996,N_4552);
or U5392 (N_5392,N_941,N_1958);
xnor U5393 (N_5393,N_3077,N_686);
nor U5394 (N_5394,N_2617,N_52);
and U5395 (N_5395,N_4227,N_3385);
nor U5396 (N_5396,N_1296,N_3606);
and U5397 (N_5397,N_4653,N_1220);
nand U5398 (N_5398,N_3128,N_2501);
xnor U5399 (N_5399,N_4011,N_2615);
and U5400 (N_5400,N_2003,N_3189);
or U5401 (N_5401,N_3266,N_2097);
nor U5402 (N_5402,N_3566,N_408);
or U5403 (N_5403,N_569,N_3286);
xnor U5404 (N_5404,N_848,N_3309);
nor U5405 (N_5405,N_611,N_4495);
xnor U5406 (N_5406,N_2417,N_1356);
xor U5407 (N_5407,N_1773,N_3985);
or U5408 (N_5408,N_2688,N_246);
xnor U5409 (N_5409,N_4259,N_662);
or U5410 (N_5410,N_4924,N_4090);
and U5411 (N_5411,N_148,N_1340);
xor U5412 (N_5412,N_2837,N_3563);
or U5413 (N_5413,N_4678,N_1289);
nor U5414 (N_5414,N_4092,N_4813);
nand U5415 (N_5415,N_1235,N_2915);
nand U5416 (N_5416,N_4881,N_4014);
and U5417 (N_5417,N_634,N_3053);
nor U5418 (N_5418,N_4506,N_965);
nor U5419 (N_5419,N_1799,N_1946);
or U5420 (N_5420,N_2296,N_4677);
xnor U5421 (N_5421,N_1095,N_3740);
nand U5422 (N_5422,N_1932,N_4804);
or U5423 (N_5423,N_456,N_1823);
nand U5424 (N_5424,N_461,N_2502);
nand U5425 (N_5425,N_264,N_3413);
and U5426 (N_5426,N_1904,N_1542);
nor U5427 (N_5427,N_300,N_3350);
nor U5428 (N_5428,N_3067,N_4643);
nor U5429 (N_5429,N_3601,N_2595);
nor U5430 (N_5430,N_1151,N_1684);
and U5431 (N_5431,N_1711,N_4228);
xnor U5432 (N_5432,N_4026,N_3876);
xnor U5433 (N_5433,N_3555,N_2747);
xnor U5434 (N_5434,N_4752,N_2997);
nand U5435 (N_5435,N_4192,N_2024);
nor U5436 (N_5436,N_3195,N_1225);
nand U5437 (N_5437,N_3841,N_4242);
and U5438 (N_5438,N_3227,N_4231);
and U5439 (N_5439,N_4450,N_2883);
and U5440 (N_5440,N_3447,N_1258);
nor U5441 (N_5441,N_437,N_59);
xnor U5442 (N_5442,N_2155,N_1103);
nor U5443 (N_5443,N_888,N_3855);
xor U5444 (N_5444,N_2980,N_3757);
or U5445 (N_5445,N_1147,N_868);
xnor U5446 (N_5446,N_2521,N_4147);
nor U5447 (N_5447,N_171,N_3003);
xor U5448 (N_5448,N_4931,N_2037);
xor U5449 (N_5449,N_1738,N_1341);
nor U5450 (N_5450,N_2192,N_4911);
and U5451 (N_5451,N_3432,N_2827);
xnor U5452 (N_5452,N_3287,N_1355);
nor U5453 (N_5453,N_412,N_296);
nand U5454 (N_5454,N_3993,N_975);
or U5455 (N_5455,N_2641,N_3221);
nor U5456 (N_5456,N_3656,N_533);
nor U5457 (N_5457,N_4914,N_2069);
nor U5458 (N_5458,N_1284,N_4756);
nand U5459 (N_5459,N_3645,N_1104);
and U5460 (N_5460,N_100,N_2209);
or U5461 (N_5461,N_3044,N_2117);
nor U5462 (N_5462,N_917,N_4252);
xor U5463 (N_5463,N_3872,N_1605);
and U5464 (N_5464,N_1137,N_4046);
xor U5465 (N_5465,N_940,N_115);
and U5466 (N_5466,N_3835,N_3659);
nand U5467 (N_5467,N_3916,N_1928);
xor U5468 (N_5468,N_4183,N_4020);
xnor U5469 (N_5469,N_4527,N_3176);
xor U5470 (N_5470,N_2920,N_738);
or U5471 (N_5471,N_247,N_4690);
and U5472 (N_5472,N_3509,N_2874);
xor U5473 (N_5473,N_2471,N_1094);
or U5474 (N_5474,N_4879,N_1135);
or U5475 (N_5475,N_615,N_1621);
nand U5476 (N_5476,N_1314,N_4894);
and U5477 (N_5477,N_4326,N_581);
and U5478 (N_5478,N_4832,N_3929);
and U5479 (N_5479,N_3800,N_2174);
and U5480 (N_5480,N_3134,N_2131);
and U5481 (N_5481,N_1918,N_4791);
and U5482 (N_5482,N_2828,N_3940);
or U5483 (N_5483,N_3083,N_224);
and U5484 (N_5484,N_3153,N_2974);
nor U5485 (N_5485,N_1603,N_4904);
xor U5486 (N_5486,N_3590,N_2514);
nor U5487 (N_5487,N_896,N_4158);
and U5488 (N_5488,N_469,N_2055);
or U5489 (N_5489,N_4412,N_3198);
and U5490 (N_5490,N_1853,N_3878);
or U5491 (N_5491,N_4463,N_4077);
or U5492 (N_5492,N_3051,N_2558);
nand U5493 (N_5493,N_3837,N_2530);
or U5494 (N_5494,N_995,N_1572);
nand U5495 (N_5495,N_3575,N_309);
nand U5496 (N_5496,N_2256,N_2264);
and U5497 (N_5497,N_3388,N_2930);
or U5498 (N_5498,N_3853,N_4994);
or U5499 (N_5499,N_3937,N_2746);
nor U5500 (N_5500,N_1022,N_1161);
or U5501 (N_5501,N_3100,N_3285);
nor U5502 (N_5502,N_3809,N_3329);
xor U5503 (N_5503,N_2691,N_4172);
nor U5504 (N_5504,N_537,N_350);
or U5505 (N_5505,N_3884,N_1630);
nor U5506 (N_5506,N_3099,N_2846);
and U5507 (N_5507,N_3926,N_1036);
nand U5508 (N_5508,N_2378,N_1446);
nor U5509 (N_5509,N_1306,N_4247);
nor U5510 (N_5510,N_2001,N_1105);
and U5511 (N_5511,N_77,N_2929);
and U5512 (N_5512,N_4404,N_813);
and U5513 (N_5513,N_3478,N_1513);
nand U5514 (N_5514,N_4646,N_156);
and U5515 (N_5515,N_3691,N_379);
or U5516 (N_5516,N_4033,N_1840);
nor U5517 (N_5517,N_2717,N_2601);
and U5518 (N_5518,N_1442,N_2393);
nor U5519 (N_5519,N_1389,N_1856);
and U5520 (N_5520,N_3209,N_1588);
and U5521 (N_5521,N_745,N_4165);
nor U5522 (N_5522,N_3554,N_1406);
or U5523 (N_5523,N_415,N_4580);
nand U5524 (N_5524,N_1559,N_1750);
xor U5525 (N_5525,N_1748,N_664);
or U5526 (N_5526,N_3407,N_2822);
or U5527 (N_5527,N_2661,N_2635);
or U5528 (N_5528,N_88,N_1043);
nand U5529 (N_5529,N_232,N_1521);
nor U5530 (N_5530,N_3545,N_1038);
nor U5531 (N_5531,N_2957,N_986);
nor U5532 (N_5532,N_4803,N_2561);
nand U5533 (N_5533,N_1992,N_1201);
or U5534 (N_5534,N_332,N_1961);
and U5535 (N_5535,N_942,N_1566);
xor U5536 (N_5536,N_3455,N_1648);
or U5537 (N_5537,N_1251,N_1889);
xnor U5538 (N_5538,N_1025,N_3588);
nand U5539 (N_5539,N_4762,N_3737);
nor U5540 (N_5540,N_1782,N_4822);
nor U5541 (N_5541,N_3782,N_2035);
nand U5542 (N_5542,N_2171,N_319);
xor U5543 (N_5543,N_373,N_839);
nand U5544 (N_5544,N_3047,N_4826);
nand U5545 (N_5545,N_3967,N_3975);
nor U5546 (N_5546,N_2416,N_4237);
nand U5547 (N_5547,N_4234,N_508);
nand U5548 (N_5548,N_2587,N_400);
xnor U5549 (N_5549,N_856,N_1308);
nor U5550 (N_5550,N_2111,N_969);
or U5551 (N_5551,N_2239,N_1875);
nor U5552 (N_5552,N_2956,N_4027);
nor U5553 (N_5553,N_320,N_531);
nand U5554 (N_5554,N_683,N_3631);
xor U5555 (N_5555,N_4044,N_900);
or U5556 (N_5556,N_82,N_1456);
xnor U5557 (N_5557,N_619,N_3310);
or U5558 (N_5558,N_2311,N_3370);
xor U5559 (N_5559,N_3406,N_2797);
and U5560 (N_5560,N_4694,N_273);
nand U5561 (N_5561,N_4189,N_3155);
and U5562 (N_5562,N_2573,N_916);
or U5563 (N_5563,N_1628,N_317);
nand U5564 (N_5564,N_4981,N_4045);
nor U5565 (N_5565,N_3306,N_613);
nand U5566 (N_5566,N_4660,N_1280);
and U5567 (N_5567,N_2847,N_2419);
and U5568 (N_5568,N_1056,N_1078);
xor U5569 (N_5569,N_2968,N_1535);
xnor U5570 (N_5570,N_4842,N_4703);
and U5571 (N_5571,N_3112,N_3292);
and U5572 (N_5572,N_1860,N_2178);
nand U5573 (N_5573,N_3854,N_4315);
nor U5574 (N_5574,N_385,N_2962);
nor U5575 (N_5575,N_1877,N_3428);
nor U5576 (N_5576,N_2468,N_1195);
and U5577 (N_5577,N_4193,N_673);
and U5578 (N_5578,N_3834,N_4489);
xor U5579 (N_5579,N_4457,N_270);
xor U5580 (N_5580,N_775,N_4631);
nor U5581 (N_5581,N_640,N_4796);
or U5582 (N_5582,N_475,N_1109);
or U5583 (N_5583,N_3391,N_1599);
and U5584 (N_5584,N_2076,N_959);
and U5585 (N_5585,N_582,N_659);
and U5586 (N_5586,N_1519,N_4927);
nor U5587 (N_5587,N_983,N_4254);
or U5588 (N_5588,N_4572,N_3906);
nand U5589 (N_5589,N_142,N_3234);
or U5590 (N_5590,N_4743,N_2475);
and U5591 (N_5591,N_3485,N_1966);
or U5592 (N_5592,N_3766,N_979);
nand U5593 (N_5593,N_4775,N_257);
nor U5594 (N_5594,N_912,N_4988);
xnor U5595 (N_5595,N_3543,N_421);
nor U5596 (N_5596,N_2537,N_4695);
nor U5597 (N_5597,N_1849,N_4088);
or U5598 (N_5598,N_4824,N_3986);
xnor U5599 (N_5599,N_4100,N_3552);
and U5600 (N_5600,N_1647,N_4613);
nand U5601 (N_5601,N_1064,N_1334);
xor U5602 (N_5602,N_2044,N_3461);
nand U5603 (N_5603,N_2011,N_1745);
and U5604 (N_5604,N_3319,N_968);
or U5605 (N_5605,N_4091,N_2535);
xnor U5606 (N_5606,N_4115,N_526);
nor U5607 (N_5607,N_4665,N_1598);
or U5608 (N_5608,N_1351,N_706);
nand U5609 (N_5609,N_610,N_4777);
and U5610 (N_5610,N_3648,N_1476);
or U5611 (N_5611,N_3866,N_3795);
or U5612 (N_5612,N_2309,N_1679);
xnor U5613 (N_5613,N_4184,N_4840);
nor U5614 (N_5614,N_4663,N_4148);
or U5615 (N_5615,N_3743,N_2328);
and U5616 (N_5616,N_3403,N_381);
or U5617 (N_5617,N_2318,N_1939);
or U5618 (N_5618,N_549,N_1948);
and U5619 (N_5619,N_1175,N_2046);
nor U5620 (N_5620,N_3583,N_2153);
nand U5621 (N_5621,N_3651,N_3280);
xnor U5622 (N_5622,N_3676,N_847);
and U5623 (N_5623,N_4037,N_557);
nor U5624 (N_5624,N_1098,N_2036);
or U5625 (N_5625,N_1126,N_889);
xor U5626 (N_5626,N_3232,N_4566);
or U5627 (N_5627,N_4225,N_4304);
nor U5628 (N_5628,N_4836,N_1528);
nand U5629 (N_5629,N_3118,N_614);
or U5630 (N_5630,N_2569,N_3504);
nor U5631 (N_5631,N_930,N_26);
xor U5632 (N_5632,N_1088,N_3206);
nand U5633 (N_5633,N_3658,N_1869);
nor U5634 (N_5634,N_4530,N_2210);
and U5635 (N_5635,N_1558,N_4785);
and U5636 (N_5636,N_2992,N_2807);
nand U5637 (N_5637,N_869,N_2424);
and U5638 (N_5638,N_2581,N_2112);
nor U5639 (N_5639,N_3536,N_4432);
and U5640 (N_5640,N_4636,N_799);
or U5641 (N_5641,N_3812,N_2248);
and U5642 (N_5642,N_2425,N_1253);
nor U5643 (N_5643,N_346,N_2643);
nor U5644 (N_5644,N_1643,N_50);
xor U5645 (N_5645,N_1204,N_4093);
nand U5646 (N_5646,N_4713,N_4249);
xnor U5647 (N_5647,N_2756,N_3673);
xnor U5648 (N_5648,N_538,N_4851);
nand U5649 (N_5649,N_3852,N_991);
and U5650 (N_5650,N_2052,N_3333);
or U5651 (N_5651,N_2034,N_4893);
or U5652 (N_5652,N_4086,N_3452);
nand U5653 (N_5653,N_1194,N_3172);
nand U5654 (N_5654,N_4626,N_744);
or U5655 (N_5655,N_2234,N_2574);
nand U5656 (N_5656,N_378,N_2026);
or U5657 (N_5657,N_4153,N_424);
nor U5658 (N_5658,N_4137,N_2138);
and U5659 (N_5659,N_2513,N_780);
or U5660 (N_5660,N_511,N_4976);
nor U5661 (N_5661,N_770,N_3080);
nor U5662 (N_5662,N_121,N_267);
or U5663 (N_5663,N_1995,N_1514);
nand U5664 (N_5664,N_3277,N_205);
nand U5665 (N_5665,N_2472,N_3415);
nor U5666 (N_5666,N_3466,N_1291);
nand U5667 (N_5667,N_3712,N_4279);
and U5668 (N_5668,N_186,N_321);
xnor U5669 (N_5669,N_2964,N_4714);
nor U5670 (N_5670,N_4615,N_4557);
nand U5671 (N_5671,N_2205,N_3612);
or U5672 (N_5672,N_4792,N_1892);
nor U5673 (N_5673,N_3968,N_3472);
xor U5674 (N_5674,N_2761,N_543);
nor U5675 (N_5675,N_2445,N_2167);
xnor U5676 (N_5676,N_519,N_2079);
nand U5677 (N_5677,N_4602,N_1852);
xor U5678 (N_5678,N_436,N_349);
nor U5679 (N_5679,N_2338,N_2486);
and U5680 (N_5680,N_2892,N_1724);
nand U5681 (N_5681,N_837,N_120);
xnor U5682 (N_5682,N_3726,N_2912);
nand U5683 (N_5683,N_3146,N_4688);
xnor U5684 (N_5684,N_4363,N_1326);
nor U5685 (N_5685,N_3842,N_189);
xor U5686 (N_5686,N_222,N_796);
or U5687 (N_5687,N_3817,N_1287);
or U5688 (N_5688,N_2611,N_1271);
nand U5689 (N_5689,N_4841,N_1759);
nor U5690 (N_5690,N_2363,N_3768);
and U5691 (N_5691,N_4782,N_4816);
nor U5692 (N_5692,N_266,N_252);
nand U5693 (N_5693,N_3412,N_2474);
nor U5694 (N_5694,N_3015,N_881);
nand U5695 (N_5695,N_2759,N_1792);
xnor U5696 (N_5696,N_2498,N_3271);
and U5697 (N_5697,N_4837,N_491);
and U5698 (N_5698,N_606,N_1595);
or U5699 (N_5699,N_752,N_899);
or U5700 (N_5700,N_3989,N_4686);
and U5701 (N_5701,N_962,N_1469);
and U5702 (N_5702,N_1288,N_4264);
and U5703 (N_5703,N_2546,N_2734);
nand U5704 (N_5704,N_3701,N_1981);
nand U5705 (N_5705,N_3196,N_1473);
nand U5706 (N_5706,N_2579,N_2972);
and U5707 (N_5707,N_4972,N_4126);
or U5708 (N_5708,N_230,N_4715);
or U5709 (N_5709,N_4909,N_325);
nor U5710 (N_5710,N_1479,N_3952);
nor U5711 (N_5711,N_1583,N_2479);
or U5712 (N_5712,N_4975,N_2083);
nand U5713 (N_5713,N_3923,N_1574);
xnor U5714 (N_5714,N_175,N_445);
or U5715 (N_5715,N_3900,N_3072);
and U5716 (N_5716,N_1509,N_2598);
nor U5717 (N_5717,N_1430,N_1425);
nor U5718 (N_5718,N_1023,N_1967);
xor U5719 (N_5719,N_2790,N_2027);
xor U5720 (N_5720,N_1353,N_2944);
xnor U5721 (N_5721,N_1191,N_1207);
or U5722 (N_5722,N_4788,N_3300);
nand U5723 (N_5723,N_79,N_80);
nand U5724 (N_5724,N_4807,N_976);
nand U5725 (N_5725,N_354,N_3249);
xnor U5726 (N_5726,N_2560,N_4272);
xor U5727 (N_5727,N_4818,N_2588);
and U5728 (N_5728,N_4067,N_1736);
xor U5729 (N_5729,N_2096,N_1386);
nor U5730 (N_5730,N_4722,N_2120);
nand U5731 (N_5731,N_3208,N_4431);
and U5732 (N_5732,N_536,N_2664);
nand U5733 (N_5733,N_46,N_3194);
or U5734 (N_5734,N_2557,N_2023);
or U5735 (N_5735,N_1731,N_2924);
nand U5736 (N_5736,N_3849,N_2908);
nand U5737 (N_5737,N_3330,N_2856);
xnor U5738 (N_5738,N_1441,N_750);
or U5739 (N_5739,N_195,N_783);
or U5740 (N_5740,N_4136,N_1554);
and U5741 (N_5741,N_2379,N_226);
nor U5742 (N_5742,N_2753,N_2666);
nand U5743 (N_5743,N_1437,N_784);
and U5744 (N_5744,N_2890,N_702);
nand U5745 (N_5745,N_4711,N_1429);
and U5746 (N_5746,N_2388,N_1798);
or U5747 (N_5747,N_4,N_4396);
xnor U5748 (N_5748,N_3058,N_2285);
and U5749 (N_5749,N_4453,N_395);
nor U5750 (N_5750,N_1144,N_3558);
or U5751 (N_5751,N_1474,N_878);
or U5752 (N_5752,N_4339,N_3689);
xnor U5753 (N_5753,N_4787,N_2638);
xnor U5754 (N_5754,N_1891,N_884);
nor U5755 (N_5755,N_1770,N_1659);
or U5756 (N_5756,N_631,N_789);
nor U5757 (N_5757,N_2005,N_4581);
nand U5758 (N_5758,N_2389,N_3382);
or U5759 (N_5759,N_3088,N_1774);
or U5760 (N_5760,N_3600,N_3514);
or U5761 (N_5761,N_360,N_527);
nor U5762 (N_5762,N_4052,N_1228);
or U5763 (N_5763,N_4668,N_1589);
and U5764 (N_5764,N_1074,N_1131);
nand U5765 (N_5765,N_4130,N_3245);
or U5766 (N_5766,N_3484,N_1138);
and U5767 (N_5767,N_2618,N_4017);
or U5768 (N_5768,N_398,N_785);
or U5769 (N_5769,N_3481,N_2516);
nor U5770 (N_5770,N_2728,N_3394);
nand U5771 (N_5771,N_2300,N_1255);
or U5772 (N_5772,N_4595,N_674);
xnor U5773 (N_5773,N_4699,N_3698);
nor U5774 (N_5774,N_3037,N_3516);
and U5775 (N_5775,N_3177,N_1331);
and U5776 (N_5776,N_1178,N_2088);
xnor U5777 (N_5777,N_1197,N_3408);
xnor U5778 (N_5778,N_2685,N_1885);
or U5779 (N_5779,N_2359,N_74);
nor U5780 (N_5780,N_4220,N_4871);
nand U5781 (N_5781,N_1646,N_3984);
nand U5782 (N_5782,N_4963,N_1652);
nand U5783 (N_5783,N_539,N_130);
nor U5784 (N_5784,N_2340,N_1618);
or U5785 (N_5785,N_4550,N_3668);
xor U5786 (N_5786,N_1846,N_3607);
and U5787 (N_5787,N_155,N_4028);
or U5788 (N_5788,N_284,N_1252);
or U5789 (N_5789,N_2793,N_1906);
or U5790 (N_5790,N_4731,N_34);
xor U5791 (N_5791,N_4122,N_4750);
and U5792 (N_5792,N_3727,N_2403);
and U5793 (N_5793,N_71,N_2431);
or U5794 (N_5794,N_1494,N_1209);
and U5795 (N_5795,N_2724,N_534);
and U5796 (N_5796,N_2405,N_2675);
and U5797 (N_5797,N_1008,N_10);
xor U5798 (N_5798,N_740,N_4043);
xnor U5799 (N_5799,N_2877,N_2321);
and U5800 (N_5800,N_3722,N_4348);
xor U5801 (N_5801,N_822,N_4674);
nand U5802 (N_5802,N_3742,N_1316);
and U5803 (N_5803,N_1693,N_291);
and U5804 (N_5804,N_1905,N_3787);
xnor U5805 (N_5805,N_3879,N_3367);
nor U5806 (N_5806,N_3816,N_707);
nor U5807 (N_5807,N_9,N_4598);
nand U5808 (N_5808,N_3824,N_2722);
and U5809 (N_5809,N_45,N_1668);
nand U5810 (N_5810,N_1168,N_2676);
or U5811 (N_5811,N_3928,N_3774);
and U5812 (N_5812,N_2391,N_2660);
xor U5813 (N_5813,N_4738,N_3813);
xnor U5814 (N_5814,N_2469,N_2299);
and U5815 (N_5815,N_2028,N_551);
and U5816 (N_5816,N_3264,N_3948);
xnor U5817 (N_5817,N_2603,N_1149);
nand U5818 (N_5818,N_2947,N_4764);
xor U5819 (N_5819,N_4654,N_1061);
and U5820 (N_5820,N_2351,N_2872);
or U5821 (N_5821,N_2295,N_1976);
xnor U5822 (N_5822,N_3215,N_4305);
nor U5823 (N_5823,N_4330,N_2191);
and U5824 (N_5824,N_2121,N_219);
and U5825 (N_5825,N_3056,N_2198);
nand U5826 (N_5826,N_3109,N_1179);
and U5827 (N_5827,N_2522,N_1678);
nand U5828 (N_5828,N_1349,N_407);
and U5829 (N_5829,N_4239,N_1297);
nand U5830 (N_5830,N_3888,N_4150);
or U5831 (N_5831,N_3493,N_3238);
nand U5832 (N_5832,N_1274,N_3273);
xnor U5833 (N_5833,N_1117,N_4144);
nor U5834 (N_5834,N_3863,N_4862);
nand U5835 (N_5835,N_3613,N_3846);
xor U5836 (N_5836,N_4197,N_433);
nor U5837 (N_5837,N_97,N_2358);
or U5838 (N_5838,N_4936,N_3440);
nand U5839 (N_5839,N_1644,N_1060);
or U5840 (N_5840,N_4066,N_1066);
xnor U5841 (N_5841,N_2476,N_638);
nor U5842 (N_5842,N_4265,N_4479);
nor U5843 (N_5843,N_2105,N_2713);
nor U5844 (N_5844,N_1994,N_4341);
nand U5845 (N_5845,N_520,N_2861);
and U5846 (N_5846,N_4426,N_1245);
nor U5847 (N_5847,N_4238,N_2773);
xor U5848 (N_5848,N_4493,N_1027);
xnor U5849 (N_5849,N_1596,N_1164);
and U5850 (N_5850,N_880,N_710);
or U5851 (N_5851,N_2818,N_1872);
xor U5852 (N_5852,N_3345,N_2152);
nor U5853 (N_5853,N_1382,N_4917);
nand U5854 (N_5854,N_4617,N_1672);
or U5855 (N_5855,N_4525,N_76);
or U5856 (N_5856,N_3826,N_3120);
or U5857 (N_5857,N_2015,N_3404);
xor U5858 (N_5858,N_426,N_1309);
nor U5859 (N_5859,N_1811,N_1874);
or U5860 (N_5860,N_3216,N_1564);
or U5861 (N_5861,N_3304,N_4629);
or U5862 (N_5862,N_2397,N_1680);
and U5863 (N_5863,N_4389,N_2911);
and U5864 (N_5864,N_3457,N_2876);
or U5865 (N_5865,N_2550,N_1501);
nor U5866 (N_5866,N_739,N_2094);
xnor U5867 (N_5867,N_1720,N_4300);
xor U5868 (N_5868,N_4118,N_1665);
nor U5869 (N_5869,N_1390,N_657);
nand U5870 (N_5870,N_3105,N_1257);
nand U5871 (N_5871,N_4500,N_1725);
nand U5872 (N_5872,N_573,N_3628);
nand U5873 (N_5873,N_4716,N_980);
and U5874 (N_5874,N_1004,N_2700);
xor U5875 (N_5875,N_648,N_1671);
nor U5876 (N_5876,N_4850,N_2160);
nor U5877 (N_5877,N_1781,N_1982);
xnor U5878 (N_5878,N_167,N_1884);
nand U5879 (N_5879,N_3317,N_3570);
xor U5880 (N_5880,N_3716,N_723);
and U5881 (N_5881,N_8,N_1551);
xnor U5882 (N_5882,N_2806,N_3561);
or U5883 (N_5883,N_85,N_3602);
xor U5884 (N_5884,N_4828,N_2272);
nor U5885 (N_5885,N_249,N_2898);
nand U5886 (N_5886,N_4926,N_4355);
xnor U5887 (N_5887,N_2375,N_4425);
nor U5888 (N_5888,N_4209,N_2921);
and U5889 (N_5889,N_1130,N_302);
nand U5890 (N_5890,N_493,N_180);
and U5891 (N_5891,N_4268,N_2882);
and U5892 (N_5892,N_4719,N_299);
or U5893 (N_5893,N_3182,N_2706);
nor U5894 (N_5894,N_787,N_2201);
xnor U5895 (N_5895,N_3518,N_3425);
xor U5896 (N_5896,N_2776,N_4119);
xor U5897 (N_5897,N_817,N_4257);
xor U5898 (N_5898,N_3235,N_1145);
xor U5899 (N_5899,N_139,N_382);
nand U5900 (N_5900,N_4652,N_1650);
xor U5901 (N_5901,N_1878,N_835);
xnor U5902 (N_5902,N_3963,N_4610);
nor U5903 (N_5903,N_3704,N_1428);
nand U5904 (N_5904,N_4554,N_2841);
nor U5905 (N_5905,N_1115,N_4876);
nand U5906 (N_5906,N_3380,N_777);
and U5907 (N_5907,N_210,N_4510);
nand U5908 (N_5908,N_4319,N_3203);
and U5909 (N_5909,N_4563,N_1350);
and U5910 (N_5910,N_2750,N_1833);
and U5911 (N_5911,N_3094,N_860);
nand U5912 (N_5912,N_192,N_4206);
or U5913 (N_5913,N_4381,N_4367);
or U5914 (N_5914,N_4138,N_2410);
nor U5915 (N_5915,N_4684,N_1917);
nor U5916 (N_5916,N_3749,N_3971);
or U5917 (N_5917,N_1682,N_3839);
xnor U5918 (N_5918,N_4657,N_3007);
xor U5919 (N_5919,N_2423,N_4084);
nor U5920 (N_5920,N_4683,N_87);
nor U5921 (N_5921,N_2032,N_3283);
nand U5922 (N_5922,N_2278,N_372);
or U5923 (N_5923,N_1338,N_2659);
and U5924 (N_5924,N_748,N_4918);
nor U5925 (N_5925,N_251,N_3907);
nand U5926 (N_5926,N_562,N_4882);
xor U5927 (N_5927,N_823,N_4492);
nor U5928 (N_5928,N_369,N_743);
and U5929 (N_5929,N_1416,N_4233);
xor U5930 (N_5930,N_1654,N_794);
nor U5931 (N_5931,N_3881,N_2916);
nand U5932 (N_5932,N_4258,N_1125);
or U5933 (N_5933,N_4608,N_1769);
nor U5934 (N_5934,N_572,N_250);
xor U5935 (N_5935,N_1757,N_460);
or U5936 (N_5936,N_4465,N_1018);
and U5937 (N_5937,N_3932,N_3123);
and U5938 (N_5938,N_4635,N_3349);
and U5939 (N_5939,N_3771,N_1529);
nand U5940 (N_5940,N_4000,N_2442);
xor U5941 (N_5941,N_1890,N_3564);
or U5942 (N_5942,N_4082,N_2854);
nor U5943 (N_5943,N_4496,N_3887);
nor U5944 (N_5944,N_2441,N_2030);
nor U5945 (N_5945,N_2341,N_3856);
and U5946 (N_5946,N_1113,N_3050);
xnor U5947 (N_5947,N_3347,N_3845);
and U5948 (N_5948,N_2166,N_2973);
nor U5949 (N_5949,N_3360,N_3323);
or U5950 (N_5950,N_4877,N_987);
xor U5951 (N_5951,N_2711,N_3621);
nand U5952 (N_5952,N_4338,N_1063);
nor U5953 (N_5953,N_3390,N_1047);
or U5954 (N_5954,N_3302,N_1949);
nand U5955 (N_5955,N_3366,N_1694);
nor U5956 (N_5956,N_523,N_2214);
nand U5957 (N_5957,N_4853,N_1916);
xnor U5958 (N_5958,N_725,N_708);
and U5959 (N_5959,N_4142,N_3786);
and U5960 (N_5960,N_4223,N_1058);
xor U5961 (N_5961,N_2184,N_3009);
xor U5962 (N_5962,N_4102,N_4384);
xor U5963 (N_5963,N_4729,N_160);
nor U5964 (N_5964,N_1108,N_440);
xnor U5965 (N_5965,N_718,N_4484);
xnor U5966 (N_5966,N_1743,N_524);
nor U5967 (N_5967,N_1804,N_4947);
or U5968 (N_5968,N_1039,N_3491);
xnor U5969 (N_5969,N_303,N_827);
nand U5970 (N_5970,N_2142,N_1943);
nand U5971 (N_5971,N_3625,N_892);
xor U5972 (N_5972,N_4362,N_1828);
and U5973 (N_5973,N_1279,N_1962);
nand U5974 (N_5974,N_4864,N_2602);
nor U5975 (N_5975,N_1041,N_2653);
or U5976 (N_5976,N_416,N_4309);
nand U5977 (N_5977,N_564,N_3469);
nor U5978 (N_5978,N_2367,N_3548);
and U5979 (N_5979,N_3334,N_550);
or U5980 (N_5980,N_2553,N_334);
or U5981 (N_5981,N_3513,N_2817);
or U5982 (N_5982,N_2701,N_3870);
xnor U5983 (N_5983,N_4212,N_4376);
and U5984 (N_5984,N_3998,N_1483);
xnor U5985 (N_5985,N_4188,N_3192);
or U5986 (N_5986,N_4124,N_3178);
nor U5987 (N_5987,N_2240,N_3288);
nand U5988 (N_5988,N_3780,N_3785);
nand U5989 (N_5989,N_410,N_2324);
or U5990 (N_5990,N_3396,N_4053);
and U5991 (N_5991,N_1937,N_1439);
and U5992 (N_5992,N_905,N_1477);
nand U5993 (N_5993,N_2357,N_3140);
xor U5994 (N_5994,N_1744,N_4312);
xor U5995 (N_5995,N_3076,N_4191);
xnor U5996 (N_5996,N_3919,N_4548);
nand U5997 (N_5997,N_2211,N_2104);
xor U5998 (N_5998,N_1110,N_4112);
xor U5999 (N_5999,N_1606,N_4761);
xor U6000 (N_6000,N_528,N_3729);
nor U6001 (N_6001,N_1489,N_4650);
nand U6002 (N_6002,N_4442,N_3885);
or U6003 (N_6003,N_376,N_1637);
nor U6004 (N_6004,N_1015,N_1607);
or U6005 (N_6005,N_3375,N_1409);
nor U6006 (N_6006,N_1706,N_4502);
and U6007 (N_6007,N_3133,N_2116);
xor U6008 (N_6008,N_1873,N_778);
xnor U6009 (N_6009,N_1581,N_3979);
nand U6010 (N_6010,N_4892,N_1805);
and U6011 (N_6011,N_697,N_2428);
and U6012 (N_6012,N_111,N_3496);
nor U6013 (N_6013,N_2765,N_1096);
or U6014 (N_6014,N_2763,N_1926);
nor U6015 (N_6015,N_2322,N_234);
xor U6016 (N_6016,N_3124,N_3106);
and U6017 (N_6017,N_4103,N_190);
or U6018 (N_6018,N_4830,N_29);
nand U6019 (N_6019,N_1159,N_2065);
xor U6020 (N_6020,N_43,N_1717);
or U6021 (N_6021,N_679,N_1985);
nand U6022 (N_6022,N_4480,N_3149);
xnor U6023 (N_6023,N_4771,N_129);
xor U6024 (N_6024,N_1996,N_3594);
nand U6025 (N_6025,N_1503,N_194);
nor U6026 (N_6026,N_4452,N_1302);
and U6027 (N_6027,N_2868,N_3355);
nor U6028 (N_6028,N_977,N_310);
xnor U6029 (N_6029,N_4462,N_598);
nor U6030 (N_6030,N_3873,N_2194);
nand U6031 (N_6031,N_3449,N_2878);
and U6032 (N_6032,N_3035,N_3647);
nand U6033 (N_6033,N_3789,N_696);
and U6034 (N_6034,N_4768,N_3479);
xor U6035 (N_6035,N_866,N_358);
and U6036 (N_6036,N_3164,N_1573);
and U6037 (N_6037,N_1808,N_2009);
nor U6038 (N_6038,N_3358,N_4414);
nor U6039 (N_6039,N_2221,N_2740);
xnor U6040 (N_6040,N_1229,N_2785);
xor U6041 (N_6041,N_330,N_19);
xor U6042 (N_6042,N_2958,N_1728);
xor U6043 (N_6043,N_1907,N_931);
or U6044 (N_6044,N_2650,N_4647);
and U6045 (N_6045,N_4814,N_2577);
or U6046 (N_6046,N_329,N_1705);
and U6047 (N_6047,N_1154,N_128);
nand U6048 (N_6048,N_4760,N_1676);
nand U6049 (N_6049,N_274,N_1273);
and U6050 (N_6050,N_4261,N_2466);
nor U6051 (N_6051,N_212,N_2780);
xor U6052 (N_6052,N_177,N_1172);
or U6053 (N_6053,N_1107,N_1198);
or U6054 (N_6054,N_454,N_3914);
nor U6055 (N_6055,N_2845,N_1541);
nor U6056 (N_6056,N_4863,N_2580);
or U6057 (N_6057,N_4282,N_733);
nor U6058 (N_6058,N_1079,N_4013);
and U6059 (N_6059,N_2435,N_2613);
xor U6060 (N_6060,N_639,N_2137);
and U6061 (N_6061,N_2150,N_2080);
nand U6062 (N_6062,N_4848,N_3122);
nor U6063 (N_6063,N_4415,N_4098);
or U6064 (N_6064,N_2503,N_3829);
and U6065 (N_6065,N_4819,N_2193);
xnor U6066 (N_6066,N_1369,N_3295);
or U6067 (N_6067,N_2422,N_1667);
and U6068 (N_6068,N_2118,N_2933);
xor U6069 (N_6069,N_2555,N_4200);
or U6070 (N_6070,N_4905,N_1945);
nand U6071 (N_6071,N_1346,N_578);
xor U6072 (N_6072,N_1286,N_393);
and U6073 (N_6073,N_4080,N_3803);
nor U6074 (N_6074,N_1360,N_2250);
or U6075 (N_6075,N_4278,N_2764);
or U6076 (N_6076,N_2985,N_4995);
nand U6077 (N_6077,N_1223,N_1912);
and U6078 (N_6078,N_1555,N_1243);
and U6079 (N_6079,N_1908,N_3401);
or U6080 (N_6080,N_4658,N_4151);
or U6081 (N_6081,N_2161,N_4898);
xnor U6082 (N_6082,N_2608,N_2294);
and U6083 (N_6083,N_1040,N_4145);
and U6084 (N_6084,N_3233,N_2042);
nand U6085 (N_6085,N_3683,N_3955);
or U6086 (N_6086,N_587,N_590);
or U6087 (N_6087,N_810,N_4474);
nand U6088 (N_6088,N_3661,N_3775);
nor U6089 (N_6089,N_3016,N_3381);
nand U6090 (N_6090,N_1611,N_803);
and U6091 (N_6091,N_1304,N_2230);
or U6092 (N_6092,N_4861,N_1162);
and U6093 (N_6093,N_1330,N_1119);
nand U6094 (N_6094,N_2982,N_3132);
nor U6095 (N_6095,N_2177,N_4064);
or U6096 (N_6096,N_2025,N_368);
xor U6097 (N_6097,N_3437,N_3204);
or U6098 (N_6098,N_3303,N_1656);
or U6099 (N_6099,N_2732,N_1664);
or U6100 (N_6100,N_4405,N_1205);
nand U6101 (N_6101,N_1839,N_1940);
nor U6102 (N_6102,N_213,N_1368);
or U6103 (N_6103,N_2251,N_2848);
or U6104 (N_6104,N_2524,N_1264);
and U6105 (N_6105,N_4298,N_2187);
nand U6106 (N_6106,N_661,N_914);
or U6107 (N_6107,N_3761,N_3383);
and U6108 (N_6108,N_1512,N_2767);
and U6109 (N_6109,N_3580,N_751);
or U6110 (N_6110,N_6,N_4275);
xor U6111 (N_6111,N_2216,N_4601);
and U6112 (N_6112,N_3364,N_3808);
xor U6113 (N_6113,N_4669,N_3427);
and U6114 (N_6114,N_126,N_1681);
nor U6115 (N_6115,N_370,N_4979);
or U6116 (N_6116,N_2745,N_2304);
nor U6117 (N_6117,N_4143,N_2165);
or U6118 (N_6118,N_2237,N_4324);
xnor U6119 (N_6119,N_1383,N_182);
or U6120 (N_6120,N_3687,N_4815);
xor U6121 (N_6121,N_1797,N_3010);
nor U6122 (N_6122,N_4398,N_2273);
and U6123 (N_6123,N_1931,N_4565);
xor U6124 (N_6124,N_1862,N_452);
xor U6125 (N_6125,N_4961,N_4128);
nand U6126 (N_6126,N_967,N_3418);
nand U6127 (N_6127,N_3062,N_3402);
or U6128 (N_6128,N_1800,N_4420);
and U6129 (N_6129,N_2652,N_4301);
nand U6130 (N_6130,N_4478,N_2777);
nand U6131 (N_6131,N_1269,N_1440);
or U6132 (N_6132,N_669,N_4329);
nand U6133 (N_6133,N_1772,N_3444);
and U6134 (N_6134,N_3474,N_678);
or U6135 (N_6135,N_441,N_2064);
xor U6136 (N_6136,N_105,N_1460);
xnor U6137 (N_6137,N_1420,N_3618);
xnor U6138 (N_6138,N_1232,N_2672);
and U6139 (N_6139,N_3610,N_894);
xor U6140 (N_6140,N_1408,N_4123);
nand U6141 (N_6141,N_243,N_4968);
nor U6142 (N_6142,N_851,N_3547);
xor U6143 (N_6143,N_4436,N_3168);
nand U6144 (N_6144,N_1318,N_2122);
nor U6145 (N_6145,N_4110,N_2556);
nand U6146 (N_6146,N_3694,N_396);
nand U6147 (N_6147,N_3604,N_4523);
xor U6148 (N_6148,N_3875,N_1335);
xor U6149 (N_6149,N_3964,N_964);
nor U6150 (N_6150,N_4382,N_1898);
xor U6151 (N_6151,N_2781,N_1636);
xnor U6152 (N_6152,N_1388,N_4352);
nor U6153 (N_6153,N_3144,N_3042);
or U6154 (N_6154,N_4883,N_4002);
nand U6155 (N_6155,N_3102,N_2729);
nand U6156 (N_6156,N_3338,N_4010);
nand U6157 (N_6157,N_184,N_1259);
xnor U6158 (N_6158,N_3379,N_711);
nor U6159 (N_6159,N_3951,N_3987);
and U6160 (N_6160,N_2430,N_2605);
nand U6161 (N_6161,N_1432,N_4140);
nor U6162 (N_6162,N_1834,N_887);
nand U6163 (N_6163,N_2332,N_1464);
nand U6164 (N_6164,N_2000,N_3108);
nor U6165 (N_6165,N_2280,N_3008);
and U6166 (N_6166,N_3270,N_282);
xor U6167 (N_6167,N_1763,N_1929);
nor U6168 (N_6168,N_4740,N_1050);
xor U6169 (N_6169,N_4125,N_2951);
or U6170 (N_6170,N_955,N_3905);
nor U6171 (N_6171,N_2220,N_776);
xor U6172 (N_6172,N_1788,N_1776);
nand U6173 (N_6173,N_327,N_2305);
xnor U6174 (N_6174,N_1051,N_3419);
nand U6175 (N_6175,N_4322,N_4250);
nand U6176 (N_6176,N_4569,N_3325);
xor U6177 (N_6177,N_923,N_935);
nor U6178 (N_6178,N_1972,N_353);
and U6179 (N_6179,N_57,N_3622);
nand U6180 (N_6180,N_1275,N_2490);
xnor U6181 (N_6181,N_3282,N_2426);
xnor U6182 (N_6182,N_4042,N_4476);
or U6183 (N_6183,N_3744,N_1171);
and U6184 (N_6184,N_315,N_196);
and U6185 (N_6185,N_2227,N_3117);
or U6186 (N_6186,N_2021,N_298);
nand U6187 (N_6187,N_4490,N_2542);
xor U6188 (N_6188,N_3920,N_3991);
nor U6189 (N_6189,N_485,N_2427);
and U6190 (N_6190,N_1810,N_4560);
or U6191 (N_6191,N_3063,N_4810);
and U6192 (N_6192,N_1924,N_736);
xnor U6193 (N_6193,N_1612,N_1585);
nor U6194 (N_6194,N_1397,N_3291);
nand U6195 (N_6195,N_471,N_1963);
nand U6196 (N_6196,N_918,N_2619);
and U6197 (N_6197,N_3041,N_1570);
nand U6198 (N_6198,N_3281,N_1052);
and U6199 (N_6199,N_588,N_4944);
nand U6200 (N_6200,N_468,N_1954);
nor U6201 (N_6201,N_305,N_566);
xnor U6202 (N_6202,N_1735,N_3307);
nand U6203 (N_6203,N_490,N_2508);
nor U6204 (N_6204,N_3623,N_1);
and U6205 (N_6205,N_3751,N_901);
and U6206 (N_6206,N_3116,N_845);
or U6207 (N_6207,N_2723,N_3463);
xnor U6208 (N_6208,N_1044,N_4464);
nor U6209 (N_6209,N_2144,N_4985);
or U6210 (N_6210,N_1002,N_2387);
or U6211 (N_6211,N_874,N_4108);
nor U6212 (N_6212,N_4246,N_4632);
and U6213 (N_6213,N_110,N_3414);
nor U6214 (N_6214,N_4758,N_3965);
xor U6215 (N_6215,N_693,N_3943);
xnor U6216 (N_6216,N_4980,N_1698);
and U6217 (N_6217,N_54,N_1969);
and U6218 (N_6218,N_3533,N_1819);
nand U6219 (N_6219,N_809,N_3681);
xnor U6220 (N_6220,N_2792,N_616);
and U6221 (N_6221,N_3973,N_950);
xor U6222 (N_6222,N_3495,N_910);
nand U6223 (N_6223,N_3844,N_3927);
nor U6224 (N_6224,N_2590,N_185);
xor U6225 (N_6225,N_4256,N_4366);
nand U6226 (N_6226,N_1925,N_3719);
nor U6227 (N_6227,N_1827,N_1217);
and U6228 (N_6228,N_4852,N_3847);
and U6229 (N_6229,N_3486,N_2862);
xor U6230 (N_6230,N_4116,N_4960);
or U6231 (N_6231,N_4651,N_865);
or U6232 (N_6232,N_3890,N_4620);
and U6233 (N_6233,N_3537,N_3897);
and U6234 (N_6234,N_1342,N_4997);
and U6235 (N_6235,N_3501,N_1075);
or U6236 (N_6236,N_1930,N_388);
and U6237 (N_6237,N_4354,N_3019);
nor U6238 (N_6238,N_102,N_64);
xnor U6239 (N_6239,N_3372,N_3251);
or U6240 (N_6240,N_4021,N_1277);
or U6241 (N_6241,N_1365,N_2687);
nand U6242 (N_6242,N_108,N_3446);
nor U6243 (N_6243,N_216,N_3130);
or U6244 (N_6244,N_1825,N_2421);
nor U6245 (N_6245,N_351,N_1387);
nand U6246 (N_6246,N_4880,N_4105);
or U6247 (N_6247,N_1683,N_2520);
nor U6248 (N_6248,N_2606,N_1357);
nand U6249 (N_6249,N_1267,N_759);
xor U6250 (N_6250,N_3336,N_1524);
nand U6251 (N_6251,N_994,N_4127);
xnor U6252 (N_6252,N_4707,N_3136);
and U6253 (N_6253,N_3843,N_3883);
nor U6254 (N_6254,N_32,N_113);
and U6255 (N_6255,N_4019,N_496);
or U6256 (N_6256,N_375,N_2162);
and U6257 (N_6257,N_3174,N_1511);
nor U6258 (N_6258,N_4542,N_1373);
and U6259 (N_6259,N_307,N_946);
or U6260 (N_6260,N_3910,N_575);
nor U6261 (N_6261,N_3022,N_1594);
xnor U6262 (N_6262,N_3459,N_546);
xnor U6263 (N_6263,N_1964,N_2970);
nand U6264 (N_6264,N_92,N_1049);
and U6265 (N_6265,N_4406,N_341);
xor U6266 (N_6266,N_1449,N_31);
and U6267 (N_6267,N_1701,N_2988);
nand U6268 (N_6268,N_658,N_253);
or U6269 (N_6269,N_1777,N_3958);
nand U6270 (N_6270,N_2277,N_2033);
nand U6271 (N_6271,N_2018,N_4161);
and U6272 (N_6272,N_199,N_4645);
and U6273 (N_6273,N_2938,N_1445);
nor U6274 (N_6274,N_3098,N_599);
nor U6275 (N_6275,N_146,N_293);
and U6276 (N_6276,N_726,N_4599);
or U6277 (N_6277,N_2527,N_4056);
nand U6278 (N_6278,N_2362,N_288);
or U6279 (N_6279,N_201,N_3197);
and U6280 (N_6280,N_4568,N_2984);
nand U6281 (N_6281,N_1858,N_2528);
xor U6282 (N_6282,N_2154,N_841);
nand U6283 (N_6283,N_2434,N_3790);
nand U6284 (N_6284,N_4201,N_4941);
and U6285 (N_6285,N_2197,N_1212);
nand U6286 (N_6286,N_3143,N_4730);
xor U6287 (N_6287,N_3434,N_2048);
nand U6288 (N_6288,N_2219,N_2098);
xnor U6289 (N_6289,N_4741,N_2547);
or U6290 (N_6290,N_2545,N_4316);
and U6291 (N_6291,N_1443,N_3068);
nand U6292 (N_6292,N_1806,N_4167);
or U6293 (N_6293,N_629,N_552);
nand U6294 (N_6294,N_2510,N_3236);
nor U6295 (N_6295,N_2353,N_3032);
xnor U6296 (N_6296,N_4323,N_4965);
xor U6297 (N_6297,N_3354,N_2365);
or U6298 (N_6298,N_3640,N_2497);
and U6299 (N_6299,N_667,N_2695);
or U6300 (N_6300,N_1609,N_3511);
nor U6301 (N_6301,N_4410,N_4969);
nor U6302 (N_6302,N_3690,N_3508);
xor U6303 (N_6303,N_198,N_593);
nor U6304 (N_6304,N_3568,N_301);
nor U6305 (N_6305,N_1790,N_2671);
nor U6306 (N_6306,N_1843,N_1584);
or U6307 (N_6307,N_644,N_450);
nand U6308 (N_6308,N_4248,N_3903);
nand U6309 (N_6309,N_2987,N_4675);
nor U6310 (N_6310,N_1478,N_2222);
and U6311 (N_6311,N_1375,N_4779);
or U6312 (N_6312,N_2900,N_3301);
xnor U6313 (N_6313,N_3498,N_3229);
nand U6314 (N_6314,N_479,N_4321);
nand U6315 (N_6315,N_1152,N_63);
nand U6316 (N_6316,N_2986,N_522);
and U6317 (N_6317,N_2087,N_1495);
or U6318 (N_6318,N_525,N_3868);
and U6319 (N_6319,N_2420,N_4612);
nor U6320 (N_6320,N_3523,N_4203);
and U6321 (N_6321,N_1730,N_547);
and U6322 (N_6322,N_4393,N_3642);
nand U6323 (N_6323,N_1505,N_3754);
and U6324 (N_6324,N_1697,N_2725);
or U6325 (N_6325,N_1651,N_4299);
xor U6326 (N_6326,N_4856,N_1374);
nor U6327 (N_6327,N_4766,N_2241);
nor U6328 (N_6328,N_2407,N_1634);
xor U6329 (N_6329,N_2858,N_1237);
nor U6330 (N_6330,N_951,N_3941);
and U6331 (N_6331,N_2478,N_1414);
xor U6332 (N_6332,N_3865,N_1045);
nor U6333 (N_6333,N_3318,N_1984);
nor U6334 (N_6334,N_316,N_3435);
xor U6335 (N_6335,N_4948,N_4867);
nor U6336 (N_6336,N_1046,N_1626);
xor U6337 (N_6337,N_2190,N_1786);
nand U6338 (N_6338,N_2914,N_3934);
xnor U6339 (N_6339,N_4870,N_3369);
or U6340 (N_6340,N_4920,N_356);
nand U6341 (N_6341,N_1699,N_1739);
nor U6342 (N_6342,N_4618,N_3445);
nor U6343 (N_6343,N_996,N_4886);
nand U6344 (N_6344,N_1139,N_844);
and U6345 (N_6345,N_269,N_1158);
nand U6346 (N_6346,N_800,N_2127);
and U6347 (N_6347,N_4177,N_1540);
or U6348 (N_6348,N_1344,N_1006);
and U6349 (N_6349,N_2401,N_4131);
nand U6350 (N_6350,N_656,N_3524);
xnor U6351 (N_6351,N_3848,N_2850);
and U6352 (N_6352,N_3014,N_279);
xnor U6353 (N_6353,N_699,N_4718);
and U6354 (N_6354,N_654,N_1163);
or U6355 (N_6355,N_3763,N_448);
nand U6356 (N_6356,N_1669,N_1123);
nand U6357 (N_6357,N_1156,N_500);
and U6358 (N_6358,N_676,N_3095);
xnor U6359 (N_6359,N_4368,N_4833);
nor U6360 (N_6360,N_2384,N_3728);
nand U6361 (N_6361,N_2262,N_3904);
nor U6362 (N_6362,N_413,N_4835);
or U6363 (N_6363,N_885,N_2960);
nor U6364 (N_6364,N_259,N_1415);
nand U6365 (N_6365,N_2625,N_1213);
nor U6366 (N_6366,N_501,N_3311);
nor U6367 (N_6367,N_352,N_1490);
xnor U6368 (N_6368,N_3697,N_3901);
or U6369 (N_6369,N_1268,N_4372);
nor U6370 (N_6370,N_2020,N_242);
nor U6371 (N_6371,N_4171,N_3483);
or U6372 (N_6372,N_632,N_187);
or U6373 (N_6373,N_4984,N_3240);
nor U6374 (N_6374,N_600,N_4327);
nor U6375 (N_6375,N_4742,N_4812);
and U6376 (N_6376,N_2485,N_4501);
nand U6377 (N_6377,N_1249,N_3166);
and U6378 (N_6378,N_2568,N_367);
nand U6379 (N_6379,N_4637,N_653);
nand U6380 (N_6380,N_3458,N_1292);
xnor U6381 (N_6381,N_2826,N_2719);
or U6382 (N_6382,N_1578,N_30);
and U6383 (N_6383,N_3794,N_4546);
xor U6384 (N_6384,N_2100,N_4285);
nand U6385 (N_6385,N_3313,N_2518);
and U6386 (N_6386,N_2186,N_1076);
nand U6387 (N_6387,N_2415,N_4954);
xor U6388 (N_6388,N_3279,N_2019);
nand U6389 (N_6389,N_4343,N_2786);
nor U6390 (N_6390,N_444,N_2313);
xor U6391 (N_6391,N_4616,N_3373);
nor U6392 (N_6392,N_3969,N_3956);
or U6393 (N_6393,N_3777,N_3930);
or U6394 (N_6394,N_4522,N_2931);
nand U6395 (N_6395,N_2670,N_1639);
nand U6396 (N_6396,N_1602,N_3139);
and U6397 (N_6397,N_2529,N_383);
or U6398 (N_6398,N_482,N_3034);
xor U6399 (N_6399,N_4585,N_728);
xor U6400 (N_6400,N_3859,N_2130);
or U6401 (N_6401,N_2983,N_1143);
nand U6402 (N_6402,N_4380,N_2511);
xnor U6403 (N_6403,N_99,N_4507);
xnor U6404 (N_6404,N_2805,N_44);
nor U6405 (N_6405,N_4712,N_481);
xnor U6406 (N_6406,N_3747,N_4720);
or U6407 (N_6407,N_3572,N_4214);
nand U6408 (N_6408,N_4866,N_1332);
nor U6409 (N_6409,N_1486,N_3046);
and U6410 (N_6410,N_4932,N_3141);
and U6411 (N_6411,N_4293,N_3091);
and U6412 (N_6412,N_3585,N_3703);
and U6413 (N_6413,N_1080,N_3574);
xor U6414 (N_6414,N_311,N_795);
and U6415 (N_6415,N_1482,N_1871);
or U6416 (N_6416,N_4009,N_768);
nor U6417 (N_6417,N_3494,N_1913);
or U6418 (N_6418,N_902,N_1084);
nor U6419 (N_6419,N_921,N_3156);
xor U6420 (N_6420,N_3411,N_2402);
nand U6421 (N_6421,N_2582,N_3735);
nand U6422 (N_6422,N_2040,N_1703);
or U6423 (N_6423,N_1492,N_608);
or U6424 (N_6424,N_4481,N_812);
and U6425 (N_6425,N_592,N_1734);
nor U6426 (N_6426,N_828,N_1150);
nand U6427 (N_6427,N_1438,N_178);
nand U6428 (N_6428,N_1185,N_3550);
nor U6429 (N_6429,N_1062,N_1649);
or U6430 (N_6430,N_1325,N_3711);
or U6431 (N_6431,N_1960,N_3188);
nor U6432 (N_6432,N_2090,N_2134);
or U6433 (N_6433,N_3324,N_3595);
xnor U6434 (N_6434,N_4593,N_4403);
or U6435 (N_6435,N_2132,N_4325);
nor U6436 (N_6436,N_1450,N_277);
nand U6437 (N_6437,N_626,N_4786);
nand U6438 (N_6438,N_3223,N_937);
nor U6439 (N_6439,N_4065,N_4725);
nand U6440 (N_6440,N_3505,N_1324);
and U6441 (N_6441,N_476,N_1242);
xor U6442 (N_6442,N_4681,N_170);
nand U6443 (N_6443,N_4273,N_3039);
and U6444 (N_6444,N_51,N_814);
nand U6445 (N_6445,N_145,N_1481);
nor U6446 (N_6446,N_984,N_1563);
nor U6447 (N_6447,N_2377,N_2149);
or U6448 (N_6448,N_3362,N_2310);
xor U6449 (N_6449,N_3460,N_819);
nand U6450 (N_6450,N_3646,N_286);
nor U6451 (N_6451,N_684,N_928);
xor U6452 (N_6452,N_4516,N_3332);
and U6453 (N_6453,N_4915,N_3489);
xnor U6454 (N_6454,N_2231,N_3925);
xnor U6455 (N_6455,N_2049,N_17);
xnor U6456 (N_6456,N_206,N_891);
xnor U6457 (N_6457,N_2885,N_1463);
nand U6458 (N_6458,N_2247,N_2213);
xnor U6459 (N_6459,N_4547,N_3999);
xor U6460 (N_6460,N_671,N_2693);
or U6461 (N_6461,N_1087,N_502);
xnor U6462 (N_6462,N_3079,N_761);
nor U6463 (N_6463,N_2200,N_1370);
nand U6464 (N_6464,N_3150,N_4698);
and U6465 (N_6465,N_4164,N_3183);
nor U6466 (N_6466,N_4933,N_1758);
xnor U6467 (N_6467,N_3465,N_2062);
xnor U6468 (N_6468,N_804,N_907);
or U6469 (N_6469,N_1238,N_3171);
or U6470 (N_6470,N_2855,N_4421);
or U6471 (N_6471,N_4353,N_4989);
nor U6472 (N_6472,N_2255,N_2572);
and U6473 (N_6473,N_974,N_227);
or U6474 (N_6474,N_882,N_4971);
nand U6475 (N_6475,N_3954,N_280);
and U6476 (N_6476,N_4083,N_504);
nand U6477 (N_6477,N_4993,N_159);
nor U6478 (N_6478,N_2157,N_3706);
xnor U6479 (N_6479,N_3087,N_3520);
nor U6480 (N_6480,N_1317,N_4400);
or U6481 (N_6481,N_1459,N_1026);
and U6482 (N_6482,N_3,N_1580);
and U6483 (N_6483,N_4857,N_1696);
nand U6484 (N_6484,N_2293,N_3190);
and U6485 (N_6485,N_1733,N_957);
nand U6486 (N_6486,N_1662,N_3624);
nor U6487 (N_6487,N_2151,N_4267);
xor U6488 (N_6488,N_1067,N_4543);
and U6489 (N_6489,N_2859,N_4005);
nand U6490 (N_6490,N_781,N_2148);
nor U6491 (N_6491,N_1399,N_1866);
nor U6492 (N_6492,N_1613,N_2172);
nor U6493 (N_6493,N_2291,N_1347);
or U6494 (N_6494,N_2054,N_1543);
xor U6495 (N_6495,N_2844,N_3250);
and U6496 (N_6496,N_695,N_628);
or U6497 (N_6497,N_516,N_392);
nand U6498 (N_6498,N_3256,N_3666);
nor U6499 (N_6499,N_4364,N_755);
and U6500 (N_6500,N_1550,N_698);
nor U6501 (N_6501,N_2778,N_3092);
nand U6502 (N_6502,N_4391,N_2853);
nand U6503 (N_6503,N_3464,N_709);
and U6504 (N_6504,N_3320,N_3664);
or U6505 (N_6505,N_2893,N_2228);
or U6506 (N_6506,N_1624,N_477);
and U6507 (N_6507,N_2074,N_1708);
nor U6508 (N_6508,N_713,N_2604);
or U6509 (N_6509,N_2315,N_2487);
nand U6510 (N_6510,N_1716,N_347);
or U6511 (N_6511,N_1272,N_1028);
or U6512 (N_6512,N_879,N_1468);
nor U6513 (N_6513,N_2674,N_1549);
xor U6514 (N_6514,N_2991,N_4956);
nand U6515 (N_6515,N_2287,N_3257);
nand U6516 (N_6516,N_2314,N_2217);
nor U6517 (N_6517,N_620,N_3810);
or U6518 (N_6518,N_1377,N_4555);
and U6519 (N_6519,N_331,N_2819);
or U6520 (N_6520,N_3147,N_2816);
and U6521 (N_6521,N_2554,N_1633);
or U6522 (N_6522,N_2113,N_3603);
xor U6523 (N_6523,N_2268,N_4271);
xnor U6524 (N_6524,N_2298,N_495);
nor U6525 (N_6525,N_4477,N_4292);
xor U6526 (N_6526,N_2830,N_3576);
nor U6527 (N_6527,N_28,N_2196);
nor U6528 (N_6528,N_4078,N_2124);
nor U6529 (N_6529,N_4922,N_1565);
xnor U6530 (N_6530,N_4407,N_4710);
xnor U6531 (N_6531,N_20,N_2433);
nor U6532 (N_6532,N_2694,N_3731);
xor U6533 (N_6533,N_1082,N_1760);
xnor U6534 (N_6534,N_2798,N_1756);
xor U6535 (N_6535,N_1321,N_2051);
nor U6536 (N_6536,N_1009,N_3947);
and U6537 (N_6537,N_2346,N_3584);
and U6538 (N_6538,N_919,N_4222);
or U6539 (N_6539,N_4622,N_4524);
and U6540 (N_6540,N_3055,N_2812);
nor U6541 (N_6541,N_24,N_403);
or U6542 (N_6542,N_4628,N_677);
nor U6543 (N_6543,N_4378,N_4288);
xor U6544 (N_6544,N_4358,N_2549);
and U6545 (N_6545,N_389,N_2282);
and U6546 (N_6546,N_1007,N_3976);
or U6547 (N_6547,N_3992,N_1250);
and U6548 (N_6548,N_3230,N_4308);
and U6549 (N_6549,N_4606,N_4790);
and U6550 (N_6550,N_514,N_4897);
nand U6551 (N_6551,N_568,N_2045);
and U6552 (N_6552,N_961,N_4106);
nor U6553 (N_6553,N_4728,N_1177);
or U6554 (N_6554,N_1631,N_3224);
nand U6555 (N_6555,N_3371,N_3730);
nand U6556 (N_6556,N_1142,N_1741);
nand U6557 (N_6557,N_1419,N_735);
and U6558 (N_6558,N_3700,N_1953);
nor U6559 (N_6559,N_4195,N_4659);
or U6560 (N_6560,N_3125,N_439);
nand U6561 (N_6561,N_2164,N_4318);
xor U6562 (N_6562,N_3191,N_4770);
nor U6563 (N_6563,N_1077,N_2089);
nand U6564 (N_6564,N_2678,N_2185);
xnor U6565 (N_6565,N_2758,N_473);
or U6566 (N_6566,N_972,N_904);
nor U6567 (N_6567,N_3297,N_340);
nor U6568 (N_6568,N_1303,N_3851);
xor U6569 (N_6569,N_1533,N_2567);
nor U6570 (N_6570,N_1791,N_858);
or U6571 (N_6571,N_470,N_924);
nor U6572 (N_6572,N_4455,N_2133);
xnor U6573 (N_6573,N_2895,N_4283);
nand U6574 (N_6574,N_4902,N_3231);
nor U6575 (N_6575,N_1231,N_2443);
nor U6576 (N_6576,N_133,N_911);
or U6577 (N_6577,N_2515,N_4166);
xnor U6578 (N_6578,N_4038,N_2242);
nor U6579 (N_6579,N_3160,N_603);
and U6580 (N_6580,N_361,N_2480);
nor U6581 (N_6581,N_2783,N_633);
xnor U6582 (N_6582,N_2292,N_4175);
nand U6583 (N_6583,N_404,N_3531);
nand U6584 (N_6584,N_1900,N_1746);
xor U6585 (N_6585,N_1402,N_1822);
and U6586 (N_6586,N_1965,N_4245);
nor U6587 (N_6587,N_1395,N_2954);
or U6588 (N_6588,N_3121,N_4470);
nand U6589 (N_6589,N_2136,N_4310);
nand U6590 (N_6590,N_2235,N_3679);
or U6591 (N_6591,N_3717,N_3356);
and U6592 (N_6592,N_366,N_4289);
and U6593 (N_6593,N_1412,N_1134);
or U6594 (N_6594,N_2831,N_3321);
nor U6595 (N_6595,N_2063,N_3792);
or U6596 (N_6596,N_3405,N_4517);
nand U6597 (N_6597,N_4196,N_2998);
or U6598 (N_6598,N_3158,N_458);
or U6599 (N_6599,N_1240,N_2543);
nor U6600 (N_6600,N_2692,N_3592);
xnor U6601 (N_6601,N_2811,N_1993);
nand U6602 (N_6602,N_2072,N_3858);
nor U6603 (N_6603,N_4559,N_3983);
or U6604 (N_6604,N_4520,N_4611);
nor U6605 (N_6605,N_1785,N_3217);
nand U6606 (N_6606,N_4928,N_4291);
nor U6607 (N_6607,N_107,N_1903);
and U6608 (N_6608,N_2800,N_791);
nand U6609 (N_6609,N_245,N_3244);
or U6610 (N_6610,N_4574,N_2396);
or U6611 (N_6611,N_2411,N_2667);
nand U6612 (N_6612,N_4025,N_4532);
or U6613 (N_6613,N_2224,N_4075);
nor U6614 (N_6614,N_895,N_4374);
xor U6615 (N_6615,N_1401,N_371);
or U6616 (N_6616,N_1582,N_3103);
nand U6617 (N_6617,N_4173,N_1577);
or U6618 (N_6618,N_1301,N_601);
nor U6619 (N_6619,N_769,N_3126);
or U6620 (N_6620,N_453,N_1729);
and U6621 (N_6621,N_4692,N_3811);
xnor U6622 (N_6622,N_4269,N_324);
or U6623 (N_6623,N_1832,N_2766);
or U6624 (N_6624,N_390,N_2932);
and U6625 (N_6625,N_123,N_4644);
and U6626 (N_6626,N_3540,N_1530);
and U6627 (N_6627,N_61,N_1148);
or U6628 (N_6628,N_4217,N_2496);
xnor U6629 (N_6629,N_1610,N_3821);
and U6630 (N_6630,N_3165,N_2886);
nor U6631 (N_6631,N_2342,N_1470);
or U6632 (N_6632,N_4806,N_4219);
xor U6633 (N_6633,N_1836,N_855);
and U6634 (N_6634,N_2760,N_1887);
and U6635 (N_6635,N_2366,N_3974);
and U6636 (N_6636,N_585,N_4939);
and U6637 (N_6637,N_2948,N_2731);
xnor U6638 (N_6638,N_4641,N_1641);
xnor U6639 (N_6639,N_2768,N_1141);
xnor U6640 (N_6640,N_4375,N_2276);
and U6641 (N_6641,N_2937,N_672);
or U6642 (N_6642,N_4784,N_1687);
or U6643 (N_6643,N_3738,N_612);
nand U6644 (N_6644,N_3131,N_2533);
or U6645 (N_6645,N_4661,N_4745);
xor U6646 (N_6646,N_4213,N_3154);
or U6647 (N_6647,N_3649,N_3151);
and U6648 (N_6648,N_4655,N_418);
xor U6649 (N_6649,N_3542,N_774);
nor U6650 (N_6650,N_2644,N_4682);
nor U6651 (N_6651,N_3252,N_2748);
or U6652 (N_6652,N_3632,N_2891);
xor U6653 (N_6653,N_2232,N_1019);
nand U6654 (N_6654,N_4459,N_1484);
nor U6655 (N_6655,N_3657,N_236);
nor U6656 (N_6656,N_3840,N_4885);
nor U6657 (N_6657,N_405,N_4726);
xnor U6658 (N_6658,N_1560,N_4133);
or U6659 (N_6659,N_1765,N_83);
or U6660 (N_6660,N_990,N_312);
nor U6661 (N_6661,N_3180,N_3977);
nor U6662 (N_6662,N_1070,N_380);
xor U6663 (N_6663,N_3670,N_149);
nand U6664 (N_6664,N_1980,N_953);
xor U6665 (N_6665,N_1615,N_488);
or U6666 (N_6666,N_4281,N_4656);
nand U6667 (N_6667,N_3348,N_4556);
nand U6668 (N_6668,N_1498,N_4513);
and U6669 (N_6669,N_183,N_1640);
nand U6670 (N_6670,N_2317,N_2925);
nand U6671 (N_6671,N_561,N_1184);
and U6672 (N_6672,N_3869,N_3159);
or U6673 (N_6673,N_3939,N_4801);
nand U6674 (N_6674,N_2538,N_2934);
nand U6675 (N_6675,N_2484,N_1534);
or U6676 (N_6676,N_4567,N_3535);
and U6677 (N_6677,N_394,N_4600);
nor U6678 (N_6678,N_3423,N_4226);
xnor U6679 (N_6679,N_830,N_3871);
xnor U6680 (N_6680,N_2955,N_3641);
nor U6681 (N_6681,N_3467,N_945);
and U6682 (N_6682,N_2492,N_4838);
xor U6683 (N_6683,N_4413,N_4587);
and U6684 (N_6684,N_1407,N_2114);
xor U6685 (N_6685,N_2626,N_104);
nand U6686 (N_6686,N_1895,N_478);
nand U6687 (N_6687,N_2779,N_1367);
or U6688 (N_6688,N_2259,N_1629);
and U6689 (N_6689,N_94,N_3579);
nand U6690 (N_6690,N_263,N_4578);
xor U6691 (N_6691,N_225,N_1829);
and U6692 (N_6692,N_3066,N_2086);
or U6693 (N_6693,N_67,N_2935);
nand U6694 (N_6694,N_3765,N_797);
and U6695 (N_6695,N_4024,N_3714);
xor U6696 (N_6696,N_4679,N_4081);
xnor U6697 (N_6697,N_3442,N_1423);
nand U6698 (N_6698,N_244,N_512);
nand U6699 (N_6699,N_3200,N_161);
and U6700 (N_6700,N_3278,N_326);
xnor U6701 (N_6701,N_4071,N_2941);
and U6702 (N_6702,N_2286,N_4104);
xnor U6703 (N_6703,N_4096,N_2654);
xnor U6704 (N_6704,N_1381,N_3344);
nor U6705 (N_6705,N_314,N_2875);
nand U6706 (N_6706,N_4430,N_4068);
nor U6707 (N_6707,N_4445,N_2456);
nor U6708 (N_6708,N_220,N_4047);
nand U6709 (N_6709,N_2252,N_1848);
or U6710 (N_6710,N_1870,N_2801);
xor U6711 (N_6711,N_3004,N_2716);
nor U6712 (N_6712,N_584,N_3253);
xor U6713 (N_6713,N_3043,N_4449);
xnor U6714 (N_6714,N_4054,N_3110);
and U6715 (N_6715,N_3424,N_109);
and U6716 (N_6716,N_3376,N_2849);
and U6717 (N_6717,N_3081,N_2953);
or U6718 (N_6718,N_42,N_2534);
or U6719 (N_6719,N_4408,N_166);
and U6720 (N_6720,N_489,N_1404);
or U6721 (N_6721,N_4921,N_1124);
xnor U6722 (N_6722,N_4538,N_2835);
nand U6723 (N_6723,N_3807,N_134);
nor U6724 (N_6724,N_2887,N_3748);
and U6725 (N_6725,N_4423,N_4409);
nand U6726 (N_6726,N_3525,N_3938);
nand U6727 (N_6727,N_701,N_3438);
and U6728 (N_6728,N_4035,N_4469);
nand U6729 (N_6729,N_1436,N_4800);
xnor U6730 (N_6730,N_1952,N_336);
xor U6731 (N_6731,N_2576,N_2593);
nand U6732 (N_6732,N_861,N_2742);
and U6733 (N_6733,N_3686,N_2680);
nand U6734 (N_6734,N_3788,N_4120);
nand U6735 (N_6735,N_4369,N_1012);
or U6736 (N_6736,N_292,N_4018);
and U6737 (N_6737,N_4755,N_2078);
xnor U6738 (N_6738,N_3935,N_3502);
and U6739 (N_6739,N_3567,N_4221);
or U6740 (N_6740,N_4757,N_1090);
nand U6741 (N_6741,N_1378,N_1121);
and U6742 (N_6742,N_18,N_2614);
xor U6743 (N_6743,N_4767,N_4614);
or U6744 (N_6744,N_364,N_1957);
nand U6745 (N_6745,N_1072,N_591);
nor U6746 (N_6746,N_2334,N_3619);
nor U6747 (N_6747,N_2458,N_357);
and U6748 (N_6748,N_4633,N_2814);
or U6749 (N_6749,N_4903,N_647);
or U6750 (N_6750,N_4946,N_1794);
and U6751 (N_6751,N_2897,N_3675);
nor U6752 (N_6752,N_1294,N_682);
and U6753 (N_6753,N_4187,N_724);
nand U6754 (N_6754,N_3335,N_4970);
or U6755 (N_6755,N_749,N_3298);
and U6756 (N_6756,N_805,N_152);
and U6757 (N_6757,N_2623,N_2575);
nor U6758 (N_6758,N_1506,N_1821);
and U6759 (N_6759,N_625,N_933);
xor U6760 (N_6760,N_3705,N_365);
or U6761 (N_6761,N_3629,N_3269);
xnor U6762 (N_6762,N_4174,N_2414);
nand U6763 (N_6763,N_3732,N_3615);
or U6764 (N_6764,N_765,N_2050);
nand U6765 (N_6765,N_1883,N_1988);
nand U6766 (N_6766,N_1337,N_2880);
xor U6767 (N_6767,N_3089,N_2990);
nand U6768 (N_6768,N_4676,N_1299);
nor U6769 (N_6769,N_4607,N_518);
nor U6770 (N_6770,N_1435,N_1973);
nor U6771 (N_6771,N_4401,N_1881);
or U6772 (N_6772,N_1517,N_2103);
nand U6773 (N_6773,N_806,N_3707);
or U6774 (N_6774,N_3002,N_650);
and U6775 (N_6775,N_66,N_428);
or U6776 (N_6776,N_2145,N_1034);
or U6777 (N_6777,N_927,N_3665);
nor U6778 (N_6778,N_22,N_1897);
xnor U6779 (N_6779,N_1298,N_86);
nand U6780 (N_6780,N_399,N_3636);
and U6781 (N_6781,N_4351,N_1522);
xnor U6782 (N_6782,N_623,N_218);
and U6783 (N_6783,N_1112,N_4402);
and U6784 (N_6784,N_2940,N_4487);
nor U6785 (N_6785,N_542,N_256);
and U6786 (N_6786,N_3185,N_1553);
xnor U6787 (N_6787,N_3237,N_4016);
xnor U6788 (N_6788,N_3488,N_449);
and U6789 (N_6789,N_1174,N_157);
nand U6790 (N_6790,N_47,N_4448);
nand U6791 (N_6791,N_1488,N_4178);
xor U6792 (N_6792,N_3519,N_176);
or U6793 (N_6793,N_1673,N_1311);
xnor U6794 (N_6794,N_2101,N_359);
nand U6795 (N_6795,N_2447,N_4472);
or U6796 (N_6796,N_4823,N_2500);
and U6797 (N_6797,N_4076,N_833);
xnor U6798 (N_6798,N_1021,N_4701);
or U6799 (N_6799,N_541,N_2491);
nand U6800 (N_6800,N_117,N_2004);
nor U6801 (N_6801,N_576,N_2966);
nand U6802 (N_6802,N_1592,N_3368);
nand U6803 (N_6803,N_2901,N_1538);
and U6804 (N_6804,N_3605,N_4207);
xor U6805 (N_6805,N_4896,N_3420);
and U6806 (N_6806,N_4454,N_4672);
or U6807 (N_6807,N_886,N_285);
xor U6808 (N_6808,N_4868,N_3933);
nor U6809 (N_6809,N_1627,N_1666);
nor U6810 (N_6810,N_1616,N_4094);
nand U6811 (N_6811,N_2720,N_95);
and U6812 (N_6812,N_992,N_2212);
and U6813 (N_6813,N_925,N_2108);
nor U6814 (N_6814,N_3861,N_2339);
and U6815 (N_6815,N_3263,N_4778);
and U6816 (N_6816,N_214,N_2110);
xor U6817 (N_6817,N_922,N_829);
xor U6818 (N_6818,N_802,N_3101);
and U6819 (N_6819,N_4255,N_4007);
nand U6820 (N_6820,N_4544,N_2621);
nand U6821 (N_6821,N_3945,N_4460);
and U6822 (N_6822,N_1715,N_3832);
nand U6823 (N_6823,N_3893,N_3577);
and U6824 (N_6824,N_4287,N_2715);
nor U6825 (N_6825,N_3220,N_4700);
xor U6826 (N_6826,N_1915,N_4794);
nor U6827 (N_6827,N_764,N_1208);
xnor U6828 (N_6828,N_3596,N_2270);
or U6829 (N_6829,N_116,N_877);
or U6830 (N_6830,N_2450,N_4359);
or U6831 (N_6831,N_1003,N_548);
nand U6832 (N_6832,N_2156,N_2743);
nand U6833 (N_6833,N_3040,N_618);
nor U6834 (N_6834,N_4640,N_4331);
nor U6835 (N_6835,N_2888,N_4443);
nor U6836 (N_6836,N_4780,N_3528);
nor U6837 (N_6837,N_3833,N_3296);
nand U6838 (N_6838,N_2066,N_746);
xnor U6839 (N_6839,N_158,N_4416);
or U6840 (N_6840,N_2699,N_1801);
nand U6841 (N_6841,N_2225,N_306);
or U6842 (N_6842,N_556,N_3036);
and U6843 (N_6843,N_1181,N_2665);
xnor U6844 (N_6844,N_248,N_3114);
xor U6845 (N_6845,N_3911,N_2884);
and U6846 (N_6846,N_3359,N_1835);
or U6847 (N_6847,N_3060,N_422);
xor U6848 (N_6848,N_3745,N_3210);
or U6849 (N_6849,N_871,N_1983);
nand U6850 (N_6850,N_1601,N_2395);
and U6851 (N_6851,N_1215,N_2499);
nor U6852 (N_6852,N_1591,N_4099);
or U6853 (N_6853,N_3268,N_4666);
nand U6854 (N_6854,N_3443,N_4437);
xor U6855 (N_6855,N_3741,N_164);
nor U6856 (N_6856,N_4241,N_897);
xnor U6857 (N_6857,N_3346,N_1816);
nand U6858 (N_6858,N_1146,N_229);
and U6859 (N_6859,N_4008,N_2350);
nand U6860 (N_6860,N_4673,N_3451);
or U6861 (N_6861,N_3895,N_1032);
or U6862 (N_6862,N_3021,N_141);
nand U6863 (N_6863,N_4055,N_169);
nor U6864 (N_6864,N_2710,N_2813);
nand U6865 (N_6865,N_4982,N_2686);
and U6866 (N_6866,N_173,N_906);
and U6867 (N_6867,N_497,N_36);
nor U6868 (N_6868,N_4751,N_989);
nor U6869 (N_6869,N_4855,N_1200);
xor U6870 (N_6870,N_507,N_4727);
and U6871 (N_6871,N_1938,N_4180);
and U6872 (N_6872,N_3454,N_3804);
nor U6873 (N_6873,N_3980,N_2494);
xor U6874 (N_6874,N_2245,N_4579);
xor U6875 (N_6875,N_3793,N_3981);
or U6876 (N_6876,N_2869,N_2682);
xor U6877 (N_6877,N_2095,N_1270);
nor U6878 (N_6878,N_1230,N_1452);
xor U6879 (N_6879,N_652,N_4704);
nand U6880 (N_6880,N_1216,N_4276);
nor U6881 (N_6881,N_3882,N_3718);
nor U6882 (N_6882,N_3499,N_435);
xnor U6883 (N_6883,N_2002,N_1276);
nand U6884 (N_6884,N_1844,N_1413);
nor U6885 (N_6885,N_2126,N_2226);
or U6886 (N_6886,N_2107,N_2769);
nand U6887 (N_6887,N_271,N_1934);
and U6888 (N_6888,N_4638,N_834);
nor U6889 (N_6889,N_3473,N_2360);
or U6890 (N_6890,N_846,N_3045);
nand U6891 (N_6891,N_849,N_1227);
and U6892 (N_6892,N_1657,N_2168);
nand U6893 (N_6893,N_3127,N_432);
and U6894 (N_6894,N_929,N_4347);
or U6895 (N_6895,N_3982,N_2646);
or U6896 (N_6896,N_4937,N_3616);
nand U6897 (N_6897,N_304,N_3758);
nor U6898 (N_6898,N_2662,N_660);
nor U6899 (N_6899,N_2902,N_3569);
nor U6900 (N_6900,N_4702,N_112);
nand U6901 (N_6901,N_2591,N_4846);
nand U6902 (N_6902,N_4313,N_3626);
or U6903 (N_6903,N_3071,N_3796);
or U6904 (N_6904,N_93,N_3521);
nand U6905 (N_6905,N_3482,N_275);
xor U6906 (N_6906,N_1742,N_2115);
and U6907 (N_6907,N_3724,N_3342);
nor U6908 (N_6908,N_2564,N_3398);
nand U6909 (N_6909,N_1721,N_4514);
nand U6910 (N_6910,N_1099,N_2333);
and U6911 (N_6911,N_2173,N_579);
or U6912 (N_6912,N_3783,N_15);
xor U6913 (N_6913,N_75,N_4753);
nor U6914 (N_6914,N_4858,N_1723);
or U6915 (N_6915,N_2628,N_1471);
xor U6916 (N_6916,N_4957,N_3517);
xnor U6917 (N_6917,N_3894,N_3090);
nor U6918 (N_6918,N_58,N_1660);
or U6919 (N_6919,N_2727,N_1847);
nor U6920 (N_6920,N_4135,N_2279);
xnor U6921 (N_6921,N_3357,N_3760);
and U6922 (N_6922,N_2649,N_3480);
nor U6923 (N_6923,N_1155,N_2736);
nand U6924 (N_6924,N_1086,N_188);
nand U6925 (N_6925,N_589,N_3896);
or U6926 (N_6926,N_3328,N_3175);
nor U6927 (N_6927,N_3773,N_13);
and U6928 (N_6928,N_565,N_228);
or U6929 (N_6929,N_758,N_2374);
nand U6930 (N_6930,N_2012,N_2636);
xnor U6931 (N_6931,N_2452,N_3961);
nand U6932 (N_6932,N_532,N_73);
or U6933 (N_6933,N_2249,N_480);
or U6934 (N_6934,N_609,N_2429);
or U6935 (N_6935,N_4159,N_339);
and U6936 (N_6936,N_4793,N_3827);
nand U6937 (N_6937,N_1901,N_4074);
or U6938 (N_6938,N_4772,N_462);
and U6939 (N_6939,N_2829,N_151);
or U6940 (N_6940,N_2467,N_790);
nor U6941 (N_6941,N_1747,N_4689);
or U6942 (N_6942,N_4141,N_3096);
or U6943 (N_6943,N_1083,N_4333);
nor U6944 (N_6944,N_3163,N_2541);
and U6945 (N_6945,N_1328,N_207);
or U6946 (N_6946,N_763,N_1986);
xnor U6947 (N_6947,N_2336,N_1265);
or U6948 (N_6948,N_2969,N_3549);
nor U6949 (N_6949,N_1122,N_7);
nor U6950 (N_6950,N_1830,N_3565);
nand U6951 (N_6951,N_1689,N_1385);
nand U6952 (N_6952,N_818,N_1290);
nand U6953 (N_6953,N_261,N_2229);
nor U6954 (N_6954,N_2648,N_3889);
and U6955 (N_6955,N_1789,N_65);
nor U6956 (N_6956,N_2927,N_690);
nand U6957 (N_6957,N_2583,N_4483);
xor U6958 (N_6958,N_4817,N_2400);
or U6959 (N_6959,N_2158,N_3387);
or U6960 (N_6960,N_3343,N_694);
and U6961 (N_6961,N_4132,N_3468);
or U6962 (N_6962,N_4736,N_1686);
xnor U6963 (N_6963,N_235,N_4095);
nand U6964 (N_6964,N_2061,N_4545);
and U6965 (N_6965,N_4036,N_1865);
or U6966 (N_6966,N_2437,N_4721);
or U6967 (N_6967,N_4887,N_3912);
xnor U6968 (N_6968,N_1293,N_1081);
and U6969 (N_6969,N_852,N_2302);
and U6970 (N_6970,N_3643,N_4847);
and U6971 (N_6971,N_21,N_2820);
and U6972 (N_6972,N_3267,N_705);
nor U6973 (N_6973,N_1586,N_4458);
nand U6974 (N_6974,N_982,N_2994);
or U6975 (N_6975,N_4723,N_451);
nor U6976 (N_6976,N_4379,N_2918);
and U6977 (N_6977,N_3248,N_645);
xnor U6978 (N_6978,N_2372,N_963);
xnor U6979 (N_6979,N_215,N_2681);
and U6980 (N_6980,N_3065,N_3061);
nand U6981 (N_6981,N_4512,N_3005);
and U6982 (N_6982,N_3510,N_4999);
xnor U6983 (N_6983,N_2077,N_3138);
and U6984 (N_6984,N_2448,N_4705);
or U6985 (N_6985,N_2842,N_3970);
xor U6986 (N_6986,N_2355,N_1210);
or U6987 (N_6987,N_1556,N_2655);
nor U6988 (N_6988,N_4737,N_3966);
and U6989 (N_6989,N_838,N_872);
and U6990 (N_6990,N_1160,N_363);
xor U6991 (N_6991,N_1841,N_2316);
and U6992 (N_6992,N_4878,N_3351);
xor U6993 (N_6993,N_3429,N_4003);
and U6994 (N_6994,N_1562,N_3393);
nor U6995 (N_6995,N_55,N_782);
xnor U6996 (N_6996,N_1933,N_4583);
nor U6997 (N_6997,N_3085,N_377);
nand U6998 (N_6998,N_3173,N_4211);
or U6999 (N_6999,N_2803,N_1677);
nand U7000 (N_7000,N_3680,N_3815);
nand U7001 (N_7001,N_2922,N_33);
and U7002 (N_7002,N_1472,N_2175);
nor U7003 (N_7003,N_37,N_717);
and U7004 (N_7004,N_3522,N_1879);
nor U7005 (N_7005,N_484,N_642);
nand U7006 (N_7006,N_3049,N_3111);
nand U7007 (N_7007,N_1919,N_4051);
xnor U7008 (N_7008,N_1775,N_62);
or U7009 (N_7009,N_4561,N_4533);
or U7010 (N_7010,N_3259,N_1815);
nand U7011 (N_7011,N_1199,N_3137);
nand U7012 (N_7012,N_2696,N_594);
and U7013 (N_7013,N_3725,N_1354);
nand U7014 (N_7014,N_1764,N_3997);
nor U7015 (N_7015,N_4168,N_4943);
or U7016 (N_7016,N_1568,N_1400);
and U7017 (N_7017,N_3284,N_3721);
nor U7018 (N_7018,N_3609,N_1909);
nor U7019 (N_7019,N_801,N_1526);
nor U7020 (N_7020,N_4012,N_767);
nand U7021 (N_7021,N_4605,N_757);
xnor U7022 (N_7022,N_3733,N_3205);
and U7023 (N_7023,N_4185,N_2);
xor U7024 (N_7024,N_165,N_1575);
xnor U7025 (N_7025,N_4317,N_3978);
nor U7026 (N_7026,N_355,N_1100);
or U7027 (N_7027,N_815,N_4302);
and U7028 (N_7028,N_2738,N_3152);
xor U7029 (N_7029,N_4290,N_2446);
xnor U7030 (N_7030,N_1169,N_4949);
nand U7031 (N_7031,N_4872,N_2047);
and U7032 (N_7032,N_4831,N_715);
xor U7033 (N_7033,N_1714,N_1310);
and U7034 (N_7034,N_1991,N_3599);
and U7035 (N_7035,N_4111,N_1030);
nand U7036 (N_7036,N_574,N_4754);
and U7037 (N_7037,N_3450,N_338);
nand U7038 (N_7038,N_2865,N_2698);
and U7039 (N_7039,N_197,N_2141);
nand U7040 (N_7040,N_4466,N_3315);
or U7041 (N_7041,N_3246,N_2836);
xnor U7042 (N_7042,N_1263,N_3199);
xnor U7043 (N_7043,N_4451,N_1576);
nand U7044 (N_7044,N_3093,N_472);
and U7045 (N_7045,N_4041,N_938);
xnor U7046 (N_7046,N_2373,N_3025);
or U7047 (N_7047,N_2910,N_4955);
and U7048 (N_7048,N_555,N_2838);
or U7049 (N_7049,N_3226,N_4732);
xnor U7050 (N_7050,N_3477,N_2010);
nor U7051 (N_7051,N_943,N_1974);
and U7052 (N_7052,N_3392,N_2519);
and U7053 (N_7053,N_1132,N_4923);
nor U7054 (N_7054,N_2936,N_4586);
nand U7055 (N_7055,N_4190,N_1411);
nor U7056 (N_7056,N_4345,N_3057);
xnor U7057 (N_7057,N_627,N_4419);
xor U7058 (N_7058,N_4170,N_4440);
and U7059 (N_7059,N_260,N_4934);
or U7060 (N_7060,N_4916,N_712);
or U7061 (N_7061,N_2755,N_106);
nand U7062 (N_7062,N_2610,N_409);
or U7063 (N_7063,N_140,N_4575);
nand U7064 (N_7064,N_665,N_1029);
nor U7065 (N_7065,N_3753,N_4328);
and U7066 (N_7066,N_1520,N_2775);
nand U7067 (N_7067,N_2233,N_1911);
and U7068 (N_7068,N_2762,N_1813);
and U7069 (N_7069,N_4216,N_397);
nor U7070 (N_7070,N_2271,N_2707);
nor U7071 (N_7071,N_3006,N_3475);
nor U7072 (N_7072,N_3439,N_233);
nor U7073 (N_7073,N_4619,N_1691);
and U7074 (N_7074,N_4919,N_162);
nand U7075 (N_7075,N_4332,N_2562);
and U7076 (N_7076,N_529,N_2123);
nor U7077 (N_7077,N_1922,N_322);
nor U7078 (N_7078,N_4973,N_2451);
nand U7079 (N_7079,N_2714,N_4365);
nor U7080 (N_7080,N_4079,N_3211);
or U7081 (N_7081,N_2624,N_2297);
and U7082 (N_7082,N_4117,N_1136);
nand U7083 (N_7083,N_4808,N_731);
nand U7084 (N_7084,N_517,N_3988);
nand U7085 (N_7085,N_2323,N_4888);
nor U7086 (N_7086,N_2119,N_2326);
xnor U7087 (N_7087,N_3801,N_1824);
nand U7088 (N_7088,N_1783,N_772);
nor U7089 (N_7089,N_402,N_2335);
and U7090 (N_7090,N_2483,N_2380);
nor U7091 (N_7091,N_4383,N_2771);
or U7092 (N_7092,N_3353,N_4023);
or U7093 (N_7093,N_3476,N_2585);
or U7094 (N_7094,N_4182,N_4537);
nor U7095 (N_7095,N_4435,N_3115);
nor U7096 (N_7096,N_3936,N_1226);
nor U7097 (N_7097,N_4485,N_3784);
or U7098 (N_7098,N_3902,N_35);
nand U7099 (N_7099,N_2290,N_3456);
nor U7100 (N_7100,N_3573,N_2369);
nand U7101 (N_7101,N_3361,N_4154);
xnor U7102 (N_7102,N_3696,N_1838);
xor U7103 (N_7103,N_2784,N_3142);
nor U7104 (N_7104,N_4486,N_4573);
or U7105 (N_7105,N_281,N_3326);
nand U7106 (N_7106,N_1426,N_908);
and U7107 (N_7107,N_2733,N_2993);
nor U7108 (N_7108,N_4059,N_4891);
xor U7109 (N_7109,N_958,N_4109);
nor U7110 (N_7110,N_1285,N_4526);
nand U7111 (N_7111,N_3909,N_4284);
nand U7112 (N_7112,N_875,N_1732);
or U7113 (N_7113,N_3254,N_3421);
xor U7114 (N_7114,N_1818,N_262);
or U7115 (N_7115,N_3582,N_1950);
or U7116 (N_7116,N_2085,N_427);
nor U7117 (N_7117,N_208,N_56);
nor U7118 (N_7118,N_3290,N_1886);
or U7119 (N_7119,N_4001,N_2809);
and U7120 (N_7120,N_530,N_2971);
xnor U7121 (N_7121,N_4208,N_554);
nor U7122 (N_7122,N_72,N_3417);
and U7123 (N_7123,N_753,N_1454);
nor U7124 (N_7124,N_3212,N_2038);
nor U7125 (N_7125,N_2284,N_2961);
nor U7126 (N_7126,N_3877,N_859);
or U7127 (N_7127,N_3202,N_4901);
nor U7128 (N_7128,N_1863,N_3654);
and U7129 (N_7129,N_1544,N_2634);
and U7130 (N_7130,N_4964,N_1920);
nor U7131 (N_7131,N_4987,N_137);
nand U7132 (N_7132,N_4802,N_1561);
nand U7133 (N_7133,N_2404,N_3953);
xor U7134 (N_7134,N_4473,N_915);
and U7135 (N_7135,N_4070,N_3655);
nand U7136 (N_7136,N_4040,N_3532);
nand U7137 (N_7137,N_3512,N_3529);
nor U7138 (N_7138,N_1362,N_788);
nand U7139 (N_7139,N_3186,N_2041);
nand U7140 (N_7140,N_3017,N_374);
or U7141 (N_7141,N_3515,N_2329);
nand U7142 (N_7142,N_2176,N_3672);
or U7143 (N_7143,N_4825,N_1837);
xnor U7144 (N_7144,N_2999,N_4444);
or U7145 (N_7145,N_760,N_559);
xor U7146 (N_7146,N_1364,N_1071);
or U7147 (N_7147,N_4687,N_1539);
and U7148 (N_7148,N_2013,N_2566);
xor U7149 (N_7149,N_4910,N_2438);
xnor U7150 (N_7150,N_2504,N_2923);
or U7151 (N_7151,N_3399,N_966);
nand U7152 (N_7152,N_1453,N_4667);
and U7153 (N_7153,N_2919,N_2253);
or U7154 (N_7154,N_2343,N_4357);
xnor U7155 (N_7155,N_1418,N_792);
nor U7156 (N_7156,N_3608,N_3546);
and U7157 (N_7157,N_1661,N_2663);
nand U7158 (N_7158,N_4908,N_1941);
nand U7159 (N_7159,N_1690,N_1190);
nand U7160 (N_7160,N_4235,N_1579);
and U7161 (N_7161,N_700,N_3272);
nor U7162 (N_7162,N_2093,N_2782);
nand U7163 (N_7163,N_1358,N_4418);
nor U7164 (N_7164,N_4630,N_2073);
and U7165 (N_7165,N_486,N_209);
or U7166 (N_7166,N_689,N_1307);
xnor U7167 (N_7167,N_4834,N_27);
or U7168 (N_7168,N_4634,N_3598);
nor U7169 (N_7169,N_3593,N_1281);
and U7170 (N_7170,N_2140,N_4536);
nand U7171 (N_7171,N_2889,N_1978);
or U7172 (N_7172,N_391,N_3059);
or U7173 (N_7173,N_2823,N_832);
or U7174 (N_7174,N_498,N_1254);
nor U7175 (N_7175,N_843,N_240);
xor U7176 (N_7176,N_876,N_2283);
xor U7177 (N_7177,N_2243,N_3710);
or U7178 (N_7178,N_1767,N_4199);
nor U7179 (N_7179,N_3597,N_16);
nand U7180 (N_7180,N_4774,N_3639);
or U7181 (N_7181,N_2493,N_2810);
nor U7182 (N_7182,N_3038,N_3819);
nand U7183 (N_7183,N_3559,N_3020);
nor U7184 (N_7184,N_38,N_297);
nand U7185 (N_7185,N_3448,N_913);
nand U7186 (N_7186,N_4434,N_2607);
and U7187 (N_7187,N_3107,N_4388);
and U7188 (N_7188,N_4860,N_3316);
or U7189 (N_7189,N_2708,N_1398);
and U7190 (N_7190,N_3723,N_2125);
nand U7191 (N_7191,N_3538,N_4739);
nand U7192 (N_7192,N_4597,N_1059);
and U7193 (N_7193,N_4198,N_4945);
nand U7194 (N_7194,N_1864,N_2512);
and U7195 (N_7195,N_3416,N_1282);
nor U7196 (N_7196,N_714,N_150);
and U7197 (N_7197,N_1312,N_1001);
nand U7198 (N_7198,N_3589,N_2394);
nand U7199 (N_7199,N_1868,N_2135);
and U7200 (N_7200,N_3441,N_4229);
xnor U7201 (N_7201,N_3996,N_348);
or U7202 (N_7202,N_4977,N_3892);
nand U7203 (N_7203,N_308,N_217);
nand U7204 (N_7204,N_4032,N_4162);
or U7205 (N_7205,N_4385,N_2563);
xnor U7206 (N_7206,N_890,N_4194);
xor U7207 (N_7207,N_202,N_3874);
or U7208 (N_7208,N_3886,N_4061);
or U7209 (N_7209,N_1809,N_1133);
nor U7210 (N_7210,N_1262,N_816);
nor U7211 (N_7211,N_3275,N_3340);
and U7212 (N_7212,N_2879,N_1011);
nor U7213 (N_7213,N_920,N_4799);
nor U7214 (N_7214,N_727,N_1461);
nand U7215 (N_7215,N_2589,N_1845);
or U7216 (N_7216,N_2390,N_1755);
and U7217 (N_7217,N_3526,N_3867);
nor U7218 (N_7218,N_2658,N_2381);
nor U7219 (N_7219,N_1987,N_40);
and U7220 (N_7220,N_4843,N_793);
xnor U7221 (N_7221,N_4553,N_3539);
nand U7222 (N_7222,N_1359,N_2059);
nand U7223 (N_7223,N_1557,N_4952);
nand U7224 (N_7224,N_2627,N_4050);
nor U7225 (N_7225,N_411,N_2327);
nand U7226 (N_7226,N_926,N_4210);
xnor U7227 (N_7227,N_680,N_1510);
nor U7228 (N_7228,N_1170,N_3490);
nand U7229 (N_7229,N_2352,N_560);
nor U7230 (N_7230,N_3663,N_2312);
xor U7231 (N_7231,N_2509,N_4441);
and U7232 (N_7232,N_1959,N_2139);
or U7233 (N_7233,N_4603,N_1434);
nand U7234 (N_7234,N_3720,N_898);
xnor U7235 (N_7235,N_122,N_1704);
nand U7236 (N_7236,N_1186,N_4303);
and U7237 (N_7237,N_1189,N_1244);
or U7238 (N_7238,N_1065,N_4992);
xor U7239 (N_7239,N_3942,N_2669);
nor U7240 (N_7240,N_1278,N_893);
nand U7241 (N_7241,N_2802,N_333);
xnor U7242 (N_7242,N_4805,N_515);
nor U7243 (N_7243,N_3677,N_2578);
nand U7244 (N_7244,N_981,N_78);
nor U7245 (N_7245,N_3239,N_3562);
nor U7246 (N_7246,N_4350,N_3962);
nand U7247 (N_7247,N_1211,N_997);
nor U7248 (N_7248,N_1831,N_1999);
or U7249 (N_7249,N_2382,N_4373);
xnor U7250 (N_7250,N_3693,N_1192);
or U7251 (N_7251,N_3578,N_1480);
or U7252 (N_7252,N_4399,N_535);
nor U7253 (N_7253,N_2461,N_4625);
nor U7254 (N_7254,N_3627,N_4356);
nor U7255 (N_7255,N_3000,N_4286);
nor U7256 (N_7256,N_3779,N_2571);
nor U7257 (N_7257,N_4811,N_521);
nand U7258 (N_7258,N_3086,N_278);
and U7259 (N_7259,N_1990,N_2946);
xor U7260 (N_7260,N_3030,N_4958);
or U7261 (N_7261,N_4558,N_3814);
or U7262 (N_7262,N_655,N_4482);
xor U7263 (N_7263,N_1600,N_2081);
nor U7264 (N_7264,N_3614,N_204);
nand U7265 (N_7265,N_1710,N_836);
and U7266 (N_7266,N_1515,N_651);
or U7267 (N_7267,N_1234,N_119);
nand U7268 (N_7268,N_3715,N_2008);
or U7269 (N_7269,N_174,N_200);
xnor U7270 (N_7270,N_4642,N_2620);
nand U7271 (N_7271,N_3635,N_1979);
or U7272 (N_7272,N_1035,N_3791);
or U7273 (N_7273,N_1754,N_3949);
and U7274 (N_7274,N_2683,N_1458);
and U7275 (N_7275,N_1702,N_4539);
nor U7276 (N_7276,N_1851,N_1248);
xnor U7277 (N_7277,N_3660,N_563);
or U7278 (N_7278,N_98,N_2147);
or U7279 (N_7279,N_2029,N_779);
or U7280 (N_7280,N_687,N_2825);
nor U7281 (N_7281,N_417,N_3400);
nor U7282 (N_7282,N_3331,N_4708);
xor U7283 (N_7283,N_1153,N_3397);
and U7284 (N_7284,N_289,N_2739);
nor U7285 (N_7285,N_3799,N_883);
nor U7286 (N_7286,N_1403,N_2067);
nand U7287 (N_7287,N_2349,N_3001);
xor U7288 (N_7288,N_636,N_2261);
nor U7289 (N_7289,N_2905,N_3946);
and U7290 (N_7290,N_1807,N_756);
and U7291 (N_7291,N_570,N_434);
or U7292 (N_7292,N_2223,N_646);
xor U7293 (N_7293,N_1102,N_4488);
nand U7294 (N_7294,N_3265,N_2647);
or U7295 (N_7295,N_3772,N_2903);
and U7296 (N_7296,N_1817,N_3560);
nor U7297 (N_7297,N_342,N_1391);
and U7298 (N_7298,N_2215,N_1372);
or U7299 (N_7299,N_4176,N_577);
nand U7300 (N_7300,N_4670,N_4015);
or U7301 (N_7301,N_1880,N_604);
and U7302 (N_7302,N_3113,N_2863);
nor U7303 (N_7303,N_3027,N_1005);
and U7304 (N_7304,N_1236,N_4467);
and U7305 (N_7305,N_69,N_1749);
nand U7306 (N_7306,N_1523,N_595);
nand U7307 (N_7307,N_2068,N_2082);
and U7308 (N_7308,N_4913,N_2673);
and U7309 (N_7309,N_510,N_1552);
xnor U7310 (N_7310,N_238,N_3802);
xnor U7311 (N_7311,N_1740,N_3097);
xnor U7312 (N_7312,N_4562,N_1779);
xnor U7313 (N_7313,N_2376,N_1855);
xor U7314 (N_7314,N_4624,N_3305);
or U7315 (N_7315,N_2526,N_4950);
nand U7316 (N_7316,N_2202,N_1329);
xnor U7317 (N_7317,N_1802,N_3994);
xor U7318 (N_7318,N_4529,N_1977);
nor U7319 (N_7319,N_850,N_3308);
nor U7320 (N_7320,N_1068,N_3028);
xor U7321 (N_7321,N_2408,N_4765);
and U7322 (N_7322,N_2645,N_1548);
or U7323 (N_7323,N_762,N_4959);
xor U7324 (N_7324,N_3591,N_2749);
nor U7325 (N_7325,N_4062,N_3918);
xor U7326 (N_7326,N_3662,N_138);
xnor U7327 (N_7327,N_1888,N_1894);
xor U7328 (N_7328,N_4101,N_1127);
nor U7329 (N_7329,N_25,N_2440);
or U7330 (N_7330,N_754,N_1955);
or U7331 (N_7331,N_4974,N_3746);
nor U7332 (N_7332,N_643,N_446);
nand U7333 (N_7333,N_4849,N_3806);
or U7334 (N_7334,N_2943,N_132);
nand U7335 (N_7335,N_1780,N_3167);
xnor U7336 (N_7336,N_4535,N_1256);
nor U7337 (N_7337,N_2267,N_4230);
nor U7338 (N_7338,N_4942,N_1499);
nand U7339 (N_7339,N_624,N_3633);
and U7340 (N_7340,N_3762,N_4029);
or U7341 (N_7341,N_580,N_1547);
nand U7342 (N_7342,N_4623,N_3492);
nand U7343 (N_7343,N_2368,N_1635);
nor U7344 (N_7344,N_4734,N_1000);
xnor U7345 (N_7345,N_1111,N_4744);
nand U7346 (N_7346,N_2548,N_1944);
or U7347 (N_7347,N_4519,N_2857);
xor U7348 (N_7348,N_4006,N_3586);
or U7349 (N_7349,N_4996,N_2444);
and U7350 (N_7350,N_544,N_1447);
nand U7351 (N_7351,N_487,N_136);
or U7352 (N_7352,N_4696,N_4270);
and U7353 (N_7353,N_842,N_3653);
nand U7354 (N_7354,N_1713,N_3778);
nand U7355 (N_7355,N_3181,N_1379);
nor U7356 (N_7356,N_1597,N_988);
and U7357 (N_7357,N_2182,N_3243);
nand U7358 (N_7358,N_971,N_2833);
or U7359 (N_7359,N_1218,N_1193);
nor U7360 (N_7360,N_464,N_1010);
or U7361 (N_7361,N_4498,N_509);
nor U7362 (N_7362,N_3913,N_4845);
xnor U7363 (N_7363,N_4344,N_2637);
or U7364 (N_7364,N_2257,N_4417);
nor U7365 (N_7365,N_1771,N_4251);
nand U7366 (N_7366,N_811,N_4048);
nor U7367 (N_7367,N_4371,N_3012);
and U7368 (N_7368,N_840,N_4809);
xor U7369 (N_7369,N_4594,N_1167);
and U7370 (N_7370,N_668,N_1500);
and U7371 (N_7371,N_2791,N_903);
or U7372 (N_7372,N_1069,N_3031);
or U7373 (N_7373,N_1761,N_2789);
or U7374 (N_7374,N_2586,N_742);
xor U7375 (N_7375,N_3213,N_1814);
nor U7376 (N_7376,N_3327,N_4783);
nor U7377 (N_7377,N_2640,N_4859);
nor U7378 (N_7378,N_3823,N_1166);
nand U7379 (N_7379,N_2834,N_675);
and U7380 (N_7380,N_1455,N_344);
or U7381 (N_7381,N_4471,N_90);
or U7382 (N_7382,N_4990,N_221);
and U7383 (N_7383,N_4639,N_4494);
or U7384 (N_7384,N_127,N_1614);
nor U7385 (N_7385,N_2926,N_258);
nor U7386 (N_7386,N_4609,N_3378);
and U7387 (N_7387,N_1762,N_1604);
nor U7388 (N_7388,N_734,N_287);
or U7389 (N_7389,N_4709,N_1219);
nor U7390 (N_7390,N_1345,N_3638);
or U7391 (N_7391,N_2616,N_4935);
and U7392 (N_7392,N_2657,N_4540);
nor U7393 (N_7393,N_586,N_873);
nand U7394 (N_7394,N_1632,N_499);
nand U7395 (N_7395,N_4447,N_2689);
or U7396 (N_7396,N_2821,N_3341);
and U7397 (N_7397,N_4763,N_2730);
or U7398 (N_7398,N_766,N_999);
or U7399 (N_7399,N_2642,N_4564);
nor U7400 (N_7400,N_3247,N_2084);
or U7401 (N_7401,N_1188,N_4297);
xnor U7402 (N_7402,N_3018,N_954);
nor U7403 (N_7403,N_4534,N_2794);
or U7404 (N_7404,N_3436,N_1183);
nor U7405 (N_7405,N_1504,N_4865);
or U7406 (N_7406,N_4336,N_1233);
and U7407 (N_7407,N_1507,N_4397);
and U7408 (N_7408,N_2507,N_4215);
nand U7409 (N_7409,N_807,N_1033);
xor U7410 (N_7410,N_423,N_3069);
and U7411 (N_7411,N_4156,N_124);
and U7412 (N_7412,N_2871,N_2406);
or U7413 (N_7413,N_4063,N_3314);
and U7414 (N_7414,N_2347,N_2274);
or U7415 (N_7415,N_867,N_237);
nand U7416 (N_7416,N_4169,N_3052);
nor U7417 (N_7417,N_2690,N_3644);
and U7418 (N_7418,N_1545,N_1531);
and U7419 (N_7419,N_4925,N_96);
or U7420 (N_7420,N_4204,N_2712);
and U7421 (N_7421,N_4146,N_153);
nand U7422 (N_7422,N_3860,N_3145);
xor U7423 (N_7423,N_2697,N_4584);
and U7424 (N_7424,N_1751,N_2995);
nand U7425 (N_7425,N_2824,N_4039);
or U7426 (N_7426,N_3798,N_3990);
or U7427 (N_7427,N_1396,N_1246);
nand U7428 (N_7428,N_1322,N_4334);
and U7429 (N_7429,N_2832,N_3339);
nor U7430 (N_7430,N_2418,N_2735);
nor U7431 (N_7431,N_2109,N_0);
nand U7432 (N_7432,N_2896,N_2370);
and U7433 (N_7433,N_3838,N_1718);
and U7434 (N_7434,N_1315,N_2439);
and U7435 (N_7435,N_3261,N_48);
nand U7436 (N_7436,N_1266,N_3048);
nand U7437 (N_7437,N_4149,N_2477);
nand U7438 (N_7438,N_691,N_4022);
or U7439 (N_7439,N_2718,N_2967);
or U7440 (N_7440,N_2726,N_1923);
or U7441 (N_7441,N_2306,N_3759);
nor U7442 (N_7442,N_4576,N_1670);
nand U7443 (N_7443,N_1073,N_936);
nand U7444 (N_7444,N_1619,N_1882);
or U7445 (N_7445,N_821,N_3950);
or U7446 (N_7446,N_3026,N_567);
and U7447 (N_7447,N_2596,N_635);
nor U7448 (N_7448,N_4439,N_323);
xor U7449 (N_7449,N_3431,N_1727);
nor U7450 (N_7450,N_3617,N_2536);
or U7451 (N_7451,N_2459,N_4827);
nor U7452 (N_7452,N_3276,N_2702);
nand U7453 (N_7453,N_2959,N_948);
xor U7454 (N_7454,N_4797,N_2552);
or U7455 (N_7455,N_3825,N_4962);
nand U7456 (N_7456,N_3161,N_3135);
or U7457 (N_7457,N_1688,N_3219);
xnor U7458 (N_7458,N_4991,N_1042);
nor U7459 (N_7459,N_1444,N_1867);
nand U7460 (N_7460,N_688,N_3831);
and U7461 (N_7461,N_4724,N_3312);
xnor U7462 (N_7462,N_1753,N_1348);
xnor U7463 (N_7463,N_4181,N_663);
nand U7464 (N_7464,N_1366,N_1054);
nand U7465 (N_7465,N_571,N_3218);
nand U7466 (N_7466,N_3023,N_4789);
or U7467 (N_7467,N_14,N_630);
xor U7468 (N_7468,N_430,N_4427);
nand U7469 (N_7469,N_956,N_4160);
nand U7470 (N_7470,N_254,N_4411);
and U7471 (N_7471,N_4664,N_3864);
xor U7472 (N_7472,N_2206,N_459);
xnor U7473 (N_7473,N_3931,N_3064);
nor U7474 (N_7474,N_605,N_2455);
and U7475 (N_7475,N_1914,N_3674);
and U7476 (N_7476,N_3453,N_1300);
xnor U7477 (N_7477,N_4295,N_1653);
or U7478 (N_7478,N_4429,N_4277);
nor U7479 (N_7479,N_4748,N_131);
and U7480 (N_7480,N_4428,N_89);
nor U7481 (N_7481,N_438,N_3274);
xor U7482 (N_7482,N_3767,N_135);
or U7483 (N_7483,N_4821,N_1421);
and U7484 (N_7484,N_2795,N_4912);
nor U7485 (N_7485,N_1921,N_1101);
or U7486 (N_7486,N_2597,N_3011);
or U7487 (N_7487,N_1645,N_4236);
and U7488 (N_7488,N_1947,N_4468);
or U7489 (N_7489,N_1617,N_414);
nand U7490 (N_7490,N_193,N_2744);
nand U7491 (N_7491,N_583,N_947);
nand U7492 (N_7492,N_2331,N_179);
nand U7493 (N_7493,N_2071,N_3587);
xnor U7494 (N_7494,N_4890,N_2787);
xnor U7495 (N_7495,N_4967,N_147);
nor U7496 (N_7496,N_2679,N_2482);
and U7497 (N_7497,N_4461,N_2203);
and U7498 (N_7498,N_732,N_4244);
nand U7499 (N_7499,N_4340,N_3828);
and U7500 (N_7500,N_3686,N_3190);
and U7501 (N_7501,N_4166,N_2693);
or U7502 (N_7502,N_4489,N_4375);
nor U7503 (N_7503,N_4671,N_593);
nor U7504 (N_7504,N_2876,N_995);
xnor U7505 (N_7505,N_4863,N_2602);
nor U7506 (N_7506,N_4709,N_2136);
nor U7507 (N_7507,N_1221,N_1382);
xnor U7508 (N_7508,N_1029,N_4289);
nand U7509 (N_7509,N_14,N_1953);
and U7510 (N_7510,N_565,N_1753);
nand U7511 (N_7511,N_225,N_3601);
xnor U7512 (N_7512,N_2351,N_1392);
xnor U7513 (N_7513,N_4146,N_2177);
and U7514 (N_7514,N_3516,N_4907);
xnor U7515 (N_7515,N_3486,N_2671);
or U7516 (N_7516,N_4813,N_257);
nor U7517 (N_7517,N_4484,N_3363);
or U7518 (N_7518,N_4053,N_2360);
nand U7519 (N_7519,N_812,N_1095);
xnor U7520 (N_7520,N_2700,N_4407);
or U7521 (N_7521,N_4098,N_4320);
and U7522 (N_7522,N_4172,N_343);
and U7523 (N_7523,N_2462,N_2067);
xnor U7524 (N_7524,N_2053,N_910);
nand U7525 (N_7525,N_1622,N_4195);
nand U7526 (N_7526,N_546,N_84);
nand U7527 (N_7527,N_3897,N_1714);
xnor U7528 (N_7528,N_2584,N_2345);
and U7529 (N_7529,N_4500,N_1694);
nand U7530 (N_7530,N_2586,N_2528);
or U7531 (N_7531,N_629,N_1184);
xnor U7532 (N_7532,N_607,N_1740);
nand U7533 (N_7533,N_1238,N_3051);
and U7534 (N_7534,N_4943,N_4929);
nor U7535 (N_7535,N_1179,N_4810);
or U7536 (N_7536,N_1498,N_1502);
or U7537 (N_7537,N_4539,N_3411);
and U7538 (N_7538,N_3117,N_2620);
xor U7539 (N_7539,N_4145,N_1697);
xnor U7540 (N_7540,N_2879,N_4890);
and U7541 (N_7541,N_4829,N_1462);
xnor U7542 (N_7542,N_684,N_4857);
xnor U7543 (N_7543,N_3473,N_2526);
or U7544 (N_7544,N_4067,N_3366);
xnor U7545 (N_7545,N_2598,N_1786);
xor U7546 (N_7546,N_4177,N_2271);
or U7547 (N_7547,N_286,N_1977);
nor U7548 (N_7548,N_2795,N_868);
or U7549 (N_7549,N_474,N_4358);
xor U7550 (N_7550,N_4906,N_2609);
and U7551 (N_7551,N_3102,N_3708);
xor U7552 (N_7552,N_3290,N_986);
and U7553 (N_7553,N_663,N_3646);
or U7554 (N_7554,N_4951,N_2287);
nor U7555 (N_7555,N_260,N_4876);
nand U7556 (N_7556,N_361,N_4177);
nor U7557 (N_7557,N_920,N_1126);
xor U7558 (N_7558,N_3046,N_4109);
nor U7559 (N_7559,N_4113,N_2155);
or U7560 (N_7560,N_2472,N_1271);
nand U7561 (N_7561,N_3660,N_1350);
nand U7562 (N_7562,N_2594,N_3828);
nor U7563 (N_7563,N_4542,N_779);
nand U7564 (N_7564,N_4704,N_1382);
or U7565 (N_7565,N_3795,N_3535);
xnor U7566 (N_7566,N_3146,N_301);
xor U7567 (N_7567,N_67,N_439);
nor U7568 (N_7568,N_3986,N_1714);
nand U7569 (N_7569,N_4619,N_2843);
nand U7570 (N_7570,N_1253,N_789);
nand U7571 (N_7571,N_3687,N_800);
nor U7572 (N_7572,N_3694,N_4211);
nand U7573 (N_7573,N_2608,N_244);
or U7574 (N_7574,N_3448,N_4645);
nor U7575 (N_7575,N_349,N_3033);
nand U7576 (N_7576,N_1649,N_3214);
nand U7577 (N_7577,N_1464,N_1397);
or U7578 (N_7578,N_3090,N_2353);
xor U7579 (N_7579,N_4064,N_472);
or U7580 (N_7580,N_4652,N_3303);
nor U7581 (N_7581,N_1774,N_237);
nor U7582 (N_7582,N_3829,N_4344);
or U7583 (N_7583,N_212,N_3083);
xor U7584 (N_7584,N_2145,N_2754);
or U7585 (N_7585,N_3345,N_3645);
nor U7586 (N_7586,N_3815,N_1199);
nor U7587 (N_7587,N_856,N_3935);
nor U7588 (N_7588,N_263,N_313);
or U7589 (N_7589,N_3053,N_4548);
and U7590 (N_7590,N_409,N_4552);
nor U7591 (N_7591,N_3557,N_4438);
and U7592 (N_7592,N_3571,N_32);
or U7593 (N_7593,N_2614,N_2357);
xnor U7594 (N_7594,N_3174,N_4892);
nor U7595 (N_7595,N_159,N_267);
and U7596 (N_7596,N_4103,N_2905);
or U7597 (N_7597,N_3155,N_2676);
nor U7598 (N_7598,N_1232,N_1046);
xnor U7599 (N_7599,N_3800,N_1619);
xnor U7600 (N_7600,N_2809,N_2765);
or U7601 (N_7601,N_4404,N_679);
nor U7602 (N_7602,N_3660,N_1039);
and U7603 (N_7603,N_2495,N_3436);
nor U7604 (N_7604,N_1161,N_808);
xnor U7605 (N_7605,N_572,N_2800);
or U7606 (N_7606,N_2474,N_2567);
nor U7607 (N_7607,N_2488,N_736);
nor U7608 (N_7608,N_539,N_2505);
nand U7609 (N_7609,N_2759,N_4123);
xor U7610 (N_7610,N_4108,N_4814);
xnor U7611 (N_7611,N_3205,N_4516);
and U7612 (N_7612,N_2393,N_2814);
and U7613 (N_7613,N_1514,N_3514);
xor U7614 (N_7614,N_233,N_4498);
nor U7615 (N_7615,N_1052,N_57);
and U7616 (N_7616,N_1309,N_408);
xor U7617 (N_7617,N_1593,N_2583);
xnor U7618 (N_7618,N_3544,N_4051);
or U7619 (N_7619,N_4851,N_4421);
or U7620 (N_7620,N_54,N_73);
nand U7621 (N_7621,N_3674,N_2258);
xor U7622 (N_7622,N_4738,N_850);
xnor U7623 (N_7623,N_3397,N_1516);
nor U7624 (N_7624,N_2099,N_4993);
xor U7625 (N_7625,N_17,N_2649);
xnor U7626 (N_7626,N_1188,N_4516);
nand U7627 (N_7627,N_2267,N_1947);
and U7628 (N_7628,N_2136,N_3080);
xor U7629 (N_7629,N_959,N_4101);
nand U7630 (N_7630,N_1362,N_490);
xor U7631 (N_7631,N_1480,N_1475);
xnor U7632 (N_7632,N_2927,N_800);
xor U7633 (N_7633,N_1523,N_653);
nand U7634 (N_7634,N_2662,N_551);
xnor U7635 (N_7635,N_1936,N_3980);
nor U7636 (N_7636,N_2223,N_4925);
nand U7637 (N_7637,N_4828,N_2414);
and U7638 (N_7638,N_1676,N_638);
nand U7639 (N_7639,N_1801,N_2168);
or U7640 (N_7640,N_1576,N_1538);
xnor U7641 (N_7641,N_2555,N_4367);
nand U7642 (N_7642,N_3012,N_4241);
xor U7643 (N_7643,N_4733,N_1568);
or U7644 (N_7644,N_2880,N_4876);
nor U7645 (N_7645,N_3677,N_3206);
xor U7646 (N_7646,N_4552,N_2772);
and U7647 (N_7647,N_4700,N_3890);
nand U7648 (N_7648,N_846,N_3381);
or U7649 (N_7649,N_2187,N_4237);
nor U7650 (N_7650,N_586,N_4439);
xor U7651 (N_7651,N_3869,N_4076);
nand U7652 (N_7652,N_2569,N_668);
and U7653 (N_7653,N_3466,N_424);
and U7654 (N_7654,N_2906,N_4081);
or U7655 (N_7655,N_1112,N_4656);
nand U7656 (N_7656,N_2900,N_4519);
nor U7657 (N_7657,N_2047,N_3017);
xor U7658 (N_7658,N_3678,N_4760);
or U7659 (N_7659,N_4985,N_3042);
xor U7660 (N_7660,N_92,N_402);
nor U7661 (N_7661,N_378,N_3967);
nand U7662 (N_7662,N_437,N_2974);
xor U7663 (N_7663,N_53,N_2977);
xnor U7664 (N_7664,N_4881,N_541);
and U7665 (N_7665,N_1021,N_1243);
nand U7666 (N_7666,N_2683,N_563);
xor U7667 (N_7667,N_2942,N_2152);
or U7668 (N_7668,N_1927,N_4873);
and U7669 (N_7669,N_1204,N_4225);
and U7670 (N_7670,N_610,N_1117);
xnor U7671 (N_7671,N_1100,N_3826);
and U7672 (N_7672,N_2276,N_4871);
nor U7673 (N_7673,N_2054,N_4167);
nand U7674 (N_7674,N_2600,N_4052);
nand U7675 (N_7675,N_3676,N_4515);
nand U7676 (N_7676,N_2966,N_3621);
or U7677 (N_7677,N_3157,N_3822);
and U7678 (N_7678,N_1514,N_3196);
nor U7679 (N_7679,N_2293,N_4801);
or U7680 (N_7680,N_2613,N_2072);
and U7681 (N_7681,N_4942,N_765);
and U7682 (N_7682,N_1962,N_4196);
and U7683 (N_7683,N_437,N_2395);
or U7684 (N_7684,N_1972,N_1748);
or U7685 (N_7685,N_4165,N_249);
xor U7686 (N_7686,N_2179,N_541);
nand U7687 (N_7687,N_2192,N_229);
or U7688 (N_7688,N_4604,N_2988);
nand U7689 (N_7689,N_502,N_1166);
and U7690 (N_7690,N_330,N_2645);
nor U7691 (N_7691,N_1134,N_2374);
and U7692 (N_7692,N_1353,N_3395);
nand U7693 (N_7693,N_4777,N_4774);
and U7694 (N_7694,N_988,N_3058);
nand U7695 (N_7695,N_249,N_2882);
or U7696 (N_7696,N_1689,N_2604);
and U7697 (N_7697,N_1527,N_1477);
xor U7698 (N_7698,N_2515,N_2985);
or U7699 (N_7699,N_2728,N_1688);
nor U7700 (N_7700,N_161,N_3030);
xnor U7701 (N_7701,N_4007,N_492);
or U7702 (N_7702,N_3193,N_1199);
nand U7703 (N_7703,N_245,N_1602);
and U7704 (N_7704,N_1894,N_1216);
or U7705 (N_7705,N_3692,N_4046);
xor U7706 (N_7706,N_12,N_1971);
nand U7707 (N_7707,N_4059,N_4863);
nor U7708 (N_7708,N_4686,N_3874);
nand U7709 (N_7709,N_4543,N_59);
xor U7710 (N_7710,N_3525,N_1200);
or U7711 (N_7711,N_2750,N_1629);
and U7712 (N_7712,N_1365,N_626);
nand U7713 (N_7713,N_586,N_495);
xnor U7714 (N_7714,N_3127,N_3694);
and U7715 (N_7715,N_1791,N_4447);
nand U7716 (N_7716,N_3933,N_2254);
nor U7717 (N_7717,N_221,N_1143);
and U7718 (N_7718,N_1833,N_899);
and U7719 (N_7719,N_1374,N_1136);
or U7720 (N_7720,N_2447,N_204);
nand U7721 (N_7721,N_3171,N_1869);
xnor U7722 (N_7722,N_3569,N_2008);
nand U7723 (N_7723,N_3510,N_3789);
xnor U7724 (N_7724,N_1788,N_4170);
nor U7725 (N_7725,N_4876,N_3827);
nor U7726 (N_7726,N_4599,N_268);
nand U7727 (N_7727,N_3766,N_1393);
or U7728 (N_7728,N_3673,N_3670);
xor U7729 (N_7729,N_1567,N_2328);
and U7730 (N_7730,N_1222,N_3860);
or U7731 (N_7731,N_525,N_1998);
and U7732 (N_7732,N_3238,N_2013);
or U7733 (N_7733,N_769,N_2930);
nand U7734 (N_7734,N_2002,N_1963);
and U7735 (N_7735,N_1521,N_3759);
nor U7736 (N_7736,N_4502,N_2124);
and U7737 (N_7737,N_3690,N_3996);
nor U7738 (N_7738,N_2052,N_4192);
nor U7739 (N_7739,N_4505,N_2695);
and U7740 (N_7740,N_4007,N_1210);
nand U7741 (N_7741,N_286,N_2311);
or U7742 (N_7742,N_1713,N_3581);
nand U7743 (N_7743,N_4033,N_2997);
nor U7744 (N_7744,N_4012,N_3149);
and U7745 (N_7745,N_350,N_1147);
nor U7746 (N_7746,N_4743,N_3863);
or U7747 (N_7747,N_248,N_3821);
xor U7748 (N_7748,N_604,N_2767);
and U7749 (N_7749,N_3052,N_2882);
or U7750 (N_7750,N_3593,N_1811);
or U7751 (N_7751,N_3391,N_4355);
nor U7752 (N_7752,N_2282,N_2269);
or U7753 (N_7753,N_182,N_4202);
nand U7754 (N_7754,N_4180,N_1069);
and U7755 (N_7755,N_1957,N_2609);
or U7756 (N_7756,N_3769,N_3426);
and U7757 (N_7757,N_884,N_4503);
and U7758 (N_7758,N_2403,N_1719);
and U7759 (N_7759,N_325,N_1281);
or U7760 (N_7760,N_3970,N_1006);
xor U7761 (N_7761,N_917,N_3019);
xor U7762 (N_7762,N_3677,N_3143);
and U7763 (N_7763,N_4524,N_1164);
and U7764 (N_7764,N_4254,N_3110);
nand U7765 (N_7765,N_3493,N_2505);
and U7766 (N_7766,N_4455,N_1003);
and U7767 (N_7767,N_1772,N_155);
xor U7768 (N_7768,N_3038,N_1429);
or U7769 (N_7769,N_1382,N_1083);
xnor U7770 (N_7770,N_1897,N_4689);
nand U7771 (N_7771,N_3994,N_691);
and U7772 (N_7772,N_3055,N_3643);
nor U7773 (N_7773,N_1475,N_4738);
xor U7774 (N_7774,N_1368,N_766);
and U7775 (N_7775,N_3081,N_2242);
nand U7776 (N_7776,N_2080,N_1202);
or U7777 (N_7777,N_3331,N_3362);
xnor U7778 (N_7778,N_3273,N_2222);
and U7779 (N_7779,N_855,N_2923);
or U7780 (N_7780,N_4372,N_1628);
nand U7781 (N_7781,N_2603,N_2102);
and U7782 (N_7782,N_1183,N_726);
nor U7783 (N_7783,N_2940,N_1277);
nor U7784 (N_7784,N_4973,N_1994);
and U7785 (N_7785,N_1361,N_2604);
nand U7786 (N_7786,N_2935,N_3006);
xnor U7787 (N_7787,N_4658,N_1282);
or U7788 (N_7788,N_3236,N_4231);
or U7789 (N_7789,N_1421,N_4141);
nor U7790 (N_7790,N_3518,N_4508);
and U7791 (N_7791,N_2909,N_1573);
nor U7792 (N_7792,N_2894,N_3982);
or U7793 (N_7793,N_317,N_846);
or U7794 (N_7794,N_3139,N_1645);
nand U7795 (N_7795,N_1401,N_3412);
or U7796 (N_7796,N_2032,N_3431);
xor U7797 (N_7797,N_2242,N_4801);
nand U7798 (N_7798,N_163,N_2164);
nor U7799 (N_7799,N_1598,N_910);
nor U7800 (N_7800,N_2098,N_2345);
or U7801 (N_7801,N_1377,N_510);
and U7802 (N_7802,N_3654,N_4789);
or U7803 (N_7803,N_2112,N_1965);
xnor U7804 (N_7804,N_730,N_4976);
xor U7805 (N_7805,N_2979,N_1989);
nor U7806 (N_7806,N_4677,N_4214);
and U7807 (N_7807,N_4223,N_2711);
nor U7808 (N_7808,N_4329,N_4055);
or U7809 (N_7809,N_3977,N_2760);
xor U7810 (N_7810,N_1050,N_2053);
and U7811 (N_7811,N_4063,N_1396);
or U7812 (N_7812,N_2681,N_2953);
xor U7813 (N_7813,N_4728,N_2779);
nand U7814 (N_7814,N_4907,N_1294);
xor U7815 (N_7815,N_1709,N_1559);
or U7816 (N_7816,N_65,N_848);
and U7817 (N_7817,N_2569,N_1391);
xor U7818 (N_7818,N_4891,N_4921);
nand U7819 (N_7819,N_112,N_3568);
nor U7820 (N_7820,N_2318,N_3914);
and U7821 (N_7821,N_833,N_3769);
xnor U7822 (N_7822,N_4482,N_4955);
and U7823 (N_7823,N_2746,N_2681);
nand U7824 (N_7824,N_3343,N_4305);
nand U7825 (N_7825,N_4817,N_4122);
and U7826 (N_7826,N_4305,N_745);
or U7827 (N_7827,N_1479,N_3361);
xnor U7828 (N_7828,N_4162,N_4241);
and U7829 (N_7829,N_2711,N_2098);
nor U7830 (N_7830,N_3049,N_3830);
nor U7831 (N_7831,N_4173,N_1595);
and U7832 (N_7832,N_4584,N_4697);
or U7833 (N_7833,N_2772,N_4800);
nand U7834 (N_7834,N_3386,N_311);
and U7835 (N_7835,N_2352,N_3709);
nor U7836 (N_7836,N_222,N_3969);
nor U7837 (N_7837,N_2679,N_1083);
nor U7838 (N_7838,N_1452,N_3486);
or U7839 (N_7839,N_155,N_1856);
xnor U7840 (N_7840,N_4680,N_2591);
and U7841 (N_7841,N_3866,N_1491);
nand U7842 (N_7842,N_4707,N_1605);
nand U7843 (N_7843,N_664,N_4785);
or U7844 (N_7844,N_398,N_3589);
xnor U7845 (N_7845,N_3570,N_3310);
nand U7846 (N_7846,N_1786,N_263);
nand U7847 (N_7847,N_861,N_1726);
or U7848 (N_7848,N_1423,N_3828);
or U7849 (N_7849,N_4813,N_3484);
or U7850 (N_7850,N_2407,N_2903);
and U7851 (N_7851,N_3450,N_2881);
nor U7852 (N_7852,N_4100,N_4268);
nand U7853 (N_7853,N_492,N_2094);
nor U7854 (N_7854,N_2488,N_3240);
and U7855 (N_7855,N_1346,N_2196);
and U7856 (N_7856,N_1073,N_4568);
xor U7857 (N_7857,N_1468,N_3056);
nor U7858 (N_7858,N_751,N_781);
nor U7859 (N_7859,N_3409,N_771);
nor U7860 (N_7860,N_2139,N_4044);
xnor U7861 (N_7861,N_4571,N_1918);
and U7862 (N_7862,N_990,N_3658);
xor U7863 (N_7863,N_1791,N_4431);
xor U7864 (N_7864,N_4997,N_572);
or U7865 (N_7865,N_2241,N_1858);
and U7866 (N_7866,N_4257,N_4018);
nor U7867 (N_7867,N_3040,N_1132);
nor U7868 (N_7868,N_1604,N_4572);
or U7869 (N_7869,N_4113,N_1948);
or U7870 (N_7870,N_701,N_610);
nor U7871 (N_7871,N_4441,N_610);
and U7872 (N_7872,N_3271,N_1551);
xnor U7873 (N_7873,N_699,N_3348);
and U7874 (N_7874,N_1226,N_2368);
nor U7875 (N_7875,N_431,N_4657);
nand U7876 (N_7876,N_4496,N_3051);
nor U7877 (N_7877,N_2815,N_3072);
xnor U7878 (N_7878,N_2042,N_4935);
or U7879 (N_7879,N_1668,N_2614);
nand U7880 (N_7880,N_1231,N_922);
and U7881 (N_7881,N_2810,N_964);
xor U7882 (N_7882,N_3180,N_2048);
or U7883 (N_7883,N_3732,N_1209);
or U7884 (N_7884,N_3217,N_1686);
xnor U7885 (N_7885,N_2275,N_593);
and U7886 (N_7886,N_2760,N_460);
nor U7887 (N_7887,N_2099,N_4654);
nand U7888 (N_7888,N_1410,N_3733);
and U7889 (N_7889,N_188,N_1727);
and U7890 (N_7890,N_3133,N_328);
or U7891 (N_7891,N_532,N_2721);
nand U7892 (N_7892,N_4279,N_801);
or U7893 (N_7893,N_2323,N_4031);
nor U7894 (N_7894,N_3835,N_4724);
nor U7895 (N_7895,N_3209,N_283);
nand U7896 (N_7896,N_576,N_3968);
nor U7897 (N_7897,N_4309,N_114);
xnor U7898 (N_7898,N_722,N_924);
nor U7899 (N_7899,N_2504,N_1747);
xnor U7900 (N_7900,N_1669,N_1528);
or U7901 (N_7901,N_119,N_4132);
and U7902 (N_7902,N_3913,N_829);
or U7903 (N_7903,N_1678,N_3991);
or U7904 (N_7904,N_2681,N_3057);
nand U7905 (N_7905,N_3276,N_3452);
nor U7906 (N_7906,N_3674,N_3750);
nor U7907 (N_7907,N_4088,N_4926);
and U7908 (N_7908,N_3915,N_4695);
xor U7909 (N_7909,N_1601,N_1029);
or U7910 (N_7910,N_516,N_3450);
nor U7911 (N_7911,N_4404,N_151);
or U7912 (N_7912,N_4458,N_4992);
nand U7913 (N_7913,N_1690,N_1515);
nand U7914 (N_7914,N_3624,N_3415);
nor U7915 (N_7915,N_514,N_3516);
or U7916 (N_7916,N_3176,N_4698);
xnor U7917 (N_7917,N_3896,N_4866);
nor U7918 (N_7918,N_173,N_1987);
and U7919 (N_7919,N_36,N_3612);
or U7920 (N_7920,N_4505,N_3803);
nand U7921 (N_7921,N_2763,N_3197);
xor U7922 (N_7922,N_4953,N_1580);
xor U7923 (N_7923,N_3093,N_161);
nand U7924 (N_7924,N_4153,N_1020);
xor U7925 (N_7925,N_3361,N_1458);
nand U7926 (N_7926,N_2513,N_2264);
xnor U7927 (N_7927,N_1866,N_46);
xnor U7928 (N_7928,N_4417,N_546);
or U7929 (N_7929,N_1110,N_4707);
nand U7930 (N_7930,N_4604,N_1346);
xor U7931 (N_7931,N_4433,N_1893);
or U7932 (N_7932,N_1670,N_831);
xnor U7933 (N_7933,N_1582,N_1985);
xnor U7934 (N_7934,N_4443,N_2083);
and U7935 (N_7935,N_1644,N_4859);
and U7936 (N_7936,N_2332,N_517);
and U7937 (N_7937,N_62,N_1688);
nand U7938 (N_7938,N_3795,N_2021);
xnor U7939 (N_7939,N_4200,N_4656);
nor U7940 (N_7940,N_2357,N_2349);
xnor U7941 (N_7941,N_19,N_2030);
nor U7942 (N_7942,N_1281,N_4700);
and U7943 (N_7943,N_3486,N_2425);
and U7944 (N_7944,N_3014,N_2179);
nand U7945 (N_7945,N_3688,N_3725);
and U7946 (N_7946,N_3475,N_3364);
xnor U7947 (N_7947,N_1013,N_4196);
nand U7948 (N_7948,N_2822,N_3257);
xor U7949 (N_7949,N_4501,N_2352);
nor U7950 (N_7950,N_467,N_4999);
and U7951 (N_7951,N_3375,N_1825);
nand U7952 (N_7952,N_3872,N_4210);
nor U7953 (N_7953,N_2691,N_823);
nand U7954 (N_7954,N_1033,N_2491);
xor U7955 (N_7955,N_1790,N_3579);
and U7956 (N_7956,N_280,N_737);
xnor U7957 (N_7957,N_3628,N_1533);
and U7958 (N_7958,N_2559,N_4202);
and U7959 (N_7959,N_4153,N_3401);
nor U7960 (N_7960,N_1921,N_1567);
nand U7961 (N_7961,N_2515,N_957);
xor U7962 (N_7962,N_726,N_714);
nor U7963 (N_7963,N_4707,N_4973);
and U7964 (N_7964,N_489,N_3168);
nor U7965 (N_7965,N_4407,N_314);
xnor U7966 (N_7966,N_2078,N_1673);
or U7967 (N_7967,N_639,N_673);
or U7968 (N_7968,N_2885,N_430);
nor U7969 (N_7969,N_2390,N_3702);
and U7970 (N_7970,N_1066,N_3253);
and U7971 (N_7971,N_3285,N_1403);
nor U7972 (N_7972,N_2764,N_974);
nor U7973 (N_7973,N_426,N_3177);
nor U7974 (N_7974,N_2647,N_3348);
nor U7975 (N_7975,N_4656,N_3365);
nor U7976 (N_7976,N_1005,N_3778);
nor U7977 (N_7977,N_1224,N_2610);
and U7978 (N_7978,N_345,N_3544);
xnor U7979 (N_7979,N_2954,N_665);
xor U7980 (N_7980,N_4736,N_2280);
or U7981 (N_7981,N_790,N_39);
xor U7982 (N_7982,N_3081,N_3347);
nor U7983 (N_7983,N_1973,N_1695);
xnor U7984 (N_7984,N_1011,N_2235);
or U7985 (N_7985,N_3704,N_2603);
nor U7986 (N_7986,N_1712,N_490);
and U7987 (N_7987,N_3147,N_4655);
and U7988 (N_7988,N_4867,N_974);
or U7989 (N_7989,N_4366,N_1286);
nor U7990 (N_7990,N_3047,N_4355);
nor U7991 (N_7991,N_3497,N_1413);
or U7992 (N_7992,N_1663,N_1295);
xnor U7993 (N_7993,N_11,N_2187);
nand U7994 (N_7994,N_4394,N_1836);
and U7995 (N_7995,N_943,N_621);
or U7996 (N_7996,N_2442,N_1551);
xnor U7997 (N_7997,N_2309,N_3840);
and U7998 (N_7998,N_638,N_803);
and U7999 (N_7999,N_1133,N_2409);
nor U8000 (N_8000,N_4040,N_3940);
and U8001 (N_8001,N_1027,N_1673);
nor U8002 (N_8002,N_3469,N_403);
nor U8003 (N_8003,N_998,N_2086);
nor U8004 (N_8004,N_4091,N_449);
nor U8005 (N_8005,N_474,N_3720);
or U8006 (N_8006,N_4208,N_2710);
or U8007 (N_8007,N_2988,N_1044);
xnor U8008 (N_8008,N_4416,N_1275);
and U8009 (N_8009,N_4869,N_259);
nand U8010 (N_8010,N_1356,N_4368);
and U8011 (N_8011,N_1036,N_1720);
and U8012 (N_8012,N_4345,N_4777);
and U8013 (N_8013,N_105,N_4194);
and U8014 (N_8014,N_909,N_626);
nand U8015 (N_8015,N_413,N_1673);
and U8016 (N_8016,N_4654,N_4637);
nor U8017 (N_8017,N_567,N_1121);
nor U8018 (N_8018,N_3472,N_783);
nor U8019 (N_8019,N_280,N_1126);
and U8020 (N_8020,N_3624,N_1395);
nor U8021 (N_8021,N_3337,N_4425);
or U8022 (N_8022,N_4753,N_364);
and U8023 (N_8023,N_4776,N_2510);
and U8024 (N_8024,N_954,N_4464);
nand U8025 (N_8025,N_2521,N_663);
nand U8026 (N_8026,N_4874,N_4229);
and U8027 (N_8027,N_3367,N_4477);
and U8028 (N_8028,N_3828,N_2029);
xor U8029 (N_8029,N_659,N_660);
nor U8030 (N_8030,N_1156,N_1946);
nor U8031 (N_8031,N_3920,N_3009);
xnor U8032 (N_8032,N_1331,N_515);
xor U8033 (N_8033,N_2711,N_2206);
or U8034 (N_8034,N_449,N_3723);
nand U8035 (N_8035,N_2732,N_4897);
nor U8036 (N_8036,N_1132,N_4324);
nor U8037 (N_8037,N_1696,N_1705);
and U8038 (N_8038,N_4915,N_2837);
nor U8039 (N_8039,N_303,N_3827);
xor U8040 (N_8040,N_3224,N_2890);
or U8041 (N_8041,N_4833,N_3776);
and U8042 (N_8042,N_571,N_2620);
nor U8043 (N_8043,N_479,N_3741);
or U8044 (N_8044,N_4845,N_4378);
or U8045 (N_8045,N_2391,N_1512);
nor U8046 (N_8046,N_99,N_1618);
nor U8047 (N_8047,N_2987,N_1502);
and U8048 (N_8048,N_385,N_3183);
or U8049 (N_8049,N_1160,N_4451);
nand U8050 (N_8050,N_663,N_3157);
and U8051 (N_8051,N_4575,N_655);
or U8052 (N_8052,N_1774,N_812);
or U8053 (N_8053,N_1478,N_2813);
or U8054 (N_8054,N_1921,N_3189);
nand U8055 (N_8055,N_134,N_264);
or U8056 (N_8056,N_4141,N_3068);
nor U8057 (N_8057,N_4077,N_645);
nor U8058 (N_8058,N_1817,N_2357);
nor U8059 (N_8059,N_3221,N_954);
nor U8060 (N_8060,N_544,N_2879);
nor U8061 (N_8061,N_2798,N_2318);
nand U8062 (N_8062,N_4054,N_2186);
or U8063 (N_8063,N_3597,N_4539);
or U8064 (N_8064,N_474,N_4543);
xor U8065 (N_8065,N_2155,N_3078);
xor U8066 (N_8066,N_4666,N_1621);
or U8067 (N_8067,N_2414,N_4575);
nor U8068 (N_8068,N_2599,N_3611);
and U8069 (N_8069,N_1639,N_3943);
nand U8070 (N_8070,N_1463,N_613);
or U8071 (N_8071,N_966,N_4830);
nand U8072 (N_8072,N_2196,N_2488);
or U8073 (N_8073,N_4740,N_4341);
and U8074 (N_8074,N_4361,N_409);
nor U8075 (N_8075,N_643,N_346);
xnor U8076 (N_8076,N_2913,N_559);
nor U8077 (N_8077,N_4555,N_1212);
or U8078 (N_8078,N_3679,N_2519);
or U8079 (N_8079,N_2243,N_3151);
and U8080 (N_8080,N_3284,N_4053);
nand U8081 (N_8081,N_2017,N_1636);
nor U8082 (N_8082,N_3355,N_3333);
and U8083 (N_8083,N_1511,N_1685);
or U8084 (N_8084,N_1154,N_531);
nand U8085 (N_8085,N_4222,N_4995);
xor U8086 (N_8086,N_1923,N_416);
nor U8087 (N_8087,N_2622,N_2153);
or U8088 (N_8088,N_2621,N_4874);
or U8089 (N_8089,N_2846,N_4781);
or U8090 (N_8090,N_1653,N_3221);
nand U8091 (N_8091,N_2731,N_3351);
nor U8092 (N_8092,N_1600,N_2463);
and U8093 (N_8093,N_905,N_4999);
nand U8094 (N_8094,N_2744,N_4191);
xor U8095 (N_8095,N_955,N_834);
nand U8096 (N_8096,N_398,N_1129);
nor U8097 (N_8097,N_3348,N_1951);
nor U8098 (N_8098,N_4195,N_216);
nand U8099 (N_8099,N_1528,N_2032);
xnor U8100 (N_8100,N_1600,N_4926);
xnor U8101 (N_8101,N_2910,N_879);
nand U8102 (N_8102,N_4530,N_1301);
and U8103 (N_8103,N_1059,N_1252);
nor U8104 (N_8104,N_3301,N_4562);
or U8105 (N_8105,N_4530,N_2414);
nor U8106 (N_8106,N_316,N_1876);
or U8107 (N_8107,N_1627,N_1041);
nand U8108 (N_8108,N_4897,N_3181);
xnor U8109 (N_8109,N_1187,N_3852);
xnor U8110 (N_8110,N_3905,N_801);
or U8111 (N_8111,N_2976,N_3068);
nand U8112 (N_8112,N_628,N_2201);
xnor U8113 (N_8113,N_4150,N_1492);
and U8114 (N_8114,N_1924,N_996);
and U8115 (N_8115,N_1392,N_4887);
or U8116 (N_8116,N_1521,N_245);
nor U8117 (N_8117,N_963,N_870);
xor U8118 (N_8118,N_1522,N_4384);
or U8119 (N_8119,N_3078,N_2124);
nor U8120 (N_8120,N_4794,N_3529);
nand U8121 (N_8121,N_579,N_3773);
or U8122 (N_8122,N_1648,N_3151);
and U8123 (N_8123,N_3005,N_2572);
or U8124 (N_8124,N_2255,N_3356);
and U8125 (N_8125,N_1561,N_428);
nor U8126 (N_8126,N_4578,N_3341);
nor U8127 (N_8127,N_3666,N_1885);
xor U8128 (N_8128,N_1449,N_1322);
nand U8129 (N_8129,N_4035,N_379);
and U8130 (N_8130,N_3665,N_2028);
xnor U8131 (N_8131,N_3142,N_3246);
or U8132 (N_8132,N_2620,N_813);
nor U8133 (N_8133,N_4576,N_552);
and U8134 (N_8134,N_2407,N_1587);
or U8135 (N_8135,N_2732,N_4565);
or U8136 (N_8136,N_839,N_2916);
and U8137 (N_8137,N_1852,N_2446);
or U8138 (N_8138,N_172,N_2000);
nor U8139 (N_8139,N_1478,N_3325);
and U8140 (N_8140,N_3202,N_3680);
or U8141 (N_8141,N_829,N_2246);
nor U8142 (N_8142,N_39,N_1912);
xnor U8143 (N_8143,N_652,N_3389);
xor U8144 (N_8144,N_1373,N_3675);
xnor U8145 (N_8145,N_1020,N_4280);
nand U8146 (N_8146,N_1146,N_2315);
or U8147 (N_8147,N_1184,N_1933);
nand U8148 (N_8148,N_1984,N_1295);
or U8149 (N_8149,N_4044,N_4571);
or U8150 (N_8150,N_4656,N_302);
and U8151 (N_8151,N_1012,N_2910);
nor U8152 (N_8152,N_318,N_3645);
xnor U8153 (N_8153,N_2880,N_1924);
xnor U8154 (N_8154,N_1926,N_2672);
xor U8155 (N_8155,N_2480,N_4423);
and U8156 (N_8156,N_1431,N_2187);
nand U8157 (N_8157,N_1878,N_2428);
nand U8158 (N_8158,N_270,N_334);
and U8159 (N_8159,N_1536,N_1106);
xnor U8160 (N_8160,N_3164,N_2715);
xnor U8161 (N_8161,N_583,N_4806);
or U8162 (N_8162,N_2897,N_1246);
nor U8163 (N_8163,N_4283,N_1242);
nand U8164 (N_8164,N_745,N_4806);
or U8165 (N_8165,N_533,N_1218);
and U8166 (N_8166,N_4840,N_2149);
nand U8167 (N_8167,N_3936,N_4714);
nand U8168 (N_8168,N_494,N_2095);
or U8169 (N_8169,N_4307,N_2157);
xnor U8170 (N_8170,N_1038,N_4571);
or U8171 (N_8171,N_1340,N_3948);
xor U8172 (N_8172,N_3007,N_2806);
xnor U8173 (N_8173,N_935,N_3865);
or U8174 (N_8174,N_3261,N_1327);
or U8175 (N_8175,N_1273,N_1475);
xnor U8176 (N_8176,N_3060,N_2807);
nand U8177 (N_8177,N_3054,N_4871);
and U8178 (N_8178,N_320,N_3944);
nand U8179 (N_8179,N_3423,N_3487);
or U8180 (N_8180,N_1440,N_2285);
and U8181 (N_8181,N_4363,N_3710);
xor U8182 (N_8182,N_1881,N_1032);
and U8183 (N_8183,N_1508,N_771);
and U8184 (N_8184,N_2407,N_1325);
nor U8185 (N_8185,N_4127,N_932);
nor U8186 (N_8186,N_1946,N_3709);
and U8187 (N_8187,N_272,N_3140);
xor U8188 (N_8188,N_4309,N_2907);
and U8189 (N_8189,N_3716,N_1752);
nor U8190 (N_8190,N_2203,N_1203);
nand U8191 (N_8191,N_4022,N_1147);
nand U8192 (N_8192,N_3682,N_247);
and U8193 (N_8193,N_2501,N_2709);
or U8194 (N_8194,N_630,N_4388);
or U8195 (N_8195,N_1332,N_464);
and U8196 (N_8196,N_855,N_1394);
nand U8197 (N_8197,N_1613,N_1897);
or U8198 (N_8198,N_3934,N_3633);
xor U8199 (N_8199,N_447,N_3604);
or U8200 (N_8200,N_514,N_3271);
nor U8201 (N_8201,N_3303,N_2152);
or U8202 (N_8202,N_275,N_3987);
or U8203 (N_8203,N_2733,N_600);
nand U8204 (N_8204,N_2227,N_4718);
nand U8205 (N_8205,N_3436,N_4919);
and U8206 (N_8206,N_3202,N_4917);
nand U8207 (N_8207,N_3452,N_1514);
xor U8208 (N_8208,N_2869,N_4964);
nor U8209 (N_8209,N_2089,N_1753);
or U8210 (N_8210,N_4685,N_2396);
or U8211 (N_8211,N_1412,N_4818);
or U8212 (N_8212,N_2571,N_3340);
nor U8213 (N_8213,N_2364,N_4892);
and U8214 (N_8214,N_1974,N_3402);
nor U8215 (N_8215,N_1312,N_4551);
nand U8216 (N_8216,N_1193,N_2544);
nor U8217 (N_8217,N_1812,N_4392);
xnor U8218 (N_8218,N_3317,N_2342);
and U8219 (N_8219,N_4646,N_1103);
and U8220 (N_8220,N_1832,N_4931);
and U8221 (N_8221,N_2997,N_2091);
and U8222 (N_8222,N_4848,N_754);
xor U8223 (N_8223,N_545,N_2360);
or U8224 (N_8224,N_2779,N_2099);
xnor U8225 (N_8225,N_538,N_2616);
nand U8226 (N_8226,N_1539,N_1118);
or U8227 (N_8227,N_3143,N_3616);
nand U8228 (N_8228,N_1935,N_4973);
or U8229 (N_8229,N_1947,N_1536);
or U8230 (N_8230,N_888,N_3269);
nor U8231 (N_8231,N_1760,N_3534);
or U8232 (N_8232,N_2786,N_602);
nor U8233 (N_8233,N_158,N_3252);
nor U8234 (N_8234,N_4206,N_3108);
and U8235 (N_8235,N_252,N_3376);
and U8236 (N_8236,N_4557,N_725);
nand U8237 (N_8237,N_3229,N_4957);
and U8238 (N_8238,N_3873,N_1234);
nand U8239 (N_8239,N_3483,N_940);
nor U8240 (N_8240,N_1318,N_1359);
xnor U8241 (N_8241,N_3522,N_4449);
nand U8242 (N_8242,N_1661,N_4288);
nor U8243 (N_8243,N_222,N_2444);
or U8244 (N_8244,N_1047,N_2600);
nand U8245 (N_8245,N_4206,N_1677);
xnor U8246 (N_8246,N_2651,N_3101);
and U8247 (N_8247,N_2618,N_3945);
nand U8248 (N_8248,N_4655,N_1884);
or U8249 (N_8249,N_3535,N_993);
nor U8250 (N_8250,N_3487,N_3947);
xnor U8251 (N_8251,N_1798,N_3323);
nand U8252 (N_8252,N_1843,N_3187);
xnor U8253 (N_8253,N_1544,N_3148);
nor U8254 (N_8254,N_2907,N_1490);
nand U8255 (N_8255,N_2023,N_1588);
nand U8256 (N_8256,N_3180,N_1772);
nor U8257 (N_8257,N_3205,N_3688);
or U8258 (N_8258,N_2056,N_3688);
and U8259 (N_8259,N_2514,N_3325);
or U8260 (N_8260,N_841,N_3696);
nor U8261 (N_8261,N_2282,N_1286);
xnor U8262 (N_8262,N_1547,N_3599);
nor U8263 (N_8263,N_66,N_4501);
and U8264 (N_8264,N_755,N_3864);
xnor U8265 (N_8265,N_3419,N_3728);
nand U8266 (N_8266,N_1363,N_1196);
and U8267 (N_8267,N_2501,N_4524);
or U8268 (N_8268,N_2154,N_4849);
and U8269 (N_8269,N_1810,N_1086);
xor U8270 (N_8270,N_2888,N_4236);
or U8271 (N_8271,N_178,N_4821);
nand U8272 (N_8272,N_2422,N_621);
nand U8273 (N_8273,N_59,N_2729);
or U8274 (N_8274,N_274,N_1973);
or U8275 (N_8275,N_656,N_4716);
nand U8276 (N_8276,N_2070,N_3829);
nand U8277 (N_8277,N_901,N_3291);
or U8278 (N_8278,N_4639,N_3233);
and U8279 (N_8279,N_4387,N_2117);
nand U8280 (N_8280,N_3506,N_4514);
xnor U8281 (N_8281,N_3607,N_2522);
xnor U8282 (N_8282,N_1734,N_2767);
and U8283 (N_8283,N_1660,N_1907);
or U8284 (N_8284,N_1894,N_1871);
nor U8285 (N_8285,N_4932,N_1687);
nor U8286 (N_8286,N_2278,N_3149);
xnor U8287 (N_8287,N_3423,N_2295);
nand U8288 (N_8288,N_1118,N_1577);
and U8289 (N_8289,N_1421,N_235);
nor U8290 (N_8290,N_269,N_2432);
or U8291 (N_8291,N_2022,N_18);
nand U8292 (N_8292,N_4501,N_3952);
nor U8293 (N_8293,N_1610,N_2674);
xor U8294 (N_8294,N_2334,N_3821);
nor U8295 (N_8295,N_4855,N_2684);
nor U8296 (N_8296,N_2713,N_1224);
and U8297 (N_8297,N_3248,N_2853);
nand U8298 (N_8298,N_3090,N_4906);
nor U8299 (N_8299,N_3492,N_3286);
nor U8300 (N_8300,N_900,N_2510);
and U8301 (N_8301,N_2900,N_4525);
nor U8302 (N_8302,N_2488,N_86);
and U8303 (N_8303,N_3924,N_28);
nand U8304 (N_8304,N_2231,N_2047);
xnor U8305 (N_8305,N_3523,N_3);
nand U8306 (N_8306,N_2965,N_79);
nor U8307 (N_8307,N_3663,N_1734);
nand U8308 (N_8308,N_2586,N_1557);
and U8309 (N_8309,N_2101,N_4529);
and U8310 (N_8310,N_2535,N_969);
nand U8311 (N_8311,N_4738,N_4879);
or U8312 (N_8312,N_4243,N_271);
nor U8313 (N_8313,N_3505,N_3608);
nor U8314 (N_8314,N_2735,N_1948);
and U8315 (N_8315,N_3966,N_4567);
nor U8316 (N_8316,N_766,N_670);
or U8317 (N_8317,N_896,N_3091);
and U8318 (N_8318,N_4176,N_2711);
or U8319 (N_8319,N_4836,N_3484);
and U8320 (N_8320,N_4339,N_3500);
xnor U8321 (N_8321,N_3020,N_4117);
xor U8322 (N_8322,N_2905,N_2415);
nand U8323 (N_8323,N_859,N_2849);
xnor U8324 (N_8324,N_4290,N_4416);
nor U8325 (N_8325,N_1439,N_4929);
or U8326 (N_8326,N_2319,N_4890);
or U8327 (N_8327,N_1216,N_4778);
nor U8328 (N_8328,N_2506,N_3129);
or U8329 (N_8329,N_4999,N_1366);
and U8330 (N_8330,N_3139,N_2779);
or U8331 (N_8331,N_2252,N_1649);
xor U8332 (N_8332,N_1993,N_4901);
or U8333 (N_8333,N_4532,N_4861);
nor U8334 (N_8334,N_859,N_1718);
xor U8335 (N_8335,N_3579,N_4572);
and U8336 (N_8336,N_4418,N_4675);
nand U8337 (N_8337,N_2533,N_2727);
nor U8338 (N_8338,N_3635,N_2763);
xnor U8339 (N_8339,N_3080,N_1154);
nor U8340 (N_8340,N_3085,N_1791);
and U8341 (N_8341,N_2893,N_1747);
xor U8342 (N_8342,N_3366,N_4723);
nand U8343 (N_8343,N_2568,N_2935);
and U8344 (N_8344,N_3148,N_3674);
and U8345 (N_8345,N_20,N_2486);
and U8346 (N_8346,N_1758,N_691);
nor U8347 (N_8347,N_1603,N_2141);
or U8348 (N_8348,N_4462,N_3060);
nand U8349 (N_8349,N_4702,N_3488);
or U8350 (N_8350,N_288,N_2669);
nor U8351 (N_8351,N_4656,N_1119);
xnor U8352 (N_8352,N_3392,N_4371);
and U8353 (N_8353,N_3024,N_2631);
and U8354 (N_8354,N_2129,N_2801);
or U8355 (N_8355,N_3831,N_449);
or U8356 (N_8356,N_2543,N_4247);
nor U8357 (N_8357,N_525,N_698);
and U8358 (N_8358,N_2372,N_1496);
or U8359 (N_8359,N_2867,N_1600);
or U8360 (N_8360,N_361,N_2175);
and U8361 (N_8361,N_2252,N_4071);
xor U8362 (N_8362,N_1515,N_3088);
nand U8363 (N_8363,N_4,N_3568);
nand U8364 (N_8364,N_2951,N_500);
nor U8365 (N_8365,N_2877,N_4851);
or U8366 (N_8366,N_473,N_4136);
and U8367 (N_8367,N_405,N_238);
xor U8368 (N_8368,N_825,N_2422);
xnor U8369 (N_8369,N_92,N_3137);
nand U8370 (N_8370,N_700,N_1886);
nand U8371 (N_8371,N_3116,N_874);
or U8372 (N_8372,N_4693,N_4142);
or U8373 (N_8373,N_3615,N_3327);
or U8374 (N_8374,N_1450,N_3501);
nand U8375 (N_8375,N_1890,N_2087);
or U8376 (N_8376,N_3595,N_1785);
xor U8377 (N_8377,N_845,N_1512);
xnor U8378 (N_8378,N_1482,N_3980);
nand U8379 (N_8379,N_2332,N_853);
and U8380 (N_8380,N_1772,N_2853);
nand U8381 (N_8381,N_674,N_1216);
nor U8382 (N_8382,N_1878,N_4383);
or U8383 (N_8383,N_3327,N_2614);
nor U8384 (N_8384,N_2209,N_368);
xnor U8385 (N_8385,N_3613,N_3282);
nor U8386 (N_8386,N_4971,N_3222);
xnor U8387 (N_8387,N_3039,N_2670);
xnor U8388 (N_8388,N_3144,N_3146);
or U8389 (N_8389,N_3016,N_4284);
nor U8390 (N_8390,N_2945,N_1766);
or U8391 (N_8391,N_532,N_4434);
nor U8392 (N_8392,N_1652,N_4014);
nand U8393 (N_8393,N_2149,N_1283);
xor U8394 (N_8394,N_1152,N_3676);
xor U8395 (N_8395,N_4257,N_4571);
or U8396 (N_8396,N_2200,N_4056);
nor U8397 (N_8397,N_3670,N_2661);
nor U8398 (N_8398,N_2050,N_3349);
or U8399 (N_8399,N_3466,N_3295);
nand U8400 (N_8400,N_520,N_1335);
xor U8401 (N_8401,N_2257,N_3880);
and U8402 (N_8402,N_4009,N_2558);
xor U8403 (N_8403,N_2430,N_3675);
nor U8404 (N_8404,N_3417,N_556);
nand U8405 (N_8405,N_2149,N_4435);
or U8406 (N_8406,N_2568,N_1639);
or U8407 (N_8407,N_519,N_774);
nor U8408 (N_8408,N_1182,N_2909);
and U8409 (N_8409,N_283,N_1433);
and U8410 (N_8410,N_4657,N_1781);
or U8411 (N_8411,N_1202,N_831);
nand U8412 (N_8412,N_1531,N_50);
nand U8413 (N_8413,N_1065,N_1768);
nor U8414 (N_8414,N_1902,N_310);
and U8415 (N_8415,N_731,N_1081);
and U8416 (N_8416,N_2434,N_3123);
xor U8417 (N_8417,N_1942,N_1826);
or U8418 (N_8418,N_4246,N_1821);
nor U8419 (N_8419,N_2834,N_4960);
and U8420 (N_8420,N_2888,N_1258);
nand U8421 (N_8421,N_4183,N_3120);
xnor U8422 (N_8422,N_1727,N_922);
xor U8423 (N_8423,N_880,N_4543);
or U8424 (N_8424,N_2871,N_1727);
nand U8425 (N_8425,N_1023,N_2802);
nand U8426 (N_8426,N_2767,N_4048);
nor U8427 (N_8427,N_1449,N_3031);
and U8428 (N_8428,N_4214,N_4317);
or U8429 (N_8429,N_4444,N_4750);
xnor U8430 (N_8430,N_930,N_4721);
and U8431 (N_8431,N_3971,N_3806);
xnor U8432 (N_8432,N_1184,N_2482);
or U8433 (N_8433,N_733,N_2614);
nor U8434 (N_8434,N_1340,N_1935);
nand U8435 (N_8435,N_4839,N_3478);
nor U8436 (N_8436,N_2632,N_1541);
nor U8437 (N_8437,N_4346,N_1537);
nand U8438 (N_8438,N_4292,N_3332);
or U8439 (N_8439,N_4460,N_2327);
and U8440 (N_8440,N_492,N_1455);
nand U8441 (N_8441,N_3775,N_3368);
or U8442 (N_8442,N_3625,N_867);
nand U8443 (N_8443,N_819,N_4112);
or U8444 (N_8444,N_1805,N_3399);
or U8445 (N_8445,N_768,N_539);
or U8446 (N_8446,N_238,N_1104);
or U8447 (N_8447,N_4772,N_1004);
or U8448 (N_8448,N_3640,N_2453);
nor U8449 (N_8449,N_3610,N_3325);
and U8450 (N_8450,N_2425,N_404);
xnor U8451 (N_8451,N_3252,N_1779);
nor U8452 (N_8452,N_1645,N_468);
or U8453 (N_8453,N_1390,N_473);
or U8454 (N_8454,N_668,N_2188);
nor U8455 (N_8455,N_1330,N_2350);
nand U8456 (N_8456,N_1892,N_187);
or U8457 (N_8457,N_3855,N_3771);
nor U8458 (N_8458,N_4870,N_188);
xor U8459 (N_8459,N_2768,N_1190);
and U8460 (N_8460,N_351,N_832);
nor U8461 (N_8461,N_2998,N_914);
nand U8462 (N_8462,N_2141,N_2803);
xor U8463 (N_8463,N_2720,N_2280);
and U8464 (N_8464,N_3167,N_2201);
nor U8465 (N_8465,N_1962,N_3598);
and U8466 (N_8466,N_2901,N_323);
nand U8467 (N_8467,N_77,N_2139);
nand U8468 (N_8468,N_1444,N_4218);
or U8469 (N_8469,N_2258,N_1558);
xnor U8470 (N_8470,N_2118,N_4406);
or U8471 (N_8471,N_4088,N_4620);
and U8472 (N_8472,N_1253,N_466);
xor U8473 (N_8473,N_3766,N_3398);
nand U8474 (N_8474,N_1852,N_2827);
nor U8475 (N_8475,N_3463,N_4541);
and U8476 (N_8476,N_3493,N_3435);
xnor U8477 (N_8477,N_747,N_2701);
and U8478 (N_8478,N_3986,N_1330);
or U8479 (N_8479,N_4773,N_2119);
xor U8480 (N_8480,N_2561,N_4519);
and U8481 (N_8481,N_2798,N_2278);
nand U8482 (N_8482,N_1285,N_2461);
nand U8483 (N_8483,N_244,N_422);
xnor U8484 (N_8484,N_2294,N_236);
xnor U8485 (N_8485,N_218,N_4668);
nand U8486 (N_8486,N_2422,N_523);
nor U8487 (N_8487,N_839,N_4879);
nand U8488 (N_8488,N_2699,N_3951);
or U8489 (N_8489,N_1307,N_2854);
nand U8490 (N_8490,N_3273,N_1773);
or U8491 (N_8491,N_4743,N_3120);
nand U8492 (N_8492,N_3459,N_1360);
nand U8493 (N_8493,N_3131,N_935);
and U8494 (N_8494,N_2735,N_265);
and U8495 (N_8495,N_4722,N_91);
xnor U8496 (N_8496,N_1346,N_4712);
and U8497 (N_8497,N_4778,N_4418);
or U8498 (N_8498,N_995,N_3350);
or U8499 (N_8499,N_3516,N_835);
nor U8500 (N_8500,N_1721,N_3978);
nor U8501 (N_8501,N_3322,N_1322);
nor U8502 (N_8502,N_1558,N_2283);
nand U8503 (N_8503,N_2855,N_2863);
nor U8504 (N_8504,N_4029,N_4817);
or U8505 (N_8505,N_3135,N_1027);
xor U8506 (N_8506,N_1348,N_380);
nor U8507 (N_8507,N_3398,N_3796);
or U8508 (N_8508,N_3920,N_3238);
xnor U8509 (N_8509,N_3132,N_1256);
nand U8510 (N_8510,N_4063,N_806);
xnor U8511 (N_8511,N_3450,N_2790);
or U8512 (N_8512,N_4515,N_3415);
nor U8513 (N_8513,N_1230,N_4465);
or U8514 (N_8514,N_2117,N_338);
xor U8515 (N_8515,N_707,N_153);
and U8516 (N_8516,N_1597,N_2128);
nor U8517 (N_8517,N_4669,N_4046);
nor U8518 (N_8518,N_2682,N_1674);
nand U8519 (N_8519,N_198,N_462);
and U8520 (N_8520,N_201,N_1833);
nor U8521 (N_8521,N_511,N_351);
xor U8522 (N_8522,N_3254,N_4871);
and U8523 (N_8523,N_4950,N_4092);
or U8524 (N_8524,N_3758,N_2344);
and U8525 (N_8525,N_3759,N_3361);
and U8526 (N_8526,N_4477,N_2915);
nand U8527 (N_8527,N_1439,N_954);
and U8528 (N_8528,N_579,N_3534);
or U8529 (N_8529,N_3106,N_320);
or U8530 (N_8530,N_1198,N_322);
nor U8531 (N_8531,N_4609,N_581);
xor U8532 (N_8532,N_872,N_3713);
and U8533 (N_8533,N_4737,N_89);
or U8534 (N_8534,N_1692,N_2483);
nor U8535 (N_8535,N_1733,N_4469);
and U8536 (N_8536,N_4553,N_662);
xnor U8537 (N_8537,N_1234,N_234);
nand U8538 (N_8538,N_2246,N_1724);
nor U8539 (N_8539,N_1590,N_4099);
and U8540 (N_8540,N_4338,N_4764);
or U8541 (N_8541,N_2263,N_4482);
and U8542 (N_8542,N_140,N_1686);
nand U8543 (N_8543,N_1909,N_1516);
xor U8544 (N_8544,N_379,N_4436);
and U8545 (N_8545,N_4189,N_2479);
and U8546 (N_8546,N_4330,N_1247);
nor U8547 (N_8547,N_4339,N_1726);
nor U8548 (N_8548,N_3657,N_1210);
xnor U8549 (N_8549,N_2436,N_3907);
and U8550 (N_8550,N_2546,N_2004);
or U8551 (N_8551,N_2894,N_133);
xor U8552 (N_8552,N_959,N_4169);
and U8553 (N_8553,N_3556,N_1163);
xor U8554 (N_8554,N_156,N_2512);
or U8555 (N_8555,N_842,N_617);
and U8556 (N_8556,N_3968,N_4886);
and U8557 (N_8557,N_2664,N_3498);
xnor U8558 (N_8558,N_1764,N_1763);
nand U8559 (N_8559,N_3331,N_3173);
nor U8560 (N_8560,N_4016,N_89);
or U8561 (N_8561,N_2518,N_1352);
nor U8562 (N_8562,N_3683,N_2619);
nand U8563 (N_8563,N_3130,N_41);
xor U8564 (N_8564,N_4810,N_1839);
nand U8565 (N_8565,N_3648,N_4560);
nand U8566 (N_8566,N_569,N_1113);
nand U8567 (N_8567,N_1784,N_4010);
nor U8568 (N_8568,N_2146,N_2932);
or U8569 (N_8569,N_707,N_2786);
nor U8570 (N_8570,N_1627,N_3717);
or U8571 (N_8571,N_4966,N_4917);
or U8572 (N_8572,N_1774,N_2581);
nand U8573 (N_8573,N_2244,N_148);
nand U8574 (N_8574,N_4030,N_4091);
xnor U8575 (N_8575,N_3294,N_4817);
nand U8576 (N_8576,N_4946,N_4296);
xnor U8577 (N_8577,N_4883,N_2043);
nor U8578 (N_8578,N_2092,N_343);
nor U8579 (N_8579,N_190,N_1870);
nand U8580 (N_8580,N_142,N_224);
or U8581 (N_8581,N_3843,N_843);
xnor U8582 (N_8582,N_2134,N_4007);
nor U8583 (N_8583,N_2091,N_4656);
xor U8584 (N_8584,N_4258,N_4452);
nor U8585 (N_8585,N_3468,N_4261);
xnor U8586 (N_8586,N_782,N_2181);
nor U8587 (N_8587,N_3050,N_3480);
xnor U8588 (N_8588,N_3133,N_1521);
and U8589 (N_8589,N_686,N_4383);
or U8590 (N_8590,N_1214,N_2877);
xor U8591 (N_8591,N_598,N_1120);
xnor U8592 (N_8592,N_936,N_3263);
and U8593 (N_8593,N_1293,N_2009);
and U8594 (N_8594,N_3893,N_2427);
nor U8595 (N_8595,N_465,N_958);
nand U8596 (N_8596,N_4720,N_4245);
nor U8597 (N_8597,N_917,N_4601);
xnor U8598 (N_8598,N_3199,N_4911);
and U8599 (N_8599,N_1705,N_406);
and U8600 (N_8600,N_4042,N_4000);
nand U8601 (N_8601,N_1205,N_1030);
or U8602 (N_8602,N_1271,N_1449);
xor U8603 (N_8603,N_2829,N_2918);
nor U8604 (N_8604,N_1867,N_559);
nand U8605 (N_8605,N_933,N_2133);
nor U8606 (N_8606,N_17,N_3615);
nor U8607 (N_8607,N_135,N_228);
and U8608 (N_8608,N_2262,N_4038);
nand U8609 (N_8609,N_2348,N_3074);
xor U8610 (N_8610,N_4714,N_2676);
or U8611 (N_8611,N_4555,N_1146);
nand U8612 (N_8612,N_1718,N_4136);
xnor U8613 (N_8613,N_3962,N_3705);
nor U8614 (N_8614,N_767,N_4150);
or U8615 (N_8615,N_1576,N_2159);
nor U8616 (N_8616,N_4789,N_4748);
nor U8617 (N_8617,N_2248,N_490);
xnor U8618 (N_8618,N_3122,N_666);
xnor U8619 (N_8619,N_2672,N_2957);
and U8620 (N_8620,N_3972,N_1038);
nor U8621 (N_8621,N_2594,N_1757);
nor U8622 (N_8622,N_911,N_4570);
and U8623 (N_8623,N_319,N_2037);
and U8624 (N_8624,N_2838,N_2781);
or U8625 (N_8625,N_869,N_1322);
nand U8626 (N_8626,N_1143,N_3524);
nand U8627 (N_8627,N_1054,N_2949);
and U8628 (N_8628,N_2590,N_63);
xnor U8629 (N_8629,N_4505,N_1874);
xnor U8630 (N_8630,N_3634,N_538);
nand U8631 (N_8631,N_4643,N_2711);
and U8632 (N_8632,N_3676,N_4725);
nor U8633 (N_8633,N_1733,N_854);
xnor U8634 (N_8634,N_383,N_329);
xor U8635 (N_8635,N_1890,N_922);
xnor U8636 (N_8636,N_479,N_2067);
or U8637 (N_8637,N_1046,N_35);
or U8638 (N_8638,N_4705,N_3476);
or U8639 (N_8639,N_456,N_2871);
nor U8640 (N_8640,N_4282,N_1398);
nand U8641 (N_8641,N_3323,N_573);
xor U8642 (N_8642,N_2833,N_614);
nor U8643 (N_8643,N_4305,N_3914);
and U8644 (N_8644,N_1027,N_2762);
nor U8645 (N_8645,N_2646,N_3918);
xnor U8646 (N_8646,N_3619,N_1495);
or U8647 (N_8647,N_2628,N_4009);
and U8648 (N_8648,N_1701,N_3995);
nor U8649 (N_8649,N_4658,N_2600);
and U8650 (N_8650,N_2283,N_4196);
nand U8651 (N_8651,N_3337,N_2895);
xor U8652 (N_8652,N_1494,N_2805);
xnor U8653 (N_8653,N_2661,N_3244);
nand U8654 (N_8654,N_4845,N_4321);
and U8655 (N_8655,N_884,N_4749);
nand U8656 (N_8656,N_3511,N_2007);
xor U8657 (N_8657,N_4648,N_3243);
nand U8658 (N_8658,N_3866,N_3873);
or U8659 (N_8659,N_3644,N_2810);
nor U8660 (N_8660,N_24,N_4016);
and U8661 (N_8661,N_2742,N_3051);
or U8662 (N_8662,N_2648,N_3563);
nand U8663 (N_8663,N_1106,N_33);
or U8664 (N_8664,N_883,N_716);
nand U8665 (N_8665,N_4847,N_1811);
xor U8666 (N_8666,N_3724,N_2841);
xor U8667 (N_8667,N_3499,N_3277);
nor U8668 (N_8668,N_2074,N_4551);
nand U8669 (N_8669,N_1050,N_4853);
or U8670 (N_8670,N_4056,N_4924);
nor U8671 (N_8671,N_1155,N_3579);
or U8672 (N_8672,N_114,N_1492);
nor U8673 (N_8673,N_1741,N_1663);
and U8674 (N_8674,N_805,N_3761);
nor U8675 (N_8675,N_1101,N_4429);
nor U8676 (N_8676,N_964,N_772);
or U8677 (N_8677,N_3052,N_1173);
nand U8678 (N_8678,N_4337,N_4019);
or U8679 (N_8679,N_405,N_4606);
and U8680 (N_8680,N_2298,N_3412);
or U8681 (N_8681,N_4905,N_309);
and U8682 (N_8682,N_2479,N_2848);
xnor U8683 (N_8683,N_1749,N_1156);
and U8684 (N_8684,N_2740,N_2325);
or U8685 (N_8685,N_2980,N_3297);
and U8686 (N_8686,N_2101,N_2703);
and U8687 (N_8687,N_1846,N_3126);
and U8688 (N_8688,N_1497,N_2906);
nand U8689 (N_8689,N_2605,N_4779);
and U8690 (N_8690,N_3877,N_285);
nand U8691 (N_8691,N_1867,N_1316);
and U8692 (N_8692,N_794,N_864);
nand U8693 (N_8693,N_3399,N_1843);
and U8694 (N_8694,N_102,N_557);
xor U8695 (N_8695,N_3504,N_1135);
or U8696 (N_8696,N_3168,N_1022);
and U8697 (N_8697,N_4963,N_2489);
and U8698 (N_8698,N_3891,N_245);
nand U8699 (N_8699,N_1587,N_1259);
xor U8700 (N_8700,N_4835,N_4393);
nand U8701 (N_8701,N_784,N_3021);
nor U8702 (N_8702,N_660,N_3034);
nor U8703 (N_8703,N_224,N_1968);
xor U8704 (N_8704,N_1463,N_411);
xnor U8705 (N_8705,N_2568,N_2919);
xor U8706 (N_8706,N_3201,N_1293);
or U8707 (N_8707,N_1419,N_3084);
and U8708 (N_8708,N_2076,N_3363);
or U8709 (N_8709,N_605,N_4933);
xor U8710 (N_8710,N_1894,N_837);
nor U8711 (N_8711,N_4718,N_2382);
nor U8712 (N_8712,N_931,N_739);
and U8713 (N_8713,N_1047,N_4129);
and U8714 (N_8714,N_2874,N_1346);
nor U8715 (N_8715,N_256,N_4225);
xor U8716 (N_8716,N_3892,N_3439);
nand U8717 (N_8717,N_1618,N_1559);
xor U8718 (N_8718,N_739,N_3733);
nor U8719 (N_8719,N_791,N_4317);
and U8720 (N_8720,N_4380,N_190);
and U8721 (N_8721,N_954,N_1948);
nor U8722 (N_8722,N_3706,N_3406);
nor U8723 (N_8723,N_160,N_3451);
or U8724 (N_8724,N_4149,N_256);
or U8725 (N_8725,N_848,N_2121);
nand U8726 (N_8726,N_3160,N_414);
and U8727 (N_8727,N_2161,N_2853);
nor U8728 (N_8728,N_2697,N_2274);
or U8729 (N_8729,N_579,N_2363);
and U8730 (N_8730,N_1432,N_297);
xnor U8731 (N_8731,N_4683,N_807);
and U8732 (N_8732,N_176,N_13);
or U8733 (N_8733,N_3434,N_690);
xnor U8734 (N_8734,N_1748,N_3447);
and U8735 (N_8735,N_1416,N_3813);
nand U8736 (N_8736,N_1337,N_4409);
xor U8737 (N_8737,N_898,N_1242);
or U8738 (N_8738,N_4842,N_1358);
xnor U8739 (N_8739,N_549,N_3987);
or U8740 (N_8740,N_1116,N_316);
and U8741 (N_8741,N_2168,N_3604);
nor U8742 (N_8742,N_4675,N_1137);
xnor U8743 (N_8743,N_1079,N_4619);
or U8744 (N_8744,N_2914,N_4752);
and U8745 (N_8745,N_2962,N_4414);
and U8746 (N_8746,N_3390,N_4482);
nor U8747 (N_8747,N_2521,N_1690);
xnor U8748 (N_8748,N_739,N_2499);
and U8749 (N_8749,N_377,N_2773);
nand U8750 (N_8750,N_4559,N_589);
xor U8751 (N_8751,N_1022,N_1975);
xor U8752 (N_8752,N_2167,N_4014);
xor U8753 (N_8753,N_2969,N_4264);
xnor U8754 (N_8754,N_1547,N_1813);
and U8755 (N_8755,N_1978,N_2298);
or U8756 (N_8756,N_1199,N_4014);
and U8757 (N_8757,N_603,N_3448);
nand U8758 (N_8758,N_836,N_808);
and U8759 (N_8759,N_1504,N_2086);
nand U8760 (N_8760,N_3454,N_4534);
nor U8761 (N_8761,N_2657,N_4922);
or U8762 (N_8762,N_4178,N_1592);
or U8763 (N_8763,N_2811,N_740);
nor U8764 (N_8764,N_4234,N_1354);
nand U8765 (N_8765,N_1828,N_337);
nand U8766 (N_8766,N_1589,N_3818);
nand U8767 (N_8767,N_1394,N_2098);
nor U8768 (N_8768,N_3772,N_2131);
xnor U8769 (N_8769,N_4936,N_4016);
and U8770 (N_8770,N_418,N_4057);
xnor U8771 (N_8771,N_3867,N_1342);
or U8772 (N_8772,N_4829,N_10);
or U8773 (N_8773,N_1365,N_3653);
and U8774 (N_8774,N_3399,N_4242);
nand U8775 (N_8775,N_3614,N_1425);
nand U8776 (N_8776,N_3494,N_3968);
nand U8777 (N_8777,N_4793,N_1766);
and U8778 (N_8778,N_1097,N_1681);
or U8779 (N_8779,N_3784,N_2863);
or U8780 (N_8780,N_3069,N_1113);
or U8781 (N_8781,N_1212,N_275);
or U8782 (N_8782,N_4135,N_2975);
or U8783 (N_8783,N_1508,N_4874);
and U8784 (N_8784,N_408,N_2412);
and U8785 (N_8785,N_2501,N_4841);
nor U8786 (N_8786,N_4929,N_2580);
nand U8787 (N_8787,N_2799,N_1587);
xnor U8788 (N_8788,N_4557,N_1117);
nand U8789 (N_8789,N_3797,N_608);
nand U8790 (N_8790,N_483,N_2854);
nor U8791 (N_8791,N_3289,N_2335);
nor U8792 (N_8792,N_2119,N_611);
and U8793 (N_8793,N_421,N_2466);
nor U8794 (N_8794,N_2572,N_463);
or U8795 (N_8795,N_3904,N_605);
xor U8796 (N_8796,N_1676,N_2624);
or U8797 (N_8797,N_4394,N_4258);
nand U8798 (N_8798,N_4247,N_69);
and U8799 (N_8799,N_365,N_4726);
nand U8800 (N_8800,N_4184,N_65);
or U8801 (N_8801,N_1928,N_2310);
nand U8802 (N_8802,N_1277,N_2727);
or U8803 (N_8803,N_4195,N_3303);
nand U8804 (N_8804,N_3412,N_1887);
and U8805 (N_8805,N_3650,N_2802);
and U8806 (N_8806,N_3989,N_1495);
or U8807 (N_8807,N_4878,N_1606);
nand U8808 (N_8808,N_22,N_564);
and U8809 (N_8809,N_988,N_877);
nor U8810 (N_8810,N_2817,N_3594);
and U8811 (N_8811,N_712,N_44);
nor U8812 (N_8812,N_2902,N_1713);
nand U8813 (N_8813,N_4021,N_4556);
xor U8814 (N_8814,N_2174,N_2526);
or U8815 (N_8815,N_2753,N_2732);
xor U8816 (N_8816,N_1160,N_4543);
or U8817 (N_8817,N_901,N_2895);
nand U8818 (N_8818,N_4230,N_2013);
or U8819 (N_8819,N_1049,N_2627);
nor U8820 (N_8820,N_898,N_2746);
xor U8821 (N_8821,N_1614,N_3355);
nand U8822 (N_8822,N_190,N_2052);
nand U8823 (N_8823,N_747,N_3607);
nand U8824 (N_8824,N_4839,N_1673);
xor U8825 (N_8825,N_984,N_4931);
nand U8826 (N_8826,N_4519,N_666);
or U8827 (N_8827,N_3719,N_3782);
xor U8828 (N_8828,N_2718,N_214);
nand U8829 (N_8829,N_402,N_1037);
and U8830 (N_8830,N_2144,N_1137);
and U8831 (N_8831,N_4992,N_2538);
and U8832 (N_8832,N_1304,N_3832);
and U8833 (N_8833,N_2904,N_407);
nand U8834 (N_8834,N_4419,N_1560);
xor U8835 (N_8835,N_3143,N_276);
xnor U8836 (N_8836,N_2419,N_720);
or U8837 (N_8837,N_3605,N_2005);
and U8838 (N_8838,N_2208,N_297);
and U8839 (N_8839,N_2946,N_3444);
nor U8840 (N_8840,N_531,N_1138);
xnor U8841 (N_8841,N_2719,N_2933);
nand U8842 (N_8842,N_3799,N_4965);
or U8843 (N_8843,N_1519,N_4275);
nor U8844 (N_8844,N_2280,N_1493);
nor U8845 (N_8845,N_167,N_2506);
and U8846 (N_8846,N_857,N_480);
xor U8847 (N_8847,N_226,N_4472);
xnor U8848 (N_8848,N_4917,N_1052);
or U8849 (N_8849,N_1619,N_4768);
and U8850 (N_8850,N_2942,N_1834);
nor U8851 (N_8851,N_3033,N_3921);
or U8852 (N_8852,N_3931,N_165);
or U8853 (N_8853,N_3886,N_4408);
nand U8854 (N_8854,N_1106,N_4659);
and U8855 (N_8855,N_4319,N_3599);
nand U8856 (N_8856,N_2960,N_844);
and U8857 (N_8857,N_3756,N_2848);
or U8858 (N_8858,N_3993,N_389);
and U8859 (N_8859,N_4521,N_532);
nor U8860 (N_8860,N_86,N_553);
xor U8861 (N_8861,N_3324,N_4811);
and U8862 (N_8862,N_629,N_2915);
nand U8863 (N_8863,N_389,N_1449);
nand U8864 (N_8864,N_1483,N_2455);
and U8865 (N_8865,N_1591,N_1823);
and U8866 (N_8866,N_2422,N_4945);
and U8867 (N_8867,N_1425,N_4889);
nor U8868 (N_8868,N_4660,N_3122);
and U8869 (N_8869,N_807,N_781);
xor U8870 (N_8870,N_1310,N_1089);
and U8871 (N_8871,N_824,N_3792);
nand U8872 (N_8872,N_2151,N_3939);
and U8873 (N_8873,N_4729,N_4012);
nand U8874 (N_8874,N_3672,N_263);
or U8875 (N_8875,N_4983,N_1502);
nand U8876 (N_8876,N_2145,N_3805);
and U8877 (N_8877,N_2739,N_160);
and U8878 (N_8878,N_475,N_3752);
and U8879 (N_8879,N_3457,N_980);
or U8880 (N_8880,N_3881,N_1071);
or U8881 (N_8881,N_673,N_4298);
or U8882 (N_8882,N_3528,N_1009);
nor U8883 (N_8883,N_1084,N_3780);
nand U8884 (N_8884,N_1140,N_249);
and U8885 (N_8885,N_2196,N_2214);
nor U8886 (N_8886,N_4511,N_2902);
nor U8887 (N_8887,N_4989,N_223);
xnor U8888 (N_8888,N_4908,N_2280);
and U8889 (N_8889,N_3674,N_3051);
nand U8890 (N_8890,N_209,N_4482);
or U8891 (N_8891,N_3697,N_1886);
xor U8892 (N_8892,N_4924,N_1122);
xor U8893 (N_8893,N_4677,N_4884);
xnor U8894 (N_8894,N_1428,N_81);
or U8895 (N_8895,N_3900,N_2852);
nor U8896 (N_8896,N_3626,N_4793);
nand U8897 (N_8897,N_502,N_4347);
and U8898 (N_8898,N_3438,N_70);
xnor U8899 (N_8899,N_2647,N_1803);
or U8900 (N_8900,N_628,N_2790);
nand U8901 (N_8901,N_4006,N_1228);
or U8902 (N_8902,N_2012,N_1695);
nor U8903 (N_8903,N_2448,N_4083);
and U8904 (N_8904,N_3913,N_1615);
nand U8905 (N_8905,N_3930,N_3501);
nand U8906 (N_8906,N_1705,N_2800);
and U8907 (N_8907,N_2000,N_4736);
or U8908 (N_8908,N_389,N_2747);
or U8909 (N_8909,N_4199,N_83);
xor U8910 (N_8910,N_3504,N_3381);
xnor U8911 (N_8911,N_156,N_2065);
nor U8912 (N_8912,N_1128,N_3011);
and U8913 (N_8913,N_1770,N_4120);
and U8914 (N_8914,N_2392,N_264);
and U8915 (N_8915,N_383,N_1419);
and U8916 (N_8916,N_321,N_1700);
and U8917 (N_8917,N_2585,N_119);
xor U8918 (N_8918,N_2380,N_2097);
nor U8919 (N_8919,N_3529,N_3422);
xor U8920 (N_8920,N_146,N_2376);
or U8921 (N_8921,N_4250,N_1318);
or U8922 (N_8922,N_4023,N_3770);
nand U8923 (N_8923,N_4021,N_4549);
xnor U8924 (N_8924,N_1783,N_303);
or U8925 (N_8925,N_3723,N_1382);
nor U8926 (N_8926,N_1385,N_2402);
or U8927 (N_8927,N_3920,N_3222);
and U8928 (N_8928,N_304,N_734);
xnor U8929 (N_8929,N_4199,N_2953);
nand U8930 (N_8930,N_3708,N_2533);
xor U8931 (N_8931,N_4782,N_3467);
or U8932 (N_8932,N_688,N_2843);
and U8933 (N_8933,N_689,N_1487);
nand U8934 (N_8934,N_1578,N_1943);
nand U8935 (N_8935,N_3956,N_2056);
xnor U8936 (N_8936,N_4460,N_1009);
nand U8937 (N_8937,N_485,N_2373);
xor U8938 (N_8938,N_1428,N_3286);
and U8939 (N_8939,N_542,N_4653);
and U8940 (N_8940,N_2844,N_361);
nor U8941 (N_8941,N_2937,N_3879);
xor U8942 (N_8942,N_2182,N_4418);
nor U8943 (N_8943,N_4802,N_1407);
and U8944 (N_8944,N_642,N_3939);
nand U8945 (N_8945,N_3558,N_4418);
or U8946 (N_8946,N_3803,N_4807);
nand U8947 (N_8947,N_388,N_1540);
nor U8948 (N_8948,N_1917,N_4528);
nor U8949 (N_8949,N_3740,N_1326);
and U8950 (N_8950,N_4282,N_2734);
nor U8951 (N_8951,N_3147,N_4378);
xor U8952 (N_8952,N_434,N_290);
xor U8953 (N_8953,N_3782,N_2714);
and U8954 (N_8954,N_4892,N_2491);
and U8955 (N_8955,N_4256,N_4907);
or U8956 (N_8956,N_3465,N_1310);
nor U8957 (N_8957,N_2376,N_3424);
or U8958 (N_8958,N_2377,N_3351);
and U8959 (N_8959,N_1667,N_837);
nor U8960 (N_8960,N_4819,N_4438);
xor U8961 (N_8961,N_2869,N_1810);
nand U8962 (N_8962,N_1456,N_4683);
xnor U8963 (N_8963,N_642,N_4141);
nand U8964 (N_8964,N_4875,N_1876);
xor U8965 (N_8965,N_3445,N_1883);
xnor U8966 (N_8966,N_2741,N_3663);
nand U8967 (N_8967,N_4192,N_1624);
nand U8968 (N_8968,N_816,N_1832);
xnor U8969 (N_8969,N_1914,N_3427);
and U8970 (N_8970,N_1350,N_920);
and U8971 (N_8971,N_801,N_1417);
xor U8972 (N_8972,N_3212,N_2790);
and U8973 (N_8973,N_4046,N_538);
nand U8974 (N_8974,N_4709,N_2727);
xor U8975 (N_8975,N_143,N_3149);
xor U8976 (N_8976,N_4430,N_784);
or U8977 (N_8977,N_4369,N_351);
nor U8978 (N_8978,N_749,N_1352);
nor U8979 (N_8979,N_274,N_4643);
nand U8980 (N_8980,N_2890,N_2998);
or U8981 (N_8981,N_1894,N_4067);
and U8982 (N_8982,N_1642,N_3210);
nand U8983 (N_8983,N_2244,N_3650);
and U8984 (N_8984,N_1264,N_135);
nor U8985 (N_8985,N_4364,N_1399);
nor U8986 (N_8986,N_574,N_1826);
nand U8987 (N_8987,N_3444,N_1602);
or U8988 (N_8988,N_2532,N_1502);
and U8989 (N_8989,N_2984,N_982);
or U8990 (N_8990,N_3868,N_390);
and U8991 (N_8991,N_29,N_2340);
xnor U8992 (N_8992,N_486,N_3052);
nand U8993 (N_8993,N_139,N_4412);
and U8994 (N_8994,N_4840,N_2862);
xnor U8995 (N_8995,N_3618,N_708);
or U8996 (N_8996,N_2,N_3659);
and U8997 (N_8997,N_323,N_1356);
nand U8998 (N_8998,N_2323,N_2795);
nand U8999 (N_8999,N_736,N_730);
and U9000 (N_9000,N_1483,N_240);
or U9001 (N_9001,N_4797,N_1333);
nand U9002 (N_9002,N_4165,N_3541);
nor U9003 (N_9003,N_3061,N_465);
nor U9004 (N_9004,N_2617,N_4976);
nand U9005 (N_9005,N_2641,N_87);
nor U9006 (N_9006,N_1230,N_3234);
xor U9007 (N_9007,N_2941,N_3435);
nor U9008 (N_9008,N_1886,N_1201);
or U9009 (N_9009,N_4457,N_1969);
and U9010 (N_9010,N_1222,N_2160);
and U9011 (N_9011,N_4061,N_651);
or U9012 (N_9012,N_1188,N_2861);
xor U9013 (N_9013,N_1021,N_2828);
and U9014 (N_9014,N_2828,N_496);
and U9015 (N_9015,N_4836,N_1484);
nand U9016 (N_9016,N_3542,N_109);
xor U9017 (N_9017,N_2061,N_3137);
nor U9018 (N_9018,N_3488,N_2171);
or U9019 (N_9019,N_2197,N_2553);
nor U9020 (N_9020,N_2770,N_870);
nor U9021 (N_9021,N_1999,N_4999);
nor U9022 (N_9022,N_1883,N_3538);
nor U9023 (N_9023,N_1073,N_1410);
and U9024 (N_9024,N_4623,N_822);
nor U9025 (N_9025,N_4366,N_2144);
and U9026 (N_9026,N_1112,N_430);
and U9027 (N_9027,N_2338,N_3441);
nor U9028 (N_9028,N_74,N_3545);
or U9029 (N_9029,N_4056,N_2312);
nor U9030 (N_9030,N_16,N_21);
or U9031 (N_9031,N_897,N_3969);
xor U9032 (N_9032,N_3901,N_4810);
or U9033 (N_9033,N_2451,N_2827);
xnor U9034 (N_9034,N_707,N_659);
and U9035 (N_9035,N_4395,N_4592);
nand U9036 (N_9036,N_2851,N_2554);
nor U9037 (N_9037,N_1221,N_1752);
or U9038 (N_9038,N_1731,N_4586);
or U9039 (N_9039,N_3557,N_4641);
xor U9040 (N_9040,N_595,N_1156);
nor U9041 (N_9041,N_4903,N_4657);
or U9042 (N_9042,N_256,N_2627);
or U9043 (N_9043,N_3937,N_4669);
or U9044 (N_9044,N_181,N_4268);
nand U9045 (N_9045,N_2735,N_1006);
xnor U9046 (N_9046,N_3930,N_3343);
and U9047 (N_9047,N_1717,N_4232);
or U9048 (N_9048,N_1448,N_2686);
nand U9049 (N_9049,N_1420,N_1106);
xor U9050 (N_9050,N_3443,N_3644);
or U9051 (N_9051,N_1341,N_4062);
xor U9052 (N_9052,N_1009,N_541);
or U9053 (N_9053,N_4022,N_959);
nor U9054 (N_9054,N_3240,N_584);
nand U9055 (N_9055,N_1307,N_3338);
or U9056 (N_9056,N_432,N_769);
and U9057 (N_9057,N_203,N_338);
nor U9058 (N_9058,N_3556,N_1803);
and U9059 (N_9059,N_606,N_3111);
and U9060 (N_9060,N_1588,N_3028);
nor U9061 (N_9061,N_3162,N_4671);
nand U9062 (N_9062,N_1448,N_2769);
or U9063 (N_9063,N_1820,N_4714);
and U9064 (N_9064,N_4495,N_14);
xnor U9065 (N_9065,N_4941,N_1100);
nand U9066 (N_9066,N_1333,N_4782);
or U9067 (N_9067,N_4622,N_767);
nor U9068 (N_9068,N_2914,N_1918);
and U9069 (N_9069,N_3119,N_423);
or U9070 (N_9070,N_2489,N_2929);
and U9071 (N_9071,N_2732,N_4792);
xor U9072 (N_9072,N_1346,N_2036);
nor U9073 (N_9073,N_3582,N_4687);
nor U9074 (N_9074,N_3306,N_3532);
nor U9075 (N_9075,N_316,N_4840);
and U9076 (N_9076,N_4535,N_4997);
nand U9077 (N_9077,N_3360,N_4651);
xor U9078 (N_9078,N_1039,N_1998);
xnor U9079 (N_9079,N_4626,N_2979);
and U9080 (N_9080,N_1532,N_3175);
nand U9081 (N_9081,N_2627,N_648);
nor U9082 (N_9082,N_1544,N_1110);
nand U9083 (N_9083,N_4590,N_2607);
and U9084 (N_9084,N_4910,N_3695);
and U9085 (N_9085,N_472,N_2657);
or U9086 (N_9086,N_3350,N_3794);
nor U9087 (N_9087,N_2551,N_974);
or U9088 (N_9088,N_2478,N_2966);
nor U9089 (N_9089,N_2518,N_3792);
xnor U9090 (N_9090,N_613,N_115);
nor U9091 (N_9091,N_2577,N_3767);
xor U9092 (N_9092,N_1046,N_3795);
nor U9093 (N_9093,N_3784,N_1824);
and U9094 (N_9094,N_1312,N_715);
nand U9095 (N_9095,N_3600,N_3633);
nor U9096 (N_9096,N_3934,N_1118);
xnor U9097 (N_9097,N_2408,N_559);
and U9098 (N_9098,N_4454,N_2649);
nand U9099 (N_9099,N_1490,N_3843);
nand U9100 (N_9100,N_4090,N_2124);
nand U9101 (N_9101,N_2920,N_1181);
and U9102 (N_9102,N_1103,N_2858);
xnor U9103 (N_9103,N_349,N_718);
nor U9104 (N_9104,N_2265,N_316);
and U9105 (N_9105,N_4197,N_2511);
xor U9106 (N_9106,N_4251,N_1793);
xor U9107 (N_9107,N_929,N_4050);
and U9108 (N_9108,N_2543,N_2414);
and U9109 (N_9109,N_1110,N_1989);
xor U9110 (N_9110,N_1885,N_1632);
nor U9111 (N_9111,N_4741,N_4105);
nand U9112 (N_9112,N_4518,N_3348);
xnor U9113 (N_9113,N_3609,N_2564);
and U9114 (N_9114,N_3860,N_2478);
or U9115 (N_9115,N_2790,N_2191);
xor U9116 (N_9116,N_2327,N_256);
nand U9117 (N_9117,N_3965,N_4030);
nand U9118 (N_9118,N_1706,N_4700);
xnor U9119 (N_9119,N_3180,N_1584);
nand U9120 (N_9120,N_4622,N_369);
xor U9121 (N_9121,N_1453,N_4459);
xor U9122 (N_9122,N_2778,N_820);
xor U9123 (N_9123,N_1492,N_4800);
or U9124 (N_9124,N_1007,N_817);
and U9125 (N_9125,N_2297,N_874);
nand U9126 (N_9126,N_3186,N_4390);
xor U9127 (N_9127,N_663,N_4008);
or U9128 (N_9128,N_1754,N_2870);
and U9129 (N_9129,N_1360,N_2566);
xnor U9130 (N_9130,N_626,N_3375);
and U9131 (N_9131,N_1422,N_1934);
and U9132 (N_9132,N_1623,N_703);
and U9133 (N_9133,N_4285,N_1374);
or U9134 (N_9134,N_832,N_3885);
and U9135 (N_9135,N_3158,N_2429);
or U9136 (N_9136,N_4502,N_1735);
and U9137 (N_9137,N_2390,N_654);
nand U9138 (N_9138,N_1230,N_4384);
nor U9139 (N_9139,N_343,N_3309);
nand U9140 (N_9140,N_3419,N_4060);
and U9141 (N_9141,N_17,N_1627);
xnor U9142 (N_9142,N_542,N_1603);
and U9143 (N_9143,N_4320,N_1876);
nor U9144 (N_9144,N_634,N_812);
nor U9145 (N_9145,N_477,N_172);
xor U9146 (N_9146,N_3570,N_2470);
nand U9147 (N_9147,N_1961,N_677);
xor U9148 (N_9148,N_1254,N_1783);
nor U9149 (N_9149,N_4920,N_4888);
or U9150 (N_9150,N_3940,N_520);
xnor U9151 (N_9151,N_2417,N_2359);
and U9152 (N_9152,N_2623,N_1260);
nor U9153 (N_9153,N_249,N_4916);
or U9154 (N_9154,N_569,N_2651);
or U9155 (N_9155,N_2256,N_3789);
nand U9156 (N_9156,N_4795,N_4005);
nand U9157 (N_9157,N_4719,N_4042);
nand U9158 (N_9158,N_3533,N_1400);
or U9159 (N_9159,N_3790,N_116);
nand U9160 (N_9160,N_4250,N_46);
or U9161 (N_9161,N_4892,N_3842);
nand U9162 (N_9162,N_4718,N_863);
xnor U9163 (N_9163,N_1950,N_3751);
or U9164 (N_9164,N_3688,N_3293);
and U9165 (N_9165,N_2313,N_2108);
xnor U9166 (N_9166,N_1041,N_1212);
or U9167 (N_9167,N_3769,N_342);
xor U9168 (N_9168,N_3230,N_3491);
xnor U9169 (N_9169,N_4552,N_2588);
and U9170 (N_9170,N_1609,N_2255);
nor U9171 (N_9171,N_2306,N_3986);
and U9172 (N_9172,N_2770,N_2794);
xnor U9173 (N_9173,N_2865,N_3540);
and U9174 (N_9174,N_3537,N_2381);
xor U9175 (N_9175,N_3448,N_1055);
xnor U9176 (N_9176,N_993,N_2908);
and U9177 (N_9177,N_3949,N_566);
or U9178 (N_9178,N_1364,N_333);
nand U9179 (N_9179,N_2904,N_896);
nand U9180 (N_9180,N_2456,N_4800);
nand U9181 (N_9181,N_345,N_987);
or U9182 (N_9182,N_1604,N_3369);
nand U9183 (N_9183,N_1081,N_648);
or U9184 (N_9184,N_4215,N_2752);
or U9185 (N_9185,N_4631,N_32);
nand U9186 (N_9186,N_4486,N_1567);
nor U9187 (N_9187,N_1099,N_3417);
nor U9188 (N_9188,N_2103,N_2133);
nand U9189 (N_9189,N_1517,N_3853);
nor U9190 (N_9190,N_1606,N_3577);
or U9191 (N_9191,N_637,N_1064);
or U9192 (N_9192,N_1093,N_1762);
or U9193 (N_9193,N_999,N_1988);
and U9194 (N_9194,N_4768,N_3478);
or U9195 (N_9195,N_1164,N_2225);
xor U9196 (N_9196,N_19,N_102);
nor U9197 (N_9197,N_2169,N_1549);
nand U9198 (N_9198,N_1678,N_4165);
nor U9199 (N_9199,N_791,N_3825);
nand U9200 (N_9200,N_1684,N_1381);
and U9201 (N_9201,N_349,N_1362);
nor U9202 (N_9202,N_2880,N_2169);
xor U9203 (N_9203,N_3525,N_1043);
and U9204 (N_9204,N_2031,N_3431);
or U9205 (N_9205,N_341,N_4859);
or U9206 (N_9206,N_2591,N_3555);
xnor U9207 (N_9207,N_4112,N_3567);
or U9208 (N_9208,N_4623,N_4035);
and U9209 (N_9209,N_4280,N_3418);
and U9210 (N_9210,N_4672,N_851);
nor U9211 (N_9211,N_2581,N_995);
nor U9212 (N_9212,N_3421,N_785);
and U9213 (N_9213,N_409,N_1174);
nor U9214 (N_9214,N_1024,N_266);
and U9215 (N_9215,N_1130,N_3633);
and U9216 (N_9216,N_663,N_4365);
nor U9217 (N_9217,N_1044,N_591);
or U9218 (N_9218,N_1091,N_2828);
and U9219 (N_9219,N_2526,N_3759);
and U9220 (N_9220,N_2843,N_2258);
nor U9221 (N_9221,N_2609,N_655);
or U9222 (N_9222,N_1409,N_4874);
xor U9223 (N_9223,N_353,N_1245);
nor U9224 (N_9224,N_1756,N_4395);
xnor U9225 (N_9225,N_646,N_2014);
nor U9226 (N_9226,N_3075,N_1480);
and U9227 (N_9227,N_1504,N_1677);
nor U9228 (N_9228,N_1411,N_4819);
nor U9229 (N_9229,N_2756,N_1496);
nor U9230 (N_9230,N_4610,N_2992);
or U9231 (N_9231,N_447,N_94);
and U9232 (N_9232,N_1548,N_629);
nand U9233 (N_9233,N_297,N_2953);
nor U9234 (N_9234,N_1132,N_3835);
or U9235 (N_9235,N_4072,N_1025);
nand U9236 (N_9236,N_674,N_69);
nor U9237 (N_9237,N_1338,N_548);
and U9238 (N_9238,N_2846,N_1968);
xnor U9239 (N_9239,N_2451,N_3617);
nand U9240 (N_9240,N_2405,N_3679);
nor U9241 (N_9241,N_2271,N_508);
and U9242 (N_9242,N_428,N_1257);
xor U9243 (N_9243,N_2469,N_1808);
nor U9244 (N_9244,N_2726,N_2018);
or U9245 (N_9245,N_151,N_3443);
and U9246 (N_9246,N_15,N_3015);
and U9247 (N_9247,N_711,N_4734);
and U9248 (N_9248,N_4553,N_1373);
nor U9249 (N_9249,N_1239,N_3715);
and U9250 (N_9250,N_1686,N_4794);
nor U9251 (N_9251,N_1006,N_3992);
and U9252 (N_9252,N_2306,N_2560);
xor U9253 (N_9253,N_322,N_1348);
xnor U9254 (N_9254,N_4000,N_889);
nor U9255 (N_9255,N_3783,N_3104);
nor U9256 (N_9256,N_2628,N_3559);
and U9257 (N_9257,N_3899,N_1247);
or U9258 (N_9258,N_1671,N_1580);
and U9259 (N_9259,N_1281,N_4105);
nand U9260 (N_9260,N_3289,N_903);
and U9261 (N_9261,N_2089,N_2015);
nand U9262 (N_9262,N_444,N_4726);
or U9263 (N_9263,N_3678,N_788);
and U9264 (N_9264,N_4627,N_2221);
or U9265 (N_9265,N_3919,N_3528);
nor U9266 (N_9266,N_2465,N_1628);
xnor U9267 (N_9267,N_683,N_3648);
xnor U9268 (N_9268,N_4959,N_1509);
nand U9269 (N_9269,N_653,N_1068);
nand U9270 (N_9270,N_1657,N_1675);
nor U9271 (N_9271,N_1434,N_3283);
nor U9272 (N_9272,N_4134,N_4806);
and U9273 (N_9273,N_4290,N_52);
and U9274 (N_9274,N_1250,N_423);
xnor U9275 (N_9275,N_4944,N_1619);
xor U9276 (N_9276,N_4435,N_4932);
xor U9277 (N_9277,N_4647,N_3075);
xnor U9278 (N_9278,N_1750,N_3590);
xnor U9279 (N_9279,N_320,N_2258);
nor U9280 (N_9280,N_4342,N_2239);
or U9281 (N_9281,N_801,N_2278);
nor U9282 (N_9282,N_1504,N_2875);
nor U9283 (N_9283,N_1897,N_41);
nor U9284 (N_9284,N_696,N_1475);
nor U9285 (N_9285,N_2398,N_4871);
nand U9286 (N_9286,N_4870,N_3469);
and U9287 (N_9287,N_4738,N_146);
nor U9288 (N_9288,N_2819,N_4051);
nor U9289 (N_9289,N_2998,N_1270);
and U9290 (N_9290,N_1532,N_1889);
xor U9291 (N_9291,N_4879,N_229);
nand U9292 (N_9292,N_3752,N_1589);
nor U9293 (N_9293,N_2764,N_3205);
or U9294 (N_9294,N_2412,N_1912);
or U9295 (N_9295,N_4245,N_71);
or U9296 (N_9296,N_4631,N_3630);
xnor U9297 (N_9297,N_1939,N_3266);
and U9298 (N_9298,N_4598,N_3506);
nor U9299 (N_9299,N_2006,N_4181);
or U9300 (N_9300,N_3580,N_174);
nand U9301 (N_9301,N_468,N_108);
xnor U9302 (N_9302,N_959,N_889);
and U9303 (N_9303,N_225,N_4387);
xor U9304 (N_9304,N_3756,N_3570);
and U9305 (N_9305,N_3840,N_3460);
xor U9306 (N_9306,N_4221,N_3716);
nor U9307 (N_9307,N_4810,N_3940);
xnor U9308 (N_9308,N_4131,N_2271);
xnor U9309 (N_9309,N_4093,N_3012);
or U9310 (N_9310,N_1244,N_727);
xor U9311 (N_9311,N_1136,N_99);
nor U9312 (N_9312,N_451,N_3878);
nor U9313 (N_9313,N_4345,N_1477);
xor U9314 (N_9314,N_3009,N_3270);
nor U9315 (N_9315,N_26,N_4469);
xnor U9316 (N_9316,N_3324,N_2855);
nor U9317 (N_9317,N_1932,N_415);
nand U9318 (N_9318,N_1361,N_404);
nor U9319 (N_9319,N_2379,N_2913);
nor U9320 (N_9320,N_4572,N_8);
xnor U9321 (N_9321,N_3128,N_4060);
and U9322 (N_9322,N_1083,N_3059);
or U9323 (N_9323,N_4296,N_2909);
xor U9324 (N_9324,N_4514,N_2135);
nor U9325 (N_9325,N_3403,N_4375);
or U9326 (N_9326,N_201,N_2440);
and U9327 (N_9327,N_3972,N_793);
and U9328 (N_9328,N_1792,N_4619);
or U9329 (N_9329,N_1722,N_4177);
xor U9330 (N_9330,N_511,N_4633);
xnor U9331 (N_9331,N_2385,N_710);
or U9332 (N_9332,N_3951,N_2509);
nand U9333 (N_9333,N_2520,N_3625);
nor U9334 (N_9334,N_2306,N_290);
nand U9335 (N_9335,N_4356,N_4441);
or U9336 (N_9336,N_2921,N_3948);
or U9337 (N_9337,N_3206,N_2778);
and U9338 (N_9338,N_4575,N_2244);
or U9339 (N_9339,N_3168,N_1795);
nand U9340 (N_9340,N_1100,N_1322);
nor U9341 (N_9341,N_3304,N_3398);
and U9342 (N_9342,N_4638,N_1081);
nor U9343 (N_9343,N_755,N_4823);
nor U9344 (N_9344,N_2579,N_1068);
nand U9345 (N_9345,N_2516,N_2631);
or U9346 (N_9346,N_1227,N_382);
nor U9347 (N_9347,N_1178,N_78);
or U9348 (N_9348,N_643,N_4745);
and U9349 (N_9349,N_1205,N_2989);
nor U9350 (N_9350,N_427,N_4004);
and U9351 (N_9351,N_2375,N_3463);
nor U9352 (N_9352,N_4622,N_1022);
xnor U9353 (N_9353,N_729,N_2653);
xnor U9354 (N_9354,N_3432,N_2665);
nor U9355 (N_9355,N_4724,N_2928);
xnor U9356 (N_9356,N_874,N_1866);
and U9357 (N_9357,N_4156,N_3618);
nor U9358 (N_9358,N_1562,N_609);
xor U9359 (N_9359,N_491,N_4993);
and U9360 (N_9360,N_212,N_3669);
or U9361 (N_9361,N_4874,N_3887);
nor U9362 (N_9362,N_168,N_713);
or U9363 (N_9363,N_1730,N_2227);
and U9364 (N_9364,N_3990,N_2886);
and U9365 (N_9365,N_3486,N_1875);
and U9366 (N_9366,N_3221,N_1195);
nor U9367 (N_9367,N_1724,N_3244);
or U9368 (N_9368,N_2494,N_3054);
xnor U9369 (N_9369,N_3691,N_2649);
nor U9370 (N_9370,N_2685,N_3065);
xnor U9371 (N_9371,N_3597,N_2124);
nand U9372 (N_9372,N_1954,N_3499);
and U9373 (N_9373,N_1973,N_1447);
nand U9374 (N_9374,N_1433,N_4707);
nor U9375 (N_9375,N_2014,N_1378);
xnor U9376 (N_9376,N_1469,N_4351);
or U9377 (N_9377,N_4922,N_2502);
xor U9378 (N_9378,N_2600,N_2499);
and U9379 (N_9379,N_366,N_2579);
nand U9380 (N_9380,N_255,N_344);
nor U9381 (N_9381,N_2845,N_2774);
and U9382 (N_9382,N_2868,N_2044);
xnor U9383 (N_9383,N_4570,N_227);
or U9384 (N_9384,N_156,N_1220);
nor U9385 (N_9385,N_211,N_4949);
or U9386 (N_9386,N_1597,N_1647);
or U9387 (N_9387,N_509,N_3667);
nand U9388 (N_9388,N_3226,N_2079);
and U9389 (N_9389,N_4056,N_2302);
or U9390 (N_9390,N_660,N_4888);
and U9391 (N_9391,N_2314,N_1432);
xnor U9392 (N_9392,N_1170,N_4832);
and U9393 (N_9393,N_838,N_1292);
xor U9394 (N_9394,N_2795,N_1154);
and U9395 (N_9395,N_204,N_4879);
nand U9396 (N_9396,N_4906,N_958);
nand U9397 (N_9397,N_3153,N_2323);
xor U9398 (N_9398,N_1734,N_2031);
xor U9399 (N_9399,N_772,N_595);
xnor U9400 (N_9400,N_4135,N_379);
and U9401 (N_9401,N_3747,N_1863);
and U9402 (N_9402,N_4403,N_2102);
and U9403 (N_9403,N_36,N_646);
xor U9404 (N_9404,N_792,N_3242);
nor U9405 (N_9405,N_3773,N_4224);
nand U9406 (N_9406,N_613,N_2297);
and U9407 (N_9407,N_4698,N_1698);
nand U9408 (N_9408,N_1293,N_3876);
nand U9409 (N_9409,N_2236,N_3874);
xnor U9410 (N_9410,N_942,N_995);
and U9411 (N_9411,N_1199,N_3080);
or U9412 (N_9412,N_1329,N_1062);
xnor U9413 (N_9413,N_4579,N_4682);
xor U9414 (N_9414,N_1498,N_3261);
or U9415 (N_9415,N_3073,N_371);
and U9416 (N_9416,N_2995,N_2619);
xnor U9417 (N_9417,N_4519,N_2619);
xnor U9418 (N_9418,N_4652,N_1578);
or U9419 (N_9419,N_1980,N_3367);
and U9420 (N_9420,N_4262,N_2048);
xnor U9421 (N_9421,N_51,N_4801);
nor U9422 (N_9422,N_3691,N_1565);
nor U9423 (N_9423,N_2253,N_4585);
nand U9424 (N_9424,N_3327,N_2164);
nor U9425 (N_9425,N_3856,N_4598);
or U9426 (N_9426,N_3706,N_4399);
and U9427 (N_9427,N_2418,N_4073);
nor U9428 (N_9428,N_1264,N_290);
nand U9429 (N_9429,N_3258,N_2775);
xnor U9430 (N_9430,N_1512,N_4186);
nand U9431 (N_9431,N_1525,N_1463);
xor U9432 (N_9432,N_1075,N_534);
xor U9433 (N_9433,N_2835,N_155);
nor U9434 (N_9434,N_2034,N_3650);
or U9435 (N_9435,N_2437,N_388);
nor U9436 (N_9436,N_2908,N_589);
nand U9437 (N_9437,N_2707,N_951);
and U9438 (N_9438,N_4954,N_2777);
xor U9439 (N_9439,N_2,N_2496);
nor U9440 (N_9440,N_3757,N_1967);
or U9441 (N_9441,N_3836,N_4487);
nor U9442 (N_9442,N_2111,N_2057);
nor U9443 (N_9443,N_1164,N_4870);
nor U9444 (N_9444,N_3580,N_852);
nand U9445 (N_9445,N_3459,N_1172);
or U9446 (N_9446,N_547,N_1686);
and U9447 (N_9447,N_4009,N_3753);
nand U9448 (N_9448,N_2977,N_2720);
nor U9449 (N_9449,N_2848,N_3762);
and U9450 (N_9450,N_4606,N_4152);
and U9451 (N_9451,N_903,N_4053);
nand U9452 (N_9452,N_2947,N_2838);
and U9453 (N_9453,N_4604,N_2839);
or U9454 (N_9454,N_4149,N_3146);
xnor U9455 (N_9455,N_4259,N_1757);
xor U9456 (N_9456,N_1872,N_1187);
and U9457 (N_9457,N_3340,N_418);
or U9458 (N_9458,N_4237,N_1157);
nor U9459 (N_9459,N_257,N_304);
or U9460 (N_9460,N_2468,N_2158);
xnor U9461 (N_9461,N_2378,N_4629);
nand U9462 (N_9462,N_3461,N_4969);
and U9463 (N_9463,N_4883,N_3224);
and U9464 (N_9464,N_2939,N_2776);
and U9465 (N_9465,N_3823,N_1087);
and U9466 (N_9466,N_2621,N_1842);
and U9467 (N_9467,N_2471,N_708);
nor U9468 (N_9468,N_2817,N_496);
or U9469 (N_9469,N_2698,N_315);
xor U9470 (N_9470,N_266,N_1266);
nor U9471 (N_9471,N_4608,N_4259);
nor U9472 (N_9472,N_4761,N_4588);
and U9473 (N_9473,N_3798,N_4599);
nor U9474 (N_9474,N_2251,N_4207);
or U9475 (N_9475,N_2507,N_2272);
or U9476 (N_9476,N_3781,N_3313);
xor U9477 (N_9477,N_719,N_4490);
nor U9478 (N_9478,N_3938,N_191);
and U9479 (N_9479,N_2735,N_1461);
and U9480 (N_9480,N_2767,N_430);
nor U9481 (N_9481,N_4562,N_22);
and U9482 (N_9482,N_2593,N_2053);
nor U9483 (N_9483,N_3772,N_3996);
nand U9484 (N_9484,N_4620,N_879);
nand U9485 (N_9485,N_4410,N_1529);
and U9486 (N_9486,N_4570,N_2469);
xnor U9487 (N_9487,N_1146,N_407);
nor U9488 (N_9488,N_1213,N_536);
xnor U9489 (N_9489,N_2445,N_3881);
xnor U9490 (N_9490,N_1124,N_2385);
and U9491 (N_9491,N_1929,N_2124);
or U9492 (N_9492,N_1788,N_2405);
or U9493 (N_9493,N_4753,N_480);
xnor U9494 (N_9494,N_1379,N_1039);
nand U9495 (N_9495,N_3894,N_792);
nand U9496 (N_9496,N_1126,N_3544);
and U9497 (N_9497,N_1942,N_2431);
xnor U9498 (N_9498,N_1946,N_3939);
nand U9499 (N_9499,N_647,N_3934);
and U9500 (N_9500,N_211,N_4187);
and U9501 (N_9501,N_64,N_634);
and U9502 (N_9502,N_2191,N_2071);
nor U9503 (N_9503,N_4112,N_3016);
or U9504 (N_9504,N_4430,N_365);
nor U9505 (N_9505,N_712,N_990);
or U9506 (N_9506,N_4575,N_427);
nor U9507 (N_9507,N_2488,N_3640);
xnor U9508 (N_9508,N_4170,N_3178);
and U9509 (N_9509,N_1220,N_1170);
or U9510 (N_9510,N_2730,N_3777);
and U9511 (N_9511,N_1641,N_3783);
and U9512 (N_9512,N_4451,N_267);
nand U9513 (N_9513,N_185,N_2626);
xor U9514 (N_9514,N_848,N_1697);
nor U9515 (N_9515,N_1897,N_3140);
nor U9516 (N_9516,N_2197,N_1069);
and U9517 (N_9517,N_1047,N_859);
or U9518 (N_9518,N_547,N_1125);
nand U9519 (N_9519,N_3702,N_3215);
nor U9520 (N_9520,N_3457,N_572);
or U9521 (N_9521,N_1995,N_1624);
nand U9522 (N_9522,N_4591,N_2512);
and U9523 (N_9523,N_1003,N_4616);
or U9524 (N_9524,N_2944,N_4907);
xor U9525 (N_9525,N_2577,N_3901);
or U9526 (N_9526,N_3092,N_2328);
or U9527 (N_9527,N_741,N_3989);
and U9528 (N_9528,N_1627,N_3750);
and U9529 (N_9529,N_4404,N_101);
nor U9530 (N_9530,N_1606,N_179);
nor U9531 (N_9531,N_3916,N_3619);
and U9532 (N_9532,N_938,N_4953);
and U9533 (N_9533,N_2883,N_184);
or U9534 (N_9534,N_294,N_1213);
nor U9535 (N_9535,N_1902,N_2390);
and U9536 (N_9536,N_4200,N_3840);
nor U9537 (N_9537,N_2881,N_342);
or U9538 (N_9538,N_2111,N_2661);
and U9539 (N_9539,N_1732,N_2674);
xor U9540 (N_9540,N_1079,N_1727);
nand U9541 (N_9541,N_1280,N_1395);
xnor U9542 (N_9542,N_319,N_4449);
xor U9543 (N_9543,N_275,N_4211);
nand U9544 (N_9544,N_1981,N_2115);
nand U9545 (N_9545,N_4284,N_3816);
nand U9546 (N_9546,N_4569,N_3046);
and U9547 (N_9547,N_1577,N_2940);
nor U9548 (N_9548,N_112,N_3986);
or U9549 (N_9549,N_4748,N_4538);
nand U9550 (N_9550,N_3910,N_2919);
and U9551 (N_9551,N_4725,N_3130);
nand U9552 (N_9552,N_4076,N_1766);
nor U9553 (N_9553,N_2730,N_1316);
nand U9554 (N_9554,N_4110,N_225);
nor U9555 (N_9555,N_3607,N_4589);
nor U9556 (N_9556,N_169,N_2541);
nand U9557 (N_9557,N_4200,N_2399);
and U9558 (N_9558,N_1684,N_3119);
or U9559 (N_9559,N_1573,N_4540);
nor U9560 (N_9560,N_2884,N_4650);
or U9561 (N_9561,N_1571,N_3702);
nand U9562 (N_9562,N_1432,N_4973);
xnor U9563 (N_9563,N_3855,N_4265);
nand U9564 (N_9564,N_405,N_2412);
and U9565 (N_9565,N_1807,N_10);
xor U9566 (N_9566,N_917,N_2812);
nor U9567 (N_9567,N_2906,N_31);
nor U9568 (N_9568,N_3065,N_2578);
and U9569 (N_9569,N_515,N_3824);
xor U9570 (N_9570,N_1721,N_3495);
or U9571 (N_9571,N_4688,N_1638);
xor U9572 (N_9572,N_898,N_4776);
nor U9573 (N_9573,N_2131,N_1671);
and U9574 (N_9574,N_371,N_4025);
nor U9575 (N_9575,N_1980,N_1355);
nand U9576 (N_9576,N_1109,N_1972);
xnor U9577 (N_9577,N_1219,N_963);
nand U9578 (N_9578,N_1429,N_1032);
nand U9579 (N_9579,N_149,N_248);
and U9580 (N_9580,N_1638,N_277);
nor U9581 (N_9581,N_794,N_2324);
xor U9582 (N_9582,N_3175,N_1291);
or U9583 (N_9583,N_1174,N_1959);
xnor U9584 (N_9584,N_1410,N_3651);
or U9585 (N_9585,N_554,N_1210);
or U9586 (N_9586,N_4478,N_3670);
nor U9587 (N_9587,N_3080,N_707);
nand U9588 (N_9588,N_901,N_4546);
nand U9589 (N_9589,N_3367,N_2464);
nand U9590 (N_9590,N_2384,N_4656);
nand U9591 (N_9591,N_3408,N_3111);
nor U9592 (N_9592,N_2573,N_1967);
nor U9593 (N_9593,N_1363,N_1898);
nor U9594 (N_9594,N_3899,N_2720);
nor U9595 (N_9595,N_4200,N_3032);
xor U9596 (N_9596,N_303,N_2497);
or U9597 (N_9597,N_2379,N_673);
nand U9598 (N_9598,N_1732,N_4443);
or U9599 (N_9599,N_1816,N_3932);
or U9600 (N_9600,N_4278,N_2005);
or U9601 (N_9601,N_4892,N_2920);
nand U9602 (N_9602,N_395,N_1541);
nor U9603 (N_9603,N_1566,N_1777);
nand U9604 (N_9604,N_518,N_4695);
nor U9605 (N_9605,N_1542,N_1697);
and U9606 (N_9606,N_890,N_1641);
nor U9607 (N_9607,N_2623,N_3537);
and U9608 (N_9608,N_2630,N_4964);
xnor U9609 (N_9609,N_2457,N_865);
nor U9610 (N_9610,N_787,N_664);
nand U9611 (N_9611,N_1629,N_3795);
nor U9612 (N_9612,N_1935,N_1590);
or U9613 (N_9613,N_4986,N_2795);
or U9614 (N_9614,N_3384,N_515);
nand U9615 (N_9615,N_915,N_1295);
nand U9616 (N_9616,N_1405,N_4611);
and U9617 (N_9617,N_4403,N_1286);
nand U9618 (N_9618,N_1616,N_1844);
xnor U9619 (N_9619,N_1765,N_3515);
xnor U9620 (N_9620,N_3596,N_3232);
nor U9621 (N_9621,N_2892,N_11);
or U9622 (N_9622,N_1551,N_3581);
and U9623 (N_9623,N_1533,N_4615);
and U9624 (N_9624,N_315,N_4952);
xnor U9625 (N_9625,N_4215,N_4048);
or U9626 (N_9626,N_1330,N_854);
xor U9627 (N_9627,N_839,N_852);
xor U9628 (N_9628,N_2234,N_1632);
and U9629 (N_9629,N_4647,N_1805);
xnor U9630 (N_9630,N_2576,N_2722);
nor U9631 (N_9631,N_4778,N_405);
nand U9632 (N_9632,N_446,N_1632);
nor U9633 (N_9633,N_294,N_4770);
and U9634 (N_9634,N_518,N_2133);
or U9635 (N_9635,N_2809,N_456);
and U9636 (N_9636,N_4728,N_4810);
nor U9637 (N_9637,N_1948,N_3930);
nand U9638 (N_9638,N_3907,N_1290);
and U9639 (N_9639,N_2960,N_4986);
or U9640 (N_9640,N_4720,N_1544);
nand U9641 (N_9641,N_2111,N_1814);
xor U9642 (N_9642,N_1258,N_1280);
nand U9643 (N_9643,N_962,N_1841);
nor U9644 (N_9644,N_3525,N_1838);
nand U9645 (N_9645,N_4905,N_3869);
xnor U9646 (N_9646,N_2109,N_3450);
xnor U9647 (N_9647,N_4551,N_4544);
xor U9648 (N_9648,N_2456,N_28);
or U9649 (N_9649,N_274,N_3516);
nand U9650 (N_9650,N_3597,N_4390);
nand U9651 (N_9651,N_3314,N_4159);
xnor U9652 (N_9652,N_4469,N_3967);
or U9653 (N_9653,N_1125,N_4120);
and U9654 (N_9654,N_2013,N_3533);
or U9655 (N_9655,N_1108,N_1768);
and U9656 (N_9656,N_395,N_507);
nand U9657 (N_9657,N_2546,N_1226);
or U9658 (N_9658,N_398,N_3120);
nor U9659 (N_9659,N_3028,N_1547);
nor U9660 (N_9660,N_4854,N_396);
or U9661 (N_9661,N_2186,N_4237);
and U9662 (N_9662,N_4574,N_1901);
xor U9663 (N_9663,N_1860,N_4892);
nor U9664 (N_9664,N_191,N_517);
xor U9665 (N_9665,N_1190,N_1279);
or U9666 (N_9666,N_3924,N_1012);
nor U9667 (N_9667,N_3603,N_260);
xor U9668 (N_9668,N_1782,N_1816);
nand U9669 (N_9669,N_656,N_3941);
nor U9670 (N_9670,N_2503,N_4652);
nor U9671 (N_9671,N_619,N_2819);
xnor U9672 (N_9672,N_781,N_1896);
or U9673 (N_9673,N_3872,N_3153);
nor U9674 (N_9674,N_3978,N_189);
and U9675 (N_9675,N_2784,N_2735);
nor U9676 (N_9676,N_4483,N_2464);
or U9677 (N_9677,N_4652,N_4157);
or U9678 (N_9678,N_900,N_2286);
nand U9679 (N_9679,N_3684,N_1679);
or U9680 (N_9680,N_2069,N_3282);
xnor U9681 (N_9681,N_1686,N_3203);
nand U9682 (N_9682,N_4805,N_4999);
and U9683 (N_9683,N_2505,N_524);
or U9684 (N_9684,N_2719,N_2286);
and U9685 (N_9685,N_2476,N_2328);
xnor U9686 (N_9686,N_1556,N_162);
or U9687 (N_9687,N_3583,N_4564);
and U9688 (N_9688,N_1791,N_4467);
and U9689 (N_9689,N_306,N_2605);
nand U9690 (N_9690,N_4362,N_600);
nand U9691 (N_9691,N_3305,N_161);
and U9692 (N_9692,N_1337,N_5);
or U9693 (N_9693,N_3012,N_2227);
nand U9694 (N_9694,N_4691,N_1602);
or U9695 (N_9695,N_2364,N_138);
xor U9696 (N_9696,N_2188,N_3044);
nor U9697 (N_9697,N_1397,N_3605);
and U9698 (N_9698,N_3698,N_1580);
and U9699 (N_9699,N_2754,N_3967);
or U9700 (N_9700,N_833,N_610);
nand U9701 (N_9701,N_585,N_4519);
and U9702 (N_9702,N_312,N_4774);
xnor U9703 (N_9703,N_2461,N_670);
xor U9704 (N_9704,N_2525,N_3409);
nor U9705 (N_9705,N_2461,N_2381);
nor U9706 (N_9706,N_3412,N_510);
and U9707 (N_9707,N_1583,N_77);
nor U9708 (N_9708,N_2637,N_4459);
xnor U9709 (N_9709,N_2096,N_4324);
nand U9710 (N_9710,N_2320,N_3016);
nand U9711 (N_9711,N_444,N_2426);
and U9712 (N_9712,N_4219,N_820);
nor U9713 (N_9713,N_1936,N_347);
or U9714 (N_9714,N_3566,N_3288);
nor U9715 (N_9715,N_2277,N_1818);
nand U9716 (N_9716,N_1272,N_2402);
and U9717 (N_9717,N_1083,N_3163);
and U9718 (N_9718,N_4009,N_1378);
nand U9719 (N_9719,N_4015,N_2489);
or U9720 (N_9720,N_2310,N_3275);
xnor U9721 (N_9721,N_2324,N_3325);
and U9722 (N_9722,N_2104,N_1780);
nand U9723 (N_9723,N_859,N_2509);
or U9724 (N_9724,N_4784,N_1509);
nand U9725 (N_9725,N_4662,N_3293);
or U9726 (N_9726,N_1455,N_4201);
or U9727 (N_9727,N_2259,N_3428);
nand U9728 (N_9728,N_1280,N_3773);
xnor U9729 (N_9729,N_980,N_1557);
or U9730 (N_9730,N_2688,N_3937);
nand U9731 (N_9731,N_3545,N_3828);
or U9732 (N_9732,N_4093,N_269);
and U9733 (N_9733,N_4499,N_597);
or U9734 (N_9734,N_896,N_2541);
xor U9735 (N_9735,N_4872,N_3364);
and U9736 (N_9736,N_4616,N_2544);
xnor U9737 (N_9737,N_3534,N_739);
and U9738 (N_9738,N_4608,N_4257);
nor U9739 (N_9739,N_4248,N_1671);
or U9740 (N_9740,N_4071,N_1483);
nor U9741 (N_9741,N_738,N_694);
nor U9742 (N_9742,N_2793,N_1585);
or U9743 (N_9743,N_2062,N_1440);
nand U9744 (N_9744,N_974,N_2194);
nor U9745 (N_9745,N_3164,N_1330);
or U9746 (N_9746,N_2022,N_1713);
and U9747 (N_9747,N_4963,N_1013);
nor U9748 (N_9748,N_428,N_4972);
nor U9749 (N_9749,N_779,N_2928);
xnor U9750 (N_9750,N_4815,N_1421);
xnor U9751 (N_9751,N_2226,N_4309);
nor U9752 (N_9752,N_4060,N_290);
or U9753 (N_9753,N_1657,N_4388);
xor U9754 (N_9754,N_783,N_1897);
nand U9755 (N_9755,N_2436,N_3278);
or U9756 (N_9756,N_3288,N_3737);
nor U9757 (N_9757,N_2528,N_316);
or U9758 (N_9758,N_2623,N_3227);
and U9759 (N_9759,N_1803,N_179);
and U9760 (N_9760,N_2673,N_1626);
nor U9761 (N_9761,N_1999,N_2042);
nand U9762 (N_9762,N_979,N_632);
or U9763 (N_9763,N_1455,N_1259);
nand U9764 (N_9764,N_3950,N_1755);
or U9765 (N_9765,N_1010,N_3021);
and U9766 (N_9766,N_3815,N_36);
xnor U9767 (N_9767,N_1986,N_4849);
nand U9768 (N_9768,N_2087,N_4623);
nor U9769 (N_9769,N_3788,N_4143);
and U9770 (N_9770,N_3756,N_1491);
or U9771 (N_9771,N_4102,N_1189);
nor U9772 (N_9772,N_3145,N_3304);
and U9773 (N_9773,N_2098,N_620);
nand U9774 (N_9774,N_1772,N_1735);
or U9775 (N_9775,N_857,N_2631);
or U9776 (N_9776,N_3230,N_2970);
nor U9777 (N_9777,N_569,N_3101);
xnor U9778 (N_9778,N_4435,N_4764);
and U9779 (N_9779,N_1762,N_2224);
or U9780 (N_9780,N_4146,N_1560);
and U9781 (N_9781,N_3397,N_2376);
nand U9782 (N_9782,N_3593,N_1537);
and U9783 (N_9783,N_3954,N_1367);
nand U9784 (N_9784,N_2932,N_2377);
nor U9785 (N_9785,N_2877,N_2987);
nor U9786 (N_9786,N_3811,N_4859);
nor U9787 (N_9787,N_4148,N_3823);
or U9788 (N_9788,N_2414,N_3951);
and U9789 (N_9789,N_994,N_384);
nand U9790 (N_9790,N_3430,N_2038);
nand U9791 (N_9791,N_4181,N_2458);
and U9792 (N_9792,N_4583,N_2288);
or U9793 (N_9793,N_1439,N_1484);
and U9794 (N_9794,N_1869,N_702);
xor U9795 (N_9795,N_899,N_4819);
nand U9796 (N_9796,N_536,N_698);
xnor U9797 (N_9797,N_3563,N_3937);
nor U9798 (N_9798,N_2066,N_2019);
nand U9799 (N_9799,N_4522,N_2195);
xor U9800 (N_9800,N_4640,N_3923);
nand U9801 (N_9801,N_2704,N_3958);
nor U9802 (N_9802,N_2921,N_1365);
nor U9803 (N_9803,N_4299,N_1538);
and U9804 (N_9804,N_3672,N_1883);
or U9805 (N_9805,N_281,N_1518);
or U9806 (N_9806,N_1723,N_3440);
nand U9807 (N_9807,N_1996,N_1308);
or U9808 (N_9808,N_1507,N_686);
nand U9809 (N_9809,N_2102,N_4853);
and U9810 (N_9810,N_4201,N_919);
xor U9811 (N_9811,N_492,N_1945);
and U9812 (N_9812,N_3824,N_492);
xor U9813 (N_9813,N_3247,N_1920);
or U9814 (N_9814,N_322,N_2471);
and U9815 (N_9815,N_2743,N_3887);
or U9816 (N_9816,N_2120,N_4348);
and U9817 (N_9817,N_1762,N_2268);
or U9818 (N_9818,N_403,N_1992);
nor U9819 (N_9819,N_2847,N_3686);
and U9820 (N_9820,N_2086,N_3659);
or U9821 (N_9821,N_1937,N_304);
or U9822 (N_9822,N_2119,N_886);
nand U9823 (N_9823,N_2485,N_1558);
nor U9824 (N_9824,N_662,N_2421);
nor U9825 (N_9825,N_246,N_995);
nand U9826 (N_9826,N_3580,N_2123);
or U9827 (N_9827,N_4363,N_3799);
xnor U9828 (N_9828,N_4500,N_3477);
or U9829 (N_9829,N_1704,N_1490);
nor U9830 (N_9830,N_4345,N_4647);
or U9831 (N_9831,N_1894,N_1858);
nand U9832 (N_9832,N_1447,N_2427);
nand U9833 (N_9833,N_3997,N_1723);
nor U9834 (N_9834,N_4776,N_4313);
or U9835 (N_9835,N_2455,N_1224);
xor U9836 (N_9836,N_4550,N_286);
nand U9837 (N_9837,N_1321,N_2391);
nor U9838 (N_9838,N_4869,N_975);
and U9839 (N_9839,N_2228,N_1030);
xnor U9840 (N_9840,N_4504,N_3719);
xor U9841 (N_9841,N_69,N_2513);
or U9842 (N_9842,N_4236,N_1003);
or U9843 (N_9843,N_2853,N_971);
xor U9844 (N_9844,N_3060,N_2442);
xor U9845 (N_9845,N_4690,N_2183);
nand U9846 (N_9846,N_3473,N_627);
xor U9847 (N_9847,N_4519,N_1422);
and U9848 (N_9848,N_994,N_4368);
and U9849 (N_9849,N_997,N_3131);
nor U9850 (N_9850,N_3350,N_4651);
xnor U9851 (N_9851,N_3276,N_966);
or U9852 (N_9852,N_254,N_443);
xor U9853 (N_9853,N_3100,N_362);
nor U9854 (N_9854,N_2837,N_1501);
or U9855 (N_9855,N_2645,N_4153);
nor U9856 (N_9856,N_3379,N_3567);
or U9857 (N_9857,N_866,N_2785);
xor U9858 (N_9858,N_3201,N_654);
nor U9859 (N_9859,N_3769,N_2915);
nor U9860 (N_9860,N_2710,N_2951);
xnor U9861 (N_9861,N_1067,N_3888);
xor U9862 (N_9862,N_4045,N_3228);
nor U9863 (N_9863,N_4486,N_3064);
xor U9864 (N_9864,N_740,N_4305);
and U9865 (N_9865,N_1826,N_531);
nand U9866 (N_9866,N_837,N_4254);
xor U9867 (N_9867,N_2050,N_218);
nor U9868 (N_9868,N_658,N_2379);
nand U9869 (N_9869,N_1888,N_953);
nand U9870 (N_9870,N_3999,N_2756);
and U9871 (N_9871,N_4334,N_3011);
and U9872 (N_9872,N_4780,N_4989);
nand U9873 (N_9873,N_3159,N_3797);
and U9874 (N_9874,N_3998,N_2938);
or U9875 (N_9875,N_3461,N_3784);
or U9876 (N_9876,N_4851,N_1183);
nor U9877 (N_9877,N_1003,N_1027);
or U9878 (N_9878,N_1706,N_2050);
and U9879 (N_9879,N_3087,N_3766);
and U9880 (N_9880,N_2807,N_3057);
or U9881 (N_9881,N_3823,N_666);
nor U9882 (N_9882,N_4463,N_3686);
and U9883 (N_9883,N_3255,N_3028);
xnor U9884 (N_9884,N_2926,N_4473);
or U9885 (N_9885,N_1922,N_918);
nand U9886 (N_9886,N_4349,N_1765);
and U9887 (N_9887,N_4388,N_500);
nand U9888 (N_9888,N_3461,N_3646);
nand U9889 (N_9889,N_2050,N_112);
xnor U9890 (N_9890,N_1205,N_941);
or U9891 (N_9891,N_3620,N_2040);
nor U9892 (N_9892,N_1966,N_903);
xnor U9893 (N_9893,N_561,N_1141);
nor U9894 (N_9894,N_2768,N_1597);
and U9895 (N_9895,N_335,N_2960);
nand U9896 (N_9896,N_2953,N_939);
nand U9897 (N_9897,N_809,N_3415);
or U9898 (N_9898,N_1846,N_3152);
nor U9899 (N_9899,N_975,N_1654);
xor U9900 (N_9900,N_2170,N_2702);
and U9901 (N_9901,N_889,N_3998);
xnor U9902 (N_9902,N_531,N_3294);
nand U9903 (N_9903,N_4203,N_1138);
nand U9904 (N_9904,N_2209,N_3800);
and U9905 (N_9905,N_3116,N_2786);
nand U9906 (N_9906,N_1057,N_3070);
or U9907 (N_9907,N_2017,N_697);
nand U9908 (N_9908,N_4313,N_3931);
nand U9909 (N_9909,N_3513,N_4630);
nand U9910 (N_9910,N_4258,N_496);
and U9911 (N_9911,N_899,N_3023);
or U9912 (N_9912,N_1633,N_1239);
xor U9913 (N_9913,N_1190,N_3973);
and U9914 (N_9914,N_981,N_3549);
and U9915 (N_9915,N_541,N_4324);
nand U9916 (N_9916,N_4839,N_0);
or U9917 (N_9917,N_781,N_3642);
and U9918 (N_9918,N_340,N_2884);
xnor U9919 (N_9919,N_463,N_3390);
xor U9920 (N_9920,N_2385,N_3197);
nand U9921 (N_9921,N_2512,N_3695);
xnor U9922 (N_9922,N_2698,N_3145);
or U9923 (N_9923,N_3212,N_4331);
or U9924 (N_9924,N_669,N_3708);
and U9925 (N_9925,N_4791,N_1674);
nor U9926 (N_9926,N_3302,N_4978);
and U9927 (N_9927,N_2253,N_874);
and U9928 (N_9928,N_3667,N_2687);
or U9929 (N_9929,N_3044,N_4488);
or U9930 (N_9930,N_4062,N_798);
nor U9931 (N_9931,N_2642,N_2244);
nor U9932 (N_9932,N_3557,N_2325);
and U9933 (N_9933,N_262,N_3137);
and U9934 (N_9934,N_1717,N_3173);
xnor U9935 (N_9935,N_2400,N_731);
nand U9936 (N_9936,N_1540,N_2136);
xor U9937 (N_9937,N_3221,N_3783);
and U9938 (N_9938,N_4784,N_1521);
nand U9939 (N_9939,N_3817,N_2940);
nor U9940 (N_9940,N_3595,N_1430);
nand U9941 (N_9941,N_4813,N_844);
or U9942 (N_9942,N_2280,N_1114);
nor U9943 (N_9943,N_2930,N_4707);
nand U9944 (N_9944,N_258,N_2060);
nand U9945 (N_9945,N_1643,N_2381);
or U9946 (N_9946,N_2918,N_2140);
nand U9947 (N_9947,N_2894,N_4137);
nand U9948 (N_9948,N_2792,N_165);
xor U9949 (N_9949,N_401,N_4618);
or U9950 (N_9950,N_3781,N_2492);
and U9951 (N_9951,N_213,N_3857);
nand U9952 (N_9952,N_3365,N_2747);
and U9953 (N_9953,N_4181,N_4630);
nand U9954 (N_9954,N_859,N_3724);
nand U9955 (N_9955,N_1346,N_228);
nand U9956 (N_9956,N_4275,N_82);
nand U9957 (N_9957,N_1912,N_831);
nor U9958 (N_9958,N_3825,N_4753);
and U9959 (N_9959,N_3828,N_1068);
and U9960 (N_9960,N_460,N_2302);
or U9961 (N_9961,N_2594,N_203);
and U9962 (N_9962,N_3204,N_4847);
or U9963 (N_9963,N_1603,N_1831);
nand U9964 (N_9964,N_733,N_2324);
and U9965 (N_9965,N_763,N_522);
xnor U9966 (N_9966,N_3591,N_4175);
nor U9967 (N_9967,N_11,N_4127);
and U9968 (N_9968,N_2059,N_2383);
or U9969 (N_9969,N_2244,N_2431);
and U9970 (N_9970,N_260,N_2464);
xor U9971 (N_9971,N_4803,N_4892);
nand U9972 (N_9972,N_3876,N_1113);
nor U9973 (N_9973,N_857,N_81);
xor U9974 (N_9974,N_3548,N_2341);
xor U9975 (N_9975,N_753,N_2666);
nor U9976 (N_9976,N_318,N_2471);
or U9977 (N_9977,N_2494,N_1561);
nor U9978 (N_9978,N_4613,N_1780);
nor U9979 (N_9979,N_3276,N_3995);
or U9980 (N_9980,N_1506,N_2807);
and U9981 (N_9981,N_4700,N_1466);
or U9982 (N_9982,N_4753,N_1284);
nand U9983 (N_9983,N_553,N_2052);
nor U9984 (N_9984,N_4754,N_3101);
or U9985 (N_9985,N_1910,N_1749);
nand U9986 (N_9986,N_981,N_3020);
and U9987 (N_9987,N_980,N_4952);
and U9988 (N_9988,N_726,N_2480);
nor U9989 (N_9989,N_2491,N_284);
nand U9990 (N_9990,N_1362,N_1291);
nor U9991 (N_9991,N_4326,N_4250);
nand U9992 (N_9992,N_2052,N_3535);
nand U9993 (N_9993,N_3546,N_1725);
or U9994 (N_9994,N_1940,N_1531);
and U9995 (N_9995,N_4383,N_1760);
and U9996 (N_9996,N_2418,N_2716);
nor U9997 (N_9997,N_306,N_4228);
xnor U9998 (N_9998,N_2864,N_3685);
xnor U9999 (N_9999,N_4563,N_3785);
or U10000 (N_10000,N_9533,N_9690);
xor U10001 (N_10001,N_6815,N_7789);
and U10002 (N_10002,N_8514,N_6883);
and U10003 (N_10003,N_6438,N_8019);
nand U10004 (N_10004,N_5220,N_8814);
nand U10005 (N_10005,N_6732,N_7055);
nor U10006 (N_10006,N_9752,N_8887);
and U10007 (N_10007,N_6402,N_5058);
xor U10008 (N_10008,N_5834,N_9857);
nand U10009 (N_10009,N_6631,N_8707);
nand U10010 (N_10010,N_9045,N_8842);
xor U10011 (N_10011,N_6670,N_6326);
and U10012 (N_10012,N_7728,N_8780);
xor U10013 (N_10013,N_5630,N_7568);
xor U10014 (N_10014,N_5318,N_9260);
and U10015 (N_10015,N_5144,N_5176);
nand U10016 (N_10016,N_9021,N_7649);
xnor U10017 (N_10017,N_8025,N_7888);
nor U10018 (N_10018,N_9273,N_8954);
nor U10019 (N_10019,N_6575,N_7735);
xor U10020 (N_10020,N_8477,N_7667);
xnor U10021 (N_10021,N_8429,N_7493);
or U10022 (N_10022,N_5773,N_9854);
xnor U10023 (N_10023,N_6268,N_6070);
nor U10024 (N_10024,N_9839,N_5407);
nor U10025 (N_10025,N_7379,N_8447);
or U10026 (N_10026,N_5118,N_6618);
nor U10027 (N_10027,N_7634,N_7793);
xor U10028 (N_10028,N_9562,N_5725);
nand U10029 (N_10029,N_8028,N_9284);
or U10030 (N_10030,N_8096,N_9984);
nor U10031 (N_10031,N_6408,N_7841);
nor U10032 (N_10032,N_6876,N_6581);
nor U10033 (N_10033,N_6279,N_7441);
nor U10034 (N_10034,N_7121,N_7617);
nor U10035 (N_10035,N_5526,N_5676);
nand U10036 (N_10036,N_9244,N_8748);
nor U10037 (N_10037,N_7037,N_7541);
xor U10038 (N_10038,N_7264,N_5071);
nor U10039 (N_10039,N_7343,N_9873);
or U10040 (N_10040,N_7699,N_5518);
nor U10041 (N_10041,N_9238,N_6629);
nor U10042 (N_10042,N_9830,N_8679);
and U10043 (N_10043,N_7756,N_8844);
or U10044 (N_10044,N_6170,N_6640);
nor U10045 (N_10045,N_6867,N_8967);
and U10046 (N_10046,N_8457,N_8758);
nand U10047 (N_10047,N_7399,N_7713);
nand U10048 (N_10048,N_8008,N_5499);
nor U10049 (N_10049,N_6582,N_8724);
or U10050 (N_10050,N_9859,N_8589);
or U10051 (N_10051,N_8878,N_5788);
nor U10052 (N_10052,N_7350,N_5736);
and U10053 (N_10053,N_6156,N_8284);
nor U10054 (N_10054,N_5020,N_9052);
xor U10055 (N_10055,N_5158,N_7676);
or U10056 (N_10056,N_7389,N_8868);
and U10057 (N_10057,N_8393,N_9787);
or U10058 (N_10058,N_9982,N_8975);
or U10059 (N_10059,N_8643,N_8932);
xnor U10060 (N_10060,N_7895,N_5771);
or U10061 (N_10061,N_8599,N_6101);
or U10062 (N_10062,N_6941,N_6298);
and U10063 (N_10063,N_9082,N_9347);
or U10064 (N_10064,N_5816,N_5899);
xnor U10065 (N_10065,N_5049,N_6263);
xor U10066 (N_10066,N_8093,N_7693);
nor U10067 (N_10067,N_6793,N_8017);
or U10068 (N_10068,N_8247,N_5939);
and U10069 (N_10069,N_6313,N_6009);
xor U10070 (N_10070,N_7831,N_5243);
nor U10071 (N_10071,N_8164,N_7301);
xnor U10072 (N_10072,N_9832,N_7336);
nand U10073 (N_10073,N_6538,N_5821);
xor U10074 (N_10074,N_7886,N_5219);
and U10075 (N_10075,N_6634,N_9644);
and U10076 (N_10076,N_9774,N_7276);
or U10077 (N_10077,N_9550,N_5187);
or U10078 (N_10078,N_6537,N_5491);
xnor U10079 (N_10079,N_9462,N_5803);
xnor U10080 (N_10080,N_6801,N_7365);
nand U10081 (N_10081,N_7603,N_9889);
and U10082 (N_10082,N_8836,N_7280);
and U10083 (N_10083,N_6451,N_7746);
or U10084 (N_10084,N_6820,N_9215);
and U10085 (N_10085,N_8580,N_7885);
nand U10086 (N_10086,N_7712,N_8060);
nor U10087 (N_10087,N_8896,N_7443);
and U10088 (N_10088,N_9812,N_8181);
and U10089 (N_10089,N_9996,N_8144);
or U10090 (N_10090,N_7013,N_7259);
nand U10091 (N_10091,N_5321,N_8658);
and U10092 (N_10092,N_6990,N_6118);
xor U10093 (N_10093,N_8491,N_9331);
and U10094 (N_10094,N_9039,N_8249);
and U10095 (N_10095,N_9521,N_8980);
xor U10096 (N_10096,N_8466,N_8108);
nand U10097 (N_10097,N_5201,N_6217);
xnor U10098 (N_10098,N_6223,N_8979);
xor U10099 (N_10099,N_8610,N_5983);
nor U10100 (N_10100,N_7230,N_9910);
or U10101 (N_10101,N_6973,N_6863);
or U10102 (N_10102,N_6977,N_5864);
or U10103 (N_10103,N_6129,N_9792);
nor U10104 (N_10104,N_7088,N_8867);
and U10105 (N_10105,N_9921,N_5808);
or U10106 (N_10106,N_8297,N_6744);
and U10107 (N_10107,N_8823,N_9038);
nand U10108 (N_10108,N_6940,N_9168);
and U10109 (N_10109,N_6355,N_9934);
xnor U10110 (N_10110,N_5610,N_5712);
or U10111 (N_10111,N_8890,N_7976);
nor U10112 (N_10112,N_9738,N_5211);
nor U10113 (N_10113,N_8485,N_7854);
xnor U10114 (N_10114,N_8224,N_7318);
xor U10115 (N_10115,N_6910,N_9141);
or U10116 (N_10116,N_9416,N_9256);
or U10117 (N_10117,N_8331,N_9085);
and U10118 (N_10118,N_7560,N_5358);
xnor U10119 (N_10119,N_9335,N_7265);
and U10120 (N_10120,N_8227,N_7559);
or U10121 (N_10121,N_5578,N_7434);
or U10122 (N_10122,N_8791,N_8808);
or U10123 (N_10123,N_8433,N_5165);
and U10124 (N_10124,N_9708,N_9618);
nor U10125 (N_10125,N_5238,N_5730);
nand U10126 (N_10126,N_9295,N_5598);
nand U10127 (N_10127,N_6092,N_9578);
nor U10128 (N_10128,N_8322,N_9504);
and U10129 (N_10129,N_6344,N_7966);
or U10130 (N_10130,N_8766,N_7381);
nand U10131 (N_10131,N_9376,N_5533);
nor U10132 (N_10132,N_5625,N_7144);
and U10133 (N_10133,N_6844,N_7754);
nor U10134 (N_10134,N_9123,N_7557);
xnor U10135 (N_10135,N_7120,N_7372);
xnor U10136 (N_10136,N_5404,N_7353);
nor U10137 (N_10137,N_5822,N_8973);
nand U10138 (N_10138,N_6405,N_9140);
nand U10139 (N_10139,N_7812,N_5599);
or U10140 (N_10140,N_6703,N_7476);
xnor U10141 (N_10141,N_6446,N_7583);
nor U10142 (N_10142,N_5953,N_8609);
or U10143 (N_10143,N_5589,N_6672);
nand U10144 (N_10144,N_5095,N_6248);
nor U10145 (N_10145,N_7995,N_6544);
or U10146 (N_10146,N_5979,N_7190);
or U10147 (N_10147,N_9214,N_8186);
nor U10148 (N_10148,N_9239,N_9429);
nand U10149 (N_10149,N_5690,N_5539);
xor U10150 (N_10150,N_6783,N_8551);
nand U10151 (N_10151,N_5796,N_5760);
and U10152 (N_10152,N_5591,N_5437);
nand U10153 (N_10153,N_8966,N_8061);
or U10154 (N_10154,N_6122,N_9961);
and U10155 (N_10155,N_7149,N_6680);
or U10156 (N_10156,N_9636,N_5500);
or U10157 (N_10157,N_8441,N_6262);
nand U10158 (N_10158,N_7123,N_5570);
or U10159 (N_10159,N_6816,N_6964);
nor U10160 (N_10160,N_9553,N_9303);
and U10161 (N_10161,N_5141,N_9699);
xnor U10162 (N_10162,N_7141,N_6418);
nor U10163 (N_10163,N_7707,N_5868);
nor U10164 (N_10164,N_7802,N_7354);
and U10165 (N_10165,N_8696,N_8112);
or U10166 (N_10166,N_6585,N_5643);
xor U10167 (N_10167,N_9795,N_6578);
nor U10168 (N_10168,N_7852,N_7824);
xnor U10169 (N_10169,N_6315,N_6623);
nand U10170 (N_10170,N_9131,N_9970);
and U10171 (N_10171,N_7239,N_8291);
or U10172 (N_10172,N_6372,N_7578);
and U10173 (N_10173,N_7352,N_9374);
or U10174 (N_10174,N_7509,N_6958);
nor U10175 (N_10175,N_7504,N_5913);
and U10176 (N_10176,N_8330,N_9081);
nand U10177 (N_10177,N_8194,N_5915);
nor U10178 (N_10178,N_8241,N_5584);
and U10179 (N_10179,N_9664,N_5726);
nor U10180 (N_10180,N_8238,N_9298);
or U10181 (N_10181,N_5932,N_7075);
xor U10182 (N_10182,N_6561,N_5546);
or U10183 (N_10183,N_7142,N_5278);
nor U10184 (N_10184,N_7759,N_6887);
and U10185 (N_10185,N_9978,N_8803);
and U10186 (N_10186,N_5798,N_7705);
xor U10187 (N_10187,N_8257,N_6157);
xor U10188 (N_10188,N_9304,N_6955);
xnor U10189 (N_10189,N_7018,N_5448);
or U10190 (N_10190,N_8732,N_5799);
or U10191 (N_10191,N_5964,N_5000);
nor U10192 (N_10192,N_7737,N_6567);
and U10193 (N_10193,N_8911,N_8290);
nand U10194 (N_10194,N_7813,N_5950);
nor U10195 (N_10195,N_7192,N_9451);
or U10196 (N_10196,N_6753,N_6603);
nand U10197 (N_10197,N_9422,N_7956);
xnor U10198 (N_10198,N_6385,N_7105);
xnor U10199 (N_10199,N_5093,N_5752);
xor U10200 (N_10200,N_8346,N_5860);
and U10201 (N_10201,N_5743,N_7471);
and U10202 (N_10202,N_8901,N_7223);
nor U10203 (N_10203,N_8571,N_9975);
or U10204 (N_10204,N_6764,N_8719);
nor U10205 (N_10205,N_6025,N_9761);
nand U10206 (N_10206,N_5172,N_6758);
nand U10207 (N_10207,N_8588,N_8212);
and U10208 (N_10208,N_6879,N_9296);
or U10209 (N_10209,N_7401,N_6574);
nor U10210 (N_10210,N_5421,N_9108);
or U10211 (N_10211,N_8948,N_6008);
nand U10212 (N_10212,N_5096,N_8461);
or U10213 (N_10213,N_8745,N_9243);
nand U10214 (N_10214,N_5360,N_7270);
nor U10215 (N_10215,N_8215,N_8971);
nand U10216 (N_10216,N_8851,N_9166);
nand U10217 (N_10217,N_6282,N_5253);
nor U10218 (N_10218,N_7134,N_9345);
or U10219 (N_10219,N_5431,N_7781);
nand U10220 (N_10220,N_7536,N_7216);
or U10221 (N_10221,N_8459,N_6570);
xnor U10222 (N_10222,N_6205,N_5588);
xnor U10223 (N_10223,N_5716,N_8360);
and U10224 (N_10224,N_7009,N_6023);
nor U10225 (N_10225,N_9440,N_9765);
nand U10226 (N_10226,N_5128,N_9363);
xor U10227 (N_10227,N_7889,N_9925);
nand U10228 (N_10228,N_5449,N_7650);
nand U10229 (N_10229,N_8970,N_5345);
or U10230 (N_10230,N_6461,N_5368);
nor U10231 (N_10231,N_7774,N_9145);
nand U10232 (N_10232,N_7939,N_7750);
nand U10233 (N_10233,N_6305,N_6192);
xor U10234 (N_10234,N_8933,N_6102);
nand U10235 (N_10235,N_9734,N_9588);
and U10236 (N_10236,N_6474,N_8796);
or U10237 (N_10237,N_8993,N_9788);
nor U10238 (N_10238,N_8286,N_8147);
nor U10239 (N_10239,N_8757,N_5889);
or U10240 (N_10240,N_6889,N_6925);
xor U10241 (N_10241,N_9223,N_7309);
and U10242 (N_10242,N_9778,N_8114);
or U10243 (N_10243,N_9005,N_5981);
and U10244 (N_10244,N_5818,N_7256);
xor U10245 (N_10245,N_8462,N_8509);
or U10246 (N_10246,N_9030,N_6151);
nor U10247 (N_10247,N_6416,N_7883);
nor U10248 (N_10248,N_9790,N_5522);
nand U10249 (N_10249,N_7522,N_9515);
nor U10250 (N_10250,N_6447,N_6004);
nand U10251 (N_10251,N_5907,N_5848);
or U10252 (N_10252,N_9603,N_7106);
nor U10253 (N_10253,N_8914,N_8098);
xnor U10254 (N_10254,N_8770,N_6518);
xor U10255 (N_10255,N_5579,N_7954);
nand U10256 (N_10256,N_6286,N_9130);
nor U10257 (N_10257,N_9027,N_5363);
nor U10258 (N_10258,N_6614,N_6909);
nor U10259 (N_10259,N_5855,N_9084);
or U10260 (N_10260,N_9763,N_7537);
and U10261 (N_10261,N_6633,N_6987);
or U10262 (N_10262,N_8103,N_6699);
and U10263 (N_10263,N_9330,N_7618);
xnor U10264 (N_10264,N_7472,N_7539);
nand U10265 (N_10265,N_9139,N_9217);
xnor U10266 (N_10266,N_8591,N_5662);
or U10267 (N_10267,N_7874,N_9877);
nand U10268 (N_10268,N_6558,N_9770);
nor U10269 (N_10269,N_9104,N_6245);
and U10270 (N_10270,N_6865,N_8774);
or U10271 (N_10271,N_7506,N_6836);
nor U10272 (N_10272,N_8526,N_8334);
xnor U10273 (N_10273,N_7971,N_5688);
or U10274 (N_10274,N_8006,N_7589);
or U10275 (N_10275,N_5426,N_7411);
xor U10276 (N_10276,N_6254,N_8986);
xnor U10277 (N_10277,N_6420,N_7101);
nor U10278 (N_10278,N_5530,N_9360);
and U10279 (N_10279,N_9871,N_7292);
and U10280 (N_10280,N_9173,N_9319);
xor U10281 (N_10281,N_6334,N_7868);
and U10282 (N_10282,N_8064,N_9418);
nand U10283 (N_10283,N_9261,N_7273);
nor U10284 (N_10284,N_5543,N_8573);
nor U10285 (N_10285,N_6267,N_9133);
nand U10286 (N_10286,N_6682,N_5346);
xor U10287 (N_10287,N_9758,N_8964);
xnor U10288 (N_10288,N_9268,N_8128);
nor U10289 (N_10289,N_8501,N_6924);
xor U10290 (N_10290,N_5621,N_5463);
nor U10291 (N_10291,N_5721,N_6845);
or U10292 (N_10292,N_9643,N_9764);
and U10293 (N_10293,N_6596,N_6087);
or U10294 (N_10294,N_9674,N_5664);
nand U10295 (N_10295,N_6123,N_7428);
or U10296 (N_10296,N_8208,N_6110);
xor U10297 (N_10297,N_7905,N_6178);
and U10298 (N_10298,N_8261,N_7054);
and U10299 (N_10299,N_9829,N_9035);
nor U10300 (N_10300,N_6899,N_7688);
and U10301 (N_10301,N_6489,N_7201);
nor U10302 (N_10302,N_8176,N_7990);
xor U10303 (N_10303,N_7810,N_6880);
xnor U10304 (N_10304,N_7394,N_5971);
nand U10305 (N_10305,N_9118,N_9164);
or U10306 (N_10306,N_7546,N_5099);
nand U10307 (N_10307,N_9019,N_6382);
nor U10308 (N_10308,N_5405,N_5677);
or U10309 (N_10309,N_6505,N_8513);
nand U10310 (N_10310,N_7588,N_5215);
xor U10311 (N_10311,N_6183,N_8192);
or U10312 (N_10312,N_6919,N_7770);
nand U10313 (N_10313,N_9836,N_6549);
nand U10314 (N_10314,N_8529,N_5954);
or U10315 (N_10315,N_9658,N_8549);
and U10316 (N_10316,N_5438,N_5890);
or U10317 (N_10317,N_5135,N_9291);
or U10318 (N_10318,N_9097,N_6806);
or U10319 (N_10319,N_6525,N_6077);
nor U10320 (N_10320,N_5371,N_7507);
and U10321 (N_10321,N_7156,N_6652);
xor U10322 (N_10322,N_8772,N_8062);
xor U10323 (N_10323,N_6520,N_6463);
xor U10324 (N_10324,N_8036,N_6789);
or U10325 (N_10325,N_6821,N_7042);
nor U10326 (N_10326,N_5347,N_6908);
nor U10327 (N_10327,N_6177,N_6540);
nor U10328 (N_10328,N_7732,N_7277);
nor U10329 (N_10329,N_5858,N_5381);
or U10330 (N_10330,N_9736,N_5683);
nand U10331 (N_10331,N_5393,N_6551);
or U10332 (N_10332,N_7489,N_5657);
xnor U10333 (N_10333,N_6340,N_8155);
or U10334 (N_10334,N_5654,N_6220);
or U10335 (N_10335,N_7154,N_8005);
nor U10336 (N_10336,N_7016,N_8534);
and U10337 (N_10337,N_5309,N_9604);
nor U10338 (N_10338,N_7425,N_8039);
nor U10339 (N_10339,N_9348,N_8618);
or U10340 (N_10340,N_6454,N_9968);
nand U10341 (N_10341,N_6215,N_5949);
nand U10342 (N_10342,N_8219,N_8422);
xnor U10343 (N_10343,N_9182,N_8502);
nand U10344 (N_10344,N_6602,N_5432);
nand U10345 (N_10345,N_9258,N_9635);
or U10346 (N_10346,N_5602,N_9138);
xor U10347 (N_10347,N_5638,N_8515);
or U10348 (N_10348,N_6565,N_6516);
or U10349 (N_10349,N_7143,N_7116);
and U10350 (N_10350,N_8166,N_8439);
and U10351 (N_10351,N_7753,N_5446);
nor U10352 (N_10352,N_5264,N_6460);
nand U10353 (N_10353,N_5227,N_9638);
xor U10354 (N_10354,N_6094,N_5606);
nand U10355 (N_10355,N_9385,N_8455);
or U10356 (N_10356,N_5778,N_5424);
xnor U10357 (N_10357,N_8382,N_8188);
nor U10358 (N_10358,N_8734,N_7605);
xnor U10359 (N_10359,N_5733,N_7168);
and U10360 (N_10360,N_7330,N_7175);
xnor U10361 (N_10361,N_7591,N_8220);
and U10362 (N_10362,N_8184,N_7020);
nor U10363 (N_10363,N_6819,N_6259);
nor U10364 (N_10364,N_5877,N_7656);
nand U10365 (N_10365,N_8628,N_5772);
and U10366 (N_10366,N_6349,N_7729);
xnor U10367 (N_10367,N_5383,N_8945);
xor U10368 (N_10368,N_5998,N_5356);
xor U10369 (N_10369,N_6466,N_8657);
and U10370 (N_10370,N_8804,N_6452);
nor U10371 (N_10371,N_7659,N_6788);
or U10372 (N_10372,N_9179,N_5952);
or U10373 (N_10373,N_5078,N_7950);
nand U10374 (N_10374,N_7654,N_9611);
and U10375 (N_10375,N_7238,N_8169);
or U10376 (N_10376,N_8812,N_8396);
xnor U10377 (N_10377,N_7674,N_9648);
and U10378 (N_10378,N_7136,N_5836);
nand U10379 (N_10379,N_6529,N_7968);
nor U10380 (N_10380,N_5751,N_8448);
xnor U10381 (N_10381,N_6960,N_9887);
nor U10382 (N_10382,N_8044,N_8495);
xnor U10383 (N_10383,N_8582,N_5089);
nor U10384 (N_10384,N_6506,N_8034);
nor U10385 (N_10385,N_7677,N_6932);
xor U10386 (N_10386,N_7241,N_6576);
nor U10387 (N_10387,N_9438,N_8689);
nand U10388 (N_10388,N_7046,N_7010);
nor U10389 (N_10389,N_7269,N_5273);
nor U10390 (N_10390,N_9373,N_9435);
and U10391 (N_10391,N_6056,N_6892);
nand U10392 (N_10392,N_5919,N_9405);
or U10393 (N_10393,N_7700,N_9403);
and U10394 (N_10394,N_5854,N_6795);
nor U10395 (N_10395,N_5682,N_7978);
and U10396 (N_10396,N_8314,N_7725);
and U10397 (N_10397,N_5109,N_8715);
or U10398 (N_10398,N_6841,N_7943);
or U10399 (N_10399,N_9436,N_8225);
xor U10400 (N_10400,N_8626,N_5047);
and U10401 (N_10401,N_9053,N_7487);
nand U10402 (N_10402,N_6513,N_8872);
and U10403 (N_10403,N_6666,N_5221);
or U10404 (N_10404,N_8996,N_8517);
and U10405 (N_10405,N_7347,N_6329);
or U10406 (N_10406,N_9264,N_5857);
xnor U10407 (N_10407,N_6415,N_9819);
nand U10408 (N_10408,N_9977,N_5299);
xnor U10409 (N_10409,N_8403,N_9060);
xnor U10410 (N_10410,N_5254,N_9411);
and U10411 (N_10411,N_5113,N_8743);
and U10412 (N_10412,N_6969,N_7017);
nor U10413 (N_10413,N_7570,N_8962);
nor U10414 (N_10414,N_9883,N_5988);
or U10415 (N_10415,N_9063,N_9806);
and U10416 (N_10416,N_7421,N_9647);
and U10417 (N_10417,N_7069,N_7179);
or U10418 (N_10418,N_7930,N_8400);
nor U10419 (N_10419,N_9419,N_8856);
xnor U10420 (N_10420,N_6626,N_7207);
or U10421 (N_10421,N_8827,N_9686);
and U10422 (N_10422,N_6979,N_7111);
nor U10423 (N_10423,N_9320,N_9392);
nor U10424 (N_10424,N_7417,N_8793);
nor U10425 (N_10425,N_8700,N_6822);
nor U10426 (N_10426,N_8443,N_6697);
nor U10427 (N_10427,N_5520,N_5251);
and U10428 (N_10428,N_5317,N_5171);
or U10429 (N_10429,N_5642,N_9912);
or U10430 (N_10430,N_6046,N_7043);
and U10431 (N_10431,N_7349,N_7283);
xnor U10432 (N_10432,N_7479,N_9904);
and U10433 (N_10433,N_8671,N_8771);
nand U10434 (N_10434,N_7552,N_5314);
and U10435 (N_10435,N_9576,N_8881);
nand U10436 (N_10436,N_6342,N_7368);
or U10437 (N_10437,N_6162,N_6972);
xor U10438 (N_10438,N_6957,N_9058);
and U10439 (N_10439,N_6384,N_5138);
nand U10440 (N_10440,N_8635,N_6661);
xnor U10441 (N_10441,N_6470,N_5486);
and U10442 (N_10442,N_6061,N_9154);
xor U10443 (N_10443,N_6113,N_9126);
nor U10444 (N_10444,N_9971,N_5250);
nand U10445 (N_10445,N_9152,N_9353);
nand U10446 (N_10446,N_6556,N_7373);
nand U10447 (N_10447,N_6115,N_7152);
nand U10448 (N_10448,N_5908,N_8059);
xnor U10449 (N_10449,N_8325,N_8148);
or U10450 (N_10450,N_8199,N_8577);
nor U10451 (N_10451,N_8251,N_8998);
xor U10452 (N_10452,N_5892,N_9443);
xnor U10453 (N_10453,N_8106,N_7337);
xnor U10454 (N_10454,N_7052,N_7364);
xor U10455 (N_10455,N_9008,N_5717);
or U10456 (N_10456,N_9383,N_5006);
nor U10457 (N_10457,N_5633,N_5029);
xnor U10458 (N_10458,N_8388,N_6920);
nand U10459 (N_10459,N_6807,N_8412);
xor U10460 (N_10460,N_5240,N_9809);
and U10461 (N_10461,N_6428,N_6900);
nor U10462 (N_10462,N_7795,N_8737);
nand U10463 (N_10463,N_5521,N_8828);
xor U10464 (N_10464,N_7528,N_8058);
nand U10465 (N_10465,N_7334,N_7569);
xnor U10466 (N_10466,N_9776,N_7922);
or U10467 (N_10467,N_6098,N_7220);
or U10468 (N_10468,N_5829,N_5162);
and U10469 (N_10469,N_5134,N_9653);
or U10470 (N_10470,N_5761,N_9370);
and U10471 (N_10471,N_7520,N_7908);
nand U10472 (N_10472,N_9870,N_7550);
nand U10473 (N_10473,N_9573,N_7548);
nand U10474 (N_10474,N_6124,N_5618);
and U10475 (N_10475,N_7717,N_6103);
and U10476 (N_10476,N_9449,N_6981);
nor U10477 (N_10477,N_9208,N_9190);
xor U10478 (N_10478,N_8556,N_7483);
nor U10479 (N_10479,N_8145,N_8370);
nand U10480 (N_10480,N_8922,N_8554);
and U10481 (N_10481,N_8539,N_7384);
and U10482 (N_10482,N_6874,N_8099);
nand U10483 (N_10483,N_6174,N_5157);
nand U10484 (N_10484,N_5884,N_5204);
xor U10485 (N_10485,N_5624,N_7374);
nor U10486 (N_10486,N_9941,N_7442);
xnor U10487 (N_10487,N_9297,N_7184);
nand U10488 (N_10488,N_9953,N_6696);
nand U10489 (N_10489,N_5989,N_6278);
nor U10490 (N_10490,N_8533,N_6060);
nand U10491 (N_10491,N_6299,N_5376);
or U10492 (N_10492,N_7387,N_9651);
and U10493 (N_10493,N_9279,N_8389);
nand U10494 (N_10494,N_8611,N_6750);
xor U10495 (N_10495,N_9659,N_7919);
nor U10496 (N_10496,N_9973,N_5795);
nand U10497 (N_10497,N_7576,N_7481);
nor U10498 (N_10498,N_9885,N_7612);
xnor U10499 (N_10499,N_6541,N_6361);
and U10500 (N_10500,N_8693,N_8444);
nor U10501 (N_10501,N_9584,N_7408);
and U10502 (N_10502,N_6280,N_6642);
or U10503 (N_10503,N_8951,N_9619);
or U10504 (N_10504,N_9597,N_5420);
nor U10505 (N_10505,N_6982,N_7474);
or U10506 (N_10506,N_7780,N_8710);
nand U10507 (N_10507,N_5337,N_9900);
and U10508 (N_10508,N_8295,N_6588);
xor U10509 (N_10509,N_5659,N_9022);
nand U10510 (N_10510,N_8230,N_6169);
xnor U10511 (N_10511,N_7150,N_5814);
nand U10512 (N_10512,N_7687,N_5107);
and U10513 (N_10513,N_5439,N_7495);
and U10514 (N_10514,N_7931,N_8323);
or U10515 (N_10515,N_6126,N_6096);
nand U10516 (N_10516,N_5958,N_9799);
or U10517 (N_10517,N_5484,N_8264);
and U10518 (N_10518,N_7665,N_8525);
nand U10519 (N_10519,N_5985,N_6546);
and U10520 (N_10520,N_8978,N_5759);
and U10521 (N_10521,N_6921,N_6208);
or U10522 (N_10522,N_7718,N_8375);
or U10523 (N_10523,N_8740,N_6471);
or U10524 (N_10524,N_5851,N_9516);
xor U10525 (N_10525,N_8730,N_6097);
and U10526 (N_10526,N_9029,N_9276);
nand U10527 (N_10527,N_5838,N_9471);
or U10528 (N_10528,N_8999,N_6199);
nor U10529 (N_10529,N_9055,N_9151);
nand U10530 (N_10530,N_9427,N_6376);
nand U10531 (N_10531,N_9423,N_5259);
nand U10532 (N_10532,N_5531,N_6371);
xor U10533 (N_10533,N_7253,N_8566);
nand U10534 (N_10534,N_7405,N_5558);
nor U10535 (N_10535,N_8153,N_9537);
nor U10536 (N_10536,N_7170,N_7926);
nand U10537 (N_10537,N_5362,N_5596);
nor U10538 (N_10538,N_8486,N_9564);
xnor U10539 (N_10539,N_9178,N_6748);
and U10540 (N_10540,N_7574,N_9224);
nor U10541 (N_10541,N_8568,N_5088);
or U10542 (N_10542,N_9204,N_5027);
nor U10543 (N_10543,N_8163,N_7800);
nand U10544 (N_10544,N_8759,N_5747);
and U10545 (N_10545,N_5957,N_8110);
nand U10546 (N_10546,N_9113,N_8742);
nor U10547 (N_10547,N_8256,N_5178);
xor U10548 (N_10548,N_6677,N_6441);
nand U10549 (N_10549,N_7279,N_6586);
xor U10550 (N_10550,N_7772,N_6018);
and U10551 (N_10551,N_5490,N_5460);
nor U10552 (N_10552,N_7686,N_7103);
xnor U10553 (N_10553,N_7530,N_5656);
or U10554 (N_10554,N_6503,N_7983);
and U10555 (N_10555,N_8031,N_9400);
nor U10556 (N_10556,N_9768,N_8981);
xnor U10557 (N_10557,N_9315,N_7015);
or U10558 (N_10558,N_8320,N_5626);
nand U10559 (N_10559,N_5781,N_8862);
xnor U10560 (N_10560,N_8175,N_5607);
xnor U10561 (N_10561,N_9800,N_7206);
or U10562 (N_10562,N_8047,N_8493);
nand U10563 (N_10563,N_6811,N_8801);
and U10564 (N_10564,N_9474,N_7701);
nand U10565 (N_10565,N_9623,N_7115);
nand U10566 (N_10566,N_8081,N_7345);
and U10567 (N_10567,N_5079,N_8865);
or U10568 (N_10568,N_9632,N_8469);
and U10569 (N_10569,N_9514,N_9020);
xnor U10570 (N_10570,N_6636,N_9987);
xor U10571 (N_10571,N_5731,N_7249);
nor U10572 (N_10572,N_7388,N_5505);
nor U10573 (N_10573,N_9072,N_9199);
xnor U10574 (N_10574,N_6885,N_6171);
nor U10575 (N_10575,N_7580,N_5945);
nor U10576 (N_10576,N_5469,N_9101);
xor U10577 (N_10577,N_7409,N_5035);
xor U10578 (N_10578,N_6784,N_8160);
or U10579 (N_10579,N_5617,N_9233);
xor U10580 (N_10580,N_7323,N_7366);
or U10581 (N_10581,N_5557,N_5445);
nand U10582 (N_10582,N_8273,N_5594);
nand U10583 (N_10583,N_8744,N_8458);
and U10584 (N_10584,N_5070,N_5323);
nor U10585 (N_10585,N_6155,N_7980);
nand U10586 (N_10586,N_5501,N_9660);
xor U10587 (N_10587,N_5104,N_5051);
xor U10588 (N_10588,N_9649,N_8394);
xnor U10589 (N_10589,N_8311,N_6198);
or U10590 (N_10590,N_9575,N_6269);
and U10591 (N_10591,N_8703,N_6107);
xnor U10592 (N_10592,N_6358,N_9200);
nand U10593 (N_10593,N_7669,N_8417);
nand U10594 (N_10594,N_6119,N_8930);
xor U10595 (N_10595,N_9503,N_9026);
nand U10596 (N_10596,N_8779,N_8348);
nand U10597 (N_10597,N_8956,N_7794);
and U10598 (N_10598,N_5931,N_8222);
xor U10599 (N_10599,N_8535,N_5161);
nor U10600 (N_10600,N_5327,N_6436);
nor U10601 (N_10601,N_7174,N_6759);
nand U10602 (N_10602,N_5639,N_5425);
nor U10603 (N_10603,N_7523,N_5871);
xor U10604 (N_10604,N_6706,N_8133);
nand U10605 (N_10605,N_9929,N_8864);
and U10606 (N_10606,N_8029,N_5665);
or U10607 (N_10607,N_8839,N_7453);
or U10608 (N_10608,N_8091,N_9881);
nand U10609 (N_10609,N_9450,N_8102);
and U10610 (N_10610,N_6196,N_8624);
or U10611 (N_10611,N_9300,N_7429);
or U10612 (N_10612,N_7525,N_7177);
nor U10613 (N_10613,N_8521,N_6616);
and U10614 (N_10614,N_5698,N_5033);
and U10615 (N_10615,N_5196,N_7455);
or U10616 (N_10616,N_8123,N_7491);
or U10617 (N_10617,N_7161,N_8992);
xnor U10618 (N_10618,N_7290,N_5496);
and U10619 (N_10619,N_8385,N_9913);
nor U10620 (N_10620,N_8200,N_9479);
and U10621 (N_10621,N_5832,N_8874);
or U10622 (N_10622,N_5480,N_5366);
and U10623 (N_10623,N_8917,N_5668);
or U10624 (N_10624,N_6099,N_8645);
xor U10625 (N_10625,N_9456,N_7697);
nor U10626 (N_10626,N_9948,N_7932);
nor U10627 (N_10627,N_9779,N_9046);
or U10628 (N_10628,N_6809,N_8904);
and U10629 (N_10629,N_5707,N_9952);
xor U10630 (N_10630,N_9976,N_6055);
nand U10631 (N_10631,N_6287,N_9444);
or U10632 (N_10632,N_9538,N_9007);
and U10633 (N_10633,N_9078,N_7755);
or U10634 (N_10634,N_8731,N_5693);
nor U10635 (N_10635,N_8708,N_5252);
nor U10636 (N_10636,N_7477,N_5968);
or U10637 (N_10637,N_8543,N_5385);
and U10638 (N_10638,N_7806,N_7915);
nor U10639 (N_10639,N_6047,N_7285);
nand U10640 (N_10640,N_7558,N_9717);
nor U10641 (N_10641,N_9511,N_9967);
nand U10642 (N_10642,N_9501,N_5236);
or U10643 (N_10643,N_5956,N_7432);
and U10644 (N_10644,N_5470,N_6735);
xnor U10645 (N_10645,N_9566,N_9212);
and U10646 (N_10646,N_6741,N_7287);
nand U10647 (N_10647,N_5228,N_5436);
or U10648 (N_10648,N_7566,N_9122);
xnor U10649 (N_10649,N_5234,N_6147);
or U10650 (N_10650,N_5441,N_7825);
and U10651 (N_10651,N_7632,N_9316);
or U10652 (N_10652,N_6226,N_5865);
or U10653 (N_10653,N_8860,N_7726);
and U10654 (N_10654,N_9476,N_7935);
and U10655 (N_10655,N_5544,N_8158);
xnor U10656 (N_10656,N_8843,N_5255);
or U10657 (N_10657,N_7457,N_5072);
nand U10658 (N_10658,N_8299,N_5467);
nand U10659 (N_10659,N_6090,N_8590);
nand U10660 (N_10660,N_8677,N_8185);
or U10661 (N_10661,N_8987,N_6674);
or U10662 (N_10662,N_7126,N_7077);
nand U10663 (N_10663,N_7938,N_5031);
nor U10664 (N_10664,N_7085,N_6519);
xor U10665 (N_10665,N_5635,N_5492);
xor U10666 (N_10666,N_5282,N_7370);
xor U10667 (N_10667,N_5302,N_9234);
xor U10668 (N_10668,N_6104,N_7475);
and U10669 (N_10669,N_6728,N_6045);
nor U10670 (N_10670,N_9517,N_9942);
nor U10671 (N_10671,N_5205,N_9093);
nor U10672 (N_10672,N_7312,N_6849);
xor U10673 (N_10673,N_6133,N_9432);
nor U10674 (N_10674,N_9074,N_8274);
or U10675 (N_10675,N_5422,N_6679);
nor U10676 (N_10676,N_7501,N_7597);
or U10677 (N_10677,N_5519,N_9037);
nor U10678 (N_10678,N_8880,N_7247);
or U10679 (N_10679,N_5784,N_5713);
and U10680 (N_10680,N_7929,N_9979);
nor U10681 (N_10681,N_8935,N_8381);
and U10682 (N_10682,N_5997,N_7288);
and U10683 (N_10683,N_8907,N_7340);
or U10684 (N_10684,N_8545,N_9355);
and U10685 (N_10685,N_6894,N_6181);
xnor U10686 (N_10686,N_7551,N_6031);
nand U10687 (N_10687,N_7801,N_9109);
nor U10688 (N_10688,N_9949,N_7060);
or U10689 (N_10689,N_9525,N_7736);
nor U10690 (N_10690,N_6803,N_9783);
nand U10691 (N_10691,N_7071,N_7221);
or U10692 (N_10692,N_5209,N_5127);
xor U10693 (N_10693,N_8272,N_7333);
and U10694 (N_10694,N_7579,N_6504);
nor U10695 (N_10695,N_6901,N_8928);
or U10696 (N_10696,N_6648,N_5561);
xor U10697 (N_10697,N_6598,N_8324);
nand U10698 (N_10698,N_8173,N_7321);
and U10699 (N_10699,N_5727,N_8617);
xor U10700 (N_10700,N_9302,N_5343);
xnor U10701 (N_10701,N_8594,N_9465);
and U10702 (N_10702,N_9455,N_9683);
or U10703 (N_10703,N_9524,N_7893);
xor U10704 (N_10704,N_7397,N_6481);
nor U10705 (N_10705,N_8406,N_9067);
and U10706 (N_10706,N_8283,N_7414);
nand U10707 (N_10707,N_9692,N_7182);
or U10708 (N_10708,N_9011,N_6695);
and U10709 (N_10709,N_7313,N_8695);
and U10710 (N_10710,N_6407,N_5791);
or U10711 (N_10711,N_7846,N_9784);
nor U10712 (N_10712,N_5380,N_7315);
nor U10713 (N_10713,N_8204,N_5455);
nor U10714 (N_10714,N_6656,N_9554);
or U10715 (N_10715,N_9112,N_6427);
or U10716 (N_10716,N_6937,N_9669);
nand U10717 (N_10717,N_6041,N_6188);
nor U10718 (N_10718,N_7996,N_6241);
and U10719 (N_10719,N_8078,N_9995);
xor U10720 (N_10720,N_9727,N_6778);
or U10721 (N_10721,N_5023,N_9879);
nor U10722 (N_10722,N_6072,N_8705);
and U10723 (N_10723,N_9205,N_6444);
xnor U10724 (N_10724,N_7611,N_6952);
nor U10725 (N_10725,N_5615,N_8454);
and U10726 (N_10726,N_8511,N_9430);
nand U10727 (N_10727,N_7672,N_7505);
or U10728 (N_10728,N_6433,N_6945);
nand U10729 (N_10729,N_8410,N_6563);
and U10730 (N_10730,N_9188,N_5177);
or U10731 (N_10731,N_9426,N_6476);
nor U10732 (N_10732,N_5429,N_8810);
or U10733 (N_10733,N_5289,N_6688);
nor U10734 (N_10734,N_9452,N_5349);
nor U10735 (N_10735,N_7446,N_9472);
and U10736 (N_10736,N_6738,N_8046);
xnor U10737 (N_10737,N_6347,N_9789);
nand U10738 (N_10738,N_6777,N_7928);
nor U10739 (N_10739,N_7470,N_5325);
and U10740 (N_10740,N_7842,N_8399);
xor U10741 (N_10741,N_6212,N_9117);
or U10742 (N_10742,N_6637,N_9732);
nand U10743 (N_10743,N_6745,N_6423);
xnor U10744 (N_10744,N_6792,N_8305);
and U10745 (N_10745,N_8189,N_5444);
or U10746 (N_10746,N_7164,N_9731);
xor U10747 (N_10747,N_5335,N_9475);
and U10748 (N_10748,N_9380,N_7622);
xnor U10749 (N_10749,N_9467,N_8910);
and U10750 (N_10750,N_8831,N_8321);
and U10751 (N_10751,N_5472,N_6968);
xor U10752 (N_10752,N_8507,N_8409);
xnor U10753 (N_10753,N_5370,N_8023);
and U10754 (N_10754,N_9997,N_5581);
nor U10755 (N_10755,N_6027,N_5697);
nand U10756 (N_10756,N_8929,N_7675);
nor U10757 (N_10757,N_7571,N_7531);
and U10758 (N_10758,N_7563,N_6496);
xor U10759 (N_10759,N_8678,N_9349);
xor U10760 (N_10760,N_5372,N_8209);
nor U10761 (N_10761,N_5040,N_6896);
nor U10762 (N_10762,N_8482,N_8352);
xor U10763 (N_10763,N_5306,N_5194);
or U10764 (N_10764,N_6465,N_7704);
nor U10765 (N_10765,N_6144,N_8587);
xor U10766 (N_10766,N_9482,N_7361);
nand U10767 (N_10767,N_8627,N_6377);
nor U10768 (N_10768,N_8090,N_5293);
or U10769 (N_10769,N_7827,N_7616);
xor U10770 (N_10770,N_6175,N_9852);
or U10771 (N_10771,N_5050,N_5019);
and U10772 (N_10772,N_8407,N_5680);
xnor U10773 (N_10773,N_7140,N_6594);
xor U10774 (N_10774,N_6569,N_9454);
or U10775 (N_10775,N_8353,N_6521);
or U10776 (N_10776,N_6609,N_6393);
and U10777 (N_10777,N_6638,N_9327);
or U10778 (N_10778,N_5670,N_7655);
nand U10779 (N_10779,N_5433,N_7748);
nor U10780 (N_10780,N_9721,N_5573);
and U10781 (N_10781,N_8319,N_7004);
xnor U10782 (N_10782,N_5770,N_7203);
nand U10783 (N_10783,N_6911,N_8014);
nand U10784 (N_10784,N_9808,N_9802);
xor U10785 (N_10785,N_6028,N_6232);
xor U10786 (N_10786,N_9928,N_8236);
nor U10787 (N_10787,N_5002,N_8009);
and U10788 (N_10788,N_8925,N_8873);
and U10789 (N_10789,N_6266,N_6780);
and U10790 (N_10790,N_6462,N_9757);
or U10791 (N_10791,N_7331,N_7720);
xor U10792 (N_10792,N_5755,N_5767);
xnor U10793 (N_10793,N_9753,N_7527);
or U10794 (N_10794,N_6325,N_9811);
or U10795 (N_10795,N_9630,N_9986);
nor U10796 (N_10796,N_5286,N_5967);
or U10797 (N_10797,N_9391,N_9951);
nor U10798 (N_10798,N_9652,N_6966);
xnor U10799 (N_10799,N_7843,N_6526);
and U10800 (N_10800,N_6253,N_5671);
nand U10801 (N_10801,N_7740,N_5125);
xor U10802 (N_10802,N_9710,N_5540);
xor U10803 (N_10803,N_5825,N_6201);
nand U10804 (N_10804,N_7991,N_5493);
xnor U10805 (N_10805,N_9620,N_5565);
nor U10806 (N_10806,N_9061,N_5775);
and U10807 (N_10807,N_8465,N_7113);
or U10808 (N_10808,N_5344,N_5940);
nand U10809 (N_10809,N_9064,N_9098);
and U10810 (N_10810,N_7959,N_8268);
nand U10811 (N_10811,N_5080,N_7920);
nand U10812 (N_10812,N_9163,N_7002);
and U10813 (N_10813,N_5239,N_7599);
nor U10814 (N_10814,N_7092,N_6271);
or U10815 (N_10815,N_9285,N_9894);
nand U10816 (N_10816,N_7652,N_9641);
nor U10817 (N_10817,N_8318,N_5701);
nor U10818 (N_10818,N_7715,N_8681);
xor U10819 (N_10819,N_9079,N_8765);
or U10820 (N_10820,N_5653,N_5878);
nand U10821 (N_10821,N_9369,N_8056);
xor U10822 (N_10822,N_5922,N_7023);
nor U10823 (N_10823,N_7593,N_9485);
xnor U10824 (N_10824,N_5875,N_7447);
and U10825 (N_10825,N_6399,N_8480);
xor U10826 (N_10826,N_5900,N_8397);
and U10827 (N_10827,N_8038,N_7989);
or U10828 (N_10828,N_7775,N_9492);
and U10829 (N_10829,N_7741,N_6258);
nand U10830 (N_10830,N_9637,N_9329);
and U10831 (N_10831,N_5435,N_7329);
or U10832 (N_10832,N_7496,N_9161);
or U10833 (N_10833,N_5903,N_9557);
or U10834 (N_10834,N_5136,N_5200);
or U10835 (N_10835,N_8947,N_8271);
nor U10836 (N_10836,N_9044,N_8214);
nand U10837 (N_10837,N_5790,N_7653);
and U10838 (N_10838,N_6034,N_6650);
or U10839 (N_10839,N_8988,N_8282);
nand U10840 (N_10840,N_5068,N_5231);
or U10841 (N_10841,N_7875,N_5400);
nand U10842 (N_10842,N_8020,N_5198);
xor U10843 (N_10843,N_5819,N_5651);
nand U10844 (N_10844,N_6145,N_7584);
or U10845 (N_10845,N_7856,N_5324);
nor U10846 (N_10846,N_8372,N_7840);
nor U10847 (N_10847,N_6319,N_9704);
nand U10848 (N_10848,N_6121,N_6085);
nor U10849 (N_10849,N_6069,N_7488);
nor U10850 (N_10850,N_9488,N_5394);
or U10851 (N_10851,N_5398,N_6032);
or U10852 (N_10852,N_5545,N_7961);
nand U10853 (N_10853,N_9751,N_8387);
xor U10854 (N_10854,N_9013,N_7439);
nor U10855 (N_10855,N_7639,N_7271);
xor U10856 (N_10856,N_7214,N_7641);
or U10857 (N_10857,N_9582,N_7631);
or U10858 (N_10858,N_8234,N_9201);
xnor U10859 (N_10859,N_7378,N_8440);
nand U10860 (N_10860,N_5996,N_7877);
nand U10861 (N_10861,N_7625,N_6417);
and U10862 (N_10862,N_5813,N_5297);
and U10863 (N_10863,N_6019,N_9498);
nand U10864 (N_10864,N_7380,N_5925);
nand U10865 (N_10865,N_5757,N_6089);
xor U10866 (N_10866,N_7796,N_5091);
nand U10867 (N_10867,N_8775,N_9962);
xnor U10868 (N_10868,N_9608,N_6225);
xor U10869 (N_10869,N_8722,N_8634);
nand U10870 (N_10870,N_5587,N_9805);
xor U10871 (N_10871,N_9634,N_9446);
and U10872 (N_10872,N_5525,N_9102);
or U10873 (N_10873,N_7033,N_6016);
xnor U10874 (N_10874,N_5974,N_5184);
and U10875 (N_10875,N_7751,N_6593);
nor U10876 (N_10876,N_5987,N_6036);
xor U10877 (N_10877,N_8421,N_9157);
or U10878 (N_10878,N_7308,N_9032);
or U10879 (N_10879,N_5962,N_9433);
or U10880 (N_10880,N_5896,N_9715);
xnor U10881 (N_10881,N_6468,N_6701);
or U10882 (N_10882,N_7714,N_6779);
and U10883 (N_10883,N_7832,N_5413);
nor U10884 (N_10884,N_5308,N_6234);
nor U10885 (N_10885,N_6412,N_5806);
xor U10886 (N_10886,N_8076,N_5005);
or U10887 (N_10887,N_5528,N_8989);
nor U10888 (N_10888,N_9092,N_5663);
nand U10889 (N_10889,N_9933,N_8682);
nand U10890 (N_10890,N_8363,N_7749);
nor U10891 (N_10891,N_9197,N_8340);
or U10892 (N_10892,N_6681,N_9733);
or U10893 (N_10893,N_6997,N_6628);
nor U10894 (N_10894,N_9057,N_7424);
nand U10895 (N_10895,N_9095,N_8615);
or U10896 (N_10896,N_9237,N_6146);
and U10897 (N_10897,N_9415,N_6663);
and U10898 (N_10898,N_9886,N_9909);
and U10899 (N_10899,N_7577,N_5199);
nand U10900 (N_10900,N_6043,N_8629);
nor U10901 (N_10901,N_9593,N_7621);
xnor U10902 (N_10902,N_7284,N_8540);
nor U10903 (N_10903,N_9902,N_8304);
and U10904 (N_10904,N_6856,N_6172);
nand U10905 (N_10905,N_7902,N_7643);
nor U10906 (N_10906,N_6622,N_8605);
or U10907 (N_10907,N_5320,N_5452);
nand U10908 (N_10908,N_5794,N_9235);
xnor U10909 (N_10909,N_5296,N_8541);
xor U10910 (N_10910,N_9936,N_7703);
nor U10911 (N_10911,N_7147,N_5869);
and U10912 (N_10912,N_5880,N_9431);
or U10913 (N_10913,N_7438,N_8126);
xnor U10914 (N_10914,N_5386,N_7598);
or U10915 (N_10915,N_8415,N_8326);
and U10916 (N_10916,N_6543,N_9719);
and U10917 (N_10917,N_7835,N_5719);
and U10918 (N_10918,N_8776,N_5673);
xor U10919 (N_10919,N_7623,N_6410);
xor U10920 (N_10920,N_9705,N_5402);
nor U10921 (N_10921,N_8712,N_5028);
xor U10922 (N_10922,N_5655,N_5704);
nand U10923 (N_10923,N_5936,N_8649);
and U10924 (N_10924,N_5745,N_7153);
nand U10925 (N_10925,N_6591,N_8650);
nor U10926 (N_10926,N_6950,N_5053);
nand U10927 (N_10927,N_8132,N_9621);
and U10928 (N_10928,N_8179,N_9526);
xnor U10929 (N_10929,N_7859,N_6392);
and U10930 (N_10930,N_8769,N_6063);
or U10931 (N_10931,N_6721,N_6704);
nand U10932 (N_10932,N_6495,N_8728);
xor U10933 (N_10933,N_5649,N_6184);
or U10934 (N_10934,N_7232,N_9614);
xor U10935 (N_10935,N_6015,N_7314);
and U10936 (N_10936,N_9531,N_9943);
and U10937 (N_10937,N_6904,N_5774);
nand U10938 (N_10938,N_9769,N_7187);
or U10939 (N_10939,N_6512,N_5559);
nor U10940 (N_10940,N_9530,N_6013);
or U10941 (N_10941,N_7912,N_9916);
nand U10942 (N_10942,N_7193,N_7744);
nand U10943 (N_10943,N_6206,N_9760);
nor U10944 (N_10944,N_7532,N_5453);
nand U10945 (N_10945,N_6665,N_7681);
xnor U10946 (N_10946,N_7993,N_8496);
and U10947 (N_10947,N_7837,N_5036);
xor U10948 (N_10948,N_5166,N_9023);
xor U10949 (N_10949,N_5123,N_7178);
or U10950 (N_10950,N_8280,N_6757);
and U10951 (N_10951,N_6774,N_8760);
or U10952 (N_10952,N_6834,N_9378);
xor U10953 (N_10953,N_8702,N_8900);
nand U10954 (N_10954,N_9631,N_5210);
nand U10955 (N_10955,N_5011,N_6499);
nor U10956 (N_10956,N_8701,N_5955);
xor U10957 (N_10957,N_9693,N_6510);
nand U10958 (N_10958,N_6353,N_7339);
xnor U10959 (N_10959,N_8789,N_9080);
nand U10960 (N_10960,N_7752,N_6289);
or U10961 (N_10961,N_6323,N_7209);
and U10962 (N_10962,N_9059,N_9944);
nand U10963 (N_10963,N_6692,N_6397);
and U10964 (N_10964,N_8908,N_7460);
nand U10965 (N_10965,N_6273,N_7820);
nor U10966 (N_10966,N_6429,N_8303);
nand U10967 (N_10967,N_7181,N_8632);
nand U10968 (N_10968,N_9310,N_8655);
nor U10969 (N_10969,N_7942,N_6296);
xnor U10970 (N_10970,N_8337,N_5340);
and U10971 (N_10971,N_9505,N_7516);
nand U10972 (N_10972,N_7838,N_6003);
nor U10973 (N_10973,N_6837,N_6457);
nor U10974 (N_10974,N_9172,N_6413);
xnor U10975 (N_10975,N_6890,N_9354);
xnor U10976 (N_10976,N_9939,N_6523);
or U10977 (N_10977,N_6203,N_7246);
nand U10978 (N_10978,N_8139,N_5423);
or U10979 (N_10979,N_7773,N_6163);
nand U10980 (N_10980,N_9219,N_5013);
nor U10981 (N_10981,N_7860,N_8888);
xor U10982 (N_10982,N_5266,N_6459);
xnor U10983 (N_10983,N_5946,N_5928);
or U10984 (N_10984,N_5536,N_8007);
and U10985 (N_10985,N_5143,N_8313);
or U10986 (N_10986,N_8067,N_9866);
nor U10987 (N_10987,N_6775,N_8994);
nor U10988 (N_10988,N_5616,N_7198);
nand U10989 (N_10989,N_8013,N_5992);
xnor U10990 (N_10990,N_7899,N_9323);
nand U10991 (N_10991,N_5249,N_8838);
and U10992 (N_10992,N_7784,N_9701);
nand U10993 (N_10993,N_8464,N_8802);
and U10994 (N_10994,N_7685,N_8167);
or U10995 (N_10995,N_8500,N_9317);
nand U10996 (N_10996,N_6005,N_8593);
and U10997 (N_10997,N_6180,N_7293);
nand U10998 (N_10998,N_9040,N_9959);
or U10999 (N_10999,N_8478,N_6646);
or U11000 (N_11000,N_9677,N_5246);
xor U11001 (N_11001,N_8246,N_8310);
nand U11002 (N_11002,N_9230,N_7808);
xnor U11003 (N_11003,N_8983,N_6088);
xor U11004 (N_11004,N_9691,N_5430);
xnor U11005 (N_11005,N_7586,N_7076);
nand U11006 (N_11006,N_8263,N_6173);
or U11007 (N_11007,N_5622,N_6022);
nand U11008 (N_11008,N_5564,N_5924);
nor U11009 (N_11009,N_9226,N_9569);
and U11010 (N_11010,N_8216,N_6838);
xnor U11011 (N_11011,N_5315,N_9305);
nor U11012 (N_11012,N_5728,N_7906);
xnor U11013 (N_11013,N_5510,N_9834);
xnor U11014 (N_11014,N_8049,N_6740);
xnor U11015 (N_11015,N_6294,N_8423);
or U11016 (N_11016,N_9286,N_6716);
or U11017 (N_11017,N_5661,N_7272);
nor U11018 (N_11018,N_7229,N_9236);
nand U11019 (N_11019,N_8287,N_7680);
xor U11020 (N_11020,N_6772,N_5442);
and U11021 (N_11021,N_5415,N_7375);
xor U11022 (N_11022,N_5692,N_6875);
nand U11023 (N_11023,N_5762,N_6364);
or U11024 (N_11024,N_5850,N_5710);
or U11025 (N_11025,N_8129,N_6401);
xnor U11026 (N_11026,N_6448,N_9922);
xnor U11027 (N_11027,N_9028,N_6848);
nand U11028 (N_11028,N_7490,N_7035);
xor U11029 (N_11029,N_8328,N_8416);
or U11030 (N_11030,N_9864,N_8694);
nor U11031 (N_11031,N_8845,N_7172);
xnor U11032 (N_11032,N_8356,N_9372);
or U11033 (N_11033,N_7044,N_5004);
or U11034 (N_11034,N_7430,N_5052);
nand U11035 (N_11035,N_5145,N_6639);
and U11036 (N_11036,N_8055,N_8885);
xnor U11037 (N_11037,N_8673,N_8171);
nand U11038 (N_11038,N_7864,N_6943);
and U11039 (N_11039,N_6307,N_5748);
nor U11040 (N_11040,N_7385,N_9610);
nand U11041 (N_11041,N_8764,N_6435);
and U11042 (N_11042,N_8142,N_6078);
nand U11043 (N_11043,N_6134,N_6580);
or U11044 (N_11044,N_5959,N_9845);
nor U11045 (N_11045,N_5567,N_7392);
and U11046 (N_11046,N_5060,N_7148);
or U11047 (N_11047,N_8733,N_8065);
nand U11048 (N_11048,N_8829,N_6366);
nor U11049 (N_11049,N_7900,N_6587);
xor U11050 (N_11050,N_5097,N_8651);
and U11051 (N_11051,N_6093,N_9189);
xnor U11052 (N_11052,N_5257,N_9847);
and U11053 (N_11053,N_8883,N_9709);
or U11054 (N_11054,N_8248,N_6729);
xnor U11055 (N_11055,N_8680,N_7440);
xnor U11056 (N_11056,N_5817,N_5292);
and U11057 (N_11057,N_6386,N_9281);
and U11058 (N_11058,N_5303,N_7629);
nand U11059 (N_11059,N_8470,N_5310);
nand U11060 (N_11060,N_6923,N_7628);
and U11061 (N_11061,N_6796,N_5995);
and U11062 (N_11062,N_7668,N_9183);
nor U11063 (N_11063,N_5001,N_7212);
and U11064 (N_11064,N_8069,N_8921);
nand U11065 (N_11065,N_9211,N_7038);
or U11066 (N_11066,N_8562,N_5853);
and U11067 (N_11067,N_9626,N_8644);
or U11068 (N_11068,N_6507,N_5930);
or U11069 (N_11069,N_9306,N_7413);
nand U11070 (N_11070,N_7320,N_6324);
nand U11071 (N_11071,N_9512,N_8349);
nor U11072 (N_11072,N_7955,N_8674);
or U11073 (N_11073,N_6195,N_9739);
nor U11074 (N_11074,N_5294,N_8919);
and U11075 (N_11075,N_9560,N_7826);
xnor U11076 (N_11076,N_6112,N_6878);
nor U11077 (N_11077,N_6257,N_8531);
xor U11078 (N_11078,N_6649,N_7219);
xnor U11079 (N_11079,N_8358,N_7804);
nand U11080 (N_11080,N_9294,N_7089);
nand U11081 (N_11081,N_7666,N_7861);
or U11082 (N_11082,N_9850,N_6348);
or U11083 (N_11083,N_9519,N_6455);
xor U11084 (N_11084,N_5100,N_8293);
or U11085 (N_11085,N_9983,N_8798);
xor U11086 (N_11086,N_9266,N_9445);
and U11087 (N_11087,N_5043,N_6871);
nand U11088 (N_11088,N_5841,N_6001);
or U11089 (N_11089,N_9175,N_5287);
nor U11090 (N_11090,N_5164,N_8120);
xor U11091 (N_11091,N_9195,N_8196);
and U11092 (N_11092,N_5975,N_6675);
xor U11093 (N_11093,N_5920,N_5319);
nor U11094 (N_11094,N_8720,N_9666);
nand U11095 (N_11095,N_5410,N_9827);
xor U11096 (N_11096,N_8863,N_8121);
and U11097 (N_11097,N_6482,N_9478);
or U11098 (N_11098,N_6012,N_5336);
nor U11099 (N_11099,N_9459,N_7464);
and U11100 (N_11100,N_6645,N_6010);
nor U11101 (N_11101,N_9570,N_7048);
nor U11102 (N_11102,N_5631,N_9685);
nor U11103 (N_11103,N_7698,N_9389);
nand U11104 (N_11104,N_5375,N_9714);
xor U11105 (N_11105,N_9410,N_8522);
or U11106 (N_11106,N_7169,N_7510);
nand U11107 (N_11107,N_7573,N_8141);
nor U11108 (N_11108,N_8210,N_7311);
nand U11109 (N_11109,N_8364,N_9740);
and U11110 (N_11110,N_8232,N_5904);
xor U11111 (N_11111,N_5572,N_8436);
nor U11112 (N_11112,N_6754,N_5810);
nand U11113 (N_11113,N_9742,N_9004);
xnor U11114 (N_11114,N_9868,N_8154);
xnor U11115 (N_11115,N_6437,N_7969);
nor U11116 (N_11116,N_9186,N_9539);
nor U11117 (N_11117,N_6139,N_5699);
or U11118 (N_11118,N_8205,N_8168);
nand U11119 (N_11119,N_8359,N_6389);
nand U11120 (N_11120,N_8490,N_8451);
and U11121 (N_11121,N_8616,N_7268);
and U11122 (N_11122,N_6532,N_9338);
xor U11123 (N_11123,N_8253,N_5628);
or U11124 (N_11124,N_9831,N_9990);
nor U11125 (N_11125,N_5032,N_9880);
nor U11126 (N_11126,N_7262,N_9613);
and U11127 (N_11127,N_5785,N_7739);
and U11128 (N_11128,N_8217,N_6655);
xor U11129 (N_11129,N_9707,N_6914);
xor U11130 (N_11130,N_8484,N_6431);
nor U11131 (N_11131,N_7607,N_5740);
and U11132 (N_11132,N_5634,N_8072);
and U11133 (N_11133,N_7114,N_5479);
or U11134 (N_11134,N_6464,N_7940);
or U11135 (N_11135,N_8195,N_9225);
or U11136 (N_11136,N_7845,N_8909);
and U11137 (N_11137,N_8411,N_9875);
nor U11138 (N_11138,N_8718,N_5541);
nor U11139 (N_11139,N_9615,N_7068);
xnor U11140 (N_11140,N_5506,N_8068);
and U11141 (N_11141,N_7400,N_8137);
nor U11142 (N_11142,N_6687,N_8923);
nand U11143 (N_11143,N_9390,N_8266);
nor U11144 (N_11144,N_5192,N_6852);
nor U11145 (N_11145,N_7335,N_9840);
nor U11146 (N_11146,N_9908,N_9523);
xnor U11147 (N_11147,N_8894,N_8647);
xnor U11148 (N_11148,N_9633,N_9357);
nand U11149 (N_11149,N_8218,N_7129);
nor U11150 (N_11150,N_6768,N_5623);
or U11151 (N_11151,N_8004,N_5856);
and U11152 (N_11152,N_7127,N_6210);
or U11153 (N_11153,N_8092,N_8269);
xnor U11154 (N_11154,N_6823,N_9180);
xnor U11155 (N_11155,N_7828,N_6425);
nor U11156 (N_11156,N_8183,N_6611);
and U11157 (N_11157,N_8276,N_7689);
nand U11158 (N_11158,N_8052,N_8054);
nor U11159 (N_11159,N_9534,N_6959);
and U11160 (N_11160,N_6238,N_5906);
nand U11161 (N_11161,N_9213,N_8898);
nor U11162 (N_11162,N_5746,N_7694);
and U11163 (N_11163,N_9974,N_8095);
nor U11164 (N_11164,N_9206,N_9655);
nor U11165 (N_11165,N_7967,N_5645);
nand U11166 (N_11166,N_5729,N_9105);
or U11167 (N_11167,N_9252,N_5122);
and U11168 (N_11168,N_8686,N_7243);
xnor U11169 (N_11169,N_5703,N_8621);
nor U11170 (N_11170,N_7102,N_7099);
and U11171 (N_11171,N_5156,N_7007);
xnor U11172 (N_11172,N_8884,N_8361);
or U11173 (N_11173,N_8854,N_6686);
nand U11174 (N_11174,N_9616,N_9568);
nor U11175 (N_11175,N_5180,N_9711);
xor U11176 (N_11176,N_7303,N_7823);
or U11177 (N_11177,N_9600,N_7678);
nand U11178 (N_11178,N_6106,N_6277);
xnor U11179 (N_11179,N_6630,N_9160);
and U11180 (N_11180,N_7360,N_7851);
nor U11181 (N_11181,N_9414,N_8223);
xnor U11182 (N_11182,N_6037,N_6667);
nor U11183 (N_11183,N_7070,N_9087);
nor U11184 (N_11184,N_9507,N_9009);
nand U11185 (N_11185,N_9957,N_8553);
nor U11186 (N_11186,N_7210,N_6128);
xor U11187 (N_11187,N_6717,N_9250);
nand U11188 (N_11188,N_9272,N_9394);
nand U11189 (N_11189,N_5098,N_7406);
nor U11190 (N_11190,N_7664,N_6424);
and U11191 (N_11191,N_8738,N_8602);
nor U11192 (N_11192,N_7945,N_7291);
xor U11193 (N_11193,N_9194,N_9283);
nor U11194 (N_11194,N_8557,N_9956);
nor U11195 (N_11195,N_6817,N_7567);
xor U11196 (N_11196,N_5408,N_5111);
nor U11197 (N_11197,N_5888,N_9086);
or U11198 (N_11198,N_8015,N_7006);
and U11199 (N_11199,N_8662,N_6362);
or U11200 (N_11200,N_8434,N_8452);
nand U11201 (N_11201,N_9318,N_6723);
and U11202 (N_11202,N_8243,N_7286);
xnor U11203 (N_11203,N_6847,N_7063);
or U11204 (N_11204,N_7001,N_7927);
nor U11205 (N_11205,N_7758,N_6021);
nor U11206 (N_11206,N_5146,N_5290);
and U11207 (N_11207,N_6770,N_9246);
or U11208 (N_11208,N_9483,N_8335);
nand U11209 (N_11209,N_7062,N_7036);
nand U11210 (N_11210,N_7393,N_7786);
or U11211 (N_11211,N_7419,N_6014);
or U11212 (N_11212,N_9362,N_8000);
or U11213 (N_11213,N_5304,N_7171);
or U11214 (N_11214,N_6873,N_7706);
xor U11215 (N_11215,N_5416,N_5207);
nand U11216 (N_11216,N_5862,N_7878);
or U11217 (N_11217,N_6396,N_8613);
or U11218 (N_11218,N_9018,N_8239);
or U11219 (N_11219,N_7670,N_7398);
nand U11220 (N_11220,N_8048,N_7724);
and U11221 (N_11221,N_5652,N_6483);
nand U11222 (N_11222,N_8117,N_8051);
nor U11223 (N_11223,N_9529,N_7587);
xnor U11224 (N_11224,N_6387,N_6166);
or U11225 (N_11225,N_5339,N_8152);
or U11226 (N_11226,N_5465,N_9723);
nand U11227 (N_11227,N_6771,N_6024);
nor U11228 (N_11228,N_8790,N_9307);
or U11229 (N_11229,N_5873,N_5660);
or U11230 (N_11230,N_6942,N_8419);
nor U11231 (N_11231,N_9654,N_7809);
nor U11232 (N_11232,N_8050,N_9119);
and U11233 (N_11233,N_8445,N_6346);
xor U11234 (N_11234,N_6458,N_7798);
nor U11235 (N_11235,N_8033,N_6829);
nor U11236 (N_11236,N_8561,N_7721);
or U11237 (N_11237,N_8584,N_8082);
xnor U11238 (N_11238,N_9407,N_7792);
nor U11239 (N_11239,N_6204,N_9047);
nand U11240 (N_11240,N_9169,N_6414);
nand U11241 (N_11241,N_5411,N_5556);
xor U11242 (N_11242,N_8698,N_6832);
nand U11243 (N_11243,N_5092,N_7186);
xnor U11244 (N_11244,N_7604,N_5669);
nor U11245 (N_11245,N_9490,N_6531);
and U11246 (N_11246,N_6105,N_9499);
xnor U11247 (N_11247,N_6722,N_8398);
nand U11248 (N_11248,N_7582,N_5265);
xor U11249 (N_11249,N_7082,N_7848);
xnor U11250 (N_11250,N_8518,N_8229);
nand U11251 (N_11251,N_5632,N_6991);
or U11252 (N_11252,N_5478,N_9628);
nand U11253 (N_11253,N_7690,N_8565);
xor U11254 (N_11254,N_9066,N_8032);
nor U11255 (N_11255,N_9216,N_6522);
and U11256 (N_11256,N_5641,N_9777);
xnor U11257 (N_11257,N_6862,N_9207);
nor U11258 (N_11258,N_8312,N_9548);
xnor U11259 (N_11259,N_6592,N_6379);
nand U11260 (N_11260,N_6373,N_9469);
xor U11261 (N_11261,N_7619,N_8254);
nor U11262 (N_11262,N_7923,N_6330);
xor U11263 (N_11263,N_6595,N_6644);
or U11264 (N_11264,N_8378,N_8667);
and U11265 (N_11265,N_5941,N_7514);
nor U11266 (N_11266,N_5326,N_9814);
and U11267 (N_11267,N_9843,N_6292);
or U11268 (N_11268,N_8855,N_6515);
and U11269 (N_11269,N_5233,N_9861);
nor U11270 (N_11270,N_8786,N_8782);
and U11271 (N_11271,N_5681,N_6866);
or U11272 (N_11272,N_8876,N_9599);
and U11273 (N_11273,N_5022,N_9049);
nor U11274 (N_11274,N_9425,N_6075);
or U11275 (N_11275,N_6606,N_6755);
xnor U11276 (N_11276,N_8315,N_5859);
nand U11277 (N_11277,N_7817,N_5102);
nand U11278 (N_11278,N_5793,N_7449);
xnor U11279 (N_11279,N_6933,N_5131);
nand U11280 (N_11280,N_5328,N_9906);
and U11281 (N_11281,N_7248,N_9867);
xor U11282 (N_11282,N_6320,N_8660);
xnor U11283 (N_11283,N_7594,N_8661);
xor U11284 (N_11284,N_9397,N_7924);
xor U11285 (N_11285,N_6264,N_8281);
and U11286 (N_11286,N_8685,N_6949);
or U11287 (N_11287,N_9412,N_8583);
nor U11288 (N_11288,N_7947,N_6550);
nand U11289 (N_11289,N_9447,N_8614);
nand U11290 (N_11290,N_6256,N_7815);
nor U11291 (N_11291,N_5511,N_5593);
and U11292 (N_11292,N_6073,N_7145);
nor U11293 (N_11293,N_5695,N_6062);
nor U11294 (N_11294,N_7167,N_7620);
xor U11295 (N_11295,N_9100,N_8709);
xnor U11296 (N_11296,N_9202,N_7517);
nand U11297 (N_11297,N_5474,N_8235);
xnor U11298 (N_11298,N_7555,N_7371);
nor U11299 (N_11299,N_7743,N_6168);
nor U11300 (N_11300,N_5674,N_7624);
nand U11301 (N_11301,N_5513,N_8084);
and U11302 (N_11302,N_7382,N_8260);
xnor U11303 (N_11303,N_5700,N_7418);
xor U11304 (N_11304,N_6992,N_5312);
nor U11305 (N_11305,N_7857,N_5473);
xnor U11306 (N_11306,N_8558,N_5758);
and U11307 (N_11307,N_9544,N_5756);
nand U11308 (N_11308,N_9622,N_6995);
and U11309 (N_11309,N_9893,N_8985);
and U11310 (N_11310,N_8974,N_7180);
and U11311 (N_11311,N_9463,N_6694);
nand U11312 (N_11312,N_6456,N_8113);
xnor U11313 (N_11313,N_5369,N_6352);
or U11314 (N_11314,N_6150,N_7194);
xor U11315 (N_11315,N_6141,N_6625);
nor U11316 (N_11316,N_9565,N_7757);
nand U11317 (N_11317,N_8683,N_9627);
and U11318 (N_11318,N_9365,N_6600);
xnor U11319 (N_11319,N_6426,N_5568);
nor U11320 (N_11320,N_7289,N_9803);
or U11321 (N_11321,N_7911,N_7356);
and U11322 (N_11322,N_5965,N_6338);
and U11323 (N_11323,N_6050,N_9148);
xor U11324 (N_11324,N_8848,N_5235);
xor U11325 (N_11325,N_8245,N_8203);
nor U11326 (N_11326,N_6493,N_9848);
nand U11327 (N_11327,N_6590,N_6530);
xnor U11328 (N_11328,N_6568,N_9437);
nor U11329 (N_11329,N_5353,N_9954);
nand U11330 (N_11330,N_7767,N_5406);
nor U11331 (N_11331,N_8066,N_9137);
nand U11332 (N_11332,N_7012,N_5650);
or U11333 (N_11333,N_9042,N_7245);
nor U11334 (N_11334,N_5191,N_9171);
nand U11335 (N_11335,N_9043,N_5417);
or U11336 (N_11336,N_5150,N_6187);
and U11337 (N_11337,N_9862,N_8623);
nor U11338 (N_11338,N_8294,N_9388);
xor U11339 (N_11339,N_6430,N_9607);
nor U11340 (N_11340,N_5999,N_5277);
and U11341 (N_11341,N_9865,N_6207);
and U11342 (N_11342,N_9551,N_9090);
and U11343 (N_11343,N_5769,N_9174);
nand U11344 (N_11344,N_8585,N_7963);
and U11345 (N_11345,N_5190,N_8853);
nand U11346 (N_11346,N_6477,N_6159);
xnor U11347 (N_11347,N_8637,N_9073);
nand U11348 (N_11348,N_7916,N_9629);
nand U11349 (N_11349,N_5580,N_5026);
and U11350 (N_11350,N_5921,N_6691);
nand U11351 (N_11351,N_6333,N_7377);
nand U11352 (N_11352,N_9496,N_7691);
nor U11353 (N_11353,N_6176,N_6913);
xnor U11354 (N_11354,N_5414,N_7556);
or U11355 (N_11355,N_5597,N_6641);
nand U11356 (N_11356,N_5675,N_8079);
nand U11357 (N_11357,N_6805,N_6247);
nor U11358 (N_11358,N_8902,N_5154);
nor U11359 (N_11359,N_9807,N_7322);
nand U11360 (N_11360,N_6194,N_6479);
or U11361 (N_11361,N_5397,N_5298);
nand U11362 (N_11362,N_7640,N_7627);
nand U11363 (N_11363,N_8298,N_7651);
xnor U11364 (N_11364,N_7045,N_7734);
and U11365 (N_11365,N_5061,N_9780);
nand U11366 (N_11366,N_8669,N_7056);
nor U11367 (N_11367,N_9595,N_7663);
nor U11368 (N_11368,N_5137,N_9417);
and U11369 (N_11369,N_9232,N_5459);
or U11370 (N_11370,N_6375,N_9146);
and U11371 (N_11371,N_8597,N_9860);
and U11372 (N_11372,N_6130,N_7524);
nand U11373 (N_11373,N_5188,N_9989);
and U11374 (N_11374,N_8563,N_7437);
or U11375 (N_11375,N_6501,N_7818);
nand U11376 (N_11376,N_5224,N_9343);
and U11377 (N_11377,N_6142,N_6566);
nor U11378 (N_11378,N_6251,N_5182);
nor U11379 (N_11379,N_6956,N_9592);
and U11380 (N_11380,N_6743,N_5181);
or U11381 (N_11381,N_5392,N_7711);
xnor U11382 (N_11382,N_8027,N_7614);
nand U11383 (N_11383,N_9842,N_6135);
nor U11384 (N_11384,N_6065,N_7642);
or U11385 (N_11385,N_9267,N_5275);
and U11386 (N_11386,N_7040,N_6548);
nand U11387 (N_11387,N_7199,N_9312);
or U11388 (N_11388,N_8278,N_9606);
or U11389 (N_11389,N_6318,N_8761);
nor U11390 (N_11390,N_9676,N_8473);
or U11391 (N_11391,N_9817,N_6048);
or U11392 (N_11392,N_8806,N_9497);
and U11393 (N_11393,N_5112,N_8021);
and U11394 (N_11394,N_9099,N_9326);
nor U11395 (N_11395,N_7716,N_7252);
nand U11396 (N_11396,N_6029,N_8161);
and U11397 (N_11397,N_8425,N_7982);
xnor U11398 (N_11398,N_5083,N_6971);
nor U11399 (N_11399,N_5483,N_9247);
xor U11400 (N_11400,N_7561,N_9903);
nand U11401 (N_11401,N_7683,N_9598);
nor U11402 (N_11402,N_9601,N_6042);
xnor U11403 (N_11403,N_9254,N_6485);
nand U11404 (N_11404,N_6794,N_9170);
or U11405 (N_11405,N_7601,N_8045);
and U11406 (N_11406,N_9935,N_5517);
nand U11407 (N_11407,N_7281,N_9675);
and U11408 (N_11408,N_6480,N_5288);
or U11409 (N_11409,N_6711,N_5504);
xnor U11410 (N_11410,N_6954,N_5990);
nand U11411 (N_11411,N_7155,N_6781);
nand U11412 (N_11412,N_7157,N_8706);
or U11413 (N_11413,N_5694,N_5120);
and U11414 (N_11414,N_5313,N_6231);
nor U11415 (N_11415,N_8475,N_9193);
nand U11416 (N_11416,N_8631,N_8690);
nand U11417 (N_11417,N_9014,N_5037);
nor U11418 (N_11418,N_9901,N_8471);
xor U11419 (N_11419,N_9221,N_9833);
nor U11420 (N_11420,N_6006,N_6660);
and U11421 (N_11421,N_6310,N_7862);
and U11422 (N_11422,N_7644,N_6368);
nor U11423 (N_11423,N_8575,N_7135);
nand U11424 (N_11424,N_5537,N_6929);
and U11425 (N_11425,N_9625,N_9682);
nor U11426 (N_11426,N_8198,N_6316);
nand U11427 (N_11427,N_6617,N_7890);
xnor U11428 (N_11428,N_5377,N_7093);
xor U11429 (N_11429,N_9743,N_5149);
xnor U11430 (N_11430,N_7266,N_6202);
or U11431 (N_11431,N_8746,N_7494);
nand U11432 (N_11432,N_7952,N_8506);
or U11433 (N_11433,N_9299,N_9001);
nand U11434 (N_11434,N_9958,N_5667);
nand U11435 (N_11435,N_7452,N_5732);
nand U11436 (N_11436,N_9434,N_7779);
nand U11437 (N_11437,N_6936,N_7061);
nor U11438 (N_11438,N_6864,N_9884);
or U11439 (N_11439,N_6213,N_6868);
nand U11440 (N_11440,N_8150,N_8749);
and U11441 (N_11441,N_9926,N_9371);
nor U11442 (N_11442,N_8941,N_8202);
and U11443 (N_11443,N_8333,N_6066);
or U11444 (N_11444,N_7326,N_7237);
or U11445 (N_11445,N_6058,N_9825);
nor U11446 (N_11446,N_7988,N_7498);
xor U11447 (N_11447,N_8472,N_7722);
or U11448 (N_11448,N_7872,N_5130);
nand U11449 (N_11449,N_9846,N_8976);
xor U11450 (N_11450,N_6547,N_6020);
xor U11451 (N_11451,N_8074,N_7047);
or U11452 (N_11452,N_9033,N_6337);
xor U11453 (N_11453,N_9153,N_5837);
nor U11454 (N_11454,N_9420,N_9136);
xnor U11455 (N_11455,N_8532,N_5056);
nor U11456 (N_11456,N_9129,N_7608);
nand U11457 (N_11457,N_6149,N_8316);
nor U11458 (N_11458,N_5116,N_9191);
and U11459 (N_11459,N_6702,N_6922);
xnor U11460 (N_11460,N_6312,N_6511);
xor U11461 (N_11461,N_9050,N_7816);
nor U11462 (N_11462,N_8879,N_5361);
nand U11463 (N_11463,N_5212,N_8244);
nor U11464 (N_11464,N_9680,N_5497);
nor U11465 (N_11465,N_5333,N_8721);
nor U11466 (N_11466,N_9116,N_9341);
nor U11467 (N_11467,N_6276,N_9718);
nor U11468 (N_11468,N_7545,N_9024);
and U11469 (N_11469,N_7165,N_6252);
and U11470 (N_11470,N_6946,N_6707);
nand U11471 (N_11471,N_7159,N_8805);
xnor U11472 (N_11472,N_6651,N_8002);
nand U11473 (N_11473,N_8995,N_7564);
and U11474 (N_11474,N_6994,N_5203);
xnor U11475 (N_11475,N_5562,N_6302);
nor U11476 (N_11476,N_5475,N_7359);
nor U11477 (N_11477,N_6980,N_5067);
xnor U11478 (N_11478,N_9923,N_8723);
xor U11479 (N_11479,N_6309,N_5905);
xor U11480 (N_11480,N_7191,N_9301);
xnor U11481 (N_11481,N_7117,N_5689);
or U11482 (N_11482,N_7975,N_9159);
xnor U11483 (N_11483,N_7836,N_9265);
nor U11484 (N_11484,N_9461,N_8300);
and U11485 (N_11485,N_7107,N_7011);
and U11486 (N_11486,N_8530,N_5447);
nand U11487 (N_11487,N_6261,N_7300);
xnor U11488 (N_11488,N_5268,N_8965);
xor U11489 (N_11489,N_8960,N_5768);
xor U11490 (N_11490,N_8094,N_6301);
and U11491 (N_11491,N_9439,N_8538);
and U11492 (N_11492,N_7658,N_8317);
nand U11493 (N_11493,N_5629,N_8713);
and U11494 (N_11494,N_8818,N_9931);
xnor U11495 (N_11495,N_9720,N_7540);
and U11496 (N_11496,N_6076,N_7166);
and U11497 (N_11497,N_9502,N_6132);
or U11498 (N_11498,N_8997,N_9775);
and U11499 (N_11499,N_8875,N_6388);
xor U11500 (N_11500,N_7769,N_9366);
nor U11501 (N_11501,N_7662,N_6938);
xor U11502 (N_11502,N_5374,N_7904);
and U11503 (N_11503,N_5891,N_6281);
xor U11504 (N_11504,N_5972,N_6209);
nand U11505 (N_11505,N_8912,N_6140);
nor U11506 (N_11506,N_7204,N_6762);
and U11507 (N_11507,N_8550,N_9821);
nand U11508 (N_11508,N_9513,N_7244);
nand U11509 (N_11509,N_8670,N_9969);
xnor U11510 (N_11510,N_7499,N_5454);
or U11511 (N_11511,N_5812,N_5542);
nor U11512 (N_11512,N_7709,N_7797);
or U11513 (N_11513,N_8018,N_5081);
and U11514 (N_11514,N_6439,N_8131);
and U11515 (N_11515,N_5586,N_9220);
nor U11516 (N_11516,N_8010,N_5495);
or U11517 (N_11517,N_8338,N_5933);
and U11518 (N_11518,N_8711,N_6610);
xnor U11519 (N_11519,N_6799,N_7014);
or U11520 (N_11520,N_6700,N_5969);
nor U11521 (N_11521,N_7325,N_9905);
or U11522 (N_11522,N_6804,N_9289);
and U11523 (N_11523,N_8697,N_6306);
and U11524 (N_11524,N_5886,N_5476);
xor U11525 (N_11525,N_8886,N_6400);
and U11526 (N_11526,N_7395,N_9874);
and U11527 (N_11527,N_7319,N_8920);
or U11528 (N_11528,N_8343,N_8542);
nand U11529 (N_11529,N_5284,N_5115);
or U11530 (N_11530,N_9495,N_8498);
xor U11531 (N_11531,N_8850,N_5901);
nor U11532 (N_11532,N_5160,N_6747);
nand U11533 (N_11533,N_5461,N_6886);
or U11534 (N_11534,N_9773,N_6751);
or U11535 (N_11535,N_5824,N_6767);
and U11536 (N_11536,N_8972,N_9387);
and U11537 (N_11537,N_9222,N_7348);
nor U11538 (N_11538,N_5148,N_8813);
or U11539 (N_11539,N_8134,N_8924);
xnor U11540 (N_11540,N_8834,N_9702);
xnor U11541 (N_11541,N_9546,N_9121);
and U11542 (N_11542,N_5984,N_9198);
xnor U11543 (N_11543,N_9489,N_7324);
xor U11544 (N_11544,N_6293,N_6411);
and U11545 (N_11545,N_9470,N_9413);
or U11546 (N_11546,N_6356,N_6394);
or U11547 (N_11547,N_5515,N_7468);
or U11548 (N_11548,N_9181,N_7830);
or U11549 (N_11549,N_5801,N_9114);
and U11550 (N_11550,N_9580,N_8351);
xnor U11551 (N_11551,N_9749,N_8140);
or U11552 (N_11552,N_5489,N_5087);
nor U11553 (N_11553,N_5468,N_9981);
or U11554 (N_11554,N_5373,N_9031);
xor U11555 (N_11555,N_9668,N_7833);
nand U11556 (N_11556,N_5571,N_6350);
or U11557 (N_11557,N_5274,N_6572);
nor U11558 (N_11558,N_5428,N_9259);
and U11559 (N_11559,N_7880,N_7226);
or U11560 (N_11560,N_5101,N_6843);
and U11561 (N_11561,N_6374,N_9346);
nand U11562 (N_11562,N_6930,N_9972);
xnor U11563 (N_11563,N_8476,N_5754);
nand U11564 (N_11564,N_9076,N_8395);
nand U11565 (N_11565,N_6143,N_8279);
nor U11566 (N_11566,N_8213,N_6690);
and U11567 (N_11567,N_6497,N_5139);
and U11568 (N_11568,N_8952,N_9325);
xor U11569 (N_11569,N_6327,N_7346);
xnor U11570 (N_11570,N_8797,N_9796);
xor U11571 (N_11571,N_5509,N_9899);
or U11572 (N_11572,N_6808,N_6961);
nand U11573 (N_11573,N_6536,N_5443);
and U11574 (N_11574,N_9645,N_9270);
xor U11575 (N_11575,N_9679,N_8289);
or U11576 (N_11576,N_7390,N_8428);
xor U11577 (N_11577,N_9187,N_7719);
and U11578 (N_11578,N_7917,N_5927);
nand U11579 (N_11579,N_5811,N_5846);
nor U11580 (N_11580,N_9955,N_6828);
nor U11581 (N_11581,N_8170,N_6643);
nand U11582 (N_11582,N_8570,N_8109);
nor U11583 (N_11583,N_7351,N_9750);
and U11584 (N_11584,N_8905,N_7867);
nor U11585 (N_11585,N_6189,N_8420);
xor U11586 (N_11586,N_9746,N_5063);
and U11587 (N_11587,N_7901,N_5637);
and U11588 (N_11588,N_7267,N_7733);
and U11589 (N_11589,N_7974,N_5849);
nor U11590 (N_11590,N_9697,N_5951);
nor U11591 (N_11591,N_8125,N_9590);
or U11592 (N_11592,N_8143,N_9586);
and U11593 (N_11593,N_8957,N_6984);
and U11594 (N_11594,N_9000,N_5603);
nor U11595 (N_11595,N_7213,N_8892);
nand U11596 (N_11596,N_9695,N_5258);
xnor U11597 (N_11597,N_7814,N_8528);
or U11598 (N_11598,N_6002,N_6370);
or U11599 (N_11599,N_5553,N_8371);
xor U11600 (N_11600,N_8835,N_9585);
nand U11601 (N_11601,N_8692,N_5069);
nor U11602 (N_11602,N_8785,N_8177);
or U11603 (N_11603,N_8510,N_6487);
or U11604 (N_11604,N_6673,N_5218);
or U11605 (N_11605,N_5765,N_9556);
nand U11606 (N_11606,N_5488,N_6331);
and U11607 (N_11607,N_7992,N_6693);
and U11608 (N_11608,N_7782,N_8336);
or U11609 (N_11609,N_5943,N_7484);
nand U11610 (N_11610,N_5711,N_6730);
xor U11611 (N_11611,N_7304,N_6138);
or U11612 (N_11612,N_8350,N_9278);
nand U11613 (N_11613,N_7999,N_5262);
xor U11614 (N_11614,N_8953,N_8384);
nand U11615 (N_11615,N_7083,N_6855);
or U11616 (N_11616,N_6557,N_7909);
nand U11617 (N_11617,N_5753,N_7130);
nor U11618 (N_11618,N_9421,N_8704);
xor U11619 (N_11619,N_7673,N_5276);
nor U11620 (N_11620,N_9468,N_8193);
nor U11621 (N_11621,N_5419,N_9844);
nand U11622 (N_11622,N_9581,N_9404);
and U11623 (N_11623,N_7444,N_6117);
nand U11624 (N_11624,N_7459,N_9025);
nor U11625 (N_11625,N_9477,N_5870);
nand U11626 (N_11626,N_9006,N_9089);
xor U11627 (N_11627,N_6528,N_6434);
xnor U11628 (N_11628,N_8736,N_6354);
nand U11629 (N_11629,N_6733,N_6583);
nor U11630 (N_11630,N_8467,N_7242);
xor U11631 (N_11631,N_9135,N_6079);
xnor U11632 (N_11632,N_6555,N_6120);
and U11633 (N_11633,N_8035,N_5382);
nor U11634 (N_11634,N_9687,N_8820);
nor U11635 (N_11635,N_5451,N_7255);
or U11636 (N_11636,N_7307,N_7657);
and U11637 (N_11637,N_9368,N_7296);
and U11638 (N_11638,N_8104,N_5295);
or U11639 (N_11639,N_8481,N_8595);
nand U11640 (N_11640,N_8414,N_8308);
xor U11641 (N_11641,N_8955,N_6939);
nor U11642 (N_11642,N_5267,N_8768);
or U11643 (N_11643,N_9012,N_7132);
xnor U11644 (N_11644,N_5833,N_6167);
or U11645 (N_11645,N_9269,N_5763);
nand U11646 (N_11646,N_5947,N_7933);
nor U11647 (N_11647,N_9915,N_9466);
and U11648 (N_11648,N_9744,N_8739);
xnor U11649 (N_11649,N_8877,N_6785);
or U11650 (N_11650,N_5384,N_8825);
or U11651 (N_11651,N_8807,N_8489);
or U11652 (N_11652,N_5039,N_8365);
nor U11653 (N_11653,N_7383,N_8620);
nor U11654 (N_11654,N_6219,N_7869);
nor U11655 (N_11655,N_8725,N_5706);
xor U11656 (N_11656,N_5742,N_9851);
nand U11657 (N_11657,N_8811,N_9016);
xor U11658 (N_11658,N_5170,N_5831);
xnor U11659 (N_11659,N_5911,N_6297);
nand U11660 (N_11660,N_7513,N_9491);
nor U11661 (N_11661,N_6577,N_9142);
xor U11662 (N_11662,N_7200,N_5391);
and U11663 (N_11663,N_9158,N_6486);
xor U11664 (N_11664,N_9863,N_9041);
nand U11665 (N_11665,N_6514,N_8073);
or U11666 (N_11666,N_5042,N_5066);
or U11667 (N_11667,N_7030,N_7039);
or U11668 (N_11668,N_6488,N_5009);
and U11669 (N_11669,N_9820,N_9054);
or U11670 (N_11670,N_6798,N_5261);
and U11671 (N_11671,N_8516,N_9287);
and U11672 (N_11672,N_5232,N_9336);
or U11673 (N_11673,N_5976,N_9798);
and U11674 (N_11674,N_6684,N_8408);
nand U11675 (N_11675,N_6450,N_8934);
xnor U11676 (N_11676,N_7258,N_8413);
or U11677 (N_11677,N_6057,N_5270);
nor U11678 (N_11678,N_6842,N_8285);
nor U11679 (N_11679,N_9290,N_9964);
xnor U11680 (N_11680,N_7543,N_5944);
or U11681 (N_11681,N_9077,N_6304);
nor U11682 (N_11682,N_6947,N_6453);
xnor U11683 (N_11683,N_8961,N_6737);
xnor U11684 (N_11684,N_6539,N_8463);
and U11685 (N_11685,N_6554,N_6000);
nor U11686 (N_11686,N_5978,N_7003);
xor U11687 (N_11687,N_6242,N_6668);
or U11688 (N_11688,N_8089,N_9911);
and U11689 (N_11689,N_6445,N_5202);
nand U11690 (N_11690,N_6676,N_9508);
xor U11691 (N_11691,N_8165,N_7465);
or U11692 (N_11692,N_8822,N_6599);
xnor U11693 (N_11693,N_8228,N_7776);
xnor U11694 (N_11694,N_8688,N_8504);
and U11695 (N_11695,N_7058,N_6627);
nor U11696 (N_11696,N_8157,N_5672);
nand U11697 (N_11697,N_6870,N_6978);
or U11698 (N_11698,N_8592,N_7661);
and U11699 (N_11699,N_8327,N_8438);
or U11700 (N_11700,N_7702,N_5966);
and U11701 (N_11701,N_9132,N_7025);
nand U11702 (N_11702,N_7080,N_7420);
nand U11703 (N_11703,N_5086,N_5678);
and U11704 (N_11704,N_8201,N_9509);
nand U11705 (N_11705,N_9567,N_9381);
and U11706 (N_11706,N_7051,N_6490);
xnor U11707 (N_11707,N_8237,N_6742);
or U11708 (N_11708,N_7602,N_6787);
nor U11709 (N_11709,N_7422,N_5183);
nor U11710 (N_11710,N_9878,N_9110);
xor U11711 (N_11711,N_6011,N_5457);
nor U11712 (N_11712,N_8794,N_5867);
or U11713 (N_11713,N_6051,N_7263);
and U11714 (N_11714,N_7970,N_5185);
xor U11715 (N_11715,N_5986,N_6839);
xor U11716 (N_11716,N_6658,N_9339);
xnor U11717 (N_11717,N_8991,N_5782);
and U11718 (N_11718,N_9068,N_5206);
xor U11719 (N_11719,N_7805,N_5750);
nand U11720 (N_11720,N_5427,N_7850);
nand U11721 (N_11721,N_5702,N_9907);
xnor U11722 (N_11722,N_9872,N_5658);
and U11723 (N_11723,N_8567,N_6931);
and U11724 (N_11724,N_8392,N_5179);
and U11725 (N_11725,N_5471,N_5418);
and U11726 (N_11726,N_7829,N_8446);
xnor U11727 (N_11727,N_5074,N_5627);
nor U11728 (N_11728,N_8071,N_7454);
and U11729 (N_11729,N_7302,N_5331);
and U11730 (N_11730,N_7637,N_5399);
nor U11731 (N_11731,N_7542,N_9545);
nand U11732 (N_11732,N_7646,N_7613);
nor U11733 (N_11733,N_7344,N_6492);
nor U11734 (N_11734,N_6724,N_5367);
nand U11735 (N_11735,N_6898,N_8668);
nor U11736 (N_11736,N_8386,N_6935);
nor U11737 (N_11737,N_7994,N_6054);
nand U11738 (N_11738,N_5223,N_6619);
nor U11739 (N_11739,N_7450,N_6953);
or U11740 (N_11740,N_5574,N_7410);
nor U11741 (N_11741,N_6763,N_9998);
nand U11742 (N_11742,N_6749,N_8259);
nand U11743 (N_11743,N_6612,N_6249);
nand U11744 (N_11744,N_5898,N_8537);
and U11745 (N_11745,N_5330,N_7074);
and U11746 (N_11746,N_9858,N_9662);
xor U11747 (N_11747,N_8097,N_9520);
nor U11748 (N_11748,N_8927,N_5263);
nand U11749 (N_11749,N_5132,N_9083);
and U11750 (N_11750,N_5516,N_6773);
xor U11751 (N_11751,N_6390,N_5777);
and U11752 (N_11752,N_6328,N_7445);
xnor U11753 (N_11753,N_8754,N_8946);
and U11754 (N_11754,N_5942,N_6288);
or U11755 (N_11755,N_9156,N_9322);
and U11756 (N_11756,N_6091,N_7783);
xnor U11757 (N_11757,N_7533,N_8172);
nand U11758 (N_11758,N_5222,N_7195);
nor U11759 (N_11759,N_6734,N_6049);
or U11760 (N_11760,N_7727,N_5640);
nor U11761 (N_11761,N_7095,N_9352);
nor U11762 (N_11762,N_7019,N_6615);
and U11763 (N_11763,N_7233,N_8487);
xnor U11764 (N_11764,N_7217,N_7914);
and U11765 (N_11765,N_7738,N_5800);
nor U11766 (N_11766,N_9980,N_5827);
nand U11767 (N_11767,N_6351,N_5021);
xor U11768 (N_11768,N_6083,N_7791);
and U11769 (N_11769,N_8675,N_8138);
nor U11770 (N_11770,N_8119,N_7645);
xor U11771 (N_11771,N_9106,N_7362);
nor U11772 (N_11772,N_6084,N_7892);
and U11773 (N_11773,N_5329,N_6620);
or U11774 (N_11774,N_8639,N_9107);
xnor U11775 (N_11775,N_8547,N_5017);
nand U11776 (N_11776,N_6533,N_7977);
or U11777 (N_11777,N_8063,N_7957);
nand U11778 (N_11778,N_6341,N_9036);
or U11779 (N_11779,N_8329,N_5401);
and U11780 (N_11780,N_6893,N_6897);
and U11781 (N_11781,N_7480,N_9251);
xnor U11782 (N_11782,N_8405,N_5894);
nand U11783 (N_11783,N_6243,N_5554);
and U11784 (N_11784,N_6657,N_8544);
or U11785 (N_11785,N_7034,N_8373);
nor U11786 (N_11786,N_6756,N_5551);
or U11787 (N_11787,N_9056,N_9924);
xor U11788 (N_11788,N_6802,N_7151);
nor U11789 (N_11789,N_7761,N_6746);
nor U11790 (N_11790,N_6491,N_5316);
or U11791 (N_11791,N_8753,N_5647);
and U11792 (N_11792,N_6607,N_5644);
nand U11793 (N_11793,N_8858,N_8895);
nor U11794 (N_11794,N_9248,N_5075);
xor U11795 (N_11795,N_8578,N_5503);
and U11796 (N_11796,N_7158,N_6186);
and U11797 (N_11797,N_5600,N_6685);
xor U11798 (N_11798,N_8306,N_7338);
xnor U11799 (N_11799,N_6818,N_5893);
or U11800 (N_11800,N_5173,N_5839);
and U11801 (N_11801,N_7462,N_7376);
nand U11802 (N_11802,N_6726,N_7907);
nor U11803 (N_11803,N_6179,N_9663);
nor U11804 (N_11804,N_6604,N_9741);
nand U11805 (N_11805,N_9332,N_6359);
nand U11806 (N_11806,N_6654,N_5991);
nand U11807 (N_11807,N_7396,N_7765);
nor U11808 (N_11808,N_6237,N_5498);
and U11809 (N_11809,N_6290,N_6193);
xor U11810 (N_11810,N_8783,N_7799);
nor U11811 (N_11811,N_8250,N_8344);
and U11812 (N_11812,N_7807,N_8646);
nor U11813 (N_11813,N_8601,N_9785);
or U11814 (N_11814,N_9728,N_6285);
or U11815 (N_11815,N_8075,N_7423);
xor U11816 (N_11816,N_8088,N_6067);
nor U11817 (N_11817,N_8086,N_7451);
or U11818 (N_11818,N_6190,N_9464);
and U11819 (N_11819,N_5077,N_8800);
and U11820 (N_11820,N_6272,N_6127);
nand U11821 (N_11821,N_7254,N_5741);
and U11822 (N_11822,N_8676,N_8345);
nand U11823 (N_11823,N_8916,N_5590);
nand U11824 (N_11824,N_7865,N_8778);
xor U11825 (N_11825,N_7671,N_9816);
xor U11826 (N_11826,N_8717,N_9574);
xor U11827 (N_11827,N_7225,N_5153);
and U11828 (N_11828,N_9837,N_5830);
and U11829 (N_11829,N_8756,N_6369);
nand U11830 (N_11830,N_7485,N_9361);
xor U11831 (N_11831,N_6560,N_6621);
or U11832 (N_11832,N_6398,N_8641);
or U11833 (N_11833,N_9124,N_6882);
nor U11834 (N_11834,N_7695,N_9441);
nand U11835 (N_11835,N_5948,N_9384);
nor U11836 (N_11836,N_9646,N_6872);
or U11837 (N_11837,N_5961,N_8784);
nor U11838 (N_11838,N_8969,N_9722);
xnor U11839 (N_11839,N_9096,N_7066);
nor U11840 (N_11840,N_5685,N_8362);
nor U11841 (N_11841,N_6114,N_8548);
nand U11842 (N_11842,N_5256,N_7027);
xnor U11843 (N_11843,N_9241,N_9203);
nor U11844 (N_11844,N_6317,N_6116);
or U11845 (N_11845,N_6962,N_5119);
or U11846 (N_11846,N_8156,N_8275);
nor U11847 (N_11847,N_7222,N_8380);
nor U11848 (N_11848,N_5852,N_5409);
and U11849 (N_11849,N_5084,N_6824);
or U11850 (N_11850,N_6853,N_5705);
nor U11851 (N_11851,N_5691,N_6494);
nand U11852 (N_11852,N_5062,N_5114);
xnor U11853 (N_11853,N_8391,N_9914);
and U11854 (N_11854,N_7951,N_5605);
nor U11855 (N_11855,N_7118,N_6813);
xnor U11856 (N_11856,N_5129,N_6108);
nand U11857 (N_11857,N_8755,N_7679);
nand U11858 (N_11858,N_6052,N_9518);
xnor U11859 (N_11859,N_9681,N_9927);
nand U11860 (N_11860,N_7529,N_8162);
nor U11861 (N_11861,N_9876,N_8442);
nand U11862 (N_11862,N_9838,N_8559);
xor U11863 (N_11863,N_7137,N_6367);
nor U11864 (N_11864,N_9689,N_5786);
and U11865 (N_11865,N_9896,N_7762);
nor U11866 (N_11866,N_6053,N_7526);
nor U11867 (N_11867,N_7332,N_8437);
or U11868 (N_11868,N_5283,N_8432);
nor U11869 (N_11869,N_9535,N_8653);
or U11870 (N_11870,N_9257,N_8159);
nand U11871 (N_11871,N_8468,N_8861);
nor U11872 (N_11872,N_6760,N_6227);
and U11873 (N_11873,N_9919,N_8115);
or U11874 (N_11874,N_7275,N_8401);
and U11875 (N_11875,N_5307,N_8596);
or U11876 (N_11876,N_6542,N_6944);
or U11877 (N_11877,N_7600,N_8939);
nand U11878 (N_11878,N_5739,N_6211);
xnor U11879 (N_11879,N_7708,N_7050);
nor U11880 (N_11880,N_5272,N_5687);
nor U11881 (N_11881,N_9364,N_6291);
xor U11882 (N_11882,N_7098,N_7972);
and U11883 (N_11883,N_7402,N_7565);
nor U11884 (N_11884,N_8366,N_8950);
nand U11885 (N_11885,N_6988,N_5378);
nand U11886 (N_11886,N_8512,N_8374);
or U11887 (N_11887,N_5648,N_8270);
xnor U11888 (N_11888,N_9794,N_8777);
xor U11889 (N_11889,N_6498,N_7412);
nor U11890 (N_11890,N_9424,N_6951);
or U11891 (N_11891,N_8937,N_6903);
nor U11892 (N_11892,N_7898,N_6509);
or U11893 (N_11893,N_7984,N_9460);
nand U11894 (N_11894,N_5155,N_5024);
xnor U11895 (N_11895,N_7125,N_6152);
xnor U11896 (N_11896,N_6761,N_6275);
xnor U11897 (N_11897,N_7183,N_8118);
or U11898 (N_11898,N_8944,N_8959);
xor U11899 (N_11899,N_5883,N_6500);
xor U11900 (N_11900,N_7585,N_6948);
and U11901 (N_11901,N_6081,N_5802);
xor U11902 (N_11902,N_9017,N_8135);
nor U11903 (N_11903,N_9946,N_7122);
and U11904 (N_11904,N_6709,N_5174);
or U11905 (N_11905,N_9162,N_9698);
and U11906 (N_11906,N_6905,N_6579);
and U11907 (N_11907,N_9015,N_9453);
nor U11908 (N_11908,N_8037,N_9356);
nor U11909 (N_11909,N_7960,N_9724);
nor U11910 (N_11910,N_9920,N_8342);
or U11911 (N_11911,N_8663,N_6222);
nand U11912 (N_11912,N_6478,N_7032);
xor U11913 (N_11913,N_8080,N_9280);
nand U11914 (N_11914,N_7819,N_5993);
nor U11915 (N_11915,N_7873,N_8729);
nand U11916 (N_11916,N_6068,N_8792);
nor U11917 (N_11917,N_9493,N_7072);
and U11918 (N_11918,N_7024,N_5842);
nor U11919 (N_11919,N_9401,N_7855);
or U11920 (N_11920,N_5916,N_7433);
or U11921 (N_11921,N_6664,N_9071);
nor U11922 (N_11922,N_6712,N_9255);
and U11923 (N_11923,N_6970,N_9640);
and U11924 (N_11924,N_8146,N_6404);
xnor U11925 (N_11925,N_8826,N_9577);
xnor U11926 (N_11926,N_6303,N_7630);
or U11927 (N_11927,N_7119,N_7811);
xor U11928 (N_11928,N_6553,N_8187);
or U11929 (N_11929,N_5458,N_5364);
xor U11930 (N_11930,N_5064,N_6963);
nor U11931 (N_11931,N_8840,N_5552);
or U11932 (N_11932,N_6831,N_5555);
or U11933 (N_11933,N_7785,N_8869);
xor U11934 (N_11934,N_9818,N_7078);
or U11935 (N_11935,N_5030,N_5046);
or U11936 (N_11936,N_5592,N_8357);
nand U11937 (N_11937,N_9988,N_6517);
nor U11938 (N_11938,N_8012,N_5342);
nor U11939 (N_11939,N_9786,N_7575);
nand U11940 (N_11940,N_8821,N_6260);
xnor U11941 (N_11941,N_6906,N_7768);
and U11942 (N_11942,N_5477,N_7317);
or U11943 (N_11943,N_9993,N_7847);
and U11944 (N_11944,N_7463,N_7416);
nor U11945 (N_11945,N_6449,N_7228);
nand U11946 (N_11946,N_8726,N_8292);
xnor U11947 (N_11947,N_9898,N_8915);
xor U11948 (N_11948,N_9793,N_9176);
nor U11949 (N_11949,N_5395,N_8968);
xor U11950 (N_11950,N_9671,N_8488);
xor U11951 (N_11951,N_6311,N_6739);
xnor U11952 (N_11952,N_7005,N_7469);
or U11953 (N_11953,N_7367,N_9561);
or U11954 (N_11954,N_5805,N_5807);
xnor U11955 (N_11955,N_9713,N_8001);
xnor U11956 (N_11956,N_9522,N_7777);
nand U11957 (N_11957,N_7173,N_5980);
or U11958 (N_11958,N_5048,N_8296);
nand U11959 (N_11959,N_5105,N_7822);
nor U11960 (N_11960,N_6986,N_9070);
nand U11961 (N_11961,N_5038,N_8672);
xnor U11962 (N_11962,N_8847,N_9134);
and U11963 (N_11963,N_9835,N_6332);
xnor U11964 (N_11964,N_9144,N_6216);
xor U11965 (N_11965,N_5566,N_8659);
or U11966 (N_11966,N_9351,N_5152);
xor U11967 (N_11967,N_7112,N_9253);
xor U11968 (N_11968,N_8435,N_7710);
or U11969 (N_11969,N_7261,N_6365);
or U11970 (N_11970,N_5357,N_6321);
and U11971 (N_11971,N_5708,N_7592);
or U11972 (N_11972,N_9313,N_8889);
or U11973 (N_11973,N_5809,N_5912);
xnor U11974 (N_11974,N_8931,N_9745);
or U11975 (N_11975,N_5609,N_8207);
nor U11976 (N_11976,N_6158,N_7298);
and U11977 (N_11977,N_9275,N_9918);
xor U11978 (N_11978,N_5576,N_9263);
nor U11979 (N_11979,N_8341,N_8100);
and U11980 (N_11980,N_9288,N_8267);
and U11981 (N_11981,N_5548,N_7965);
and U11982 (N_11982,N_8377,N_5547);
xor U11983 (N_11983,N_8494,N_8574);
nor U11984 (N_11984,N_5535,N_6214);
nand U11985 (N_11985,N_6653,N_6467);
and U11986 (N_11986,N_6825,N_9688);
xor U11987 (N_11987,N_7882,N_8497);
or U11988 (N_11988,N_8527,N_7215);
nor U11989 (N_11989,N_5734,N_7745);
or U11990 (N_11990,N_9558,N_7363);
nor U11991 (N_11991,N_9726,N_9826);
or U11992 (N_11992,N_9103,N_6926);
nor U11993 (N_11993,N_5247,N_6830);
xor U11994 (N_11994,N_6153,N_8870);
or U11995 (N_11995,N_5604,N_7124);
and U11996 (N_11996,N_5714,N_7163);
and U11997 (N_11997,N_6800,N_5885);
xnor U11998 (N_11998,N_5970,N_9111);
and U11999 (N_11999,N_8262,N_7185);
nand U12000 (N_12000,N_7328,N_8042);
and U12001 (N_12001,N_9670,N_7278);
nand U12002 (N_12002,N_7467,N_8642);
nand U12003 (N_12003,N_9892,N_8354);
nor U12004 (N_12004,N_8552,N_5466);
nand U12005 (N_12005,N_8122,N_8841);
or U12006 (N_12006,N_5082,N_9147);
nand U12007 (N_12007,N_5529,N_5923);
nor U12008 (N_12008,N_9344,N_6322);
and U12009 (N_12009,N_5797,N_8809);
and U12010 (N_12010,N_7084,N_5612);
and U12011 (N_12011,N_9377,N_7086);
nand U12012 (N_12012,N_7934,N_7250);
xor U12013 (N_12013,N_7771,N_9756);
xnor U12014 (N_12014,N_9650,N_9228);
or U12015 (N_12015,N_6752,N_9797);
nor U12016 (N_12016,N_7369,N_5379);
and U12017 (N_12017,N_7097,N_5334);
nor U12018 (N_12018,N_8190,N_5396);
nand U12019 (N_12019,N_7894,N_5861);
nor U12020 (N_12020,N_6797,N_7021);
xnor U12021 (N_12021,N_9309,N_9540);
and U12022 (N_12022,N_6662,N_5167);
or U12023 (N_12023,N_6236,N_5514);
or U12024 (N_12024,N_5440,N_8024);
nand U12025 (N_12025,N_8221,N_5217);
and U12026 (N_12026,N_6274,N_6907);
or U12027 (N_12027,N_8418,N_8302);
or U12028 (N_12028,N_6765,N_7189);
nor U12029 (N_12029,N_6534,N_6974);
and U12030 (N_12030,N_5764,N_5776);
or U12031 (N_12031,N_7723,N_8041);
or U12032 (N_12032,N_8206,N_9985);
and U12033 (N_12033,N_6197,N_9822);
nand U12034 (N_12034,N_7094,N_5686);
or U12035 (N_12035,N_6810,N_7562);
xnor U12036 (N_12036,N_5789,N_9494);
and U12037 (N_12037,N_7160,N_8111);
xor U12038 (N_12038,N_7041,N_6391);
xnor U12039 (N_12039,N_8656,N_5106);
or U12040 (N_12040,N_9500,N_7274);
nor U12041 (N_12041,N_8404,N_9127);
and U12042 (N_12042,N_6017,N_5197);
nand U12043 (N_12043,N_9917,N_5982);
nand U12044 (N_12044,N_9737,N_6071);
nand U12045 (N_12045,N_6928,N_5434);
nor U12046 (N_12046,N_8376,N_8926);
or U12047 (N_12047,N_9937,N_9767);
and U12048 (N_12048,N_5636,N_5462);
and U12049 (N_12049,N_7110,N_6545);
nand U12050 (N_12050,N_7231,N_9271);
nand U12051 (N_12051,N_5549,N_6335);
or U12052 (N_12052,N_9609,N_5524);
xor U12053 (N_12053,N_8178,N_9612);
xnor U12054 (N_12054,N_7763,N_5820);
nand U12055 (N_12055,N_6869,N_7684);
nand U12056 (N_12056,N_7590,N_6776);
nor U12057 (N_12057,N_9781,N_7870);
or U12058 (N_12058,N_5456,N_5355);
and U12059 (N_12059,N_7436,N_5041);
or U12060 (N_12060,N_6030,N_9888);
nor U12061 (N_12061,N_5874,N_5879);
nor U12062 (N_12062,N_8124,N_9966);
or U12063 (N_12063,N_5737,N_8977);
nor U12064 (N_12064,N_9069,N_9359);
xor U12065 (N_12065,N_8815,N_7535);
and U12066 (N_12066,N_8767,N_5722);
xnor U12067 (N_12067,N_8265,N_5973);
and U12068 (N_12068,N_6766,N_5241);
nand U12069 (N_12069,N_5619,N_9855);
and U12070 (N_12070,N_9184,N_9448);
and U12071 (N_12071,N_8763,N_8684);
or U12072 (N_12072,N_7609,N_5938);
and U12073 (N_12073,N_8648,N_7188);
xnor U12074 (N_12074,N_8936,N_7131);
xnor U12075 (N_12075,N_9328,N_7029);
nor U12076 (N_12076,N_9150,N_6934);
nor U12077 (N_12077,N_5054,N_6858);
or U12078 (N_12078,N_5960,N_8849);
or U12079 (N_12079,N_5723,N_9994);
xor U12080 (N_12080,N_7778,N_9665);
xnor U12081 (N_12081,N_9406,N_7887);
xnor U12082 (N_12082,N_9218,N_8913);
and U12083 (N_12083,N_8897,N_6562);
nor U12084 (N_12084,N_6601,N_8918);
nand U12085 (N_12085,N_7497,N_5507);
xor U12086 (N_12086,N_7342,N_5389);
xor U12087 (N_12087,N_9051,N_9542);
and U12088 (N_12088,N_9813,N_9002);
nor U12089 (N_12089,N_6608,N_6395);
or U12090 (N_12090,N_8057,N_8307);
or U12091 (N_12091,N_6026,N_9409);
nand U12092 (N_12092,N_5550,N_5352);
and U12093 (N_12093,N_7059,N_7636);
xnor U12094 (N_12094,N_5724,N_9532);
nor U12095 (N_12095,N_8332,N_6185);
nand U12096 (N_12096,N_5305,N_5926);
or U12097 (N_12097,N_7208,N_8633);
or U12098 (N_12098,N_8699,N_7647);
or U12099 (N_12099,N_7096,N_8963);
or U12100 (N_12100,N_6559,N_8586);
and U12101 (N_12101,N_7478,N_7260);
xnor U12102 (N_12102,N_5608,N_9510);
xor U12103 (N_12103,N_7431,N_8893);
or U12104 (N_12104,N_9771,N_5230);
nand U12105 (N_12105,N_7913,N_6902);
xnor U12106 (N_12106,N_9992,N_5914);
or U12107 (N_12107,N_6229,N_5214);
xnor U12108 (N_12108,N_7073,N_5260);
nand U12109 (N_12109,N_9841,N_7884);
nand U12110 (N_12110,N_5508,N_7108);
nor U12111 (N_12111,N_5749,N_9484);
and U12112 (N_12112,N_6228,N_5844);
xnor U12113 (N_12113,N_5485,N_7987);
nor U12114 (N_12114,N_6632,N_6659);
or U12115 (N_12115,N_8483,N_5271);
or U12116 (N_12116,N_9642,N_6605);
nor U12117 (N_12117,N_8383,N_9408);
nor U12118 (N_12118,N_7519,N_7448);
xor U12119 (N_12119,N_6314,N_9667);
xnor U12120 (N_12120,N_8191,N_6221);
nand U12121 (N_12121,N_9065,N_6283);
or U12122 (N_12122,N_8762,N_8735);
and U12123 (N_12123,N_8819,N_9559);
and U12124 (N_12124,N_7803,N_8116);
xor U12125 (N_12125,N_7766,N_9572);
nor U12126 (N_12126,N_7844,N_8347);
and U12127 (N_12127,N_9541,N_5365);
or U12128 (N_12128,N_7764,N_6790);
or U12129 (N_12129,N_8622,N_9242);
nand U12130 (N_12130,N_7297,N_9897);
nor U12131 (N_12131,N_6769,N_8508);
nor U12132 (N_12132,N_9062,N_5412);
or U12133 (N_12133,N_9999,N_7866);
xor U12134 (N_12134,N_8520,N_6877);
or U12135 (N_12135,N_7435,N_5934);
nand U12136 (N_12136,N_5787,N_9227);
xnor U12137 (N_12137,N_6161,N_8242);
and U12138 (N_12138,N_7834,N_7554);
and U12139 (N_12139,N_5902,N_5186);
nand U12140 (N_12140,N_5140,N_9766);
or U12141 (N_12141,N_8741,N_8211);
or U12142 (N_12142,N_7953,N_8101);
xor U12143 (N_12143,N_7503,N_8016);
or U12144 (N_12144,N_7881,N_8022);
and U12145 (N_12145,N_9748,N_8984);
or U12146 (N_12146,N_6137,N_8379);
nor U12147 (N_12147,N_7305,N_7391);
and U12148 (N_12148,N_9755,N_9891);
nand U12149 (N_12149,N_6613,N_8846);
or U12150 (N_12150,N_9801,N_9930);
and U12151 (N_12151,N_7218,N_6881);
nor U12152 (N_12152,N_6422,N_7486);
xor U12153 (N_12153,N_6814,N_9386);
and U12154 (N_12154,N_9716,N_8070);
nor U12155 (N_12155,N_8982,N_9571);
nor U12156 (N_12156,N_5242,N_7925);
xnor U12157 (N_12157,N_5613,N_7295);
nand U12158 (N_12158,N_7081,N_8003);
and U12159 (N_12159,N_6999,N_8402);
or U12160 (N_12160,N_7964,N_5684);
and U12161 (N_12161,N_5216,N_9395);
and U12162 (N_12162,N_9815,N_9367);
and U12163 (N_12163,N_9624,N_7427);
nand U12164 (N_12164,N_6165,N_8026);
or U12165 (N_12165,N_8174,N_7747);
and U12166 (N_12166,N_7986,N_5866);
xnor U12167 (N_12167,N_6131,N_5918);
or U12168 (N_12168,N_8536,N_6059);
nand U12169 (N_12169,N_8938,N_7282);
nand U12170 (N_12170,N_9091,N_6884);
xor U12171 (N_12171,N_7638,N_9337);
or U12172 (N_12172,N_8011,N_8747);
and U12173 (N_12173,N_8857,N_9282);
nor U12174 (N_12174,N_5117,N_5847);
or U12175 (N_12175,N_7205,N_9703);
xor U12176 (N_12176,N_7696,N_6100);
or U12177 (N_12177,N_5237,N_7341);
xnor U12178 (N_12178,N_6535,N_8180);
xnor U12179 (N_12179,N_8030,N_5843);
nand U12180 (N_12180,N_9034,N_8625);
nand U12181 (N_12181,N_6308,N_7948);
xor U12182 (N_12182,N_7606,N_5792);
and U12183 (N_12183,N_7985,N_7998);
and U12184 (N_12184,N_9963,N_6708);
or U12185 (N_12185,N_6039,N_7294);
nand U12186 (N_12186,N_6983,N_8355);
nand U12187 (N_12187,N_9730,N_7310);
xnor U12188 (N_12188,N_7316,N_8630);
nand U12189 (N_12189,N_5872,N_8456);
nand U12190 (N_12190,N_6624,N_5804);
or U12191 (N_12191,N_9700,N_6250);
nand U12192 (N_12192,N_8606,N_9125);
or U12193 (N_12193,N_7234,N_7235);
nor U12194 (N_12194,N_7251,N_7458);
nand U12195 (N_12195,N_9210,N_5110);
or U12196 (N_12196,N_7760,N_6380);
xnor U12197 (N_12197,N_9321,N_7065);
or U12198 (N_12198,N_6564,N_5720);
xnor U12199 (N_12199,N_6270,N_5482);
and U12200 (N_12200,N_7876,N_8087);
nor U12201 (N_12201,N_9589,N_5718);
or U12202 (N_12202,N_5229,N_5338);
nor U12203 (N_12203,N_7941,N_9965);
nand U12204 (N_12204,N_9350,N_7635);
xor U12205 (N_12205,N_7139,N_9402);
nor U12206 (N_12206,N_8799,N_5193);
and U12207 (N_12207,N_7962,N_6095);
or U12208 (N_12208,N_5348,N_5585);
nand U12209 (N_12209,N_8604,N_6671);
xnor U12210 (N_12210,N_9672,N_5994);
nor U12211 (N_12211,N_7633,N_5225);
nand U12212 (N_12212,N_8990,N_5151);
xor U12213 (N_12213,N_6295,N_6705);
or U12214 (N_12214,N_7879,N_8942);
nor U12215 (N_12215,N_5582,N_9639);
or U12216 (N_12216,N_6967,N_8833);
or U12217 (N_12217,N_7949,N_6265);
nand U12218 (N_12218,N_8369,N_8136);
nand U12219 (N_12219,N_9128,N_7500);
nand U12220 (N_12220,N_6965,N_8367);
xor U12221 (N_12221,N_9382,N_9596);
and U12222 (N_12222,N_5341,N_8560);
or U12223 (N_12223,N_9684,N_9823);
nand U12224 (N_12224,N_7133,N_6715);
nor U12225 (N_12225,N_9506,N_5715);
or U12226 (N_12226,N_6895,N_6678);
nand U12227 (N_12227,N_9209,N_8579);
or U12228 (N_12228,N_9579,N_5569);
or U12229 (N_12229,N_7534,N_7973);
and U12230 (N_12230,N_9192,N_6975);
and U12231 (N_12231,N_9583,N_7596);
xor U12232 (N_12232,N_8752,N_8085);
nor U12233 (N_12233,N_7821,N_8368);
and U12234 (N_12234,N_6246,N_9229);
and U12235 (N_12235,N_8891,N_6421);
nor U12236 (N_12236,N_5055,N_6989);
xnor U12237 (N_12237,N_8714,N_7788);
nor U12238 (N_12238,N_9882,N_8524);
and U12239 (N_12239,N_6040,N_8576);
nor U12240 (N_12240,N_5354,N_9240);
xnor U12241 (N_12241,N_6524,N_5560);
xnor U12242 (N_12242,N_7918,N_5523);
nand U12243 (N_12243,N_6861,N_7227);
nand U12244 (N_12244,N_5464,N_6473);
and U12245 (N_12245,N_5481,N_6714);
nand U12246 (N_12246,N_7240,N_8581);
and U12247 (N_12247,N_6082,N_5245);
and U12248 (N_12248,N_8431,N_6846);
nor U12249 (N_12249,N_9782,N_5073);
or U12250 (N_12250,N_8555,N_8751);
nand U12251 (N_12251,N_8612,N_8773);
nor U12252 (N_12252,N_9856,N_6915);
and U12253 (N_12253,N_5076,N_5147);
nand U12254 (N_12254,N_8824,N_9379);
xnor U12255 (N_12255,N_6244,N_5059);
nand U12256 (N_12256,N_9853,N_7057);
nor U12257 (N_12257,N_9115,N_8077);
and U12258 (N_12258,N_9308,N_6993);
nor U12259 (N_12259,N_7404,N_7521);
and U12260 (N_12260,N_7511,N_8852);
xor U12261 (N_12261,N_7839,N_9393);
and U12262 (N_12262,N_7403,N_5142);
nand U12263 (N_12263,N_6927,N_5387);
nand U12264 (N_12264,N_6647,N_9938);
nor U12265 (N_12265,N_8424,N_8903);
nor U12266 (N_12266,N_8664,N_5057);
nor U12267 (N_12267,N_7224,N_6007);
or U12268 (N_12268,N_5937,N_6125);
and U12269 (N_12269,N_7863,N_5735);
nor U12270 (N_12270,N_9587,N_6584);
nand U12271 (N_12271,N_5085,N_6725);
nor U12272 (N_12272,N_6826,N_6111);
or U12273 (N_12273,N_7572,N_9249);
or U12274 (N_12274,N_6472,N_8226);
and U12275 (N_12275,N_7937,N_8233);
or U12276 (N_12276,N_6033,N_5169);
xor U12277 (N_12277,N_6284,N_8151);
nand U12278 (N_12278,N_5007,N_6403);
xor U12279 (N_12279,N_8665,N_9185);
xor U12280 (N_12280,N_6812,N_8492);
xor U12281 (N_12281,N_6996,N_5065);
nand U12282 (N_12282,N_7979,N_7742);
nand U12283 (N_12283,N_5018,N_9706);
or U12284 (N_12284,N_9735,N_5696);
nand U12285 (N_12285,N_5280,N_6669);
and U12286 (N_12286,N_8619,N_5910);
and U12287 (N_12287,N_9824,N_9549);
and U12288 (N_12288,N_8788,N_6200);
xor U12289 (N_12289,N_5783,N_7049);
and U12290 (N_12290,N_6835,N_5090);
or U12291 (N_12291,N_6857,N_5666);
nor U12292 (N_12292,N_5014,N_9563);
or U12293 (N_12293,N_5512,N_5285);
nor U12294 (N_12294,N_9094,N_6854);
and U12295 (N_12295,N_7236,N_5300);
nor U12296 (N_12296,N_8479,N_7581);
nor U12297 (N_12297,N_8240,N_7358);
nor U12298 (N_12298,N_6360,N_9849);
xor U12299 (N_12299,N_7547,N_7891);
nor U12300 (N_12300,N_9869,N_7615);
or U12301 (N_12301,N_7997,N_7910);
or U12302 (N_12302,N_8503,N_9293);
nand U12303 (N_12303,N_9712,N_7128);
nor U12304 (N_12304,N_6240,N_9661);
and U12305 (N_12305,N_5388,N_8107);
nand U12306 (N_12306,N_5780,N_8339);
nor U12307 (N_12307,N_6912,N_5189);
or U12308 (N_12308,N_8871,N_8958);
xnor U12309 (N_12309,N_6419,N_7903);
or U12310 (N_12310,N_5168,N_5244);
nand U12311 (N_12311,N_8040,N_6917);
or U12312 (N_12312,N_7426,N_9747);
nor U12313 (N_12313,N_6635,N_9088);
nand U12314 (N_12314,N_5538,N_9555);
or U12315 (N_12315,N_5450,N_7202);
and U12316 (N_12316,N_9696,N_8687);
or U12317 (N_12317,N_6589,N_6406);
nor U12318 (N_12318,N_5779,N_5108);
xor U12319 (N_12319,N_7515,N_8449);
xor U12320 (N_12320,N_7787,N_5815);
and U12321 (N_12321,N_9895,N_8182);
and U12322 (N_12322,N_6916,N_5534);
or U12323 (N_12323,N_7176,N_7682);
nor U12324 (N_12324,N_9810,N_6064);
nor U12325 (N_12325,N_6339,N_6164);
xor U12326 (N_12326,N_8949,N_5175);
or U12327 (N_12327,N_5744,N_6918);
xnor U12328 (N_12328,N_7502,N_9457);
or U12329 (N_12329,N_9940,N_5213);
or U12330 (N_12330,N_8781,N_6851);
xnor U12331 (N_12331,N_8832,N_5620);
nor U12332 (N_12332,N_7196,N_8795);
or U12333 (N_12333,N_8859,N_6233);
xor U12334 (N_12334,N_6224,N_9340);
nand U12335 (N_12335,N_8301,N_7053);
xor U12336 (N_12336,N_7730,N_7461);
nor U12337 (N_12337,N_8460,N_7257);
nor U12338 (N_12338,N_8149,N_6469);
or U12339 (N_12339,N_6683,N_8608);
xnor U12340 (N_12340,N_7162,N_7028);
or U12341 (N_12341,N_8043,N_9528);
or U12342 (N_12342,N_5895,N_6985);
and U12343 (N_12343,N_5359,N_8277);
xnor U12344 (N_12344,N_8816,N_8546);
xnor U12345 (N_12345,N_5840,N_9487);
nand U12346 (N_12346,N_5595,N_9527);
nand U12347 (N_12347,N_6698,N_5195);
nand U12348 (N_12348,N_8837,N_6191);
xnor U12349 (N_12349,N_5646,N_6833);
nor U12350 (N_12350,N_9292,N_9804);
nor U12351 (N_12351,N_6484,N_8572);
xor U12352 (N_12352,N_9591,N_7731);
or U12353 (N_12353,N_9231,N_6827);
nor U12354 (N_12354,N_6891,N_5121);
nand U12355 (N_12355,N_9725,N_7492);
nand U12356 (N_12356,N_9791,N_6443);
and U12357 (N_12357,N_6710,N_7692);
and U12358 (N_12358,N_8474,N_5034);
or U12359 (N_12359,N_9155,N_7849);
nor U12360 (N_12360,N_6508,N_7197);
nor U12361 (N_12361,N_7871,N_6239);
or U12362 (N_12362,N_7921,N_9010);
and U12363 (N_12363,N_8258,N_6218);
and U12364 (N_12364,N_6160,N_7306);
and U12365 (N_12365,N_7473,N_9277);
or U12366 (N_12366,N_6235,N_5881);
or U12367 (N_12367,N_7000,N_6074);
nor U12368 (N_12368,N_8654,N_8603);
and U12369 (N_12369,N_9945,N_7553);
or U12370 (N_12370,N_6713,N_9605);
xnor U12371 (N_12371,N_8866,N_7944);
xnor U12372 (N_12372,N_8427,N_7544);
xor U12373 (N_12373,N_9245,N_7090);
nor U12374 (N_12374,N_8640,N_5863);
nand U12375 (N_12375,N_7064,N_5577);
or U12376 (N_12376,N_9167,N_8288);
and U12377 (N_12377,N_5103,N_7104);
or U12378 (N_12378,N_5226,N_8899);
xor U12379 (N_12379,N_6378,N_7146);
nor U12380 (N_12380,N_8750,N_6300);
or U12381 (N_12381,N_5601,N_7790);
and U12382 (N_12382,N_7211,N_6255);
nor U12383 (N_12383,N_9149,N_9950);
and U12384 (N_12384,N_8105,N_8598);
nand U12385 (N_12385,N_9428,N_6719);
and U12386 (N_12386,N_7087,N_5291);
or U12387 (N_12387,N_8499,N_6573);
or U12388 (N_12388,N_7853,N_5527);
nand U12389 (N_12389,N_5563,N_5301);
and U12390 (N_12390,N_6136,N_7031);
or U12391 (N_12391,N_8523,N_8691);
and U12392 (N_12392,N_8127,N_5897);
nor U12393 (N_12393,N_5835,N_8197);
xor U12394 (N_12394,N_9143,N_8426);
xnor U12395 (N_12395,N_9314,N_9396);
nor U12396 (N_12396,N_6850,N_9694);
xor U12397 (N_12397,N_7936,N_6860);
xor U12398 (N_12398,N_8830,N_5003);
or U12399 (N_12399,N_5010,N_8666);
nor U12400 (N_12400,N_5159,N_8309);
or U12401 (N_12401,N_9536,N_8453);
xnor U12402 (N_12402,N_7518,N_7508);
or U12403 (N_12403,N_6718,N_6782);
nand U12404 (N_12404,N_5709,N_5350);
or U12405 (N_12405,N_6080,N_8943);
or U12406 (N_12406,N_5679,N_9828);
or U12407 (N_12407,N_9552,N_6336);
or U12408 (N_12408,N_7299,N_7648);
and U12409 (N_12409,N_8607,N_6859);
and U12410 (N_12410,N_5269,N_5876);
and U12411 (N_12411,N_7897,N_6148);
or U12412 (N_12412,N_6791,N_8564);
xnor U12413 (N_12413,N_7357,N_5311);
or U12414 (N_12414,N_8727,N_9594);
nor U12415 (N_12415,N_5738,N_7100);
nor U12416 (N_12416,N_9486,N_9375);
and U12417 (N_12417,N_5322,N_8882);
xnor U12418 (N_12418,N_9311,N_5583);
xnor U12419 (N_12419,N_8652,N_6976);
and U12420 (N_12420,N_5016,N_9617);
xor U12421 (N_12421,N_6571,N_9442);
nand U12422 (N_12422,N_5390,N_6230);
or U12423 (N_12423,N_6786,N_6475);
nor U12424 (N_12424,N_8519,N_5845);
nand U12425 (N_12425,N_5351,N_7109);
or U12426 (N_12426,N_6552,N_9334);
xnor U12427 (N_12427,N_6502,N_6383);
xor U12428 (N_12428,N_8787,N_9481);
nor U12429 (N_12429,N_6109,N_5163);
nand U12430 (N_12430,N_9262,N_8817);
xor U12431 (N_12431,N_5826,N_5279);
and U12432 (N_12432,N_5015,N_9480);
nor U12433 (N_12433,N_5487,N_8252);
nand U12434 (N_12434,N_9762,N_6527);
and U12435 (N_12435,N_7946,N_5281);
or U12436 (N_12436,N_7008,N_7981);
and U12437 (N_12437,N_5977,N_5008);
nor U12438 (N_12438,N_5332,N_9458);
xor U12439 (N_12439,N_5025,N_9602);
or U12440 (N_12440,N_8430,N_5887);
nor U12441 (N_12441,N_7022,N_5045);
xnor U12442 (N_12442,N_9274,N_9177);
xnor U12443 (N_12443,N_7355,N_7482);
nand U12444 (N_12444,N_5935,N_6409);
nand U12445 (N_12445,N_6154,N_6182);
or U12446 (N_12446,N_6086,N_5124);
or U12447 (N_12447,N_7327,N_8716);
and U12448 (N_12448,N_9543,N_9399);
and U12449 (N_12449,N_7538,N_5614);
and U12450 (N_12450,N_7079,N_6731);
nor U12451 (N_12451,N_7958,N_6689);
xnor U12452 (N_12452,N_5248,N_9547);
nor U12453 (N_12453,N_6597,N_6432);
or U12454 (N_12454,N_6345,N_5044);
xnor U12455 (N_12455,N_6038,N_9656);
nand U12456 (N_12456,N_6363,N_6440);
or U12457 (N_12457,N_9932,N_5929);
or U12458 (N_12458,N_5963,N_5532);
nand U12459 (N_12459,N_9473,N_7512);
xor U12460 (N_12460,N_8053,N_7858);
nand U12461 (N_12461,N_6381,N_9890);
or U12462 (N_12462,N_9342,N_5494);
or U12463 (N_12463,N_9003,N_5823);
or U12464 (N_12464,N_8940,N_6442);
xor U12465 (N_12465,N_5611,N_7138);
nand U12466 (N_12466,N_6035,N_9165);
xor U12467 (N_12467,N_9678,N_7415);
nor U12468 (N_12468,N_9754,N_6888);
and U12469 (N_12469,N_8450,N_5126);
and U12470 (N_12470,N_5828,N_9196);
nand U12471 (N_12471,N_8231,N_6044);
or U12472 (N_12472,N_7610,N_5766);
and U12473 (N_12473,N_6727,N_6357);
nand U12474 (N_12474,N_7386,N_7549);
xor U12475 (N_12475,N_9759,N_9398);
and U12476 (N_12476,N_9075,N_8636);
nand U12477 (N_12477,N_7026,N_7626);
xnor U12478 (N_12478,N_8505,N_9358);
xor U12479 (N_12479,N_8638,N_5094);
xnor U12480 (N_12480,N_5403,N_5208);
xor U12481 (N_12481,N_6736,N_9947);
nor U12482 (N_12482,N_9120,N_9991);
xor U12483 (N_12483,N_6720,N_9324);
nand U12484 (N_12484,N_6840,N_9657);
and U12485 (N_12485,N_7595,N_7067);
and U12486 (N_12486,N_7466,N_8906);
xnor U12487 (N_12487,N_9960,N_8600);
nor U12488 (N_12488,N_7896,N_7660);
xor U12489 (N_12489,N_5012,N_6343);
and U12490 (N_12490,N_6998,N_5882);
and U12491 (N_12491,N_8130,N_5502);
or U12492 (N_12492,N_5909,N_7456);
nand U12493 (N_12493,N_8569,N_7091);
nand U12494 (N_12494,N_8255,N_9772);
and U12495 (N_12495,N_5917,N_9673);
nand U12496 (N_12496,N_8390,N_7407);
or U12497 (N_12497,N_8083,N_9048);
nor U12498 (N_12498,N_9333,N_5133);
and U12499 (N_12499,N_5575,N_9729);
nor U12500 (N_12500,N_8012,N_6229);
or U12501 (N_12501,N_8661,N_6851);
or U12502 (N_12502,N_8558,N_8744);
and U12503 (N_12503,N_8761,N_8431);
nor U12504 (N_12504,N_5332,N_9463);
and U12505 (N_12505,N_9688,N_7351);
or U12506 (N_12506,N_5413,N_7505);
xor U12507 (N_12507,N_7914,N_7619);
and U12508 (N_12508,N_9800,N_5937);
or U12509 (N_12509,N_7707,N_6395);
xor U12510 (N_12510,N_7437,N_6973);
nor U12511 (N_12511,N_5686,N_7851);
nor U12512 (N_12512,N_9901,N_9389);
and U12513 (N_12513,N_5604,N_7168);
or U12514 (N_12514,N_6015,N_6234);
xor U12515 (N_12515,N_6984,N_6701);
nand U12516 (N_12516,N_6473,N_7046);
xnor U12517 (N_12517,N_7951,N_5889);
and U12518 (N_12518,N_6472,N_7058);
and U12519 (N_12519,N_7237,N_9863);
xnor U12520 (N_12520,N_7268,N_7820);
and U12521 (N_12521,N_5403,N_7672);
xor U12522 (N_12522,N_7009,N_7436);
nand U12523 (N_12523,N_7963,N_5796);
and U12524 (N_12524,N_9142,N_9077);
nand U12525 (N_12525,N_9599,N_7655);
nand U12526 (N_12526,N_5331,N_9629);
and U12527 (N_12527,N_5507,N_9923);
and U12528 (N_12528,N_7286,N_7488);
nand U12529 (N_12529,N_6717,N_7639);
and U12530 (N_12530,N_5050,N_7565);
xnor U12531 (N_12531,N_5621,N_6261);
nand U12532 (N_12532,N_6810,N_7067);
and U12533 (N_12533,N_5248,N_9535);
nand U12534 (N_12534,N_6686,N_5834);
or U12535 (N_12535,N_9675,N_5438);
and U12536 (N_12536,N_8101,N_6348);
nor U12537 (N_12537,N_9140,N_6152);
nor U12538 (N_12538,N_5625,N_7082);
or U12539 (N_12539,N_9064,N_9054);
nor U12540 (N_12540,N_7144,N_5390);
and U12541 (N_12541,N_6284,N_6154);
xor U12542 (N_12542,N_5346,N_8350);
nand U12543 (N_12543,N_5123,N_6065);
xor U12544 (N_12544,N_5129,N_6709);
nand U12545 (N_12545,N_5126,N_5165);
and U12546 (N_12546,N_5540,N_8362);
and U12547 (N_12547,N_6554,N_7040);
nor U12548 (N_12548,N_9060,N_8129);
or U12549 (N_12549,N_8495,N_8105);
or U12550 (N_12550,N_5019,N_5113);
nand U12551 (N_12551,N_8341,N_7201);
xnor U12552 (N_12552,N_8992,N_6652);
nand U12553 (N_12553,N_6311,N_5798);
or U12554 (N_12554,N_7171,N_5609);
or U12555 (N_12555,N_5878,N_8169);
and U12556 (N_12556,N_6401,N_6961);
xnor U12557 (N_12557,N_6494,N_8382);
nand U12558 (N_12558,N_9282,N_7608);
nor U12559 (N_12559,N_9823,N_8684);
xnor U12560 (N_12560,N_9166,N_7446);
nor U12561 (N_12561,N_8652,N_6828);
or U12562 (N_12562,N_6724,N_5353);
and U12563 (N_12563,N_6677,N_6865);
nor U12564 (N_12564,N_9655,N_9090);
xnor U12565 (N_12565,N_7346,N_7962);
or U12566 (N_12566,N_8578,N_6685);
and U12567 (N_12567,N_7275,N_5834);
or U12568 (N_12568,N_7846,N_9903);
and U12569 (N_12569,N_5124,N_7380);
nor U12570 (N_12570,N_9701,N_7009);
nand U12571 (N_12571,N_5270,N_6120);
and U12572 (N_12572,N_9461,N_8421);
xor U12573 (N_12573,N_5655,N_7044);
xnor U12574 (N_12574,N_8213,N_8550);
nor U12575 (N_12575,N_6268,N_6652);
and U12576 (N_12576,N_9259,N_8811);
xnor U12577 (N_12577,N_6701,N_8517);
and U12578 (N_12578,N_5602,N_8213);
and U12579 (N_12579,N_6624,N_7979);
xnor U12580 (N_12580,N_8436,N_6854);
or U12581 (N_12581,N_5965,N_5950);
and U12582 (N_12582,N_5635,N_7555);
xor U12583 (N_12583,N_7404,N_5688);
and U12584 (N_12584,N_9884,N_7891);
nand U12585 (N_12585,N_6869,N_5855);
and U12586 (N_12586,N_9013,N_5483);
and U12587 (N_12587,N_6056,N_8904);
and U12588 (N_12588,N_5896,N_6802);
or U12589 (N_12589,N_9839,N_6980);
and U12590 (N_12590,N_9027,N_5569);
nor U12591 (N_12591,N_6183,N_9779);
nand U12592 (N_12592,N_8588,N_6373);
and U12593 (N_12593,N_8867,N_7756);
xnor U12594 (N_12594,N_8745,N_5912);
and U12595 (N_12595,N_6985,N_9741);
nand U12596 (N_12596,N_9945,N_8554);
xnor U12597 (N_12597,N_9038,N_7439);
xnor U12598 (N_12598,N_5290,N_5703);
nor U12599 (N_12599,N_8530,N_8860);
nor U12600 (N_12600,N_7568,N_7674);
nand U12601 (N_12601,N_6701,N_8462);
and U12602 (N_12602,N_9942,N_5209);
xor U12603 (N_12603,N_6800,N_9638);
nor U12604 (N_12604,N_9910,N_7781);
and U12605 (N_12605,N_7532,N_7787);
and U12606 (N_12606,N_8959,N_5148);
nand U12607 (N_12607,N_6892,N_9606);
xor U12608 (N_12608,N_5131,N_7360);
and U12609 (N_12609,N_7583,N_8912);
nand U12610 (N_12610,N_8680,N_8052);
or U12611 (N_12611,N_9255,N_7714);
and U12612 (N_12612,N_7444,N_8286);
nand U12613 (N_12613,N_9306,N_7524);
nand U12614 (N_12614,N_6178,N_8670);
nor U12615 (N_12615,N_9483,N_5532);
nor U12616 (N_12616,N_8791,N_7555);
or U12617 (N_12617,N_7631,N_6998);
and U12618 (N_12618,N_6244,N_5610);
and U12619 (N_12619,N_5479,N_7092);
nor U12620 (N_12620,N_7995,N_8843);
or U12621 (N_12621,N_7037,N_7286);
nor U12622 (N_12622,N_8321,N_7115);
or U12623 (N_12623,N_8335,N_8351);
or U12624 (N_12624,N_5984,N_5306);
or U12625 (N_12625,N_9548,N_8078);
and U12626 (N_12626,N_7413,N_7414);
nor U12627 (N_12627,N_6645,N_8119);
and U12628 (N_12628,N_8738,N_8506);
and U12629 (N_12629,N_7016,N_7114);
xor U12630 (N_12630,N_6602,N_9777);
or U12631 (N_12631,N_8291,N_8021);
nand U12632 (N_12632,N_8246,N_5841);
nor U12633 (N_12633,N_7143,N_7382);
nor U12634 (N_12634,N_8160,N_8726);
or U12635 (N_12635,N_6637,N_9785);
or U12636 (N_12636,N_9470,N_6750);
nand U12637 (N_12637,N_6212,N_5235);
nor U12638 (N_12638,N_9702,N_7127);
nor U12639 (N_12639,N_6432,N_9212);
xor U12640 (N_12640,N_6534,N_8390);
nor U12641 (N_12641,N_9896,N_6552);
or U12642 (N_12642,N_7108,N_8127);
xnor U12643 (N_12643,N_5793,N_8485);
xor U12644 (N_12644,N_6480,N_9860);
nand U12645 (N_12645,N_6585,N_9632);
and U12646 (N_12646,N_7859,N_8024);
nor U12647 (N_12647,N_8463,N_8482);
nor U12648 (N_12648,N_7015,N_9974);
or U12649 (N_12649,N_7323,N_9369);
or U12650 (N_12650,N_5421,N_7943);
or U12651 (N_12651,N_5749,N_6463);
or U12652 (N_12652,N_9140,N_5756);
xor U12653 (N_12653,N_5151,N_9158);
and U12654 (N_12654,N_9172,N_5886);
nand U12655 (N_12655,N_7807,N_9075);
and U12656 (N_12656,N_6182,N_6782);
nor U12657 (N_12657,N_8118,N_5526);
or U12658 (N_12658,N_5389,N_7159);
nor U12659 (N_12659,N_6703,N_6381);
and U12660 (N_12660,N_9394,N_5952);
and U12661 (N_12661,N_6024,N_5755);
nor U12662 (N_12662,N_6806,N_6286);
and U12663 (N_12663,N_8998,N_5770);
xnor U12664 (N_12664,N_7578,N_6822);
nand U12665 (N_12665,N_7407,N_7904);
nand U12666 (N_12666,N_9339,N_7466);
xnor U12667 (N_12667,N_9957,N_5695);
or U12668 (N_12668,N_6743,N_7411);
and U12669 (N_12669,N_8143,N_6380);
nor U12670 (N_12670,N_9382,N_8223);
or U12671 (N_12671,N_8534,N_9391);
or U12672 (N_12672,N_5239,N_8822);
nor U12673 (N_12673,N_7247,N_9047);
nor U12674 (N_12674,N_6651,N_8955);
nand U12675 (N_12675,N_8498,N_7121);
and U12676 (N_12676,N_5990,N_7911);
xor U12677 (N_12677,N_9440,N_9035);
or U12678 (N_12678,N_6044,N_5524);
or U12679 (N_12679,N_6525,N_7700);
nor U12680 (N_12680,N_9354,N_5863);
nor U12681 (N_12681,N_9354,N_9276);
nand U12682 (N_12682,N_9857,N_6829);
or U12683 (N_12683,N_6645,N_5909);
xnor U12684 (N_12684,N_8365,N_7181);
or U12685 (N_12685,N_5233,N_8277);
and U12686 (N_12686,N_9475,N_6725);
xnor U12687 (N_12687,N_5952,N_5622);
and U12688 (N_12688,N_6215,N_5827);
nand U12689 (N_12689,N_9874,N_7863);
xnor U12690 (N_12690,N_8749,N_5992);
nand U12691 (N_12691,N_6011,N_5766);
or U12692 (N_12692,N_8007,N_8907);
nor U12693 (N_12693,N_6228,N_9768);
and U12694 (N_12694,N_7295,N_9212);
xnor U12695 (N_12695,N_9977,N_9140);
nor U12696 (N_12696,N_9809,N_8846);
nand U12697 (N_12697,N_7392,N_6016);
nand U12698 (N_12698,N_6753,N_7471);
xor U12699 (N_12699,N_7108,N_7055);
nand U12700 (N_12700,N_7908,N_7067);
nand U12701 (N_12701,N_6163,N_6526);
or U12702 (N_12702,N_9197,N_8803);
xnor U12703 (N_12703,N_9843,N_9907);
or U12704 (N_12704,N_9454,N_6012);
xnor U12705 (N_12705,N_7309,N_5246);
or U12706 (N_12706,N_5433,N_6274);
nor U12707 (N_12707,N_5812,N_5655);
nand U12708 (N_12708,N_6657,N_5522);
nand U12709 (N_12709,N_6630,N_5563);
xnor U12710 (N_12710,N_5003,N_9847);
or U12711 (N_12711,N_6125,N_7485);
nor U12712 (N_12712,N_6486,N_8062);
nor U12713 (N_12713,N_9818,N_7350);
or U12714 (N_12714,N_8971,N_5922);
or U12715 (N_12715,N_7266,N_5062);
nor U12716 (N_12716,N_6841,N_9482);
nor U12717 (N_12717,N_7478,N_7406);
and U12718 (N_12718,N_6954,N_5414);
nor U12719 (N_12719,N_9539,N_6120);
nor U12720 (N_12720,N_8264,N_9506);
nand U12721 (N_12721,N_9341,N_8433);
and U12722 (N_12722,N_7770,N_9997);
xnor U12723 (N_12723,N_7829,N_5664);
nand U12724 (N_12724,N_7975,N_7751);
nand U12725 (N_12725,N_7824,N_9746);
xor U12726 (N_12726,N_5120,N_8236);
nand U12727 (N_12727,N_9640,N_5616);
xnor U12728 (N_12728,N_9146,N_5888);
and U12729 (N_12729,N_8822,N_9342);
and U12730 (N_12730,N_7157,N_7337);
xnor U12731 (N_12731,N_5958,N_8001);
nor U12732 (N_12732,N_8492,N_5446);
nand U12733 (N_12733,N_9245,N_8330);
and U12734 (N_12734,N_5704,N_5339);
nand U12735 (N_12735,N_8359,N_5263);
and U12736 (N_12736,N_7092,N_7661);
xnor U12737 (N_12737,N_7487,N_6020);
nor U12738 (N_12738,N_8061,N_8526);
or U12739 (N_12739,N_8134,N_8437);
and U12740 (N_12740,N_8188,N_8695);
nand U12741 (N_12741,N_9957,N_6032);
xnor U12742 (N_12742,N_6954,N_7105);
xnor U12743 (N_12743,N_5721,N_8192);
or U12744 (N_12744,N_9942,N_7152);
and U12745 (N_12745,N_7648,N_7485);
nor U12746 (N_12746,N_7719,N_8998);
or U12747 (N_12747,N_7777,N_5784);
nand U12748 (N_12748,N_6131,N_8425);
and U12749 (N_12749,N_8263,N_9192);
and U12750 (N_12750,N_7666,N_7595);
or U12751 (N_12751,N_5396,N_6474);
and U12752 (N_12752,N_6355,N_5977);
xor U12753 (N_12753,N_5949,N_6968);
xnor U12754 (N_12754,N_6266,N_7907);
xor U12755 (N_12755,N_6811,N_9029);
xor U12756 (N_12756,N_9182,N_5478);
nand U12757 (N_12757,N_5997,N_9651);
nand U12758 (N_12758,N_6023,N_7825);
or U12759 (N_12759,N_6474,N_9333);
nand U12760 (N_12760,N_9876,N_7135);
nor U12761 (N_12761,N_7528,N_5450);
and U12762 (N_12762,N_7939,N_9331);
xor U12763 (N_12763,N_6024,N_7400);
nor U12764 (N_12764,N_6593,N_5714);
and U12765 (N_12765,N_5891,N_5876);
nor U12766 (N_12766,N_7514,N_9992);
and U12767 (N_12767,N_8944,N_8136);
nand U12768 (N_12768,N_7321,N_7331);
nor U12769 (N_12769,N_7924,N_5189);
or U12770 (N_12770,N_8660,N_5134);
xnor U12771 (N_12771,N_6247,N_5234);
and U12772 (N_12772,N_8618,N_7765);
or U12773 (N_12773,N_9449,N_6935);
nand U12774 (N_12774,N_5669,N_9181);
and U12775 (N_12775,N_7895,N_5106);
nor U12776 (N_12776,N_8773,N_9782);
or U12777 (N_12777,N_9566,N_9914);
and U12778 (N_12778,N_8289,N_7031);
and U12779 (N_12779,N_6521,N_9796);
and U12780 (N_12780,N_8217,N_8952);
nor U12781 (N_12781,N_6507,N_8503);
or U12782 (N_12782,N_8666,N_8567);
or U12783 (N_12783,N_7500,N_7365);
or U12784 (N_12784,N_5439,N_5465);
and U12785 (N_12785,N_8484,N_6949);
nand U12786 (N_12786,N_9272,N_8181);
nor U12787 (N_12787,N_9717,N_7382);
nor U12788 (N_12788,N_9499,N_7636);
and U12789 (N_12789,N_7445,N_8146);
and U12790 (N_12790,N_7596,N_6181);
or U12791 (N_12791,N_7279,N_9412);
nand U12792 (N_12792,N_5483,N_6910);
nor U12793 (N_12793,N_6043,N_7982);
and U12794 (N_12794,N_8916,N_7126);
nor U12795 (N_12795,N_8806,N_6463);
and U12796 (N_12796,N_8692,N_6852);
xnor U12797 (N_12797,N_7750,N_7608);
or U12798 (N_12798,N_6602,N_5929);
or U12799 (N_12799,N_9224,N_5252);
xnor U12800 (N_12800,N_7060,N_6762);
nand U12801 (N_12801,N_7888,N_9715);
nor U12802 (N_12802,N_7178,N_6108);
xnor U12803 (N_12803,N_5714,N_5175);
and U12804 (N_12804,N_5404,N_6957);
and U12805 (N_12805,N_5053,N_9733);
or U12806 (N_12806,N_9711,N_6433);
and U12807 (N_12807,N_9789,N_9291);
nand U12808 (N_12808,N_8116,N_5401);
nor U12809 (N_12809,N_8018,N_8044);
nand U12810 (N_12810,N_9166,N_6236);
xor U12811 (N_12811,N_8863,N_7700);
or U12812 (N_12812,N_7540,N_7720);
or U12813 (N_12813,N_5006,N_9499);
nor U12814 (N_12814,N_9792,N_7685);
or U12815 (N_12815,N_9529,N_7962);
and U12816 (N_12816,N_6471,N_8316);
or U12817 (N_12817,N_7590,N_5610);
and U12818 (N_12818,N_5612,N_7519);
nor U12819 (N_12819,N_5798,N_6754);
nor U12820 (N_12820,N_8214,N_6970);
or U12821 (N_12821,N_6117,N_6902);
and U12822 (N_12822,N_8031,N_5943);
nand U12823 (N_12823,N_6830,N_9381);
nand U12824 (N_12824,N_6641,N_6478);
nand U12825 (N_12825,N_8787,N_8991);
nand U12826 (N_12826,N_7182,N_8946);
and U12827 (N_12827,N_6484,N_8449);
and U12828 (N_12828,N_6340,N_9296);
xor U12829 (N_12829,N_7024,N_6315);
nor U12830 (N_12830,N_5828,N_5364);
or U12831 (N_12831,N_7866,N_5561);
or U12832 (N_12832,N_6356,N_5333);
nor U12833 (N_12833,N_5443,N_5133);
xor U12834 (N_12834,N_7827,N_7800);
or U12835 (N_12835,N_6179,N_8752);
nand U12836 (N_12836,N_7411,N_8094);
or U12837 (N_12837,N_5869,N_7885);
nor U12838 (N_12838,N_7161,N_9726);
xor U12839 (N_12839,N_5324,N_9862);
and U12840 (N_12840,N_7789,N_8193);
nor U12841 (N_12841,N_8689,N_8789);
xor U12842 (N_12842,N_6720,N_8943);
and U12843 (N_12843,N_7091,N_7748);
nand U12844 (N_12844,N_6433,N_7242);
nor U12845 (N_12845,N_6286,N_7388);
nand U12846 (N_12846,N_9687,N_6605);
nand U12847 (N_12847,N_6085,N_7320);
nor U12848 (N_12848,N_9773,N_9410);
or U12849 (N_12849,N_6105,N_9896);
xor U12850 (N_12850,N_9136,N_5395);
and U12851 (N_12851,N_7757,N_6610);
and U12852 (N_12852,N_6181,N_9873);
nor U12853 (N_12853,N_5520,N_5700);
or U12854 (N_12854,N_5268,N_7003);
or U12855 (N_12855,N_9325,N_9638);
nor U12856 (N_12856,N_9953,N_5820);
nor U12857 (N_12857,N_6884,N_6246);
xor U12858 (N_12858,N_8876,N_7690);
or U12859 (N_12859,N_8123,N_7796);
nand U12860 (N_12860,N_6096,N_9306);
xnor U12861 (N_12861,N_8936,N_6350);
xor U12862 (N_12862,N_8832,N_7811);
nand U12863 (N_12863,N_5739,N_9103);
xor U12864 (N_12864,N_6767,N_5834);
nor U12865 (N_12865,N_9724,N_7090);
or U12866 (N_12866,N_7217,N_5255);
xnor U12867 (N_12867,N_8419,N_5103);
nor U12868 (N_12868,N_9315,N_6266);
xnor U12869 (N_12869,N_7842,N_8811);
or U12870 (N_12870,N_9042,N_5381);
xor U12871 (N_12871,N_6912,N_5695);
or U12872 (N_12872,N_6937,N_5885);
and U12873 (N_12873,N_6373,N_8039);
xor U12874 (N_12874,N_6396,N_9318);
nor U12875 (N_12875,N_5203,N_9782);
nand U12876 (N_12876,N_6322,N_5411);
and U12877 (N_12877,N_7469,N_5248);
or U12878 (N_12878,N_8222,N_9618);
or U12879 (N_12879,N_6601,N_8275);
xor U12880 (N_12880,N_8684,N_7239);
nor U12881 (N_12881,N_8039,N_9054);
or U12882 (N_12882,N_7539,N_8464);
xor U12883 (N_12883,N_8120,N_8732);
nor U12884 (N_12884,N_8585,N_8248);
nand U12885 (N_12885,N_7893,N_7558);
nand U12886 (N_12886,N_9730,N_9822);
or U12887 (N_12887,N_5964,N_5782);
xor U12888 (N_12888,N_6863,N_9118);
or U12889 (N_12889,N_5078,N_6157);
xor U12890 (N_12890,N_9081,N_9741);
nor U12891 (N_12891,N_7038,N_8540);
and U12892 (N_12892,N_9363,N_9119);
or U12893 (N_12893,N_7452,N_6358);
or U12894 (N_12894,N_7706,N_8613);
or U12895 (N_12895,N_5830,N_8093);
or U12896 (N_12896,N_7825,N_5922);
nand U12897 (N_12897,N_7621,N_6266);
xor U12898 (N_12898,N_9479,N_6979);
or U12899 (N_12899,N_6842,N_8044);
xnor U12900 (N_12900,N_8471,N_8411);
xnor U12901 (N_12901,N_9203,N_7229);
nand U12902 (N_12902,N_5879,N_6104);
xnor U12903 (N_12903,N_8302,N_5243);
nor U12904 (N_12904,N_6935,N_5847);
nor U12905 (N_12905,N_9503,N_7026);
nor U12906 (N_12906,N_9316,N_5338);
or U12907 (N_12907,N_7839,N_7997);
nor U12908 (N_12908,N_9773,N_6943);
and U12909 (N_12909,N_7358,N_5674);
and U12910 (N_12910,N_8991,N_8748);
nand U12911 (N_12911,N_8374,N_9065);
and U12912 (N_12912,N_8852,N_8738);
and U12913 (N_12913,N_9763,N_8564);
or U12914 (N_12914,N_8007,N_6923);
nand U12915 (N_12915,N_9049,N_8240);
nor U12916 (N_12916,N_9546,N_7277);
xor U12917 (N_12917,N_6223,N_5065);
nand U12918 (N_12918,N_6622,N_6722);
nand U12919 (N_12919,N_7915,N_7132);
xnor U12920 (N_12920,N_6778,N_7606);
or U12921 (N_12921,N_9175,N_8351);
and U12922 (N_12922,N_7304,N_5590);
and U12923 (N_12923,N_8271,N_6914);
and U12924 (N_12924,N_8101,N_8673);
nor U12925 (N_12925,N_6320,N_7170);
xor U12926 (N_12926,N_7019,N_7863);
xor U12927 (N_12927,N_6241,N_5998);
or U12928 (N_12928,N_9326,N_8225);
nor U12929 (N_12929,N_5806,N_7173);
nand U12930 (N_12930,N_5909,N_9780);
xnor U12931 (N_12931,N_5215,N_9792);
or U12932 (N_12932,N_8649,N_5644);
nor U12933 (N_12933,N_8774,N_6769);
nand U12934 (N_12934,N_5286,N_7771);
or U12935 (N_12935,N_8554,N_5632);
and U12936 (N_12936,N_8710,N_6310);
nor U12937 (N_12937,N_6932,N_8797);
xnor U12938 (N_12938,N_8037,N_7734);
and U12939 (N_12939,N_5578,N_6019);
and U12940 (N_12940,N_8780,N_6930);
nand U12941 (N_12941,N_7791,N_5260);
xnor U12942 (N_12942,N_9050,N_8367);
nand U12943 (N_12943,N_5961,N_6544);
and U12944 (N_12944,N_6240,N_8102);
nand U12945 (N_12945,N_8276,N_8848);
or U12946 (N_12946,N_6791,N_6276);
and U12947 (N_12947,N_7604,N_5011);
nor U12948 (N_12948,N_6359,N_5272);
nand U12949 (N_12949,N_7029,N_6447);
xor U12950 (N_12950,N_9359,N_8491);
or U12951 (N_12951,N_9475,N_8364);
nor U12952 (N_12952,N_6788,N_5123);
nor U12953 (N_12953,N_9230,N_9055);
nor U12954 (N_12954,N_6216,N_7147);
xnor U12955 (N_12955,N_6635,N_6195);
nand U12956 (N_12956,N_6154,N_5197);
and U12957 (N_12957,N_6809,N_8347);
xnor U12958 (N_12958,N_6819,N_5416);
xnor U12959 (N_12959,N_8541,N_7737);
or U12960 (N_12960,N_8730,N_6057);
nand U12961 (N_12961,N_8665,N_9109);
and U12962 (N_12962,N_8423,N_8631);
xor U12963 (N_12963,N_8186,N_9515);
and U12964 (N_12964,N_5368,N_9325);
xor U12965 (N_12965,N_5188,N_6668);
nand U12966 (N_12966,N_9234,N_9750);
or U12967 (N_12967,N_7550,N_5415);
nand U12968 (N_12968,N_7297,N_9427);
or U12969 (N_12969,N_6976,N_8180);
nand U12970 (N_12970,N_6624,N_5051);
xor U12971 (N_12971,N_6081,N_5024);
and U12972 (N_12972,N_7312,N_9833);
nor U12973 (N_12973,N_5487,N_6044);
xor U12974 (N_12974,N_7755,N_9248);
and U12975 (N_12975,N_8384,N_9048);
nor U12976 (N_12976,N_7428,N_7571);
or U12977 (N_12977,N_6324,N_6938);
nand U12978 (N_12978,N_5684,N_5889);
nor U12979 (N_12979,N_8177,N_9052);
nor U12980 (N_12980,N_9421,N_5501);
nand U12981 (N_12981,N_7279,N_5484);
nor U12982 (N_12982,N_8678,N_9595);
and U12983 (N_12983,N_7880,N_8378);
xnor U12984 (N_12984,N_6500,N_5247);
nand U12985 (N_12985,N_8009,N_5939);
nand U12986 (N_12986,N_7484,N_7357);
xor U12987 (N_12987,N_7796,N_6342);
nor U12988 (N_12988,N_5792,N_9985);
and U12989 (N_12989,N_8263,N_8235);
nand U12990 (N_12990,N_5256,N_6485);
nor U12991 (N_12991,N_8225,N_7189);
and U12992 (N_12992,N_7523,N_9433);
xnor U12993 (N_12993,N_7939,N_5301);
nand U12994 (N_12994,N_6498,N_8698);
nor U12995 (N_12995,N_9360,N_8818);
and U12996 (N_12996,N_5377,N_6017);
nand U12997 (N_12997,N_9195,N_5684);
nand U12998 (N_12998,N_6419,N_9028);
or U12999 (N_12999,N_8850,N_6417);
nand U13000 (N_13000,N_8827,N_5834);
nor U13001 (N_13001,N_7407,N_8942);
nor U13002 (N_13002,N_9487,N_5331);
nor U13003 (N_13003,N_5694,N_8289);
and U13004 (N_13004,N_5158,N_9750);
and U13005 (N_13005,N_7827,N_7913);
and U13006 (N_13006,N_5044,N_9152);
xor U13007 (N_13007,N_9185,N_8423);
or U13008 (N_13008,N_6650,N_8513);
or U13009 (N_13009,N_5173,N_5068);
or U13010 (N_13010,N_6181,N_7866);
nand U13011 (N_13011,N_9200,N_7750);
and U13012 (N_13012,N_8288,N_8207);
xnor U13013 (N_13013,N_9878,N_5359);
nand U13014 (N_13014,N_8202,N_7568);
and U13015 (N_13015,N_8783,N_9594);
nor U13016 (N_13016,N_7687,N_6438);
and U13017 (N_13017,N_7542,N_5336);
nand U13018 (N_13018,N_8879,N_5049);
nand U13019 (N_13019,N_6474,N_6212);
xnor U13020 (N_13020,N_7996,N_9298);
nand U13021 (N_13021,N_5238,N_5912);
xor U13022 (N_13022,N_9776,N_9919);
xor U13023 (N_13023,N_5716,N_9365);
nand U13024 (N_13024,N_5210,N_6188);
or U13025 (N_13025,N_7326,N_8130);
xnor U13026 (N_13026,N_9354,N_9976);
nor U13027 (N_13027,N_5598,N_5952);
nand U13028 (N_13028,N_7506,N_6438);
nor U13029 (N_13029,N_7664,N_6328);
nor U13030 (N_13030,N_9565,N_9271);
xor U13031 (N_13031,N_5752,N_7150);
xnor U13032 (N_13032,N_5153,N_8033);
nor U13033 (N_13033,N_6067,N_9037);
xor U13034 (N_13034,N_5085,N_7079);
nor U13035 (N_13035,N_7732,N_5350);
nand U13036 (N_13036,N_5827,N_6844);
xnor U13037 (N_13037,N_5920,N_9587);
or U13038 (N_13038,N_9006,N_8835);
and U13039 (N_13039,N_7073,N_6562);
xor U13040 (N_13040,N_5836,N_7001);
or U13041 (N_13041,N_6783,N_9892);
nor U13042 (N_13042,N_8011,N_5315);
xor U13043 (N_13043,N_5801,N_8300);
nor U13044 (N_13044,N_8740,N_8945);
nor U13045 (N_13045,N_5785,N_8430);
xnor U13046 (N_13046,N_7794,N_5915);
nand U13047 (N_13047,N_8199,N_5794);
nand U13048 (N_13048,N_8397,N_7445);
nand U13049 (N_13049,N_8123,N_6722);
nand U13050 (N_13050,N_5771,N_7588);
nor U13051 (N_13051,N_6352,N_9019);
nand U13052 (N_13052,N_5207,N_7071);
nor U13053 (N_13053,N_5871,N_8881);
and U13054 (N_13054,N_8550,N_9809);
or U13055 (N_13055,N_5867,N_5032);
nand U13056 (N_13056,N_7123,N_7655);
and U13057 (N_13057,N_9273,N_5102);
and U13058 (N_13058,N_8625,N_5554);
or U13059 (N_13059,N_9515,N_5308);
nand U13060 (N_13060,N_5768,N_7533);
or U13061 (N_13061,N_8743,N_7684);
xor U13062 (N_13062,N_9309,N_5825);
or U13063 (N_13063,N_5618,N_6569);
nand U13064 (N_13064,N_5731,N_6937);
or U13065 (N_13065,N_7844,N_6511);
and U13066 (N_13066,N_9641,N_5550);
or U13067 (N_13067,N_5424,N_9028);
xor U13068 (N_13068,N_6074,N_9165);
nor U13069 (N_13069,N_6315,N_6576);
or U13070 (N_13070,N_5984,N_6389);
xnor U13071 (N_13071,N_9614,N_5046);
or U13072 (N_13072,N_5053,N_7440);
or U13073 (N_13073,N_8045,N_7513);
and U13074 (N_13074,N_7387,N_5272);
or U13075 (N_13075,N_7352,N_9665);
or U13076 (N_13076,N_6174,N_9988);
xor U13077 (N_13077,N_5693,N_9275);
or U13078 (N_13078,N_6384,N_9837);
nand U13079 (N_13079,N_6625,N_7915);
and U13080 (N_13080,N_7463,N_7616);
nor U13081 (N_13081,N_6590,N_6554);
nand U13082 (N_13082,N_7115,N_5734);
nand U13083 (N_13083,N_5392,N_9622);
nand U13084 (N_13084,N_9074,N_8067);
nand U13085 (N_13085,N_5906,N_8601);
or U13086 (N_13086,N_7538,N_5385);
nor U13087 (N_13087,N_6576,N_9544);
or U13088 (N_13088,N_8816,N_9118);
nor U13089 (N_13089,N_5849,N_8131);
xnor U13090 (N_13090,N_9796,N_5019);
and U13091 (N_13091,N_8935,N_8622);
xor U13092 (N_13092,N_6986,N_9766);
xnor U13093 (N_13093,N_6150,N_7963);
and U13094 (N_13094,N_9142,N_8505);
nand U13095 (N_13095,N_7140,N_6859);
and U13096 (N_13096,N_5825,N_9869);
nand U13097 (N_13097,N_6401,N_6220);
nand U13098 (N_13098,N_8259,N_8216);
nand U13099 (N_13099,N_7307,N_9975);
or U13100 (N_13100,N_7583,N_7326);
xnor U13101 (N_13101,N_5223,N_8642);
or U13102 (N_13102,N_6652,N_9410);
or U13103 (N_13103,N_5155,N_6087);
and U13104 (N_13104,N_5492,N_8145);
nand U13105 (N_13105,N_6384,N_6329);
nor U13106 (N_13106,N_5703,N_5252);
or U13107 (N_13107,N_7940,N_7107);
and U13108 (N_13108,N_5669,N_8465);
and U13109 (N_13109,N_5164,N_8993);
xnor U13110 (N_13110,N_8584,N_6766);
nand U13111 (N_13111,N_6396,N_5804);
and U13112 (N_13112,N_6201,N_8245);
or U13113 (N_13113,N_5152,N_5369);
and U13114 (N_13114,N_7700,N_6027);
nand U13115 (N_13115,N_5301,N_9287);
xnor U13116 (N_13116,N_7407,N_5235);
nor U13117 (N_13117,N_8690,N_6474);
xor U13118 (N_13118,N_9353,N_6579);
xor U13119 (N_13119,N_5184,N_9623);
xor U13120 (N_13120,N_8198,N_9538);
xor U13121 (N_13121,N_9361,N_8396);
xnor U13122 (N_13122,N_6357,N_7617);
nand U13123 (N_13123,N_6208,N_6693);
nand U13124 (N_13124,N_6777,N_9320);
and U13125 (N_13125,N_8220,N_8718);
and U13126 (N_13126,N_7027,N_8297);
xnor U13127 (N_13127,N_8920,N_8994);
xor U13128 (N_13128,N_5164,N_8108);
nor U13129 (N_13129,N_9059,N_6077);
nand U13130 (N_13130,N_8214,N_7877);
xnor U13131 (N_13131,N_8664,N_7103);
xor U13132 (N_13132,N_5344,N_8852);
nor U13133 (N_13133,N_9113,N_7046);
nor U13134 (N_13134,N_5038,N_6190);
nor U13135 (N_13135,N_8804,N_8333);
and U13136 (N_13136,N_5668,N_8166);
nand U13137 (N_13137,N_7669,N_9766);
xor U13138 (N_13138,N_8489,N_9075);
and U13139 (N_13139,N_6785,N_5010);
nand U13140 (N_13140,N_8803,N_7165);
and U13141 (N_13141,N_9623,N_6852);
nor U13142 (N_13142,N_8002,N_9226);
xnor U13143 (N_13143,N_9278,N_7741);
nor U13144 (N_13144,N_5302,N_9722);
xor U13145 (N_13145,N_8824,N_5872);
nor U13146 (N_13146,N_8164,N_7790);
or U13147 (N_13147,N_5778,N_5140);
or U13148 (N_13148,N_7963,N_7920);
xor U13149 (N_13149,N_6853,N_8797);
or U13150 (N_13150,N_7913,N_8517);
nor U13151 (N_13151,N_8221,N_6354);
or U13152 (N_13152,N_8473,N_5674);
and U13153 (N_13153,N_8803,N_7738);
and U13154 (N_13154,N_5101,N_8787);
nor U13155 (N_13155,N_8911,N_7063);
or U13156 (N_13156,N_8347,N_9553);
nor U13157 (N_13157,N_8230,N_6779);
nor U13158 (N_13158,N_6981,N_8042);
nor U13159 (N_13159,N_8487,N_5458);
nand U13160 (N_13160,N_8813,N_8591);
or U13161 (N_13161,N_6625,N_7241);
or U13162 (N_13162,N_5008,N_5485);
or U13163 (N_13163,N_9306,N_5682);
xnor U13164 (N_13164,N_7039,N_7728);
or U13165 (N_13165,N_6640,N_7526);
nand U13166 (N_13166,N_6651,N_6764);
and U13167 (N_13167,N_7444,N_5481);
xor U13168 (N_13168,N_9814,N_8651);
nor U13169 (N_13169,N_5128,N_6665);
or U13170 (N_13170,N_5006,N_6463);
nor U13171 (N_13171,N_5153,N_5378);
and U13172 (N_13172,N_7522,N_5741);
and U13173 (N_13173,N_8950,N_9422);
xor U13174 (N_13174,N_6477,N_5742);
nand U13175 (N_13175,N_7686,N_9021);
nand U13176 (N_13176,N_6361,N_9845);
or U13177 (N_13177,N_7066,N_8029);
xor U13178 (N_13178,N_8308,N_8381);
nand U13179 (N_13179,N_5425,N_8897);
nor U13180 (N_13180,N_6769,N_9066);
nand U13181 (N_13181,N_8175,N_5876);
or U13182 (N_13182,N_7433,N_6619);
and U13183 (N_13183,N_7930,N_7439);
nand U13184 (N_13184,N_5080,N_5257);
and U13185 (N_13185,N_7230,N_5593);
or U13186 (N_13186,N_7334,N_7228);
or U13187 (N_13187,N_7368,N_5442);
and U13188 (N_13188,N_5442,N_9166);
xnor U13189 (N_13189,N_8264,N_8001);
xnor U13190 (N_13190,N_6958,N_5417);
xnor U13191 (N_13191,N_8528,N_6856);
or U13192 (N_13192,N_8407,N_7958);
and U13193 (N_13193,N_7936,N_5034);
nor U13194 (N_13194,N_6004,N_9417);
xor U13195 (N_13195,N_6443,N_8300);
nand U13196 (N_13196,N_8455,N_9444);
and U13197 (N_13197,N_5692,N_8028);
nor U13198 (N_13198,N_9053,N_7883);
and U13199 (N_13199,N_7374,N_6038);
nor U13200 (N_13200,N_8035,N_5219);
nand U13201 (N_13201,N_7651,N_5852);
or U13202 (N_13202,N_9875,N_6286);
and U13203 (N_13203,N_9710,N_5918);
and U13204 (N_13204,N_9566,N_5278);
xor U13205 (N_13205,N_6232,N_7732);
xor U13206 (N_13206,N_9198,N_7684);
nand U13207 (N_13207,N_9824,N_7976);
nand U13208 (N_13208,N_8710,N_5984);
nand U13209 (N_13209,N_5684,N_6555);
xor U13210 (N_13210,N_7897,N_5554);
nand U13211 (N_13211,N_8075,N_7516);
and U13212 (N_13212,N_5209,N_5873);
nor U13213 (N_13213,N_9143,N_7730);
or U13214 (N_13214,N_7785,N_8793);
nand U13215 (N_13215,N_7044,N_7152);
nor U13216 (N_13216,N_5623,N_6513);
and U13217 (N_13217,N_7234,N_9225);
nand U13218 (N_13218,N_6093,N_9341);
nor U13219 (N_13219,N_5087,N_9081);
nor U13220 (N_13220,N_9795,N_9711);
nand U13221 (N_13221,N_6129,N_8019);
nand U13222 (N_13222,N_6270,N_8339);
or U13223 (N_13223,N_6905,N_8945);
xor U13224 (N_13224,N_6781,N_8256);
and U13225 (N_13225,N_9805,N_6322);
xnor U13226 (N_13226,N_9200,N_8081);
xor U13227 (N_13227,N_9964,N_6089);
nor U13228 (N_13228,N_5952,N_6930);
nand U13229 (N_13229,N_6676,N_6662);
nand U13230 (N_13230,N_5079,N_5776);
or U13231 (N_13231,N_7044,N_5310);
or U13232 (N_13232,N_7973,N_7888);
and U13233 (N_13233,N_7080,N_7743);
nand U13234 (N_13234,N_7928,N_7372);
nor U13235 (N_13235,N_8230,N_7853);
xor U13236 (N_13236,N_9993,N_9050);
nand U13237 (N_13237,N_7366,N_5486);
nor U13238 (N_13238,N_7491,N_9401);
or U13239 (N_13239,N_6234,N_7344);
nand U13240 (N_13240,N_5938,N_9345);
or U13241 (N_13241,N_9244,N_7276);
nor U13242 (N_13242,N_9364,N_9311);
and U13243 (N_13243,N_8287,N_9109);
and U13244 (N_13244,N_7614,N_9090);
nand U13245 (N_13245,N_6636,N_6240);
xor U13246 (N_13246,N_5887,N_9815);
nor U13247 (N_13247,N_9725,N_6569);
xnor U13248 (N_13248,N_9821,N_7128);
or U13249 (N_13249,N_5683,N_9447);
nor U13250 (N_13250,N_8684,N_8219);
nand U13251 (N_13251,N_7156,N_6033);
nor U13252 (N_13252,N_7801,N_6824);
or U13253 (N_13253,N_8915,N_5322);
or U13254 (N_13254,N_8309,N_8256);
and U13255 (N_13255,N_5996,N_9879);
nand U13256 (N_13256,N_8418,N_7060);
and U13257 (N_13257,N_6332,N_8526);
nand U13258 (N_13258,N_5635,N_5698);
nand U13259 (N_13259,N_5496,N_9335);
nand U13260 (N_13260,N_5791,N_5216);
and U13261 (N_13261,N_6787,N_7590);
and U13262 (N_13262,N_9051,N_5068);
nand U13263 (N_13263,N_9356,N_7037);
nand U13264 (N_13264,N_7432,N_5466);
xor U13265 (N_13265,N_6990,N_9094);
xnor U13266 (N_13266,N_7650,N_9375);
xor U13267 (N_13267,N_7778,N_5144);
nand U13268 (N_13268,N_8612,N_8326);
xnor U13269 (N_13269,N_7171,N_9181);
nand U13270 (N_13270,N_5931,N_5726);
or U13271 (N_13271,N_5184,N_7576);
or U13272 (N_13272,N_6944,N_7447);
xor U13273 (N_13273,N_7351,N_5017);
or U13274 (N_13274,N_5134,N_6939);
xnor U13275 (N_13275,N_6757,N_5752);
xnor U13276 (N_13276,N_7184,N_5886);
nand U13277 (N_13277,N_8054,N_7051);
and U13278 (N_13278,N_6568,N_8547);
xnor U13279 (N_13279,N_6019,N_7234);
and U13280 (N_13280,N_8485,N_9298);
nor U13281 (N_13281,N_5595,N_5246);
nand U13282 (N_13282,N_5919,N_5149);
xnor U13283 (N_13283,N_6924,N_7490);
or U13284 (N_13284,N_8899,N_5956);
and U13285 (N_13285,N_9552,N_7367);
nor U13286 (N_13286,N_7889,N_8122);
or U13287 (N_13287,N_5109,N_9184);
nor U13288 (N_13288,N_5356,N_5310);
or U13289 (N_13289,N_6089,N_6602);
or U13290 (N_13290,N_8606,N_8698);
or U13291 (N_13291,N_6966,N_5056);
xor U13292 (N_13292,N_7656,N_9164);
or U13293 (N_13293,N_7972,N_7063);
nand U13294 (N_13294,N_5482,N_7158);
nand U13295 (N_13295,N_7155,N_5709);
or U13296 (N_13296,N_8110,N_9328);
nor U13297 (N_13297,N_6413,N_9156);
and U13298 (N_13298,N_9104,N_9898);
and U13299 (N_13299,N_5704,N_5261);
nand U13300 (N_13300,N_8115,N_9867);
xnor U13301 (N_13301,N_6986,N_9274);
or U13302 (N_13302,N_8772,N_7763);
and U13303 (N_13303,N_6120,N_6961);
or U13304 (N_13304,N_7512,N_8927);
nand U13305 (N_13305,N_5066,N_6986);
xor U13306 (N_13306,N_6628,N_9506);
nor U13307 (N_13307,N_9389,N_6255);
nand U13308 (N_13308,N_5712,N_5811);
xor U13309 (N_13309,N_8285,N_9736);
and U13310 (N_13310,N_9881,N_7080);
nand U13311 (N_13311,N_7731,N_7521);
or U13312 (N_13312,N_5783,N_6441);
xor U13313 (N_13313,N_9418,N_8200);
or U13314 (N_13314,N_5079,N_9724);
xnor U13315 (N_13315,N_8015,N_6826);
xnor U13316 (N_13316,N_5260,N_6365);
and U13317 (N_13317,N_9491,N_5237);
xnor U13318 (N_13318,N_8496,N_5226);
and U13319 (N_13319,N_5034,N_9656);
or U13320 (N_13320,N_6391,N_9366);
nand U13321 (N_13321,N_5823,N_5916);
or U13322 (N_13322,N_8843,N_6236);
xor U13323 (N_13323,N_5984,N_6343);
nor U13324 (N_13324,N_5929,N_7271);
nand U13325 (N_13325,N_6865,N_6637);
and U13326 (N_13326,N_5000,N_5723);
nand U13327 (N_13327,N_9604,N_6648);
or U13328 (N_13328,N_8276,N_9990);
nor U13329 (N_13329,N_5922,N_9218);
or U13330 (N_13330,N_5996,N_9640);
xnor U13331 (N_13331,N_7518,N_5136);
or U13332 (N_13332,N_6322,N_9493);
nor U13333 (N_13333,N_7217,N_7853);
nor U13334 (N_13334,N_5032,N_9019);
or U13335 (N_13335,N_6432,N_5642);
nor U13336 (N_13336,N_6058,N_6090);
xor U13337 (N_13337,N_9754,N_9842);
or U13338 (N_13338,N_7104,N_9292);
nand U13339 (N_13339,N_8457,N_5350);
and U13340 (N_13340,N_7565,N_5476);
and U13341 (N_13341,N_9765,N_9961);
nand U13342 (N_13342,N_6293,N_8620);
nand U13343 (N_13343,N_6526,N_6092);
xor U13344 (N_13344,N_6220,N_8827);
or U13345 (N_13345,N_9183,N_5279);
and U13346 (N_13346,N_9256,N_9500);
nand U13347 (N_13347,N_9959,N_7977);
nor U13348 (N_13348,N_6588,N_8236);
nor U13349 (N_13349,N_5735,N_6039);
or U13350 (N_13350,N_5880,N_6991);
nand U13351 (N_13351,N_6026,N_6102);
or U13352 (N_13352,N_5572,N_8472);
and U13353 (N_13353,N_7928,N_5145);
nand U13354 (N_13354,N_8642,N_6620);
and U13355 (N_13355,N_5057,N_9863);
and U13356 (N_13356,N_8450,N_8602);
and U13357 (N_13357,N_6605,N_7801);
xor U13358 (N_13358,N_6932,N_8585);
nor U13359 (N_13359,N_5056,N_9452);
and U13360 (N_13360,N_9036,N_8261);
xnor U13361 (N_13361,N_9342,N_9626);
nand U13362 (N_13362,N_7709,N_7829);
nand U13363 (N_13363,N_9743,N_5796);
and U13364 (N_13364,N_6938,N_7396);
and U13365 (N_13365,N_6638,N_9314);
or U13366 (N_13366,N_8937,N_8453);
nor U13367 (N_13367,N_8180,N_8441);
nor U13368 (N_13368,N_7369,N_7908);
xor U13369 (N_13369,N_6636,N_5024);
xnor U13370 (N_13370,N_8597,N_8988);
or U13371 (N_13371,N_5809,N_5586);
nand U13372 (N_13372,N_5204,N_6987);
nor U13373 (N_13373,N_9980,N_5637);
or U13374 (N_13374,N_8612,N_7991);
or U13375 (N_13375,N_8000,N_5265);
and U13376 (N_13376,N_5956,N_5291);
xor U13377 (N_13377,N_5461,N_9788);
or U13378 (N_13378,N_9707,N_8958);
nand U13379 (N_13379,N_8595,N_6200);
nor U13380 (N_13380,N_5449,N_7965);
or U13381 (N_13381,N_5364,N_8764);
and U13382 (N_13382,N_8943,N_7343);
xnor U13383 (N_13383,N_5171,N_5983);
and U13384 (N_13384,N_6026,N_8799);
and U13385 (N_13385,N_7864,N_8548);
or U13386 (N_13386,N_8759,N_8177);
xnor U13387 (N_13387,N_5629,N_8895);
nor U13388 (N_13388,N_7725,N_8468);
and U13389 (N_13389,N_5635,N_9616);
nor U13390 (N_13390,N_6236,N_6128);
xor U13391 (N_13391,N_9474,N_7902);
and U13392 (N_13392,N_8982,N_8278);
nand U13393 (N_13393,N_8688,N_6053);
or U13394 (N_13394,N_5643,N_7537);
nand U13395 (N_13395,N_5169,N_6321);
nor U13396 (N_13396,N_7915,N_9026);
and U13397 (N_13397,N_6218,N_7436);
and U13398 (N_13398,N_7429,N_6874);
nor U13399 (N_13399,N_9954,N_8189);
or U13400 (N_13400,N_8579,N_6214);
and U13401 (N_13401,N_8945,N_6024);
and U13402 (N_13402,N_6044,N_9731);
and U13403 (N_13403,N_6763,N_7032);
nand U13404 (N_13404,N_7904,N_7969);
xnor U13405 (N_13405,N_7918,N_7846);
nand U13406 (N_13406,N_6805,N_9201);
or U13407 (N_13407,N_8751,N_6828);
or U13408 (N_13408,N_7256,N_9971);
xnor U13409 (N_13409,N_5879,N_6379);
or U13410 (N_13410,N_9654,N_9619);
or U13411 (N_13411,N_8293,N_6515);
xnor U13412 (N_13412,N_8488,N_6611);
xnor U13413 (N_13413,N_8279,N_9832);
nor U13414 (N_13414,N_7678,N_5251);
or U13415 (N_13415,N_9958,N_5270);
or U13416 (N_13416,N_7875,N_7917);
nor U13417 (N_13417,N_8343,N_7107);
or U13418 (N_13418,N_8351,N_9980);
or U13419 (N_13419,N_5412,N_7690);
nor U13420 (N_13420,N_5180,N_9601);
nand U13421 (N_13421,N_9015,N_7829);
xor U13422 (N_13422,N_8635,N_8501);
nand U13423 (N_13423,N_8441,N_9812);
or U13424 (N_13424,N_5790,N_8412);
nand U13425 (N_13425,N_7548,N_8908);
xor U13426 (N_13426,N_6424,N_5031);
xor U13427 (N_13427,N_6105,N_8467);
or U13428 (N_13428,N_6266,N_5404);
nand U13429 (N_13429,N_9762,N_7789);
nor U13430 (N_13430,N_9810,N_7951);
nor U13431 (N_13431,N_8789,N_7592);
or U13432 (N_13432,N_9885,N_7692);
xnor U13433 (N_13433,N_6006,N_6474);
or U13434 (N_13434,N_5991,N_8225);
or U13435 (N_13435,N_5930,N_8838);
and U13436 (N_13436,N_7830,N_5656);
nand U13437 (N_13437,N_6010,N_5990);
xor U13438 (N_13438,N_9012,N_6916);
nor U13439 (N_13439,N_5698,N_6650);
xor U13440 (N_13440,N_8119,N_5299);
xnor U13441 (N_13441,N_8558,N_6380);
and U13442 (N_13442,N_7730,N_9948);
or U13443 (N_13443,N_6867,N_5950);
nand U13444 (N_13444,N_8843,N_7769);
xnor U13445 (N_13445,N_5888,N_9594);
nor U13446 (N_13446,N_6660,N_9630);
or U13447 (N_13447,N_9566,N_7570);
or U13448 (N_13448,N_8695,N_6985);
nand U13449 (N_13449,N_9840,N_6699);
nand U13450 (N_13450,N_9759,N_5729);
nor U13451 (N_13451,N_6759,N_6483);
nand U13452 (N_13452,N_6657,N_8202);
nand U13453 (N_13453,N_9083,N_5079);
xor U13454 (N_13454,N_6371,N_8848);
xor U13455 (N_13455,N_5488,N_5143);
nor U13456 (N_13456,N_8914,N_7774);
and U13457 (N_13457,N_7956,N_9838);
or U13458 (N_13458,N_7341,N_8912);
nand U13459 (N_13459,N_6955,N_9970);
xor U13460 (N_13460,N_9105,N_6351);
nand U13461 (N_13461,N_9608,N_8688);
xor U13462 (N_13462,N_6676,N_8844);
nand U13463 (N_13463,N_9098,N_6839);
nand U13464 (N_13464,N_6988,N_9870);
or U13465 (N_13465,N_7346,N_8167);
or U13466 (N_13466,N_8117,N_7724);
nor U13467 (N_13467,N_5457,N_7607);
nor U13468 (N_13468,N_7479,N_7982);
xnor U13469 (N_13469,N_7480,N_7249);
nor U13470 (N_13470,N_9441,N_7155);
nand U13471 (N_13471,N_5030,N_6871);
nand U13472 (N_13472,N_7684,N_7382);
and U13473 (N_13473,N_7930,N_6676);
xnor U13474 (N_13474,N_7973,N_6980);
and U13475 (N_13475,N_5332,N_6345);
nor U13476 (N_13476,N_9108,N_6744);
nand U13477 (N_13477,N_5809,N_5197);
or U13478 (N_13478,N_8774,N_5893);
nand U13479 (N_13479,N_7088,N_7423);
nor U13480 (N_13480,N_7371,N_9546);
nor U13481 (N_13481,N_8285,N_6630);
nand U13482 (N_13482,N_5342,N_9798);
xnor U13483 (N_13483,N_5310,N_7349);
xnor U13484 (N_13484,N_9612,N_8719);
or U13485 (N_13485,N_7510,N_7927);
and U13486 (N_13486,N_8221,N_6506);
and U13487 (N_13487,N_5106,N_7047);
xor U13488 (N_13488,N_7224,N_8689);
nor U13489 (N_13489,N_9056,N_6267);
and U13490 (N_13490,N_9509,N_7778);
xor U13491 (N_13491,N_5924,N_8248);
and U13492 (N_13492,N_7793,N_9233);
and U13493 (N_13493,N_8386,N_6828);
and U13494 (N_13494,N_5656,N_8109);
or U13495 (N_13495,N_8986,N_8397);
nand U13496 (N_13496,N_6950,N_5175);
nor U13497 (N_13497,N_5421,N_5200);
or U13498 (N_13498,N_5443,N_6833);
nand U13499 (N_13499,N_7514,N_9568);
xnor U13500 (N_13500,N_9044,N_8227);
xnor U13501 (N_13501,N_7131,N_7934);
xor U13502 (N_13502,N_9946,N_9076);
nand U13503 (N_13503,N_6263,N_5247);
or U13504 (N_13504,N_6836,N_8067);
and U13505 (N_13505,N_6674,N_9343);
nand U13506 (N_13506,N_6937,N_9904);
xor U13507 (N_13507,N_6258,N_9732);
or U13508 (N_13508,N_6080,N_6477);
xor U13509 (N_13509,N_8937,N_7365);
xor U13510 (N_13510,N_6683,N_9354);
nand U13511 (N_13511,N_7550,N_5134);
xor U13512 (N_13512,N_8777,N_5734);
nor U13513 (N_13513,N_6161,N_7100);
nand U13514 (N_13514,N_8953,N_6173);
xnor U13515 (N_13515,N_8267,N_6127);
nor U13516 (N_13516,N_8774,N_7885);
and U13517 (N_13517,N_9836,N_9978);
and U13518 (N_13518,N_5572,N_5641);
xnor U13519 (N_13519,N_7396,N_6555);
nor U13520 (N_13520,N_7554,N_5916);
nor U13521 (N_13521,N_6061,N_5153);
nor U13522 (N_13522,N_5029,N_7023);
nor U13523 (N_13523,N_7247,N_7555);
and U13524 (N_13524,N_5221,N_6198);
nor U13525 (N_13525,N_7657,N_9681);
xor U13526 (N_13526,N_9068,N_5043);
or U13527 (N_13527,N_5008,N_8525);
xnor U13528 (N_13528,N_9788,N_9397);
nor U13529 (N_13529,N_6781,N_9608);
and U13530 (N_13530,N_8952,N_7554);
or U13531 (N_13531,N_9979,N_7648);
or U13532 (N_13532,N_5677,N_7697);
xor U13533 (N_13533,N_6935,N_7753);
nand U13534 (N_13534,N_9123,N_5552);
nand U13535 (N_13535,N_9350,N_5384);
xnor U13536 (N_13536,N_6143,N_9126);
xnor U13537 (N_13537,N_6148,N_8787);
or U13538 (N_13538,N_6800,N_7489);
nor U13539 (N_13539,N_9734,N_9599);
nor U13540 (N_13540,N_9294,N_9085);
and U13541 (N_13541,N_7482,N_9849);
nand U13542 (N_13542,N_5672,N_9192);
nor U13543 (N_13543,N_7608,N_7224);
or U13544 (N_13544,N_5494,N_9941);
or U13545 (N_13545,N_5889,N_7855);
xnor U13546 (N_13546,N_9401,N_8994);
or U13547 (N_13547,N_9072,N_6157);
or U13548 (N_13548,N_5793,N_7133);
nor U13549 (N_13549,N_5214,N_5786);
xor U13550 (N_13550,N_8639,N_5172);
nand U13551 (N_13551,N_6427,N_5186);
xnor U13552 (N_13552,N_8876,N_6269);
nor U13553 (N_13553,N_7793,N_9136);
nor U13554 (N_13554,N_9942,N_9987);
nor U13555 (N_13555,N_9277,N_6915);
or U13556 (N_13556,N_8723,N_7775);
xnor U13557 (N_13557,N_8994,N_5900);
and U13558 (N_13558,N_8848,N_8709);
nand U13559 (N_13559,N_5596,N_7860);
nor U13560 (N_13560,N_5850,N_8868);
and U13561 (N_13561,N_6714,N_5468);
or U13562 (N_13562,N_8869,N_6180);
or U13563 (N_13563,N_5482,N_8166);
nor U13564 (N_13564,N_9856,N_7126);
xor U13565 (N_13565,N_5386,N_6544);
nand U13566 (N_13566,N_7883,N_5479);
or U13567 (N_13567,N_6662,N_6413);
nor U13568 (N_13568,N_9189,N_5254);
xor U13569 (N_13569,N_5389,N_8174);
or U13570 (N_13570,N_6652,N_8399);
and U13571 (N_13571,N_9091,N_5475);
nand U13572 (N_13572,N_9180,N_8051);
and U13573 (N_13573,N_9993,N_8566);
or U13574 (N_13574,N_7792,N_5610);
nand U13575 (N_13575,N_9452,N_9051);
nand U13576 (N_13576,N_6524,N_8703);
nand U13577 (N_13577,N_9754,N_5945);
nand U13578 (N_13578,N_7355,N_5538);
nand U13579 (N_13579,N_9414,N_8585);
and U13580 (N_13580,N_7742,N_6583);
xnor U13581 (N_13581,N_6212,N_6400);
and U13582 (N_13582,N_7125,N_5411);
nor U13583 (N_13583,N_8938,N_7780);
nand U13584 (N_13584,N_6981,N_5109);
nor U13585 (N_13585,N_7214,N_5762);
or U13586 (N_13586,N_5809,N_6493);
and U13587 (N_13587,N_6375,N_8707);
nor U13588 (N_13588,N_6090,N_7975);
nor U13589 (N_13589,N_6515,N_6230);
nor U13590 (N_13590,N_5108,N_6680);
nand U13591 (N_13591,N_8020,N_8256);
xnor U13592 (N_13592,N_5709,N_9556);
or U13593 (N_13593,N_5995,N_6630);
and U13594 (N_13594,N_9653,N_6844);
xnor U13595 (N_13595,N_7665,N_7428);
nor U13596 (N_13596,N_6733,N_5310);
nor U13597 (N_13597,N_8877,N_6574);
and U13598 (N_13598,N_9975,N_6186);
or U13599 (N_13599,N_9780,N_7671);
and U13600 (N_13600,N_6108,N_8373);
xnor U13601 (N_13601,N_6301,N_6856);
or U13602 (N_13602,N_9209,N_9691);
or U13603 (N_13603,N_6696,N_8744);
xor U13604 (N_13604,N_5605,N_6285);
xnor U13605 (N_13605,N_6523,N_6088);
nand U13606 (N_13606,N_5864,N_7062);
and U13607 (N_13607,N_8295,N_5694);
nand U13608 (N_13608,N_5619,N_6633);
or U13609 (N_13609,N_9861,N_8418);
or U13610 (N_13610,N_6315,N_6574);
nand U13611 (N_13611,N_5598,N_9337);
nor U13612 (N_13612,N_5243,N_7807);
and U13613 (N_13613,N_9379,N_8787);
nand U13614 (N_13614,N_5502,N_8565);
xor U13615 (N_13615,N_8406,N_8345);
nand U13616 (N_13616,N_8263,N_6585);
nand U13617 (N_13617,N_7516,N_5030);
xnor U13618 (N_13618,N_5769,N_7791);
nor U13619 (N_13619,N_5435,N_9866);
and U13620 (N_13620,N_6593,N_5283);
nand U13621 (N_13621,N_9730,N_6030);
nand U13622 (N_13622,N_9094,N_6617);
and U13623 (N_13623,N_8235,N_7133);
nor U13624 (N_13624,N_5061,N_7920);
xnor U13625 (N_13625,N_7823,N_9737);
xor U13626 (N_13626,N_8912,N_9347);
xor U13627 (N_13627,N_5015,N_8959);
and U13628 (N_13628,N_6301,N_6945);
or U13629 (N_13629,N_8322,N_6896);
nand U13630 (N_13630,N_9361,N_8441);
and U13631 (N_13631,N_9514,N_8156);
or U13632 (N_13632,N_8873,N_6309);
nand U13633 (N_13633,N_7544,N_8480);
xor U13634 (N_13634,N_5443,N_7524);
nand U13635 (N_13635,N_8154,N_5477);
or U13636 (N_13636,N_7310,N_5148);
nor U13637 (N_13637,N_9139,N_6457);
nand U13638 (N_13638,N_8505,N_9781);
or U13639 (N_13639,N_5276,N_7939);
or U13640 (N_13640,N_9933,N_8257);
nand U13641 (N_13641,N_9813,N_7603);
xor U13642 (N_13642,N_6147,N_7191);
and U13643 (N_13643,N_5292,N_7026);
nand U13644 (N_13644,N_6969,N_9841);
xor U13645 (N_13645,N_8435,N_5860);
nor U13646 (N_13646,N_5979,N_5036);
nor U13647 (N_13647,N_7017,N_8138);
nand U13648 (N_13648,N_9509,N_6775);
xor U13649 (N_13649,N_7414,N_5485);
xnor U13650 (N_13650,N_9688,N_9553);
xor U13651 (N_13651,N_6318,N_5339);
or U13652 (N_13652,N_8087,N_5222);
and U13653 (N_13653,N_7832,N_5076);
nor U13654 (N_13654,N_5157,N_8964);
nor U13655 (N_13655,N_5609,N_5955);
nand U13656 (N_13656,N_7319,N_9247);
or U13657 (N_13657,N_6040,N_5065);
nor U13658 (N_13658,N_7249,N_7784);
nand U13659 (N_13659,N_8745,N_9854);
xnor U13660 (N_13660,N_9649,N_5313);
or U13661 (N_13661,N_9485,N_8006);
and U13662 (N_13662,N_7053,N_6359);
or U13663 (N_13663,N_6437,N_5248);
and U13664 (N_13664,N_7036,N_7830);
nand U13665 (N_13665,N_6509,N_9097);
nand U13666 (N_13666,N_5637,N_5670);
and U13667 (N_13667,N_7325,N_7318);
and U13668 (N_13668,N_7969,N_5199);
nor U13669 (N_13669,N_6223,N_9067);
or U13670 (N_13670,N_9605,N_5557);
or U13671 (N_13671,N_7468,N_6660);
nand U13672 (N_13672,N_6590,N_9946);
and U13673 (N_13673,N_7057,N_7023);
or U13674 (N_13674,N_5715,N_8239);
nand U13675 (N_13675,N_5740,N_7586);
nor U13676 (N_13676,N_6439,N_5611);
and U13677 (N_13677,N_6652,N_8822);
or U13678 (N_13678,N_5407,N_6827);
nor U13679 (N_13679,N_9802,N_7071);
or U13680 (N_13680,N_5764,N_6210);
and U13681 (N_13681,N_9603,N_6253);
or U13682 (N_13682,N_6999,N_8458);
and U13683 (N_13683,N_9468,N_7553);
nor U13684 (N_13684,N_8927,N_9698);
nand U13685 (N_13685,N_6046,N_5550);
nand U13686 (N_13686,N_8186,N_5535);
or U13687 (N_13687,N_8909,N_8360);
nor U13688 (N_13688,N_7246,N_6271);
xnor U13689 (N_13689,N_6232,N_9999);
and U13690 (N_13690,N_9480,N_7792);
nor U13691 (N_13691,N_7136,N_9943);
or U13692 (N_13692,N_7469,N_8324);
nand U13693 (N_13693,N_6005,N_6170);
or U13694 (N_13694,N_8457,N_8545);
nand U13695 (N_13695,N_7435,N_8850);
and U13696 (N_13696,N_8561,N_8726);
or U13697 (N_13697,N_5847,N_9174);
xor U13698 (N_13698,N_7101,N_8138);
nand U13699 (N_13699,N_5112,N_5511);
or U13700 (N_13700,N_8210,N_8928);
nand U13701 (N_13701,N_5382,N_5992);
nor U13702 (N_13702,N_8202,N_9953);
and U13703 (N_13703,N_6340,N_7657);
and U13704 (N_13704,N_8118,N_9058);
xnor U13705 (N_13705,N_8723,N_7101);
or U13706 (N_13706,N_7151,N_8848);
nor U13707 (N_13707,N_6192,N_6467);
and U13708 (N_13708,N_9317,N_8204);
or U13709 (N_13709,N_6378,N_5674);
nor U13710 (N_13710,N_7141,N_9582);
nand U13711 (N_13711,N_7230,N_5609);
nor U13712 (N_13712,N_7948,N_8183);
nand U13713 (N_13713,N_6384,N_6039);
or U13714 (N_13714,N_9019,N_7678);
and U13715 (N_13715,N_5579,N_9267);
nor U13716 (N_13716,N_9851,N_5573);
and U13717 (N_13717,N_7187,N_7544);
nand U13718 (N_13718,N_7283,N_7661);
and U13719 (N_13719,N_5153,N_9925);
or U13720 (N_13720,N_6978,N_6772);
and U13721 (N_13721,N_7209,N_5683);
nand U13722 (N_13722,N_8134,N_9526);
or U13723 (N_13723,N_5998,N_6716);
or U13724 (N_13724,N_6895,N_8717);
xor U13725 (N_13725,N_7646,N_6944);
nor U13726 (N_13726,N_6375,N_6950);
nand U13727 (N_13727,N_8198,N_8447);
or U13728 (N_13728,N_7292,N_7813);
and U13729 (N_13729,N_5103,N_8632);
nor U13730 (N_13730,N_5864,N_6715);
or U13731 (N_13731,N_5074,N_5967);
nor U13732 (N_13732,N_9014,N_8501);
nor U13733 (N_13733,N_7914,N_9062);
and U13734 (N_13734,N_5166,N_5856);
nand U13735 (N_13735,N_5557,N_9550);
nor U13736 (N_13736,N_8209,N_8004);
nand U13737 (N_13737,N_6089,N_5662);
nand U13738 (N_13738,N_6343,N_5468);
xnor U13739 (N_13739,N_7358,N_8155);
nor U13740 (N_13740,N_7115,N_7574);
and U13741 (N_13741,N_9557,N_6310);
and U13742 (N_13742,N_6617,N_6958);
nand U13743 (N_13743,N_6908,N_5164);
xnor U13744 (N_13744,N_8742,N_5878);
and U13745 (N_13745,N_7725,N_5595);
nand U13746 (N_13746,N_9221,N_5011);
and U13747 (N_13747,N_7131,N_5212);
xor U13748 (N_13748,N_7276,N_9886);
and U13749 (N_13749,N_5963,N_7613);
and U13750 (N_13750,N_5100,N_9714);
nand U13751 (N_13751,N_9308,N_5195);
xor U13752 (N_13752,N_8288,N_8382);
nor U13753 (N_13753,N_8961,N_6001);
nor U13754 (N_13754,N_8212,N_7371);
and U13755 (N_13755,N_6870,N_8106);
xor U13756 (N_13756,N_7210,N_8608);
or U13757 (N_13757,N_6581,N_9440);
or U13758 (N_13758,N_9595,N_5696);
xor U13759 (N_13759,N_6633,N_7211);
nor U13760 (N_13760,N_5820,N_5231);
nand U13761 (N_13761,N_6095,N_7481);
and U13762 (N_13762,N_9006,N_9403);
and U13763 (N_13763,N_5660,N_8695);
xnor U13764 (N_13764,N_8524,N_7077);
and U13765 (N_13765,N_6845,N_9819);
nand U13766 (N_13766,N_5200,N_7583);
nor U13767 (N_13767,N_5046,N_8905);
xnor U13768 (N_13768,N_7150,N_9601);
nor U13769 (N_13769,N_9531,N_6964);
or U13770 (N_13770,N_9323,N_9008);
nor U13771 (N_13771,N_9288,N_6696);
and U13772 (N_13772,N_8813,N_5440);
xor U13773 (N_13773,N_8904,N_6394);
nand U13774 (N_13774,N_5213,N_8875);
xor U13775 (N_13775,N_6293,N_8803);
and U13776 (N_13776,N_8521,N_8094);
or U13777 (N_13777,N_6151,N_7557);
and U13778 (N_13778,N_9672,N_7929);
and U13779 (N_13779,N_7723,N_7074);
xnor U13780 (N_13780,N_8645,N_7149);
xnor U13781 (N_13781,N_7799,N_7617);
or U13782 (N_13782,N_8219,N_5053);
or U13783 (N_13783,N_5120,N_7810);
xor U13784 (N_13784,N_5684,N_8395);
xor U13785 (N_13785,N_8804,N_6345);
and U13786 (N_13786,N_6985,N_9061);
and U13787 (N_13787,N_8714,N_5471);
nand U13788 (N_13788,N_5150,N_9636);
or U13789 (N_13789,N_9921,N_7949);
and U13790 (N_13790,N_9747,N_7600);
xor U13791 (N_13791,N_8095,N_5794);
and U13792 (N_13792,N_6102,N_5140);
nand U13793 (N_13793,N_6863,N_8875);
nor U13794 (N_13794,N_7945,N_8523);
nor U13795 (N_13795,N_9440,N_9547);
or U13796 (N_13796,N_5740,N_7401);
xor U13797 (N_13797,N_5110,N_7833);
nand U13798 (N_13798,N_8945,N_9833);
or U13799 (N_13799,N_6988,N_9876);
nand U13800 (N_13800,N_6071,N_6993);
and U13801 (N_13801,N_5653,N_5489);
nand U13802 (N_13802,N_7664,N_8859);
nand U13803 (N_13803,N_5923,N_6374);
xor U13804 (N_13804,N_9407,N_8574);
nand U13805 (N_13805,N_5182,N_5000);
nand U13806 (N_13806,N_8951,N_7487);
nand U13807 (N_13807,N_7062,N_7829);
or U13808 (N_13808,N_8223,N_8065);
or U13809 (N_13809,N_6156,N_8640);
nand U13810 (N_13810,N_8546,N_5853);
or U13811 (N_13811,N_7062,N_8472);
nor U13812 (N_13812,N_7157,N_6910);
or U13813 (N_13813,N_5436,N_6003);
nor U13814 (N_13814,N_9223,N_9003);
nand U13815 (N_13815,N_6023,N_7968);
nand U13816 (N_13816,N_9823,N_8817);
and U13817 (N_13817,N_9042,N_6586);
nand U13818 (N_13818,N_9854,N_5282);
nor U13819 (N_13819,N_5056,N_5418);
nor U13820 (N_13820,N_8273,N_9076);
or U13821 (N_13821,N_9296,N_7032);
nand U13822 (N_13822,N_7441,N_9865);
nor U13823 (N_13823,N_9128,N_5638);
and U13824 (N_13824,N_8605,N_5382);
or U13825 (N_13825,N_5999,N_6625);
nor U13826 (N_13826,N_6167,N_9624);
and U13827 (N_13827,N_9294,N_8694);
xnor U13828 (N_13828,N_5987,N_9736);
nand U13829 (N_13829,N_5038,N_6632);
and U13830 (N_13830,N_9602,N_5568);
nor U13831 (N_13831,N_5847,N_8538);
or U13832 (N_13832,N_6667,N_6333);
nor U13833 (N_13833,N_6681,N_9647);
or U13834 (N_13834,N_5683,N_6001);
xor U13835 (N_13835,N_9188,N_5498);
xnor U13836 (N_13836,N_7158,N_8684);
or U13837 (N_13837,N_8958,N_8739);
nor U13838 (N_13838,N_6115,N_6046);
or U13839 (N_13839,N_9851,N_6945);
xnor U13840 (N_13840,N_7011,N_7704);
nor U13841 (N_13841,N_6957,N_9552);
and U13842 (N_13842,N_7743,N_8606);
nor U13843 (N_13843,N_5432,N_8787);
or U13844 (N_13844,N_7240,N_8009);
nand U13845 (N_13845,N_9027,N_6208);
xor U13846 (N_13846,N_6389,N_5598);
or U13847 (N_13847,N_5277,N_6773);
nor U13848 (N_13848,N_9094,N_7037);
nand U13849 (N_13849,N_7616,N_6019);
nor U13850 (N_13850,N_7277,N_8871);
and U13851 (N_13851,N_9565,N_5755);
and U13852 (N_13852,N_6020,N_9765);
nand U13853 (N_13853,N_6867,N_7414);
and U13854 (N_13854,N_6250,N_7123);
or U13855 (N_13855,N_6936,N_7361);
or U13856 (N_13856,N_8938,N_8991);
nand U13857 (N_13857,N_7666,N_6054);
nor U13858 (N_13858,N_5153,N_7272);
nand U13859 (N_13859,N_6462,N_5241);
and U13860 (N_13860,N_7994,N_7692);
or U13861 (N_13861,N_5895,N_7591);
or U13862 (N_13862,N_5353,N_7289);
or U13863 (N_13863,N_9095,N_5979);
nand U13864 (N_13864,N_8332,N_6953);
and U13865 (N_13865,N_7391,N_7042);
xnor U13866 (N_13866,N_7831,N_5589);
or U13867 (N_13867,N_5112,N_9886);
xor U13868 (N_13868,N_9821,N_7977);
xor U13869 (N_13869,N_8220,N_9266);
or U13870 (N_13870,N_7152,N_5186);
and U13871 (N_13871,N_6378,N_5826);
or U13872 (N_13872,N_6260,N_9287);
or U13873 (N_13873,N_5213,N_9638);
nor U13874 (N_13874,N_8367,N_5307);
xnor U13875 (N_13875,N_5189,N_8096);
xnor U13876 (N_13876,N_5773,N_5484);
xor U13877 (N_13877,N_8133,N_8060);
or U13878 (N_13878,N_5241,N_6519);
and U13879 (N_13879,N_5895,N_9798);
nand U13880 (N_13880,N_9146,N_7457);
and U13881 (N_13881,N_9630,N_8218);
and U13882 (N_13882,N_8488,N_7899);
or U13883 (N_13883,N_9571,N_5435);
nor U13884 (N_13884,N_8628,N_7695);
xnor U13885 (N_13885,N_5321,N_7446);
xor U13886 (N_13886,N_9139,N_5870);
nand U13887 (N_13887,N_8537,N_5484);
and U13888 (N_13888,N_7444,N_6067);
nor U13889 (N_13889,N_8716,N_9508);
xnor U13890 (N_13890,N_9484,N_9128);
and U13891 (N_13891,N_7966,N_6837);
xor U13892 (N_13892,N_9377,N_6436);
or U13893 (N_13893,N_8400,N_5152);
nor U13894 (N_13894,N_5662,N_8203);
nand U13895 (N_13895,N_5467,N_8973);
and U13896 (N_13896,N_7041,N_8832);
or U13897 (N_13897,N_6218,N_7194);
xor U13898 (N_13898,N_9286,N_6221);
nand U13899 (N_13899,N_8890,N_6528);
xor U13900 (N_13900,N_7237,N_8379);
and U13901 (N_13901,N_8569,N_7922);
nor U13902 (N_13902,N_7919,N_9173);
nor U13903 (N_13903,N_8806,N_9585);
xnor U13904 (N_13904,N_5159,N_7340);
nor U13905 (N_13905,N_5142,N_8374);
nand U13906 (N_13906,N_8723,N_6528);
or U13907 (N_13907,N_8204,N_9975);
or U13908 (N_13908,N_9780,N_9408);
xor U13909 (N_13909,N_9202,N_7767);
xor U13910 (N_13910,N_5264,N_6867);
xnor U13911 (N_13911,N_8866,N_7446);
xor U13912 (N_13912,N_7553,N_7317);
nor U13913 (N_13913,N_7408,N_7951);
or U13914 (N_13914,N_7379,N_9851);
nor U13915 (N_13915,N_5526,N_8382);
nor U13916 (N_13916,N_9643,N_8696);
or U13917 (N_13917,N_5673,N_9144);
or U13918 (N_13918,N_5881,N_6261);
xor U13919 (N_13919,N_7800,N_9497);
nor U13920 (N_13920,N_6673,N_8570);
and U13921 (N_13921,N_7525,N_6481);
or U13922 (N_13922,N_9555,N_6764);
nand U13923 (N_13923,N_8193,N_7606);
and U13924 (N_13924,N_7812,N_9978);
xor U13925 (N_13925,N_8870,N_6473);
and U13926 (N_13926,N_6778,N_7221);
xnor U13927 (N_13927,N_5532,N_9328);
nand U13928 (N_13928,N_5659,N_5692);
nor U13929 (N_13929,N_7434,N_5272);
nor U13930 (N_13930,N_6266,N_7615);
nor U13931 (N_13931,N_6223,N_6863);
nor U13932 (N_13932,N_7564,N_6163);
and U13933 (N_13933,N_7099,N_9629);
and U13934 (N_13934,N_8347,N_8626);
and U13935 (N_13935,N_5059,N_9181);
and U13936 (N_13936,N_6669,N_9190);
nor U13937 (N_13937,N_9599,N_6250);
nand U13938 (N_13938,N_6400,N_5432);
xor U13939 (N_13939,N_7294,N_7112);
or U13940 (N_13940,N_5454,N_7572);
xnor U13941 (N_13941,N_7571,N_6563);
and U13942 (N_13942,N_8659,N_9892);
xor U13943 (N_13943,N_9698,N_6713);
nand U13944 (N_13944,N_6385,N_9122);
nor U13945 (N_13945,N_6216,N_9174);
and U13946 (N_13946,N_5883,N_5793);
nor U13947 (N_13947,N_6793,N_9174);
nor U13948 (N_13948,N_7157,N_7926);
or U13949 (N_13949,N_6150,N_6906);
xnor U13950 (N_13950,N_7475,N_8268);
and U13951 (N_13951,N_7586,N_6524);
or U13952 (N_13952,N_5084,N_5417);
or U13953 (N_13953,N_7715,N_6936);
or U13954 (N_13954,N_5926,N_9366);
xor U13955 (N_13955,N_9915,N_9854);
and U13956 (N_13956,N_5762,N_9240);
nand U13957 (N_13957,N_6845,N_9003);
nor U13958 (N_13958,N_5631,N_6000);
nor U13959 (N_13959,N_6636,N_5687);
xor U13960 (N_13960,N_7068,N_8875);
nor U13961 (N_13961,N_7275,N_8875);
and U13962 (N_13962,N_8001,N_5636);
nand U13963 (N_13963,N_8655,N_5850);
xor U13964 (N_13964,N_9929,N_7548);
or U13965 (N_13965,N_5832,N_9226);
and U13966 (N_13966,N_5686,N_9762);
and U13967 (N_13967,N_7684,N_5781);
nor U13968 (N_13968,N_9296,N_8986);
nand U13969 (N_13969,N_7000,N_6109);
nor U13970 (N_13970,N_9394,N_5865);
nand U13971 (N_13971,N_6505,N_6367);
and U13972 (N_13972,N_5016,N_6840);
xnor U13973 (N_13973,N_7525,N_5490);
nor U13974 (N_13974,N_6312,N_7352);
nor U13975 (N_13975,N_7133,N_7393);
or U13976 (N_13976,N_5215,N_7685);
or U13977 (N_13977,N_6786,N_5159);
nor U13978 (N_13978,N_8775,N_8346);
and U13979 (N_13979,N_9226,N_5266);
xor U13980 (N_13980,N_5175,N_6433);
nor U13981 (N_13981,N_6120,N_8043);
and U13982 (N_13982,N_5131,N_9743);
and U13983 (N_13983,N_8746,N_8443);
xor U13984 (N_13984,N_6769,N_9192);
or U13985 (N_13985,N_9920,N_9073);
and U13986 (N_13986,N_7357,N_6252);
and U13987 (N_13987,N_7207,N_8590);
and U13988 (N_13988,N_8092,N_5500);
nor U13989 (N_13989,N_5249,N_6088);
and U13990 (N_13990,N_9751,N_7555);
xor U13991 (N_13991,N_9968,N_8611);
nand U13992 (N_13992,N_6514,N_9368);
nor U13993 (N_13993,N_7719,N_6831);
or U13994 (N_13994,N_7536,N_7023);
and U13995 (N_13995,N_9514,N_7993);
and U13996 (N_13996,N_5154,N_9554);
xor U13997 (N_13997,N_5398,N_6800);
and U13998 (N_13998,N_5174,N_5722);
and U13999 (N_13999,N_6703,N_6504);
nand U14000 (N_14000,N_5050,N_8016);
xor U14001 (N_14001,N_5665,N_5563);
nand U14002 (N_14002,N_9894,N_5767);
and U14003 (N_14003,N_8907,N_8336);
and U14004 (N_14004,N_7132,N_8384);
xnor U14005 (N_14005,N_6862,N_7024);
nand U14006 (N_14006,N_7857,N_7810);
or U14007 (N_14007,N_8287,N_9941);
nor U14008 (N_14008,N_7793,N_7391);
and U14009 (N_14009,N_9527,N_5984);
xnor U14010 (N_14010,N_7682,N_8886);
or U14011 (N_14011,N_6804,N_6699);
nand U14012 (N_14012,N_9276,N_8159);
nor U14013 (N_14013,N_9395,N_7436);
and U14014 (N_14014,N_8635,N_7775);
nor U14015 (N_14015,N_5759,N_9215);
nand U14016 (N_14016,N_6129,N_7969);
xnor U14017 (N_14017,N_9183,N_5790);
nand U14018 (N_14018,N_8946,N_8820);
and U14019 (N_14019,N_9147,N_7131);
and U14020 (N_14020,N_9919,N_8426);
nand U14021 (N_14021,N_6019,N_7592);
nor U14022 (N_14022,N_8890,N_8694);
and U14023 (N_14023,N_9607,N_8837);
xor U14024 (N_14024,N_7694,N_5415);
nand U14025 (N_14025,N_5238,N_6559);
xnor U14026 (N_14026,N_8327,N_9112);
xnor U14027 (N_14027,N_5922,N_8923);
or U14028 (N_14028,N_8655,N_6126);
and U14029 (N_14029,N_7451,N_5135);
xnor U14030 (N_14030,N_7325,N_6025);
xnor U14031 (N_14031,N_5996,N_7999);
and U14032 (N_14032,N_6296,N_5362);
xor U14033 (N_14033,N_5923,N_7164);
and U14034 (N_14034,N_9818,N_5823);
xnor U14035 (N_14035,N_5881,N_7673);
xnor U14036 (N_14036,N_8650,N_9398);
or U14037 (N_14037,N_7840,N_7362);
xor U14038 (N_14038,N_7846,N_9610);
nor U14039 (N_14039,N_5433,N_6374);
nand U14040 (N_14040,N_9376,N_8298);
or U14041 (N_14041,N_7897,N_9130);
and U14042 (N_14042,N_8038,N_9309);
xnor U14043 (N_14043,N_8878,N_6965);
xnor U14044 (N_14044,N_7282,N_9127);
or U14045 (N_14045,N_9762,N_9000);
and U14046 (N_14046,N_5666,N_6111);
nand U14047 (N_14047,N_8005,N_8106);
or U14048 (N_14048,N_7072,N_6962);
xnor U14049 (N_14049,N_7842,N_6411);
nand U14050 (N_14050,N_5189,N_8050);
and U14051 (N_14051,N_6839,N_9260);
and U14052 (N_14052,N_7928,N_6224);
and U14053 (N_14053,N_8911,N_5558);
or U14054 (N_14054,N_5886,N_6406);
xor U14055 (N_14055,N_6626,N_7206);
or U14056 (N_14056,N_9164,N_7396);
or U14057 (N_14057,N_7526,N_6623);
nand U14058 (N_14058,N_5814,N_6330);
and U14059 (N_14059,N_7101,N_8423);
or U14060 (N_14060,N_5210,N_7167);
and U14061 (N_14061,N_9612,N_7944);
and U14062 (N_14062,N_7024,N_6477);
and U14063 (N_14063,N_8140,N_8023);
nand U14064 (N_14064,N_6402,N_8670);
xnor U14065 (N_14065,N_5015,N_9722);
xnor U14066 (N_14066,N_7981,N_9067);
or U14067 (N_14067,N_7704,N_7052);
and U14068 (N_14068,N_6351,N_9801);
nand U14069 (N_14069,N_5703,N_8291);
xor U14070 (N_14070,N_7337,N_9140);
xnor U14071 (N_14071,N_7202,N_5572);
or U14072 (N_14072,N_6391,N_6925);
and U14073 (N_14073,N_6830,N_7579);
nand U14074 (N_14074,N_8979,N_6485);
and U14075 (N_14075,N_8218,N_9187);
and U14076 (N_14076,N_7578,N_8493);
nor U14077 (N_14077,N_6168,N_5037);
or U14078 (N_14078,N_7060,N_7832);
nor U14079 (N_14079,N_8466,N_6969);
xor U14080 (N_14080,N_8245,N_5589);
or U14081 (N_14081,N_9035,N_9714);
xor U14082 (N_14082,N_6853,N_9703);
nand U14083 (N_14083,N_8942,N_8400);
or U14084 (N_14084,N_7025,N_7558);
nor U14085 (N_14085,N_9837,N_5988);
and U14086 (N_14086,N_8993,N_6478);
nand U14087 (N_14087,N_8222,N_8726);
nand U14088 (N_14088,N_6778,N_6056);
nand U14089 (N_14089,N_6705,N_5275);
xor U14090 (N_14090,N_6714,N_7912);
or U14091 (N_14091,N_5832,N_9214);
or U14092 (N_14092,N_9531,N_6806);
nand U14093 (N_14093,N_9317,N_5062);
and U14094 (N_14094,N_8806,N_8752);
or U14095 (N_14095,N_6549,N_9710);
nand U14096 (N_14096,N_5989,N_5332);
or U14097 (N_14097,N_6624,N_6977);
xnor U14098 (N_14098,N_9671,N_7572);
nand U14099 (N_14099,N_7451,N_6549);
or U14100 (N_14100,N_5496,N_7526);
or U14101 (N_14101,N_7671,N_6550);
nand U14102 (N_14102,N_9049,N_8594);
or U14103 (N_14103,N_6115,N_8226);
nand U14104 (N_14104,N_6369,N_9212);
and U14105 (N_14105,N_8374,N_9489);
or U14106 (N_14106,N_7556,N_9141);
xnor U14107 (N_14107,N_6260,N_5696);
xnor U14108 (N_14108,N_9254,N_9291);
and U14109 (N_14109,N_9796,N_9108);
nor U14110 (N_14110,N_5465,N_8711);
or U14111 (N_14111,N_9213,N_8592);
nor U14112 (N_14112,N_8600,N_6990);
and U14113 (N_14113,N_8057,N_6637);
and U14114 (N_14114,N_6381,N_5205);
xor U14115 (N_14115,N_8341,N_7361);
nand U14116 (N_14116,N_7240,N_6185);
and U14117 (N_14117,N_9373,N_9551);
xor U14118 (N_14118,N_9089,N_7522);
nand U14119 (N_14119,N_5003,N_8379);
nand U14120 (N_14120,N_6049,N_8859);
nor U14121 (N_14121,N_6604,N_9197);
nand U14122 (N_14122,N_6198,N_8713);
or U14123 (N_14123,N_5385,N_5319);
and U14124 (N_14124,N_7655,N_9942);
or U14125 (N_14125,N_7317,N_6380);
and U14126 (N_14126,N_9093,N_9360);
and U14127 (N_14127,N_6746,N_9064);
and U14128 (N_14128,N_9677,N_7816);
xnor U14129 (N_14129,N_9610,N_7598);
nand U14130 (N_14130,N_9703,N_5229);
xor U14131 (N_14131,N_7677,N_8390);
nor U14132 (N_14132,N_8689,N_5015);
nand U14133 (N_14133,N_5447,N_7693);
nor U14134 (N_14134,N_9912,N_9901);
or U14135 (N_14135,N_5708,N_8540);
and U14136 (N_14136,N_6366,N_7609);
and U14137 (N_14137,N_7206,N_7590);
and U14138 (N_14138,N_8705,N_7133);
xor U14139 (N_14139,N_7004,N_6772);
xnor U14140 (N_14140,N_6820,N_6810);
nor U14141 (N_14141,N_6353,N_6628);
nor U14142 (N_14142,N_9415,N_7177);
or U14143 (N_14143,N_8810,N_8287);
nand U14144 (N_14144,N_5055,N_7937);
xor U14145 (N_14145,N_6141,N_5571);
or U14146 (N_14146,N_6034,N_5751);
nand U14147 (N_14147,N_8176,N_7747);
and U14148 (N_14148,N_7069,N_6193);
nor U14149 (N_14149,N_7384,N_9586);
nor U14150 (N_14150,N_5761,N_7533);
xor U14151 (N_14151,N_7377,N_6569);
nand U14152 (N_14152,N_6691,N_9199);
nand U14153 (N_14153,N_8813,N_8132);
or U14154 (N_14154,N_9725,N_5058);
xor U14155 (N_14155,N_9477,N_6145);
xor U14156 (N_14156,N_5208,N_7999);
nor U14157 (N_14157,N_5218,N_9099);
nand U14158 (N_14158,N_7090,N_9720);
nand U14159 (N_14159,N_7258,N_6193);
nor U14160 (N_14160,N_6004,N_5357);
nand U14161 (N_14161,N_6104,N_6023);
nand U14162 (N_14162,N_8064,N_8451);
or U14163 (N_14163,N_9727,N_7587);
xor U14164 (N_14164,N_8929,N_8674);
and U14165 (N_14165,N_9051,N_8282);
nand U14166 (N_14166,N_5423,N_7310);
and U14167 (N_14167,N_7950,N_7859);
and U14168 (N_14168,N_9792,N_7416);
nand U14169 (N_14169,N_7164,N_5121);
xor U14170 (N_14170,N_7451,N_9400);
and U14171 (N_14171,N_5495,N_6636);
nand U14172 (N_14172,N_6859,N_6846);
and U14173 (N_14173,N_6623,N_8197);
and U14174 (N_14174,N_9949,N_8514);
xor U14175 (N_14175,N_7417,N_8195);
nor U14176 (N_14176,N_5984,N_5995);
xor U14177 (N_14177,N_9424,N_7876);
nand U14178 (N_14178,N_8031,N_6632);
and U14179 (N_14179,N_9767,N_6694);
xor U14180 (N_14180,N_8441,N_5773);
xor U14181 (N_14181,N_5420,N_5330);
nand U14182 (N_14182,N_5694,N_8777);
nor U14183 (N_14183,N_9224,N_9703);
or U14184 (N_14184,N_9096,N_7272);
or U14185 (N_14185,N_5567,N_7777);
and U14186 (N_14186,N_7702,N_7802);
xnor U14187 (N_14187,N_5130,N_7226);
nor U14188 (N_14188,N_7793,N_9258);
xnor U14189 (N_14189,N_8621,N_8023);
xor U14190 (N_14190,N_8900,N_6824);
nor U14191 (N_14191,N_9906,N_9164);
nand U14192 (N_14192,N_5262,N_5432);
nand U14193 (N_14193,N_6832,N_8275);
or U14194 (N_14194,N_9680,N_5971);
nor U14195 (N_14195,N_5560,N_7883);
or U14196 (N_14196,N_5239,N_8326);
nor U14197 (N_14197,N_5001,N_8421);
and U14198 (N_14198,N_9622,N_9384);
nor U14199 (N_14199,N_9686,N_9019);
nor U14200 (N_14200,N_5598,N_9303);
nor U14201 (N_14201,N_7741,N_7894);
xnor U14202 (N_14202,N_9824,N_5169);
and U14203 (N_14203,N_9544,N_6509);
xor U14204 (N_14204,N_5031,N_7354);
and U14205 (N_14205,N_7903,N_6364);
nand U14206 (N_14206,N_9512,N_9055);
xor U14207 (N_14207,N_5314,N_6521);
nand U14208 (N_14208,N_9131,N_8141);
or U14209 (N_14209,N_7808,N_5708);
or U14210 (N_14210,N_7223,N_5848);
nand U14211 (N_14211,N_6613,N_7129);
xnor U14212 (N_14212,N_6349,N_7251);
xor U14213 (N_14213,N_7312,N_9563);
xnor U14214 (N_14214,N_7858,N_7860);
and U14215 (N_14215,N_7999,N_5974);
nand U14216 (N_14216,N_6148,N_9587);
and U14217 (N_14217,N_6127,N_7044);
or U14218 (N_14218,N_7504,N_9512);
nand U14219 (N_14219,N_7888,N_6453);
nand U14220 (N_14220,N_6853,N_7300);
nor U14221 (N_14221,N_9950,N_5459);
xnor U14222 (N_14222,N_8058,N_6302);
nand U14223 (N_14223,N_7683,N_5416);
xnor U14224 (N_14224,N_7176,N_6761);
xor U14225 (N_14225,N_9972,N_7344);
or U14226 (N_14226,N_8539,N_5884);
and U14227 (N_14227,N_6689,N_8303);
xnor U14228 (N_14228,N_8513,N_8609);
nand U14229 (N_14229,N_6264,N_5211);
or U14230 (N_14230,N_5146,N_6689);
xnor U14231 (N_14231,N_7379,N_6171);
nor U14232 (N_14232,N_9760,N_9114);
or U14233 (N_14233,N_8813,N_6924);
nor U14234 (N_14234,N_9151,N_8337);
nor U14235 (N_14235,N_8334,N_6552);
xnor U14236 (N_14236,N_6390,N_5751);
or U14237 (N_14237,N_9939,N_9863);
and U14238 (N_14238,N_6454,N_9160);
xnor U14239 (N_14239,N_8508,N_7281);
nand U14240 (N_14240,N_9554,N_8343);
and U14241 (N_14241,N_6330,N_9428);
nor U14242 (N_14242,N_8606,N_7106);
or U14243 (N_14243,N_6891,N_8721);
nand U14244 (N_14244,N_6588,N_5019);
or U14245 (N_14245,N_8658,N_6813);
or U14246 (N_14246,N_8422,N_6728);
xor U14247 (N_14247,N_8814,N_6604);
nand U14248 (N_14248,N_9815,N_5505);
nor U14249 (N_14249,N_5683,N_7493);
or U14250 (N_14250,N_8536,N_8349);
nor U14251 (N_14251,N_6119,N_8592);
nor U14252 (N_14252,N_6272,N_7550);
xor U14253 (N_14253,N_7242,N_7535);
and U14254 (N_14254,N_9770,N_8614);
nand U14255 (N_14255,N_9640,N_6598);
nor U14256 (N_14256,N_7455,N_9052);
xnor U14257 (N_14257,N_5099,N_5650);
and U14258 (N_14258,N_8886,N_7705);
and U14259 (N_14259,N_9123,N_6486);
nor U14260 (N_14260,N_5683,N_6916);
or U14261 (N_14261,N_9467,N_9922);
xor U14262 (N_14262,N_7396,N_7500);
nand U14263 (N_14263,N_7292,N_9276);
nor U14264 (N_14264,N_7492,N_9551);
and U14265 (N_14265,N_7387,N_7014);
nand U14266 (N_14266,N_6374,N_5280);
xor U14267 (N_14267,N_5925,N_9051);
or U14268 (N_14268,N_8936,N_8197);
xnor U14269 (N_14269,N_5266,N_8707);
or U14270 (N_14270,N_6301,N_7940);
nand U14271 (N_14271,N_9865,N_8375);
nor U14272 (N_14272,N_5159,N_6346);
and U14273 (N_14273,N_5225,N_5922);
nand U14274 (N_14274,N_7114,N_8639);
nand U14275 (N_14275,N_7810,N_9622);
nand U14276 (N_14276,N_8362,N_5535);
or U14277 (N_14277,N_9338,N_7707);
nor U14278 (N_14278,N_6799,N_9658);
nand U14279 (N_14279,N_9701,N_6339);
nand U14280 (N_14280,N_8125,N_6306);
or U14281 (N_14281,N_8507,N_8795);
xnor U14282 (N_14282,N_7221,N_6843);
nor U14283 (N_14283,N_5736,N_5404);
or U14284 (N_14284,N_7260,N_5401);
or U14285 (N_14285,N_8265,N_5090);
nand U14286 (N_14286,N_8820,N_7438);
xnor U14287 (N_14287,N_5113,N_6560);
xor U14288 (N_14288,N_5894,N_6744);
and U14289 (N_14289,N_9404,N_7200);
or U14290 (N_14290,N_7200,N_6712);
or U14291 (N_14291,N_8922,N_7787);
nand U14292 (N_14292,N_8021,N_6040);
nor U14293 (N_14293,N_9267,N_9371);
xnor U14294 (N_14294,N_6270,N_8723);
xnor U14295 (N_14295,N_8823,N_9154);
or U14296 (N_14296,N_6641,N_5239);
nor U14297 (N_14297,N_5044,N_8942);
xnor U14298 (N_14298,N_6540,N_9612);
and U14299 (N_14299,N_6677,N_7638);
or U14300 (N_14300,N_6154,N_9956);
nand U14301 (N_14301,N_5292,N_9516);
and U14302 (N_14302,N_8219,N_7336);
xor U14303 (N_14303,N_7543,N_5286);
nor U14304 (N_14304,N_7299,N_9967);
xor U14305 (N_14305,N_5011,N_8943);
or U14306 (N_14306,N_8731,N_5532);
xor U14307 (N_14307,N_9067,N_8485);
nand U14308 (N_14308,N_8930,N_6055);
and U14309 (N_14309,N_5354,N_7776);
xnor U14310 (N_14310,N_7383,N_7949);
xnor U14311 (N_14311,N_5282,N_6189);
and U14312 (N_14312,N_6858,N_6643);
or U14313 (N_14313,N_7282,N_7391);
and U14314 (N_14314,N_8667,N_8651);
and U14315 (N_14315,N_5371,N_5696);
nand U14316 (N_14316,N_6770,N_6134);
nand U14317 (N_14317,N_6003,N_9896);
or U14318 (N_14318,N_8604,N_6198);
nand U14319 (N_14319,N_5263,N_8636);
and U14320 (N_14320,N_9463,N_7982);
or U14321 (N_14321,N_7839,N_9692);
xnor U14322 (N_14322,N_7700,N_7969);
xnor U14323 (N_14323,N_8248,N_6039);
xnor U14324 (N_14324,N_9294,N_9754);
nor U14325 (N_14325,N_6631,N_7436);
nor U14326 (N_14326,N_9068,N_7617);
and U14327 (N_14327,N_9816,N_7895);
nand U14328 (N_14328,N_5286,N_6171);
xor U14329 (N_14329,N_9226,N_8193);
nor U14330 (N_14330,N_9261,N_6375);
nor U14331 (N_14331,N_8657,N_5788);
and U14332 (N_14332,N_8574,N_8537);
nor U14333 (N_14333,N_5921,N_6516);
nor U14334 (N_14334,N_5169,N_9471);
xnor U14335 (N_14335,N_5937,N_7608);
nand U14336 (N_14336,N_8652,N_6423);
or U14337 (N_14337,N_9341,N_5421);
or U14338 (N_14338,N_5994,N_5237);
xnor U14339 (N_14339,N_8709,N_6622);
nor U14340 (N_14340,N_5988,N_9920);
nor U14341 (N_14341,N_9385,N_9910);
or U14342 (N_14342,N_6737,N_8477);
xor U14343 (N_14343,N_7101,N_9961);
xnor U14344 (N_14344,N_6155,N_6677);
and U14345 (N_14345,N_5257,N_8012);
nand U14346 (N_14346,N_5396,N_7895);
nor U14347 (N_14347,N_7293,N_7522);
and U14348 (N_14348,N_8905,N_6502);
and U14349 (N_14349,N_6563,N_5446);
and U14350 (N_14350,N_6344,N_9580);
and U14351 (N_14351,N_6133,N_5420);
nor U14352 (N_14352,N_7856,N_8501);
and U14353 (N_14353,N_6423,N_8857);
nand U14354 (N_14354,N_9736,N_7861);
or U14355 (N_14355,N_8481,N_9245);
xor U14356 (N_14356,N_5886,N_6154);
xnor U14357 (N_14357,N_7023,N_8825);
nand U14358 (N_14358,N_5483,N_5111);
xor U14359 (N_14359,N_6538,N_9399);
and U14360 (N_14360,N_9153,N_5582);
and U14361 (N_14361,N_6339,N_8184);
or U14362 (N_14362,N_6740,N_9877);
xnor U14363 (N_14363,N_8936,N_9288);
nor U14364 (N_14364,N_9807,N_5357);
xnor U14365 (N_14365,N_8900,N_7572);
or U14366 (N_14366,N_5309,N_6307);
or U14367 (N_14367,N_5150,N_6341);
nand U14368 (N_14368,N_8693,N_9846);
or U14369 (N_14369,N_6732,N_7667);
nand U14370 (N_14370,N_7907,N_5237);
and U14371 (N_14371,N_5088,N_8866);
or U14372 (N_14372,N_7052,N_5170);
or U14373 (N_14373,N_6460,N_5600);
nor U14374 (N_14374,N_8337,N_5741);
nor U14375 (N_14375,N_6085,N_8848);
or U14376 (N_14376,N_7730,N_5091);
and U14377 (N_14377,N_7807,N_9259);
xor U14378 (N_14378,N_8315,N_8600);
xor U14379 (N_14379,N_6430,N_7446);
nor U14380 (N_14380,N_7335,N_7922);
or U14381 (N_14381,N_8709,N_7985);
and U14382 (N_14382,N_6445,N_6810);
and U14383 (N_14383,N_5023,N_9890);
and U14384 (N_14384,N_9955,N_6164);
nor U14385 (N_14385,N_7508,N_9497);
and U14386 (N_14386,N_7557,N_7889);
nand U14387 (N_14387,N_6096,N_7928);
nand U14388 (N_14388,N_9374,N_8964);
xor U14389 (N_14389,N_6258,N_6606);
nor U14390 (N_14390,N_6158,N_6676);
nand U14391 (N_14391,N_7587,N_8955);
nor U14392 (N_14392,N_6483,N_9242);
or U14393 (N_14393,N_5810,N_5067);
nor U14394 (N_14394,N_8963,N_6561);
nand U14395 (N_14395,N_9354,N_5257);
and U14396 (N_14396,N_9385,N_9181);
nor U14397 (N_14397,N_7519,N_7523);
nor U14398 (N_14398,N_9191,N_9482);
nor U14399 (N_14399,N_5931,N_5383);
nand U14400 (N_14400,N_5084,N_7852);
xor U14401 (N_14401,N_8810,N_7748);
and U14402 (N_14402,N_6692,N_6913);
xnor U14403 (N_14403,N_7242,N_6924);
and U14404 (N_14404,N_6554,N_6663);
or U14405 (N_14405,N_5226,N_5135);
nand U14406 (N_14406,N_8262,N_8503);
and U14407 (N_14407,N_6933,N_8206);
nor U14408 (N_14408,N_6898,N_8451);
or U14409 (N_14409,N_9661,N_6007);
nand U14410 (N_14410,N_6544,N_8846);
nor U14411 (N_14411,N_9568,N_6344);
or U14412 (N_14412,N_7252,N_9206);
nor U14413 (N_14413,N_6234,N_7789);
and U14414 (N_14414,N_7656,N_8974);
nand U14415 (N_14415,N_8859,N_5877);
nor U14416 (N_14416,N_8595,N_9609);
and U14417 (N_14417,N_8587,N_6421);
nand U14418 (N_14418,N_6095,N_7415);
and U14419 (N_14419,N_7442,N_9913);
or U14420 (N_14420,N_5959,N_5130);
and U14421 (N_14421,N_9914,N_9458);
or U14422 (N_14422,N_7726,N_7037);
and U14423 (N_14423,N_8235,N_8966);
xor U14424 (N_14424,N_7146,N_9716);
nand U14425 (N_14425,N_6651,N_9780);
xnor U14426 (N_14426,N_6677,N_5482);
or U14427 (N_14427,N_6251,N_8501);
nor U14428 (N_14428,N_5983,N_6080);
nand U14429 (N_14429,N_7834,N_8407);
or U14430 (N_14430,N_9130,N_9872);
or U14431 (N_14431,N_5626,N_9272);
or U14432 (N_14432,N_6845,N_5106);
nand U14433 (N_14433,N_9233,N_7084);
or U14434 (N_14434,N_9652,N_7447);
xnor U14435 (N_14435,N_8492,N_8868);
or U14436 (N_14436,N_9990,N_9708);
nand U14437 (N_14437,N_5738,N_9913);
or U14438 (N_14438,N_7568,N_8662);
or U14439 (N_14439,N_9311,N_5459);
and U14440 (N_14440,N_8324,N_7492);
or U14441 (N_14441,N_7970,N_5392);
xor U14442 (N_14442,N_8035,N_7243);
xor U14443 (N_14443,N_7585,N_5495);
nor U14444 (N_14444,N_9228,N_6481);
nand U14445 (N_14445,N_7428,N_5924);
or U14446 (N_14446,N_6299,N_5280);
nor U14447 (N_14447,N_7501,N_7046);
xnor U14448 (N_14448,N_5355,N_5767);
and U14449 (N_14449,N_5587,N_7273);
nand U14450 (N_14450,N_8494,N_5429);
xor U14451 (N_14451,N_8626,N_5296);
and U14452 (N_14452,N_8514,N_5411);
xnor U14453 (N_14453,N_8524,N_7365);
nand U14454 (N_14454,N_7807,N_7980);
xor U14455 (N_14455,N_7093,N_5675);
xor U14456 (N_14456,N_7227,N_7543);
nand U14457 (N_14457,N_6534,N_9114);
nand U14458 (N_14458,N_7733,N_7646);
and U14459 (N_14459,N_5507,N_6790);
xnor U14460 (N_14460,N_9964,N_5956);
nor U14461 (N_14461,N_9586,N_5710);
and U14462 (N_14462,N_7084,N_8078);
or U14463 (N_14463,N_9273,N_5591);
and U14464 (N_14464,N_8073,N_9439);
and U14465 (N_14465,N_7290,N_8139);
and U14466 (N_14466,N_6884,N_6735);
nor U14467 (N_14467,N_7235,N_8044);
and U14468 (N_14468,N_5699,N_8120);
xnor U14469 (N_14469,N_9245,N_7766);
nand U14470 (N_14470,N_9353,N_5045);
nor U14471 (N_14471,N_5970,N_5500);
nand U14472 (N_14472,N_5250,N_7724);
nand U14473 (N_14473,N_8579,N_9966);
and U14474 (N_14474,N_7360,N_9248);
or U14475 (N_14475,N_7321,N_8977);
xnor U14476 (N_14476,N_9203,N_8064);
and U14477 (N_14477,N_6787,N_9298);
nand U14478 (N_14478,N_7093,N_6236);
nand U14479 (N_14479,N_5662,N_7893);
xor U14480 (N_14480,N_6431,N_5593);
nor U14481 (N_14481,N_7356,N_8837);
nand U14482 (N_14482,N_6225,N_8991);
or U14483 (N_14483,N_6260,N_7545);
and U14484 (N_14484,N_9111,N_7761);
xnor U14485 (N_14485,N_7106,N_8536);
nor U14486 (N_14486,N_8999,N_9783);
xnor U14487 (N_14487,N_9881,N_9034);
or U14488 (N_14488,N_8207,N_9076);
nand U14489 (N_14489,N_7822,N_9182);
nor U14490 (N_14490,N_5174,N_9385);
nand U14491 (N_14491,N_8141,N_6748);
and U14492 (N_14492,N_9904,N_8451);
and U14493 (N_14493,N_5076,N_6409);
and U14494 (N_14494,N_6795,N_6868);
and U14495 (N_14495,N_9706,N_6968);
and U14496 (N_14496,N_9008,N_5431);
and U14497 (N_14497,N_8558,N_6567);
nor U14498 (N_14498,N_6100,N_9962);
and U14499 (N_14499,N_5226,N_7018);
nand U14500 (N_14500,N_5016,N_8593);
or U14501 (N_14501,N_6606,N_9996);
xnor U14502 (N_14502,N_8171,N_8446);
nand U14503 (N_14503,N_7494,N_9929);
nor U14504 (N_14504,N_5583,N_5290);
or U14505 (N_14505,N_7008,N_5339);
nor U14506 (N_14506,N_7918,N_5857);
xnor U14507 (N_14507,N_9205,N_6809);
xnor U14508 (N_14508,N_5326,N_8332);
xor U14509 (N_14509,N_8318,N_7536);
nor U14510 (N_14510,N_7541,N_6659);
xnor U14511 (N_14511,N_6245,N_9288);
and U14512 (N_14512,N_8819,N_8162);
xor U14513 (N_14513,N_6449,N_9817);
nor U14514 (N_14514,N_6443,N_8471);
xor U14515 (N_14515,N_7473,N_6956);
nor U14516 (N_14516,N_6795,N_5463);
or U14517 (N_14517,N_7925,N_6175);
xnor U14518 (N_14518,N_6508,N_8184);
nor U14519 (N_14519,N_5043,N_5459);
or U14520 (N_14520,N_8504,N_6530);
xor U14521 (N_14521,N_6071,N_8494);
and U14522 (N_14522,N_6926,N_7323);
and U14523 (N_14523,N_9090,N_9167);
nor U14524 (N_14524,N_7202,N_7412);
xor U14525 (N_14525,N_8965,N_7083);
and U14526 (N_14526,N_6310,N_8558);
nor U14527 (N_14527,N_9975,N_6013);
or U14528 (N_14528,N_6321,N_5666);
xor U14529 (N_14529,N_8421,N_6705);
nand U14530 (N_14530,N_8475,N_9529);
nand U14531 (N_14531,N_9315,N_8353);
and U14532 (N_14532,N_8508,N_9147);
and U14533 (N_14533,N_7191,N_6779);
or U14534 (N_14534,N_5460,N_9736);
or U14535 (N_14535,N_8080,N_7676);
nor U14536 (N_14536,N_8696,N_7648);
nand U14537 (N_14537,N_6026,N_9290);
nand U14538 (N_14538,N_6973,N_6172);
and U14539 (N_14539,N_7828,N_8537);
nand U14540 (N_14540,N_5713,N_5648);
or U14541 (N_14541,N_8077,N_9170);
nand U14542 (N_14542,N_8474,N_5157);
and U14543 (N_14543,N_5509,N_8486);
and U14544 (N_14544,N_9811,N_8633);
or U14545 (N_14545,N_7404,N_5347);
nand U14546 (N_14546,N_9013,N_6896);
or U14547 (N_14547,N_6541,N_5751);
nand U14548 (N_14548,N_7353,N_8294);
nand U14549 (N_14549,N_6595,N_9489);
xor U14550 (N_14550,N_8299,N_9408);
nor U14551 (N_14551,N_9014,N_6878);
and U14552 (N_14552,N_8969,N_6338);
xnor U14553 (N_14553,N_5993,N_9229);
nand U14554 (N_14554,N_7049,N_8417);
xor U14555 (N_14555,N_7521,N_6587);
nor U14556 (N_14556,N_9361,N_8861);
nand U14557 (N_14557,N_5532,N_9212);
nand U14558 (N_14558,N_9054,N_5498);
nor U14559 (N_14559,N_7610,N_7996);
and U14560 (N_14560,N_6122,N_9264);
and U14561 (N_14561,N_6737,N_6213);
xor U14562 (N_14562,N_6116,N_9862);
or U14563 (N_14563,N_5345,N_6628);
nor U14564 (N_14564,N_9960,N_5073);
xor U14565 (N_14565,N_6132,N_8684);
xor U14566 (N_14566,N_7843,N_5484);
nor U14567 (N_14567,N_6641,N_7313);
nand U14568 (N_14568,N_7698,N_7561);
nor U14569 (N_14569,N_8404,N_7299);
nand U14570 (N_14570,N_5758,N_7907);
and U14571 (N_14571,N_7213,N_5370);
and U14572 (N_14572,N_9055,N_7273);
nand U14573 (N_14573,N_5035,N_7833);
xnor U14574 (N_14574,N_5021,N_7599);
and U14575 (N_14575,N_9498,N_8256);
nor U14576 (N_14576,N_8844,N_9287);
or U14577 (N_14577,N_6064,N_6543);
nand U14578 (N_14578,N_6086,N_7404);
nor U14579 (N_14579,N_8041,N_5515);
or U14580 (N_14580,N_7041,N_6649);
nand U14581 (N_14581,N_7887,N_6640);
xor U14582 (N_14582,N_5470,N_8168);
nor U14583 (N_14583,N_7512,N_5043);
or U14584 (N_14584,N_8455,N_7414);
nand U14585 (N_14585,N_7586,N_8314);
or U14586 (N_14586,N_5347,N_5889);
or U14587 (N_14587,N_6068,N_6883);
nor U14588 (N_14588,N_9053,N_9441);
and U14589 (N_14589,N_8538,N_6382);
nor U14590 (N_14590,N_8768,N_8198);
or U14591 (N_14591,N_6973,N_5197);
and U14592 (N_14592,N_7447,N_5604);
nor U14593 (N_14593,N_5842,N_5987);
xor U14594 (N_14594,N_5909,N_6692);
nand U14595 (N_14595,N_8049,N_5684);
or U14596 (N_14596,N_8735,N_9690);
nand U14597 (N_14597,N_6009,N_5165);
xor U14598 (N_14598,N_5150,N_9726);
and U14599 (N_14599,N_8199,N_5434);
nor U14600 (N_14600,N_6165,N_7381);
xnor U14601 (N_14601,N_9382,N_9720);
and U14602 (N_14602,N_8426,N_7809);
xor U14603 (N_14603,N_8733,N_5279);
and U14604 (N_14604,N_9589,N_6058);
nand U14605 (N_14605,N_8956,N_9144);
or U14606 (N_14606,N_6908,N_9822);
and U14607 (N_14607,N_9540,N_6059);
and U14608 (N_14608,N_6608,N_9917);
and U14609 (N_14609,N_8040,N_5462);
nor U14610 (N_14610,N_8177,N_7647);
nor U14611 (N_14611,N_6507,N_6122);
nor U14612 (N_14612,N_7390,N_7694);
or U14613 (N_14613,N_9387,N_7668);
nor U14614 (N_14614,N_5300,N_6917);
nor U14615 (N_14615,N_5934,N_9276);
nand U14616 (N_14616,N_5911,N_8812);
nand U14617 (N_14617,N_6640,N_9519);
xor U14618 (N_14618,N_7950,N_7341);
nand U14619 (N_14619,N_9924,N_5212);
and U14620 (N_14620,N_8423,N_6748);
and U14621 (N_14621,N_7850,N_5178);
and U14622 (N_14622,N_7714,N_7318);
nand U14623 (N_14623,N_5436,N_6597);
nor U14624 (N_14624,N_8668,N_6067);
nor U14625 (N_14625,N_8782,N_6633);
nand U14626 (N_14626,N_6231,N_6631);
nor U14627 (N_14627,N_5404,N_9679);
and U14628 (N_14628,N_9155,N_9686);
or U14629 (N_14629,N_6937,N_5781);
and U14630 (N_14630,N_9322,N_7168);
nand U14631 (N_14631,N_7500,N_5826);
xor U14632 (N_14632,N_7321,N_8306);
and U14633 (N_14633,N_7385,N_8505);
nand U14634 (N_14634,N_7284,N_6908);
and U14635 (N_14635,N_6509,N_9827);
and U14636 (N_14636,N_7047,N_7179);
xor U14637 (N_14637,N_5641,N_8785);
xnor U14638 (N_14638,N_8989,N_8289);
xor U14639 (N_14639,N_6805,N_5205);
and U14640 (N_14640,N_6389,N_6041);
or U14641 (N_14641,N_6231,N_6263);
or U14642 (N_14642,N_9443,N_8610);
xor U14643 (N_14643,N_5387,N_5826);
or U14644 (N_14644,N_8412,N_9732);
nand U14645 (N_14645,N_9315,N_9916);
xnor U14646 (N_14646,N_8404,N_6123);
or U14647 (N_14647,N_5712,N_7690);
xor U14648 (N_14648,N_7622,N_8723);
or U14649 (N_14649,N_5422,N_5633);
and U14650 (N_14650,N_5530,N_8363);
xor U14651 (N_14651,N_8543,N_5098);
xor U14652 (N_14652,N_8568,N_5091);
nor U14653 (N_14653,N_5517,N_8105);
xnor U14654 (N_14654,N_6750,N_9191);
xor U14655 (N_14655,N_7059,N_5164);
xor U14656 (N_14656,N_8925,N_6638);
nor U14657 (N_14657,N_8044,N_8662);
xor U14658 (N_14658,N_8930,N_7262);
nor U14659 (N_14659,N_9873,N_9680);
nor U14660 (N_14660,N_6516,N_8103);
and U14661 (N_14661,N_9218,N_8493);
nand U14662 (N_14662,N_9981,N_9989);
nand U14663 (N_14663,N_6786,N_7007);
nand U14664 (N_14664,N_9301,N_9355);
xnor U14665 (N_14665,N_5897,N_6736);
or U14666 (N_14666,N_6801,N_7153);
nand U14667 (N_14667,N_9107,N_7758);
nor U14668 (N_14668,N_5921,N_5502);
or U14669 (N_14669,N_8571,N_9069);
and U14670 (N_14670,N_5521,N_5725);
and U14671 (N_14671,N_5534,N_5246);
xor U14672 (N_14672,N_5814,N_9948);
nor U14673 (N_14673,N_5078,N_9974);
and U14674 (N_14674,N_9370,N_6148);
and U14675 (N_14675,N_7356,N_6818);
and U14676 (N_14676,N_5413,N_8012);
nand U14677 (N_14677,N_8328,N_9170);
and U14678 (N_14678,N_6907,N_7850);
or U14679 (N_14679,N_8743,N_5255);
or U14680 (N_14680,N_8171,N_6909);
or U14681 (N_14681,N_8396,N_6905);
xnor U14682 (N_14682,N_5558,N_6015);
or U14683 (N_14683,N_7492,N_7927);
and U14684 (N_14684,N_6519,N_8377);
nor U14685 (N_14685,N_8139,N_5211);
nor U14686 (N_14686,N_6917,N_8998);
xor U14687 (N_14687,N_6348,N_6586);
nor U14688 (N_14688,N_5578,N_9964);
and U14689 (N_14689,N_8510,N_5280);
and U14690 (N_14690,N_6983,N_7279);
xor U14691 (N_14691,N_8526,N_5262);
or U14692 (N_14692,N_9361,N_6512);
nand U14693 (N_14693,N_5692,N_8328);
nor U14694 (N_14694,N_8591,N_7905);
nor U14695 (N_14695,N_6001,N_7452);
or U14696 (N_14696,N_9963,N_8857);
and U14697 (N_14697,N_8006,N_8353);
or U14698 (N_14698,N_8841,N_6719);
nand U14699 (N_14699,N_9520,N_7770);
nand U14700 (N_14700,N_7386,N_9466);
xnor U14701 (N_14701,N_8535,N_6607);
or U14702 (N_14702,N_6783,N_9202);
xnor U14703 (N_14703,N_8691,N_9837);
xnor U14704 (N_14704,N_9429,N_8647);
nand U14705 (N_14705,N_9955,N_8090);
xor U14706 (N_14706,N_6186,N_5225);
and U14707 (N_14707,N_5898,N_8839);
and U14708 (N_14708,N_5526,N_8333);
or U14709 (N_14709,N_9831,N_5774);
and U14710 (N_14710,N_6491,N_5656);
and U14711 (N_14711,N_7845,N_5983);
and U14712 (N_14712,N_7786,N_5506);
and U14713 (N_14713,N_5649,N_7868);
and U14714 (N_14714,N_9751,N_7046);
nor U14715 (N_14715,N_5467,N_6143);
nor U14716 (N_14716,N_9659,N_6194);
or U14717 (N_14717,N_8359,N_7343);
and U14718 (N_14718,N_7687,N_9673);
or U14719 (N_14719,N_6758,N_9982);
xnor U14720 (N_14720,N_6843,N_5867);
nand U14721 (N_14721,N_6328,N_6138);
or U14722 (N_14722,N_7375,N_5612);
and U14723 (N_14723,N_9831,N_9298);
or U14724 (N_14724,N_8748,N_8744);
nand U14725 (N_14725,N_5981,N_9682);
nand U14726 (N_14726,N_6586,N_9574);
and U14727 (N_14727,N_5369,N_8127);
xor U14728 (N_14728,N_9870,N_9565);
or U14729 (N_14729,N_7379,N_9030);
or U14730 (N_14730,N_6525,N_6130);
xnor U14731 (N_14731,N_5418,N_8576);
and U14732 (N_14732,N_6365,N_8319);
xor U14733 (N_14733,N_6850,N_6174);
and U14734 (N_14734,N_5622,N_5831);
nor U14735 (N_14735,N_8418,N_6906);
or U14736 (N_14736,N_8513,N_6613);
nor U14737 (N_14737,N_5794,N_8622);
nand U14738 (N_14738,N_9977,N_9928);
nand U14739 (N_14739,N_7080,N_9783);
xor U14740 (N_14740,N_8101,N_6700);
nor U14741 (N_14741,N_7766,N_7110);
and U14742 (N_14742,N_8520,N_8073);
xnor U14743 (N_14743,N_8805,N_6980);
nand U14744 (N_14744,N_5675,N_9957);
and U14745 (N_14745,N_8486,N_9995);
and U14746 (N_14746,N_5203,N_9298);
nor U14747 (N_14747,N_9145,N_9271);
or U14748 (N_14748,N_6763,N_8024);
nor U14749 (N_14749,N_7870,N_7424);
nor U14750 (N_14750,N_5908,N_6861);
xnor U14751 (N_14751,N_5752,N_7834);
nand U14752 (N_14752,N_5411,N_7462);
nand U14753 (N_14753,N_6391,N_9893);
xnor U14754 (N_14754,N_7771,N_6551);
or U14755 (N_14755,N_7465,N_9330);
and U14756 (N_14756,N_6138,N_5202);
nand U14757 (N_14757,N_5167,N_8505);
nor U14758 (N_14758,N_5949,N_8155);
or U14759 (N_14759,N_6190,N_5781);
and U14760 (N_14760,N_5887,N_5114);
or U14761 (N_14761,N_6418,N_6697);
or U14762 (N_14762,N_6559,N_8244);
or U14763 (N_14763,N_5568,N_6140);
or U14764 (N_14764,N_6483,N_8941);
nand U14765 (N_14765,N_9522,N_5581);
xor U14766 (N_14766,N_5559,N_6676);
and U14767 (N_14767,N_6257,N_6331);
xnor U14768 (N_14768,N_6368,N_7013);
or U14769 (N_14769,N_5642,N_5702);
nor U14770 (N_14770,N_9941,N_8503);
and U14771 (N_14771,N_7337,N_6410);
or U14772 (N_14772,N_7081,N_9185);
and U14773 (N_14773,N_8355,N_8859);
and U14774 (N_14774,N_6745,N_9522);
and U14775 (N_14775,N_9082,N_9191);
and U14776 (N_14776,N_7802,N_6020);
or U14777 (N_14777,N_7955,N_8389);
and U14778 (N_14778,N_7652,N_9046);
nand U14779 (N_14779,N_6602,N_7247);
or U14780 (N_14780,N_6894,N_6083);
xnor U14781 (N_14781,N_8021,N_5449);
nand U14782 (N_14782,N_5123,N_7511);
or U14783 (N_14783,N_5251,N_9143);
or U14784 (N_14784,N_6191,N_9029);
nor U14785 (N_14785,N_5814,N_8418);
nor U14786 (N_14786,N_6542,N_5574);
and U14787 (N_14787,N_7832,N_9651);
xor U14788 (N_14788,N_9497,N_7806);
nor U14789 (N_14789,N_6913,N_6187);
xor U14790 (N_14790,N_7664,N_5462);
xor U14791 (N_14791,N_6316,N_9116);
and U14792 (N_14792,N_9047,N_6923);
nand U14793 (N_14793,N_9200,N_7944);
nor U14794 (N_14794,N_9683,N_8818);
nor U14795 (N_14795,N_5348,N_5867);
xor U14796 (N_14796,N_8561,N_7923);
or U14797 (N_14797,N_8769,N_7334);
or U14798 (N_14798,N_7613,N_8814);
xor U14799 (N_14799,N_7520,N_9022);
nand U14800 (N_14800,N_7901,N_9435);
nand U14801 (N_14801,N_6319,N_7845);
nand U14802 (N_14802,N_5393,N_8898);
nor U14803 (N_14803,N_8881,N_9749);
or U14804 (N_14804,N_7030,N_7369);
or U14805 (N_14805,N_7530,N_7642);
nand U14806 (N_14806,N_8626,N_7535);
or U14807 (N_14807,N_6252,N_6391);
xnor U14808 (N_14808,N_8893,N_9738);
and U14809 (N_14809,N_9216,N_9751);
xor U14810 (N_14810,N_5016,N_5319);
nor U14811 (N_14811,N_8853,N_9937);
nor U14812 (N_14812,N_6551,N_5834);
nor U14813 (N_14813,N_5296,N_8005);
nand U14814 (N_14814,N_6783,N_9458);
xor U14815 (N_14815,N_7524,N_5685);
xor U14816 (N_14816,N_5889,N_8326);
nand U14817 (N_14817,N_7176,N_9839);
nor U14818 (N_14818,N_9020,N_9482);
nand U14819 (N_14819,N_8998,N_5255);
nor U14820 (N_14820,N_6976,N_7079);
nand U14821 (N_14821,N_9733,N_5421);
xnor U14822 (N_14822,N_6048,N_7727);
nand U14823 (N_14823,N_5578,N_8341);
xor U14824 (N_14824,N_7236,N_6824);
nand U14825 (N_14825,N_8454,N_7618);
xor U14826 (N_14826,N_8932,N_9940);
nor U14827 (N_14827,N_5743,N_5876);
and U14828 (N_14828,N_6380,N_7464);
xnor U14829 (N_14829,N_5320,N_5574);
nor U14830 (N_14830,N_9159,N_8652);
nand U14831 (N_14831,N_7582,N_6803);
or U14832 (N_14832,N_9169,N_5639);
nor U14833 (N_14833,N_9894,N_6405);
nor U14834 (N_14834,N_5646,N_6591);
nand U14835 (N_14835,N_7960,N_7938);
or U14836 (N_14836,N_5090,N_5082);
or U14837 (N_14837,N_5528,N_7383);
or U14838 (N_14838,N_8439,N_6917);
xor U14839 (N_14839,N_7291,N_9319);
and U14840 (N_14840,N_7047,N_5193);
and U14841 (N_14841,N_5275,N_8690);
nor U14842 (N_14842,N_5255,N_9179);
and U14843 (N_14843,N_8320,N_6304);
or U14844 (N_14844,N_7651,N_9780);
nor U14845 (N_14845,N_5559,N_8380);
or U14846 (N_14846,N_9113,N_6805);
or U14847 (N_14847,N_5752,N_6439);
nor U14848 (N_14848,N_7483,N_9079);
nand U14849 (N_14849,N_5878,N_7574);
or U14850 (N_14850,N_9275,N_7580);
nand U14851 (N_14851,N_7720,N_6162);
or U14852 (N_14852,N_8290,N_7522);
or U14853 (N_14853,N_8597,N_9367);
nand U14854 (N_14854,N_6211,N_5738);
nand U14855 (N_14855,N_7791,N_9712);
xnor U14856 (N_14856,N_7820,N_9299);
nor U14857 (N_14857,N_6962,N_7533);
and U14858 (N_14858,N_6318,N_6688);
or U14859 (N_14859,N_7590,N_6422);
or U14860 (N_14860,N_7705,N_6797);
and U14861 (N_14861,N_5545,N_9774);
or U14862 (N_14862,N_5678,N_5791);
nand U14863 (N_14863,N_8984,N_9514);
nor U14864 (N_14864,N_8983,N_8795);
nand U14865 (N_14865,N_5128,N_7547);
or U14866 (N_14866,N_6727,N_5392);
nand U14867 (N_14867,N_7475,N_5155);
xnor U14868 (N_14868,N_7871,N_8348);
nor U14869 (N_14869,N_5742,N_6331);
xnor U14870 (N_14870,N_6702,N_8192);
and U14871 (N_14871,N_9180,N_8062);
nor U14872 (N_14872,N_5475,N_6974);
nand U14873 (N_14873,N_6928,N_5274);
and U14874 (N_14874,N_9196,N_9620);
or U14875 (N_14875,N_7857,N_6158);
xnor U14876 (N_14876,N_7330,N_6478);
nor U14877 (N_14877,N_9630,N_6800);
and U14878 (N_14878,N_5600,N_8124);
nor U14879 (N_14879,N_8566,N_5313);
and U14880 (N_14880,N_5812,N_6170);
and U14881 (N_14881,N_9297,N_5422);
or U14882 (N_14882,N_6298,N_9898);
nor U14883 (N_14883,N_9189,N_7206);
and U14884 (N_14884,N_8220,N_5531);
xor U14885 (N_14885,N_6666,N_7891);
nand U14886 (N_14886,N_7044,N_5038);
and U14887 (N_14887,N_5387,N_6630);
or U14888 (N_14888,N_8182,N_9352);
nor U14889 (N_14889,N_9552,N_5409);
or U14890 (N_14890,N_6450,N_7484);
or U14891 (N_14891,N_9270,N_6851);
and U14892 (N_14892,N_5853,N_8498);
xnor U14893 (N_14893,N_8683,N_9073);
nor U14894 (N_14894,N_8015,N_5815);
and U14895 (N_14895,N_5442,N_5011);
nand U14896 (N_14896,N_9012,N_5574);
or U14897 (N_14897,N_5823,N_8188);
xnor U14898 (N_14898,N_5343,N_6015);
or U14899 (N_14899,N_9737,N_8376);
and U14900 (N_14900,N_7833,N_9480);
and U14901 (N_14901,N_7851,N_9470);
and U14902 (N_14902,N_6712,N_6055);
nor U14903 (N_14903,N_5840,N_9518);
or U14904 (N_14904,N_8519,N_6010);
or U14905 (N_14905,N_9647,N_8506);
or U14906 (N_14906,N_7282,N_5643);
nand U14907 (N_14907,N_7476,N_8177);
and U14908 (N_14908,N_9923,N_9755);
or U14909 (N_14909,N_6817,N_7548);
nand U14910 (N_14910,N_8715,N_5191);
and U14911 (N_14911,N_7154,N_6443);
and U14912 (N_14912,N_8590,N_7236);
and U14913 (N_14913,N_7050,N_5682);
or U14914 (N_14914,N_6617,N_7216);
and U14915 (N_14915,N_6778,N_9719);
xor U14916 (N_14916,N_8900,N_7306);
nor U14917 (N_14917,N_5941,N_8729);
xnor U14918 (N_14918,N_7776,N_7156);
nor U14919 (N_14919,N_9442,N_7421);
xor U14920 (N_14920,N_9479,N_7647);
nor U14921 (N_14921,N_5633,N_7506);
or U14922 (N_14922,N_8572,N_9869);
xnor U14923 (N_14923,N_9967,N_8329);
xnor U14924 (N_14924,N_8963,N_6922);
nand U14925 (N_14925,N_9389,N_9923);
and U14926 (N_14926,N_8297,N_5884);
xor U14927 (N_14927,N_6836,N_9747);
nand U14928 (N_14928,N_8548,N_7098);
and U14929 (N_14929,N_8469,N_6641);
nand U14930 (N_14930,N_5263,N_6148);
nand U14931 (N_14931,N_6618,N_8846);
nand U14932 (N_14932,N_7885,N_7312);
or U14933 (N_14933,N_5354,N_7764);
and U14934 (N_14934,N_7954,N_9078);
and U14935 (N_14935,N_9138,N_7740);
xor U14936 (N_14936,N_9117,N_9792);
nand U14937 (N_14937,N_7362,N_6110);
nand U14938 (N_14938,N_6050,N_6098);
xor U14939 (N_14939,N_9313,N_8827);
nand U14940 (N_14940,N_7819,N_6640);
or U14941 (N_14941,N_8897,N_8167);
and U14942 (N_14942,N_7132,N_9837);
nor U14943 (N_14943,N_5556,N_8412);
and U14944 (N_14944,N_6016,N_8976);
nand U14945 (N_14945,N_6576,N_9422);
or U14946 (N_14946,N_8574,N_5672);
or U14947 (N_14947,N_7232,N_6671);
nor U14948 (N_14948,N_7813,N_5353);
nand U14949 (N_14949,N_9726,N_5383);
nand U14950 (N_14950,N_6736,N_5626);
nand U14951 (N_14951,N_7779,N_8702);
xnor U14952 (N_14952,N_7856,N_9064);
xor U14953 (N_14953,N_9987,N_8383);
and U14954 (N_14954,N_5811,N_8696);
xnor U14955 (N_14955,N_7338,N_7943);
xor U14956 (N_14956,N_5361,N_9412);
xor U14957 (N_14957,N_6947,N_7836);
or U14958 (N_14958,N_8276,N_5298);
xor U14959 (N_14959,N_9882,N_7536);
and U14960 (N_14960,N_6951,N_7679);
and U14961 (N_14961,N_5331,N_5996);
xnor U14962 (N_14962,N_7031,N_9755);
and U14963 (N_14963,N_6652,N_9585);
or U14964 (N_14964,N_8556,N_6324);
nor U14965 (N_14965,N_6918,N_9663);
nor U14966 (N_14966,N_5822,N_6952);
and U14967 (N_14967,N_7565,N_9501);
xnor U14968 (N_14968,N_9914,N_9174);
or U14969 (N_14969,N_6793,N_5123);
xnor U14970 (N_14970,N_8892,N_7630);
xnor U14971 (N_14971,N_8751,N_6736);
nand U14972 (N_14972,N_5929,N_6363);
nor U14973 (N_14973,N_9715,N_6615);
nor U14974 (N_14974,N_6835,N_7473);
nor U14975 (N_14975,N_7046,N_6430);
and U14976 (N_14976,N_7475,N_7858);
xor U14977 (N_14977,N_9691,N_7035);
xor U14978 (N_14978,N_5727,N_8373);
xor U14979 (N_14979,N_5791,N_5914);
and U14980 (N_14980,N_9353,N_9756);
or U14981 (N_14981,N_7561,N_5093);
and U14982 (N_14982,N_7000,N_9975);
and U14983 (N_14983,N_6352,N_5000);
nand U14984 (N_14984,N_8609,N_8385);
nor U14985 (N_14985,N_9330,N_5003);
xor U14986 (N_14986,N_9752,N_9785);
nand U14987 (N_14987,N_8231,N_6070);
nor U14988 (N_14988,N_9698,N_6441);
nand U14989 (N_14989,N_7198,N_7304);
or U14990 (N_14990,N_6657,N_6584);
and U14991 (N_14991,N_9975,N_9235);
xor U14992 (N_14992,N_6698,N_9083);
xnor U14993 (N_14993,N_9789,N_8716);
xnor U14994 (N_14994,N_5588,N_7740);
nand U14995 (N_14995,N_9767,N_7646);
nand U14996 (N_14996,N_6772,N_5155);
nand U14997 (N_14997,N_5297,N_5241);
or U14998 (N_14998,N_5456,N_6182);
and U14999 (N_14999,N_9669,N_5779);
xnor UO_0 (O_0,N_14979,N_12777);
or UO_1 (O_1,N_14083,N_12542);
nor UO_2 (O_2,N_13168,N_12370);
nor UO_3 (O_3,N_12006,N_11228);
xor UO_4 (O_4,N_11312,N_10131);
nand UO_5 (O_5,N_11360,N_11324);
or UO_6 (O_6,N_13307,N_14832);
xnor UO_7 (O_7,N_10461,N_13067);
or UO_8 (O_8,N_11636,N_10211);
or UO_9 (O_9,N_14715,N_11529);
or UO_10 (O_10,N_13691,N_14171);
or UO_11 (O_11,N_14022,N_13896);
nand UO_12 (O_12,N_10778,N_11987);
xnor UO_13 (O_13,N_12819,N_13811);
xnor UO_14 (O_14,N_12228,N_13281);
nor UO_15 (O_15,N_14438,N_11980);
and UO_16 (O_16,N_12417,N_10314);
nor UO_17 (O_17,N_11180,N_10873);
nand UO_18 (O_18,N_11532,N_14904);
nand UO_19 (O_19,N_13618,N_14709);
and UO_20 (O_20,N_14454,N_11280);
and UO_21 (O_21,N_14426,N_11771);
nand UO_22 (O_22,N_10229,N_13620);
and UO_23 (O_23,N_10212,N_11624);
or UO_24 (O_24,N_13006,N_13016);
nand UO_25 (O_25,N_13101,N_13419);
xor UO_26 (O_26,N_14017,N_12199);
xor UO_27 (O_27,N_14195,N_14146);
or UO_28 (O_28,N_10750,N_12571);
xnor UO_29 (O_29,N_11459,N_12580);
and UO_30 (O_30,N_10444,N_14530);
nor UO_31 (O_31,N_11752,N_14970);
nand UO_32 (O_32,N_10071,N_10440);
and UO_33 (O_33,N_10107,N_14977);
and UO_34 (O_34,N_14114,N_14916);
or UO_35 (O_35,N_10341,N_14285);
or UO_36 (O_36,N_13424,N_12014);
nor UO_37 (O_37,N_11340,N_14663);
xor UO_38 (O_38,N_14096,N_10259);
xnor UO_39 (O_39,N_14913,N_11145);
or UO_40 (O_40,N_11817,N_10089);
and UO_41 (O_41,N_11622,N_13624);
nor UO_42 (O_42,N_13169,N_13868);
nand UO_43 (O_43,N_11387,N_10953);
nand UO_44 (O_44,N_10180,N_11538);
or UO_45 (O_45,N_11179,N_11915);
and UO_46 (O_46,N_12755,N_13496);
nand UO_47 (O_47,N_10017,N_11720);
nor UO_48 (O_48,N_10985,N_10906);
nand UO_49 (O_49,N_12793,N_14876);
nor UO_50 (O_50,N_13011,N_12357);
xnor UO_51 (O_51,N_12943,N_12154);
nand UO_52 (O_52,N_13999,N_14945);
xor UO_53 (O_53,N_14359,N_12535);
nand UO_54 (O_54,N_10464,N_14814);
nor UO_55 (O_55,N_14166,N_10082);
xor UO_56 (O_56,N_12207,N_10132);
nor UO_57 (O_57,N_11286,N_13909);
nand UO_58 (O_58,N_14725,N_10365);
nor UO_59 (O_59,N_14552,N_14445);
xor UO_60 (O_60,N_10226,N_13209);
nand UO_61 (O_61,N_13435,N_10401);
xnor UO_62 (O_62,N_14013,N_14626);
xor UO_63 (O_63,N_13605,N_14273);
xor UO_64 (O_64,N_12654,N_14525);
xor UO_65 (O_65,N_10659,N_10407);
or UO_66 (O_66,N_13702,N_14401);
nand UO_67 (O_67,N_12056,N_13747);
or UO_68 (O_68,N_13386,N_11645);
nor UO_69 (O_69,N_10821,N_12843);
xnor UO_70 (O_70,N_11036,N_12108);
xnor UO_71 (O_71,N_10110,N_13870);
and UO_72 (O_72,N_12776,N_12817);
nand UO_73 (O_73,N_11380,N_12497);
or UO_74 (O_74,N_10503,N_12834);
or UO_75 (O_75,N_14194,N_14356);
nor UO_76 (O_76,N_13364,N_13692);
nand UO_77 (O_77,N_13196,N_11059);
nand UO_78 (O_78,N_13544,N_14380);
xor UO_79 (O_79,N_12021,N_11982);
nand UO_80 (O_80,N_11735,N_12670);
nor UO_81 (O_81,N_13619,N_13256);
or UO_82 (O_82,N_11164,N_12892);
or UO_83 (O_83,N_12442,N_10342);
and UO_84 (O_84,N_13222,N_12951);
or UO_85 (O_85,N_14631,N_14211);
xor UO_86 (O_86,N_14065,N_10404);
xnor UO_87 (O_87,N_10125,N_12925);
xnor UO_88 (O_88,N_10427,N_14217);
nand UO_89 (O_89,N_12087,N_11253);
xnor UO_90 (O_90,N_12074,N_13672);
and UO_91 (O_91,N_14117,N_13321);
nand UO_92 (O_92,N_11346,N_10742);
or UO_93 (O_93,N_14005,N_13369);
or UO_94 (O_94,N_13934,N_12227);
xnor UO_95 (O_95,N_14960,N_11182);
or UO_96 (O_96,N_13684,N_14707);
nand UO_97 (O_97,N_12059,N_14115);
nor UO_98 (O_98,N_14405,N_10710);
and UO_99 (O_99,N_14125,N_12416);
nor UO_100 (O_100,N_11329,N_10815);
and UO_101 (O_101,N_13028,N_12893);
or UO_102 (O_102,N_13714,N_12932);
or UO_103 (O_103,N_12184,N_10679);
and UO_104 (O_104,N_13629,N_11582);
nor UO_105 (O_105,N_10773,N_12183);
nand UO_106 (O_106,N_13122,N_10391);
and UO_107 (O_107,N_13211,N_13856);
nand UO_108 (O_108,N_11745,N_11561);
xnor UO_109 (O_109,N_11569,N_11239);
or UO_110 (O_110,N_12725,N_10292);
nand UO_111 (O_111,N_12239,N_10465);
xor UO_112 (O_112,N_14705,N_10516);
or UO_113 (O_113,N_10301,N_11860);
nand UO_114 (O_114,N_10797,N_12702);
nor UO_115 (O_115,N_10002,N_14299);
xor UO_116 (O_116,N_11226,N_11090);
and UO_117 (O_117,N_13184,N_11251);
nand UO_118 (O_118,N_11306,N_11434);
nand UO_119 (O_119,N_11402,N_13349);
xnor UO_120 (O_120,N_12274,N_13189);
xnor UO_121 (O_121,N_14771,N_11767);
nand UO_122 (O_122,N_11870,N_11707);
and UO_123 (O_123,N_13442,N_13834);
nor UO_124 (O_124,N_12582,N_14233);
nand UO_125 (O_125,N_10696,N_14357);
nor UO_126 (O_126,N_10103,N_11456);
xor UO_127 (O_127,N_14752,N_13267);
or UO_128 (O_128,N_14720,N_11399);
and UO_129 (O_129,N_11833,N_10267);
nor UO_130 (O_130,N_12393,N_11323);
or UO_131 (O_131,N_12447,N_13363);
and UO_132 (O_132,N_14122,N_12944);
and UO_133 (O_133,N_11259,N_11295);
xor UO_134 (O_134,N_13855,N_12996);
xor UO_135 (O_135,N_14774,N_13548);
and UO_136 (O_136,N_11152,N_14089);
or UO_137 (O_137,N_12315,N_14662);
or UO_138 (O_138,N_12898,N_13495);
xnor UO_139 (O_139,N_13402,N_13697);
nor UO_140 (O_140,N_12909,N_12837);
xnor UO_141 (O_141,N_11773,N_11689);
and UO_142 (O_142,N_11025,N_12858);
xor UO_143 (O_143,N_10702,N_14883);
nor UO_144 (O_144,N_10166,N_14740);
xnor UO_145 (O_145,N_10854,N_11520);
nand UO_146 (O_146,N_10571,N_12999);
and UO_147 (O_147,N_11102,N_10263);
or UO_148 (O_148,N_13262,N_11045);
or UO_149 (O_149,N_10045,N_11785);
and UO_150 (O_150,N_10884,N_11037);
nand UO_151 (O_151,N_14926,N_11186);
and UO_152 (O_152,N_13054,N_11000);
or UO_153 (O_153,N_10044,N_10338);
or UO_154 (O_154,N_11511,N_11886);
and UO_155 (O_155,N_10435,N_14778);
and UO_156 (O_156,N_10540,N_13872);
or UO_157 (O_157,N_14834,N_12166);
nor UO_158 (O_158,N_10237,N_11921);
xnor UO_159 (O_159,N_10429,N_12242);
and UO_160 (O_160,N_10383,N_10526);
or UO_161 (O_161,N_11831,N_12450);
xnor UO_162 (O_162,N_11680,N_13205);
xor UO_163 (O_163,N_12591,N_12623);
or UO_164 (O_164,N_14566,N_10069);
and UO_165 (O_165,N_13430,N_14140);
or UO_166 (O_166,N_12729,N_14598);
and UO_167 (O_167,N_13833,N_10892);
nand UO_168 (O_168,N_10327,N_10294);
and UO_169 (O_169,N_10672,N_14290);
and UO_170 (O_170,N_11417,N_10923);
nor UO_171 (O_171,N_11033,N_14646);
nand UO_172 (O_172,N_11801,N_13270);
or UO_173 (O_173,N_10496,N_14579);
or UO_174 (O_174,N_14372,N_14167);
nand UO_175 (O_175,N_11082,N_14753);
xnor UO_176 (O_176,N_13533,N_14655);
nand UO_177 (O_177,N_12002,N_10618);
and UO_178 (O_178,N_14796,N_10645);
and UO_179 (O_179,N_12356,N_13519);
or UO_180 (O_180,N_13193,N_10802);
or UO_181 (O_181,N_13073,N_13686);
or UO_182 (O_182,N_14414,N_12413);
nand UO_183 (O_183,N_12480,N_10153);
and UO_184 (O_184,N_14717,N_13465);
and UO_185 (O_185,N_11461,N_10330);
xor UO_186 (O_186,N_12500,N_10369);
or UO_187 (O_187,N_14370,N_10991);
and UO_188 (O_188,N_11264,N_14982);
nand UO_189 (O_189,N_10978,N_13569);
and UO_190 (O_190,N_14345,N_11614);
nand UO_191 (O_191,N_10922,N_13542);
or UO_192 (O_192,N_13118,N_12386);
and UO_193 (O_193,N_14657,N_10176);
and UO_194 (O_194,N_11502,N_12699);
nand UO_195 (O_195,N_12621,N_13780);
nor UO_196 (O_196,N_10587,N_12853);
nor UO_197 (O_197,N_10971,N_13177);
xnor UO_198 (O_198,N_14640,N_11178);
nor UO_199 (O_199,N_11495,N_11026);
nor UO_200 (O_200,N_12887,N_12738);
and UO_201 (O_201,N_12923,N_11499);
nor UO_202 (O_202,N_11221,N_13514);
xnor UO_203 (O_203,N_12915,N_10860);
xor UO_204 (O_204,N_13730,N_11855);
nor UO_205 (O_205,N_13339,N_10996);
or UO_206 (O_206,N_14212,N_12380);
xnor UO_207 (O_207,N_10345,N_10049);
xor UO_208 (O_208,N_10782,N_10683);
and UO_209 (O_209,N_12201,N_11976);
nand UO_210 (O_210,N_10517,N_11054);
xnor UO_211 (O_211,N_10916,N_14928);
and UO_212 (O_212,N_10939,N_10812);
xor UO_213 (O_213,N_12489,N_10962);
nor UO_214 (O_214,N_12515,N_10572);
xor UO_215 (O_215,N_10631,N_10870);
nor UO_216 (O_216,N_13634,N_12363);
xor UO_217 (O_217,N_10373,N_11476);
xor UO_218 (O_218,N_10143,N_11258);
xnor UO_219 (O_219,N_10533,N_10480);
nand UO_220 (O_220,N_11302,N_11104);
nor UO_221 (O_221,N_10626,N_11255);
nand UO_222 (O_222,N_13788,N_13763);
xnor UO_223 (O_223,N_14809,N_13245);
or UO_224 (O_224,N_10570,N_14493);
and UO_225 (O_225,N_10300,N_14676);
nand UO_226 (O_226,N_13494,N_11269);
nor UO_227 (O_227,N_11115,N_13089);
xor UO_228 (O_228,N_12305,N_12409);
or UO_229 (O_229,N_14563,N_11047);
or UO_230 (O_230,N_14209,N_10515);
and UO_231 (O_231,N_11601,N_10989);
and UO_232 (O_232,N_11487,N_14489);
nor UO_233 (O_233,N_14637,N_10960);
xnor UO_234 (O_234,N_12773,N_14344);
and UO_235 (O_235,N_11917,N_14653);
nand UO_236 (O_236,N_13334,N_13188);
nand UO_237 (O_237,N_11074,N_11512);
nand UO_238 (O_238,N_13457,N_13756);
nand UO_239 (O_239,N_11204,N_10251);
or UO_240 (O_240,N_11687,N_14365);
or UO_241 (O_241,N_10690,N_11249);
xor UO_242 (O_242,N_10108,N_10956);
or UO_243 (O_243,N_12815,N_13475);
nand UO_244 (O_244,N_13461,N_14594);
nand UO_245 (O_245,N_11393,N_12096);
nand UO_246 (O_246,N_14902,N_10518);
nor UO_247 (O_247,N_12790,N_14784);
or UO_248 (O_248,N_13047,N_12960);
or UO_249 (O_249,N_11741,N_10935);
nand UO_250 (O_250,N_14284,N_14815);
nand UO_251 (O_251,N_13963,N_11382);
nand UO_252 (O_252,N_14549,N_11589);
nand UO_253 (O_253,N_11028,N_12237);
nor UO_254 (O_254,N_14072,N_10586);
nor UO_255 (O_255,N_12100,N_11523);
nor UO_256 (O_256,N_11130,N_12524);
and UO_257 (O_257,N_10832,N_10899);
or UO_258 (O_258,N_13796,N_12433);
or UO_259 (O_259,N_13058,N_11408);
nor UO_260 (O_260,N_12401,N_11001);
nand UO_261 (O_261,N_13317,N_10550);
nand UO_262 (O_262,N_11604,N_10177);
nand UO_263 (O_263,N_10824,N_14564);
nor UO_264 (O_264,N_10012,N_12816);
nand UO_265 (O_265,N_10336,N_12164);
and UO_266 (O_266,N_13035,N_12176);
xnor UO_267 (O_267,N_13652,N_10768);
or UO_268 (O_268,N_13421,N_11401);
and UO_269 (O_269,N_10312,N_12998);
or UO_270 (O_270,N_12446,N_11660);
and UO_271 (O_271,N_11057,N_13366);
and UO_272 (O_272,N_10183,N_10455);
and UO_273 (O_273,N_11658,N_11425);
xor UO_274 (O_274,N_11365,N_13335);
nand UO_275 (O_275,N_14839,N_14785);
or UO_276 (O_276,N_13023,N_12040);
nand UO_277 (O_277,N_10350,N_13264);
nand UO_278 (O_278,N_13647,N_12781);
nor UO_279 (O_279,N_11613,N_12663);
and UO_280 (O_280,N_12003,N_12089);
and UO_281 (O_281,N_10332,N_10741);
xor UO_282 (O_282,N_10561,N_11933);
or UO_283 (O_283,N_12029,N_10547);
nand UO_284 (O_284,N_10262,N_12309);
nor UO_285 (O_285,N_11681,N_14487);
xnor UO_286 (O_286,N_14110,N_14367);
and UO_287 (O_287,N_12402,N_10433);
nand UO_288 (O_288,N_12389,N_14739);
nor UO_289 (O_289,N_12861,N_10622);
and UO_290 (O_290,N_10412,N_10675);
or UO_291 (O_291,N_12831,N_12624);
nand UO_292 (O_292,N_13947,N_14260);
and UO_293 (O_293,N_10254,N_12655);
xor UO_294 (O_294,N_10296,N_14429);
nand UO_295 (O_295,N_12737,N_14817);
nor UO_296 (O_296,N_13219,N_13815);
nor UO_297 (O_297,N_12338,N_11804);
and UO_298 (O_298,N_14906,N_14931);
and UO_299 (O_299,N_10029,N_13832);
nand UO_300 (O_300,N_11042,N_13762);
nand UO_301 (O_301,N_13485,N_14136);
xor UO_302 (O_302,N_13125,N_13394);
nor UO_303 (O_303,N_12300,N_10168);
and UO_304 (O_304,N_12253,N_11939);
or UO_305 (O_305,N_11023,N_14079);
xor UO_306 (O_306,N_13809,N_13766);
or UO_307 (O_307,N_12522,N_14193);
xnor UO_308 (O_308,N_12764,N_10370);
and UO_309 (O_309,N_10459,N_12196);
nand UO_310 (O_310,N_14866,N_10646);
xor UO_311 (O_311,N_14342,N_13604);
nor UO_312 (O_312,N_14247,N_10390);
nor UO_313 (O_313,N_14292,N_14965);
xnor UO_314 (O_314,N_11270,N_14045);
nor UO_315 (O_315,N_10175,N_14840);
nand UO_316 (O_316,N_14302,N_12607);
xnor UO_317 (O_317,N_13466,N_12200);
xnor UO_318 (O_318,N_10420,N_13013);
or UO_319 (O_319,N_10806,N_10232);
xnor UO_320 (O_320,N_14076,N_10452);
or UO_321 (O_321,N_14607,N_14387);
nor UO_322 (O_322,N_14295,N_10167);
nor UO_323 (O_323,N_11814,N_14270);
and UO_324 (O_324,N_14205,N_10904);
or UO_325 (O_325,N_10919,N_11567);
nor UO_326 (O_326,N_12611,N_10719);
nor UO_327 (O_327,N_10780,N_14035);
nand UO_328 (O_328,N_13083,N_11547);
and UO_329 (O_329,N_10781,N_12286);
xor UO_330 (O_330,N_13113,N_13260);
nor UO_331 (O_331,N_14844,N_12523);
xnor UO_332 (O_332,N_11826,N_10559);
nor UO_333 (O_333,N_12826,N_10328);
xnor UO_334 (O_334,N_14777,N_12516);
nand UO_335 (O_335,N_11568,N_11682);
xor UO_336 (O_336,N_11637,N_13354);
and UO_337 (O_337,N_10952,N_12246);
or UO_338 (O_338,N_13857,N_13153);
and UO_339 (O_339,N_14148,N_12365);
nor UO_340 (O_340,N_14080,N_14239);
and UO_341 (O_341,N_12874,N_14573);
nand UO_342 (O_342,N_11667,N_11918);
and UO_343 (O_343,N_12374,N_11010);
xnor UO_344 (O_344,N_13900,N_11555);
xor UO_345 (O_345,N_13358,N_12634);
or UO_346 (O_346,N_14541,N_12175);
nand UO_347 (O_347,N_14128,N_10134);
and UO_348 (O_348,N_10475,N_10275);
and UO_349 (O_349,N_13899,N_10823);
or UO_350 (O_350,N_14716,N_11384);
nor UO_351 (O_351,N_11428,N_10026);
or UO_352 (O_352,N_12855,N_12529);
nor UO_353 (O_353,N_12674,N_11595);
nor UO_354 (O_354,N_10621,N_14461);
or UO_355 (O_355,N_10640,N_12977);
nor UO_356 (O_356,N_12366,N_14729);
nand UO_357 (O_357,N_11311,N_14535);
nand UO_358 (O_358,N_14410,N_12209);
nand UO_359 (O_359,N_11652,N_14590);
and UO_360 (O_360,N_11992,N_13266);
nor UO_361 (O_361,N_11677,N_11034);
nor UO_362 (O_362,N_14813,N_14519);
nand UO_363 (O_363,N_10510,N_12602);
xor UO_364 (O_364,N_13156,N_14320);
xor UO_365 (O_365,N_10054,N_10963);
nand UO_366 (O_366,N_12323,N_14313);
and UO_367 (O_367,N_14828,N_11800);
xnor UO_368 (O_368,N_14944,N_12035);
xnor UO_369 (O_369,N_12851,N_14693);
nand UO_370 (O_370,N_10616,N_14862);
or UO_371 (O_371,N_12839,N_10743);
or UO_372 (O_372,N_13426,N_10499);
nor UO_373 (O_373,N_14231,N_10717);
nand UO_374 (O_374,N_11430,N_10076);
or UO_375 (O_375,N_14742,N_12313);
nor UO_376 (O_376,N_11247,N_10654);
nor UO_377 (O_377,N_10067,N_13477);
nor UO_378 (O_378,N_13994,N_12260);
and UO_379 (O_379,N_14789,N_14491);
or UO_380 (O_380,N_14517,N_14923);
or UO_381 (O_381,N_10446,N_13926);
nand UO_382 (O_382,N_12197,N_11156);
nand UO_383 (O_383,N_14173,N_12660);
nand UO_384 (O_384,N_13212,N_13649);
and UO_385 (O_385,N_11497,N_10170);
nor UO_386 (O_386,N_10508,N_10347);
and UO_387 (O_387,N_10228,N_10399);
xnor UO_388 (O_388,N_10593,N_10633);
nand UO_389 (O_389,N_13302,N_11548);
or UO_390 (O_390,N_14240,N_10439);
nand UO_391 (O_391,N_12727,N_13464);
nor UO_392 (O_392,N_10008,N_12597);
xnor UO_393 (O_393,N_12712,N_11849);
or UO_394 (O_394,N_13094,N_12949);
xnor UO_395 (O_395,N_14137,N_13803);
or UO_396 (O_396,N_13659,N_11278);
nand UO_397 (O_397,N_11978,N_10409);
xor UO_398 (O_398,N_14388,N_13412);
nand UO_399 (O_399,N_14836,N_12687);
xor UO_400 (O_400,N_10882,N_13888);
and UO_401 (O_401,N_11676,N_11368);
nand UO_402 (O_402,N_12517,N_14330);
nor UO_403 (O_403,N_10493,N_11513);
or UO_404 (O_404,N_14948,N_13539);
nand UO_405 (O_405,N_14722,N_14800);
nand UO_406 (O_406,N_10512,N_13395);
nand UO_407 (O_407,N_10995,N_11101);
or UO_408 (O_408,N_14097,N_13079);
xnor UO_409 (O_409,N_11443,N_13924);
nand UO_410 (O_410,N_13069,N_13187);
nand UO_411 (O_411,N_11039,N_10794);
nor UO_412 (O_412,N_11140,N_13905);
or UO_413 (O_413,N_11373,N_12107);
nor UO_414 (O_414,N_14064,N_13308);
or UO_415 (O_415,N_13032,N_11218);
nor UO_416 (O_416,N_14155,N_11193);
xnor UO_417 (O_417,N_12694,N_13824);
xor UO_418 (O_418,N_12105,N_14478);
nand UO_419 (O_419,N_14391,N_14037);
and UO_420 (O_420,N_10744,N_12440);
and UO_421 (O_421,N_13883,N_14936);
nor UO_422 (O_422,N_13432,N_10430);
or UO_423 (O_423,N_13448,N_13493);
or UO_424 (O_424,N_12102,N_11926);
and UO_425 (O_425,N_10731,N_12956);
xnor UO_426 (O_426,N_11566,N_13626);
xnor UO_427 (O_427,N_14737,N_13879);
and UO_428 (O_428,N_11799,N_14608);
and UO_429 (O_429,N_10681,N_13781);
nand UO_430 (O_430,N_12398,N_10997);
xnor UO_431 (O_431,N_12975,N_12347);
nor UO_432 (O_432,N_10657,N_14690);
xnor UO_433 (O_433,N_13148,N_13190);
and UO_434 (O_434,N_12532,N_12772);
or UO_435 (O_435,N_10596,N_13436);
and UO_436 (O_436,N_14932,N_10145);
nor UO_437 (O_437,N_10942,N_11895);
nor UO_438 (O_438,N_13850,N_11824);
and UO_439 (O_439,N_14534,N_10663);
nand UO_440 (O_440,N_11646,N_13564);
nor UO_441 (O_441,N_10306,N_11008);
xnor UO_442 (O_442,N_10257,N_11150);
nand UO_443 (O_443,N_13607,N_14484);
and UO_444 (O_444,N_14465,N_12595);
nand UO_445 (O_445,N_13473,N_13042);
and UO_446 (O_446,N_11449,N_14020);
and UO_447 (O_447,N_13852,N_11069);
or UO_448 (O_448,N_10457,N_11787);
and UO_449 (O_449,N_12866,N_11421);
nor UO_450 (O_450,N_13874,N_13330);
xnor UO_451 (O_451,N_10091,N_14886);
nand UO_452 (O_452,N_10685,N_13463);
and UO_453 (O_453,N_10015,N_13737);
xnor UO_454 (O_454,N_12069,N_14243);
and UO_455 (O_455,N_10558,N_11858);
nor UO_456 (O_456,N_14048,N_11097);
or UO_457 (O_457,N_12519,N_12275);
nand UO_458 (O_458,N_12296,N_12444);
nor UO_459 (O_459,N_11293,N_13836);
nor UO_460 (O_460,N_10410,N_11930);
nor UO_461 (O_461,N_13954,N_14085);
and UO_462 (O_462,N_11083,N_12420);
nor UO_463 (O_463,N_11431,N_13043);
or UO_464 (O_464,N_12558,N_12361);
xor UO_465 (O_465,N_10613,N_12697);
and UO_466 (O_466,N_14255,N_14569);
nand UO_467 (O_467,N_11126,N_12410);
nand UO_468 (O_468,N_10118,N_13782);
nand UO_469 (O_469,N_14130,N_13246);
nand UO_470 (O_470,N_10491,N_14529);
nor UO_471 (O_471,N_14939,N_14054);
or UO_472 (O_472,N_13490,N_14609);
nor UO_473 (O_473,N_11436,N_12526);
nor UO_474 (O_474,N_11157,N_10800);
and UO_475 (O_475,N_13746,N_12736);
or UO_476 (O_476,N_14093,N_12490);
and UO_477 (O_477,N_13038,N_12412);
or UO_478 (O_478,N_13716,N_13429);
or UO_479 (O_479,N_13526,N_14600);
nor UO_480 (O_480,N_10767,N_13090);
or UO_481 (O_481,N_11922,N_11798);
and UO_482 (O_482,N_12026,N_12862);
or UO_483 (O_483,N_14102,N_12562);
and UO_484 (O_484,N_13258,N_10915);
or UO_485 (O_485,N_11713,N_12560);
or UO_486 (O_486,N_11759,N_12474);
nor UO_487 (O_487,N_11490,N_13971);
and UO_488 (O_488,N_11406,N_14196);
nor UO_489 (O_489,N_12276,N_11943);
and UO_490 (O_490,N_13010,N_10891);
nand UO_491 (O_491,N_14523,N_14856);
xnor UO_492 (O_492,N_10691,N_13978);
xor UO_493 (O_493,N_10426,N_11363);
xnor UO_494 (O_494,N_11577,N_10466);
and UO_495 (O_495,N_13116,N_13243);
xor UO_496 (O_496,N_10129,N_13183);
xor UO_497 (O_497,N_12880,N_10274);
nand UO_498 (O_498,N_13992,N_13411);
or UO_499 (O_499,N_13995,N_12700);
and UO_500 (O_500,N_10454,N_13743);
or UO_501 (O_501,N_14287,N_12289);
or UO_502 (O_502,N_12483,N_11465);
nand UO_503 (O_503,N_10889,N_14498);
nand UO_504 (O_504,N_14221,N_12901);
or UO_505 (O_505,N_13843,N_10227);
xnor UO_506 (O_506,N_13422,N_10712);
xnor UO_507 (O_507,N_14213,N_10965);
or UO_508 (O_508,N_14891,N_14872);
nand UO_509 (O_509,N_10172,N_14066);
nor UO_510 (O_510,N_12078,N_11233);
nor UO_511 (O_511,N_13581,N_14440);
or UO_512 (O_512,N_13603,N_13009);
and UO_513 (O_513,N_10133,N_12718);
or UO_514 (O_514,N_12448,N_11349);
nor UO_515 (O_515,N_11095,N_12921);
or UO_516 (O_516,N_11794,N_10972);
nor UO_517 (O_517,N_12481,N_14603);
and UO_518 (O_518,N_14734,N_13361);
nand UO_519 (O_519,N_12954,N_11386);
xor UO_520 (O_520,N_14689,N_12377);
xor UO_521 (O_521,N_10286,N_11050);
nand UO_522 (O_522,N_13165,N_11167);
and UO_523 (O_523,N_13352,N_10438);
or UO_524 (O_524,N_14721,N_11321);
nor UO_525 (O_525,N_11112,N_10727);
nor UO_526 (O_526,N_14994,N_14003);
nor UO_527 (O_527,N_10472,N_11643);
xnor UO_528 (O_528,N_12639,N_13131);
or UO_529 (O_529,N_11928,N_14667);
nor UO_530 (O_530,N_13860,N_12011);
nand UO_531 (O_531,N_11650,N_10834);
and UO_532 (O_532,N_10243,N_10519);
and UO_533 (O_533,N_12695,N_14610);
xor UO_534 (O_534,N_14764,N_11195);
or UO_535 (O_535,N_14808,N_12742);
nand UO_536 (O_536,N_14160,N_11072);
nor UO_537 (O_537,N_10195,N_12650);
xor UO_538 (O_538,N_13606,N_10605);
xnor UO_539 (O_539,N_11942,N_10214);
and UO_540 (O_540,N_10062,N_14679);
and UO_541 (O_541,N_13044,N_12077);
and UO_542 (O_542,N_14269,N_13949);
nand UO_543 (O_543,N_14375,N_10122);
nor UO_544 (O_544,N_12939,N_14812);
nand UO_545 (O_545,N_14470,N_12995);
nand UO_546 (O_546,N_12512,N_11170);
nor UO_547 (O_547,N_11602,N_12254);
or UO_548 (O_548,N_14578,N_14111);
xor UO_549 (O_549,N_10162,N_12139);
or UO_550 (O_550,N_14431,N_13158);
or UO_551 (O_551,N_12429,N_12137);
nand UO_552 (O_552,N_10920,N_12280);
and UO_553 (O_553,N_11543,N_13797);
nand UO_554 (O_554,N_11261,N_12092);
and UO_555 (O_555,N_14559,N_12959);
xnor UO_556 (O_556,N_13980,N_11232);
or UO_557 (O_557,N_13390,N_11970);
nand UO_558 (O_558,N_14200,N_13761);
xnor UO_559 (O_559,N_11730,N_10846);
nand UO_560 (O_560,N_13972,N_13481);
and UO_561 (O_561,N_14069,N_12734);
nor UO_562 (O_562,N_12156,N_13810);
or UO_563 (O_563,N_14376,N_12933);
xnor UO_564 (O_564,N_10179,N_12608);
nor UO_565 (O_565,N_11908,N_10574);
or UO_566 (O_566,N_10056,N_13765);
xor UO_567 (O_567,N_12173,N_13142);
and UO_568 (O_568,N_13690,N_13572);
or UO_569 (O_569,N_11158,N_13878);
nand UO_570 (O_570,N_12885,N_11993);
or UO_571 (O_571,N_12544,N_13795);
and UO_572 (O_572,N_14068,N_11761);
or UO_573 (O_573,N_10458,N_13382);
nand UO_574 (O_574,N_11403,N_12924);
or UO_575 (O_575,N_10554,N_13310);
nand UO_576 (O_576,N_11884,N_12797);
and UO_577 (O_577,N_11536,N_10692);
and UO_578 (O_578,N_12080,N_14358);
and UO_579 (O_579,N_13085,N_14620);
xor UO_580 (O_580,N_13749,N_10708);
xnor UO_581 (O_581,N_14546,N_13884);
and UO_582 (O_582,N_13574,N_12701);
and UO_583 (O_583,N_10527,N_10334);
xnor UO_584 (O_584,N_11721,N_14057);
or UO_585 (O_585,N_11208,N_11829);
nor UO_586 (O_586,N_13232,N_10735);
and UO_587 (O_587,N_14700,N_11725);
xor UO_588 (O_588,N_12667,N_11108);
xnor UO_589 (O_589,N_12072,N_14539);
nor UO_590 (O_590,N_11951,N_14801);
or UO_591 (O_591,N_14855,N_11273);
xnor UO_592 (O_592,N_14369,N_13541);
xnor UO_593 (O_593,N_14918,N_10878);
nor UO_594 (O_594,N_13105,N_13055);
nand UO_595 (O_595,N_10113,N_13141);
nand UO_596 (O_596,N_14222,N_13641);
nand UO_597 (O_597,N_14857,N_12930);
nor UO_598 (O_598,N_13365,N_11277);
or UO_599 (O_599,N_14682,N_12589);
and UO_600 (O_600,N_13420,N_13751);
or UO_601 (O_601,N_13709,N_13408);
nand UO_602 (O_602,N_10661,N_11961);
and UO_603 (O_603,N_13320,N_14592);
and UO_604 (O_604,N_12635,N_12916);
or UO_605 (O_605,N_11584,N_10303);
and UO_606 (O_606,N_13826,N_13774);
or UO_607 (O_607,N_14123,N_13095);
nand UO_608 (O_608,N_12530,N_11374);
nor UO_609 (O_609,N_10666,N_10836);
or UO_610 (O_610,N_14355,N_12600);
or UO_611 (O_611,N_14001,N_13441);
or UO_612 (O_612,N_11784,N_10908);
xnor UO_613 (O_613,N_14303,N_12133);
nor UO_614 (O_614,N_10885,N_10964);
xor UO_615 (O_615,N_10694,N_11203);
nand UO_616 (O_616,N_12469,N_14185);
and UO_617 (O_617,N_13121,N_11125);
and UO_618 (O_618,N_13527,N_10667);
nor UO_619 (O_619,N_11141,N_13471);
or UO_620 (O_620,N_11089,N_13942);
nor UO_621 (O_621,N_10190,N_12267);
or UO_622 (O_622,N_11587,N_13806);
nor UO_623 (O_623,N_14134,N_14371);
or UO_624 (O_624,N_11444,N_14187);
or UO_625 (O_625,N_11751,N_13478);
and UO_626 (O_626,N_13825,N_12271);
nand UO_627 (O_627,N_11290,N_14423);
or UO_628 (O_628,N_14606,N_11958);
and UO_629 (O_629,N_12703,N_13708);
xor UO_630 (O_630,N_10238,N_12093);
xnor UO_631 (O_631,N_12550,N_11452);
nand UO_632 (O_632,N_12493,N_12626);
xnor UO_633 (O_633,N_10689,N_10219);
xor UO_634 (O_634,N_11289,N_13557);
nand UO_635 (O_635,N_10772,N_13521);
nand UO_636 (O_636,N_10470,N_12810);
nor UO_637 (O_637,N_12820,N_11129);
or UO_638 (O_638,N_13842,N_11351);
nand UO_639 (O_639,N_12032,N_12945);
and UO_640 (O_640,N_14557,N_12470);
nor UO_641 (O_641,N_13120,N_14075);
or UO_642 (O_642,N_10147,N_14047);
and UO_643 (O_643,N_10022,N_14754);
xnor UO_644 (O_644,N_11211,N_13958);
nor UO_645 (O_645,N_12958,N_10987);
and UO_646 (O_646,N_14691,N_13546);
and UO_647 (O_647,N_11729,N_10912);
xnor UO_648 (O_648,N_10386,N_12174);
or UO_649 (O_649,N_11032,N_11600);
or UO_650 (O_650,N_13917,N_11812);
xnor UO_651 (O_651,N_11537,N_12453);
nor UO_652 (O_652,N_14540,N_12691);
nor UO_653 (O_653,N_11096,N_10789);
or UO_654 (O_654,N_12037,N_11830);
nor UO_655 (O_655,N_10380,N_12645);
xnor UO_656 (O_656,N_10722,N_14018);
xnor UO_657 (O_657,N_10174,N_13162);
nand UO_658 (O_658,N_14803,N_13813);
xor UO_659 (O_659,N_11336,N_10652);
nor UO_660 (O_660,N_12301,N_12963);
or UO_661 (O_661,N_13271,N_11626);
xor UO_662 (O_662,N_11846,N_11313);
or UO_663 (O_663,N_10748,N_13964);
nand UO_664 (O_664,N_10793,N_12038);
nand UO_665 (O_665,N_14584,N_11376);
nand UO_666 (O_666,N_11791,N_12726);
xnor UO_667 (O_667,N_12989,N_10387);
and UO_668 (O_668,N_10842,N_10047);
nand UO_669 (O_669,N_12573,N_14978);
and UO_670 (O_670,N_10413,N_10253);
and UO_671 (O_671,N_11006,N_11946);
xor UO_672 (O_672,N_12510,N_12619);
nor UO_673 (O_673,N_10396,N_11891);
xnor UO_674 (O_674,N_12747,N_12706);
or UO_675 (O_675,N_14805,N_12459);
nand UO_676 (O_676,N_13739,N_14787);
xor UO_677 (O_677,N_13288,N_12328);
nand UO_678 (O_678,N_14095,N_12912);
or UO_679 (O_679,N_12213,N_12934);
nor UO_680 (O_680,N_13907,N_14379);
or UO_681 (O_681,N_13719,N_14150);
xor UO_682 (O_682,N_11136,N_11803);
xnor UO_683 (O_683,N_13586,N_11863);
and UO_684 (O_684,N_14030,N_11510);
nor UO_685 (O_685,N_12050,N_13694);
nand UO_686 (O_686,N_10567,N_13863);
nand UO_687 (O_687,N_13996,N_14373);
nor UO_688 (O_688,N_10864,N_13231);
or UO_689 (O_689,N_10907,N_13663);
or UO_690 (O_690,N_11189,N_13182);
and UO_691 (O_691,N_13476,N_12025);
nor UO_692 (O_692,N_11257,N_13946);
nand UO_693 (O_693,N_13594,N_10575);
nand UO_694 (O_694,N_11350,N_10283);
nor UO_695 (O_695,N_12863,N_12060);
nand UO_696 (O_696,N_11960,N_12770);
xnor UO_697 (O_697,N_13437,N_11719);
and UO_698 (O_698,N_11364,N_14268);
nand UO_699 (O_699,N_10389,N_10311);
or UO_700 (O_700,N_10098,N_12662);
xor UO_701 (O_701,N_11056,N_11040);
or UO_702 (O_702,N_12083,N_12596);
and UO_703 (O_703,N_13670,N_12594);
and UO_704 (O_704,N_13588,N_14458);
nand UO_705 (O_705,N_12163,N_14668);
xor UO_706 (O_706,N_11342,N_11768);
nand UO_707 (O_707,N_13129,N_10579);
xor UO_708 (O_708,N_10988,N_10351);
or UO_709 (O_709,N_12218,N_11690);
nand UO_710 (O_710,N_14781,N_14407);
xnor UO_711 (O_711,N_12479,N_12877);
xor UO_712 (O_712,N_14920,N_12145);
nor UO_713 (O_713,N_13912,N_12814);
nand UO_714 (O_714,N_13773,N_12717);
xnor UO_715 (O_715,N_13643,N_11770);
and UO_716 (O_716,N_13019,N_13237);
xnor UO_717 (O_717,N_14341,N_10867);
nand UO_718 (O_718,N_10046,N_12972);
nor UO_719 (O_719,N_13727,N_10140);
xnor UO_720 (O_720,N_11686,N_14437);
or UO_721 (O_721,N_11868,N_12929);
xnor UO_722 (O_722,N_11254,N_10425);
nor UO_723 (O_723,N_10739,N_13425);
and UO_724 (O_724,N_12900,N_11137);
xor UO_725 (O_725,N_11494,N_12657);
xnor UO_726 (O_726,N_10529,N_10447);
xnor UO_727 (O_727,N_10304,N_10932);
nand UO_728 (O_728,N_10848,N_11107);
nor UO_729 (O_729,N_13505,N_11427);
nand UO_730 (O_730,N_11688,N_13392);
and UO_731 (O_731,N_10900,N_14275);
and UO_732 (O_732,N_14133,N_13400);
or UO_733 (O_733,N_13589,N_14432);
and UO_734 (O_734,N_11337,N_12158);
or UO_735 (O_735,N_12191,N_13197);
or UO_736 (O_736,N_12167,N_12187);
or UO_737 (O_737,N_10948,N_14158);
and UO_738 (O_738,N_14002,N_10424);
and UO_739 (O_739,N_10777,N_13889);
or UO_740 (O_740,N_10097,N_14542);
nand UO_741 (O_741,N_12569,N_11931);
and UO_742 (O_742,N_12279,N_11395);
nor UO_743 (O_743,N_14683,N_14315);
nand UO_744 (O_744,N_11509,N_14650);
nand UO_745 (O_745,N_10157,N_11116);
nor UO_746 (O_746,N_11437,N_14561);
and UO_747 (O_747,N_12928,N_12149);
or UO_748 (O_748,N_11551,N_14382);
xnor UO_749 (O_749,N_12752,N_14070);
nor UO_750 (O_750,N_10418,N_10200);
and UO_751 (O_751,N_13904,N_14353);
and UO_752 (O_752,N_13528,N_10930);
or UO_753 (O_753,N_13053,N_14894);
xnor UO_754 (O_754,N_12368,N_11919);
nand UO_755 (O_755,N_13835,N_13297);
nor UO_756 (O_756,N_10024,N_11671);
xor UO_757 (O_757,N_14386,N_12907);
nor UO_758 (O_758,N_14508,N_13931);
and UO_759 (O_759,N_14642,N_12955);
xor UO_760 (O_760,N_13285,N_13837);
or UO_761 (O_761,N_12169,N_11873);
or UO_762 (O_762,N_13214,N_11880);
and UO_763 (O_763,N_13789,N_11462);
nand UO_764 (O_764,N_10437,N_12112);
or UO_765 (O_765,N_10543,N_12664);
nor UO_766 (O_766,N_11969,N_14870);
xnor UO_767 (O_767,N_11937,N_10757);
and UO_768 (O_768,N_10755,N_14168);
xor UO_769 (O_769,N_10343,N_13235);
or UO_770 (O_770,N_11563,N_14311);
or UO_771 (O_771,N_10220,N_10173);
and UO_772 (O_772,N_12787,N_13701);
xor UO_773 (O_773,N_13012,N_12642);
or UO_774 (O_774,N_14164,N_14686);
or UO_775 (O_775,N_10994,N_12762);
nand UO_776 (O_776,N_11925,N_12430);
and UO_777 (O_777,N_10265,N_10820);
nand UO_778 (O_778,N_12128,N_14572);
nor UO_779 (O_779,N_14408,N_10302);
or UO_780 (O_780,N_12856,N_11782);
and UO_781 (O_781,N_11229,N_14238);
and UO_782 (O_782,N_14450,N_11753);
and UO_783 (O_783,N_11709,N_12293);
and UO_784 (O_784,N_14029,N_10595);
or UO_785 (O_785,N_11924,N_12321);
xor UO_786 (O_786,N_11810,N_13350);
nor UO_787 (O_787,N_10406,N_13941);
nand UO_788 (O_788,N_11883,N_12606);
and UO_789 (O_789,N_11067,N_13819);
and UO_790 (O_790,N_11439,N_14976);
nand UO_791 (O_791,N_11058,N_13099);
or UO_792 (O_792,N_14937,N_12728);
xor UO_793 (O_793,N_14512,N_11727);
and UO_794 (O_794,N_10651,N_12653);
nor UO_795 (O_795,N_10171,N_11644);
xor UO_796 (O_796,N_13200,N_14232);
nor UO_797 (O_797,N_12709,N_11005);
and UO_798 (O_798,N_12298,N_14654);
or UO_799 (O_799,N_12452,N_11972);
xor UO_800 (O_800,N_13251,N_10146);
nand UO_801 (O_801,N_14266,N_13668);
nor UO_802 (O_802,N_10340,N_10753);
or UO_803 (O_803,N_13704,N_10319);
or UO_804 (O_804,N_11262,N_10033);
nor UO_805 (O_805,N_13367,N_14871);
xor UO_806 (O_806,N_14826,N_10072);
nor UO_807 (O_807,N_11556,N_13936);
or UO_808 (O_808,N_13202,N_10261);
nor UO_809 (O_809,N_11455,N_11177);
nor UO_810 (O_810,N_14163,N_13524);
nand UO_811 (O_811,N_14101,N_11453);
or UO_812 (O_812,N_10368,N_14203);
xor UO_813 (O_813,N_12974,N_11841);
nand UO_814 (O_814,N_13908,N_14460);
and UO_815 (O_815,N_11412,N_10552);
and UO_816 (O_816,N_11834,N_10423);
nand UO_817 (O_817,N_12774,N_14751);
nand UO_818 (O_818,N_12865,N_14161);
or UO_819 (O_819,N_11984,N_11017);
xnor UO_820 (O_820,N_13301,N_10144);
or UO_821 (O_821,N_13623,N_10880);
nor UO_822 (O_822,N_11748,N_10467);
nor UO_823 (O_823,N_14648,N_11766);
nand UO_824 (O_824,N_10320,N_13050);
nor UO_825 (O_825,N_10641,N_11728);
xnor UO_826 (O_826,N_14685,N_11004);
xor UO_827 (O_827,N_13720,N_11708);
and UO_828 (O_828,N_11131,N_13841);
nand UO_829 (O_829,N_12118,N_14264);
nand UO_830 (O_830,N_14567,N_13895);
xor UO_831 (O_831,N_13325,N_13025);
nor UO_832 (O_832,N_13591,N_10804);
or UO_833 (O_833,N_10382,N_12024);
nor UO_834 (O_834,N_11088,N_13385);
xor UO_835 (O_835,N_13252,N_12425);
xor UO_836 (O_836,N_12391,N_10199);
and UO_837 (O_837,N_11248,N_10609);
nor UO_838 (O_838,N_10321,N_11263);
or UO_839 (O_839,N_14040,N_12085);
nand UO_840 (O_840,N_13783,N_11084);
xnor UO_841 (O_841,N_10449,N_13208);
or UO_842 (O_842,N_12219,N_12572);
or UO_843 (O_843,N_14497,N_10436);
xor UO_844 (O_844,N_12257,N_12553);
nand UO_845 (O_845,N_13440,N_13480);
xnor UO_846 (O_846,N_10509,N_14280);
and UO_847 (O_847,N_10127,N_10866);
and UO_848 (O_848,N_14571,N_10921);
or UO_849 (O_849,N_10600,N_11504);
xor UO_850 (O_850,N_14306,N_14957);
or UO_851 (O_851,N_13845,N_13048);
or UO_852 (O_852,N_13956,N_13677);
xor UO_853 (O_853,N_10507,N_14241);
xnor UO_854 (O_854,N_14394,N_14000);
nand UO_855 (O_855,N_13096,N_11007);
nor UO_856 (O_856,N_11710,N_10537);
nand UO_857 (O_857,N_11018,N_10688);
nor UO_858 (O_858,N_12766,N_10576);
nor UO_859 (O_859,N_14746,N_11128);
and UO_860 (O_860,N_12116,N_12058);
nand UO_861 (O_861,N_13700,N_13123);
and UO_862 (O_862,N_13787,N_10326);
nand UO_863 (O_863,N_14204,N_13580);
xnor UO_864 (O_864,N_11066,N_14215);
nand UO_865 (O_865,N_14515,N_11171);
nand UO_866 (O_866,N_12171,N_11953);
nor UO_867 (O_867,N_14276,N_13397);
nor UO_868 (O_868,N_11612,N_12455);
nand UO_869 (O_869,N_12878,N_14704);
xnor UO_870 (O_870,N_13206,N_14797);
nand UO_871 (O_871,N_12036,N_13736);
xor UO_872 (O_872,N_13414,N_12099);
nand UO_873 (O_873,N_10159,N_11044);
and UO_874 (O_874,N_12981,N_12685);
xor UO_875 (O_875,N_13886,N_14043);
nand UO_876 (O_876,N_12343,N_13640);
xnor UO_877 (O_877,N_13760,N_11298);
or UO_878 (O_878,N_10986,N_14500);
or UO_879 (O_879,N_13160,N_14092);
and UO_880 (O_880,N_11916,N_11955);
and UO_881 (O_881,N_10305,N_13744);
xnor UO_882 (O_882,N_12574,N_12075);
nand UO_883 (O_883,N_14378,N_12247);
nand UO_884 (O_884,N_11634,N_11410);
and UO_885 (O_885,N_13568,N_11534);
nand UO_886 (O_886,N_10745,N_14377);
nor UO_887 (O_887,N_11716,N_10644);
nand UO_888 (O_888,N_10857,N_12796);
nand UO_889 (O_889,N_11576,N_10523);
nand UO_890 (O_890,N_12292,N_11518);
nor UO_891 (O_891,N_13119,N_14947);
nand UO_892 (O_892,N_13499,N_14651);
xor UO_893 (O_893,N_12475,N_12903);
nor UO_894 (O_894,N_11398,N_11736);
nand UO_895 (O_895,N_13407,N_12800);
or UO_896 (O_896,N_12588,N_12875);
nor UO_897 (O_897,N_14479,N_11998);
xor UO_898 (O_898,N_10375,N_14113);
and UO_899 (O_899,N_13814,N_12577);
or UO_900 (O_900,N_12964,N_14361);
nand UO_901 (O_901,N_11188,N_13145);
or UO_902 (O_902,N_14420,N_13234);
nand UO_903 (O_903,N_10169,N_12195);
nor UO_904 (O_904,N_12299,N_14518);
nor UO_905 (O_905,N_13520,N_11483);
xnor UO_906 (O_906,N_12106,N_12097);
xnor UO_907 (O_907,N_13289,N_14263);
or UO_908 (O_908,N_13977,N_11415);
or UO_909 (O_909,N_12756,N_13768);
or UO_910 (O_910,N_13304,N_13660);
nand UO_911 (O_911,N_14457,N_10414);
or UO_912 (O_912,N_14286,N_13752);
nor UO_913 (O_913,N_13331,N_13439);
or UO_914 (O_914,N_11281,N_11147);
and UO_915 (O_915,N_12644,N_12259);
nand UO_916 (O_916,N_14680,N_14711);
xor UO_917 (O_917,N_14724,N_12922);
nand UO_918 (O_918,N_10723,N_13757);
nor UO_919 (O_919,N_10270,N_11003);
or UO_920 (O_920,N_11020,N_13890);
xnor UO_921 (O_921,N_14595,N_13323);
or UO_922 (O_922,N_14183,N_11021);
nor UO_923 (O_923,N_13867,N_13117);
xnor UO_924 (O_924,N_10116,N_11482);
and UO_925 (O_925,N_10085,N_11839);
or UO_926 (O_926,N_12335,N_10359);
xor UO_927 (O_927,N_14177,N_13396);
or UO_928 (O_928,N_14439,N_13676);
nand UO_929 (O_929,N_13220,N_14820);
nor UO_930 (O_930,N_13965,N_12225);
nand UO_931 (O_931,N_13745,N_12541);
nand UO_932 (O_932,N_14425,N_14759);
or UO_933 (O_933,N_11560,N_11134);
or UO_934 (O_934,N_12017,N_12141);
or UO_935 (O_935,N_12507,N_12953);
or UO_936 (O_936,N_12503,N_11206);
or UO_937 (O_937,N_11732,N_13823);
xor UO_938 (O_938,N_14225,N_10649);
nand UO_939 (O_939,N_13065,N_13155);
xor UO_940 (O_940,N_14049,N_12426);
nor UO_941 (O_941,N_13894,N_10897);
nor UO_942 (O_942,N_14888,N_11853);
and UO_943 (O_943,N_13617,N_12696);
nand UO_944 (O_944,N_13937,N_13625);
or UO_945 (O_945,N_14580,N_13675);
nand UO_946 (O_946,N_13785,N_11896);
or UO_947 (O_947,N_13799,N_14162);
or UO_948 (O_948,N_10608,N_14505);
and UO_949 (O_949,N_10881,N_14747);
and UO_950 (O_950,N_13540,N_10505);
xor UO_951 (O_951,N_12341,N_10817);
nand UO_952 (O_952,N_12248,N_12673);
nand UO_953 (O_953,N_10925,N_10627);
xnor UO_954 (O_954,N_10463,N_14156);
and UO_955 (O_955,N_11714,N_14958);
nand UO_956 (O_956,N_10684,N_14821);
xnor UO_957 (O_957,N_11299,N_11633);
xnor UO_958 (O_958,N_14516,N_12115);
nand UO_959 (O_959,N_13170,N_14946);
and UO_960 (O_960,N_12782,N_11979);
or UO_961 (O_961,N_12540,N_10434);
and UO_962 (O_962,N_14558,N_14627);
xor UO_963 (O_963,N_11711,N_11934);
and UO_964 (O_964,N_11598,N_13866);
nand UO_965 (O_965,N_13698,N_12967);
and UO_966 (O_966,N_13387,N_11503);
nor UO_967 (O_967,N_11489,N_10548);
nor UO_968 (O_968,N_14719,N_10617);
nor UO_969 (O_969,N_11479,N_10747);
nor UO_970 (O_970,N_13238,N_14589);
or UO_971 (O_971,N_11224,N_11345);
xor UO_972 (O_972,N_12823,N_12379);
nor UO_973 (O_973,N_11593,N_11132);
nand UO_974 (O_974,N_14731,N_10698);
and UO_975 (O_975,N_11328,N_10615);
xnor UO_976 (O_976,N_12234,N_10234);
and UO_977 (O_977,N_13332,N_10090);
nor UO_978 (O_978,N_12285,N_14403);
and UO_979 (O_979,N_10276,N_12022);
and UO_980 (O_980,N_10700,N_10635);
nand UO_981 (O_981,N_14274,N_13571);
and UO_982 (O_982,N_10361,N_14402);
nand UO_983 (O_983,N_12146,N_10614);
or UO_984 (O_984,N_10239,N_12435);
and UO_985 (O_985,N_11515,N_10400);
or UO_986 (O_986,N_12857,N_13306);
and UO_987 (O_987,N_10374,N_14118);
nor UO_988 (O_988,N_11940,N_11807);
xnor UO_989 (O_989,N_12775,N_14305);
nor UO_990 (O_990,N_12232,N_14793);
and UO_991 (O_991,N_10210,N_10816);
and UO_992 (O_992,N_12270,N_10761);
and UO_993 (O_993,N_10230,N_12236);
and UO_994 (O_994,N_11162,N_12004);
and UO_995 (O_995,N_12555,N_11822);
xnor UO_996 (O_996,N_12638,N_13460);
nor UO_997 (O_997,N_14381,N_12565);
and UO_998 (O_998,N_12760,N_13021);
xnor UO_999 (O_999,N_12394,N_13989);
and UO_1000 (O_1000,N_11608,N_13662);
xor UO_1001 (O_1001,N_14779,N_12527);
nor UO_1002 (O_1002,N_11952,N_10974);
xnor UO_1003 (O_1003,N_14853,N_10203);
nand UO_1004 (O_1004,N_11903,N_11867);
and UO_1005 (O_1005,N_13015,N_14351);
nand UO_1006 (O_1006,N_11542,N_14825);
xor UO_1007 (O_1007,N_12957,N_10358);
xor UO_1008 (O_1008,N_10814,N_10876);
xor UO_1009 (O_1009,N_13902,N_13849);
xor UO_1010 (O_1010,N_14060,N_10835);
or UO_1011 (O_1011,N_14008,N_13337);
and UO_1012 (O_1012,N_10233,N_14151);
nor UO_1013 (O_1013,N_10187,N_14257);
nand UO_1014 (O_1014,N_13865,N_11400);
nand UO_1015 (O_1015,N_14838,N_14899);
or UO_1016 (O_1016,N_11856,N_13827);
or UO_1017 (O_1017,N_12879,N_11279);
nor UO_1018 (O_1018,N_13151,N_12940);
or UO_1019 (O_1019,N_14307,N_13858);
xnor UO_1020 (O_1020,N_13315,N_13503);
nor UO_1021 (O_1021,N_13489,N_11731);
or UO_1022 (O_1022,N_14390,N_12177);
nor UO_1023 (O_1023,N_13046,N_14124);
or UO_1024 (O_1024,N_13504,N_12578);
or UO_1025 (O_1025,N_11225,N_11627);
or UO_1026 (O_1026,N_12567,N_11320);
nand UO_1027 (O_1027,N_12536,N_14004);
and UO_1028 (O_1028,N_14756,N_11655);
or UO_1029 (O_1029,N_10432,N_11973);
or UO_1030 (O_1030,N_12904,N_14723);
nor UO_1031 (O_1031,N_10798,N_12590);
nand UO_1032 (O_1032,N_12984,N_12867);
nor UO_1033 (O_1033,N_12886,N_10634);
xnor UO_1034 (O_1034,N_12434,N_10095);
xnor UO_1035 (O_1035,N_13566,N_10385);
xnor UO_1036 (O_1036,N_11463,N_14281);
nand UO_1037 (O_1037,N_11223,N_13735);
nand UO_1038 (O_1038,N_14421,N_13413);
or UO_1039 (O_1039,N_10258,N_10760);
nor UO_1040 (O_1040,N_14349,N_12784);
and UO_1041 (O_1041,N_14202,N_13509);
and UO_1042 (O_1042,N_12646,N_10500);
or UO_1043 (O_1043,N_10011,N_13717);
nand UO_1044 (O_1044,N_13990,N_14780);
nand UO_1045 (O_1045,N_14537,N_11352);
nand UO_1046 (O_1046,N_13602,N_11805);
nor UO_1047 (O_1047,N_11370,N_10215);
nor UO_1048 (O_1048,N_10074,N_12486);
nand UO_1049 (O_1049,N_11718,N_10337);
and UO_1050 (O_1050,N_14822,N_13630);
or UO_1051 (O_1051,N_13322,N_13000);
xnor UO_1052 (O_1052,N_14524,N_13179);
nand UO_1053 (O_1053,N_13470,N_11519);
nor UO_1054 (O_1054,N_10279,N_12143);
nor UO_1055 (O_1055,N_11114,N_10546);
nand UO_1056 (O_1056,N_13531,N_12806);
nor UO_1057 (O_1057,N_14328,N_11015);
xor UO_1058 (O_1058,N_10803,N_11618);
xnor UO_1059 (O_1059,N_13040,N_10065);
xnor UO_1060 (O_1060,N_14383,N_13940);
nor UO_1061 (O_1061,N_13175,N_11938);
or UO_1062 (O_1062,N_10324,N_12575);
and UO_1063 (O_1063,N_11106,N_13945);
nand UO_1064 (O_1064,N_12214,N_10541);
or UO_1065 (O_1065,N_10671,N_10934);
xnor UO_1066 (O_1066,N_14318,N_10538);
nor UO_1067 (O_1067,N_12291,N_13292);
or UO_1068 (O_1068,N_13517,N_14562);
xnor UO_1069 (O_1069,N_14548,N_12125);
nand UO_1070 (O_1070,N_12948,N_12622);
and UO_1071 (O_1071,N_14874,N_14229);
nand UO_1072 (O_1072,N_12261,N_14695);
nor UO_1073 (O_1073,N_14145,N_10868);
and UO_1074 (O_1074,N_14833,N_10536);
and UO_1075 (O_1075,N_13983,N_10384);
nand UO_1076 (O_1076,N_12991,N_12238);
xnor UO_1077 (O_1077,N_11296,N_13143);
nand UO_1078 (O_1078,N_13060,N_14434);
nand UO_1079 (O_1079,N_11882,N_10310);
xnor UO_1080 (O_1080,N_10291,N_11506);
nand UO_1081 (O_1081,N_14526,N_14643);
xnor UO_1082 (O_1082,N_14577,N_14968);
nand UO_1083 (O_1083,N_11422,N_12244);
or UO_1084 (O_1084,N_14898,N_14261);
nor UO_1085 (O_1085,N_14186,N_11823);
or UO_1086 (O_1086,N_10928,N_14829);
nor UO_1087 (O_1087,N_13933,N_12241);
and UO_1088 (O_1088,N_10594,N_10751);
nor UO_1089 (O_1089,N_11836,N_13130);
nor UO_1090 (O_1090,N_12355,N_13383);
and UO_1091 (O_1091,N_10893,N_14090);
nand UO_1092 (O_1092,N_13820,N_14034);
nand UO_1093 (O_1093,N_12465,N_12561);
nor UO_1094 (O_1094,N_13844,N_13316);
or UO_1095 (O_1095,N_10732,N_12905);
nand UO_1096 (O_1096,N_13775,N_12210);
and UO_1097 (O_1097,N_11755,N_13944);
and UO_1098 (O_1098,N_13808,N_10101);
xor UO_1099 (O_1099,N_10949,N_14510);
xnor UO_1100 (O_1100,N_12255,N_11672);
and UO_1101 (O_1101,N_13573,N_11029);
or UO_1102 (O_1102,N_12679,N_11857);
nand UO_1103 (O_1103,N_11844,N_13740);
xor UO_1104 (O_1104,N_14398,N_13869);
nor UO_1105 (O_1105,N_14845,N_13758);
nand UO_1106 (O_1106,N_11763,N_13772);
and UO_1107 (O_1107,N_11143,N_13020);
and UO_1108 (O_1108,N_12339,N_13518);
nand UO_1109 (O_1109,N_10852,N_11659);
nand UO_1110 (O_1110,N_11362,N_14830);
and UO_1111 (O_1111,N_14581,N_14647);
and UO_1112 (O_1112,N_13683,N_13027);
or UO_1113 (O_1113,N_11174,N_14468);
xor UO_1114 (O_1114,N_13207,N_13922);
xnor UO_1115 (O_1115,N_11446,N_10405);
nand UO_1116 (O_1116,N_11325,N_10185);
and UO_1117 (O_1117,N_13555,N_10655);
nand UO_1118 (O_1118,N_10148,N_14818);
nand UO_1119 (O_1119,N_11902,N_10901);
xnor UO_1120 (O_1120,N_14783,N_12340);
nor UO_1121 (O_1121,N_13275,N_11859);
xnor UO_1122 (O_1122,N_14427,N_13893);
nand UO_1123 (O_1123,N_12610,N_12716);
nor UO_1124 (O_1124,N_10993,N_14364);
and UO_1125 (O_1125,N_12147,N_12375);
nand UO_1126 (O_1126,N_14333,N_11850);
or UO_1127 (O_1127,N_13608,N_12807);
nand UO_1128 (O_1128,N_12088,N_11022);
nor UO_1129 (O_1129,N_14930,N_13487);
nand UO_1130 (O_1130,N_10448,N_10398);
nand UO_1131 (O_1131,N_12395,N_10563);
or UO_1132 (O_1132,N_10317,N_11656);
nand UO_1133 (O_1133,N_10861,N_10642);
xor UO_1134 (O_1134,N_14775,N_13248);
nand UO_1135 (O_1135,N_10809,N_12990);
nor UO_1136 (O_1136,N_10756,N_11947);
and UO_1137 (O_1137,N_13276,N_12155);
nand UO_1138 (O_1138,N_14545,N_12941);
nor UO_1139 (O_1139,N_10031,N_11835);
or UO_1140 (O_1140,N_11557,N_11742);
and UO_1141 (O_1141,N_14291,N_14496);
xnor UO_1142 (O_1142,N_10701,N_10629);
or UO_1143 (O_1143,N_11815,N_12294);
or UO_1144 (O_1144,N_13741,N_13881);
nor UO_1145 (O_1145,N_11438,N_13381);
nor UO_1146 (O_1146,N_13807,N_12733);
or UO_1147 (O_1147,N_13333,N_12385);
nor UO_1148 (O_1148,N_14104,N_11617);
nor UO_1149 (O_1149,N_12054,N_14216);
xnor UO_1150 (O_1150,N_12648,N_12211);
or UO_1151 (O_1151,N_14244,N_13359);
or UO_1152 (O_1152,N_10872,N_11564);
xor UO_1153 (O_1153,N_10729,N_10715);
and UO_1154 (O_1154,N_14591,N_10680);
and UO_1155 (O_1155,N_14702,N_14768);
nor UO_1156 (O_1156,N_11071,N_14811);
nor UO_1157 (O_1157,N_12698,N_12692);
and UO_1158 (O_1158,N_12049,N_14881);
or UO_1159 (O_1159,N_10019,N_11283);
nand UO_1160 (O_1160,N_13265,N_14959);
nor UO_1161 (O_1161,N_11484,N_14322);
or UO_1162 (O_1162,N_10945,N_14593);
or UO_1163 (O_1163,N_14761,N_13877);
nor UO_1164 (O_1164,N_11588,N_14389);
nand UO_1165 (O_1165,N_12419,N_14325);
nand UO_1166 (O_1166,N_14334,N_12287);
nor UO_1167 (O_1167,N_14882,N_12647);
nor UO_1168 (O_1168,N_12405,N_10349);
and UO_1169 (O_1169,N_13927,N_11986);
and UO_1170 (O_1170,N_11594,N_12048);
xnor UO_1171 (O_1171,N_10636,N_13549);
nand UO_1172 (O_1172,N_14507,N_14614);
nand UO_1173 (O_1173,N_13462,N_12520);
or UO_1174 (O_1174,N_10362,N_11285);
nor UO_1175 (O_1175,N_11214,N_10298);
xnor UO_1176 (O_1176,N_10592,N_11485);
or UO_1177 (O_1177,N_10468,N_13498);
and UO_1178 (O_1178,N_13097,N_11562);
nor UO_1179 (O_1179,N_12367,N_13034);
or UO_1180 (O_1180,N_10379,N_10573);
nand UO_1181 (O_1181,N_11757,N_12186);
nand UO_1182 (O_1182,N_13092,N_14868);
nand UO_1183 (O_1183,N_11910,N_14152);
nand UO_1184 (O_1184,N_11113,N_13002);
xnor UO_1185 (O_1185,N_14331,N_12068);
nand UO_1186 (O_1186,N_13915,N_12836);
xor UO_1187 (O_1187,N_12123,N_12396);
nand UO_1188 (O_1188,N_10706,N_11331);
nand UO_1189 (O_1189,N_11827,N_11522);
nand UO_1190 (O_1190,N_14555,N_10639);
nand UO_1191 (O_1191,N_11297,N_10863);
and UO_1192 (O_1192,N_14061,N_13296);
nor UO_1193 (O_1193,N_12554,N_13585);
xnor UO_1194 (O_1194,N_13913,N_11241);
nand UO_1195 (O_1195,N_10209,N_10954);
and UO_1196 (O_1196,N_13848,N_13030);
or UO_1197 (O_1197,N_10589,N_11874);
and UO_1198 (O_1198,N_11073,N_11335);
xor UO_1199 (O_1199,N_10718,N_10165);
or UO_1200 (O_1200,N_12138,N_10376);
and UO_1201 (O_1201,N_10360,N_13274);
and UO_1202 (O_1202,N_11540,N_10139);
xor UO_1203 (O_1203,N_11975,N_12970);
nand UO_1204 (O_1204,N_11623,N_13673);
and UO_1205 (O_1205,N_10826,N_10099);
nand UO_1206 (O_1206,N_13371,N_12249);
or UO_1207 (O_1207,N_11780,N_14210);
nor UO_1208 (O_1208,N_12746,N_12844);
or UO_1209 (O_1209,N_14560,N_12264);
nand UO_1210 (O_1210,N_11338,N_10871);
and UO_1211 (O_1211,N_10695,N_14317);
nand UO_1212 (O_1212,N_14326,N_10838);
or UO_1213 (O_1213,N_13632,N_13939);
nor UO_1214 (O_1214,N_14975,N_10855);
or UO_1215 (O_1215,N_11155,N_13336);
or UO_1216 (O_1216,N_13303,N_12873);
and UO_1217 (O_1217,N_14697,N_11819);
xnor UO_1218 (O_1218,N_10392,N_14940);
xor UO_1219 (O_1219,N_14712,N_13114);
xor UO_1220 (O_1220,N_10476,N_13273);
xnor UO_1221 (O_1221,N_12779,N_13613);
or UO_1222 (O_1222,N_10137,N_12918);
and UO_1223 (O_1223,N_11361,N_10504);
and UO_1224 (O_1224,N_13776,N_10417);
or UO_1225 (O_1225,N_10936,N_14990);
and UO_1226 (O_1226,N_10813,N_10619);
and UO_1227 (O_1227,N_11635,N_14750);
nand UO_1228 (O_1228,N_11526,N_10686);
nand UO_1229 (O_1229,N_10021,N_14343);
xnor UO_1230 (O_1230,N_11640,N_13384);
or UO_1231 (O_1231,N_14661,N_13284);
nand UO_1232 (O_1232,N_14538,N_12612);
and UO_1233 (O_1233,N_11498,N_13326);
nand UO_1234 (O_1234,N_11704,N_10981);
nor UO_1235 (O_1235,N_11967,N_13861);
and UO_1236 (O_1236,N_10188,N_14769);
or UO_1237 (O_1237,N_10982,N_11769);
nand UO_1238 (O_1238,N_12033,N_11381);
and UO_1239 (O_1239,N_12830,N_12751);
and UO_1240 (O_1240,N_13804,N_14587);
or UO_1241 (O_1241,N_13351,N_11675);
nand UO_1242 (O_1242,N_14418,N_10217);
nor UO_1243 (O_1243,N_14159,N_10260);
and UO_1244 (O_1244,N_11866,N_12256);
nand UO_1245 (O_1245,N_12314,N_14354);
and UO_1246 (O_1246,N_13255,N_14823);
xnor UO_1247 (O_1247,N_10428,N_13106);
or UO_1248 (O_1248,N_10490,N_13221);
xnor UO_1249 (O_1249,N_10205,N_13871);
nor UO_1250 (O_1250,N_12203,N_10150);
xor UO_1251 (O_1251,N_14278,N_14462);
xor UO_1252 (O_1252,N_12749,N_12658);
nor UO_1253 (O_1253,N_11215,N_13147);
and UO_1254 (O_1254,N_14673,N_12748);
nor UO_1255 (O_1255,N_13969,N_11124);
xnor UO_1256 (O_1256,N_12400,N_11079);
and UO_1257 (O_1257,N_10032,N_13066);
xnor UO_1258 (O_1258,N_11441,N_13657);
and UO_1259 (O_1259,N_11469,N_14858);
nor UO_1260 (O_1260,N_11348,N_10471);
nor UO_1261 (O_1261,N_13750,N_13560);
or UO_1262 (O_1262,N_13875,N_12768);
or UO_1263 (O_1263,N_13962,N_14189);
nor UO_1264 (O_1264,N_13133,N_11610);
nor UO_1265 (O_1265,N_12178,N_12719);
nor UO_1266 (O_1266,N_10196,N_14480);
or UO_1267 (O_1267,N_12464,N_12165);
and UO_1268 (O_1268,N_14934,N_11260);
and UO_1269 (O_1269,N_10231,N_13656);
or UO_1270 (O_1270,N_14806,N_14954);
nand UO_1271 (O_1271,N_11472,N_14644);
and UO_1272 (O_1272,N_10397,N_10766);
and UO_1273 (O_1273,N_11488,N_14443);
or UO_1274 (O_1274,N_12902,N_10163);
nor UO_1275 (O_1275,N_12135,N_11777);
nand UO_1276 (O_1276,N_12543,N_14522);
xnor UO_1277 (O_1277,N_12882,N_14010);
and UO_1278 (O_1278,N_14835,N_11310);
xor UO_1279 (O_1279,N_10092,N_11821);
nor UO_1280 (O_1280,N_13138,N_10155);
nand UO_1281 (O_1281,N_13450,N_11521);
nor UO_1282 (O_1282,N_14042,N_10818);
and UO_1283 (O_1283,N_14911,N_11356);
and UO_1284 (O_1284,N_12327,N_12566);
nor UO_1285 (O_1285,N_14329,N_11546);
nand UO_1286 (O_1286,N_14730,N_10801);
nor UO_1287 (O_1287,N_13240,N_10123);
nand UO_1288 (O_1288,N_14021,N_10348);
nor UO_1289 (O_1289,N_11081,N_13290);
xor UO_1290 (O_1290,N_13975,N_10225);
xor UO_1291 (O_1291,N_13637,N_13590);
or UO_1292 (O_1292,N_10763,N_12860);
nand UO_1293 (O_1293,N_10653,N_14301);
nor UO_1294 (O_1294,N_14618,N_11445);
and UO_1295 (O_1295,N_13925,N_10625);
and UO_1296 (O_1296,N_11052,N_10244);
or UO_1297 (O_1297,N_13725,N_11570);
and UO_1298 (O_1298,N_13693,N_13132);
and UO_1299 (O_1299,N_10606,N_12358);
nor UO_1300 (O_1300,N_13538,N_12601);
nor UO_1301 (O_1301,N_12714,N_13223);
xnor UO_1302 (O_1302,N_11912,N_12179);
nand UO_1303 (O_1303,N_14588,N_13081);
xnor UO_1304 (O_1304,N_14188,N_13584);
nand UO_1305 (O_1305,N_13241,N_14464);
nor UO_1306 (O_1306,N_11662,N_14138);
or UO_1307 (O_1307,N_13377,N_14684);
or UO_1308 (O_1308,N_11963,N_12707);
xor UO_1309 (O_1309,N_10339,N_12005);
xnor UO_1310 (O_1310,N_13722,N_10771);
or UO_1311 (O_1311,N_13601,N_12684);
and UO_1312 (O_1312,N_14409,N_10363);
or UO_1313 (O_1313,N_11774,N_10313);
xnor UO_1314 (O_1314,N_14099,N_13713);
xor UO_1315 (O_1315,N_10787,N_11746);
or UO_1316 (O_1316,N_11553,N_10393);
or UO_1317 (O_1317,N_10299,N_13052);
xnor UO_1318 (O_1318,N_13314,N_14309);
xnor UO_1319 (O_1319,N_12079,N_12013);
nor UO_1320 (O_1320,N_13778,N_14687);
nor UO_1321 (O_1321,N_13916,N_11737);
nor UO_1322 (O_1322,N_10721,N_10282);
nand UO_1323 (O_1323,N_13706,N_12537);
nor UO_1324 (O_1324,N_13088,N_12711);
and UO_1325 (O_1325,N_12382,N_10938);
or UO_1326 (O_1326,N_12848,N_13405);
nor UO_1327 (O_1327,N_13379,N_12180);
nand UO_1328 (O_1328,N_13004,N_10060);
nor UO_1329 (O_1329,N_10862,N_12799);
and UO_1330 (O_1330,N_14324,N_13508);
nor UO_1331 (O_1331,N_12336,N_13631);
xor UO_1332 (O_1332,N_14612,N_10610);
and UO_1333 (O_1333,N_11378,N_11723);
nor UO_1334 (O_1334,N_14782,N_10178);
or UO_1335 (O_1335,N_12193,N_11467);
xnor UO_1336 (O_1336,N_12801,N_12114);
nand UO_1337 (O_1337,N_10462,N_14107);
nor UO_1338 (O_1338,N_14147,N_10331);
and UO_1339 (O_1339,N_10560,N_10005);
nor UO_1340 (O_1340,N_12473,N_11354);
and UO_1341 (O_1341,N_11665,N_14121);
xor UO_1342 (O_1342,N_11911,N_11292);
xnor UO_1343 (O_1343,N_14969,N_14062);
or UO_1344 (O_1344,N_11394,N_12427);
and UO_1345 (O_1345,N_11049,N_12333);
or UO_1346 (O_1346,N_12067,N_13488);
nand UO_1347 (O_1347,N_10808,N_11991);
xnor UO_1348 (O_1348,N_11341,N_10888);
and UO_1349 (O_1349,N_12308,N_10886);
nor UO_1350 (O_1350,N_10149,N_12350);
or UO_1351 (O_1351,N_11609,N_10704);
and UO_1352 (O_1352,N_14636,N_12871);
or UO_1353 (O_1353,N_10256,N_10764);
and UO_1354 (O_1354,N_10961,N_11877);
and UO_1355 (O_1355,N_14226,N_14413);
nand UO_1356 (O_1356,N_13817,N_14422);
nor UO_1357 (O_1357,N_13753,N_13821);
nor UO_1358 (O_1358,N_13859,N_14036);
and UO_1359 (O_1359,N_11061,N_12690);
and UO_1360 (O_1360,N_11793,N_13468);
and UO_1361 (O_1361,N_14852,N_11929);
or UO_1362 (O_1362,N_13272,N_11527);
nor UO_1363 (O_1363,N_14277,N_11854);
nand UO_1364 (O_1364,N_12204,N_13621);
or UO_1365 (O_1365,N_12785,N_10869);
xor UO_1366 (O_1366,N_11591,N_11581);
or UO_1367 (O_1367,N_13124,N_13233);
and UO_1368 (O_1368,N_12983,N_12505);
nor UO_1369 (O_1369,N_11889,N_13960);
nand UO_1370 (O_1370,N_10288,N_13449);
nor UO_1371 (O_1371,N_12757,N_13353);
or UO_1372 (O_1372,N_11326,N_14966);
xor UO_1373 (O_1373,N_13679,N_13897);
and UO_1374 (O_1374,N_13228,N_11698);
nand UO_1375 (O_1375,N_12345,N_11865);
nor UO_1376 (O_1376,N_11669,N_11514);
nor UO_1377 (O_1377,N_12704,N_13599);
or UO_1378 (O_1378,N_14486,N_11243);
xnor UO_1379 (O_1379,N_11663,N_10598);
xnor UO_1380 (O_1380,N_13734,N_11628);
xor UO_1381 (O_1381,N_12269,N_10856);
or UO_1382 (O_1382,N_11772,N_14865);
nor UO_1383 (O_1383,N_12511,N_10983);
or UO_1384 (O_1384,N_10411,N_10980);
or UO_1385 (O_1385,N_14504,N_10736);
nor UO_1386 (O_1386,N_12364,N_12265);
nand UO_1387 (O_1387,N_14999,N_10903);
nand UO_1388 (O_1388,N_11160,N_14448);
and UO_1389 (O_1389,N_11578,N_11586);
or UO_1390 (O_1390,N_11554,N_14441);
xor UO_1391 (O_1391,N_11808,N_11631);
nor UO_1392 (O_1392,N_12788,N_13059);
xnor UO_1393 (O_1393,N_10724,N_14044);
xor UO_1394 (O_1394,N_10014,N_12743);
nand UO_1395 (O_1395,N_10488,N_12428);
nor UO_1396 (O_1396,N_13553,N_14310);
xor UO_1397 (O_1397,N_10117,N_10344);
nand UO_1398 (O_1398,N_12240,N_10786);
and UO_1399 (O_1399,N_11030,N_11202);
nor UO_1400 (O_1400,N_13469,N_12869);
or UO_1401 (O_1401,N_14250,N_10714);
nand UO_1402 (O_1402,N_14455,N_14921);
nand UO_1403 (O_1403,N_14981,N_11630);
and UO_1404 (O_1404,N_13611,N_13973);
nor UO_1405 (O_1405,N_13319,N_14860);
or UO_1406 (O_1406,N_12303,N_11995);
or UO_1407 (O_1407,N_12360,N_12001);
or UO_1408 (O_1408,N_11621,N_13195);
nand UO_1409 (O_1409,N_10378,N_12192);
and UO_1410 (O_1410,N_10316,N_13230);
and UO_1411 (O_1411,N_12454,N_12614);
nand UO_1412 (O_1412,N_14533,N_13215);
nor UO_1413 (O_1413,N_12042,N_12965);
nand UO_1414 (O_1414,N_11996,N_11685);
or UO_1415 (O_1415,N_13152,N_11064);
xnor UO_1416 (O_1416,N_14745,N_12188);
xnor UO_1417 (O_1417,N_10851,N_10754);
nor UO_1418 (O_1418,N_11596,N_14615);
xor UO_1419 (O_1419,N_12034,N_11738);
and UO_1420 (O_1420,N_11500,N_14623);
or UO_1421 (O_1421,N_10947,N_14474);
nor UO_1422 (O_1422,N_14863,N_11146);
xor UO_1423 (O_1423,N_13146,N_12818);
nor UO_1424 (O_1424,N_14795,N_12304);
nand UO_1425 (O_1425,N_14135,N_13728);
nand UO_1426 (O_1426,N_13682,N_14550);
xnor UO_1427 (O_1427,N_13198,N_12615);
and UO_1428 (O_1428,N_14265,N_13080);
xnor UO_1429 (O_1429,N_10281,N_13416);
and UO_1430 (O_1430,N_10638,N_14350);
xnor UO_1431 (O_1431,N_11303,N_10443);
nor UO_1432 (O_1432,N_14234,N_10252);
or UO_1433 (O_1433,N_13935,N_10268);
nor UO_1434 (O_1434,N_14617,N_12587);
or UO_1435 (O_1435,N_14701,N_12838);
or UO_1436 (O_1436,N_10419,N_10841);
nand UO_1437 (O_1437,N_10973,N_11683);
nand UO_1438 (O_1438,N_11333,N_13667);
nor UO_1439 (O_1439,N_13293,N_13609);
nand UO_1440 (O_1440,N_12051,N_14009);
and UO_1441 (O_1441,N_14339,N_12324);
xor UO_1442 (O_1442,N_13199,N_12354);
xnor UO_1443 (O_1443,N_10006,N_12812);
nor UO_1444 (O_1444,N_12073,N_13291);
nor UO_1445 (O_1445,N_12494,N_11783);
nor UO_1446 (O_1446,N_12538,N_13082);
nor UO_1447 (O_1447,N_12198,N_14998);
xnor UO_1448 (O_1448,N_13786,N_14323);
or UO_1449 (O_1449,N_10494,N_14199);
nor UO_1450 (O_1450,N_12603,N_13444);
and UO_1451 (O_1451,N_10875,N_14854);
or UO_1452 (O_1452,N_11237,N_14297);
and UO_1453 (O_1453,N_11210,N_11287);
and UO_1454 (O_1454,N_14503,N_14502);
nand UO_1455 (O_1455,N_13627,N_13409);
and UO_1456 (O_1456,N_13404,N_12586);
nor UO_1457 (O_1457,N_11308,N_11458);
nand UO_1458 (O_1458,N_11432,N_11038);
and UO_1459 (O_1459,N_10052,N_13596);
xnor UO_1460 (O_1460,N_12620,N_10367);
or UO_1461 (O_1461,N_10315,N_12346);
xor UO_1462 (O_1462,N_14051,N_12278);
xor UO_1463 (O_1463,N_13167,N_10289);
nor UO_1464 (O_1464,N_10902,N_12605);
or UO_1465 (O_1465,N_11198,N_14956);
and UO_1466 (O_1466,N_11573,N_13558);
nor UO_1467 (O_1467,N_11899,N_13695);
xnor UO_1468 (O_1468,N_13210,N_13923);
nand UO_1469 (O_1469,N_13671,N_12046);
or UO_1470 (O_1470,N_10273,N_13329);
and UO_1471 (O_1471,N_12140,N_11181);
and UO_1472 (O_1472,N_12031,N_10833);
nor UO_1473 (O_1473,N_10124,N_14864);
and UO_1474 (O_1474,N_10138,N_12205);
nor UO_1475 (O_1475,N_10164,N_10269);
and UO_1476 (O_1476,N_12632,N_14256);
or UO_1477 (O_1477,N_13654,N_13798);
xnor UO_1478 (O_1478,N_13642,N_11505);
xnor UO_1479 (O_1479,N_11460,N_13919);
nand UO_1480 (O_1480,N_14467,N_13115);
nor UO_1481 (O_1481,N_11706,N_14611);
or UO_1482 (O_1482,N_13550,N_12795);
or UO_1483 (O_1483,N_10264,N_11451);
or UO_1484 (O_1484,N_12451,N_12110);
or UO_1485 (O_1485,N_12894,N_12316);
xor UO_1486 (O_1486,N_12705,N_14404);
nor UO_1487 (O_1487,N_12392,N_11764);
nor UO_1488 (O_1488,N_11062,N_14412);
nand UO_1489 (O_1489,N_11199,N_13348);
xnor UO_1490 (O_1490,N_14032,N_11078);
and UO_1491 (O_1491,N_12829,N_10483);
xor UO_1492 (O_1492,N_13438,N_14201);
nor UO_1493 (O_1493,N_12721,N_14624);
xnor UO_1494 (O_1494,N_10136,N_11250);
nand UO_1495 (O_1495,N_13661,N_10911);
and UO_1496 (O_1496,N_14613,N_13453);
xor UO_1497 (O_1497,N_14895,N_11103);
xor UO_1498 (O_1498,N_13447,N_12041);
nand UO_1499 (O_1499,N_12408,N_10477);
and UO_1500 (O_1500,N_14120,N_13137);
nor UO_1501 (O_1501,N_13213,N_11371);
and UO_1502 (O_1502,N_10693,N_13696);
or UO_1503 (O_1503,N_14741,N_13077);
xor UO_1504 (O_1504,N_13525,N_14116);
xnor UO_1505 (O_1505,N_13282,N_10531);
nor UO_1506 (O_1506,N_12119,N_13522);
or UO_1507 (O_1507,N_14100,N_14178);
and UO_1508 (O_1508,N_13287,N_11213);
nor UO_1509 (O_1509,N_10858,N_11200);
nand UO_1510 (O_1510,N_11266,N_12223);
and UO_1511 (O_1511,N_11454,N_14924);
xor UO_1512 (O_1512,N_10955,N_13645);
or UO_1513 (O_1513,N_13045,N_12767);
nand UO_1514 (O_1514,N_11161,N_13885);
xor UO_1515 (O_1515,N_11367,N_12421);
and UO_1516 (O_1516,N_12640,N_11492);
and UO_1517 (O_1517,N_14483,N_14770);
or UO_1518 (O_1518,N_11674,N_13299);
xor UO_1519 (O_1519,N_10670,N_14625);
nor UO_1520 (O_1520,N_13985,N_12987);
xnor UO_1521 (O_1521,N_11217,N_12082);
nor UO_1522 (O_1522,N_10111,N_11121);
and UO_1523 (O_1523,N_10346,N_11372);
and UO_1524 (O_1524,N_13951,N_10612);
or UO_1525 (O_1525,N_14873,N_13966);
nor UO_1526 (O_1526,N_14908,N_10746);
nand UO_1527 (O_1527,N_11788,N_11673);
or UO_1528 (O_1528,N_13880,N_14897);
or UO_1529 (O_1529,N_13171,N_13458);
nand UO_1530 (O_1530,N_14109,N_14743);
nand UO_1531 (O_1531,N_11334,N_12794);
or UO_1532 (O_1532,N_11893,N_11565);
and UO_1533 (O_1533,N_12926,N_11138);
and UO_1534 (O_1534,N_11480,N_14757);
xor UO_1535 (O_1535,N_14708,N_11282);
and UO_1536 (O_1536,N_12378,N_11447);
and UO_1537 (O_1537,N_13997,N_11230);
nor UO_1538 (O_1538,N_14554,N_11486);
xor UO_1539 (O_1539,N_11473,N_14028);
and UO_1540 (O_1540,N_13655,N_12683);
and UO_1541 (O_1541,N_11909,N_12066);
nor UO_1542 (O_1542,N_13948,N_13892);
or UO_1543 (O_1543,N_10513,N_14665);
and UO_1544 (O_1544,N_10236,N_13545);
and UO_1545 (O_1545,N_12506,N_11234);
or UO_1546 (O_1546,N_10603,N_10184);
and UO_1547 (O_1547,N_14059,N_12351);
nor UO_1548 (O_1548,N_11701,N_12330);
nand UO_1549 (O_1549,N_11956,N_11703);
nand UO_1550 (O_1550,N_10918,N_13279);
nor UO_1551 (O_1551,N_11985,N_11318);
nor UO_1552 (O_1552,N_11531,N_12482);
xor UO_1553 (O_1553,N_14481,N_14482);
nand UO_1554 (O_1554,N_11900,N_12854);
nor UO_1555 (O_1555,N_13636,N_12952);
nor UO_1556 (O_1556,N_13181,N_13556);
nand UO_1557 (O_1557,N_10796,N_13312);
nor UO_1558 (O_1558,N_12352,N_10853);
and UO_1559 (O_1559,N_11123,N_11240);
or UO_1560 (O_1560,N_11016,N_12485);
or UO_1561 (O_1561,N_12070,N_11776);
nor UO_1562 (O_1562,N_10388,N_11734);
and UO_1563 (O_1563,N_12432,N_10887);
and UO_1564 (O_1564,N_10555,N_10682);
nor UO_1565 (O_1565,N_14063,N_13910);
xnor UO_1566 (O_1566,N_11722,N_12656);
nand UO_1567 (O_1567,N_13022,N_11743);
nor UO_1568 (O_1568,N_14271,N_14436);
and UO_1569 (O_1569,N_12501,N_10969);
and UO_1570 (O_1570,N_14224,N_13497);
xnor UO_1571 (O_1571,N_14259,N_13914);
or UO_1572 (O_1572,N_12423,N_11176);
and UO_1573 (O_1573,N_13575,N_13911);
nor UO_1574 (O_1574,N_14348,N_10043);
or UO_1575 (O_1575,N_11294,N_11236);
nor UO_1576 (O_1576,N_13057,N_11205);
and UO_1577 (O_1577,N_12744,N_13534);
or UO_1578 (O_1578,N_14846,N_13434);
nor UO_1579 (O_1579,N_13372,N_10740);
xor UO_1580 (O_1580,N_10058,N_11433);
or UO_1581 (O_1581,N_14395,N_13086);
or UO_1582 (O_1582,N_13506,N_13523);
xnor UO_1583 (O_1583,N_12676,N_11055);
or UO_1584 (O_1584,N_14810,N_13651);
nor UO_1585 (O_1585,N_12471,N_12126);
or UO_1586 (O_1586,N_10643,N_10564);
or UO_1587 (O_1587,N_11353,N_13051);
and UO_1588 (O_1588,N_10705,N_11105);
and UO_1589 (O_1589,N_13794,N_14893);
nand UO_1590 (O_1590,N_13901,N_12913);
xnor UO_1591 (O_1591,N_12962,N_14879);
and UO_1592 (O_1592,N_14153,N_11619);
nand UO_1593 (O_1593,N_11606,N_12842);
xor UO_1594 (O_1594,N_12710,N_13710);
or UO_1595 (O_1595,N_14532,N_14453);
and UO_1596 (O_1596,N_12233,N_13374);
and UO_1597 (O_1597,N_13305,N_10055);
nor UO_1598 (O_1598,N_14433,N_13380);
nor UO_1599 (O_1599,N_11065,N_13726);
and UO_1600 (O_1600,N_10551,N_11657);
nand UO_1601 (O_1601,N_11904,N_10927);
nand UO_1602 (O_1602,N_10620,N_10068);
nand UO_1603 (O_1603,N_14703,N_11535);
xor UO_1604 (O_1604,N_11920,N_14773);
nand UO_1605 (O_1605,N_13595,N_14664);
and UO_1606 (O_1606,N_13406,N_11405);
nand UO_1607 (O_1607,N_10520,N_14360);
or UO_1608 (O_1608,N_12372,N_10895);
xnor UO_1609 (O_1609,N_13295,N_14374);
and UO_1610 (O_1610,N_12044,N_11981);
nor UO_1611 (O_1611,N_10080,N_11607);
or UO_1612 (O_1612,N_12870,N_13987);
or UO_1613 (O_1613,N_10285,N_12754);
nand UO_1614 (O_1614,N_10020,N_14282);
xor UO_1615 (O_1615,N_10662,N_14827);
nor UO_1616 (O_1616,N_10191,N_14521);
nor UO_1617 (O_1617,N_14659,N_11890);
xor UO_1618 (O_1618,N_14236,N_13298);
nor UO_1619 (O_1619,N_10030,N_10070);
nand UO_1620 (O_1620,N_14861,N_11347);
nor UO_1621 (O_1621,N_10501,N_10218);
and UO_1622 (O_1622,N_13532,N_12043);
and UO_1623 (O_1623,N_12936,N_11869);
nor UO_1624 (O_1624,N_13283,N_10088);
xnor UO_1625 (O_1625,N_14520,N_12160);
and UO_1626 (O_1626,N_12985,N_13988);
and UO_1627 (O_1627,N_12740,N_10581);
or UO_1628 (O_1628,N_12018,N_13455);
xnor UO_1629 (O_1629,N_12661,N_11122);
xor UO_1630 (O_1630,N_13582,N_12722);
xnor UO_1631 (O_1631,N_13102,N_10597);
or UO_1632 (O_1632,N_12583,N_12973);
nor UO_1633 (O_1633,N_10450,N_13770);
nand UO_1634 (O_1634,N_10637,N_12460);
and UO_1635 (O_1635,N_12669,N_12846);
nand UO_1636 (O_1636,N_14878,N_13410);
xor UO_1637 (O_1637,N_12334,N_14254);
nor UO_1638 (O_1638,N_12220,N_12579);
nor UO_1639 (O_1639,N_13388,N_12545);
xor UO_1640 (O_1640,N_10839,N_14230);
nor UO_1641 (O_1641,N_14556,N_13472);
nor UO_1642 (O_1642,N_11790,N_11165);
or UO_1643 (O_1643,N_11142,N_12399);
nand UO_1644 (O_1644,N_14417,N_11110);
xor UO_1645 (O_1645,N_14551,N_11647);
xnor UO_1646 (O_1646,N_10917,N_12935);
xnor UO_1647 (O_1647,N_11977,N_10473);
xor UO_1648 (O_1648,N_11615,N_13186);
xnor UO_1649 (O_1649,N_11694,N_10460);
xnor UO_1650 (O_1650,N_10783,N_14943);
or UO_1651 (O_1651,N_12359,N_14228);
xor UO_1652 (O_1652,N_11196,N_11369);
nand UO_1653 (O_1653,N_11887,N_11377);
and UO_1654 (O_1654,N_10034,N_10152);
and UO_1655 (O_1655,N_11024,N_14289);
xnor UO_1656 (O_1656,N_13818,N_13873);
nand UO_1657 (O_1657,N_11086,N_12514);
nor UO_1658 (O_1658,N_10255,N_13140);
and UO_1659 (O_1659,N_14253,N_12533);
or UO_1660 (O_1660,N_13056,N_11392);
and UO_1661 (O_1661,N_13759,N_14103);
nand UO_1662 (O_1662,N_13075,N_11388);
and UO_1663 (O_1663,N_10284,N_13790);
and UO_1664 (O_1664,N_10057,N_10556);
xnor UO_1665 (O_1665,N_11448,N_10590);
nor UO_1666 (O_1666,N_12910,N_14025);
or UO_1667 (O_1667,N_12502,N_12134);
and UO_1668 (O_1668,N_13828,N_12023);
nor UO_1669 (O_1669,N_13036,N_14985);
and UO_1670 (O_1670,N_10733,N_11091);
and UO_1671 (O_1671,N_11906,N_10580);
nor UO_1672 (O_1672,N_14442,N_10944);
nand UO_1673 (O_1673,N_12349,N_11528);
or UO_1674 (O_1674,N_13703,N_10194);
and UO_1675 (O_1675,N_14038,N_11875);
and UO_1676 (O_1676,N_10528,N_13536);
nand UO_1677 (O_1677,N_13370,N_10208);
nand UO_1678 (O_1678,N_11574,N_12449);
nand UO_1679 (O_1679,N_14859,N_11888);
and UO_1680 (O_1680,N_12243,N_10819);
nor UO_1681 (O_1681,N_13653,N_12616);
and UO_1682 (O_1682,N_14052,N_11307);
or UO_1683 (O_1683,N_13882,N_10051);
and UO_1684 (O_1684,N_13483,N_10707);
or UO_1685 (O_1685,N_11457,N_10946);
or UO_1686 (O_1686,N_10830,N_13345);
nand UO_1687 (O_1687,N_14748,N_11153);
xnor UO_1688 (O_1688,N_14758,N_14362);
nand UO_1689 (O_1689,N_14435,N_14696);
nand UO_1690 (O_1690,N_10272,N_12104);
nor UO_1691 (O_1691,N_14227,N_10905);
and UO_1692 (O_1692,N_12835,N_13278);
and UO_1693 (O_1693,N_14050,N_10121);
and UO_1694 (O_1694,N_10601,N_14014);
nand UO_1695 (O_1695,N_14791,N_14406);
xor UO_1696 (O_1696,N_11475,N_12332);
and UO_1697 (O_1697,N_11087,N_10914);
or UO_1698 (O_1698,N_12376,N_11558);
nor UO_1699 (O_1699,N_14699,N_14469);
and UO_1700 (O_1700,N_14071,N_12441);
nand UO_1701 (O_1701,N_13109,N_10569);
nand UO_1702 (O_1702,N_12461,N_13355);
nand UO_1703 (O_1703,N_10979,N_10335);
xnor UO_1704 (O_1704,N_12318,N_10271);
or UO_1705 (O_1705,N_10485,N_12804);
nand UO_1706 (O_1706,N_13003,N_13979);
or UO_1707 (O_1707,N_12015,N_12895);
nor UO_1708 (O_1708,N_12920,N_13635);
xnor UO_1709 (O_1709,N_12230,N_14706);
or UO_1710 (O_1710,N_10010,N_11314);
nand UO_1711 (O_1711,N_14630,N_14501);
or UO_1712 (O_1712,N_13846,N_14262);
xnor UO_1713 (O_1713,N_10492,N_13507);
nand UO_1714 (O_1714,N_11666,N_13070);
nor UO_1715 (O_1715,N_11516,N_11837);
and UO_1716 (O_1716,N_13007,N_12824);
nor UO_1717 (O_1717,N_10482,N_13764);
nand UO_1718 (O_1718,N_12950,N_12262);
and UO_1719 (O_1719,N_13938,N_13712);
or UO_1720 (O_1720,N_14073,N_12509);
and UO_1721 (O_1721,N_13104,N_14338);
or UO_1722 (O_1722,N_10668,N_13111);
xor UO_1723 (O_1723,N_12994,N_13446);
or UO_1724 (O_1724,N_10469,N_11077);
or UO_1725 (O_1725,N_11194,N_11517);
and UO_1726 (O_1726,N_13593,N_11304);
xnor UO_1727 (O_1727,N_13862,N_11375);
or UO_1728 (O_1728,N_12130,N_14129);
nor UO_1729 (O_1729,N_11754,N_10297);
xor UO_1730 (O_1730,N_13459,N_13286);
nand UO_1731 (O_1731,N_14473,N_10266);
nor UO_1732 (O_1732,N_12859,N_12534);
or UO_1733 (O_1733,N_12564,N_14451);
and UO_1734 (O_1734,N_12281,N_13451);
or UO_1735 (O_1735,N_14964,N_12000);
and UO_1736 (O_1736,N_12556,N_12833);
nand UO_1737 (O_1737,N_13998,N_13194);
nor UO_1738 (O_1738,N_12039,N_12828);
and UO_1739 (O_1739,N_13084,N_11332);
and UO_1740 (O_1740,N_12157,N_11496);
and UO_1741 (O_1741,N_12317,N_11932);
nand UO_1742 (O_1742,N_13161,N_10293);
nor UO_1743 (O_1743,N_12753,N_13204);
xor UO_1744 (O_1744,N_11109,N_12845);
nand UO_1745 (O_1745,N_12252,N_14031);
or UO_1746 (O_1746,N_10042,N_13500);
and UO_1747 (O_1747,N_11756,N_14802);
nor UO_1748 (O_1748,N_11705,N_12499);
xor UO_1749 (O_1749,N_14191,N_10913);
and UO_1750 (O_1750,N_12144,N_10193);
or UO_1751 (O_1751,N_14527,N_12809);
nor UO_1752 (O_1752,N_13974,N_12212);
or UO_1753 (O_1753,N_10883,N_12325);
nand UO_1754 (O_1754,N_13981,N_11994);
nand UO_1755 (O_1755,N_11592,N_14732);
xnor UO_1756 (O_1756,N_13906,N_10950);
nor UO_1757 (O_1757,N_14974,N_11948);
and UO_1758 (O_1758,N_10844,N_11154);
nor UO_1759 (O_1759,N_13830,N_12881);
nor UO_1760 (O_1760,N_11811,N_11715);
xnor UO_1761 (O_1761,N_12258,N_14368);
and UO_1762 (O_1762,N_10535,N_14399);
and UO_1763 (O_1763,N_11923,N_14214);
or UO_1764 (O_1764,N_11190,N_12604);
and UO_1765 (O_1765,N_13257,N_10765);
and UO_1766 (O_1766,N_10553,N_12477);
and UO_1767 (O_1767,N_14841,N_11684);
or UO_1768 (O_1768,N_11941,N_14055);
and UO_1769 (O_1769,N_11242,N_11892);
nor UO_1770 (O_1770,N_12899,N_10975);
nand UO_1771 (O_1771,N_12353,N_14925);
xor UO_1772 (O_1772,N_10478,N_14192);
nor UO_1773 (O_1773,N_11197,N_13777);
xnor UO_1774 (O_1774,N_11700,N_14912);
and UO_1775 (O_1775,N_12456,N_10403);
nor UO_1776 (O_1776,N_14347,N_11275);
and UO_1777 (O_1777,N_14536,N_14767);
nor UO_1778 (O_1778,N_14645,N_13176);
nor UO_1779 (O_1779,N_10224,N_10711);
xnor UO_1780 (O_1780,N_12643,N_12850);
xor UO_1781 (O_1781,N_11426,N_14141);
or UO_1782 (O_1782,N_13711,N_13932);
nand UO_1783 (O_1783,N_12593,N_12891);
nand UO_1784 (O_1784,N_10322,N_12094);
xor UO_1785 (O_1785,N_12552,N_11139);
xnor UO_1786 (O_1786,N_10059,N_13930);
nand UO_1787 (O_1787,N_11550,N_10514);
nand UO_1788 (O_1788,N_14180,N_12306);
and UO_1789 (O_1789,N_10248,N_12492);
and UO_1790 (O_1790,N_13921,N_11474);
nor UO_1791 (O_1791,N_11175,N_12518);
and UO_1792 (O_1792,N_10441,N_10442);
and UO_1793 (O_1793,N_11159,N_11385);
xor UO_1794 (O_1794,N_11148,N_12821);
nand UO_1795 (O_1795,N_13570,N_10822);
nor UO_1796 (O_1796,N_12508,N_12919);
or UO_1797 (O_1797,N_12780,N_11219);
and UO_1798 (O_1798,N_12771,N_13443);
or UO_1799 (O_1799,N_14799,N_12671);
and UO_1800 (O_1800,N_10182,N_13831);
nand UO_1801 (O_1801,N_10524,N_12609);
and UO_1802 (O_1802,N_13218,N_13530);
nand UO_1803 (O_1803,N_12407,N_10769);
nor UO_1804 (O_1804,N_13847,N_11871);
nand UO_1805 (O_1805,N_10728,N_12170);
and UO_1806 (O_1806,N_10086,N_12148);
xor UO_1807 (O_1807,N_10357,N_14877);
nand UO_1808 (O_1808,N_11654,N_12150);
nand UO_1809 (O_1809,N_13685,N_11818);
and UO_1810 (O_1810,N_10785,N_13993);
xor UO_1811 (O_1811,N_14694,N_13280);
nand UO_1812 (O_1812,N_14223,N_14933);
and UO_1813 (O_1813,N_10807,N_10602);
xor UO_1814 (O_1814,N_11051,N_10941);
nand UO_1815 (O_1815,N_13128,N_11629);
or UO_1816 (O_1816,N_12627,N_14294);
or UO_1817 (O_1817,N_10943,N_10160);
nor UO_1818 (O_1818,N_11043,N_11027);
nor UO_1819 (O_1819,N_13628,N_13598);
nand UO_1820 (O_1820,N_12161,N_10998);
or UO_1821 (O_1821,N_14634,N_10730);
xor UO_1822 (O_1822,N_14105,N_11945);
nand UO_1823 (O_1823,N_12348,N_14428);
and UO_1824 (O_1824,N_10829,N_13192);
nand UO_1825 (O_1825,N_11997,N_10660);
nand UO_1826 (O_1826,N_11220,N_10354);
or UO_1827 (O_1827,N_12883,N_12581);
and UO_1828 (O_1828,N_10557,N_10007);
or UO_1829 (O_1829,N_12847,N_11070);
nand UO_1830 (O_1830,N_14869,N_14635);
xnor UO_1831 (O_1831,N_10235,N_12585);
and UO_1832 (O_1832,N_14494,N_12322);
nand UO_1833 (O_1833,N_12288,N_12010);
and UO_1834 (O_1834,N_12443,N_10791);
nand UO_1835 (O_1835,N_11418,N_14967);
or UO_1836 (O_1836,N_11127,N_10096);
and UO_1837 (O_1837,N_14938,N_14619);
nand UO_1838 (O_1838,N_12741,N_13492);
or UO_1839 (O_1839,N_12172,N_13991);
xor UO_1840 (O_1840,N_12369,N_10585);
nand UO_1841 (O_1841,N_12761,N_10377);
or UO_1842 (O_1842,N_13529,N_11649);
or UO_1843 (O_1843,N_14622,N_11962);
nor UO_1844 (O_1844,N_12971,N_13313);
xnor UO_1845 (O_1845,N_14553,N_13955);
or UO_1846 (O_1846,N_13403,N_14995);
nand UO_1847 (O_1847,N_14366,N_12852);
nor UO_1848 (O_1848,N_11549,N_11974);
nand UO_1849 (O_1849,N_13554,N_10028);
nand UO_1850 (O_1850,N_14570,N_12686);
nor UO_1851 (O_1851,N_14792,N_14207);
nand UO_1852 (O_1852,N_10734,N_14649);
nor UO_1853 (O_1853,N_11133,N_13014);
xnor UO_1854 (O_1854,N_14016,N_14245);
or UO_1855 (O_1855,N_12472,N_12487);
nand UO_1856 (O_1856,N_11244,N_13486);
nor UO_1857 (O_1857,N_12978,N_10716);
and UO_1858 (O_1858,N_10894,N_11935);
or UO_1859 (O_1859,N_13072,N_11009);
and UO_1860 (O_1860,N_12938,N_10831);
or UO_1861 (O_1861,N_12132,N_13644);
nand UO_1862 (O_1862,N_10578,N_13567);
xnor UO_1863 (O_1863,N_12467,N_11256);
nor UO_1864 (O_1864,N_12065,N_12976);
and UO_1865 (O_1865,N_13024,N_14492);
nand UO_1866 (O_1866,N_12272,N_10154);
and UO_1867 (O_1867,N_13268,N_12813);
and UO_1868 (O_1868,N_12917,N_11309);
xor UO_1869 (O_1869,N_14026,N_11796);
and UO_1870 (O_1870,N_13401,N_13665);
nor UO_1871 (O_1871,N_13771,N_14583);
nor UO_1872 (O_1872,N_13150,N_10532);
xnor UO_1873 (O_1873,N_11284,N_12329);
or UO_1874 (O_1874,N_12235,N_10709);
and UO_1875 (O_1875,N_14993,N_10290);
and UO_1876 (O_1876,N_11315,N_13061);
or UO_1877 (O_1877,N_13876,N_14922);
and UO_1878 (O_1878,N_11466,N_11825);
nand UO_1879 (O_1879,N_11702,N_10810);
xor UO_1880 (O_1880,N_14672,N_12498);
nor UO_1881 (O_1881,N_13864,N_14190);
or UO_1882 (O_1882,N_11651,N_10053);
or UO_1883 (O_1883,N_11898,N_14816);
xor UO_1884 (O_1884,N_14332,N_13610);
or UO_1885 (O_1885,N_12458,N_12652);
and UO_1886 (O_1886,N_13622,N_10186);
nor UO_1887 (O_1887,N_13793,N_10084);
and UO_1888 (O_1888,N_11319,N_14197);
or UO_1889 (O_1889,N_11597,N_10142);
and UO_1890 (O_1890,N_11085,N_13648);
nand UO_1891 (O_1891,N_10795,N_10811);
or UO_1892 (O_1892,N_14509,N_14027);
xnor UO_1893 (O_1893,N_11416,N_10402);
xnor UO_1894 (O_1894,N_11075,N_14082);
nand UO_1895 (O_1895,N_11965,N_12221);
and UO_1896 (O_1896,N_14972,N_13742);
nand UO_1897 (O_1897,N_12750,N_11944);
or UO_1898 (O_1898,N_14179,N_11525);
or UO_1899 (O_1899,N_11100,N_13108);
nor UO_1900 (O_1900,N_10422,N_13259);
xor UO_1901 (O_1901,N_10588,N_12297);
or UO_1902 (O_1902,N_13418,N_14842);
nor UO_1903 (O_1903,N_10352,N_11355);
nor UO_1904 (O_1904,N_14660,N_10000);
xnor UO_1905 (O_1905,N_11692,N_13164);
and UO_1906 (O_1906,N_11571,N_12030);
or UO_1907 (O_1907,N_12805,N_12457);
or UO_1908 (O_1908,N_10898,N_14078);
nor UO_1909 (O_1909,N_12986,N_14176);
or UO_1910 (O_1910,N_14728,N_12735);
nor UO_1911 (O_1911,N_14991,N_12840);
nand UO_1912 (O_1912,N_13748,N_10063);
or UO_1913 (O_1913,N_10109,N_11845);
or UO_1914 (O_1914,N_10048,N_10078);
xnor UO_1915 (O_1915,N_14692,N_14127);
nor UO_1916 (O_1916,N_12681,N_10976);
xnor UO_1917 (O_1917,N_13294,N_14094);
nor UO_1918 (O_1918,N_14807,N_14638);
xnor UO_1919 (O_1919,N_13839,N_10016);
or UO_1920 (O_1920,N_11971,N_12613);
nor UO_1921 (O_1921,N_10416,N_11464);
or UO_1922 (O_1922,N_11697,N_10674);
or UO_1923 (O_1923,N_11440,N_13681);
nor UO_1924 (O_1924,N_12531,N_14184);
nand UO_1925 (O_1925,N_10677,N_14909);
and UO_1926 (O_1926,N_10665,N_11530);
nor UO_1927 (O_1927,N_14499,N_14710);
nand UO_1928 (O_1928,N_14169,N_12979);
xor UO_1929 (O_1929,N_12229,N_14819);
nand UO_1930 (O_1930,N_12189,N_12872);
xnor UO_1931 (O_1931,N_13816,N_13340);
xnor UO_1932 (O_1932,N_13718,N_14384);
nand UO_1933 (O_1933,N_13368,N_11135);
and UO_1934 (O_1934,N_11268,N_13903);
nor UO_1935 (O_1935,N_13076,N_12121);
nand UO_1936 (O_1936,N_13415,N_10859);
nand UO_1937 (O_1937,N_10758,N_12418);
and UO_1938 (O_1938,N_12406,N_11207);
or UO_1939 (O_1939,N_10699,N_13356);
or UO_1940 (O_1940,N_14415,N_14892);
or UO_1941 (O_1941,N_10308,N_11648);
nor UO_1942 (O_1942,N_11544,N_12090);
nand UO_1943 (O_1943,N_13658,N_13344);
nand UO_1944 (O_1944,N_10474,N_12071);
nor UO_1945 (O_1945,N_11419,N_12525);
nand UO_1946 (O_1946,N_11288,N_13791);
and UO_1947 (O_1947,N_12724,N_10958);
xor UO_1948 (O_1948,N_12422,N_12548);
nor UO_1949 (O_1949,N_13854,N_14206);
or UO_1950 (O_1950,N_10658,N_10202);
or UO_1951 (O_1951,N_11144,N_12103);
xnor UO_1952 (O_1952,N_10865,N_11012);
and UO_1953 (O_1953,N_14283,N_12549);
xnor UO_1954 (O_1954,N_10498,N_14165);
and UO_1955 (O_1955,N_13001,N_12436);
nand UO_1956 (O_1956,N_14267,N_11851);
nand UO_1957 (O_1957,N_14632,N_13535);
or UO_1958 (O_1958,N_14544,N_11927);
or UO_1959 (O_1959,N_13577,N_11864);
nand UO_1960 (O_1960,N_12504,N_13840);
nor UO_1961 (O_1961,N_12064,N_14880);
or UO_1962 (O_1962,N_14674,N_14007);
nor UO_1963 (O_1963,N_14198,N_12576);
and UO_1964 (O_1964,N_14087,N_10877);
or UO_1965 (O_1965,N_10568,N_14929);
xnor UO_1966 (O_1966,N_10607,N_14772);
nand UO_1967 (O_1967,N_11339,N_14790);
xor UO_1968 (O_1968,N_14466,N_14300);
or UO_1969 (O_1969,N_10181,N_13227);
and UO_1970 (O_1970,N_12491,N_12052);
xor UO_1971 (O_1971,N_12693,N_14602);
nor UO_1972 (O_1972,N_10004,N_12342);
and UO_1973 (O_1973,N_10050,N_14955);
nor UO_1974 (O_1974,N_13638,N_14495);
or UO_1975 (O_1975,N_14762,N_12680);
xnor UO_1976 (O_1976,N_10456,N_13216);
or UO_1977 (O_1977,N_11222,N_12495);
nand UO_1978 (O_1978,N_10664,N_13087);
xnor UO_1979 (O_1979,N_13049,N_12832);
xor UO_1980 (O_1980,N_12896,N_14675);
nor UO_1981 (O_1981,N_10604,N_13250);
xnor UO_1982 (O_1982,N_11168,N_10395);
xnor UO_1983 (O_1983,N_10192,N_14335);
and UO_1984 (O_1984,N_11936,N_10035);
and UO_1985 (O_1985,N_14139,N_12769);
nor UO_1986 (O_1986,N_10126,N_11620);
xnor UO_1987 (O_1987,N_14850,N_14847);
or UO_1988 (O_1988,N_13327,N_14251);
xor UO_1989 (O_1989,N_10788,N_13512);
xnor UO_1990 (O_1990,N_10093,N_12181);
nor UO_1991 (O_1991,N_12476,N_14506);
and UO_1992 (O_1992,N_13583,N_14727);
nor UO_1993 (O_1993,N_10630,N_10066);
and UO_1994 (O_1994,N_13597,N_10977);
or UO_1995 (O_1995,N_12397,N_12713);
nor UO_1996 (O_1996,N_13201,N_11539);
xnor UO_1997 (O_1997,N_11172,N_14755);
or UO_1998 (O_1998,N_10966,N_11235);
xor UO_1999 (O_1999,N_14393,N_13005);
endmodule