module basic_1500_15000_2000_100_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_183,In_244);
and U1 (N_1,In_1411,In_1132);
and U2 (N_2,In_1106,In_1139);
or U3 (N_3,In_630,In_616);
nor U4 (N_4,In_1112,In_323);
nor U5 (N_5,In_225,In_1170);
nor U6 (N_6,In_800,In_1074);
xnor U7 (N_7,In_9,In_1012);
or U8 (N_8,In_1459,In_1396);
or U9 (N_9,In_125,In_1449);
xnor U10 (N_10,In_1160,In_1444);
nand U11 (N_11,In_1379,In_1473);
or U12 (N_12,In_881,In_474);
nand U13 (N_13,In_1025,In_992);
nand U14 (N_14,In_1265,In_1127);
and U15 (N_15,In_1356,In_1469);
xor U16 (N_16,In_946,In_708);
xor U17 (N_17,In_1344,In_637);
xnor U18 (N_18,In_589,In_1261);
nand U19 (N_19,In_1306,In_1425);
or U20 (N_20,In_1092,In_473);
nand U21 (N_21,In_306,In_245);
nor U22 (N_22,In_1000,In_704);
xor U23 (N_23,In_1117,In_203);
or U24 (N_24,In_22,In_810);
and U25 (N_25,In_300,In_1295);
nand U26 (N_26,In_724,In_903);
xor U27 (N_27,In_251,In_858);
nand U28 (N_28,In_135,In_866);
or U29 (N_29,In_837,In_877);
nand U30 (N_30,In_108,In_1381);
or U31 (N_31,In_618,In_1049);
nor U32 (N_32,In_897,In_404);
nor U33 (N_33,In_268,In_1213);
xor U34 (N_34,In_884,In_665);
nor U35 (N_35,In_257,In_1457);
or U36 (N_36,In_845,In_408);
nand U37 (N_37,In_243,In_1342);
nand U38 (N_38,In_185,In_202);
nand U39 (N_39,In_147,In_171);
nor U40 (N_40,In_158,In_1308);
and U41 (N_41,In_1079,In_77);
or U42 (N_42,In_718,In_663);
or U43 (N_43,In_673,In_821);
nor U44 (N_44,In_740,In_462);
xor U45 (N_45,In_624,In_458);
nand U46 (N_46,In_487,In_649);
and U47 (N_47,In_594,In_33);
nand U48 (N_48,In_882,In_685);
xnor U49 (N_49,In_1369,In_1383);
nor U50 (N_50,In_689,In_394);
and U51 (N_51,In_1169,In_1482);
or U52 (N_52,In_892,In_842);
or U53 (N_53,In_94,In_558);
and U54 (N_54,In_502,In_274);
or U55 (N_55,In_525,In_1210);
nand U56 (N_56,In_1455,In_1208);
xnor U57 (N_57,In_678,In_1357);
and U58 (N_58,In_1174,In_153);
xnor U59 (N_59,In_868,In_1224);
nand U60 (N_60,In_175,In_1249);
nand U61 (N_61,In_859,In_57);
nor U62 (N_62,In_167,In_51);
xor U63 (N_63,In_517,In_709);
or U64 (N_64,In_1115,In_824);
and U65 (N_65,In_1282,In_1027);
xnor U66 (N_66,In_1166,In_694);
and U67 (N_67,In_475,In_217);
or U68 (N_68,In_1119,In_179);
and U69 (N_69,In_733,In_381);
nand U70 (N_70,In_1107,In_1296);
or U71 (N_71,In_345,In_855);
nor U72 (N_72,In_1240,In_47);
nand U73 (N_73,In_1104,In_976);
nor U74 (N_74,In_344,In_1076);
nor U75 (N_75,In_1194,In_602);
nand U76 (N_76,In_834,In_500);
nand U77 (N_77,In_1320,In_1402);
nor U78 (N_78,In_294,In_39);
and U79 (N_79,In_55,In_1324);
xor U80 (N_80,In_65,In_785);
and U81 (N_81,In_929,In_645);
nor U82 (N_82,In_468,In_852);
nand U83 (N_83,In_1195,In_1314);
nor U84 (N_84,In_1051,In_974);
nor U85 (N_85,In_849,In_1321);
xor U86 (N_86,In_794,In_1388);
or U87 (N_87,In_118,In_383);
and U88 (N_88,In_8,In_4);
and U89 (N_89,In_945,In_1220);
or U90 (N_90,In_72,In_352);
nor U91 (N_91,In_1405,In_601);
and U92 (N_92,In_1052,In_226);
xor U93 (N_93,In_36,In_885);
nand U94 (N_94,In_690,In_769);
and U95 (N_95,In_119,In_1399);
or U96 (N_96,In_819,In_947);
nand U97 (N_97,In_1222,In_755);
and U98 (N_98,In_1175,In_1346);
or U99 (N_99,In_1315,In_625);
nand U100 (N_100,In_1142,In_1275);
and U101 (N_101,In_1136,In_870);
or U102 (N_102,In_1196,In_73);
or U103 (N_103,In_1319,In_95);
xnor U104 (N_104,In_1281,In_194);
and U105 (N_105,In_1363,In_1452);
nand U106 (N_106,In_100,In_682);
xor U107 (N_107,In_1071,In_792);
nor U108 (N_108,In_122,In_638);
and U109 (N_109,In_1125,In_389);
and U110 (N_110,In_1023,In_596);
nand U111 (N_111,In_1239,In_538);
or U112 (N_112,In_980,In_715);
xor U113 (N_113,In_287,In_1029);
nor U114 (N_114,In_1011,In_409);
nor U115 (N_115,In_104,In_219);
xnor U116 (N_116,In_937,In_1272);
nand U117 (N_117,In_1299,In_727);
nor U118 (N_118,In_1391,In_944);
or U119 (N_119,In_480,In_58);
nor U120 (N_120,In_857,In_295);
xor U121 (N_121,In_363,In_451);
xor U122 (N_122,In_743,In_791);
nand U123 (N_123,In_1232,In_803);
and U124 (N_124,In_901,In_968);
and U125 (N_125,In_511,In_989);
nand U126 (N_126,In_30,In_1135);
xnor U127 (N_127,In_84,In_1191);
nor U128 (N_128,In_1002,In_959);
nand U129 (N_129,In_271,In_811);
nor U130 (N_130,In_53,In_1318);
and U131 (N_131,In_918,In_1128);
nor U132 (N_132,In_843,In_1149);
nand U133 (N_133,In_397,In_1058);
or U134 (N_134,In_664,In_463);
and U135 (N_135,In_442,In_181);
or U136 (N_136,In_1365,In_303);
nor U137 (N_137,In_1325,In_1268);
nor U138 (N_138,In_1032,In_776);
xnor U139 (N_139,In_1255,In_499);
xor U140 (N_140,In_1096,In_1326);
and U141 (N_141,In_321,In_1097);
xor U142 (N_142,In_477,In_1351);
or U143 (N_143,In_437,In_304);
nand U144 (N_144,In_711,In_120);
nor U145 (N_145,In_269,In_1233);
and U146 (N_146,In_1089,In_256);
and U147 (N_147,In_342,In_129);
xor U148 (N_148,In_60,In_206);
xor U149 (N_149,In_1088,In_176);
or U150 (N_150,In_1412,N_122);
xnor U151 (N_151,In_1018,In_748);
and U152 (N_152,N_69,In_461);
and U153 (N_153,In_433,In_695);
nor U154 (N_154,N_114,In_301);
xor U155 (N_155,In_1392,In_1238);
nor U156 (N_156,In_924,In_12);
nand U157 (N_157,In_305,In_1488);
nand U158 (N_158,In_871,In_1433);
nand U159 (N_159,In_479,In_164);
or U160 (N_160,In_156,In_913);
nor U161 (N_161,In_778,In_320);
and U162 (N_162,N_111,In_1364);
nand U163 (N_163,In_334,In_117);
and U164 (N_164,N_123,In_80);
and U165 (N_165,In_1118,In_1350);
nand U166 (N_166,In_888,In_424);
nand U167 (N_167,In_936,In_1108);
nor U168 (N_168,N_121,N_9);
nor U169 (N_169,In_1204,In_1207);
xor U170 (N_170,In_191,In_34);
nand U171 (N_171,In_13,In_841);
nor U172 (N_172,In_756,In_988);
nor U173 (N_173,In_597,In_1200);
nor U174 (N_174,In_1426,In_1167);
nand U175 (N_175,In_428,In_403);
xor U176 (N_176,In_1361,N_74);
xnor U177 (N_177,In_735,In_132);
and U178 (N_178,In_873,In_939);
nand U179 (N_179,In_1487,In_780);
nand U180 (N_180,In_832,In_288);
and U181 (N_181,N_55,In_137);
or U182 (N_182,In_338,In_264);
nor U183 (N_183,In_1436,In_311);
and U184 (N_184,In_1349,In_82);
nand U185 (N_185,In_1010,In_1408);
xor U186 (N_186,In_643,In_999);
nor U187 (N_187,In_10,In_1151);
nand U188 (N_188,In_448,N_102);
and U189 (N_189,In_703,In_143);
nor U190 (N_190,In_1086,In_1285);
xor U191 (N_191,In_591,In_169);
nand U192 (N_192,In_1267,In_355);
and U193 (N_193,In_1277,In_1338);
or U194 (N_194,N_106,In_1456);
nand U195 (N_195,In_166,In_5);
and U196 (N_196,In_152,In_476);
or U197 (N_197,N_43,In_354);
xnor U198 (N_198,In_292,In_1085);
xor U199 (N_199,In_606,In_554);
xnor U200 (N_200,In_542,In_688);
nand U201 (N_201,In_116,In_184);
and U202 (N_202,In_247,N_145);
nand U203 (N_203,In_353,In_1385);
nor U204 (N_204,In_457,In_343);
nor U205 (N_205,In_1384,In_1448);
xor U206 (N_206,N_139,In_729);
or U207 (N_207,In_46,In_782);
nor U208 (N_208,In_1123,In_1378);
and U209 (N_209,In_291,In_1437);
or U210 (N_210,N_44,In_450);
or U211 (N_211,In_779,In_1303);
nand U212 (N_212,In_380,In_406);
and U213 (N_213,In_28,In_145);
nand U214 (N_214,In_531,In_719);
nor U215 (N_215,In_81,In_585);
nor U216 (N_216,In_1226,In_812);
or U217 (N_217,In_1243,In_981);
nor U218 (N_218,In_922,In_620);
or U219 (N_219,In_214,N_67);
xnor U220 (N_220,In_931,In_805);
and U221 (N_221,In_1141,In_497);
nand U222 (N_222,In_734,In_809);
nor U223 (N_223,In_421,In_721);
nand U224 (N_224,In_1442,In_1218);
and U225 (N_225,In_1409,In_580);
nor U226 (N_226,In_1091,In_236);
or U227 (N_227,In_1276,In_1398);
or U228 (N_228,In_252,In_1168);
nand U229 (N_229,N_78,In_1090);
nor U230 (N_230,In_765,N_113);
xor U231 (N_231,In_420,In_17);
nand U232 (N_232,In_485,In_1131);
or U233 (N_233,In_1126,In_674);
nor U234 (N_234,In_905,N_103);
xnor U235 (N_235,In_199,In_712);
xor U236 (N_236,In_16,In_192);
or U237 (N_237,In_547,In_851);
or U238 (N_238,N_141,In_1355);
or U239 (N_239,In_366,In_237);
and U240 (N_240,In_211,In_666);
nand U241 (N_241,In_445,In_259);
nor U242 (N_242,In_109,In_784);
nand U243 (N_243,In_19,In_1259);
and U244 (N_244,In_846,In_1020);
and U245 (N_245,In_651,In_599);
and U246 (N_246,In_1026,In_182);
and U247 (N_247,In_59,In_565);
or U248 (N_248,N_22,In_341);
nor U249 (N_249,In_1087,In_1376);
nand U250 (N_250,In_911,In_98);
and U251 (N_251,In_262,In_1143);
nor U252 (N_252,In_446,In_969);
or U253 (N_253,In_97,In_371);
xnor U254 (N_254,In_1305,In_1124);
and U255 (N_255,In_503,In_1424);
xnor U256 (N_256,N_136,In_1337);
or U257 (N_257,In_1254,In_1245);
nand U258 (N_258,N_30,N_133);
nand U259 (N_259,In_524,In_700);
or U260 (N_260,In_1215,In_1247);
nor U261 (N_261,In_230,N_81);
nor U262 (N_262,In_646,In_1221);
or U263 (N_263,In_1418,In_56);
or U264 (N_264,In_906,In_965);
and U265 (N_265,In_826,In_796);
nor U266 (N_266,In_483,In_1333);
xnor U267 (N_267,N_134,In_279);
nand U268 (N_268,In_830,In_655);
and U269 (N_269,N_34,In_933);
xor U270 (N_270,In_557,In_818);
xor U271 (N_271,In_544,In_504);
or U272 (N_272,In_506,In_575);
and U273 (N_273,In_520,In_942);
nor U274 (N_274,In_608,In_569);
xnor U275 (N_275,In_904,In_1084);
nor U276 (N_276,In_45,In_1390);
nand U277 (N_277,In_701,In_379);
and U278 (N_278,In_1386,In_280);
nand U279 (N_279,In_836,In_435);
and U280 (N_280,In_1438,In_1317);
xnor U281 (N_281,In_1045,In_860);
xor U282 (N_282,In_691,In_86);
or U283 (N_283,N_116,In_405);
or U284 (N_284,In_32,In_996);
nor U285 (N_285,In_1053,In_1419);
nor U286 (N_286,N_10,In_510);
nor U287 (N_287,In_107,In_1256);
nor U288 (N_288,In_814,In_1188);
or U289 (N_289,In_31,In_952);
nor U290 (N_290,In_114,In_697);
or U291 (N_291,In_26,In_197);
or U292 (N_292,In_854,In_322);
xor U293 (N_293,In_1371,In_1329);
nor U294 (N_294,In_481,In_1447);
nand U295 (N_295,In_178,In_1274);
nand U296 (N_296,In_261,In_478);
and U297 (N_297,In_607,In_926);
xnor U298 (N_298,In_258,In_85);
and U299 (N_299,In_789,In_1147);
nor U300 (N_300,In_1206,In_1380);
xor U301 (N_301,In_1202,In_742);
nor U302 (N_302,N_28,In_207);
nand U303 (N_303,In_533,In_272);
xnor U304 (N_304,N_19,N_222);
and U305 (N_305,In_393,N_14);
xnor U306 (N_306,In_401,N_87);
nand U307 (N_307,In_168,In_1056);
nand U308 (N_308,In_741,In_509);
xor U309 (N_309,N_184,N_161);
and U310 (N_310,In_297,In_1260);
xor U311 (N_311,In_1273,In_1009);
and U312 (N_312,In_359,N_205);
or U313 (N_313,In_1185,N_197);
and U314 (N_314,In_263,In_610);
nand U315 (N_315,In_489,In_1284);
and U316 (N_316,N_202,N_267);
or U317 (N_317,N_278,In_1182);
nor U318 (N_318,In_339,N_129);
xor U319 (N_319,In_357,In_1413);
nand U320 (N_320,N_214,N_181);
and U321 (N_321,In_177,In_1495);
xor U322 (N_322,In_447,In_1158);
xnor U323 (N_323,In_633,In_62);
or U324 (N_324,In_1110,N_235);
and U325 (N_325,N_144,In_1353);
nand U326 (N_326,In_1030,In_516);
or U327 (N_327,In_987,In_693);
nand U328 (N_328,In_1493,N_112);
nand U329 (N_329,In_1193,In_96);
or U330 (N_330,In_308,N_33);
nand U331 (N_331,In_932,In_365);
nor U332 (N_332,In_1366,In_1022);
or U333 (N_333,In_282,In_698);
or U334 (N_334,In_1263,N_109);
nand U335 (N_335,N_173,In_1162);
and U336 (N_336,In_326,N_176);
nor U337 (N_337,In_686,N_277);
and U338 (N_338,In_970,N_26);
xor U339 (N_339,In_180,In_1257);
or U340 (N_340,In_925,N_292);
and U341 (N_341,In_210,In_1328);
or U342 (N_342,In_190,In_1001);
nor U343 (N_343,In_385,In_982);
xnor U344 (N_344,In_975,In_1013);
nand U345 (N_345,In_2,In_1031);
nand U346 (N_346,N_46,In_1393);
and U347 (N_347,In_1187,In_1227);
nand U348 (N_348,N_269,In_1146);
nand U349 (N_349,N_63,In_699);
and U350 (N_350,In_1377,In_254);
nor U351 (N_351,In_1330,In_640);
nor U352 (N_352,N_140,In_998);
nand U353 (N_353,In_66,In_731);
or U354 (N_354,In_1462,N_204);
nand U355 (N_355,In_609,In_161);
or U356 (N_356,In_1061,In_1081);
or U357 (N_357,N_50,In_351);
nor U358 (N_358,In_201,In_1434);
or U359 (N_359,In_1184,In_253);
nand U360 (N_360,In_49,In_233);
nor U361 (N_361,In_1427,In_684);
nor U362 (N_362,In_255,In_1464);
nand U363 (N_363,N_12,In_325);
or U364 (N_364,In_757,In_564);
or U365 (N_365,In_419,N_51);
xor U366 (N_366,In_612,In_1498);
and U367 (N_367,In_1102,In_89);
nand U368 (N_368,In_1279,In_537);
xor U369 (N_369,In_1219,In_1490);
and U370 (N_370,In_774,In_893);
nor U371 (N_371,N_230,N_45);
nand U372 (N_372,In_250,In_908);
xor U373 (N_373,In_839,N_201);
nor U374 (N_374,N_36,In_160);
xnor U375 (N_375,N_165,N_89);
xor U376 (N_376,In_1161,In_88);
xnor U377 (N_377,In_1179,In_472);
nor U378 (N_378,In_1105,In_221);
xnor U379 (N_379,In_386,In_1217);
or U380 (N_380,In_577,In_1038);
xor U381 (N_381,In_567,In_1252);
and U382 (N_382,In_187,In_27);
xnor U383 (N_383,In_398,In_1152);
xnor U384 (N_384,In_650,In_657);
and U385 (N_385,In_910,In_880);
and U386 (N_386,In_1080,N_15);
or U387 (N_387,In_848,In_101);
and U388 (N_388,In_286,In_349);
nand U389 (N_389,In_1294,In_647);
nor U390 (N_390,In_598,In_1138);
nand U391 (N_391,In_92,In_1075);
nor U392 (N_392,In_370,In_1236);
nand U393 (N_393,In_212,In_555);
and U394 (N_394,In_1121,In_1304);
xor U395 (N_395,In_1323,In_1015);
nor U396 (N_396,N_142,In_990);
and U397 (N_397,In_486,In_890);
nor U398 (N_398,In_1465,In_1432);
nor U399 (N_399,In_795,In_953);
and U400 (N_400,N_156,In_1262);
and U401 (N_401,N_261,In_293);
nand U402 (N_402,In_1302,In_1316);
nand U403 (N_403,In_804,In_1098);
xor U404 (N_404,In_508,In_915);
xor U405 (N_405,In_979,N_166);
and U406 (N_406,In_621,N_0);
and U407 (N_407,In_676,N_17);
or U408 (N_408,In_1485,In_592);
nand U409 (N_409,N_296,In_1439);
xor U410 (N_410,In_1415,In_559);
nor U411 (N_411,In_1060,N_180);
or U412 (N_412,In_896,N_243);
xor U413 (N_413,N_266,In_1034);
or U414 (N_414,In_1069,In_1486);
and U415 (N_415,In_613,In_1291);
or U416 (N_416,In_1230,N_248);
and U417 (N_417,In_717,In_328);
nand U418 (N_418,N_276,In_781);
xor U419 (N_419,In_204,In_955);
and U420 (N_420,In_1,In_148);
and U421 (N_421,In_441,In_928);
and U422 (N_422,In_963,In_856);
nor U423 (N_423,In_1101,N_287);
and U424 (N_424,In_984,In_566);
nor U425 (N_425,In_879,In_275);
xor U426 (N_426,N_242,In_7);
nor U427 (N_427,In_1040,In_1460);
xnor U428 (N_428,In_368,In_1078);
nor U429 (N_429,In_923,In_775);
nand U430 (N_430,In_593,N_117);
or U431 (N_431,In_422,In_1209);
nor U432 (N_432,In_1407,N_7);
or U433 (N_433,In_916,In_302);
nand U434 (N_434,N_273,In_1470);
nor U435 (N_435,N_71,In_1150);
and U436 (N_436,In_669,In_1293);
or U437 (N_437,In_138,In_822);
and U438 (N_438,N_32,In_526);
nand U439 (N_439,In_631,In_900);
or U440 (N_440,In_281,In_865);
xor U441 (N_441,N_164,In_746);
nand U442 (N_442,In_840,N_208);
xnor U443 (N_443,In_1387,N_211);
or U444 (N_444,N_147,In_494);
or U445 (N_445,In_798,In_154);
xor U446 (N_446,N_29,In_872);
and U447 (N_447,In_1290,In_747);
and U448 (N_448,In_861,In_25);
or U449 (N_449,In_490,In_707);
xor U450 (N_450,N_322,N_88);
or U451 (N_451,N_346,In_431);
or U452 (N_452,N_97,In_456);
and U453 (N_453,In_1421,N_76);
xor U454 (N_454,In_1375,In_831);
nand U455 (N_455,In_1441,In_1480);
and U456 (N_456,N_213,In_467);
xor U457 (N_457,In_1019,N_355);
nand U458 (N_458,In_330,In_808);
xor U459 (N_459,N_256,N_254);
or U460 (N_460,In_1120,N_232);
nor U461 (N_461,In_1389,In_1394);
nor U462 (N_462,In_1400,N_372);
nor U463 (N_463,In_315,N_227);
nand U464 (N_464,In_802,In_553);
or U465 (N_465,In_1177,In_788);
xnor U466 (N_466,In_276,N_75);
nand U467 (N_467,In_1403,N_146);
nor U468 (N_468,N_61,In_318);
nor U469 (N_469,In_1159,In_1322);
nand U470 (N_470,In_960,N_415);
nand U471 (N_471,In_20,N_56);
or U472 (N_472,In_1467,In_548);
nand U473 (N_473,In_1095,N_6);
or U474 (N_474,N_384,In_1474);
nand U475 (N_475,In_1137,In_290);
xnor U476 (N_476,N_163,In_964);
nor U477 (N_477,In_83,N_110);
nand U478 (N_478,In_1178,In_806);
and U479 (N_479,In_1410,N_271);
and U480 (N_480,N_21,N_259);
and U481 (N_481,In_227,In_862);
and U482 (N_482,N_420,In_954);
and U483 (N_483,In_636,In_1258);
nand U484 (N_484,In_622,N_439);
nor U485 (N_485,In_163,N_253);
nor U486 (N_486,In_360,In_87);
and U487 (N_487,In_1054,N_65);
nor U488 (N_488,N_421,In_130);
xor U489 (N_489,In_402,N_336);
and U490 (N_490,In_215,In_738);
xnor U491 (N_491,In_1203,In_412);
xnor U492 (N_492,In_745,In_127);
nand U493 (N_493,In_1401,N_335);
xnor U494 (N_494,In_93,N_189);
xnor U495 (N_495,In_78,In_1198);
and U496 (N_496,In_519,In_744);
xor U497 (N_497,In_1417,In_847);
and U498 (N_498,In_453,In_298);
nor U499 (N_499,In_772,N_127);
nand U500 (N_500,N_35,In_1047);
nand U501 (N_501,N_203,In_157);
nand U502 (N_502,In_1163,In_1360);
and U503 (N_503,N_412,In_240);
or U504 (N_504,In_1140,N_304);
xor U505 (N_505,In_1310,N_316);
xnor U506 (N_506,In_466,In_766);
and U507 (N_507,In_799,In_1343);
and U508 (N_508,N_158,In_390);
and U509 (N_509,In_737,In_777);
and U510 (N_510,In_174,N_247);
or U511 (N_511,N_334,In_828);
or U512 (N_512,In_1471,N_151);
nand U513 (N_513,N_290,N_52);
and U514 (N_514,In_310,N_285);
nand U515 (N_515,N_200,In_995);
or U516 (N_516,In_552,In_1099);
nor U517 (N_517,In_751,In_1494);
and U518 (N_518,N_101,N_178);
nand U519 (N_519,In_1481,In_681);
or U520 (N_520,In_895,In_1046);
or U521 (N_521,In_619,In_920);
xor U522 (N_522,N_375,In_867);
or U523 (N_523,In_425,N_130);
xor U524 (N_524,In_69,N_274);
nor U525 (N_525,In_962,In_823);
and U526 (N_526,In_407,In_496);
nor U527 (N_527,N_347,In_1043);
nand U528 (N_528,In_1345,In_1055);
and U529 (N_529,In_1133,N_91);
xor U530 (N_530,N_143,N_233);
and U531 (N_531,In_1212,In_570);
and U532 (N_532,In_875,In_1327);
nor U533 (N_533,In_563,N_2);
or U534 (N_534,N_342,In_605);
nor U535 (N_535,In_21,N_1);
or U536 (N_536,In_313,N_358);
xor U537 (N_537,In_455,In_102);
nor U538 (N_538,In_752,In_79);
and U539 (N_539,In_978,In_835);
nor U540 (N_540,In_518,In_316);
or U541 (N_541,In_151,In_242);
nand U542 (N_542,N_215,N_193);
nor U543 (N_543,In_115,In_535);
xor U544 (N_544,N_137,In_54);
and U545 (N_545,In_340,N_308);
xor U546 (N_546,N_337,In_1271);
or U547 (N_547,In_1339,N_206);
nor U548 (N_548,N_169,In_1048);
nand U549 (N_549,In_324,N_24);
and U550 (N_550,In_1173,N_226);
nand U551 (N_551,In_1443,In_1241);
or U552 (N_552,In_536,N_360);
nand U553 (N_553,In_1154,In_541);
nor U554 (N_554,N_385,In_1109);
nor U555 (N_555,In_1033,In_68);
xnor U556 (N_556,In_1180,N_446);
and U557 (N_557,N_218,In_1156);
nand U558 (N_558,In_377,In_238);
and U559 (N_559,N_90,N_60);
nand U560 (N_560,In_329,In_193);
nand U561 (N_561,N_170,In_1103);
or U562 (N_562,In_941,In_725);
xnor U563 (N_563,In_522,In_850);
and U564 (N_564,N_223,N_400);
or U565 (N_565,In_427,In_1445);
nor U566 (N_566,N_219,In_764);
nor U567 (N_567,In_556,In_582);
xnor U568 (N_568,N_83,In_1348);
xor U569 (N_569,In_1063,In_319);
xnor U570 (N_570,In_387,In_1017);
or U571 (N_571,N_57,In_1359);
or U572 (N_572,In_417,In_208);
nor U573 (N_573,N_80,N_321);
nand U574 (N_574,In_722,N_298);
xor U575 (N_575,N_120,N_220);
xor U576 (N_576,N_185,In_829);
xor U577 (N_577,In_951,N_96);
and U578 (N_578,N_159,In_587);
and U579 (N_579,In_560,N_245);
nor U580 (N_580,In_444,In_1111);
or U581 (N_581,In_144,N_234);
nor U582 (N_582,N_329,In_35);
nand U583 (N_583,In_392,N_3);
or U584 (N_584,In_648,In_1354);
or U585 (N_585,N_198,In_1430);
xnor U586 (N_586,N_179,In_90);
and U587 (N_587,In_696,In_838);
xor U588 (N_588,N_419,In_99);
or U589 (N_589,N_333,N_403);
and U590 (N_590,In_914,In_1082);
or U591 (N_591,N_312,In_1491);
xnor U592 (N_592,In_24,N_311);
nor U593 (N_593,In_1332,In_527);
and U594 (N_594,In_679,N_82);
and U595 (N_595,N_263,N_426);
nand U596 (N_596,In_894,In_1429);
or U597 (N_597,In_314,In_753);
and U598 (N_598,N_153,N_115);
nand U599 (N_599,N_155,In_150);
and U600 (N_600,N_590,In_590);
xnor U601 (N_601,In_1231,In_957);
or U602 (N_602,In_71,In_983);
or U603 (N_603,In_1164,In_652);
nor U604 (N_604,N_519,In_1382);
nor U605 (N_605,In_350,In_200);
xor U606 (N_606,N_162,N_291);
or U607 (N_607,In_491,In_763);
and U608 (N_608,In_436,N_578);
nor U609 (N_609,N_66,N_240);
nand U610 (N_610,In_1431,N_436);
nand U611 (N_611,In_411,N_402);
nand U612 (N_612,In_1368,N_377);
xnor U613 (N_613,In_654,N_557);
or U614 (N_614,N_448,N_39);
or U615 (N_615,N_498,In_198);
and U616 (N_616,In_754,N_338);
nand U617 (N_617,In_1176,In_1406);
nand U618 (N_618,In_656,N_480);
xnor U619 (N_619,In_126,N_416);
xnor U620 (N_620,N_177,In_787);
and U621 (N_621,N_535,N_467);
nand U622 (N_622,N_559,N_410);
and U623 (N_623,In_423,In_1072);
nand U624 (N_624,In_732,N_574);
or U625 (N_625,N_470,N_228);
and U626 (N_626,In_1006,In_583);
or U627 (N_627,N_391,N_340);
nor U628 (N_628,N_238,In_165);
xor U629 (N_629,In_584,In_384);
nand U630 (N_630,N_417,In_234);
nand U631 (N_631,In_1181,N_194);
or U632 (N_632,N_207,N_552);
xnor U633 (N_633,In_768,In_273);
xor U634 (N_634,N_453,N_560);
nand U635 (N_635,N_540,N_331);
and U636 (N_636,N_374,In_416);
nor U637 (N_637,In_1237,In_961);
nand U638 (N_638,N_239,In_1461);
nand U639 (N_639,In_123,In_886);
nor U640 (N_640,In_935,N_539);
nand U641 (N_641,In_958,N_468);
or U642 (N_642,N_317,In_820);
nand U643 (N_643,N_59,N_523);
or U644 (N_644,In_1499,N_257);
or U645 (N_645,N_212,In_1307);
nor U646 (N_646,In_546,N_270);
nand U647 (N_647,In_426,In_1440);
nand U648 (N_648,N_586,N_517);
xor U649 (N_649,In_1042,In_391);
or U650 (N_650,N_131,In_1362);
or U651 (N_651,In_574,In_15);
nand U652 (N_652,N_318,N_407);
and U653 (N_653,N_386,In_136);
and U654 (N_654,N_520,In_1250);
nand U655 (N_655,N_544,In_1094);
and U656 (N_656,In_627,N_504);
or U657 (N_657,In_1021,In_1039);
xor U658 (N_658,In_222,In_1341);
nor U659 (N_659,In_1016,In_189);
xor U660 (N_660,In_11,In_1044);
nor U661 (N_661,N_224,In_687);
xnor U662 (N_662,In_736,In_395);
nand U663 (N_663,In_710,In_1489);
and U664 (N_664,In_142,In_1497);
xnor U665 (N_665,N_105,N_530);
or U666 (N_666,In_346,N_5);
xnor U667 (N_667,In_1374,In_38);
nor U668 (N_668,N_512,In_312);
or U669 (N_669,In_443,In_907);
nor U670 (N_670,In_63,In_1155);
and U671 (N_671,N_521,In_307);
and U672 (N_672,In_267,N_454);
nor U673 (N_673,N_526,N_587);
nand U674 (N_674,In_761,N_451);
xnor U675 (N_675,In_369,In_1067);
or U676 (N_676,In_927,In_1466);
and U677 (N_677,N_395,N_356);
nand U678 (N_678,N_541,N_289);
or U679 (N_679,In_52,N_168);
nand U680 (N_680,In_658,In_14);
xnor U681 (N_681,In_188,N_599);
and U682 (N_682,In_6,In_482);
and U683 (N_683,N_551,In_1057);
and U684 (N_684,N_70,In_440);
nand U685 (N_685,In_373,N_585);
and U686 (N_686,N_409,In_579);
xor U687 (N_687,N_508,In_296);
and U688 (N_688,In_1211,In_716);
nor U689 (N_689,In_249,In_1278);
or U690 (N_690,N_547,In_1093);
and U691 (N_691,In_432,In_874);
or U692 (N_692,In_521,In_783);
nand U693 (N_693,N_461,In_807);
and U694 (N_694,N_565,N_366);
and U695 (N_695,In_1477,N_94);
or U696 (N_696,In_388,N_307);
nand U697 (N_697,In_762,N_210);
nand U698 (N_698,In_993,In_603);
or U699 (N_699,In_0,In_815);
xor U700 (N_700,N_332,N_354);
nand U701 (N_701,In_1035,N_466);
and U702 (N_702,In_429,N_505);
nand U703 (N_703,In_530,N_568);
or U704 (N_704,N_195,N_492);
xor U705 (N_705,In_1216,N_305);
nor U706 (N_706,N_516,In_1463);
nand U707 (N_707,In_739,In_1005);
nand U708 (N_708,N_534,N_4);
nor U709 (N_709,In_641,N_174);
or U710 (N_710,N_573,In_43);
nand U711 (N_711,In_1496,N_244);
or U712 (N_712,In_1028,In_611);
or U713 (N_713,N_408,N_320);
nand U714 (N_714,In_1234,N_192);
or U715 (N_715,In_1416,In_1062);
nor U716 (N_716,In_1129,N_300);
or U717 (N_717,N_528,N_533);
or U718 (N_718,In_347,N_27);
and U719 (N_719,N_84,In_105);
nor U720 (N_720,In_1223,N_462);
nand U721 (N_721,In_949,N_11);
and U722 (N_722,In_878,N_398);
and U723 (N_723,In_376,N_548);
nor U724 (N_724,N_582,N_367);
nor U725 (N_725,N_216,N_596);
and U726 (N_726,In_1297,In_1114);
and U727 (N_727,N_522,In_246);
and U728 (N_728,N_8,N_221);
xor U729 (N_729,N_483,In_1242);
nand U730 (N_730,N_246,N_348);
nand U731 (N_731,In_991,In_460);
nand U732 (N_732,N_104,N_252);
and U733 (N_733,In_1334,In_1205);
nor U734 (N_734,In_141,N_16);
or U735 (N_735,In_956,N_172);
xnor U736 (N_736,In_471,In_75);
nand U737 (N_737,In_64,N_371);
nand U738 (N_738,In_223,N_581);
nor U739 (N_739,N_138,In_128);
nand U740 (N_740,In_986,In_545);
xor U741 (N_741,In_1475,In_972);
or U742 (N_742,N_309,In_454);
nor U743 (N_743,In_495,In_213);
nand U744 (N_744,In_1024,In_415);
or U745 (N_745,N_100,N_37);
nand U746 (N_746,N_545,N_591);
or U747 (N_747,N_563,N_510);
and U748 (N_748,In_1397,N_186);
or U749 (N_749,N_199,N_431);
nor U750 (N_750,In_434,In_898);
or U751 (N_751,In_675,N_434);
or U752 (N_752,N_629,In_266);
nand U753 (N_753,N_364,N_433);
nand U754 (N_754,N_352,In_971);
or U755 (N_755,In_1253,N_399);
and U756 (N_756,In_726,In_289);
and U757 (N_757,In_902,N_739);
nand U758 (N_758,In_414,N_494);
xnor U759 (N_759,N_182,In_863);
nor U760 (N_760,In_44,N_609);
nand U761 (N_761,N_393,N_692);
xor U762 (N_762,N_554,In_1287);
and U763 (N_763,N_485,In_134);
and U764 (N_764,N_749,N_330);
nor U765 (N_765,N_717,In_940);
nand U766 (N_766,N_641,In_1484);
nand U767 (N_767,N_476,N_343);
xor U768 (N_768,In_632,In_155);
xor U769 (N_769,N_584,N_718);
nand U770 (N_770,In_515,N_640);
nand U771 (N_771,N_154,In_912);
and U772 (N_772,N_473,N_351);
xor U773 (N_773,N_737,N_496);
xor U774 (N_774,In_239,N_95);
nor U775 (N_775,N_677,In_1003);
nor U776 (N_776,N_13,N_697);
or U777 (N_777,N_598,In_103);
and U778 (N_778,N_583,N_633);
xnor U779 (N_779,N_594,N_708);
or U780 (N_780,N_418,In_550);
and U781 (N_781,In_921,N_293);
nand U782 (N_782,N_690,In_229);
or U783 (N_783,In_241,N_682);
nand U784 (N_784,In_1446,N_686);
and U785 (N_785,In_1190,In_459);
xor U786 (N_786,N_669,N_18);
or U787 (N_787,N_612,In_1288);
and U788 (N_788,N_64,N_344);
xnor U789 (N_789,N_443,In_604);
nor U790 (N_790,N_495,N_710);
and U791 (N_791,In_1372,In_1451);
nor U792 (N_792,N_264,N_663);
and U793 (N_793,N_85,In_943);
or U794 (N_794,N_642,In_917);
xor U795 (N_795,In_74,In_615);
xnor U796 (N_796,In_529,N_730);
xor U797 (N_797,In_1083,N_604);
nand U798 (N_798,N_693,In_667);
or U799 (N_799,In_40,N_423);
nor U800 (N_800,In_1286,N_597);
nor U801 (N_801,N_619,N_617);
and U802 (N_802,In_469,In_220);
or U803 (N_803,In_551,N_650);
and U804 (N_804,N_388,N_722);
xnor U805 (N_805,In_853,N_747);
xor U806 (N_806,N_23,In_1414);
and U807 (N_807,In_1492,N_225);
xor U808 (N_808,N_326,In_759);
xor U809 (N_809,N_611,In_124);
or U810 (N_810,In_139,N_580);
nand U811 (N_811,In_1352,N_275);
xor U812 (N_812,In_1065,In_749);
and U813 (N_813,N_572,In_642);
and U814 (N_814,N_694,N_258);
xnor U815 (N_815,In_1130,N_622);
xor U816 (N_816,In_1313,In_265);
and U817 (N_817,N_157,N_575);
or U818 (N_818,N_733,N_729);
nor U819 (N_819,In_1264,N_425);
xnor U820 (N_820,N_743,In_714);
xor U821 (N_821,N_427,N_696);
nor U822 (N_822,N_744,N_748);
nor U823 (N_823,N_363,N_636);
xor U824 (N_824,N_119,In_493);
and U825 (N_825,N_732,N_606);
and U826 (N_826,In_1479,N_380);
or U827 (N_827,N_707,N_126);
or U828 (N_828,N_484,In_1008);
nand U829 (N_829,N_564,N_706);
or U830 (N_830,In_113,N_324);
and U831 (N_831,In_91,N_558);
or U832 (N_832,In_534,In_372);
or U833 (N_833,In_438,N_370);
xor U834 (N_834,In_121,In_723);
or U835 (N_835,N_284,In_997);
xor U836 (N_836,N_490,N_721);
and U837 (N_837,N_713,N_621);
nor U838 (N_838,In_396,N_515);
and U839 (N_839,In_382,In_400);
or U840 (N_840,In_514,N_171);
nand U841 (N_841,N_607,In_299);
nand U842 (N_842,N_639,In_816);
and U843 (N_843,N_684,In_683);
or U844 (N_844,In_378,N_652);
and U845 (N_845,N_577,N_79);
or U846 (N_846,N_411,N_537);
xnor U847 (N_847,In_327,In_29);
or U848 (N_848,In_1004,In_364);
or U849 (N_849,N_394,In_70);
or U850 (N_850,In_635,In_1472);
xor U851 (N_851,N_628,In_173);
xnor U852 (N_852,N_680,N_553);
nor U853 (N_853,In_539,N_649);
xor U854 (N_854,N_653,In_1450);
and U855 (N_855,In_1370,In_470);
nor U856 (N_856,In_671,N_236);
and U857 (N_857,N_727,N_99);
xor U858 (N_858,N_488,N_49);
nand U859 (N_859,In_623,N_593);
nand U860 (N_860,In_771,N_698);
or U861 (N_861,N_672,N_465);
or U862 (N_862,In_786,N_310);
nor U863 (N_863,In_1165,N_282);
nand U864 (N_864,N_614,In_662);
and U865 (N_865,In_399,In_464);
nand U866 (N_866,In_817,N_382);
xnor U867 (N_867,N_705,N_673);
and U868 (N_868,N_691,N_643);
nand U869 (N_869,N_404,N_746);
nand U870 (N_870,In_985,In_948);
and U871 (N_871,In_410,N_603);
nand U872 (N_872,In_37,In_930);
nand U873 (N_873,In_670,N_440);
nor U874 (N_874,In_1483,In_677);
xnor U875 (N_875,N_477,N_679);
and U876 (N_876,In_909,N_538);
nand U877 (N_877,In_228,N_724);
nor U878 (N_878,In_449,In_1077);
and U879 (N_879,N_124,N_532);
nand U880 (N_880,In_1280,N_160);
and U881 (N_881,N_742,In_543);
nand U882 (N_882,N_301,N_514);
nand U883 (N_883,In_1225,N_183);
xnor U884 (N_884,N_579,In_232);
and U885 (N_885,In_1228,In_133);
nand U886 (N_886,N_500,N_497);
or U887 (N_887,N_474,N_478);
xnor U888 (N_888,N_562,N_735);
nand U889 (N_889,N_48,In_67);
nand U890 (N_890,N_610,In_186);
nand U891 (N_891,In_1248,In_672);
nand U892 (N_892,N_469,N_702);
nor U893 (N_893,N_373,In_1186);
xor U894 (N_894,In_375,In_586);
xnor U895 (N_895,N_543,In_1122);
nand U896 (N_896,N_73,In_1246);
or U897 (N_897,N_455,N_281);
xor U898 (N_898,N_513,In_348);
or U899 (N_899,N_725,N_357);
xor U900 (N_900,In_1144,In_76);
and U901 (N_901,In_1116,N_688);
xor U902 (N_902,N_658,N_714);
or U903 (N_903,In_887,In_899);
nand U904 (N_904,N_665,N_350);
xnor U905 (N_905,N_740,In_332);
nor U906 (N_906,In_362,N_745);
nor U907 (N_907,N_798,In_1100);
or U908 (N_908,N_438,N_771);
and U909 (N_909,N_620,N_862);
xnor U910 (N_910,N_659,N_786);
nand U911 (N_911,N_627,In_628);
and U912 (N_912,In_1050,N_840);
and U913 (N_913,N_353,N_894);
xnor U914 (N_914,N_660,In_730);
and U915 (N_915,N_40,N_836);
and U916 (N_916,N_832,In_224);
and U917 (N_917,N_306,In_439);
or U918 (N_918,N_794,N_303);
xnor U919 (N_919,N_175,N_882);
xnor U920 (N_920,N_396,N_602);
and U921 (N_921,In_561,N_229);
or U922 (N_922,In_172,N_623);
and U923 (N_923,In_1454,N_608);
or U924 (N_924,In_1270,N_757);
xor U925 (N_925,In_1312,In_889);
xor U926 (N_926,N_895,N_678);
or U927 (N_927,N_518,N_432);
nor U928 (N_928,In_1183,N_779);
nand U929 (N_929,In_1428,N_447);
xor U930 (N_930,N_812,N_750);
or U931 (N_931,In_317,N_780);
nor U932 (N_932,N_487,N_761);
xnor U933 (N_933,In_950,N_630);
nor U934 (N_934,In_1037,In_498);
and U935 (N_935,N_379,N_502);
or U936 (N_936,In_309,N_709);
and U937 (N_937,In_162,N_889);
and U938 (N_938,N_834,In_528);
xnor U939 (N_939,N_664,In_374);
and U940 (N_940,N_503,In_797);
nor U941 (N_941,N_86,N_765);
and U942 (N_942,N_796,N_635);
nand U943 (N_943,In_1113,In_1404);
nor U944 (N_944,In_1340,N_260);
xor U945 (N_945,In_532,N_661);
and U946 (N_946,N_493,In_361);
nor U947 (N_947,In_660,N_435);
xor U948 (N_948,N_863,N_58);
nand U949 (N_949,In_284,In_833);
or U950 (N_950,N_561,In_1458);
and U951 (N_951,In_218,In_706);
and U952 (N_952,N_613,In_285);
and U953 (N_953,N_445,N_511);
or U954 (N_954,N_249,In_967);
nor U955 (N_955,In_720,In_112);
nor U956 (N_956,In_23,N_827);
xor U957 (N_957,N_813,In_1309);
xnor U958 (N_958,N_362,In_140);
nand U959 (N_959,N_588,In_634);
nand U960 (N_960,N_489,In_1066);
nand U961 (N_961,N_879,In_617);
and U962 (N_962,N_589,In_728);
xor U963 (N_963,In_1367,N_638);
xnor U964 (N_964,N_806,N_760);
and U965 (N_965,N_442,N_98);
xnor U966 (N_966,In_934,N_428);
nor U967 (N_967,N_566,In_1070);
nand U968 (N_968,N_250,N_790);
xnor U969 (N_969,In_1292,In_1192);
and U970 (N_970,N_657,N_769);
or U971 (N_971,N_491,In_42);
or U972 (N_972,N_823,N_349);
xor U973 (N_973,N_31,N_685);
and U974 (N_974,N_758,N_546);
nor U975 (N_975,N_567,In_1289);
or U976 (N_976,N_464,N_390);
and U977 (N_977,In_196,N_262);
nor U978 (N_978,N_843,In_1301);
nand U979 (N_979,N_655,N_152);
nor U980 (N_980,N_716,N_818);
nor U981 (N_981,N_47,N_662);
or U982 (N_982,N_825,N_132);
nor U983 (N_983,In_48,N_644);
and U984 (N_984,N_872,N_778);
and U985 (N_985,In_523,N_865);
xor U986 (N_986,N_237,N_811);
and U987 (N_987,In_1073,In_588);
xor U988 (N_988,In_864,N_615);
xnor U989 (N_989,N_810,In_1229);
xnor U990 (N_990,N_855,In_758);
nor U991 (N_991,N_555,N_369);
and U992 (N_992,N_549,N_793);
and U993 (N_993,N_861,In_18);
nor U994 (N_994,In_1300,N_405);
nor U995 (N_995,N_42,In_938);
and U996 (N_996,In_1422,N_689);
xor U997 (N_997,In_1199,N_756);
xnor U998 (N_998,N_720,In_1335);
or U999 (N_999,N_828,N_387);
nor U1000 (N_1000,N_890,N_873);
and U1001 (N_1001,In_540,N_457);
nor U1002 (N_1002,N_667,In_653);
nor U1003 (N_1003,N_460,N_808);
and U1004 (N_1004,N_835,N_148);
nor U1005 (N_1005,In_713,In_825);
nand U1006 (N_1006,N_674,N_72);
nor U1007 (N_1007,N_576,N_327);
nor U1008 (N_1008,N_279,In_335);
and U1009 (N_1009,In_767,In_750);
and U1010 (N_1010,In_283,In_131);
nand U1011 (N_1011,N_108,N_265);
xor U1012 (N_1012,N_703,N_654);
nor U1013 (N_1013,In_562,In_661);
nand U1014 (N_1014,N_864,In_578);
or U1015 (N_1015,N_255,In_680);
nand U1016 (N_1016,N_571,In_278);
nand U1017 (N_1017,In_1157,In_501);
and U1018 (N_1018,N_20,N_251);
nand U1019 (N_1019,In_452,In_1453);
nor U1020 (N_1020,N_885,N_838);
nand U1021 (N_1021,N_845,N_92);
or U1022 (N_1022,In_705,In_1172);
xor U1023 (N_1023,N_734,In_41);
nor U1024 (N_1024,N_536,In_149);
nand U1025 (N_1025,N_870,N_68);
xor U1026 (N_1026,In_50,N_529);
and U1027 (N_1027,N_345,N_711);
nor U1028 (N_1028,In_614,N_795);
xnor U1029 (N_1029,N_525,N_441);
nor U1030 (N_1030,N_883,N_736);
nor U1031 (N_1031,In_106,In_659);
nor U1032 (N_1032,N_325,N_871);
or U1033 (N_1033,N_401,N_645);
nor U1034 (N_1034,In_973,N_361);
nand U1035 (N_1035,N_595,In_512);
or U1036 (N_1036,In_1197,In_692);
or U1037 (N_1037,N_459,In_277);
xor U1038 (N_1038,In_1171,In_869);
nand U1039 (N_1039,In_571,N_852);
nand U1040 (N_1040,In_1347,N_288);
and U1041 (N_1041,N_802,N_723);
and U1042 (N_1042,In_1201,N_381);
xor U1043 (N_1043,N_848,In_1358);
nor U1044 (N_1044,In_333,In_209);
or U1045 (N_1045,N_826,N_831);
nand U1046 (N_1046,In_568,In_883);
nand U1047 (N_1047,N_675,N_150);
nand U1048 (N_1048,N_876,N_524);
nand U1049 (N_1049,N_821,N_359);
and U1050 (N_1050,N_1033,In_418);
nor U1051 (N_1051,N_921,N_947);
and U1052 (N_1052,N_286,N_1025);
xnor U1053 (N_1053,N_570,N_905);
or U1054 (N_1054,In_595,N_915);
xor U1055 (N_1055,N_191,N_1044);
xnor U1056 (N_1056,N_880,N_797);
nor U1057 (N_1057,N_481,N_991);
or U1058 (N_1058,N_822,N_1018);
nor U1059 (N_1059,N_1032,In_1064);
nand U1060 (N_1060,N_856,N_983);
xor U1061 (N_1061,In_513,N_217);
nand U1062 (N_1062,N_328,N_302);
nor U1063 (N_1063,N_437,N_1045);
and U1064 (N_1064,N_283,N_978);
or U1065 (N_1065,N_902,N_241);
xnor U1066 (N_1066,N_471,In_331);
nor U1067 (N_1067,N_378,N_368);
and U1068 (N_1068,N_807,N_984);
nand U1069 (N_1069,N_763,In_1235);
xor U1070 (N_1070,N_314,In_1214);
or U1071 (N_1071,N_77,N_695);
nand U1072 (N_1072,In_760,N_741);
nand U1073 (N_1073,N_935,N_931);
xnor U1074 (N_1074,N_701,N_118);
and U1075 (N_1075,N_458,N_958);
nand U1076 (N_1076,N_190,N_135);
or U1077 (N_1077,In_827,N_904);
or U1078 (N_1078,N_914,In_891);
nand U1079 (N_1079,N_916,In_1476);
and U1080 (N_1080,N_605,N_860);
nand U1081 (N_1081,N_859,In_994);
and U1082 (N_1082,N_809,In_790);
and U1083 (N_1083,N_297,In_1423);
or U1084 (N_1084,N_945,N_556);
or U1085 (N_1085,N_875,N_987);
and U1086 (N_1086,N_626,N_1029);
and U1087 (N_1087,N_815,N_1034);
or U1088 (N_1088,N_550,In_146);
or U1089 (N_1089,N_752,N_846);
and U1090 (N_1090,N_1009,N_908);
nor U1091 (N_1091,N_817,N_1010);
nor U1092 (N_1092,In_248,N_853);
xor U1093 (N_1093,N_966,N_1006);
nand U1094 (N_1094,N_209,In_702);
xnor U1095 (N_1095,N_782,In_492);
nand U1096 (N_1096,N_683,N_924);
nand U1097 (N_1097,N_647,In_644);
or U1098 (N_1098,N_930,N_601);
and U1099 (N_1099,In_770,In_216);
nand U1100 (N_1100,N_456,N_800);
nand U1101 (N_1101,N_775,N_1021);
xnor U1102 (N_1102,N_920,In_484);
and U1103 (N_1103,N_937,N_444);
or U1104 (N_1104,N_781,N_851);
xnor U1105 (N_1105,N_759,N_927);
nand U1106 (N_1106,In_813,In_170);
and U1107 (N_1107,N_430,N_712);
nor U1108 (N_1108,N_936,N_479);
and U1109 (N_1109,N_231,N_1022);
or U1110 (N_1110,N_884,In_919);
nor U1111 (N_1111,N_994,N_944);
or U1112 (N_1112,N_878,N_501);
xnor U1113 (N_1113,N_452,N_499);
or U1114 (N_1114,N_1016,N_670);
xor U1115 (N_1115,In_231,N_976);
or U1116 (N_1116,N_429,N_1031);
and U1117 (N_1117,N_668,N_268);
and U1118 (N_1118,N_1049,N_857);
and U1119 (N_1119,N_422,N_943);
and U1120 (N_1120,In_1145,In_1153);
or U1121 (N_1121,N_341,In_549);
nand U1122 (N_1122,N_844,In_1036);
nand U1123 (N_1123,N_624,In_465);
xnor U1124 (N_1124,N_990,N_506);
nor U1125 (N_1125,N_819,N_634);
xnor U1126 (N_1126,N_687,N_768);
or U1127 (N_1127,In_507,N_919);
or U1128 (N_1128,N_932,In_626);
and U1129 (N_1129,N_993,In_1468);
nor U1130 (N_1130,N_569,N_933);
xnor U1131 (N_1131,N_107,In_573);
or U1132 (N_1132,N_25,In_1373);
xor U1133 (N_1133,N_1008,N_981);
xnor U1134 (N_1134,N_1042,N_866);
or U1135 (N_1135,N_1007,In_1269);
nor U1136 (N_1136,N_918,N_888);
and U1137 (N_1137,N_482,N_867);
nand U1138 (N_1138,In_1283,N_774);
or U1139 (N_1139,N_839,N_646);
or U1140 (N_1140,N_973,N_751);
xnor U1141 (N_1141,N_934,N_928);
and U1142 (N_1142,N_791,In_629);
or U1143 (N_1143,N_531,N_785);
and U1144 (N_1144,N_893,N_463);
and U1145 (N_1145,N_592,N_1003);
and U1146 (N_1146,N_486,N_974);
or U1147 (N_1147,In_639,N_909);
xor U1148 (N_1148,In_1068,N_1046);
nor U1149 (N_1149,N_979,N_389);
or U1150 (N_1150,N_849,N_125);
xor U1151 (N_1151,N_776,N_167);
nor U1152 (N_1152,N_1024,N_1015);
and U1153 (N_1153,N_939,N_392);
and U1154 (N_1154,N_93,N_449);
and U1155 (N_1155,N_41,N_824);
or U1156 (N_1156,N_820,N_600);
nor U1157 (N_1157,In_1331,N_53);
xor U1158 (N_1158,N_969,N_777);
nor U1159 (N_1159,In_581,In_260);
and U1160 (N_1160,N_874,In_430);
or U1161 (N_1161,In_358,N_959);
and U1162 (N_1162,N_789,N_949);
nor U1163 (N_1163,N_656,In_572);
and U1164 (N_1164,N_948,In_61);
nand U1165 (N_1165,N_803,N_280);
and U1166 (N_1166,In_1266,N_323);
or U1167 (N_1167,N_922,N_625);
nor U1168 (N_1168,N_637,N_450);
nand U1169 (N_1169,N_648,N_975);
nor U1170 (N_1170,N_719,In_488);
xor U1171 (N_1171,N_54,N_814);
xnor U1172 (N_1172,N_891,N_829);
xnor U1173 (N_1173,N_972,N_414);
xnor U1174 (N_1174,N_868,N_962);
nand U1175 (N_1175,N_805,N_897);
nor U1176 (N_1176,N_715,In_1244);
nand U1177 (N_1177,N_830,N_941);
and U1178 (N_1178,N_833,N_923);
nand U1179 (N_1179,N_854,N_988);
xor U1180 (N_1180,N_784,N_1036);
nor U1181 (N_1181,N_954,N_938);
nand U1182 (N_1182,N_1020,In_270);
nand U1183 (N_1183,N_1027,N_762);
nor U1184 (N_1184,N_989,N_1028);
nand U1185 (N_1185,In_1478,N_1040);
or U1186 (N_1186,N_365,In_235);
nand U1187 (N_1187,N_1043,N_1002);
nor U1188 (N_1188,N_1048,N_783);
nor U1189 (N_1189,N_965,N_952);
or U1190 (N_1190,N_898,In_801);
xnor U1191 (N_1191,N_1041,In_159);
xnor U1192 (N_1192,N_869,In_1311);
nand U1193 (N_1193,N_900,N_1030);
nor U1194 (N_1194,N_906,N_339);
nand U1195 (N_1195,N_901,N_1017);
nor U1196 (N_1196,N_1047,N_196);
nor U1197 (N_1197,N_946,N_728);
xnor U1198 (N_1198,In_1420,N_929);
xnor U1199 (N_1199,N_960,N_542);
xnor U1200 (N_1200,N_1093,N_847);
or U1201 (N_1201,N_992,N_1106);
nor U1202 (N_1202,N_1124,N_424);
nor U1203 (N_1203,N_631,In_668);
nand U1204 (N_1204,N_1037,N_1173);
and U1205 (N_1205,N_1073,N_1180);
and U1206 (N_1206,N_507,N_913);
xnor U1207 (N_1207,N_1059,N_788);
nor U1208 (N_1208,N_1068,N_681);
and U1209 (N_1209,N_877,N_397);
or U1210 (N_1210,N_1112,N_1050);
and U1211 (N_1211,N_704,N_1157);
nand U1212 (N_1212,N_1174,N_1129);
and U1213 (N_1213,N_982,N_1188);
or U1214 (N_1214,In_1336,N_1075);
nor U1215 (N_1215,N_1084,N_1161);
or U1216 (N_1216,In_337,N_700);
and U1217 (N_1217,N_472,N_1062);
nand U1218 (N_1218,N_1052,N_1145);
or U1219 (N_1219,N_1107,N_1148);
nor U1220 (N_1220,N_1194,In_773);
nor U1221 (N_1221,N_1051,N_1079);
nand U1222 (N_1222,N_1067,N_38);
nand U1223 (N_1223,N_1066,In_576);
xor U1224 (N_1224,N_997,N_1110);
or U1225 (N_1225,N_1136,N_1119);
nor U1226 (N_1226,N_1000,N_1104);
xnor U1227 (N_1227,N_1143,N_1065);
xnor U1228 (N_1228,N_986,N_899);
xnor U1229 (N_1229,N_1118,N_1153);
nand U1230 (N_1230,In_1059,N_187);
and U1231 (N_1231,N_963,N_1035);
and U1232 (N_1232,N_887,N_772);
xnor U1233 (N_1233,N_1091,N_837);
or U1234 (N_1234,N_754,N_315);
xor U1235 (N_1235,N_1102,N_787);
nor U1236 (N_1236,N_995,N_509);
nor U1237 (N_1237,N_1144,N_1094);
or U1238 (N_1238,N_1012,N_903);
and U1239 (N_1239,N_383,N_738);
nor U1240 (N_1240,N_1039,N_767);
nand U1241 (N_1241,N_1001,In_195);
nand U1242 (N_1242,N_1125,N_726);
and U1243 (N_1243,N_1183,N_967);
nor U1244 (N_1244,N_1165,In_1041);
nand U1245 (N_1245,N_1154,N_1120);
xor U1246 (N_1246,N_1014,In_793);
nor U1247 (N_1247,N_1115,N_1038);
nor U1248 (N_1248,N_886,N_1164);
nor U1249 (N_1249,N_1069,N_1086);
nand U1250 (N_1250,In_600,N_799);
xnor U1251 (N_1251,N_753,N_1082);
xor U1252 (N_1252,N_1166,N_770);
xnor U1253 (N_1253,N_1127,N_1197);
or U1254 (N_1254,N_881,N_1181);
nor U1255 (N_1255,N_801,N_1186);
nor U1256 (N_1256,N_1099,N_1070);
or U1257 (N_1257,N_764,N_1177);
nand U1258 (N_1258,N_475,N_1134);
nor U1259 (N_1259,N_1121,In_1014);
or U1260 (N_1260,N_977,N_1023);
nor U1261 (N_1261,N_1097,N_1123);
nor U1262 (N_1262,N_942,N_766);
and U1263 (N_1263,N_1061,N_792);
nand U1264 (N_1264,N_527,N_188);
nor U1265 (N_1265,N_1087,N_968);
and U1266 (N_1266,N_951,N_1063);
xnor U1267 (N_1267,N_911,N_1011);
or U1268 (N_1268,In_876,N_1117);
nor U1269 (N_1269,N_1088,N_1101);
nand U1270 (N_1270,In_1189,In_356);
nand U1271 (N_1271,N_1013,N_1163);
nand U1272 (N_1272,N_1081,N_1193);
and U1273 (N_1273,N_1055,N_917);
xor U1274 (N_1274,N_676,N_1175);
or U1275 (N_1275,N_1169,N_950);
or U1276 (N_1276,N_1159,N_299);
nand U1277 (N_1277,N_1058,N_1167);
and U1278 (N_1278,N_1085,N_1151);
and U1279 (N_1279,N_671,N_1139);
or U1280 (N_1280,N_1146,In_966);
and U1281 (N_1281,N_1155,N_1074);
and U1282 (N_1282,N_1098,N_892);
nand U1283 (N_1283,N_996,N_1056);
nor U1284 (N_1284,N_376,N_912);
nor U1285 (N_1285,N_955,In_1148);
xor U1286 (N_1286,N_971,N_842);
nor U1287 (N_1287,In_205,N_970);
xor U1288 (N_1288,N_1064,N_616);
xnor U1289 (N_1289,N_1077,N_1150);
xnor U1290 (N_1290,N_773,N_1092);
xor U1291 (N_1291,N_1116,N_1130);
xnor U1292 (N_1292,N_956,In_1134);
xnor U1293 (N_1293,N_632,N_1191);
and U1294 (N_1294,In_1007,N_294);
or U1295 (N_1295,N_910,N_850);
and U1296 (N_1296,N_1078,N_1135);
and U1297 (N_1297,N_858,N_1160);
nand U1298 (N_1298,N_1168,N_1185);
nor U1299 (N_1299,N_1072,N_1071);
xor U1300 (N_1300,In_1395,N_1147);
and U1301 (N_1301,In_110,N_1184);
nand U1302 (N_1302,N_1111,N_272);
nand U1303 (N_1303,N_1187,N_953);
and U1304 (N_1304,In_977,N_1162);
nor U1305 (N_1305,N_666,In_1298);
nor U1306 (N_1306,N_1076,N_1057);
nor U1307 (N_1307,N_1133,N_1126);
xnor U1308 (N_1308,N_1189,N_1195);
nor U1309 (N_1309,N_1170,N_1114);
nor U1310 (N_1310,N_1026,N_940);
or U1311 (N_1311,N_926,N_985);
xor U1312 (N_1312,N_1096,N_1054);
or U1313 (N_1313,N_1108,N_841);
nand U1314 (N_1314,N_1109,N_149);
and U1315 (N_1315,In_505,N_1171);
nor U1316 (N_1316,N_1122,N_295);
nand U1317 (N_1317,N_804,N_755);
or U1318 (N_1318,N_1142,N_1019);
xor U1319 (N_1319,N_907,N_699);
or U1320 (N_1320,N_618,N_651);
or U1321 (N_1321,In_3,N_1089);
or U1322 (N_1322,N_1172,N_62);
or U1323 (N_1323,N_406,N_998);
or U1324 (N_1324,N_1105,N_1100);
nor U1325 (N_1325,N_1179,N_1192);
nand U1326 (N_1326,N_1196,In_413);
nand U1327 (N_1327,N_1158,N_1053);
nor U1328 (N_1328,N_1004,N_816);
xnor U1329 (N_1329,N_1080,N_1113);
xor U1330 (N_1330,N_980,N_1131);
or U1331 (N_1331,N_128,In_111);
nor U1332 (N_1332,N_1132,N_413);
nor U1333 (N_1333,In_1251,N_1156);
nor U1334 (N_1334,N_961,N_1060);
and U1335 (N_1335,N_1083,N_313);
nor U1336 (N_1336,N_957,N_1138);
or U1337 (N_1337,N_1095,N_999);
xor U1338 (N_1338,N_1128,N_319);
nand U1339 (N_1339,N_1178,N_1005);
nor U1340 (N_1340,N_1103,N_1182);
nand U1341 (N_1341,N_1198,In_1435);
or U1342 (N_1342,N_1090,N_1149);
nor U1343 (N_1343,N_1140,N_964);
or U1344 (N_1344,N_1137,In_336);
nand U1345 (N_1345,N_1176,N_1190);
nor U1346 (N_1346,N_925,N_731);
nor U1347 (N_1347,In_844,N_1152);
or U1348 (N_1348,In_367,N_1199);
nor U1349 (N_1349,N_896,N_1141);
nand U1350 (N_1350,N_1298,N_1263);
or U1351 (N_1351,N_1305,N_1320);
nor U1352 (N_1352,N_1233,N_1343);
and U1353 (N_1353,N_1223,N_1220);
xnor U1354 (N_1354,N_1202,N_1207);
and U1355 (N_1355,N_1331,N_1313);
nor U1356 (N_1356,N_1262,N_1279);
xnor U1357 (N_1357,N_1315,N_1201);
nor U1358 (N_1358,N_1288,N_1328);
nor U1359 (N_1359,N_1286,N_1219);
nor U1360 (N_1360,N_1349,N_1230);
xnor U1361 (N_1361,N_1212,N_1200);
or U1362 (N_1362,N_1252,N_1248);
nand U1363 (N_1363,N_1275,N_1299);
nand U1364 (N_1364,N_1260,N_1303);
xor U1365 (N_1365,N_1242,N_1322);
nor U1366 (N_1366,N_1249,N_1341);
xor U1367 (N_1367,N_1325,N_1342);
and U1368 (N_1368,N_1278,N_1243);
or U1369 (N_1369,N_1256,N_1307);
and U1370 (N_1370,N_1302,N_1234);
and U1371 (N_1371,N_1336,N_1269);
xnor U1372 (N_1372,N_1290,N_1225);
and U1373 (N_1373,N_1270,N_1346);
and U1374 (N_1374,N_1257,N_1216);
nand U1375 (N_1375,N_1265,N_1314);
xor U1376 (N_1376,N_1235,N_1224);
nor U1377 (N_1377,N_1259,N_1347);
nor U1378 (N_1378,N_1335,N_1251);
and U1379 (N_1379,N_1308,N_1318);
or U1380 (N_1380,N_1291,N_1229);
or U1381 (N_1381,N_1236,N_1258);
nand U1382 (N_1382,N_1276,N_1239);
and U1383 (N_1383,N_1285,N_1254);
nor U1384 (N_1384,N_1326,N_1211);
and U1385 (N_1385,N_1245,N_1330);
or U1386 (N_1386,N_1213,N_1274);
or U1387 (N_1387,N_1319,N_1329);
or U1388 (N_1388,N_1283,N_1215);
xor U1389 (N_1389,N_1280,N_1228);
nor U1390 (N_1390,N_1272,N_1237);
xnor U1391 (N_1391,N_1301,N_1294);
nand U1392 (N_1392,N_1264,N_1324);
or U1393 (N_1393,N_1300,N_1316);
nor U1394 (N_1394,N_1287,N_1309);
or U1395 (N_1395,N_1222,N_1293);
nor U1396 (N_1396,N_1281,N_1297);
nand U1397 (N_1397,N_1232,N_1231);
nor U1398 (N_1398,N_1339,N_1282);
xnor U1399 (N_1399,N_1327,N_1277);
nand U1400 (N_1400,N_1334,N_1271);
or U1401 (N_1401,N_1206,N_1247);
or U1402 (N_1402,N_1311,N_1209);
and U1403 (N_1403,N_1338,N_1348);
xor U1404 (N_1404,N_1227,N_1296);
or U1405 (N_1405,N_1241,N_1246);
or U1406 (N_1406,N_1345,N_1317);
nand U1407 (N_1407,N_1238,N_1255);
and U1408 (N_1408,N_1273,N_1340);
nand U1409 (N_1409,N_1221,N_1321);
or U1410 (N_1410,N_1332,N_1261);
and U1411 (N_1411,N_1306,N_1266);
nor U1412 (N_1412,N_1333,N_1312);
xnor U1413 (N_1413,N_1289,N_1218);
and U1414 (N_1414,N_1292,N_1217);
nand U1415 (N_1415,N_1304,N_1310);
or U1416 (N_1416,N_1226,N_1244);
nand U1417 (N_1417,N_1337,N_1204);
xnor U1418 (N_1418,N_1253,N_1210);
nor U1419 (N_1419,N_1268,N_1295);
xnor U1420 (N_1420,N_1240,N_1214);
nor U1421 (N_1421,N_1284,N_1250);
nor U1422 (N_1422,N_1203,N_1208);
xor U1423 (N_1423,N_1205,N_1344);
xnor U1424 (N_1424,N_1323,N_1267);
xor U1425 (N_1425,N_1234,N_1279);
nand U1426 (N_1426,N_1311,N_1318);
nand U1427 (N_1427,N_1245,N_1344);
or U1428 (N_1428,N_1250,N_1225);
and U1429 (N_1429,N_1313,N_1250);
or U1430 (N_1430,N_1301,N_1314);
or U1431 (N_1431,N_1256,N_1292);
xor U1432 (N_1432,N_1241,N_1295);
xnor U1433 (N_1433,N_1226,N_1205);
xor U1434 (N_1434,N_1328,N_1244);
or U1435 (N_1435,N_1315,N_1263);
xnor U1436 (N_1436,N_1287,N_1288);
nor U1437 (N_1437,N_1203,N_1297);
nor U1438 (N_1438,N_1240,N_1254);
xor U1439 (N_1439,N_1263,N_1241);
or U1440 (N_1440,N_1244,N_1234);
nand U1441 (N_1441,N_1304,N_1243);
xor U1442 (N_1442,N_1211,N_1200);
and U1443 (N_1443,N_1299,N_1233);
and U1444 (N_1444,N_1342,N_1326);
nand U1445 (N_1445,N_1298,N_1282);
xor U1446 (N_1446,N_1227,N_1320);
or U1447 (N_1447,N_1278,N_1224);
xnor U1448 (N_1448,N_1259,N_1336);
nor U1449 (N_1449,N_1303,N_1217);
or U1450 (N_1450,N_1321,N_1320);
or U1451 (N_1451,N_1234,N_1206);
and U1452 (N_1452,N_1319,N_1334);
nor U1453 (N_1453,N_1264,N_1335);
or U1454 (N_1454,N_1235,N_1214);
and U1455 (N_1455,N_1267,N_1274);
nand U1456 (N_1456,N_1202,N_1301);
nor U1457 (N_1457,N_1252,N_1293);
nor U1458 (N_1458,N_1299,N_1229);
xnor U1459 (N_1459,N_1333,N_1269);
or U1460 (N_1460,N_1218,N_1283);
xnor U1461 (N_1461,N_1278,N_1202);
and U1462 (N_1462,N_1213,N_1321);
nor U1463 (N_1463,N_1336,N_1235);
nand U1464 (N_1464,N_1246,N_1273);
nor U1465 (N_1465,N_1260,N_1323);
or U1466 (N_1466,N_1268,N_1266);
xnor U1467 (N_1467,N_1249,N_1345);
nand U1468 (N_1468,N_1244,N_1233);
nor U1469 (N_1469,N_1231,N_1223);
nand U1470 (N_1470,N_1202,N_1243);
nor U1471 (N_1471,N_1227,N_1302);
xor U1472 (N_1472,N_1211,N_1216);
nor U1473 (N_1473,N_1315,N_1234);
nor U1474 (N_1474,N_1296,N_1201);
and U1475 (N_1475,N_1201,N_1241);
xor U1476 (N_1476,N_1294,N_1307);
and U1477 (N_1477,N_1297,N_1348);
xor U1478 (N_1478,N_1346,N_1304);
and U1479 (N_1479,N_1247,N_1224);
and U1480 (N_1480,N_1280,N_1284);
nand U1481 (N_1481,N_1282,N_1344);
xor U1482 (N_1482,N_1345,N_1324);
or U1483 (N_1483,N_1204,N_1259);
nor U1484 (N_1484,N_1205,N_1331);
and U1485 (N_1485,N_1250,N_1241);
nor U1486 (N_1486,N_1326,N_1278);
and U1487 (N_1487,N_1240,N_1244);
nand U1488 (N_1488,N_1255,N_1207);
or U1489 (N_1489,N_1276,N_1206);
or U1490 (N_1490,N_1304,N_1237);
or U1491 (N_1491,N_1312,N_1263);
or U1492 (N_1492,N_1308,N_1304);
nor U1493 (N_1493,N_1345,N_1297);
xor U1494 (N_1494,N_1259,N_1206);
and U1495 (N_1495,N_1262,N_1253);
nand U1496 (N_1496,N_1325,N_1295);
xnor U1497 (N_1497,N_1300,N_1269);
and U1498 (N_1498,N_1260,N_1265);
and U1499 (N_1499,N_1241,N_1303);
xnor U1500 (N_1500,N_1422,N_1421);
nor U1501 (N_1501,N_1419,N_1489);
and U1502 (N_1502,N_1462,N_1479);
and U1503 (N_1503,N_1366,N_1441);
xnor U1504 (N_1504,N_1395,N_1492);
nand U1505 (N_1505,N_1456,N_1491);
xnor U1506 (N_1506,N_1453,N_1386);
or U1507 (N_1507,N_1356,N_1372);
or U1508 (N_1508,N_1437,N_1448);
or U1509 (N_1509,N_1384,N_1425);
nor U1510 (N_1510,N_1402,N_1392);
and U1511 (N_1511,N_1475,N_1447);
nor U1512 (N_1512,N_1442,N_1451);
or U1513 (N_1513,N_1380,N_1400);
nor U1514 (N_1514,N_1397,N_1497);
xnor U1515 (N_1515,N_1381,N_1488);
or U1516 (N_1516,N_1438,N_1365);
xor U1517 (N_1517,N_1398,N_1495);
and U1518 (N_1518,N_1383,N_1410);
nand U1519 (N_1519,N_1490,N_1394);
and U1520 (N_1520,N_1379,N_1403);
and U1521 (N_1521,N_1393,N_1361);
and U1522 (N_1522,N_1471,N_1432);
nor U1523 (N_1523,N_1455,N_1469);
nand U1524 (N_1524,N_1466,N_1376);
nand U1525 (N_1525,N_1472,N_1358);
or U1526 (N_1526,N_1487,N_1388);
or U1527 (N_1527,N_1499,N_1485);
xnor U1528 (N_1528,N_1431,N_1414);
or U1529 (N_1529,N_1364,N_1477);
xnor U1530 (N_1530,N_1368,N_1423);
nor U1531 (N_1531,N_1353,N_1440);
nor U1532 (N_1532,N_1407,N_1468);
and U1533 (N_1533,N_1474,N_1369);
nand U1534 (N_1534,N_1424,N_1387);
nor U1535 (N_1535,N_1417,N_1415);
nand U1536 (N_1536,N_1494,N_1430);
nand U1537 (N_1537,N_1389,N_1406);
xor U1538 (N_1538,N_1426,N_1399);
xnor U1539 (N_1539,N_1473,N_1464);
and U1540 (N_1540,N_1416,N_1467);
or U1541 (N_1541,N_1390,N_1412);
nor U1542 (N_1542,N_1435,N_1405);
and U1543 (N_1543,N_1493,N_1449);
xnor U1544 (N_1544,N_1420,N_1480);
and U1545 (N_1545,N_1360,N_1378);
nor U1546 (N_1546,N_1498,N_1459);
nand U1547 (N_1547,N_1465,N_1357);
and U1548 (N_1548,N_1359,N_1434);
and U1549 (N_1549,N_1377,N_1496);
nor U1550 (N_1550,N_1486,N_1382);
and U1551 (N_1551,N_1482,N_1396);
or U1552 (N_1552,N_1443,N_1385);
nor U1553 (N_1553,N_1401,N_1460);
and U1554 (N_1554,N_1375,N_1408);
nor U1555 (N_1555,N_1484,N_1463);
and U1556 (N_1556,N_1436,N_1355);
nor U1557 (N_1557,N_1371,N_1370);
or U1558 (N_1558,N_1452,N_1391);
nand U1559 (N_1559,N_1374,N_1454);
and U1560 (N_1560,N_1418,N_1458);
and U1561 (N_1561,N_1354,N_1445);
and U1562 (N_1562,N_1457,N_1373);
nand U1563 (N_1563,N_1433,N_1362);
xor U1564 (N_1564,N_1461,N_1363);
or U1565 (N_1565,N_1483,N_1450);
nor U1566 (N_1566,N_1444,N_1351);
nor U1567 (N_1567,N_1350,N_1404);
and U1568 (N_1568,N_1367,N_1481);
or U1569 (N_1569,N_1409,N_1428);
or U1570 (N_1570,N_1413,N_1439);
and U1571 (N_1571,N_1446,N_1411);
or U1572 (N_1572,N_1478,N_1352);
nor U1573 (N_1573,N_1427,N_1429);
xor U1574 (N_1574,N_1470,N_1476);
xnor U1575 (N_1575,N_1416,N_1402);
xor U1576 (N_1576,N_1465,N_1361);
and U1577 (N_1577,N_1360,N_1462);
or U1578 (N_1578,N_1472,N_1414);
nand U1579 (N_1579,N_1440,N_1499);
nor U1580 (N_1580,N_1485,N_1452);
nor U1581 (N_1581,N_1430,N_1393);
xor U1582 (N_1582,N_1420,N_1379);
and U1583 (N_1583,N_1409,N_1459);
and U1584 (N_1584,N_1486,N_1350);
or U1585 (N_1585,N_1463,N_1443);
nor U1586 (N_1586,N_1368,N_1408);
nand U1587 (N_1587,N_1424,N_1480);
nor U1588 (N_1588,N_1439,N_1357);
nor U1589 (N_1589,N_1358,N_1471);
and U1590 (N_1590,N_1449,N_1434);
or U1591 (N_1591,N_1470,N_1412);
nand U1592 (N_1592,N_1353,N_1396);
nand U1593 (N_1593,N_1391,N_1457);
and U1594 (N_1594,N_1444,N_1428);
nand U1595 (N_1595,N_1456,N_1352);
nor U1596 (N_1596,N_1413,N_1355);
and U1597 (N_1597,N_1475,N_1381);
nor U1598 (N_1598,N_1400,N_1484);
nor U1599 (N_1599,N_1372,N_1473);
nand U1600 (N_1600,N_1448,N_1491);
or U1601 (N_1601,N_1379,N_1395);
nand U1602 (N_1602,N_1352,N_1421);
nor U1603 (N_1603,N_1494,N_1488);
xor U1604 (N_1604,N_1356,N_1393);
nand U1605 (N_1605,N_1477,N_1470);
xnor U1606 (N_1606,N_1498,N_1483);
and U1607 (N_1607,N_1459,N_1421);
nor U1608 (N_1608,N_1390,N_1427);
nand U1609 (N_1609,N_1373,N_1371);
xor U1610 (N_1610,N_1441,N_1472);
xnor U1611 (N_1611,N_1468,N_1405);
xnor U1612 (N_1612,N_1395,N_1445);
nor U1613 (N_1613,N_1496,N_1470);
or U1614 (N_1614,N_1463,N_1494);
xor U1615 (N_1615,N_1465,N_1368);
nor U1616 (N_1616,N_1397,N_1379);
xor U1617 (N_1617,N_1352,N_1446);
xor U1618 (N_1618,N_1369,N_1499);
nand U1619 (N_1619,N_1392,N_1451);
nor U1620 (N_1620,N_1463,N_1485);
and U1621 (N_1621,N_1381,N_1387);
xor U1622 (N_1622,N_1366,N_1431);
xor U1623 (N_1623,N_1368,N_1466);
or U1624 (N_1624,N_1393,N_1449);
nor U1625 (N_1625,N_1497,N_1384);
and U1626 (N_1626,N_1463,N_1351);
xor U1627 (N_1627,N_1456,N_1414);
and U1628 (N_1628,N_1414,N_1467);
and U1629 (N_1629,N_1393,N_1453);
nor U1630 (N_1630,N_1493,N_1351);
or U1631 (N_1631,N_1443,N_1389);
or U1632 (N_1632,N_1350,N_1499);
and U1633 (N_1633,N_1424,N_1385);
and U1634 (N_1634,N_1489,N_1466);
xor U1635 (N_1635,N_1430,N_1351);
or U1636 (N_1636,N_1451,N_1406);
and U1637 (N_1637,N_1445,N_1418);
xnor U1638 (N_1638,N_1450,N_1433);
xor U1639 (N_1639,N_1367,N_1399);
and U1640 (N_1640,N_1490,N_1373);
nand U1641 (N_1641,N_1479,N_1358);
nand U1642 (N_1642,N_1386,N_1364);
xnor U1643 (N_1643,N_1445,N_1373);
nor U1644 (N_1644,N_1397,N_1383);
and U1645 (N_1645,N_1434,N_1404);
nand U1646 (N_1646,N_1361,N_1480);
nor U1647 (N_1647,N_1482,N_1494);
or U1648 (N_1648,N_1438,N_1485);
xnor U1649 (N_1649,N_1362,N_1353);
nor U1650 (N_1650,N_1636,N_1647);
or U1651 (N_1651,N_1617,N_1563);
xor U1652 (N_1652,N_1638,N_1550);
nand U1653 (N_1653,N_1528,N_1512);
or U1654 (N_1654,N_1562,N_1613);
and U1655 (N_1655,N_1628,N_1625);
nand U1656 (N_1656,N_1637,N_1545);
nand U1657 (N_1657,N_1631,N_1557);
xnor U1658 (N_1658,N_1606,N_1630);
nand U1659 (N_1659,N_1588,N_1640);
nor U1660 (N_1660,N_1577,N_1569);
nor U1661 (N_1661,N_1547,N_1590);
nand U1662 (N_1662,N_1620,N_1644);
and U1663 (N_1663,N_1561,N_1535);
xnor U1664 (N_1664,N_1503,N_1529);
nand U1665 (N_1665,N_1567,N_1585);
or U1666 (N_1666,N_1523,N_1539);
nor U1667 (N_1667,N_1522,N_1548);
or U1668 (N_1668,N_1614,N_1571);
nor U1669 (N_1669,N_1621,N_1517);
or U1670 (N_1670,N_1536,N_1575);
nor U1671 (N_1671,N_1609,N_1583);
nor U1672 (N_1672,N_1627,N_1504);
or U1673 (N_1673,N_1591,N_1537);
nor U1674 (N_1674,N_1510,N_1610);
nand U1675 (N_1675,N_1532,N_1559);
xor U1676 (N_1676,N_1602,N_1632);
nand U1677 (N_1677,N_1540,N_1568);
xor U1678 (N_1678,N_1546,N_1649);
xnor U1679 (N_1679,N_1607,N_1639);
and U1680 (N_1680,N_1601,N_1576);
and U1681 (N_1681,N_1573,N_1611);
xnor U1682 (N_1682,N_1500,N_1586);
nand U1683 (N_1683,N_1584,N_1553);
and U1684 (N_1684,N_1633,N_1506);
nor U1685 (N_1685,N_1519,N_1524);
nand U1686 (N_1686,N_1518,N_1508);
or U1687 (N_1687,N_1555,N_1623);
xnor U1688 (N_1688,N_1543,N_1596);
nor U1689 (N_1689,N_1622,N_1581);
nor U1690 (N_1690,N_1578,N_1516);
or U1691 (N_1691,N_1589,N_1646);
and U1692 (N_1692,N_1641,N_1515);
nand U1693 (N_1693,N_1511,N_1530);
nand U1694 (N_1694,N_1605,N_1634);
nor U1695 (N_1695,N_1542,N_1526);
or U1696 (N_1696,N_1501,N_1648);
xnor U1697 (N_1697,N_1579,N_1635);
or U1698 (N_1698,N_1618,N_1574);
or U1699 (N_1699,N_1565,N_1538);
nor U1700 (N_1700,N_1558,N_1608);
and U1701 (N_1701,N_1593,N_1514);
nand U1702 (N_1702,N_1612,N_1592);
or U1703 (N_1703,N_1525,N_1521);
nor U1704 (N_1704,N_1509,N_1549);
and U1705 (N_1705,N_1556,N_1502);
or U1706 (N_1706,N_1552,N_1599);
nor U1707 (N_1707,N_1533,N_1624);
or U1708 (N_1708,N_1544,N_1531);
xnor U1709 (N_1709,N_1570,N_1541);
xnor U1710 (N_1710,N_1600,N_1527);
or U1711 (N_1711,N_1564,N_1580);
nor U1712 (N_1712,N_1520,N_1513);
nand U1713 (N_1713,N_1595,N_1587);
and U1714 (N_1714,N_1582,N_1604);
or U1715 (N_1715,N_1534,N_1551);
xnor U1716 (N_1716,N_1505,N_1598);
xnor U1717 (N_1717,N_1507,N_1629);
nor U1718 (N_1718,N_1619,N_1603);
and U1719 (N_1719,N_1626,N_1645);
and U1720 (N_1720,N_1566,N_1597);
and U1721 (N_1721,N_1572,N_1560);
nand U1722 (N_1722,N_1594,N_1643);
nand U1723 (N_1723,N_1642,N_1615);
xnor U1724 (N_1724,N_1554,N_1616);
xnor U1725 (N_1725,N_1506,N_1507);
xnor U1726 (N_1726,N_1582,N_1608);
and U1727 (N_1727,N_1644,N_1621);
and U1728 (N_1728,N_1637,N_1614);
and U1729 (N_1729,N_1615,N_1607);
xnor U1730 (N_1730,N_1574,N_1503);
nand U1731 (N_1731,N_1503,N_1594);
and U1732 (N_1732,N_1594,N_1579);
nor U1733 (N_1733,N_1601,N_1523);
xnor U1734 (N_1734,N_1517,N_1593);
nand U1735 (N_1735,N_1577,N_1539);
nand U1736 (N_1736,N_1634,N_1581);
nor U1737 (N_1737,N_1545,N_1552);
and U1738 (N_1738,N_1621,N_1628);
nor U1739 (N_1739,N_1554,N_1530);
and U1740 (N_1740,N_1577,N_1636);
xnor U1741 (N_1741,N_1515,N_1596);
or U1742 (N_1742,N_1506,N_1611);
or U1743 (N_1743,N_1521,N_1623);
nand U1744 (N_1744,N_1505,N_1636);
or U1745 (N_1745,N_1597,N_1507);
xor U1746 (N_1746,N_1559,N_1540);
xnor U1747 (N_1747,N_1531,N_1586);
nor U1748 (N_1748,N_1593,N_1537);
nand U1749 (N_1749,N_1597,N_1551);
nor U1750 (N_1750,N_1557,N_1518);
or U1751 (N_1751,N_1550,N_1567);
and U1752 (N_1752,N_1619,N_1632);
or U1753 (N_1753,N_1547,N_1504);
or U1754 (N_1754,N_1515,N_1643);
nand U1755 (N_1755,N_1599,N_1511);
xnor U1756 (N_1756,N_1613,N_1545);
nor U1757 (N_1757,N_1586,N_1610);
or U1758 (N_1758,N_1586,N_1570);
nand U1759 (N_1759,N_1527,N_1529);
xor U1760 (N_1760,N_1630,N_1633);
xor U1761 (N_1761,N_1581,N_1527);
nand U1762 (N_1762,N_1551,N_1520);
or U1763 (N_1763,N_1522,N_1640);
and U1764 (N_1764,N_1615,N_1567);
or U1765 (N_1765,N_1553,N_1540);
nor U1766 (N_1766,N_1599,N_1639);
and U1767 (N_1767,N_1603,N_1501);
nor U1768 (N_1768,N_1648,N_1584);
nor U1769 (N_1769,N_1577,N_1614);
xor U1770 (N_1770,N_1549,N_1648);
nand U1771 (N_1771,N_1621,N_1602);
nor U1772 (N_1772,N_1600,N_1573);
xor U1773 (N_1773,N_1647,N_1612);
and U1774 (N_1774,N_1565,N_1598);
nand U1775 (N_1775,N_1555,N_1584);
nand U1776 (N_1776,N_1506,N_1554);
nand U1777 (N_1777,N_1578,N_1551);
xor U1778 (N_1778,N_1539,N_1553);
or U1779 (N_1779,N_1609,N_1547);
and U1780 (N_1780,N_1574,N_1649);
and U1781 (N_1781,N_1584,N_1559);
nand U1782 (N_1782,N_1578,N_1632);
or U1783 (N_1783,N_1503,N_1649);
xnor U1784 (N_1784,N_1550,N_1641);
nor U1785 (N_1785,N_1520,N_1514);
nor U1786 (N_1786,N_1558,N_1575);
and U1787 (N_1787,N_1574,N_1617);
or U1788 (N_1788,N_1612,N_1566);
nand U1789 (N_1789,N_1527,N_1602);
nor U1790 (N_1790,N_1581,N_1556);
and U1791 (N_1791,N_1546,N_1611);
and U1792 (N_1792,N_1607,N_1634);
xnor U1793 (N_1793,N_1596,N_1568);
nor U1794 (N_1794,N_1572,N_1569);
and U1795 (N_1795,N_1579,N_1639);
nor U1796 (N_1796,N_1597,N_1633);
nor U1797 (N_1797,N_1577,N_1529);
xor U1798 (N_1798,N_1582,N_1539);
or U1799 (N_1799,N_1603,N_1546);
and U1800 (N_1800,N_1676,N_1757);
and U1801 (N_1801,N_1754,N_1798);
xnor U1802 (N_1802,N_1679,N_1701);
or U1803 (N_1803,N_1751,N_1716);
and U1804 (N_1804,N_1710,N_1695);
nor U1805 (N_1805,N_1731,N_1721);
xor U1806 (N_1806,N_1720,N_1660);
nand U1807 (N_1807,N_1692,N_1665);
and U1808 (N_1808,N_1683,N_1765);
nor U1809 (N_1809,N_1717,N_1699);
nand U1810 (N_1810,N_1688,N_1653);
nand U1811 (N_1811,N_1714,N_1745);
or U1812 (N_1812,N_1746,N_1680);
xnor U1813 (N_1813,N_1758,N_1666);
nand U1814 (N_1814,N_1777,N_1749);
nor U1815 (N_1815,N_1691,N_1671);
or U1816 (N_1816,N_1755,N_1743);
nand U1817 (N_1817,N_1764,N_1693);
xor U1818 (N_1818,N_1667,N_1791);
or U1819 (N_1819,N_1664,N_1654);
xor U1820 (N_1820,N_1769,N_1711);
xnor U1821 (N_1821,N_1674,N_1651);
or U1822 (N_1822,N_1744,N_1696);
and U1823 (N_1823,N_1727,N_1685);
xor U1824 (N_1824,N_1793,N_1786);
nor U1825 (N_1825,N_1737,N_1663);
xor U1826 (N_1826,N_1707,N_1787);
or U1827 (N_1827,N_1734,N_1658);
xnor U1828 (N_1828,N_1778,N_1706);
nor U1829 (N_1829,N_1713,N_1715);
nor U1830 (N_1830,N_1726,N_1760);
nor U1831 (N_1831,N_1704,N_1750);
nand U1832 (N_1832,N_1759,N_1729);
and U1833 (N_1833,N_1742,N_1681);
or U1834 (N_1834,N_1762,N_1700);
nand U1835 (N_1835,N_1669,N_1752);
or U1836 (N_1836,N_1718,N_1687);
and U1837 (N_1837,N_1738,N_1686);
or U1838 (N_1838,N_1799,N_1797);
xnor U1839 (N_1839,N_1728,N_1652);
and U1840 (N_1840,N_1668,N_1735);
and U1841 (N_1841,N_1719,N_1795);
xnor U1842 (N_1842,N_1741,N_1689);
nor U1843 (N_1843,N_1661,N_1766);
and U1844 (N_1844,N_1698,N_1672);
or U1845 (N_1845,N_1730,N_1771);
and U1846 (N_1846,N_1748,N_1781);
nor U1847 (N_1847,N_1772,N_1712);
nor U1848 (N_1848,N_1670,N_1677);
nand U1849 (N_1849,N_1723,N_1790);
xor U1850 (N_1850,N_1775,N_1767);
nor U1851 (N_1851,N_1770,N_1655);
and U1852 (N_1852,N_1656,N_1733);
or U1853 (N_1853,N_1753,N_1708);
or U1854 (N_1854,N_1794,N_1773);
nand U1855 (N_1855,N_1709,N_1784);
or U1856 (N_1856,N_1650,N_1684);
xor U1857 (N_1857,N_1739,N_1675);
and U1858 (N_1858,N_1780,N_1782);
or U1859 (N_1859,N_1705,N_1659);
or U1860 (N_1860,N_1747,N_1732);
nor U1861 (N_1861,N_1788,N_1796);
nor U1862 (N_1862,N_1756,N_1768);
nand U1863 (N_1863,N_1690,N_1761);
nor U1864 (N_1864,N_1792,N_1776);
or U1865 (N_1865,N_1662,N_1789);
nand U1866 (N_1866,N_1682,N_1722);
nor U1867 (N_1867,N_1779,N_1736);
or U1868 (N_1868,N_1657,N_1783);
or U1869 (N_1869,N_1725,N_1694);
and U1870 (N_1870,N_1785,N_1740);
and U1871 (N_1871,N_1763,N_1724);
nor U1872 (N_1872,N_1673,N_1774);
xnor U1873 (N_1873,N_1703,N_1697);
xnor U1874 (N_1874,N_1678,N_1702);
xnor U1875 (N_1875,N_1726,N_1776);
nor U1876 (N_1876,N_1691,N_1752);
nor U1877 (N_1877,N_1674,N_1700);
nor U1878 (N_1878,N_1734,N_1754);
or U1879 (N_1879,N_1718,N_1796);
xnor U1880 (N_1880,N_1724,N_1676);
or U1881 (N_1881,N_1779,N_1670);
nor U1882 (N_1882,N_1672,N_1747);
nand U1883 (N_1883,N_1697,N_1744);
and U1884 (N_1884,N_1716,N_1738);
xnor U1885 (N_1885,N_1717,N_1760);
and U1886 (N_1886,N_1665,N_1726);
and U1887 (N_1887,N_1792,N_1746);
nor U1888 (N_1888,N_1694,N_1777);
nand U1889 (N_1889,N_1709,N_1795);
xor U1890 (N_1890,N_1662,N_1749);
and U1891 (N_1891,N_1756,N_1690);
nor U1892 (N_1892,N_1782,N_1783);
or U1893 (N_1893,N_1694,N_1798);
xor U1894 (N_1894,N_1759,N_1668);
xor U1895 (N_1895,N_1714,N_1730);
xnor U1896 (N_1896,N_1794,N_1797);
nor U1897 (N_1897,N_1786,N_1664);
or U1898 (N_1898,N_1657,N_1722);
xnor U1899 (N_1899,N_1730,N_1796);
xor U1900 (N_1900,N_1668,N_1693);
nor U1901 (N_1901,N_1675,N_1790);
nand U1902 (N_1902,N_1713,N_1772);
nand U1903 (N_1903,N_1790,N_1667);
xor U1904 (N_1904,N_1779,N_1682);
or U1905 (N_1905,N_1687,N_1779);
nand U1906 (N_1906,N_1799,N_1683);
and U1907 (N_1907,N_1699,N_1698);
and U1908 (N_1908,N_1729,N_1777);
and U1909 (N_1909,N_1795,N_1686);
or U1910 (N_1910,N_1702,N_1766);
or U1911 (N_1911,N_1760,N_1707);
or U1912 (N_1912,N_1698,N_1784);
or U1913 (N_1913,N_1672,N_1721);
nor U1914 (N_1914,N_1796,N_1779);
nor U1915 (N_1915,N_1653,N_1784);
nor U1916 (N_1916,N_1740,N_1748);
nand U1917 (N_1917,N_1685,N_1745);
or U1918 (N_1918,N_1735,N_1675);
xor U1919 (N_1919,N_1721,N_1660);
or U1920 (N_1920,N_1757,N_1732);
xor U1921 (N_1921,N_1769,N_1779);
nor U1922 (N_1922,N_1790,N_1751);
xor U1923 (N_1923,N_1795,N_1769);
or U1924 (N_1924,N_1676,N_1768);
nand U1925 (N_1925,N_1712,N_1708);
nand U1926 (N_1926,N_1696,N_1699);
nor U1927 (N_1927,N_1672,N_1668);
nor U1928 (N_1928,N_1753,N_1699);
nand U1929 (N_1929,N_1683,N_1734);
nand U1930 (N_1930,N_1707,N_1690);
nand U1931 (N_1931,N_1738,N_1652);
nand U1932 (N_1932,N_1722,N_1747);
or U1933 (N_1933,N_1726,N_1656);
or U1934 (N_1934,N_1789,N_1752);
or U1935 (N_1935,N_1697,N_1767);
or U1936 (N_1936,N_1775,N_1756);
xor U1937 (N_1937,N_1795,N_1758);
nand U1938 (N_1938,N_1791,N_1676);
nor U1939 (N_1939,N_1672,N_1650);
and U1940 (N_1940,N_1695,N_1701);
xor U1941 (N_1941,N_1785,N_1745);
xor U1942 (N_1942,N_1719,N_1798);
xnor U1943 (N_1943,N_1720,N_1782);
xor U1944 (N_1944,N_1782,N_1772);
and U1945 (N_1945,N_1680,N_1716);
and U1946 (N_1946,N_1724,N_1695);
and U1947 (N_1947,N_1703,N_1685);
and U1948 (N_1948,N_1671,N_1685);
or U1949 (N_1949,N_1766,N_1724);
or U1950 (N_1950,N_1936,N_1806);
and U1951 (N_1951,N_1890,N_1938);
nor U1952 (N_1952,N_1843,N_1895);
xor U1953 (N_1953,N_1876,N_1860);
xnor U1954 (N_1954,N_1852,N_1830);
nor U1955 (N_1955,N_1865,N_1897);
xor U1956 (N_1956,N_1904,N_1811);
nor U1957 (N_1957,N_1947,N_1834);
and U1958 (N_1958,N_1882,N_1823);
or U1959 (N_1959,N_1845,N_1828);
nor U1960 (N_1960,N_1920,N_1912);
xnor U1961 (N_1961,N_1846,N_1878);
and U1962 (N_1962,N_1923,N_1937);
or U1963 (N_1963,N_1856,N_1867);
xnor U1964 (N_1964,N_1911,N_1859);
xor U1965 (N_1965,N_1939,N_1837);
or U1966 (N_1966,N_1822,N_1909);
and U1967 (N_1967,N_1864,N_1930);
xnor U1968 (N_1968,N_1941,N_1933);
xnor U1969 (N_1969,N_1889,N_1879);
or U1970 (N_1970,N_1922,N_1863);
xnor U1971 (N_1971,N_1894,N_1929);
nor U1972 (N_1972,N_1943,N_1872);
and U1973 (N_1973,N_1824,N_1841);
or U1974 (N_1974,N_1862,N_1858);
nand U1975 (N_1975,N_1942,N_1944);
nor U1976 (N_1976,N_1928,N_1807);
or U1977 (N_1977,N_1839,N_1883);
nand U1978 (N_1978,N_1836,N_1910);
and U1979 (N_1979,N_1813,N_1935);
and U1980 (N_1980,N_1926,N_1848);
xnor U1981 (N_1981,N_1888,N_1868);
nor U1982 (N_1982,N_1869,N_1857);
nand U1983 (N_1983,N_1877,N_1932);
and U1984 (N_1984,N_1840,N_1927);
and U1985 (N_1985,N_1825,N_1919);
nor U1986 (N_1986,N_1940,N_1898);
xor U1987 (N_1987,N_1908,N_1896);
or U1988 (N_1988,N_1832,N_1918);
or U1989 (N_1989,N_1853,N_1816);
xor U1990 (N_1990,N_1885,N_1916);
or U1991 (N_1991,N_1871,N_1861);
or U1992 (N_1992,N_1875,N_1847);
and U1993 (N_1993,N_1924,N_1917);
nor U1994 (N_1994,N_1945,N_1907);
and U1995 (N_1995,N_1948,N_1804);
or U1996 (N_1996,N_1854,N_1842);
nor U1997 (N_1997,N_1814,N_1906);
nand U1998 (N_1998,N_1826,N_1835);
nand U1999 (N_1999,N_1809,N_1892);
nand U2000 (N_2000,N_1902,N_1915);
nor U2001 (N_2001,N_1905,N_1866);
or U2002 (N_2002,N_1899,N_1844);
or U2003 (N_2003,N_1821,N_1913);
nand U2004 (N_2004,N_1870,N_1815);
and U2005 (N_2005,N_1817,N_1808);
xnor U2006 (N_2006,N_1874,N_1921);
nand U2007 (N_2007,N_1833,N_1802);
nand U2008 (N_2008,N_1800,N_1803);
and U2009 (N_2009,N_1886,N_1934);
or U2010 (N_2010,N_1903,N_1801);
xor U2011 (N_2011,N_1949,N_1901);
xor U2012 (N_2012,N_1812,N_1900);
xnor U2013 (N_2013,N_1925,N_1880);
xnor U2014 (N_2014,N_1851,N_1873);
or U2015 (N_2015,N_1849,N_1887);
and U2016 (N_2016,N_1881,N_1850);
or U2017 (N_2017,N_1931,N_1893);
nor U2018 (N_2018,N_1946,N_1829);
and U2019 (N_2019,N_1914,N_1827);
and U2020 (N_2020,N_1819,N_1805);
xnor U2021 (N_2021,N_1831,N_1820);
or U2022 (N_2022,N_1855,N_1818);
nand U2023 (N_2023,N_1891,N_1810);
nor U2024 (N_2024,N_1884,N_1838);
nor U2025 (N_2025,N_1825,N_1803);
nor U2026 (N_2026,N_1815,N_1823);
and U2027 (N_2027,N_1931,N_1939);
nor U2028 (N_2028,N_1866,N_1892);
nor U2029 (N_2029,N_1880,N_1855);
and U2030 (N_2030,N_1884,N_1850);
and U2031 (N_2031,N_1802,N_1901);
and U2032 (N_2032,N_1894,N_1912);
nor U2033 (N_2033,N_1914,N_1824);
or U2034 (N_2034,N_1801,N_1920);
and U2035 (N_2035,N_1943,N_1949);
nand U2036 (N_2036,N_1935,N_1850);
and U2037 (N_2037,N_1828,N_1854);
nor U2038 (N_2038,N_1826,N_1930);
or U2039 (N_2039,N_1882,N_1806);
or U2040 (N_2040,N_1899,N_1888);
nand U2041 (N_2041,N_1894,N_1938);
or U2042 (N_2042,N_1848,N_1883);
nor U2043 (N_2043,N_1902,N_1801);
xor U2044 (N_2044,N_1904,N_1882);
and U2045 (N_2045,N_1941,N_1918);
nor U2046 (N_2046,N_1889,N_1813);
xor U2047 (N_2047,N_1849,N_1848);
nor U2048 (N_2048,N_1928,N_1919);
and U2049 (N_2049,N_1825,N_1933);
nor U2050 (N_2050,N_1862,N_1868);
nor U2051 (N_2051,N_1916,N_1933);
xnor U2052 (N_2052,N_1828,N_1849);
or U2053 (N_2053,N_1821,N_1910);
or U2054 (N_2054,N_1882,N_1903);
or U2055 (N_2055,N_1908,N_1947);
nor U2056 (N_2056,N_1893,N_1812);
nand U2057 (N_2057,N_1879,N_1880);
and U2058 (N_2058,N_1829,N_1836);
nand U2059 (N_2059,N_1815,N_1873);
and U2060 (N_2060,N_1805,N_1816);
xor U2061 (N_2061,N_1888,N_1866);
nor U2062 (N_2062,N_1845,N_1807);
or U2063 (N_2063,N_1850,N_1825);
xnor U2064 (N_2064,N_1849,N_1814);
or U2065 (N_2065,N_1941,N_1807);
xnor U2066 (N_2066,N_1850,N_1810);
and U2067 (N_2067,N_1929,N_1861);
nor U2068 (N_2068,N_1876,N_1866);
or U2069 (N_2069,N_1832,N_1897);
nand U2070 (N_2070,N_1846,N_1848);
xnor U2071 (N_2071,N_1876,N_1948);
and U2072 (N_2072,N_1920,N_1862);
nor U2073 (N_2073,N_1832,N_1947);
nand U2074 (N_2074,N_1812,N_1833);
or U2075 (N_2075,N_1802,N_1889);
nand U2076 (N_2076,N_1934,N_1918);
xnor U2077 (N_2077,N_1892,N_1896);
or U2078 (N_2078,N_1807,N_1939);
nand U2079 (N_2079,N_1826,N_1875);
or U2080 (N_2080,N_1900,N_1802);
and U2081 (N_2081,N_1830,N_1939);
and U2082 (N_2082,N_1841,N_1835);
nand U2083 (N_2083,N_1941,N_1879);
and U2084 (N_2084,N_1896,N_1926);
and U2085 (N_2085,N_1838,N_1873);
xnor U2086 (N_2086,N_1833,N_1819);
and U2087 (N_2087,N_1825,N_1881);
xor U2088 (N_2088,N_1944,N_1853);
nand U2089 (N_2089,N_1872,N_1827);
xnor U2090 (N_2090,N_1821,N_1923);
xnor U2091 (N_2091,N_1862,N_1897);
and U2092 (N_2092,N_1832,N_1902);
and U2093 (N_2093,N_1944,N_1915);
nand U2094 (N_2094,N_1847,N_1893);
nor U2095 (N_2095,N_1926,N_1924);
or U2096 (N_2096,N_1874,N_1840);
and U2097 (N_2097,N_1808,N_1920);
nor U2098 (N_2098,N_1816,N_1890);
xor U2099 (N_2099,N_1933,N_1899);
nor U2100 (N_2100,N_2020,N_2008);
xnor U2101 (N_2101,N_2021,N_2040);
and U2102 (N_2102,N_2070,N_2047);
or U2103 (N_2103,N_1997,N_2050);
and U2104 (N_2104,N_1993,N_2066);
nor U2105 (N_2105,N_2005,N_2063);
or U2106 (N_2106,N_1996,N_2089);
or U2107 (N_2107,N_2095,N_2034);
xnor U2108 (N_2108,N_2011,N_2002);
xor U2109 (N_2109,N_2012,N_2004);
xor U2110 (N_2110,N_2057,N_1989);
or U2111 (N_2111,N_2019,N_2078);
or U2112 (N_2112,N_2077,N_1965);
or U2113 (N_2113,N_2056,N_2052);
xor U2114 (N_2114,N_2017,N_2069);
xnor U2115 (N_2115,N_2007,N_2053);
nor U2116 (N_2116,N_2080,N_2096);
and U2117 (N_2117,N_1950,N_2054);
and U2118 (N_2118,N_1983,N_2009);
nand U2119 (N_2119,N_2055,N_2046);
and U2120 (N_2120,N_1964,N_2068);
nor U2121 (N_2121,N_2072,N_1972);
and U2122 (N_2122,N_2093,N_1977);
nor U2123 (N_2123,N_2031,N_1969);
and U2124 (N_2124,N_2058,N_2075);
xnor U2125 (N_2125,N_2044,N_2006);
nand U2126 (N_2126,N_2028,N_2084);
nor U2127 (N_2127,N_1970,N_2082);
xnor U2128 (N_2128,N_1981,N_2092);
or U2129 (N_2129,N_1985,N_2043);
nand U2130 (N_2130,N_2045,N_1971);
and U2131 (N_2131,N_2000,N_2098);
xnor U2132 (N_2132,N_2099,N_2003);
nor U2133 (N_2133,N_2027,N_2010);
nand U2134 (N_2134,N_1952,N_1987);
nor U2135 (N_2135,N_1962,N_2024);
nor U2136 (N_2136,N_2087,N_1956);
and U2137 (N_2137,N_1973,N_1999);
nor U2138 (N_2138,N_2036,N_2064);
or U2139 (N_2139,N_1951,N_2059);
nor U2140 (N_2140,N_1998,N_1984);
xor U2141 (N_2141,N_2094,N_1995);
nor U2142 (N_2142,N_1992,N_1974);
and U2143 (N_2143,N_1958,N_1953);
and U2144 (N_2144,N_2039,N_2025);
and U2145 (N_2145,N_1982,N_2097);
nor U2146 (N_2146,N_1959,N_2014);
and U2147 (N_2147,N_2016,N_1975);
or U2148 (N_2148,N_2088,N_1967);
xor U2149 (N_2149,N_2001,N_1991);
nand U2150 (N_2150,N_2030,N_1961);
nand U2151 (N_2151,N_1980,N_1994);
nor U2152 (N_2152,N_2090,N_2065);
or U2153 (N_2153,N_2091,N_2074);
nand U2154 (N_2154,N_1966,N_2018);
or U2155 (N_2155,N_2041,N_1979);
nor U2156 (N_2156,N_1990,N_2042);
or U2157 (N_2157,N_2029,N_1955);
xor U2158 (N_2158,N_1986,N_2026);
or U2159 (N_2159,N_2022,N_2049);
xnor U2160 (N_2160,N_1960,N_1957);
or U2161 (N_2161,N_2073,N_1978);
and U2162 (N_2162,N_2081,N_2013);
xor U2163 (N_2163,N_2051,N_2085);
nand U2164 (N_2164,N_2038,N_2083);
or U2165 (N_2165,N_2076,N_2067);
nor U2166 (N_2166,N_2032,N_2033);
and U2167 (N_2167,N_1976,N_2035);
xnor U2168 (N_2168,N_2062,N_1963);
or U2169 (N_2169,N_2071,N_1954);
and U2170 (N_2170,N_2037,N_2086);
and U2171 (N_2171,N_2015,N_2060);
and U2172 (N_2172,N_1968,N_2048);
nor U2173 (N_2173,N_1988,N_2061);
or U2174 (N_2174,N_2023,N_2079);
nand U2175 (N_2175,N_1990,N_2011);
or U2176 (N_2176,N_2027,N_1990);
nor U2177 (N_2177,N_1989,N_2063);
or U2178 (N_2178,N_2069,N_1955);
and U2179 (N_2179,N_2018,N_1951);
and U2180 (N_2180,N_2028,N_2057);
nor U2181 (N_2181,N_1966,N_2079);
and U2182 (N_2182,N_1994,N_2003);
and U2183 (N_2183,N_2020,N_2070);
or U2184 (N_2184,N_1988,N_2024);
nor U2185 (N_2185,N_2041,N_1976);
or U2186 (N_2186,N_2092,N_1959);
or U2187 (N_2187,N_1976,N_2007);
and U2188 (N_2188,N_1996,N_1977);
and U2189 (N_2189,N_1970,N_2078);
nor U2190 (N_2190,N_2084,N_2017);
or U2191 (N_2191,N_2054,N_2048);
nand U2192 (N_2192,N_2068,N_2074);
or U2193 (N_2193,N_2040,N_2068);
xnor U2194 (N_2194,N_2025,N_1977);
nand U2195 (N_2195,N_2064,N_2056);
nand U2196 (N_2196,N_1996,N_2011);
xor U2197 (N_2197,N_2091,N_1992);
and U2198 (N_2198,N_1965,N_2097);
nand U2199 (N_2199,N_1954,N_1960);
xnor U2200 (N_2200,N_2041,N_2080);
xor U2201 (N_2201,N_2045,N_2048);
nand U2202 (N_2202,N_2095,N_2071);
or U2203 (N_2203,N_2044,N_1991);
nor U2204 (N_2204,N_2051,N_2039);
nor U2205 (N_2205,N_2034,N_2057);
and U2206 (N_2206,N_2036,N_2048);
nor U2207 (N_2207,N_1997,N_1952);
xnor U2208 (N_2208,N_1986,N_1962);
nand U2209 (N_2209,N_1982,N_2030);
xnor U2210 (N_2210,N_2086,N_2055);
nor U2211 (N_2211,N_2034,N_2042);
or U2212 (N_2212,N_1955,N_1975);
xor U2213 (N_2213,N_1999,N_2000);
nand U2214 (N_2214,N_1971,N_2068);
nor U2215 (N_2215,N_2030,N_2083);
or U2216 (N_2216,N_1998,N_2084);
and U2217 (N_2217,N_1990,N_2043);
or U2218 (N_2218,N_1987,N_1980);
nand U2219 (N_2219,N_1955,N_1979);
nand U2220 (N_2220,N_2049,N_2070);
nand U2221 (N_2221,N_2059,N_1999);
and U2222 (N_2222,N_2033,N_2040);
and U2223 (N_2223,N_1960,N_1981);
or U2224 (N_2224,N_1971,N_1999);
nor U2225 (N_2225,N_2061,N_2030);
nand U2226 (N_2226,N_2023,N_2092);
nand U2227 (N_2227,N_2031,N_1987);
nand U2228 (N_2228,N_2091,N_2098);
and U2229 (N_2229,N_2049,N_2078);
xnor U2230 (N_2230,N_2013,N_2098);
nand U2231 (N_2231,N_2039,N_2002);
nor U2232 (N_2232,N_2063,N_1995);
xor U2233 (N_2233,N_2059,N_2096);
xor U2234 (N_2234,N_1999,N_2077);
and U2235 (N_2235,N_1998,N_2021);
xnor U2236 (N_2236,N_1974,N_2074);
xor U2237 (N_2237,N_2021,N_2020);
nor U2238 (N_2238,N_1995,N_2011);
nand U2239 (N_2239,N_1985,N_2078);
nand U2240 (N_2240,N_1962,N_2014);
or U2241 (N_2241,N_2054,N_1970);
nor U2242 (N_2242,N_2066,N_1974);
nand U2243 (N_2243,N_2051,N_1995);
and U2244 (N_2244,N_2041,N_1972);
xnor U2245 (N_2245,N_1993,N_2016);
or U2246 (N_2246,N_2024,N_1965);
nand U2247 (N_2247,N_2073,N_2022);
xnor U2248 (N_2248,N_2068,N_1984);
or U2249 (N_2249,N_1971,N_1968);
or U2250 (N_2250,N_2166,N_2186);
xnor U2251 (N_2251,N_2122,N_2191);
nor U2252 (N_2252,N_2185,N_2106);
or U2253 (N_2253,N_2206,N_2182);
or U2254 (N_2254,N_2107,N_2142);
nand U2255 (N_2255,N_2203,N_2123);
and U2256 (N_2256,N_2118,N_2180);
nor U2257 (N_2257,N_2162,N_2226);
xnor U2258 (N_2258,N_2228,N_2225);
nand U2259 (N_2259,N_2101,N_2109);
nand U2260 (N_2260,N_2183,N_2159);
nor U2261 (N_2261,N_2113,N_2157);
and U2262 (N_2262,N_2156,N_2194);
nor U2263 (N_2263,N_2189,N_2136);
xnor U2264 (N_2264,N_2140,N_2235);
nand U2265 (N_2265,N_2120,N_2103);
and U2266 (N_2266,N_2193,N_2211);
nor U2267 (N_2267,N_2212,N_2128);
or U2268 (N_2268,N_2131,N_2223);
xor U2269 (N_2269,N_2126,N_2217);
xnor U2270 (N_2270,N_2190,N_2207);
nor U2271 (N_2271,N_2139,N_2124);
or U2272 (N_2272,N_2143,N_2213);
xnor U2273 (N_2273,N_2249,N_2174);
nor U2274 (N_2274,N_2239,N_2167);
nand U2275 (N_2275,N_2112,N_2165);
or U2276 (N_2276,N_2234,N_2192);
nor U2277 (N_2277,N_2229,N_2246);
or U2278 (N_2278,N_2148,N_2121);
nor U2279 (N_2279,N_2104,N_2222);
and U2280 (N_2280,N_2144,N_2176);
or U2281 (N_2281,N_2134,N_2154);
or U2282 (N_2282,N_2117,N_2169);
and U2283 (N_2283,N_2163,N_2153);
and U2284 (N_2284,N_2114,N_2178);
and U2285 (N_2285,N_2218,N_2237);
or U2286 (N_2286,N_2158,N_2119);
nor U2287 (N_2287,N_2138,N_2227);
xor U2288 (N_2288,N_2147,N_2108);
nor U2289 (N_2289,N_2184,N_2236);
nor U2290 (N_2290,N_2232,N_2129);
xor U2291 (N_2291,N_2146,N_2164);
nand U2292 (N_2292,N_2177,N_2132);
nor U2293 (N_2293,N_2245,N_2125);
nand U2294 (N_2294,N_2170,N_2208);
and U2295 (N_2295,N_2248,N_2155);
xnor U2296 (N_2296,N_2243,N_2205);
nand U2297 (N_2297,N_2247,N_2149);
and U2298 (N_2298,N_2102,N_2224);
and U2299 (N_2299,N_2199,N_2111);
and U2300 (N_2300,N_2116,N_2209);
or U2301 (N_2301,N_2238,N_2141);
nand U2302 (N_2302,N_2127,N_2145);
xnor U2303 (N_2303,N_2171,N_2214);
nor U2304 (N_2304,N_2150,N_2100);
nand U2305 (N_2305,N_2197,N_2220);
nor U2306 (N_2306,N_2216,N_2179);
nand U2307 (N_2307,N_2231,N_2133);
or U2308 (N_2308,N_2161,N_2233);
xor U2309 (N_2309,N_2188,N_2137);
or U2310 (N_2310,N_2196,N_2215);
and U2311 (N_2311,N_2219,N_2105);
xor U2312 (N_2312,N_2160,N_2201);
xnor U2313 (N_2313,N_2172,N_2244);
nor U2314 (N_2314,N_2241,N_2195);
nand U2315 (N_2315,N_2230,N_2135);
xor U2316 (N_2316,N_2115,N_2202);
or U2317 (N_2317,N_2240,N_2210);
nor U2318 (N_2318,N_2152,N_2187);
nor U2319 (N_2319,N_2130,N_2110);
or U2320 (N_2320,N_2221,N_2204);
nor U2321 (N_2321,N_2168,N_2200);
nor U2322 (N_2322,N_2198,N_2173);
or U2323 (N_2323,N_2242,N_2151);
and U2324 (N_2324,N_2175,N_2181);
or U2325 (N_2325,N_2242,N_2222);
nand U2326 (N_2326,N_2242,N_2202);
and U2327 (N_2327,N_2131,N_2156);
xor U2328 (N_2328,N_2188,N_2156);
and U2329 (N_2329,N_2186,N_2126);
and U2330 (N_2330,N_2108,N_2223);
and U2331 (N_2331,N_2170,N_2222);
and U2332 (N_2332,N_2198,N_2234);
xor U2333 (N_2333,N_2141,N_2112);
nor U2334 (N_2334,N_2164,N_2204);
and U2335 (N_2335,N_2226,N_2221);
nand U2336 (N_2336,N_2170,N_2102);
and U2337 (N_2337,N_2195,N_2129);
xor U2338 (N_2338,N_2153,N_2223);
nand U2339 (N_2339,N_2137,N_2178);
nor U2340 (N_2340,N_2107,N_2141);
nand U2341 (N_2341,N_2249,N_2129);
nand U2342 (N_2342,N_2183,N_2190);
nand U2343 (N_2343,N_2201,N_2195);
nand U2344 (N_2344,N_2186,N_2177);
and U2345 (N_2345,N_2188,N_2125);
and U2346 (N_2346,N_2176,N_2111);
xnor U2347 (N_2347,N_2135,N_2179);
nand U2348 (N_2348,N_2157,N_2135);
nor U2349 (N_2349,N_2118,N_2141);
xor U2350 (N_2350,N_2214,N_2225);
xnor U2351 (N_2351,N_2152,N_2226);
nor U2352 (N_2352,N_2232,N_2229);
xor U2353 (N_2353,N_2215,N_2171);
nand U2354 (N_2354,N_2150,N_2193);
and U2355 (N_2355,N_2196,N_2164);
nor U2356 (N_2356,N_2219,N_2162);
or U2357 (N_2357,N_2192,N_2196);
and U2358 (N_2358,N_2237,N_2248);
xor U2359 (N_2359,N_2141,N_2137);
or U2360 (N_2360,N_2169,N_2181);
or U2361 (N_2361,N_2208,N_2233);
xor U2362 (N_2362,N_2124,N_2147);
nor U2363 (N_2363,N_2176,N_2237);
nor U2364 (N_2364,N_2195,N_2209);
nor U2365 (N_2365,N_2134,N_2151);
or U2366 (N_2366,N_2152,N_2129);
xor U2367 (N_2367,N_2209,N_2183);
nor U2368 (N_2368,N_2123,N_2236);
xnor U2369 (N_2369,N_2101,N_2153);
or U2370 (N_2370,N_2120,N_2196);
nand U2371 (N_2371,N_2143,N_2120);
xor U2372 (N_2372,N_2132,N_2241);
nand U2373 (N_2373,N_2137,N_2198);
nand U2374 (N_2374,N_2247,N_2243);
nand U2375 (N_2375,N_2115,N_2235);
or U2376 (N_2376,N_2148,N_2110);
and U2377 (N_2377,N_2105,N_2197);
and U2378 (N_2378,N_2135,N_2207);
xnor U2379 (N_2379,N_2224,N_2121);
or U2380 (N_2380,N_2187,N_2234);
nor U2381 (N_2381,N_2136,N_2167);
nand U2382 (N_2382,N_2197,N_2141);
or U2383 (N_2383,N_2116,N_2230);
nor U2384 (N_2384,N_2194,N_2138);
or U2385 (N_2385,N_2176,N_2157);
and U2386 (N_2386,N_2185,N_2216);
nor U2387 (N_2387,N_2133,N_2202);
nand U2388 (N_2388,N_2157,N_2117);
and U2389 (N_2389,N_2200,N_2202);
and U2390 (N_2390,N_2191,N_2201);
and U2391 (N_2391,N_2190,N_2243);
xor U2392 (N_2392,N_2119,N_2130);
and U2393 (N_2393,N_2159,N_2116);
or U2394 (N_2394,N_2116,N_2224);
and U2395 (N_2395,N_2134,N_2123);
and U2396 (N_2396,N_2132,N_2108);
nor U2397 (N_2397,N_2160,N_2196);
or U2398 (N_2398,N_2188,N_2205);
or U2399 (N_2399,N_2223,N_2230);
nor U2400 (N_2400,N_2359,N_2395);
nand U2401 (N_2401,N_2355,N_2365);
nand U2402 (N_2402,N_2288,N_2335);
and U2403 (N_2403,N_2366,N_2367);
nor U2404 (N_2404,N_2311,N_2397);
xor U2405 (N_2405,N_2271,N_2361);
nand U2406 (N_2406,N_2347,N_2314);
nand U2407 (N_2407,N_2320,N_2298);
and U2408 (N_2408,N_2291,N_2300);
nand U2409 (N_2409,N_2254,N_2346);
nand U2410 (N_2410,N_2349,N_2313);
xnor U2411 (N_2411,N_2343,N_2356);
nor U2412 (N_2412,N_2334,N_2386);
xor U2413 (N_2413,N_2253,N_2284);
xnor U2414 (N_2414,N_2379,N_2357);
nor U2415 (N_2415,N_2360,N_2375);
and U2416 (N_2416,N_2387,N_2263);
nand U2417 (N_2417,N_2327,N_2285);
xnor U2418 (N_2418,N_2370,N_2280);
or U2419 (N_2419,N_2296,N_2260);
or U2420 (N_2420,N_2308,N_2369);
and U2421 (N_2421,N_2358,N_2388);
xor U2422 (N_2422,N_2276,N_2329);
nand U2423 (N_2423,N_2282,N_2268);
or U2424 (N_2424,N_2316,N_2303);
nand U2425 (N_2425,N_2341,N_2333);
xor U2426 (N_2426,N_2382,N_2325);
xor U2427 (N_2427,N_2378,N_2297);
or U2428 (N_2428,N_2261,N_2317);
nor U2429 (N_2429,N_2377,N_2339);
or U2430 (N_2430,N_2374,N_2337);
or U2431 (N_2431,N_2326,N_2272);
nand U2432 (N_2432,N_2390,N_2281);
nand U2433 (N_2433,N_2251,N_2302);
and U2434 (N_2434,N_2273,N_2287);
nor U2435 (N_2435,N_2352,N_2274);
nor U2436 (N_2436,N_2368,N_2362);
xor U2437 (N_2437,N_2289,N_2399);
nand U2438 (N_2438,N_2323,N_2262);
xnor U2439 (N_2439,N_2330,N_2265);
and U2440 (N_2440,N_2364,N_2348);
or U2441 (N_2441,N_2279,N_2381);
or U2442 (N_2442,N_2255,N_2315);
xor U2443 (N_2443,N_2342,N_2376);
nand U2444 (N_2444,N_2293,N_2384);
xor U2445 (N_2445,N_2385,N_2283);
nor U2446 (N_2446,N_2318,N_2340);
nand U2447 (N_2447,N_2306,N_2275);
nand U2448 (N_2448,N_2328,N_2267);
nor U2449 (N_2449,N_2324,N_2371);
xnor U2450 (N_2450,N_2295,N_2270);
nand U2451 (N_2451,N_2322,N_2389);
xnor U2452 (N_2452,N_2307,N_2312);
or U2453 (N_2453,N_2380,N_2383);
and U2454 (N_2454,N_2392,N_2373);
or U2455 (N_2455,N_2344,N_2277);
or U2456 (N_2456,N_2336,N_2372);
or U2457 (N_2457,N_2299,N_2304);
xnor U2458 (N_2458,N_2250,N_2310);
xor U2459 (N_2459,N_2294,N_2319);
nand U2460 (N_2460,N_2305,N_2257);
xor U2461 (N_2461,N_2264,N_2256);
xor U2462 (N_2462,N_2290,N_2278);
nor U2463 (N_2463,N_2350,N_2353);
and U2464 (N_2464,N_2266,N_2398);
xor U2465 (N_2465,N_2338,N_2394);
or U2466 (N_2466,N_2301,N_2396);
xnor U2467 (N_2467,N_2354,N_2321);
nor U2468 (N_2468,N_2252,N_2259);
nor U2469 (N_2469,N_2258,N_2292);
and U2470 (N_2470,N_2393,N_2309);
nand U2471 (N_2471,N_2351,N_2286);
nor U2472 (N_2472,N_2363,N_2345);
nor U2473 (N_2473,N_2391,N_2332);
or U2474 (N_2474,N_2269,N_2331);
and U2475 (N_2475,N_2321,N_2328);
and U2476 (N_2476,N_2309,N_2323);
nand U2477 (N_2477,N_2341,N_2290);
nor U2478 (N_2478,N_2334,N_2276);
nor U2479 (N_2479,N_2304,N_2307);
xor U2480 (N_2480,N_2374,N_2370);
and U2481 (N_2481,N_2346,N_2302);
nand U2482 (N_2482,N_2326,N_2346);
nor U2483 (N_2483,N_2392,N_2372);
xor U2484 (N_2484,N_2324,N_2291);
nor U2485 (N_2485,N_2258,N_2335);
and U2486 (N_2486,N_2289,N_2270);
xor U2487 (N_2487,N_2289,N_2275);
nor U2488 (N_2488,N_2278,N_2299);
and U2489 (N_2489,N_2368,N_2363);
nor U2490 (N_2490,N_2399,N_2369);
or U2491 (N_2491,N_2375,N_2350);
and U2492 (N_2492,N_2363,N_2350);
or U2493 (N_2493,N_2314,N_2275);
xor U2494 (N_2494,N_2281,N_2361);
and U2495 (N_2495,N_2344,N_2285);
xor U2496 (N_2496,N_2352,N_2258);
nand U2497 (N_2497,N_2281,N_2346);
and U2498 (N_2498,N_2308,N_2390);
xnor U2499 (N_2499,N_2269,N_2395);
nand U2500 (N_2500,N_2357,N_2380);
or U2501 (N_2501,N_2276,N_2299);
nand U2502 (N_2502,N_2376,N_2346);
or U2503 (N_2503,N_2261,N_2260);
xor U2504 (N_2504,N_2325,N_2298);
and U2505 (N_2505,N_2356,N_2370);
and U2506 (N_2506,N_2306,N_2278);
nand U2507 (N_2507,N_2264,N_2385);
or U2508 (N_2508,N_2296,N_2359);
or U2509 (N_2509,N_2329,N_2362);
and U2510 (N_2510,N_2261,N_2323);
or U2511 (N_2511,N_2303,N_2286);
or U2512 (N_2512,N_2289,N_2267);
or U2513 (N_2513,N_2368,N_2316);
xnor U2514 (N_2514,N_2355,N_2288);
xnor U2515 (N_2515,N_2296,N_2353);
nand U2516 (N_2516,N_2314,N_2298);
nand U2517 (N_2517,N_2285,N_2358);
xor U2518 (N_2518,N_2399,N_2273);
nor U2519 (N_2519,N_2277,N_2253);
nor U2520 (N_2520,N_2274,N_2266);
or U2521 (N_2521,N_2273,N_2323);
xor U2522 (N_2522,N_2358,N_2274);
xor U2523 (N_2523,N_2385,N_2393);
or U2524 (N_2524,N_2368,N_2324);
or U2525 (N_2525,N_2310,N_2379);
xnor U2526 (N_2526,N_2302,N_2303);
and U2527 (N_2527,N_2330,N_2333);
or U2528 (N_2528,N_2376,N_2341);
and U2529 (N_2529,N_2364,N_2399);
xor U2530 (N_2530,N_2349,N_2275);
and U2531 (N_2531,N_2307,N_2262);
or U2532 (N_2532,N_2357,N_2319);
nand U2533 (N_2533,N_2296,N_2264);
xor U2534 (N_2534,N_2389,N_2307);
or U2535 (N_2535,N_2370,N_2349);
and U2536 (N_2536,N_2321,N_2392);
nand U2537 (N_2537,N_2370,N_2354);
and U2538 (N_2538,N_2341,N_2340);
or U2539 (N_2539,N_2287,N_2251);
xnor U2540 (N_2540,N_2303,N_2307);
nand U2541 (N_2541,N_2254,N_2352);
nor U2542 (N_2542,N_2379,N_2265);
nand U2543 (N_2543,N_2376,N_2340);
or U2544 (N_2544,N_2340,N_2279);
or U2545 (N_2545,N_2387,N_2301);
xnor U2546 (N_2546,N_2399,N_2253);
nor U2547 (N_2547,N_2303,N_2324);
nand U2548 (N_2548,N_2324,N_2257);
xnor U2549 (N_2549,N_2399,N_2372);
nand U2550 (N_2550,N_2531,N_2450);
nor U2551 (N_2551,N_2411,N_2437);
and U2552 (N_2552,N_2544,N_2402);
nand U2553 (N_2553,N_2456,N_2533);
nand U2554 (N_2554,N_2468,N_2472);
or U2555 (N_2555,N_2503,N_2469);
and U2556 (N_2556,N_2481,N_2512);
and U2557 (N_2557,N_2463,N_2431);
nor U2558 (N_2558,N_2474,N_2541);
xor U2559 (N_2559,N_2415,N_2526);
and U2560 (N_2560,N_2521,N_2491);
or U2561 (N_2561,N_2419,N_2501);
or U2562 (N_2562,N_2455,N_2540);
nand U2563 (N_2563,N_2478,N_2420);
and U2564 (N_2564,N_2416,N_2543);
xor U2565 (N_2565,N_2404,N_2483);
xnor U2566 (N_2566,N_2485,N_2537);
and U2567 (N_2567,N_2487,N_2514);
xnor U2568 (N_2568,N_2459,N_2476);
or U2569 (N_2569,N_2434,N_2438);
and U2570 (N_2570,N_2532,N_2458);
nor U2571 (N_2571,N_2465,N_2406);
or U2572 (N_2572,N_2539,N_2418);
or U2573 (N_2573,N_2451,N_2433);
or U2574 (N_2574,N_2405,N_2546);
nor U2575 (N_2575,N_2517,N_2449);
xnor U2576 (N_2576,N_2498,N_2410);
nor U2577 (N_2577,N_2542,N_2409);
or U2578 (N_2578,N_2538,N_2453);
nor U2579 (N_2579,N_2427,N_2496);
or U2580 (N_2580,N_2482,N_2524);
or U2581 (N_2581,N_2506,N_2529);
and U2582 (N_2582,N_2549,N_2413);
or U2583 (N_2583,N_2445,N_2408);
xor U2584 (N_2584,N_2454,N_2421);
xnor U2585 (N_2585,N_2492,N_2477);
or U2586 (N_2586,N_2441,N_2403);
or U2587 (N_2587,N_2473,N_2426);
xor U2588 (N_2588,N_2432,N_2439);
or U2589 (N_2589,N_2475,N_2535);
xor U2590 (N_2590,N_2511,N_2467);
nor U2591 (N_2591,N_2490,N_2417);
nor U2592 (N_2592,N_2536,N_2446);
nor U2593 (N_2593,N_2457,N_2461);
nand U2594 (N_2594,N_2495,N_2519);
nor U2595 (N_2595,N_2429,N_2547);
xor U2596 (N_2596,N_2430,N_2488);
and U2597 (N_2597,N_2493,N_2530);
and U2598 (N_2598,N_2509,N_2407);
or U2599 (N_2599,N_2423,N_2443);
or U2600 (N_2600,N_2428,N_2422);
nand U2601 (N_2601,N_2507,N_2502);
nand U2602 (N_2602,N_2464,N_2480);
xnor U2603 (N_2603,N_2500,N_2494);
nor U2604 (N_2604,N_2401,N_2528);
and U2605 (N_2605,N_2534,N_2522);
nand U2606 (N_2606,N_2486,N_2516);
nor U2607 (N_2607,N_2425,N_2515);
and U2608 (N_2608,N_2440,N_2497);
nor U2609 (N_2609,N_2484,N_2548);
and U2610 (N_2610,N_2435,N_2545);
or U2611 (N_2611,N_2424,N_2499);
and U2612 (N_2612,N_2508,N_2520);
and U2613 (N_2613,N_2400,N_2448);
and U2614 (N_2614,N_2447,N_2479);
nor U2615 (N_2615,N_2523,N_2510);
or U2616 (N_2616,N_2466,N_2489);
xnor U2617 (N_2617,N_2505,N_2412);
nand U2618 (N_2618,N_2436,N_2442);
xor U2619 (N_2619,N_2513,N_2460);
and U2620 (N_2620,N_2470,N_2414);
and U2621 (N_2621,N_2471,N_2452);
and U2622 (N_2622,N_2527,N_2504);
nor U2623 (N_2623,N_2462,N_2444);
nor U2624 (N_2624,N_2518,N_2525);
nor U2625 (N_2625,N_2518,N_2420);
nor U2626 (N_2626,N_2426,N_2438);
nand U2627 (N_2627,N_2413,N_2535);
nand U2628 (N_2628,N_2412,N_2407);
xor U2629 (N_2629,N_2450,N_2470);
and U2630 (N_2630,N_2486,N_2535);
nor U2631 (N_2631,N_2468,N_2402);
nor U2632 (N_2632,N_2510,N_2460);
nor U2633 (N_2633,N_2502,N_2467);
or U2634 (N_2634,N_2480,N_2409);
and U2635 (N_2635,N_2497,N_2543);
and U2636 (N_2636,N_2518,N_2467);
nand U2637 (N_2637,N_2487,N_2496);
nand U2638 (N_2638,N_2515,N_2497);
nand U2639 (N_2639,N_2479,N_2513);
and U2640 (N_2640,N_2538,N_2527);
or U2641 (N_2641,N_2544,N_2463);
and U2642 (N_2642,N_2425,N_2430);
or U2643 (N_2643,N_2478,N_2466);
xnor U2644 (N_2644,N_2424,N_2492);
nand U2645 (N_2645,N_2408,N_2493);
or U2646 (N_2646,N_2514,N_2517);
and U2647 (N_2647,N_2447,N_2432);
nand U2648 (N_2648,N_2450,N_2439);
or U2649 (N_2649,N_2509,N_2505);
and U2650 (N_2650,N_2405,N_2518);
and U2651 (N_2651,N_2480,N_2483);
xor U2652 (N_2652,N_2486,N_2408);
and U2653 (N_2653,N_2416,N_2423);
nand U2654 (N_2654,N_2454,N_2548);
xnor U2655 (N_2655,N_2513,N_2464);
nor U2656 (N_2656,N_2424,N_2544);
and U2657 (N_2657,N_2499,N_2418);
or U2658 (N_2658,N_2539,N_2496);
xor U2659 (N_2659,N_2503,N_2484);
xor U2660 (N_2660,N_2490,N_2483);
and U2661 (N_2661,N_2454,N_2536);
xnor U2662 (N_2662,N_2418,N_2412);
nor U2663 (N_2663,N_2497,N_2507);
nand U2664 (N_2664,N_2495,N_2401);
or U2665 (N_2665,N_2517,N_2523);
nand U2666 (N_2666,N_2476,N_2538);
xor U2667 (N_2667,N_2419,N_2476);
xor U2668 (N_2668,N_2412,N_2402);
and U2669 (N_2669,N_2445,N_2519);
xor U2670 (N_2670,N_2530,N_2459);
nor U2671 (N_2671,N_2535,N_2463);
and U2672 (N_2672,N_2470,N_2422);
nor U2673 (N_2673,N_2533,N_2461);
nand U2674 (N_2674,N_2529,N_2526);
nand U2675 (N_2675,N_2541,N_2439);
xnor U2676 (N_2676,N_2435,N_2506);
and U2677 (N_2677,N_2467,N_2462);
nand U2678 (N_2678,N_2467,N_2532);
or U2679 (N_2679,N_2463,N_2510);
and U2680 (N_2680,N_2482,N_2452);
or U2681 (N_2681,N_2488,N_2412);
and U2682 (N_2682,N_2532,N_2457);
and U2683 (N_2683,N_2429,N_2421);
and U2684 (N_2684,N_2411,N_2479);
nor U2685 (N_2685,N_2460,N_2451);
xnor U2686 (N_2686,N_2407,N_2451);
xnor U2687 (N_2687,N_2543,N_2417);
nor U2688 (N_2688,N_2508,N_2450);
or U2689 (N_2689,N_2412,N_2541);
nand U2690 (N_2690,N_2463,N_2443);
nand U2691 (N_2691,N_2506,N_2534);
and U2692 (N_2692,N_2547,N_2480);
or U2693 (N_2693,N_2524,N_2486);
nor U2694 (N_2694,N_2414,N_2430);
and U2695 (N_2695,N_2404,N_2420);
xnor U2696 (N_2696,N_2460,N_2521);
or U2697 (N_2697,N_2500,N_2460);
nor U2698 (N_2698,N_2402,N_2512);
and U2699 (N_2699,N_2477,N_2472);
nor U2700 (N_2700,N_2553,N_2678);
xnor U2701 (N_2701,N_2659,N_2632);
xor U2702 (N_2702,N_2672,N_2627);
or U2703 (N_2703,N_2640,N_2697);
or U2704 (N_2704,N_2613,N_2677);
xnor U2705 (N_2705,N_2608,N_2555);
nand U2706 (N_2706,N_2664,N_2690);
xor U2707 (N_2707,N_2685,N_2581);
and U2708 (N_2708,N_2631,N_2605);
xor U2709 (N_2709,N_2626,N_2571);
nand U2710 (N_2710,N_2680,N_2556);
and U2711 (N_2711,N_2662,N_2559);
xnor U2712 (N_2712,N_2603,N_2578);
nor U2713 (N_2713,N_2569,N_2598);
xor U2714 (N_2714,N_2686,N_2649);
or U2715 (N_2715,N_2570,N_2574);
nor U2716 (N_2716,N_2643,N_2617);
or U2717 (N_2717,N_2592,N_2698);
and U2718 (N_2718,N_2667,N_2566);
nor U2719 (N_2719,N_2619,N_2567);
xor U2720 (N_2720,N_2562,N_2606);
nand U2721 (N_2721,N_2647,N_2657);
nor U2722 (N_2722,N_2642,N_2651);
or U2723 (N_2723,N_2628,N_2687);
nand U2724 (N_2724,N_2586,N_2563);
or U2725 (N_2725,N_2652,N_2577);
xnor U2726 (N_2726,N_2564,N_2573);
xnor U2727 (N_2727,N_2641,N_2621);
and U2728 (N_2728,N_2648,N_2602);
nand U2729 (N_2729,N_2666,N_2624);
and U2730 (N_2730,N_2575,N_2585);
xor U2731 (N_2731,N_2604,N_2671);
nand U2732 (N_2732,N_2669,N_2661);
and U2733 (N_2733,N_2681,N_2634);
and U2734 (N_2734,N_2695,N_2636);
xnor U2735 (N_2735,N_2607,N_2576);
and U2736 (N_2736,N_2616,N_2554);
nand U2737 (N_2737,N_2579,N_2588);
nor U2738 (N_2738,N_2637,N_2660);
or U2739 (N_2739,N_2670,N_2638);
nor U2740 (N_2740,N_2673,N_2623);
and U2741 (N_2741,N_2650,N_2552);
xnor U2742 (N_2742,N_2595,N_2609);
xnor U2743 (N_2743,N_2572,N_2699);
xnor U2744 (N_2744,N_2551,N_2593);
or U2745 (N_2745,N_2635,N_2646);
nand U2746 (N_2746,N_2618,N_2692);
and U2747 (N_2747,N_2600,N_2630);
xor U2748 (N_2748,N_2594,N_2684);
or U2749 (N_2749,N_2597,N_2633);
nor U2750 (N_2750,N_2612,N_2560);
or U2751 (N_2751,N_2656,N_2676);
and U2752 (N_2752,N_2550,N_2665);
and U2753 (N_2753,N_2653,N_2589);
xor U2754 (N_2754,N_2682,N_2584);
xnor U2755 (N_2755,N_2614,N_2558);
or U2756 (N_2756,N_2679,N_2561);
or U2757 (N_2757,N_2693,N_2645);
nor U2758 (N_2758,N_2622,N_2596);
and U2759 (N_2759,N_2611,N_2691);
nor U2760 (N_2760,N_2696,N_2683);
and U2761 (N_2761,N_2615,N_2668);
nor U2762 (N_2762,N_2689,N_2568);
nand U2763 (N_2763,N_2580,N_2625);
xnor U2764 (N_2764,N_2658,N_2582);
nor U2765 (N_2765,N_2610,N_2587);
xnor U2766 (N_2766,N_2557,N_2688);
nor U2767 (N_2767,N_2599,N_2620);
nand U2768 (N_2768,N_2674,N_2639);
nor U2769 (N_2769,N_2644,N_2601);
xor U2770 (N_2770,N_2583,N_2675);
xnor U2771 (N_2771,N_2654,N_2655);
or U2772 (N_2772,N_2663,N_2590);
or U2773 (N_2773,N_2565,N_2629);
nand U2774 (N_2774,N_2591,N_2694);
or U2775 (N_2775,N_2688,N_2654);
nor U2776 (N_2776,N_2671,N_2594);
xnor U2777 (N_2777,N_2648,N_2634);
xnor U2778 (N_2778,N_2638,N_2646);
and U2779 (N_2779,N_2605,N_2565);
nor U2780 (N_2780,N_2680,N_2655);
xor U2781 (N_2781,N_2627,N_2655);
xnor U2782 (N_2782,N_2692,N_2647);
and U2783 (N_2783,N_2687,N_2692);
nand U2784 (N_2784,N_2637,N_2686);
nor U2785 (N_2785,N_2691,N_2637);
and U2786 (N_2786,N_2664,N_2698);
and U2787 (N_2787,N_2594,N_2575);
or U2788 (N_2788,N_2581,N_2583);
nand U2789 (N_2789,N_2575,N_2612);
and U2790 (N_2790,N_2616,N_2597);
and U2791 (N_2791,N_2636,N_2673);
or U2792 (N_2792,N_2632,N_2647);
xor U2793 (N_2793,N_2653,N_2620);
nand U2794 (N_2794,N_2580,N_2587);
and U2795 (N_2795,N_2657,N_2658);
and U2796 (N_2796,N_2553,N_2686);
or U2797 (N_2797,N_2634,N_2642);
xnor U2798 (N_2798,N_2569,N_2561);
nor U2799 (N_2799,N_2644,N_2589);
or U2800 (N_2800,N_2611,N_2600);
nor U2801 (N_2801,N_2675,N_2623);
or U2802 (N_2802,N_2559,N_2624);
nor U2803 (N_2803,N_2687,N_2591);
and U2804 (N_2804,N_2698,N_2671);
and U2805 (N_2805,N_2645,N_2654);
nand U2806 (N_2806,N_2591,N_2665);
nor U2807 (N_2807,N_2564,N_2593);
nand U2808 (N_2808,N_2609,N_2658);
and U2809 (N_2809,N_2571,N_2644);
xnor U2810 (N_2810,N_2623,N_2630);
and U2811 (N_2811,N_2677,N_2572);
nor U2812 (N_2812,N_2649,N_2586);
or U2813 (N_2813,N_2607,N_2617);
xor U2814 (N_2814,N_2695,N_2647);
or U2815 (N_2815,N_2562,N_2633);
nand U2816 (N_2816,N_2690,N_2567);
and U2817 (N_2817,N_2609,N_2578);
nor U2818 (N_2818,N_2556,N_2560);
xor U2819 (N_2819,N_2609,N_2592);
nand U2820 (N_2820,N_2600,N_2590);
or U2821 (N_2821,N_2588,N_2673);
nand U2822 (N_2822,N_2637,N_2618);
nor U2823 (N_2823,N_2560,N_2624);
xor U2824 (N_2824,N_2684,N_2696);
nand U2825 (N_2825,N_2560,N_2607);
nand U2826 (N_2826,N_2672,N_2689);
nand U2827 (N_2827,N_2562,N_2622);
or U2828 (N_2828,N_2600,N_2574);
and U2829 (N_2829,N_2576,N_2582);
nand U2830 (N_2830,N_2567,N_2565);
and U2831 (N_2831,N_2615,N_2580);
xor U2832 (N_2832,N_2655,N_2568);
xor U2833 (N_2833,N_2698,N_2653);
nor U2834 (N_2834,N_2616,N_2557);
and U2835 (N_2835,N_2697,N_2617);
xnor U2836 (N_2836,N_2657,N_2612);
nor U2837 (N_2837,N_2636,N_2679);
xor U2838 (N_2838,N_2553,N_2654);
nor U2839 (N_2839,N_2622,N_2650);
or U2840 (N_2840,N_2590,N_2669);
nor U2841 (N_2841,N_2602,N_2632);
or U2842 (N_2842,N_2650,N_2697);
nor U2843 (N_2843,N_2584,N_2639);
xor U2844 (N_2844,N_2637,N_2638);
or U2845 (N_2845,N_2598,N_2597);
nor U2846 (N_2846,N_2687,N_2654);
and U2847 (N_2847,N_2583,N_2689);
or U2848 (N_2848,N_2576,N_2692);
nand U2849 (N_2849,N_2650,N_2671);
xnor U2850 (N_2850,N_2817,N_2847);
nand U2851 (N_2851,N_2738,N_2751);
and U2852 (N_2852,N_2794,N_2728);
xnor U2853 (N_2853,N_2819,N_2769);
nor U2854 (N_2854,N_2727,N_2792);
nand U2855 (N_2855,N_2789,N_2791);
or U2856 (N_2856,N_2757,N_2726);
nor U2857 (N_2857,N_2714,N_2783);
nor U2858 (N_2858,N_2836,N_2731);
and U2859 (N_2859,N_2716,N_2734);
nor U2860 (N_2860,N_2793,N_2702);
and U2861 (N_2861,N_2772,N_2780);
or U2862 (N_2862,N_2846,N_2710);
and U2863 (N_2863,N_2736,N_2740);
xnor U2864 (N_2864,N_2796,N_2730);
nand U2865 (N_2865,N_2745,N_2765);
nor U2866 (N_2866,N_2713,N_2760);
nand U2867 (N_2867,N_2763,N_2715);
and U2868 (N_2868,N_2759,N_2830);
nand U2869 (N_2869,N_2802,N_2808);
nor U2870 (N_2870,N_2803,N_2766);
nor U2871 (N_2871,N_2706,N_2776);
nor U2872 (N_2872,N_2835,N_2737);
nor U2873 (N_2873,N_2840,N_2735);
and U2874 (N_2874,N_2708,N_2767);
and U2875 (N_2875,N_2826,N_2827);
and U2876 (N_2876,N_2743,N_2717);
xor U2877 (N_2877,N_2774,N_2814);
xor U2878 (N_2878,N_2829,N_2704);
nor U2879 (N_2879,N_2754,N_2764);
xnor U2880 (N_2880,N_2805,N_2844);
nand U2881 (N_2881,N_2816,N_2810);
nand U2882 (N_2882,N_2739,N_2821);
or U2883 (N_2883,N_2747,N_2709);
nand U2884 (N_2884,N_2842,N_2721);
xnor U2885 (N_2885,N_2724,N_2822);
or U2886 (N_2886,N_2749,N_2823);
nand U2887 (N_2887,N_2839,N_2762);
nand U2888 (N_2888,N_2831,N_2752);
xnor U2889 (N_2889,N_2712,N_2729);
or U2890 (N_2890,N_2812,N_2801);
and U2891 (N_2891,N_2722,N_2742);
and U2892 (N_2892,N_2797,N_2787);
xor U2893 (N_2893,N_2790,N_2811);
nor U2894 (N_2894,N_2741,N_2786);
nor U2895 (N_2895,N_2804,N_2799);
and U2896 (N_2896,N_2725,N_2744);
and U2897 (N_2897,N_2723,N_2838);
and U2898 (N_2898,N_2746,N_2818);
nor U2899 (N_2899,N_2788,N_2711);
and U2900 (N_2900,N_2813,N_2732);
nand U2901 (N_2901,N_2837,N_2809);
and U2902 (N_2902,N_2784,N_2720);
nand U2903 (N_2903,N_2770,N_2705);
and U2904 (N_2904,N_2843,N_2785);
xor U2905 (N_2905,N_2781,N_2700);
and U2906 (N_2906,N_2771,N_2733);
or U2907 (N_2907,N_2777,N_2841);
or U2908 (N_2908,N_2806,N_2719);
and U2909 (N_2909,N_2701,N_2795);
nand U2910 (N_2910,N_2834,N_2820);
and U2911 (N_2911,N_2707,N_2748);
nand U2912 (N_2912,N_2778,N_2755);
and U2913 (N_2913,N_2825,N_2782);
nor U2914 (N_2914,N_2848,N_2833);
nand U2915 (N_2915,N_2824,N_2798);
nand U2916 (N_2916,N_2750,N_2768);
nor U2917 (N_2917,N_2807,N_2832);
xnor U2918 (N_2918,N_2718,N_2828);
and U2919 (N_2919,N_2703,N_2756);
or U2920 (N_2920,N_2775,N_2845);
or U2921 (N_2921,N_2761,N_2800);
nand U2922 (N_2922,N_2779,N_2815);
or U2923 (N_2923,N_2773,N_2753);
xor U2924 (N_2924,N_2849,N_2758);
nor U2925 (N_2925,N_2826,N_2819);
xor U2926 (N_2926,N_2848,N_2735);
nand U2927 (N_2927,N_2731,N_2752);
nand U2928 (N_2928,N_2737,N_2793);
xnor U2929 (N_2929,N_2814,N_2826);
or U2930 (N_2930,N_2765,N_2730);
and U2931 (N_2931,N_2723,N_2823);
nor U2932 (N_2932,N_2766,N_2707);
xnor U2933 (N_2933,N_2777,N_2816);
or U2934 (N_2934,N_2723,N_2785);
and U2935 (N_2935,N_2843,N_2771);
nand U2936 (N_2936,N_2751,N_2769);
or U2937 (N_2937,N_2765,N_2812);
xor U2938 (N_2938,N_2809,N_2807);
xnor U2939 (N_2939,N_2789,N_2765);
xor U2940 (N_2940,N_2805,N_2714);
and U2941 (N_2941,N_2700,N_2801);
nor U2942 (N_2942,N_2744,N_2843);
and U2943 (N_2943,N_2733,N_2759);
nor U2944 (N_2944,N_2712,N_2768);
xnor U2945 (N_2945,N_2773,N_2768);
or U2946 (N_2946,N_2796,N_2813);
nand U2947 (N_2947,N_2734,N_2846);
nor U2948 (N_2948,N_2767,N_2800);
or U2949 (N_2949,N_2807,N_2805);
xnor U2950 (N_2950,N_2711,N_2703);
xor U2951 (N_2951,N_2713,N_2740);
nand U2952 (N_2952,N_2739,N_2764);
or U2953 (N_2953,N_2770,N_2709);
or U2954 (N_2954,N_2766,N_2724);
and U2955 (N_2955,N_2821,N_2756);
or U2956 (N_2956,N_2812,N_2730);
nand U2957 (N_2957,N_2702,N_2838);
or U2958 (N_2958,N_2775,N_2735);
xnor U2959 (N_2959,N_2826,N_2840);
xor U2960 (N_2960,N_2729,N_2836);
nand U2961 (N_2961,N_2717,N_2733);
nand U2962 (N_2962,N_2749,N_2812);
nand U2963 (N_2963,N_2721,N_2755);
nor U2964 (N_2964,N_2798,N_2806);
and U2965 (N_2965,N_2801,N_2765);
or U2966 (N_2966,N_2786,N_2736);
xor U2967 (N_2967,N_2846,N_2840);
or U2968 (N_2968,N_2813,N_2797);
nor U2969 (N_2969,N_2805,N_2701);
xor U2970 (N_2970,N_2791,N_2823);
nand U2971 (N_2971,N_2744,N_2833);
nand U2972 (N_2972,N_2754,N_2842);
nor U2973 (N_2973,N_2731,N_2751);
nor U2974 (N_2974,N_2726,N_2805);
and U2975 (N_2975,N_2837,N_2797);
nor U2976 (N_2976,N_2757,N_2720);
xor U2977 (N_2977,N_2830,N_2766);
xnor U2978 (N_2978,N_2775,N_2802);
or U2979 (N_2979,N_2817,N_2702);
or U2980 (N_2980,N_2701,N_2808);
or U2981 (N_2981,N_2845,N_2784);
and U2982 (N_2982,N_2779,N_2795);
or U2983 (N_2983,N_2815,N_2795);
nand U2984 (N_2984,N_2729,N_2707);
nor U2985 (N_2985,N_2805,N_2826);
xor U2986 (N_2986,N_2749,N_2796);
and U2987 (N_2987,N_2847,N_2764);
and U2988 (N_2988,N_2764,N_2782);
nand U2989 (N_2989,N_2757,N_2774);
or U2990 (N_2990,N_2707,N_2827);
xnor U2991 (N_2991,N_2729,N_2805);
nor U2992 (N_2992,N_2747,N_2806);
and U2993 (N_2993,N_2731,N_2847);
or U2994 (N_2994,N_2741,N_2754);
and U2995 (N_2995,N_2701,N_2824);
or U2996 (N_2996,N_2707,N_2747);
and U2997 (N_2997,N_2745,N_2735);
nor U2998 (N_2998,N_2730,N_2795);
xor U2999 (N_2999,N_2712,N_2802);
nor U3000 (N_3000,N_2994,N_2934);
xor U3001 (N_3001,N_2879,N_2997);
nand U3002 (N_3002,N_2872,N_2925);
nand U3003 (N_3003,N_2853,N_2896);
or U3004 (N_3004,N_2892,N_2967);
xnor U3005 (N_3005,N_2954,N_2919);
nor U3006 (N_3006,N_2970,N_2977);
nor U3007 (N_3007,N_2902,N_2928);
nor U3008 (N_3008,N_2991,N_2929);
nor U3009 (N_3009,N_2877,N_2944);
nor U3010 (N_3010,N_2863,N_2965);
and U3011 (N_3011,N_2867,N_2958);
or U3012 (N_3012,N_2886,N_2936);
and U3013 (N_3013,N_2924,N_2948);
nand U3014 (N_3014,N_2889,N_2938);
and U3015 (N_3015,N_2895,N_2899);
xnor U3016 (N_3016,N_2971,N_2881);
nand U3017 (N_3017,N_2975,N_2859);
xor U3018 (N_3018,N_2874,N_2916);
and U3019 (N_3019,N_2900,N_2966);
nor U3020 (N_3020,N_2921,N_2969);
nand U3021 (N_3021,N_2890,N_2964);
or U3022 (N_3022,N_2945,N_2998);
nor U3023 (N_3023,N_2993,N_2891);
nand U3024 (N_3024,N_2876,N_2856);
nand U3025 (N_3025,N_2927,N_2862);
and U3026 (N_3026,N_2888,N_2941);
nor U3027 (N_3027,N_2939,N_2915);
xnor U3028 (N_3028,N_2855,N_2946);
and U3029 (N_3029,N_2981,N_2984);
and U3030 (N_3030,N_2972,N_2996);
nand U3031 (N_3031,N_2901,N_2850);
nand U3032 (N_3032,N_2912,N_2926);
and U3033 (N_3033,N_2858,N_2875);
or U3034 (N_3034,N_2983,N_2871);
and U3035 (N_3035,N_2884,N_2987);
and U3036 (N_3036,N_2990,N_2956);
nand U3037 (N_3037,N_2905,N_2898);
xor U3038 (N_3038,N_2992,N_2878);
nor U3039 (N_3039,N_2957,N_2914);
nand U3040 (N_3040,N_2962,N_2961);
nand U3041 (N_3041,N_2932,N_2897);
and U3042 (N_3042,N_2870,N_2873);
and U3043 (N_3043,N_2950,N_2989);
nor U3044 (N_3044,N_2885,N_2860);
nand U3045 (N_3045,N_2923,N_2974);
xor U3046 (N_3046,N_2880,N_2882);
nor U3047 (N_3047,N_2930,N_2988);
or U3048 (N_3048,N_2922,N_2952);
xor U3049 (N_3049,N_2973,N_2887);
nand U3050 (N_3050,N_2913,N_2866);
or U3051 (N_3051,N_2947,N_2986);
nor U3052 (N_3052,N_2869,N_2953);
nor U3053 (N_3053,N_2851,N_2852);
or U3054 (N_3054,N_2864,N_2995);
nand U3055 (N_3055,N_2976,N_2985);
and U3056 (N_3056,N_2854,N_2968);
and U3057 (N_3057,N_2865,N_2907);
nor U3058 (N_3058,N_2933,N_2918);
xor U3059 (N_3059,N_2903,N_2980);
or U3060 (N_3060,N_2949,N_2979);
nand U3061 (N_3061,N_2959,N_2935);
nand U3062 (N_3062,N_2951,N_2917);
or U3063 (N_3063,N_2894,N_2920);
nor U3064 (N_3064,N_2883,N_2893);
or U3065 (N_3065,N_2937,N_2904);
and U3066 (N_3066,N_2906,N_2910);
xnor U3067 (N_3067,N_2943,N_2963);
xor U3068 (N_3068,N_2868,N_2908);
nor U3069 (N_3069,N_2861,N_2942);
xor U3070 (N_3070,N_2940,N_2955);
xor U3071 (N_3071,N_2978,N_2999);
nor U3072 (N_3072,N_2911,N_2909);
or U3073 (N_3073,N_2857,N_2982);
or U3074 (N_3074,N_2931,N_2960);
and U3075 (N_3075,N_2982,N_2920);
and U3076 (N_3076,N_2898,N_2858);
and U3077 (N_3077,N_2902,N_2957);
nor U3078 (N_3078,N_2898,N_2984);
xor U3079 (N_3079,N_2852,N_2963);
xnor U3080 (N_3080,N_2852,N_2903);
or U3081 (N_3081,N_2991,N_2990);
nand U3082 (N_3082,N_2959,N_2941);
nor U3083 (N_3083,N_2904,N_2982);
xor U3084 (N_3084,N_2950,N_2943);
nand U3085 (N_3085,N_2892,N_2982);
xor U3086 (N_3086,N_2932,N_2906);
and U3087 (N_3087,N_2953,N_2936);
nor U3088 (N_3088,N_2913,N_2881);
nand U3089 (N_3089,N_2956,N_2959);
xor U3090 (N_3090,N_2864,N_2877);
nand U3091 (N_3091,N_2958,N_2991);
xor U3092 (N_3092,N_2969,N_2891);
and U3093 (N_3093,N_2936,N_2944);
nand U3094 (N_3094,N_2981,N_2988);
nand U3095 (N_3095,N_2943,N_2866);
and U3096 (N_3096,N_2927,N_2899);
and U3097 (N_3097,N_2962,N_2946);
nand U3098 (N_3098,N_2933,N_2903);
and U3099 (N_3099,N_2905,N_2908);
nor U3100 (N_3100,N_2866,N_2947);
xor U3101 (N_3101,N_2867,N_2928);
or U3102 (N_3102,N_2920,N_2915);
or U3103 (N_3103,N_2923,N_2991);
xnor U3104 (N_3104,N_2890,N_2973);
xor U3105 (N_3105,N_2868,N_2986);
and U3106 (N_3106,N_2967,N_2984);
and U3107 (N_3107,N_2890,N_2858);
nor U3108 (N_3108,N_2964,N_2982);
and U3109 (N_3109,N_2852,N_2910);
or U3110 (N_3110,N_2991,N_2950);
or U3111 (N_3111,N_2920,N_2964);
nand U3112 (N_3112,N_2888,N_2996);
nand U3113 (N_3113,N_2949,N_2908);
xnor U3114 (N_3114,N_2868,N_2944);
nand U3115 (N_3115,N_2960,N_2965);
xnor U3116 (N_3116,N_2975,N_2860);
xnor U3117 (N_3117,N_2858,N_2990);
nand U3118 (N_3118,N_2990,N_2873);
or U3119 (N_3119,N_2984,N_2885);
nor U3120 (N_3120,N_2925,N_2993);
nor U3121 (N_3121,N_2970,N_2859);
and U3122 (N_3122,N_2930,N_2853);
xor U3123 (N_3123,N_2902,N_2960);
xnor U3124 (N_3124,N_2875,N_2949);
nand U3125 (N_3125,N_2935,N_2869);
nor U3126 (N_3126,N_2976,N_2938);
and U3127 (N_3127,N_2892,N_2865);
nand U3128 (N_3128,N_2891,N_2927);
or U3129 (N_3129,N_2907,N_2989);
nand U3130 (N_3130,N_2875,N_2925);
xnor U3131 (N_3131,N_2986,N_2906);
or U3132 (N_3132,N_2969,N_2905);
or U3133 (N_3133,N_2857,N_2906);
nor U3134 (N_3134,N_2885,N_2886);
or U3135 (N_3135,N_2893,N_2882);
nor U3136 (N_3136,N_2924,N_2936);
nand U3137 (N_3137,N_2868,N_2869);
and U3138 (N_3138,N_2899,N_2891);
nand U3139 (N_3139,N_2951,N_2935);
or U3140 (N_3140,N_2949,N_2921);
xnor U3141 (N_3141,N_2979,N_2878);
nand U3142 (N_3142,N_2882,N_2889);
xor U3143 (N_3143,N_2937,N_2893);
and U3144 (N_3144,N_2958,N_2976);
xnor U3145 (N_3145,N_2974,N_2866);
xor U3146 (N_3146,N_2939,N_2965);
nand U3147 (N_3147,N_2972,N_2855);
and U3148 (N_3148,N_2929,N_2859);
and U3149 (N_3149,N_2976,N_2921);
or U3150 (N_3150,N_3031,N_3139);
and U3151 (N_3151,N_3034,N_3077);
nand U3152 (N_3152,N_3132,N_3125);
nand U3153 (N_3153,N_3094,N_3016);
or U3154 (N_3154,N_3030,N_3044);
nor U3155 (N_3155,N_3146,N_3058);
nor U3156 (N_3156,N_3110,N_3046);
or U3157 (N_3157,N_3023,N_3112);
nand U3158 (N_3158,N_3056,N_3127);
and U3159 (N_3159,N_3064,N_3007);
nand U3160 (N_3160,N_3065,N_3089);
nand U3161 (N_3161,N_3107,N_3081);
nand U3162 (N_3162,N_3018,N_3109);
xor U3163 (N_3163,N_3048,N_3050);
and U3164 (N_3164,N_3093,N_3011);
or U3165 (N_3165,N_3036,N_3037);
nand U3166 (N_3166,N_3114,N_3099);
nand U3167 (N_3167,N_3005,N_3010);
xor U3168 (N_3168,N_3137,N_3003);
nand U3169 (N_3169,N_3095,N_3144);
nor U3170 (N_3170,N_3013,N_3052);
or U3171 (N_3171,N_3025,N_3135);
or U3172 (N_3172,N_3067,N_3113);
nand U3173 (N_3173,N_3138,N_3103);
xnor U3174 (N_3174,N_3128,N_3075);
or U3175 (N_3175,N_3062,N_3142);
nor U3176 (N_3176,N_3119,N_3100);
xor U3177 (N_3177,N_3053,N_3105);
xor U3178 (N_3178,N_3121,N_3085);
nor U3179 (N_3179,N_3140,N_3038);
or U3180 (N_3180,N_3117,N_3054);
nor U3181 (N_3181,N_3017,N_3019);
nor U3182 (N_3182,N_3123,N_3091);
or U3183 (N_3183,N_3145,N_3028);
nor U3184 (N_3184,N_3066,N_3111);
xor U3185 (N_3185,N_3082,N_3001);
nor U3186 (N_3186,N_3087,N_3027);
or U3187 (N_3187,N_3042,N_3047);
xor U3188 (N_3188,N_3035,N_3043);
nand U3189 (N_3189,N_3120,N_3014);
xor U3190 (N_3190,N_3129,N_3057);
or U3191 (N_3191,N_3026,N_3051);
xnor U3192 (N_3192,N_3088,N_3080);
nor U3193 (N_3193,N_3074,N_3122);
or U3194 (N_3194,N_3096,N_3072);
or U3195 (N_3195,N_3124,N_3148);
or U3196 (N_3196,N_3006,N_3101);
nor U3197 (N_3197,N_3055,N_3020);
nand U3198 (N_3198,N_3008,N_3032);
nor U3199 (N_3199,N_3069,N_3083);
nand U3200 (N_3200,N_3149,N_3092);
nand U3201 (N_3201,N_3104,N_3049);
xnor U3202 (N_3202,N_3108,N_3136);
xnor U3203 (N_3203,N_3024,N_3076);
nand U3204 (N_3204,N_3033,N_3141);
nor U3205 (N_3205,N_3002,N_3116);
nand U3206 (N_3206,N_3063,N_3086);
nand U3207 (N_3207,N_3012,N_3084);
or U3208 (N_3208,N_3130,N_3073);
and U3209 (N_3209,N_3115,N_3045);
nor U3210 (N_3210,N_3068,N_3078);
or U3211 (N_3211,N_3070,N_3060);
and U3212 (N_3212,N_3097,N_3015);
nand U3213 (N_3213,N_3131,N_3143);
xnor U3214 (N_3214,N_3059,N_3004);
or U3215 (N_3215,N_3090,N_3133);
or U3216 (N_3216,N_3021,N_3009);
or U3217 (N_3217,N_3079,N_3098);
xor U3218 (N_3218,N_3039,N_3041);
nor U3219 (N_3219,N_3022,N_3134);
xor U3220 (N_3220,N_3126,N_3071);
nand U3221 (N_3221,N_3029,N_3118);
xor U3222 (N_3222,N_3040,N_3102);
nor U3223 (N_3223,N_3061,N_3106);
xnor U3224 (N_3224,N_3147,N_3000);
nand U3225 (N_3225,N_3073,N_3040);
nand U3226 (N_3226,N_3045,N_3089);
nor U3227 (N_3227,N_3024,N_3035);
and U3228 (N_3228,N_3084,N_3015);
nor U3229 (N_3229,N_3073,N_3006);
xor U3230 (N_3230,N_3123,N_3079);
xor U3231 (N_3231,N_3093,N_3136);
or U3232 (N_3232,N_3014,N_3033);
or U3233 (N_3233,N_3084,N_3008);
xnor U3234 (N_3234,N_3137,N_3045);
xor U3235 (N_3235,N_3041,N_3089);
nor U3236 (N_3236,N_3133,N_3070);
xor U3237 (N_3237,N_3014,N_3028);
nand U3238 (N_3238,N_3001,N_3112);
nor U3239 (N_3239,N_3041,N_3124);
nor U3240 (N_3240,N_3062,N_3010);
or U3241 (N_3241,N_3030,N_3022);
or U3242 (N_3242,N_3033,N_3099);
xor U3243 (N_3243,N_3042,N_3083);
or U3244 (N_3244,N_3061,N_3025);
xor U3245 (N_3245,N_3141,N_3066);
nor U3246 (N_3246,N_3069,N_3147);
or U3247 (N_3247,N_3109,N_3110);
nand U3248 (N_3248,N_3104,N_3130);
nor U3249 (N_3249,N_3063,N_3011);
nand U3250 (N_3250,N_3060,N_3124);
nor U3251 (N_3251,N_3040,N_3034);
xor U3252 (N_3252,N_3080,N_3134);
xnor U3253 (N_3253,N_3125,N_3016);
xnor U3254 (N_3254,N_3096,N_3078);
nor U3255 (N_3255,N_3110,N_3087);
xnor U3256 (N_3256,N_3025,N_3085);
nor U3257 (N_3257,N_3096,N_3095);
nand U3258 (N_3258,N_3079,N_3127);
xnor U3259 (N_3259,N_3106,N_3054);
and U3260 (N_3260,N_3120,N_3146);
xnor U3261 (N_3261,N_3098,N_3021);
xnor U3262 (N_3262,N_3100,N_3114);
or U3263 (N_3263,N_3124,N_3076);
or U3264 (N_3264,N_3132,N_3053);
and U3265 (N_3265,N_3054,N_3015);
xnor U3266 (N_3266,N_3088,N_3037);
xnor U3267 (N_3267,N_3061,N_3129);
xnor U3268 (N_3268,N_3136,N_3035);
nand U3269 (N_3269,N_3014,N_3039);
xor U3270 (N_3270,N_3034,N_3063);
xnor U3271 (N_3271,N_3108,N_3089);
nor U3272 (N_3272,N_3014,N_3040);
and U3273 (N_3273,N_3087,N_3148);
xnor U3274 (N_3274,N_3070,N_3033);
nand U3275 (N_3275,N_3108,N_3039);
nand U3276 (N_3276,N_3036,N_3050);
or U3277 (N_3277,N_3037,N_3120);
nor U3278 (N_3278,N_3106,N_3062);
nand U3279 (N_3279,N_3032,N_3135);
nor U3280 (N_3280,N_3116,N_3080);
xnor U3281 (N_3281,N_3137,N_3076);
and U3282 (N_3282,N_3067,N_3083);
or U3283 (N_3283,N_3149,N_3032);
and U3284 (N_3284,N_3053,N_3038);
nor U3285 (N_3285,N_3119,N_3078);
and U3286 (N_3286,N_3036,N_3065);
nor U3287 (N_3287,N_3120,N_3054);
and U3288 (N_3288,N_3098,N_3071);
and U3289 (N_3289,N_3015,N_3094);
nand U3290 (N_3290,N_3107,N_3019);
xnor U3291 (N_3291,N_3026,N_3066);
and U3292 (N_3292,N_3115,N_3141);
and U3293 (N_3293,N_3138,N_3076);
and U3294 (N_3294,N_3083,N_3036);
nand U3295 (N_3295,N_3005,N_3130);
nand U3296 (N_3296,N_3078,N_3100);
xnor U3297 (N_3297,N_3012,N_3080);
xnor U3298 (N_3298,N_3072,N_3051);
nand U3299 (N_3299,N_3076,N_3001);
and U3300 (N_3300,N_3289,N_3184);
nand U3301 (N_3301,N_3281,N_3228);
nor U3302 (N_3302,N_3178,N_3210);
nand U3303 (N_3303,N_3267,N_3262);
or U3304 (N_3304,N_3251,N_3249);
xnor U3305 (N_3305,N_3179,N_3218);
or U3306 (N_3306,N_3271,N_3230);
nand U3307 (N_3307,N_3292,N_3260);
and U3308 (N_3308,N_3155,N_3158);
nand U3309 (N_3309,N_3270,N_3227);
or U3310 (N_3310,N_3219,N_3159);
and U3311 (N_3311,N_3295,N_3252);
nand U3312 (N_3312,N_3239,N_3176);
xor U3313 (N_3313,N_3182,N_3231);
nand U3314 (N_3314,N_3265,N_3293);
xor U3315 (N_3315,N_3211,N_3296);
nand U3316 (N_3316,N_3183,N_3291);
xor U3317 (N_3317,N_3257,N_3152);
or U3318 (N_3318,N_3197,N_3163);
nand U3319 (N_3319,N_3151,N_3215);
xnor U3320 (N_3320,N_3234,N_3288);
and U3321 (N_3321,N_3186,N_3187);
nor U3322 (N_3322,N_3254,N_3172);
nand U3323 (N_3323,N_3225,N_3194);
xnor U3324 (N_3324,N_3195,N_3277);
or U3325 (N_3325,N_3216,N_3212);
and U3326 (N_3326,N_3196,N_3226);
xor U3327 (N_3327,N_3282,N_3276);
nand U3328 (N_3328,N_3258,N_3250);
xnor U3329 (N_3329,N_3253,N_3246);
nor U3330 (N_3330,N_3229,N_3190);
nor U3331 (N_3331,N_3272,N_3294);
xnor U3332 (N_3332,N_3165,N_3221);
or U3333 (N_3333,N_3247,N_3205);
and U3334 (N_3334,N_3177,N_3213);
or U3335 (N_3335,N_3298,N_3264);
nand U3336 (N_3336,N_3169,N_3191);
and U3337 (N_3337,N_3168,N_3201);
nand U3338 (N_3338,N_3171,N_3185);
xnor U3339 (N_3339,N_3266,N_3297);
nand U3340 (N_3340,N_3198,N_3233);
nor U3341 (N_3341,N_3263,N_3156);
or U3342 (N_3342,N_3160,N_3285);
or U3343 (N_3343,N_3268,N_3173);
nand U3344 (N_3344,N_3244,N_3243);
nor U3345 (N_3345,N_3248,N_3274);
or U3346 (N_3346,N_3188,N_3245);
nand U3347 (N_3347,N_3214,N_3299);
nand U3348 (N_3348,N_3162,N_3208);
and U3349 (N_3349,N_3259,N_3154);
and U3350 (N_3350,N_3181,N_3157);
and U3351 (N_3351,N_3206,N_3237);
xnor U3352 (N_3352,N_3153,N_3164);
xnor U3353 (N_3353,N_3280,N_3207);
nor U3354 (N_3354,N_3242,N_3286);
nand U3355 (N_3355,N_3261,N_3199);
and U3356 (N_3356,N_3232,N_3193);
nor U3357 (N_3357,N_3290,N_3223);
or U3358 (N_3358,N_3241,N_3174);
xor U3359 (N_3359,N_3287,N_3273);
and U3360 (N_3360,N_3203,N_3202);
and U3361 (N_3361,N_3170,N_3200);
or U3362 (N_3362,N_3180,N_3192);
and U3363 (N_3363,N_3150,N_3204);
xnor U3364 (N_3364,N_3217,N_3240);
and U3365 (N_3365,N_3283,N_3275);
nor U3366 (N_3366,N_3255,N_3175);
xnor U3367 (N_3367,N_3279,N_3284);
and U3368 (N_3368,N_3189,N_3209);
nand U3369 (N_3369,N_3235,N_3167);
nor U3370 (N_3370,N_3220,N_3224);
and U3371 (N_3371,N_3269,N_3161);
and U3372 (N_3372,N_3278,N_3222);
xor U3373 (N_3373,N_3236,N_3166);
and U3374 (N_3374,N_3238,N_3256);
and U3375 (N_3375,N_3211,N_3279);
nand U3376 (N_3376,N_3291,N_3292);
and U3377 (N_3377,N_3172,N_3236);
xor U3378 (N_3378,N_3260,N_3226);
nand U3379 (N_3379,N_3243,N_3161);
nand U3380 (N_3380,N_3282,N_3292);
nor U3381 (N_3381,N_3209,N_3150);
or U3382 (N_3382,N_3161,N_3240);
and U3383 (N_3383,N_3231,N_3183);
nand U3384 (N_3384,N_3294,N_3203);
or U3385 (N_3385,N_3210,N_3205);
or U3386 (N_3386,N_3254,N_3222);
nor U3387 (N_3387,N_3206,N_3191);
and U3388 (N_3388,N_3161,N_3185);
xor U3389 (N_3389,N_3179,N_3213);
or U3390 (N_3390,N_3297,N_3239);
nor U3391 (N_3391,N_3228,N_3159);
and U3392 (N_3392,N_3247,N_3233);
and U3393 (N_3393,N_3268,N_3186);
or U3394 (N_3394,N_3260,N_3234);
xor U3395 (N_3395,N_3237,N_3253);
or U3396 (N_3396,N_3289,N_3186);
nor U3397 (N_3397,N_3152,N_3286);
and U3398 (N_3398,N_3177,N_3188);
or U3399 (N_3399,N_3265,N_3152);
nor U3400 (N_3400,N_3159,N_3162);
and U3401 (N_3401,N_3291,N_3219);
and U3402 (N_3402,N_3286,N_3288);
or U3403 (N_3403,N_3293,N_3157);
or U3404 (N_3404,N_3193,N_3163);
nor U3405 (N_3405,N_3199,N_3251);
nor U3406 (N_3406,N_3240,N_3271);
xnor U3407 (N_3407,N_3165,N_3181);
nand U3408 (N_3408,N_3284,N_3246);
nand U3409 (N_3409,N_3185,N_3297);
nor U3410 (N_3410,N_3298,N_3217);
and U3411 (N_3411,N_3293,N_3296);
nor U3412 (N_3412,N_3185,N_3290);
or U3413 (N_3413,N_3289,N_3294);
nand U3414 (N_3414,N_3215,N_3248);
and U3415 (N_3415,N_3272,N_3155);
xor U3416 (N_3416,N_3268,N_3225);
xor U3417 (N_3417,N_3223,N_3273);
nand U3418 (N_3418,N_3211,N_3268);
xor U3419 (N_3419,N_3292,N_3156);
or U3420 (N_3420,N_3159,N_3262);
and U3421 (N_3421,N_3172,N_3297);
nand U3422 (N_3422,N_3216,N_3258);
nand U3423 (N_3423,N_3198,N_3159);
or U3424 (N_3424,N_3179,N_3188);
nor U3425 (N_3425,N_3243,N_3295);
nand U3426 (N_3426,N_3234,N_3198);
xnor U3427 (N_3427,N_3153,N_3183);
or U3428 (N_3428,N_3264,N_3283);
xor U3429 (N_3429,N_3160,N_3184);
nor U3430 (N_3430,N_3170,N_3239);
or U3431 (N_3431,N_3200,N_3292);
or U3432 (N_3432,N_3170,N_3222);
nand U3433 (N_3433,N_3151,N_3240);
xnor U3434 (N_3434,N_3249,N_3229);
nor U3435 (N_3435,N_3289,N_3163);
nand U3436 (N_3436,N_3176,N_3159);
xnor U3437 (N_3437,N_3178,N_3258);
and U3438 (N_3438,N_3250,N_3278);
and U3439 (N_3439,N_3274,N_3216);
nand U3440 (N_3440,N_3226,N_3291);
nand U3441 (N_3441,N_3262,N_3226);
nor U3442 (N_3442,N_3156,N_3194);
and U3443 (N_3443,N_3291,N_3166);
and U3444 (N_3444,N_3297,N_3291);
nand U3445 (N_3445,N_3205,N_3183);
xor U3446 (N_3446,N_3288,N_3202);
nor U3447 (N_3447,N_3274,N_3176);
or U3448 (N_3448,N_3183,N_3181);
nand U3449 (N_3449,N_3254,N_3189);
xor U3450 (N_3450,N_3320,N_3389);
and U3451 (N_3451,N_3380,N_3424);
or U3452 (N_3452,N_3316,N_3314);
and U3453 (N_3453,N_3415,N_3348);
nor U3454 (N_3454,N_3397,N_3334);
or U3455 (N_3455,N_3436,N_3443);
xnor U3456 (N_3456,N_3373,N_3434);
nor U3457 (N_3457,N_3416,N_3431);
nor U3458 (N_3458,N_3439,N_3386);
or U3459 (N_3459,N_3438,N_3430);
xor U3460 (N_3460,N_3336,N_3404);
xnor U3461 (N_3461,N_3433,N_3372);
or U3462 (N_3462,N_3427,N_3331);
nor U3463 (N_3463,N_3423,N_3370);
and U3464 (N_3464,N_3399,N_3401);
nor U3465 (N_3465,N_3357,N_3375);
nand U3466 (N_3466,N_3335,N_3325);
nand U3467 (N_3467,N_3418,N_3428);
or U3468 (N_3468,N_3302,N_3382);
and U3469 (N_3469,N_3394,N_3315);
and U3470 (N_3470,N_3351,N_3421);
nor U3471 (N_3471,N_3417,N_3413);
xor U3472 (N_3472,N_3381,N_3337);
nor U3473 (N_3473,N_3391,N_3383);
xor U3474 (N_3474,N_3303,N_3447);
or U3475 (N_3475,N_3445,N_3366);
and U3476 (N_3476,N_3308,N_3354);
nand U3477 (N_3477,N_3365,N_3441);
and U3478 (N_3478,N_3328,N_3367);
nand U3479 (N_3479,N_3322,N_3444);
xor U3480 (N_3480,N_3307,N_3306);
xnor U3481 (N_3481,N_3449,N_3400);
xor U3482 (N_3482,N_3368,N_3345);
nand U3483 (N_3483,N_3333,N_3311);
nand U3484 (N_3484,N_3414,N_3429);
xnor U3485 (N_3485,N_3412,N_3378);
nand U3486 (N_3486,N_3339,N_3317);
nand U3487 (N_3487,N_3385,N_3327);
nand U3488 (N_3488,N_3309,N_3338);
xnor U3489 (N_3489,N_3446,N_3324);
nor U3490 (N_3490,N_3405,N_3390);
nand U3491 (N_3491,N_3364,N_3369);
or U3492 (N_3492,N_3353,N_3321);
nor U3493 (N_3493,N_3358,N_3371);
nand U3494 (N_3494,N_3410,N_3326);
xor U3495 (N_3495,N_3305,N_3355);
xnor U3496 (N_3496,N_3300,N_3312);
xor U3497 (N_3497,N_3323,N_3313);
nor U3498 (N_3498,N_3376,N_3420);
and U3499 (N_3499,N_3425,N_3332);
or U3500 (N_3500,N_3406,N_3356);
or U3501 (N_3501,N_3422,N_3432);
nor U3502 (N_3502,N_3435,N_3442);
nor U3503 (N_3503,N_3395,N_3346);
or U3504 (N_3504,N_3361,N_3437);
nor U3505 (N_3505,N_3409,N_3304);
and U3506 (N_3506,N_3318,N_3388);
xnor U3507 (N_3507,N_3329,N_3377);
xor U3508 (N_3508,N_3374,N_3350);
xnor U3509 (N_3509,N_3408,N_3363);
nand U3510 (N_3510,N_3384,N_3393);
or U3511 (N_3511,N_3426,N_3392);
nor U3512 (N_3512,N_3360,N_3379);
xnor U3513 (N_3513,N_3407,N_3349);
and U3514 (N_3514,N_3341,N_3387);
and U3515 (N_3515,N_3319,N_3440);
nand U3516 (N_3516,N_3396,N_3359);
and U3517 (N_3517,N_3330,N_3352);
xnor U3518 (N_3518,N_3347,N_3419);
nor U3519 (N_3519,N_3402,N_3362);
xor U3520 (N_3520,N_3344,N_3403);
nor U3521 (N_3521,N_3310,N_3398);
nand U3522 (N_3522,N_3411,N_3342);
xor U3523 (N_3523,N_3343,N_3340);
and U3524 (N_3524,N_3448,N_3301);
nor U3525 (N_3525,N_3448,N_3325);
or U3526 (N_3526,N_3421,N_3376);
or U3527 (N_3527,N_3325,N_3366);
and U3528 (N_3528,N_3425,N_3366);
nand U3529 (N_3529,N_3419,N_3422);
nand U3530 (N_3530,N_3381,N_3389);
nand U3531 (N_3531,N_3360,N_3412);
nor U3532 (N_3532,N_3372,N_3366);
or U3533 (N_3533,N_3391,N_3343);
or U3534 (N_3534,N_3304,N_3337);
and U3535 (N_3535,N_3421,N_3377);
and U3536 (N_3536,N_3381,N_3351);
xnor U3537 (N_3537,N_3374,N_3333);
nor U3538 (N_3538,N_3430,N_3304);
nand U3539 (N_3539,N_3316,N_3337);
xnor U3540 (N_3540,N_3431,N_3438);
or U3541 (N_3541,N_3316,N_3365);
and U3542 (N_3542,N_3424,N_3345);
or U3543 (N_3543,N_3445,N_3412);
nor U3544 (N_3544,N_3428,N_3411);
or U3545 (N_3545,N_3391,N_3420);
and U3546 (N_3546,N_3405,N_3361);
and U3547 (N_3547,N_3423,N_3389);
xor U3548 (N_3548,N_3400,N_3310);
nand U3549 (N_3549,N_3302,N_3329);
xor U3550 (N_3550,N_3435,N_3431);
or U3551 (N_3551,N_3416,N_3445);
and U3552 (N_3552,N_3325,N_3361);
nor U3553 (N_3553,N_3403,N_3320);
nand U3554 (N_3554,N_3421,N_3325);
xnor U3555 (N_3555,N_3306,N_3319);
xnor U3556 (N_3556,N_3314,N_3442);
xor U3557 (N_3557,N_3436,N_3347);
or U3558 (N_3558,N_3324,N_3411);
nand U3559 (N_3559,N_3306,N_3311);
and U3560 (N_3560,N_3368,N_3379);
nand U3561 (N_3561,N_3309,N_3370);
and U3562 (N_3562,N_3404,N_3348);
xnor U3563 (N_3563,N_3449,N_3338);
xor U3564 (N_3564,N_3301,N_3310);
xnor U3565 (N_3565,N_3418,N_3386);
nor U3566 (N_3566,N_3410,N_3336);
nand U3567 (N_3567,N_3396,N_3386);
xor U3568 (N_3568,N_3353,N_3396);
or U3569 (N_3569,N_3430,N_3410);
and U3570 (N_3570,N_3347,N_3348);
or U3571 (N_3571,N_3405,N_3324);
nand U3572 (N_3572,N_3315,N_3321);
nor U3573 (N_3573,N_3314,N_3327);
nand U3574 (N_3574,N_3442,N_3329);
nor U3575 (N_3575,N_3413,N_3332);
and U3576 (N_3576,N_3414,N_3336);
nor U3577 (N_3577,N_3361,N_3417);
and U3578 (N_3578,N_3358,N_3412);
xnor U3579 (N_3579,N_3368,N_3363);
nor U3580 (N_3580,N_3358,N_3390);
nor U3581 (N_3581,N_3301,N_3303);
xor U3582 (N_3582,N_3355,N_3430);
xor U3583 (N_3583,N_3441,N_3443);
xor U3584 (N_3584,N_3317,N_3329);
xnor U3585 (N_3585,N_3355,N_3359);
and U3586 (N_3586,N_3343,N_3339);
nand U3587 (N_3587,N_3390,N_3395);
or U3588 (N_3588,N_3322,N_3378);
and U3589 (N_3589,N_3360,N_3340);
and U3590 (N_3590,N_3320,N_3324);
nor U3591 (N_3591,N_3321,N_3426);
and U3592 (N_3592,N_3327,N_3412);
xor U3593 (N_3593,N_3380,N_3322);
and U3594 (N_3594,N_3330,N_3360);
or U3595 (N_3595,N_3398,N_3408);
and U3596 (N_3596,N_3408,N_3443);
nand U3597 (N_3597,N_3337,N_3398);
nor U3598 (N_3598,N_3356,N_3305);
xor U3599 (N_3599,N_3352,N_3368);
xor U3600 (N_3600,N_3494,N_3574);
and U3601 (N_3601,N_3502,N_3516);
or U3602 (N_3602,N_3528,N_3543);
or U3603 (N_3603,N_3546,N_3522);
xor U3604 (N_3604,N_3515,N_3460);
or U3605 (N_3605,N_3592,N_3525);
or U3606 (N_3606,N_3567,N_3454);
or U3607 (N_3607,N_3492,N_3468);
and U3608 (N_3608,N_3536,N_3544);
xnor U3609 (N_3609,N_3566,N_3572);
and U3610 (N_3610,N_3538,N_3491);
nand U3611 (N_3611,N_3451,N_3542);
or U3612 (N_3612,N_3500,N_3456);
or U3613 (N_3613,N_3453,N_3473);
nand U3614 (N_3614,N_3485,N_3474);
nor U3615 (N_3615,N_3576,N_3475);
xor U3616 (N_3616,N_3521,N_3452);
nor U3617 (N_3617,N_3561,N_3575);
or U3618 (N_3618,N_3594,N_3462);
xor U3619 (N_3619,N_3570,N_3519);
and U3620 (N_3620,N_3508,N_3595);
nand U3621 (N_3621,N_3534,N_3551);
and U3622 (N_3622,N_3555,N_3481);
nor U3623 (N_3623,N_3487,N_3562);
xor U3624 (N_3624,N_3589,N_3556);
nor U3625 (N_3625,N_3506,N_3524);
or U3626 (N_3626,N_3466,N_3548);
nand U3627 (N_3627,N_3552,N_3455);
xnor U3628 (N_3628,N_3584,N_3531);
and U3629 (N_3629,N_3514,N_3484);
xor U3630 (N_3630,N_3590,N_3459);
and U3631 (N_3631,N_3550,N_3547);
and U3632 (N_3632,N_3493,N_3533);
nand U3633 (N_3633,N_3472,N_3591);
nor U3634 (N_3634,N_3469,N_3518);
xnor U3635 (N_3635,N_3479,N_3537);
nor U3636 (N_3636,N_3579,N_3593);
and U3637 (N_3637,N_3523,N_3558);
xor U3638 (N_3638,N_3510,N_3482);
xor U3639 (N_3639,N_3557,N_3565);
or U3640 (N_3640,N_3578,N_3461);
nor U3641 (N_3641,N_3568,N_3549);
xor U3642 (N_3642,N_3498,N_3497);
and U3643 (N_3643,N_3545,N_3509);
nand U3644 (N_3644,N_3571,N_3489);
nand U3645 (N_3645,N_3490,N_3564);
or U3646 (N_3646,N_3511,N_3458);
and U3647 (N_3647,N_3470,N_3582);
nand U3648 (N_3648,N_3480,N_3526);
and U3649 (N_3649,N_3463,N_3597);
nand U3650 (N_3650,N_3471,N_3520);
nand U3651 (N_3651,N_3553,N_3483);
xnor U3652 (N_3652,N_3580,N_3488);
and U3653 (N_3653,N_3504,N_3583);
nor U3654 (N_3654,N_3560,N_3450);
nand U3655 (N_3655,N_3527,N_3477);
xnor U3656 (N_3656,N_3599,N_3501);
and U3657 (N_3657,N_3496,N_3465);
nand U3658 (N_3658,N_3464,N_3559);
nor U3659 (N_3659,N_3569,N_3478);
nor U3660 (N_3660,N_3581,N_3467);
or U3661 (N_3661,N_3540,N_3503);
nor U3662 (N_3662,N_3532,N_3598);
xnor U3663 (N_3663,N_3486,N_3512);
and U3664 (N_3664,N_3535,N_3588);
and U3665 (N_3665,N_3541,N_3586);
or U3666 (N_3666,N_3596,N_3457);
nor U3667 (N_3667,N_3529,N_3587);
or U3668 (N_3668,N_3554,N_3517);
or U3669 (N_3669,N_3530,N_3539);
xnor U3670 (N_3670,N_3495,N_3585);
xnor U3671 (N_3671,N_3499,N_3513);
and U3672 (N_3672,N_3573,N_3563);
xnor U3673 (N_3673,N_3507,N_3505);
xor U3674 (N_3674,N_3577,N_3476);
and U3675 (N_3675,N_3506,N_3465);
or U3676 (N_3676,N_3515,N_3572);
and U3677 (N_3677,N_3535,N_3579);
xor U3678 (N_3678,N_3497,N_3533);
and U3679 (N_3679,N_3541,N_3594);
or U3680 (N_3680,N_3454,N_3492);
and U3681 (N_3681,N_3584,N_3527);
nor U3682 (N_3682,N_3460,N_3471);
nor U3683 (N_3683,N_3557,N_3502);
nand U3684 (N_3684,N_3584,N_3504);
nand U3685 (N_3685,N_3586,N_3522);
nor U3686 (N_3686,N_3486,N_3527);
and U3687 (N_3687,N_3506,N_3565);
and U3688 (N_3688,N_3526,N_3455);
and U3689 (N_3689,N_3579,N_3584);
and U3690 (N_3690,N_3489,N_3596);
and U3691 (N_3691,N_3481,N_3470);
nand U3692 (N_3692,N_3460,N_3594);
or U3693 (N_3693,N_3515,N_3552);
nor U3694 (N_3694,N_3515,N_3452);
and U3695 (N_3695,N_3473,N_3518);
and U3696 (N_3696,N_3586,N_3508);
nor U3697 (N_3697,N_3559,N_3539);
and U3698 (N_3698,N_3585,N_3482);
xnor U3699 (N_3699,N_3478,N_3562);
nor U3700 (N_3700,N_3557,N_3461);
and U3701 (N_3701,N_3490,N_3509);
xor U3702 (N_3702,N_3598,N_3537);
and U3703 (N_3703,N_3574,N_3466);
xnor U3704 (N_3704,N_3479,N_3593);
xor U3705 (N_3705,N_3481,N_3564);
nor U3706 (N_3706,N_3458,N_3474);
xor U3707 (N_3707,N_3593,N_3507);
or U3708 (N_3708,N_3499,N_3461);
nand U3709 (N_3709,N_3597,N_3501);
or U3710 (N_3710,N_3506,N_3489);
xor U3711 (N_3711,N_3502,N_3526);
nand U3712 (N_3712,N_3545,N_3515);
nand U3713 (N_3713,N_3560,N_3567);
or U3714 (N_3714,N_3536,N_3463);
xnor U3715 (N_3715,N_3450,N_3464);
and U3716 (N_3716,N_3482,N_3578);
nand U3717 (N_3717,N_3561,N_3595);
nand U3718 (N_3718,N_3515,N_3550);
nand U3719 (N_3719,N_3477,N_3501);
nor U3720 (N_3720,N_3564,N_3541);
and U3721 (N_3721,N_3549,N_3536);
or U3722 (N_3722,N_3486,N_3529);
nand U3723 (N_3723,N_3597,N_3556);
or U3724 (N_3724,N_3512,N_3579);
nand U3725 (N_3725,N_3453,N_3532);
nand U3726 (N_3726,N_3513,N_3450);
or U3727 (N_3727,N_3485,N_3477);
xor U3728 (N_3728,N_3567,N_3562);
and U3729 (N_3729,N_3531,N_3567);
xnor U3730 (N_3730,N_3562,N_3493);
and U3731 (N_3731,N_3513,N_3576);
xnor U3732 (N_3732,N_3536,N_3565);
nand U3733 (N_3733,N_3484,N_3476);
and U3734 (N_3734,N_3527,N_3461);
nor U3735 (N_3735,N_3470,N_3472);
nand U3736 (N_3736,N_3572,N_3491);
nor U3737 (N_3737,N_3591,N_3521);
or U3738 (N_3738,N_3589,N_3587);
nor U3739 (N_3739,N_3503,N_3595);
and U3740 (N_3740,N_3527,N_3572);
nand U3741 (N_3741,N_3583,N_3491);
or U3742 (N_3742,N_3512,N_3588);
xnor U3743 (N_3743,N_3560,N_3527);
or U3744 (N_3744,N_3479,N_3585);
nor U3745 (N_3745,N_3462,N_3530);
or U3746 (N_3746,N_3554,N_3515);
xor U3747 (N_3747,N_3583,N_3546);
nor U3748 (N_3748,N_3519,N_3505);
nor U3749 (N_3749,N_3479,N_3469);
nor U3750 (N_3750,N_3657,N_3644);
and U3751 (N_3751,N_3622,N_3647);
xnor U3752 (N_3752,N_3678,N_3618);
xnor U3753 (N_3753,N_3630,N_3649);
or U3754 (N_3754,N_3674,N_3613);
nor U3755 (N_3755,N_3661,N_3740);
nand U3756 (N_3756,N_3696,N_3634);
nand U3757 (N_3757,N_3608,N_3664);
or U3758 (N_3758,N_3667,N_3737);
or U3759 (N_3759,N_3689,N_3639);
xnor U3760 (N_3760,N_3706,N_3698);
nor U3761 (N_3761,N_3728,N_3628);
nor U3762 (N_3762,N_3610,N_3623);
nor U3763 (N_3763,N_3617,N_3717);
and U3764 (N_3764,N_3741,N_3645);
or U3765 (N_3765,N_3676,N_3738);
nor U3766 (N_3766,N_3609,N_3654);
nor U3767 (N_3767,N_3747,N_3725);
xor U3768 (N_3768,N_3614,N_3633);
xor U3769 (N_3769,N_3697,N_3669);
xor U3770 (N_3770,N_3611,N_3724);
and U3771 (N_3771,N_3632,N_3641);
nand U3772 (N_3772,N_3665,N_3708);
and U3773 (N_3773,N_3624,N_3694);
or U3774 (N_3774,N_3663,N_3681);
and U3775 (N_3775,N_3638,N_3686);
and U3776 (N_3776,N_3659,N_3627);
xor U3777 (N_3777,N_3606,N_3710);
nand U3778 (N_3778,N_3726,N_3746);
xnor U3779 (N_3779,N_3626,N_3736);
nor U3780 (N_3780,N_3707,N_3677);
nand U3781 (N_3781,N_3733,N_3720);
nand U3782 (N_3782,N_3643,N_3673);
nand U3783 (N_3783,N_3636,N_3684);
nor U3784 (N_3784,N_3703,N_3629);
and U3785 (N_3785,N_3642,N_3687);
nor U3786 (N_3786,N_3715,N_3704);
and U3787 (N_3787,N_3732,N_3739);
and U3788 (N_3788,N_3672,N_3668);
or U3789 (N_3789,N_3682,N_3603);
xnor U3790 (N_3790,N_3727,N_3621);
xor U3791 (N_3791,N_3619,N_3702);
nand U3792 (N_3792,N_3734,N_3713);
nor U3793 (N_3793,N_3602,N_3666);
nand U3794 (N_3794,N_3692,N_3662);
nor U3795 (N_3795,N_3607,N_3709);
and U3796 (N_3796,N_3658,N_3660);
or U3797 (N_3797,N_3721,N_3745);
nor U3798 (N_3798,N_3731,N_3651);
or U3799 (N_3799,N_3656,N_3735);
nand U3800 (N_3800,N_3716,N_3695);
or U3801 (N_3801,N_3699,N_3693);
xor U3802 (N_3802,N_3671,N_3719);
nor U3803 (N_3803,N_3712,N_3652);
or U3804 (N_3804,N_3705,N_3748);
nor U3805 (N_3805,N_3718,N_3635);
xor U3806 (N_3806,N_3729,N_3653);
nor U3807 (N_3807,N_3749,N_3616);
and U3808 (N_3808,N_3675,N_3730);
or U3809 (N_3809,N_3742,N_3679);
and U3810 (N_3810,N_3714,N_3615);
and U3811 (N_3811,N_3722,N_3688);
xnor U3812 (N_3812,N_3655,N_3744);
xor U3813 (N_3813,N_3604,N_3711);
and U3814 (N_3814,N_3648,N_3685);
nand U3815 (N_3815,N_3690,N_3680);
xor U3816 (N_3816,N_3646,N_3625);
and U3817 (N_3817,N_3691,N_3670);
nand U3818 (N_3818,N_3637,N_3650);
or U3819 (N_3819,N_3600,N_3743);
nor U3820 (N_3820,N_3683,N_3620);
and U3821 (N_3821,N_3723,N_3631);
xnor U3822 (N_3822,N_3700,N_3612);
xor U3823 (N_3823,N_3640,N_3601);
and U3824 (N_3824,N_3701,N_3605);
and U3825 (N_3825,N_3686,N_3718);
nor U3826 (N_3826,N_3659,N_3701);
nor U3827 (N_3827,N_3669,N_3628);
nor U3828 (N_3828,N_3602,N_3708);
xnor U3829 (N_3829,N_3673,N_3709);
xnor U3830 (N_3830,N_3726,N_3651);
and U3831 (N_3831,N_3665,N_3617);
xnor U3832 (N_3832,N_3706,N_3689);
or U3833 (N_3833,N_3642,N_3747);
nor U3834 (N_3834,N_3663,N_3676);
xnor U3835 (N_3835,N_3615,N_3672);
nor U3836 (N_3836,N_3639,N_3610);
or U3837 (N_3837,N_3629,N_3680);
and U3838 (N_3838,N_3742,N_3641);
or U3839 (N_3839,N_3644,N_3741);
nand U3840 (N_3840,N_3716,N_3607);
or U3841 (N_3841,N_3604,N_3665);
nand U3842 (N_3842,N_3609,N_3660);
nand U3843 (N_3843,N_3672,N_3709);
xor U3844 (N_3844,N_3634,N_3667);
nor U3845 (N_3845,N_3700,N_3678);
and U3846 (N_3846,N_3653,N_3665);
and U3847 (N_3847,N_3695,N_3706);
nand U3848 (N_3848,N_3615,N_3648);
xor U3849 (N_3849,N_3748,N_3615);
xnor U3850 (N_3850,N_3689,N_3716);
and U3851 (N_3851,N_3726,N_3696);
nor U3852 (N_3852,N_3705,N_3728);
xnor U3853 (N_3853,N_3727,N_3664);
and U3854 (N_3854,N_3622,N_3727);
nor U3855 (N_3855,N_3627,N_3628);
nor U3856 (N_3856,N_3604,N_3615);
xnor U3857 (N_3857,N_3708,N_3723);
and U3858 (N_3858,N_3717,N_3646);
nor U3859 (N_3859,N_3701,N_3653);
and U3860 (N_3860,N_3615,N_3628);
nand U3861 (N_3861,N_3667,N_3715);
nand U3862 (N_3862,N_3632,N_3630);
nor U3863 (N_3863,N_3611,N_3734);
nand U3864 (N_3864,N_3689,N_3629);
nand U3865 (N_3865,N_3633,N_3673);
and U3866 (N_3866,N_3665,N_3630);
or U3867 (N_3867,N_3657,N_3650);
and U3868 (N_3868,N_3636,N_3601);
and U3869 (N_3869,N_3735,N_3630);
and U3870 (N_3870,N_3607,N_3649);
or U3871 (N_3871,N_3623,N_3704);
nand U3872 (N_3872,N_3623,N_3613);
nand U3873 (N_3873,N_3727,N_3615);
and U3874 (N_3874,N_3716,N_3726);
or U3875 (N_3875,N_3662,N_3600);
or U3876 (N_3876,N_3651,N_3669);
xnor U3877 (N_3877,N_3696,N_3692);
xnor U3878 (N_3878,N_3706,N_3714);
and U3879 (N_3879,N_3611,N_3605);
nand U3880 (N_3880,N_3622,N_3624);
and U3881 (N_3881,N_3704,N_3713);
nor U3882 (N_3882,N_3700,N_3680);
nand U3883 (N_3883,N_3696,N_3724);
and U3884 (N_3884,N_3621,N_3605);
xor U3885 (N_3885,N_3635,N_3634);
and U3886 (N_3886,N_3637,N_3714);
xor U3887 (N_3887,N_3688,N_3623);
xnor U3888 (N_3888,N_3738,N_3679);
nor U3889 (N_3889,N_3632,N_3722);
nor U3890 (N_3890,N_3699,N_3663);
nor U3891 (N_3891,N_3688,N_3727);
and U3892 (N_3892,N_3742,N_3640);
or U3893 (N_3893,N_3631,N_3669);
and U3894 (N_3894,N_3600,N_3744);
nand U3895 (N_3895,N_3673,N_3629);
xor U3896 (N_3896,N_3662,N_3616);
xor U3897 (N_3897,N_3694,N_3639);
or U3898 (N_3898,N_3606,N_3623);
xor U3899 (N_3899,N_3611,N_3727);
xnor U3900 (N_3900,N_3774,N_3855);
nand U3901 (N_3901,N_3762,N_3876);
or U3902 (N_3902,N_3753,N_3884);
xor U3903 (N_3903,N_3798,N_3870);
or U3904 (N_3904,N_3813,N_3807);
xnor U3905 (N_3905,N_3852,N_3898);
nand U3906 (N_3906,N_3827,N_3810);
and U3907 (N_3907,N_3846,N_3819);
or U3908 (N_3908,N_3880,N_3772);
nor U3909 (N_3909,N_3869,N_3773);
nand U3910 (N_3910,N_3857,N_3808);
and U3911 (N_3911,N_3867,N_3842);
nand U3912 (N_3912,N_3801,N_3775);
nand U3913 (N_3913,N_3860,N_3838);
or U3914 (N_3914,N_3790,N_3864);
nand U3915 (N_3915,N_3851,N_3854);
and U3916 (N_3916,N_3796,N_3850);
or U3917 (N_3917,N_3766,N_3778);
nand U3918 (N_3918,N_3805,N_3763);
nor U3919 (N_3919,N_3814,N_3824);
and U3920 (N_3920,N_3868,N_3768);
nand U3921 (N_3921,N_3845,N_3820);
and U3922 (N_3922,N_3866,N_3800);
nand U3923 (N_3923,N_3887,N_3816);
or U3924 (N_3924,N_3828,N_3879);
or U3925 (N_3925,N_3761,N_3817);
nand U3926 (N_3926,N_3751,N_3750);
and U3927 (N_3927,N_3835,N_3831);
nand U3928 (N_3928,N_3878,N_3812);
nor U3929 (N_3929,N_3897,N_3840);
xnor U3930 (N_3930,N_3767,N_3765);
xor U3931 (N_3931,N_3889,N_3858);
nand U3932 (N_3932,N_3861,N_3841);
or U3933 (N_3933,N_3754,N_3795);
xnor U3934 (N_3934,N_3776,N_3797);
nand U3935 (N_3935,N_3830,N_3882);
or U3936 (N_3936,N_3883,N_3771);
and U3937 (N_3937,N_3769,N_3779);
and U3938 (N_3938,N_3781,N_3822);
or U3939 (N_3939,N_3821,N_3863);
xnor U3940 (N_3940,N_3755,N_3794);
nand U3941 (N_3941,N_3833,N_3825);
xnor U3942 (N_3942,N_3756,N_3802);
or U3943 (N_3943,N_3894,N_3764);
and U3944 (N_3944,N_3752,N_3760);
xnor U3945 (N_3945,N_3859,N_3886);
or U3946 (N_3946,N_3777,N_3865);
and U3947 (N_3947,N_3849,N_3871);
or U3948 (N_3948,N_3899,N_3892);
xor U3949 (N_3949,N_3784,N_3856);
and U3950 (N_3950,N_3823,N_3847);
nand U3951 (N_3951,N_3832,N_3792);
nor U3952 (N_3952,N_3788,N_3789);
xor U3953 (N_3953,N_3888,N_3844);
or U3954 (N_3954,N_3786,N_3829);
xnor U3955 (N_3955,N_3785,N_3834);
and U3956 (N_3956,N_3891,N_3799);
nand U3957 (N_3957,N_3896,N_3780);
nor U3958 (N_3958,N_3818,N_3836);
xnor U3959 (N_3959,N_3893,N_3895);
nor U3960 (N_3960,N_3853,N_3873);
or U3961 (N_3961,N_3885,N_3793);
nand U3962 (N_3962,N_3815,N_3787);
and U3963 (N_3963,N_3848,N_3811);
and U3964 (N_3964,N_3782,N_3875);
nand U3965 (N_3965,N_3890,N_3843);
or U3966 (N_3966,N_3809,N_3837);
nor U3967 (N_3967,N_3874,N_3783);
and U3968 (N_3968,N_3804,N_3872);
xnor U3969 (N_3969,N_3826,N_3806);
and U3970 (N_3970,N_3803,N_3881);
or U3971 (N_3971,N_3770,N_3759);
or U3972 (N_3972,N_3839,N_3758);
or U3973 (N_3973,N_3791,N_3757);
and U3974 (N_3974,N_3877,N_3862);
and U3975 (N_3975,N_3781,N_3808);
or U3976 (N_3976,N_3783,N_3831);
and U3977 (N_3977,N_3814,N_3802);
nand U3978 (N_3978,N_3838,N_3889);
nand U3979 (N_3979,N_3785,N_3814);
nor U3980 (N_3980,N_3877,N_3810);
xor U3981 (N_3981,N_3757,N_3868);
nand U3982 (N_3982,N_3798,N_3875);
and U3983 (N_3983,N_3860,N_3808);
xor U3984 (N_3984,N_3897,N_3822);
or U3985 (N_3985,N_3766,N_3780);
or U3986 (N_3986,N_3852,N_3886);
xnor U3987 (N_3987,N_3847,N_3840);
nand U3988 (N_3988,N_3784,N_3843);
xor U3989 (N_3989,N_3819,N_3779);
nor U3990 (N_3990,N_3847,N_3777);
and U3991 (N_3991,N_3836,N_3850);
xor U3992 (N_3992,N_3797,N_3829);
xor U3993 (N_3993,N_3826,N_3844);
nand U3994 (N_3994,N_3764,N_3874);
nand U3995 (N_3995,N_3768,N_3843);
xnor U3996 (N_3996,N_3802,N_3804);
nor U3997 (N_3997,N_3850,N_3767);
nand U3998 (N_3998,N_3836,N_3756);
nand U3999 (N_3999,N_3783,N_3842);
and U4000 (N_4000,N_3797,N_3835);
nor U4001 (N_4001,N_3765,N_3818);
or U4002 (N_4002,N_3814,N_3837);
and U4003 (N_4003,N_3853,N_3795);
or U4004 (N_4004,N_3878,N_3796);
nand U4005 (N_4005,N_3868,N_3880);
nor U4006 (N_4006,N_3837,N_3873);
and U4007 (N_4007,N_3797,N_3884);
nand U4008 (N_4008,N_3775,N_3777);
nor U4009 (N_4009,N_3757,N_3760);
or U4010 (N_4010,N_3802,N_3810);
nor U4011 (N_4011,N_3780,N_3750);
nand U4012 (N_4012,N_3858,N_3893);
and U4013 (N_4013,N_3801,N_3840);
xnor U4014 (N_4014,N_3861,N_3834);
or U4015 (N_4015,N_3847,N_3820);
or U4016 (N_4016,N_3836,N_3874);
and U4017 (N_4017,N_3783,N_3820);
or U4018 (N_4018,N_3817,N_3859);
or U4019 (N_4019,N_3894,N_3851);
or U4020 (N_4020,N_3823,N_3771);
and U4021 (N_4021,N_3874,N_3883);
nand U4022 (N_4022,N_3752,N_3826);
or U4023 (N_4023,N_3894,N_3823);
and U4024 (N_4024,N_3765,N_3863);
nand U4025 (N_4025,N_3772,N_3805);
and U4026 (N_4026,N_3870,N_3898);
or U4027 (N_4027,N_3784,N_3832);
xor U4028 (N_4028,N_3885,N_3856);
and U4029 (N_4029,N_3845,N_3841);
xnor U4030 (N_4030,N_3815,N_3835);
xor U4031 (N_4031,N_3784,N_3801);
nor U4032 (N_4032,N_3844,N_3879);
and U4033 (N_4033,N_3888,N_3852);
or U4034 (N_4034,N_3899,N_3874);
or U4035 (N_4035,N_3892,N_3776);
or U4036 (N_4036,N_3776,N_3804);
nor U4037 (N_4037,N_3765,N_3898);
or U4038 (N_4038,N_3882,N_3760);
or U4039 (N_4039,N_3801,N_3783);
nor U4040 (N_4040,N_3765,N_3797);
nor U4041 (N_4041,N_3827,N_3788);
or U4042 (N_4042,N_3882,N_3874);
xor U4043 (N_4043,N_3776,N_3890);
nor U4044 (N_4044,N_3766,N_3891);
xor U4045 (N_4045,N_3750,N_3831);
nor U4046 (N_4046,N_3832,N_3869);
and U4047 (N_4047,N_3861,N_3821);
nor U4048 (N_4048,N_3753,N_3792);
or U4049 (N_4049,N_3761,N_3793);
nand U4050 (N_4050,N_4026,N_3999);
nor U4051 (N_4051,N_3981,N_4043);
and U4052 (N_4052,N_3946,N_4042);
nand U4053 (N_4053,N_3955,N_3976);
nand U4054 (N_4054,N_3920,N_3959);
nand U4055 (N_4055,N_4035,N_3963);
and U4056 (N_4056,N_3915,N_3939);
xnor U4057 (N_4057,N_4005,N_3912);
and U4058 (N_4058,N_3944,N_3934);
nand U4059 (N_4059,N_4003,N_4034);
nor U4060 (N_4060,N_4041,N_3953);
nand U4061 (N_4061,N_3996,N_3991);
xnor U4062 (N_4062,N_4029,N_3913);
or U4063 (N_4063,N_4024,N_3979);
nand U4064 (N_4064,N_3970,N_4016);
or U4065 (N_4065,N_3975,N_3907);
xnor U4066 (N_4066,N_3997,N_3935);
nand U4067 (N_4067,N_3972,N_3983);
xnor U4068 (N_4068,N_3958,N_4032);
or U4069 (N_4069,N_3998,N_4006);
xnor U4070 (N_4070,N_3916,N_4038);
and U4071 (N_4071,N_3901,N_3965);
xnor U4072 (N_4072,N_4019,N_3921);
nor U4073 (N_4073,N_3966,N_3940);
or U4074 (N_4074,N_3994,N_3962);
nand U4075 (N_4075,N_4025,N_3995);
nand U4076 (N_4076,N_4046,N_3904);
nand U4077 (N_4077,N_4002,N_3984);
nor U4078 (N_4078,N_3918,N_4001);
xnor U4079 (N_4079,N_4030,N_3951);
nand U4080 (N_4080,N_4021,N_3949);
and U4081 (N_4081,N_3968,N_3914);
nand U4082 (N_4082,N_4004,N_4044);
or U4083 (N_4083,N_3993,N_3945);
and U4084 (N_4084,N_3989,N_3924);
nand U4085 (N_4085,N_4020,N_3985);
and U4086 (N_4086,N_3917,N_3988);
and U4087 (N_4087,N_3906,N_3900);
nand U4088 (N_4088,N_3971,N_3933);
xor U4089 (N_4089,N_3919,N_3908);
xnor U4090 (N_4090,N_4022,N_3909);
and U4091 (N_4091,N_4012,N_3932);
nand U4092 (N_4092,N_3936,N_4027);
nand U4093 (N_4093,N_4028,N_3957);
nand U4094 (N_4094,N_3974,N_3973);
nor U4095 (N_4095,N_3969,N_4008);
nor U4096 (N_4096,N_3905,N_4000);
or U4097 (N_4097,N_4048,N_4036);
nor U4098 (N_4098,N_3987,N_3992);
or U4099 (N_4099,N_4018,N_4023);
and U4100 (N_4100,N_3964,N_3931);
xor U4101 (N_4101,N_3947,N_3942);
nor U4102 (N_4102,N_3980,N_4039);
and U4103 (N_4103,N_4007,N_4011);
nand U4104 (N_4104,N_3938,N_3960);
or U4105 (N_4105,N_4017,N_3948);
and U4106 (N_4106,N_3922,N_4010);
nand U4107 (N_4107,N_4031,N_3937);
nor U4108 (N_4108,N_3902,N_4033);
and U4109 (N_4109,N_3978,N_4045);
nand U4110 (N_4110,N_4037,N_3943);
xor U4111 (N_4111,N_4009,N_3982);
and U4112 (N_4112,N_3910,N_4040);
nand U4113 (N_4113,N_3911,N_3954);
nor U4114 (N_4114,N_3923,N_3977);
nor U4115 (N_4115,N_3928,N_3929);
xnor U4116 (N_4116,N_3952,N_4015);
and U4117 (N_4117,N_4013,N_3967);
nand U4118 (N_4118,N_3930,N_4047);
xor U4119 (N_4119,N_3925,N_3990);
nand U4120 (N_4120,N_4014,N_3927);
or U4121 (N_4121,N_3950,N_4049);
nor U4122 (N_4122,N_3903,N_3956);
or U4123 (N_4123,N_3986,N_3941);
nand U4124 (N_4124,N_3926,N_3961);
and U4125 (N_4125,N_4042,N_3910);
nand U4126 (N_4126,N_4045,N_3999);
nand U4127 (N_4127,N_3968,N_4027);
and U4128 (N_4128,N_3928,N_3904);
or U4129 (N_4129,N_4001,N_3978);
or U4130 (N_4130,N_3911,N_3908);
or U4131 (N_4131,N_3934,N_3943);
nor U4132 (N_4132,N_3981,N_3925);
nor U4133 (N_4133,N_4047,N_4022);
xor U4134 (N_4134,N_4016,N_4047);
or U4135 (N_4135,N_4025,N_4013);
xor U4136 (N_4136,N_3929,N_3921);
or U4137 (N_4137,N_4028,N_3920);
or U4138 (N_4138,N_3969,N_3966);
xor U4139 (N_4139,N_3988,N_3991);
or U4140 (N_4140,N_3917,N_4024);
xor U4141 (N_4141,N_4010,N_3917);
xnor U4142 (N_4142,N_4015,N_3994);
nor U4143 (N_4143,N_3978,N_3986);
nor U4144 (N_4144,N_3947,N_4006);
nor U4145 (N_4145,N_3948,N_4034);
and U4146 (N_4146,N_3914,N_3946);
nor U4147 (N_4147,N_3953,N_3908);
nor U4148 (N_4148,N_3998,N_4036);
or U4149 (N_4149,N_4034,N_3946);
nand U4150 (N_4150,N_3999,N_3991);
nand U4151 (N_4151,N_3922,N_3946);
or U4152 (N_4152,N_3938,N_3979);
xor U4153 (N_4153,N_3949,N_3947);
or U4154 (N_4154,N_4021,N_4016);
nor U4155 (N_4155,N_4014,N_4046);
nor U4156 (N_4156,N_4001,N_4005);
nand U4157 (N_4157,N_3918,N_4033);
xor U4158 (N_4158,N_3941,N_3983);
nor U4159 (N_4159,N_4015,N_3944);
xnor U4160 (N_4160,N_3977,N_4046);
nand U4161 (N_4161,N_3972,N_4023);
xor U4162 (N_4162,N_3986,N_3975);
xor U4163 (N_4163,N_3916,N_3940);
nand U4164 (N_4164,N_4045,N_4049);
xor U4165 (N_4165,N_3915,N_4012);
or U4166 (N_4166,N_3919,N_4002);
nand U4167 (N_4167,N_3954,N_3921);
nand U4168 (N_4168,N_3933,N_4011);
nor U4169 (N_4169,N_3908,N_4025);
or U4170 (N_4170,N_3916,N_4023);
and U4171 (N_4171,N_3967,N_3964);
nor U4172 (N_4172,N_3933,N_3916);
or U4173 (N_4173,N_3964,N_3987);
nor U4174 (N_4174,N_3967,N_3919);
nand U4175 (N_4175,N_4037,N_3959);
xnor U4176 (N_4176,N_3902,N_3964);
xor U4177 (N_4177,N_4008,N_3976);
and U4178 (N_4178,N_4002,N_3995);
and U4179 (N_4179,N_3916,N_3986);
xnor U4180 (N_4180,N_3942,N_4025);
nor U4181 (N_4181,N_3900,N_3915);
xnor U4182 (N_4182,N_4032,N_3905);
xnor U4183 (N_4183,N_3949,N_3900);
nor U4184 (N_4184,N_4033,N_4018);
nor U4185 (N_4185,N_3910,N_3900);
xor U4186 (N_4186,N_3960,N_3923);
or U4187 (N_4187,N_4036,N_4015);
xnor U4188 (N_4188,N_3942,N_4010);
xor U4189 (N_4189,N_4034,N_3905);
and U4190 (N_4190,N_4036,N_3949);
xnor U4191 (N_4191,N_3914,N_4043);
nor U4192 (N_4192,N_4001,N_4012);
nand U4193 (N_4193,N_4047,N_3977);
and U4194 (N_4194,N_3966,N_3924);
nand U4195 (N_4195,N_3989,N_4038);
nand U4196 (N_4196,N_3901,N_4034);
nand U4197 (N_4197,N_3909,N_3944);
xor U4198 (N_4198,N_3920,N_3909);
and U4199 (N_4199,N_3998,N_3909);
xor U4200 (N_4200,N_4068,N_4053);
nand U4201 (N_4201,N_4097,N_4092);
xor U4202 (N_4202,N_4051,N_4136);
nor U4203 (N_4203,N_4098,N_4192);
nor U4204 (N_4204,N_4126,N_4179);
nand U4205 (N_4205,N_4141,N_4055);
or U4206 (N_4206,N_4195,N_4071);
nor U4207 (N_4207,N_4086,N_4165);
and U4208 (N_4208,N_4130,N_4148);
nand U4209 (N_4209,N_4105,N_4056);
nand U4210 (N_4210,N_4065,N_4103);
xor U4211 (N_4211,N_4096,N_4145);
or U4212 (N_4212,N_4158,N_4157);
nor U4213 (N_4213,N_4162,N_4111);
and U4214 (N_4214,N_4133,N_4110);
nand U4215 (N_4215,N_4134,N_4182);
or U4216 (N_4216,N_4198,N_4102);
and U4217 (N_4217,N_4135,N_4172);
xor U4218 (N_4218,N_4074,N_4109);
or U4219 (N_4219,N_4089,N_4058);
and U4220 (N_4220,N_4112,N_4164);
or U4221 (N_4221,N_4189,N_4088);
nor U4222 (N_4222,N_4142,N_4168);
nand U4223 (N_4223,N_4194,N_4095);
xor U4224 (N_4224,N_4060,N_4147);
or U4225 (N_4225,N_4197,N_4193);
nand U4226 (N_4226,N_4072,N_4069);
xor U4227 (N_4227,N_4117,N_4116);
or U4228 (N_4228,N_4090,N_4137);
nand U4229 (N_4229,N_4139,N_4191);
nor U4230 (N_4230,N_4199,N_4094);
nand U4231 (N_4231,N_4155,N_4101);
nor U4232 (N_4232,N_4064,N_4124);
xnor U4233 (N_4233,N_4087,N_4156);
nand U4234 (N_4234,N_4119,N_4067);
and U4235 (N_4235,N_4076,N_4151);
nor U4236 (N_4236,N_4099,N_4093);
nor U4237 (N_4237,N_4132,N_4140);
xor U4238 (N_4238,N_4059,N_4153);
or U4239 (N_4239,N_4079,N_4078);
and U4240 (N_4240,N_4146,N_4077);
nand U4241 (N_4241,N_4108,N_4169);
nand U4242 (N_4242,N_4122,N_4175);
xnor U4243 (N_4243,N_4063,N_4075);
xor U4244 (N_4244,N_4170,N_4129);
nand U4245 (N_4245,N_4138,N_4123);
and U4246 (N_4246,N_4161,N_4167);
nand U4247 (N_4247,N_4066,N_4100);
nand U4248 (N_4248,N_4073,N_4085);
and U4249 (N_4249,N_4106,N_4149);
nor U4250 (N_4250,N_4061,N_4176);
xor U4251 (N_4251,N_4080,N_4190);
nor U4252 (N_4252,N_4180,N_4188);
nor U4253 (N_4253,N_4062,N_4154);
nor U4254 (N_4254,N_4082,N_4125);
and U4255 (N_4255,N_4196,N_4104);
nand U4256 (N_4256,N_4091,N_4113);
nand U4257 (N_4257,N_4177,N_4181);
nand U4258 (N_4258,N_4143,N_4178);
or U4259 (N_4259,N_4083,N_4050);
nor U4260 (N_4260,N_4120,N_4121);
and U4261 (N_4261,N_4183,N_4166);
or U4262 (N_4262,N_4115,N_4159);
xnor U4263 (N_4263,N_4127,N_4081);
and U4264 (N_4264,N_4152,N_4186);
nor U4265 (N_4265,N_4171,N_4150);
xnor U4266 (N_4266,N_4128,N_4054);
and U4267 (N_4267,N_4107,N_4084);
nand U4268 (N_4268,N_4144,N_4187);
or U4269 (N_4269,N_4163,N_4118);
nor U4270 (N_4270,N_4114,N_4070);
and U4271 (N_4271,N_4057,N_4052);
xnor U4272 (N_4272,N_4174,N_4131);
xor U4273 (N_4273,N_4173,N_4160);
and U4274 (N_4274,N_4184,N_4185);
xnor U4275 (N_4275,N_4181,N_4157);
nor U4276 (N_4276,N_4136,N_4181);
nand U4277 (N_4277,N_4188,N_4076);
xnor U4278 (N_4278,N_4163,N_4170);
and U4279 (N_4279,N_4180,N_4074);
nor U4280 (N_4280,N_4181,N_4196);
or U4281 (N_4281,N_4146,N_4082);
nand U4282 (N_4282,N_4151,N_4067);
nand U4283 (N_4283,N_4169,N_4153);
nand U4284 (N_4284,N_4181,N_4113);
nand U4285 (N_4285,N_4096,N_4093);
nand U4286 (N_4286,N_4198,N_4146);
or U4287 (N_4287,N_4106,N_4060);
and U4288 (N_4288,N_4106,N_4077);
or U4289 (N_4289,N_4138,N_4181);
or U4290 (N_4290,N_4083,N_4194);
and U4291 (N_4291,N_4191,N_4192);
nand U4292 (N_4292,N_4186,N_4092);
nor U4293 (N_4293,N_4067,N_4152);
xor U4294 (N_4294,N_4178,N_4111);
nand U4295 (N_4295,N_4197,N_4082);
and U4296 (N_4296,N_4144,N_4139);
nand U4297 (N_4297,N_4183,N_4173);
and U4298 (N_4298,N_4176,N_4144);
xor U4299 (N_4299,N_4141,N_4079);
xnor U4300 (N_4300,N_4110,N_4119);
and U4301 (N_4301,N_4181,N_4182);
nor U4302 (N_4302,N_4091,N_4119);
nand U4303 (N_4303,N_4154,N_4162);
xor U4304 (N_4304,N_4072,N_4134);
or U4305 (N_4305,N_4143,N_4099);
nand U4306 (N_4306,N_4149,N_4055);
xnor U4307 (N_4307,N_4157,N_4159);
nor U4308 (N_4308,N_4168,N_4111);
and U4309 (N_4309,N_4053,N_4152);
nor U4310 (N_4310,N_4067,N_4078);
xnor U4311 (N_4311,N_4102,N_4060);
nor U4312 (N_4312,N_4077,N_4108);
xor U4313 (N_4313,N_4194,N_4075);
nor U4314 (N_4314,N_4171,N_4186);
xor U4315 (N_4315,N_4110,N_4147);
xnor U4316 (N_4316,N_4134,N_4095);
or U4317 (N_4317,N_4191,N_4193);
xor U4318 (N_4318,N_4075,N_4165);
and U4319 (N_4319,N_4065,N_4075);
nor U4320 (N_4320,N_4159,N_4183);
and U4321 (N_4321,N_4175,N_4096);
nand U4322 (N_4322,N_4196,N_4112);
xor U4323 (N_4323,N_4097,N_4085);
and U4324 (N_4324,N_4160,N_4098);
nand U4325 (N_4325,N_4114,N_4168);
nor U4326 (N_4326,N_4119,N_4139);
nor U4327 (N_4327,N_4063,N_4138);
xor U4328 (N_4328,N_4077,N_4125);
xnor U4329 (N_4329,N_4120,N_4081);
nor U4330 (N_4330,N_4078,N_4074);
xnor U4331 (N_4331,N_4075,N_4159);
nor U4332 (N_4332,N_4165,N_4097);
and U4333 (N_4333,N_4058,N_4100);
nor U4334 (N_4334,N_4111,N_4063);
or U4335 (N_4335,N_4050,N_4151);
or U4336 (N_4336,N_4134,N_4140);
or U4337 (N_4337,N_4108,N_4125);
nand U4338 (N_4338,N_4136,N_4146);
nand U4339 (N_4339,N_4126,N_4154);
nor U4340 (N_4340,N_4157,N_4077);
and U4341 (N_4341,N_4073,N_4152);
and U4342 (N_4342,N_4168,N_4184);
and U4343 (N_4343,N_4188,N_4166);
nand U4344 (N_4344,N_4081,N_4095);
xor U4345 (N_4345,N_4193,N_4062);
and U4346 (N_4346,N_4064,N_4122);
xnor U4347 (N_4347,N_4172,N_4156);
or U4348 (N_4348,N_4097,N_4186);
nand U4349 (N_4349,N_4093,N_4069);
or U4350 (N_4350,N_4243,N_4223);
and U4351 (N_4351,N_4345,N_4315);
and U4352 (N_4352,N_4284,N_4211);
or U4353 (N_4353,N_4203,N_4248);
nor U4354 (N_4354,N_4277,N_4256);
xor U4355 (N_4355,N_4282,N_4309);
nand U4356 (N_4356,N_4236,N_4327);
or U4357 (N_4357,N_4320,N_4279);
xor U4358 (N_4358,N_4251,N_4337);
and U4359 (N_4359,N_4205,N_4335);
nand U4360 (N_4360,N_4264,N_4202);
and U4361 (N_4361,N_4332,N_4340);
or U4362 (N_4362,N_4293,N_4213);
nor U4363 (N_4363,N_4275,N_4310);
or U4364 (N_4364,N_4334,N_4209);
nand U4365 (N_4365,N_4212,N_4220);
and U4366 (N_4366,N_4218,N_4253);
and U4367 (N_4367,N_4262,N_4291);
or U4368 (N_4368,N_4339,N_4246);
nor U4369 (N_4369,N_4240,N_4208);
xnor U4370 (N_4370,N_4272,N_4324);
nand U4371 (N_4371,N_4323,N_4235);
and U4372 (N_4372,N_4261,N_4299);
and U4373 (N_4373,N_4254,N_4311);
and U4374 (N_4374,N_4217,N_4244);
nand U4375 (N_4375,N_4297,N_4265);
nand U4376 (N_4376,N_4226,N_4347);
xnor U4377 (N_4377,N_4290,N_4349);
nor U4378 (N_4378,N_4319,N_4204);
nand U4379 (N_4379,N_4207,N_4329);
nand U4380 (N_4380,N_4242,N_4225);
xnor U4381 (N_4381,N_4305,N_4330);
xor U4382 (N_4382,N_4321,N_4325);
nand U4383 (N_4383,N_4214,N_4317);
and U4384 (N_4384,N_4241,N_4274);
and U4385 (N_4385,N_4318,N_4268);
nand U4386 (N_4386,N_4346,N_4287);
or U4387 (N_4387,N_4283,N_4338);
nand U4388 (N_4388,N_4331,N_4298);
nor U4389 (N_4389,N_4270,N_4238);
xnor U4390 (N_4390,N_4245,N_4234);
and U4391 (N_4391,N_4229,N_4228);
xor U4392 (N_4392,N_4210,N_4286);
xnor U4393 (N_4393,N_4322,N_4266);
xnor U4394 (N_4394,N_4271,N_4215);
or U4395 (N_4395,N_4206,N_4237);
nand U4396 (N_4396,N_4247,N_4222);
xor U4397 (N_4397,N_4280,N_4341);
xor U4398 (N_4398,N_4316,N_4255);
or U4399 (N_4399,N_4292,N_4273);
nor U4400 (N_4400,N_4239,N_4227);
nand U4401 (N_4401,N_4302,N_4296);
nand U4402 (N_4402,N_4333,N_4232);
or U4403 (N_4403,N_4257,N_4342);
and U4404 (N_4404,N_4259,N_4312);
or U4405 (N_4405,N_4278,N_4328);
or U4406 (N_4406,N_4231,N_4219);
nand U4407 (N_4407,N_4295,N_4221);
nand U4408 (N_4408,N_4267,N_4285);
and U4409 (N_4409,N_4269,N_4260);
and U4410 (N_4410,N_4303,N_4336);
nor U4411 (N_4411,N_4250,N_4304);
or U4412 (N_4412,N_4230,N_4258);
xnor U4413 (N_4413,N_4289,N_4301);
nand U4414 (N_4414,N_4344,N_4288);
nand U4415 (N_4415,N_4216,N_4348);
xnor U4416 (N_4416,N_4233,N_4343);
and U4417 (N_4417,N_4314,N_4326);
nand U4418 (N_4418,N_4294,N_4263);
nor U4419 (N_4419,N_4201,N_4252);
nand U4420 (N_4420,N_4276,N_4224);
xor U4421 (N_4421,N_4313,N_4249);
xor U4422 (N_4422,N_4200,N_4300);
xor U4423 (N_4423,N_4307,N_4306);
and U4424 (N_4424,N_4308,N_4281);
xor U4425 (N_4425,N_4267,N_4272);
xor U4426 (N_4426,N_4217,N_4245);
or U4427 (N_4427,N_4235,N_4202);
nor U4428 (N_4428,N_4291,N_4259);
nand U4429 (N_4429,N_4337,N_4289);
nand U4430 (N_4430,N_4322,N_4209);
and U4431 (N_4431,N_4223,N_4269);
or U4432 (N_4432,N_4327,N_4336);
xnor U4433 (N_4433,N_4211,N_4342);
nor U4434 (N_4434,N_4347,N_4345);
nand U4435 (N_4435,N_4240,N_4304);
xnor U4436 (N_4436,N_4207,N_4334);
nand U4437 (N_4437,N_4228,N_4304);
xnor U4438 (N_4438,N_4300,N_4303);
xor U4439 (N_4439,N_4249,N_4200);
or U4440 (N_4440,N_4338,N_4211);
nor U4441 (N_4441,N_4219,N_4280);
or U4442 (N_4442,N_4212,N_4254);
xnor U4443 (N_4443,N_4243,N_4318);
xor U4444 (N_4444,N_4254,N_4299);
nand U4445 (N_4445,N_4209,N_4264);
nand U4446 (N_4446,N_4248,N_4338);
xnor U4447 (N_4447,N_4228,N_4331);
and U4448 (N_4448,N_4308,N_4215);
nand U4449 (N_4449,N_4248,N_4226);
xnor U4450 (N_4450,N_4332,N_4303);
xor U4451 (N_4451,N_4300,N_4219);
nand U4452 (N_4452,N_4334,N_4308);
or U4453 (N_4453,N_4250,N_4230);
and U4454 (N_4454,N_4282,N_4244);
xor U4455 (N_4455,N_4249,N_4265);
xnor U4456 (N_4456,N_4211,N_4264);
and U4457 (N_4457,N_4329,N_4220);
and U4458 (N_4458,N_4317,N_4267);
xor U4459 (N_4459,N_4233,N_4239);
xor U4460 (N_4460,N_4346,N_4214);
xnor U4461 (N_4461,N_4243,N_4304);
and U4462 (N_4462,N_4279,N_4215);
or U4463 (N_4463,N_4226,N_4318);
nor U4464 (N_4464,N_4279,N_4265);
and U4465 (N_4465,N_4262,N_4213);
nand U4466 (N_4466,N_4274,N_4256);
and U4467 (N_4467,N_4271,N_4267);
nand U4468 (N_4468,N_4229,N_4210);
or U4469 (N_4469,N_4284,N_4342);
nand U4470 (N_4470,N_4334,N_4324);
or U4471 (N_4471,N_4238,N_4266);
and U4472 (N_4472,N_4268,N_4342);
nor U4473 (N_4473,N_4201,N_4266);
or U4474 (N_4474,N_4225,N_4347);
xnor U4475 (N_4475,N_4247,N_4254);
nand U4476 (N_4476,N_4220,N_4340);
nor U4477 (N_4477,N_4215,N_4219);
nor U4478 (N_4478,N_4210,N_4295);
xor U4479 (N_4479,N_4254,N_4301);
nor U4480 (N_4480,N_4286,N_4226);
and U4481 (N_4481,N_4342,N_4241);
nor U4482 (N_4482,N_4325,N_4239);
or U4483 (N_4483,N_4206,N_4302);
or U4484 (N_4484,N_4211,N_4324);
or U4485 (N_4485,N_4338,N_4217);
or U4486 (N_4486,N_4276,N_4202);
or U4487 (N_4487,N_4329,N_4209);
xnor U4488 (N_4488,N_4203,N_4283);
xnor U4489 (N_4489,N_4208,N_4269);
nand U4490 (N_4490,N_4221,N_4228);
nor U4491 (N_4491,N_4349,N_4340);
or U4492 (N_4492,N_4247,N_4259);
and U4493 (N_4493,N_4329,N_4313);
xnor U4494 (N_4494,N_4240,N_4258);
xor U4495 (N_4495,N_4320,N_4203);
nor U4496 (N_4496,N_4281,N_4232);
or U4497 (N_4497,N_4222,N_4263);
and U4498 (N_4498,N_4202,N_4288);
and U4499 (N_4499,N_4213,N_4303);
nand U4500 (N_4500,N_4423,N_4403);
xor U4501 (N_4501,N_4425,N_4475);
xnor U4502 (N_4502,N_4404,N_4440);
nor U4503 (N_4503,N_4466,N_4456);
nor U4504 (N_4504,N_4476,N_4412);
or U4505 (N_4505,N_4465,N_4426);
xnor U4506 (N_4506,N_4457,N_4387);
or U4507 (N_4507,N_4464,N_4415);
or U4508 (N_4508,N_4385,N_4473);
xnor U4509 (N_4509,N_4356,N_4454);
nand U4510 (N_4510,N_4439,N_4438);
xnor U4511 (N_4511,N_4411,N_4350);
nand U4512 (N_4512,N_4485,N_4398);
and U4513 (N_4513,N_4374,N_4396);
nand U4514 (N_4514,N_4357,N_4389);
nand U4515 (N_4515,N_4352,N_4488);
or U4516 (N_4516,N_4453,N_4397);
and U4517 (N_4517,N_4482,N_4364);
or U4518 (N_4518,N_4468,N_4498);
and U4519 (N_4519,N_4467,N_4495);
or U4520 (N_4520,N_4442,N_4407);
or U4521 (N_4521,N_4359,N_4381);
xor U4522 (N_4522,N_4471,N_4368);
nor U4523 (N_4523,N_4416,N_4420);
nand U4524 (N_4524,N_4490,N_4459);
nor U4525 (N_4525,N_4445,N_4451);
and U4526 (N_4526,N_4379,N_4372);
nor U4527 (N_4527,N_4376,N_4388);
and U4528 (N_4528,N_4401,N_4480);
nor U4529 (N_4529,N_4472,N_4455);
xnor U4530 (N_4530,N_4494,N_4417);
nand U4531 (N_4531,N_4421,N_4484);
or U4532 (N_4532,N_4441,N_4427);
xnor U4533 (N_4533,N_4400,N_4497);
nand U4534 (N_4534,N_4496,N_4499);
nand U4535 (N_4535,N_4463,N_4370);
or U4536 (N_4536,N_4478,N_4431);
nand U4537 (N_4537,N_4386,N_4371);
nand U4538 (N_4538,N_4395,N_4470);
nor U4539 (N_4539,N_4428,N_4491);
or U4540 (N_4540,N_4402,N_4469);
or U4541 (N_4541,N_4361,N_4414);
nor U4542 (N_4542,N_4353,N_4429);
xnor U4543 (N_4543,N_4432,N_4384);
or U4544 (N_4544,N_4436,N_4351);
nor U4545 (N_4545,N_4446,N_4444);
nor U4546 (N_4546,N_4378,N_4481);
nor U4547 (N_4547,N_4479,N_4477);
or U4548 (N_4548,N_4435,N_4377);
xor U4549 (N_4549,N_4354,N_4399);
nand U4550 (N_4550,N_4493,N_4382);
and U4551 (N_4551,N_4369,N_4365);
nand U4552 (N_4552,N_4487,N_4443);
or U4553 (N_4553,N_4433,N_4373);
nand U4554 (N_4554,N_4447,N_4424);
nand U4555 (N_4555,N_4460,N_4358);
xnor U4556 (N_4556,N_4380,N_4452);
nand U4557 (N_4557,N_4458,N_4462);
and U4558 (N_4558,N_4405,N_4422);
or U4559 (N_4559,N_4413,N_4430);
xnor U4560 (N_4560,N_4418,N_4360);
or U4561 (N_4561,N_4390,N_4363);
xnor U4562 (N_4562,N_4448,N_4355);
nor U4563 (N_4563,N_4474,N_4409);
or U4564 (N_4564,N_4437,N_4362);
nand U4565 (N_4565,N_4392,N_4367);
nand U4566 (N_4566,N_4486,N_4492);
xor U4567 (N_4567,N_4410,N_4366);
nand U4568 (N_4568,N_4449,N_4489);
and U4569 (N_4569,N_4383,N_4375);
xnor U4570 (N_4570,N_4450,N_4408);
or U4571 (N_4571,N_4419,N_4393);
nor U4572 (N_4572,N_4461,N_4434);
nand U4573 (N_4573,N_4394,N_4391);
or U4574 (N_4574,N_4483,N_4406);
or U4575 (N_4575,N_4433,N_4366);
nand U4576 (N_4576,N_4447,N_4451);
nand U4577 (N_4577,N_4487,N_4362);
and U4578 (N_4578,N_4452,N_4363);
nand U4579 (N_4579,N_4408,N_4481);
and U4580 (N_4580,N_4431,N_4495);
nand U4581 (N_4581,N_4433,N_4482);
nand U4582 (N_4582,N_4397,N_4468);
xnor U4583 (N_4583,N_4439,N_4445);
nand U4584 (N_4584,N_4472,N_4439);
or U4585 (N_4585,N_4404,N_4369);
and U4586 (N_4586,N_4447,N_4386);
nand U4587 (N_4587,N_4449,N_4372);
xnor U4588 (N_4588,N_4454,N_4385);
and U4589 (N_4589,N_4392,N_4422);
or U4590 (N_4590,N_4381,N_4456);
xor U4591 (N_4591,N_4373,N_4471);
nor U4592 (N_4592,N_4418,N_4416);
or U4593 (N_4593,N_4387,N_4385);
and U4594 (N_4594,N_4481,N_4449);
or U4595 (N_4595,N_4432,N_4364);
xnor U4596 (N_4596,N_4490,N_4386);
nor U4597 (N_4597,N_4378,N_4460);
and U4598 (N_4598,N_4429,N_4450);
nor U4599 (N_4599,N_4411,N_4423);
nand U4600 (N_4600,N_4457,N_4429);
xor U4601 (N_4601,N_4463,N_4361);
nand U4602 (N_4602,N_4401,N_4457);
nor U4603 (N_4603,N_4452,N_4382);
or U4604 (N_4604,N_4407,N_4432);
and U4605 (N_4605,N_4378,N_4490);
and U4606 (N_4606,N_4481,N_4369);
or U4607 (N_4607,N_4407,N_4377);
xor U4608 (N_4608,N_4405,N_4477);
or U4609 (N_4609,N_4382,N_4471);
nand U4610 (N_4610,N_4497,N_4441);
or U4611 (N_4611,N_4376,N_4378);
nor U4612 (N_4612,N_4367,N_4472);
and U4613 (N_4613,N_4406,N_4477);
nand U4614 (N_4614,N_4498,N_4461);
nor U4615 (N_4615,N_4492,N_4399);
and U4616 (N_4616,N_4465,N_4407);
nand U4617 (N_4617,N_4353,N_4411);
xnor U4618 (N_4618,N_4427,N_4472);
nand U4619 (N_4619,N_4392,N_4380);
nand U4620 (N_4620,N_4468,N_4383);
and U4621 (N_4621,N_4430,N_4454);
and U4622 (N_4622,N_4495,N_4377);
nand U4623 (N_4623,N_4409,N_4481);
nor U4624 (N_4624,N_4395,N_4475);
nand U4625 (N_4625,N_4488,N_4421);
nor U4626 (N_4626,N_4456,N_4445);
nor U4627 (N_4627,N_4462,N_4360);
nor U4628 (N_4628,N_4355,N_4473);
nand U4629 (N_4629,N_4466,N_4363);
and U4630 (N_4630,N_4497,N_4455);
and U4631 (N_4631,N_4446,N_4419);
nand U4632 (N_4632,N_4405,N_4462);
and U4633 (N_4633,N_4381,N_4494);
nand U4634 (N_4634,N_4487,N_4369);
or U4635 (N_4635,N_4455,N_4407);
nor U4636 (N_4636,N_4437,N_4364);
xor U4637 (N_4637,N_4461,N_4465);
xnor U4638 (N_4638,N_4483,N_4412);
nor U4639 (N_4639,N_4371,N_4453);
or U4640 (N_4640,N_4368,N_4398);
nor U4641 (N_4641,N_4362,N_4414);
nor U4642 (N_4642,N_4399,N_4441);
nor U4643 (N_4643,N_4498,N_4366);
nor U4644 (N_4644,N_4489,N_4498);
and U4645 (N_4645,N_4379,N_4360);
nand U4646 (N_4646,N_4459,N_4463);
nor U4647 (N_4647,N_4398,N_4456);
and U4648 (N_4648,N_4367,N_4410);
and U4649 (N_4649,N_4467,N_4360);
or U4650 (N_4650,N_4549,N_4559);
xnor U4651 (N_4651,N_4602,N_4529);
and U4652 (N_4652,N_4592,N_4630);
and U4653 (N_4653,N_4532,N_4587);
nand U4654 (N_4654,N_4611,N_4528);
nor U4655 (N_4655,N_4537,N_4627);
nand U4656 (N_4656,N_4535,N_4625);
nor U4657 (N_4657,N_4609,N_4640);
nor U4658 (N_4658,N_4544,N_4567);
xor U4659 (N_4659,N_4578,N_4606);
and U4660 (N_4660,N_4603,N_4631);
nor U4661 (N_4661,N_4585,N_4564);
nor U4662 (N_4662,N_4576,N_4605);
nor U4663 (N_4663,N_4591,N_4548);
nand U4664 (N_4664,N_4616,N_4615);
or U4665 (N_4665,N_4644,N_4522);
and U4666 (N_4666,N_4622,N_4619);
nand U4667 (N_4667,N_4506,N_4612);
nand U4668 (N_4668,N_4600,N_4572);
or U4669 (N_4669,N_4523,N_4573);
nor U4670 (N_4670,N_4524,N_4503);
and U4671 (N_4671,N_4511,N_4604);
and U4672 (N_4672,N_4552,N_4558);
nor U4673 (N_4673,N_4554,N_4596);
xnor U4674 (N_4674,N_4607,N_4513);
xnor U4675 (N_4675,N_4521,N_4595);
and U4676 (N_4676,N_4525,N_4626);
or U4677 (N_4677,N_4530,N_4641);
or U4678 (N_4678,N_4620,N_4647);
or U4679 (N_4679,N_4533,N_4569);
xor U4680 (N_4680,N_4509,N_4527);
nor U4681 (N_4681,N_4624,N_4507);
nand U4682 (N_4682,N_4555,N_4547);
xor U4683 (N_4683,N_4577,N_4565);
nor U4684 (N_4684,N_4556,N_4581);
xnor U4685 (N_4685,N_4515,N_4520);
and U4686 (N_4686,N_4504,N_4629);
nor U4687 (N_4687,N_4599,N_4594);
and U4688 (N_4688,N_4562,N_4613);
nand U4689 (N_4689,N_4571,N_4582);
xor U4690 (N_4690,N_4574,N_4583);
and U4691 (N_4691,N_4517,N_4634);
or U4692 (N_4692,N_4642,N_4531);
and U4693 (N_4693,N_4645,N_4526);
xnor U4694 (N_4694,N_4551,N_4519);
or U4695 (N_4695,N_4621,N_4561);
xnor U4696 (N_4696,N_4638,N_4568);
or U4697 (N_4697,N_4633,N_4586);
and U4698 (N_4698,N_4601,N_4566);
nor U4699 (N_4699,N_4505,N_4648);
or U4700 (N_4700,N_4553,N_4563);
nand U4701 (N_4701,N_4543,N_4632);
and U4702 (N_4702,N_4540,N_4508);
xnor U4703 (N_4703,N_4593,N_4623);
xor U4704 (N_4704,N_4610,N_4510);
and U4705 (N_4705,N_4500,N_4617);
and U4706 (N_4706,N_4628,N_4560);
and U4707 (N_4707,N_4646,N_4534);
nor U4708 (N_4708,N_4637,N_4570);
nand U4709 (N_4709,N_4614,N_4649);
xnor U4710 (N_4710,N_4636,N_4643);
or U4711 (N_4711,N_4588,N_4514);
nor U4712 (N_4712,N_4575,N_4635);
and U4713 (N_4713,N_4502,N_4539);
or U4714 (N_4714,N_4516,N_4518);
nand U4715 (N_4715,N_4501,N_4541);
nand U4716 (N_4716,N_4589,N_4545);
xor U4717 (N_4717,N_4618,N_4598);
nor U4718 (N_4718,N_4597,N_4584);
nand U4719 (N_4719,N_4512,N_4536);
nand U4720 (N_4720,N_4542,N_4579);
nor U4721 (N_4721,N_4590,N_4580);
and U4722 (N_4722,N_4557,N_4538);
and U4723 (N_4723,N_4608,N_4550);
or U4724 (N_4724,N_4639,N_4546);
xnor U4725 (N_4725,N_4520,N_4638);
xor U4726 (N_4726,N_4567,N_4631);
nand U4727 (N_4727,N_4567,N_4578);
nor U4728 (N_4728,N_4608,N_4567);
nor U4729 (N_4729,N_4519,N_4621);
nor U4730 (N_4730,N_4513,N_4604);
nor U4731 (N_4731,N_4618,N_4506);
xnor U4732 (N_4732,N_4568,N_4579);
or U4733 (N_4733,N_4620,N_4631);
nor U4734 (N_4734,N_4504,N_4514);
and U4735 (N_4735,N_4605,N_4608);
xnor U4736 (N_4736,N_4647,N_4587);
xor U4737 (N_4737,N_4503,N_4546);
xor U4738 (N_4738,N_4526,N_4501);
and U4739 (N_4739,N_4633,N_4627);
xor U4740 (N_4740,N_4644,N_4541);
and U4741 (N_4741,N_4557,N_4598);
xor U4742 (N_4742,N_4590,N_4576);
nor U4743 (N_4743,N_4558,N_4630);
nor U4744 (N_4744,N_4513,N_4599);
or U4745 (N_4745,N_4620,N_4543);
xor U4746 (N_4746,N_4502,N_4595);
xor U4747 (N_4747,N_4553,N_4591);
and U4748 (N_4748,N_4586,N_4607);
nor U4749 (N_4749,N_4514,N_4546);
or U4750 (N_4750,N_4579,N_4613);
xor U4751 (N_4751,N_4529,N_4530);
nand U4752 (N_4752,N_4548,N_4619);
and U4753 (N_4753,N_4564,N_4637);
nand U4754 (N_4754,N_4558,N_4574);
xor U4755 (N_4755,N_4582,N_4578);
and U4756 (N_4756,N_4551,N_4500);
xnor U4757 (N_4757,N_4606,N_4640);
nor U4758 (N_4758,N_4644,N_4546);
xor U4759 (N_4759,N_4631,N_4644);
or U4760 (N_4760,N_4534,N_4644);
xnor U4761 (N_4761,N_4583,N_4510);
nor U4762 (N_4762,N_4604,N_4639);
and U4763 (N_4763,N_4509,N_4629);
nor U4764 (N_4764,N_4634,N_4519);
nor U4765 (N_4765,N_4510,N_4578);
or U4766 (N_4766,N_4537,N_4619);
and U4767 (N_4767,N_4546,N_4549);
nand U4768 (N_4768,N_4577,N_4558);
xor U4769 (N_4769,N_4543,N_4585);
nand U4770 (N_4770,N_4601,N_4542);
or U4771 (N_4771,N_4583,N_4611);
nor U4772 (N_4772,N_4545,N_4577);
and U4773 (N_4773,N_4516,N_4641);
nand U4774 (N_4774,N_4565,N_4522);
and U4775 (N_4775,N_4569,N_4626);
or U4776 (N_4776,N_4562,N_4521);
nand U4777 (N_4777,N_4570,N_4641);
and U4778 (N_4778,N_4631,N_4619);
or U4779 (N_4779,N_4541,N_4639);
nand U4780 (N_4780,N_4517,N_4616);
nor U4781 (N_4781,N_4542,N_4596);
xnor U4782 (N_4782,N_4601,N_4577);
nor U4783 (N_4783,N_4617,N_4627);
or U4784 (N_4784,N_4619,N_4644);
and U4785 (N_4785,N_4508,N_4594);
nand U4786 (N_4786,N_4613,N_4611);
or U4787 (N_4787,N_4588,N_4547);
nand U4788 (N_4788,N_4613,N_4551);
or U4789 (N_4789,N_4560,N_4632);
or U4790 (N_4790,N_4542,N_4508);
or U4791 (N_4791,N_4590,N_4633);
and U4792 (N_4792,N_4558,N_4582);
and U4793 (N_4793,N_4649,N_4605);
nand U4794 (N_4794,N_4504,N_4522);
xnor U4795 (N_4795,N_4607,N_4522);
xnor U4796 (N_4796,N_4531,N_4557);
and U4797 (N_4797,N_4570,N_4605);
nor U4798 (N_4798,N_4511,N_4548);
nand U4799 (N_4799,N_4548,N_4571);
xnor U4800 (N_4800,N_4701,N_4731);
or U4801 (N_4801,N_4757,N_4709);
xnor U4802 (N_4802,N_4763,N_4666);
and U4803 (N_4803,N_4768,N_4691);
nand U4804 (N_4804,N_4664,N_4776);
and U4805 (N_4805,N_4675,N_4797);
nor U4806 (N_4806,N_4788,N_4736);
xor U4807 (N_4807,N_4782,N_4704);
nor U4808 (N_4808,N_4762,N_4681);
xor U4809 (N_4809,N_4650,N_4712);
xor U4810 (N_4810,N_4716,N_4655);
or U4811 (N_4811,N_4694,N_4656);
and U4812 (N_4812,N_4761,N_4669);
nand U4813 (N_4813,N_4651,N_4719);
nand U4814 (N_4814,N_4686,N_4737);
nor U4815 (N_4815,N_4660,N_4773);
xnor U4816 (N_4816,N_4705,N_4687);
and U4817 (N_4817,N_4678,N_4685);
and U4818 (N_4818,N_4774,N_4730);
nor U4819 (N_4819,N_4759,N_4676);
xnor U4820 (N_4820,N_4659,N_4787);
xor U4821 (N_4821,N_4696,N_4733);
xnor U4822 (N_4822,N_4785,N_4663);
nand U4823 (N_4823,N_4724,N_4740);
nand U4824 (N_4824,N_4779,N_4789);
xnor U4825 (N_4825,N_4796,N_4795);
and U4826 (N_4826,N_4743,N_4786);
xor U4827 (N_4827,N_4777,N_4784);
or U4828 (N_4828,N_4770,N_4680);
or U4829 (N_4829,N_4707,N_4741);
xor U4830 (N_4830,N_4744,N_4783);
or U4831 (N_4831,N_4749,N_4662);
and U4832 (N_4832,N_4665,N_4673);
nand U4833 (N_4833,N_4729,N_4758);
and U4834 (N_4834,N_4679,N_4799);
nor U4835 (N_4835,N_4671,N_4661);
nand U4836 (N_4836,N_4746,N_4766);
nand U4837 (N_4837,N_4710,N_4748);
and U4838 (N_4838,N_4752,N_4688);
nand U4839 (N_4839,N_4751,N_4711);
or U4840 (N_4840,N_4657,N_4690);
or U4841 (N_4841,N_4738,N_4654);
nand U4842 (N_4842,N_4755,N_4769);
nand U4843 (N_4843,N_4682,N_4765);
nor U4844 (N_4844,N_4683,N_4722);
or U4845 (N_4845,N_4715,N_4697);
and U4846 (N_4846,N_4794,N_4703);
or U4847 (N_4847,N_4745,N_4753);
nor U4848 (N_4848,N_4772,N_4767);
nor U4849 (N_4849,N_4747,N_4653);
and U4850 (N_4850,N_4699,N_4775);
nor U4851 (N_4851,N_4764,N_4677);
nand U4852 (N_4852,N_4798,N_4672);
and U4853 (N_4853,N_4721,N_4780);
or U4854 (N_4854,N_4723,N_4674);
and U4855 (N_4855,N_4706,N_4793);
nor U4856 (N_4856,N_4727,N_4713);
nor U4857 (N_4857,N_4781,N_4725);
nor U4858 (N_4858,N_4790,N_4792);
nor U4859 (N_4859,N_4778,N_4702);
or U4860 (N_4860,N_4728,N_4693);
xor U4861 (N_4861,N_4668,N_4756);
or U4862 (N_4862,N_4742,N_4735);
nand U4863 (N_4863,N_4718,N_4670);
nand U4864 (N_4864,N_4791,N_4695);
or U4865 (N_4865,N_4652,N_4732);
or U4866 (N_4866,N_4734,N_4684);
nor U4867 (N_4867,N_4771,N_4739);
nand U4868 (N_4868,N_4708,N_4698);
xnor U4869 (N_4869,N_4760,N_4754);
and U4870 (N_4870,N_4692,N_4750);
nand U4871 (N_4871,N_4717,N_4689);
xor U4872 (N_4872,N_4658,N_4726);
or U4873 (N_4873,N_4667,N_4714);
xor U4874 (N_4874,N_4700,N_4720);
or U4875 (N_4875,N_4665,N_4773);
or U4876 (N_4876,N_4721,N_4691);
and U4877 (N_4877,N_4736,N_4699);
xnor U4878 (N_4878,N_4782,N_4749);
and U4879 (N_4879,N_4784,N_4685);
nand U4880 (N_4880,N_4798,N_4679);
or U4881 (N_4881,N_4704,N_4734);
and U4882 (N_4882,N_4678,N_4674);
xor U4883 (N_4883,N_4690,N_4758);
nand U4884 (N_4884,N_4679,N_4725);
and U4885 (N_4885,N_4684,N_4730);
nor U4886 (N_4886,N_4718,N_4709);
xnor U4887 (N_4887,N_4780,N_4698);
and U4888 (N_4888,N_4694,N_4696);
or U4889 (N_4889,N_4706,N_4680);
or U4890 (N_4890,N_4696,N_4793);
xor U4891 (N_4891,N_4731,N_4711);
and U4892 (N_4892,N_4763,N_4784);
and U4893 (N_4893,N_4681,N_4723);
or U4894 (N_4894,N_4678,N_4673);
and U4895 (N_4895,N_4676,N_4699);
or U4896 (N_4896,N_4667,N_4656);
nor U4897 (N_4897,N_4743,N_4778);
and U4898 (N_4898,N_4694,N_4780);
and U4899 (N_4899,N_4729,N_4691);
nor U4900 (N_4900,N_4699,N_4793);
or U4901 (N_4901,N_4737,N_4790);
xor U4902 (N_4902,N_4666,N_4688);
xnor U4903 (N_4903,N_4729,N_4650);
nand U4904 (N_4904,N_4768,N_4751);
nand U4905 (N_4905,N_4757,N_4799);
nand U4906 (N_4906,N_4769,N_4664);
nand U4907 (N_4907,N_4794,N_4736);
nor U4908 (N_4908,N_4718,N_4678);
or U4909 (N_4909,N_4798,N_4664);
xor U4910 (N_4910,N_4661,N_4742);
nand U4911 (N_4911,N_4694,N_4684);
and U4912 (N_4912,N_4728,N_4739);
xor U4913 (N_4913,N_4667,N_4704);
and U4914 (N_4914,N_4704,N_4795);
xor U4915 (N_4915,N_4743,N_4673);
or U4916 (N_4916,N_4736,N_4797);
xor U4917 (N_4917,N_4674,N_4721);
xnor U4918 (N_4918,N_4712,N_4688);
nor U4919 (N_4919,N_4745,N_4768);
xnor U4920 (N_4920,N_4657,N_4670);
xnor U4921 (N_4921,N_4726,N_4744);
nor U4922 (N_4922,N_4737,N_4692);
nand U4923 (N_4923,N_4750,N_4734);
nand U4924 (N_4924,N_4689,N_4790);
and U4925 (N_4925,N_4789,N_4718);
xnor U4926 (N_4926,N_4768,N_4775);
nor U4927 (N_4927,N_4788,N_4765);
or U4928 (N_4928,N_4742,N_4654);
and U4929 (N_4929,N_4691,N_4778);
xor U4930 (N_4930,N_4753,N_4663);
xnor U4931 (N_4931,N_4750,N_4682);
or U4932 (N_4932,N_4793,N_4662);
nor U4933 (N_4933,N_4735,N_4754);
nand U4934 (N_4934,N_4790,N_4701);
nand U4935 (N_4935,N_4662,N_4728);
nor U4936 (N_4936,N_4720,N_4779);
xor U4937 (N_4937,N_4697,N_4661);
xor U4938 (N_4938,N_4741,N_4676);
xnor U4939 (N_4939,N_4672,N_4666);
or U4940 (N_4940,N_4659,N_4682);
xnor U4941 (N_4941,N_4777,N_4674);
nor U4942 (N_4942,N_4707,N_4695);
nor U4943 (N_4943,N_4725,N_4662);
nand U4944 (N_4944,N_4728,N_4787);
and U4945 (N_4945,N_4670,N_4753);
nand U4946 (N_4946,N_4782,N_4784);
or U4947 (N_4947,N_4766,N_4719);
nor U4948 (N_4948,N_4791,N_4738);
xnor U4949 (N_4949,N_4713,N_4782);
nand U4950 (N_4950,N_4906,N_4868);
xnor U4951 (N_4951,N_4914,N_4908);
xnor U4952 (N_4952,N_4832,N_4907);
or U4953 (N_4953,N_4836,N_4929);
xor U4954 (N_4954,N_4890,N_4840);
or U4955 (N_4955,N_4851,N_4827);
nor U4956 (N_4956,N_4911,N_4862);
nand U4957 (N_4957,N_4806,N_4826);
and U4958 (N_4958,N_4948,N_4824);
nor U4959 (N_4959,N_4820,N_4899);
xor U4960 (N_4960,N_4835,N_4813);
xnor U4961 (N_4961,N_4807,N_4822);
nor U4962 (N_4962,N_4811,N_4812);
nand U4963 (N_4963,N_4857,N_4858);
and U4964 (N_4964,N_4888,N_4947);
nand U4965 (N_4965,N_4924,N_4876);
or U4966 (N_4966,N_4875,N_4801);
nand U4967 (N_4967,N_4949,N_4918);
nand U4968 (N_4968,N_4828,N_4825);
or U4969 (N_4969,N_4889,N_4864);
xor U4970 (N_4970,N_4933,N_4938);
xor U4971 (N_4971,N_4872,N_4921);
xnor U4972 (N_4972,N_4941,N_4883);
nor U4973 (N_4973,N_4937,N_4839);
nand U4974 (N_4974,N_4861,N_4919);
or U4975 (N_4975,N_4819,N_4946);
and U4976 (N_4976,N_4860,N_4913);
nor U4977 (N_4977,N_4852,N_4939);
nor U4978 (N_4978,N_4844,N_4853);
xnor U4979 (N_4979,N_4847,N_4802);
or U4980 (N_4980,N_4936,N_4800);
or U4981 (N_4981,N_4901,N_4842);
and U4982 (N_4982,N_4894,N_4878);
or U4983 (N_4983,N_4912,N_4896);
nand U4984 (N_4984,N_4900,N_4917);
and U4985 (N_4985,N_4922,N_4885);
or U4986 (N_4986,N_4940,N_4838);
nor U4987 (N_4987,N_4915,N_4815);
or U4988 (N_4988,N_4893,N_4843);
or U4989 (N_4989,N_4923,N_4804);
or U4990 (N_4990,N_4905,N_4910);
nand U4991 (N_4991,N_4866,N_4881);
or U4992 (N_4992,N_4814,N_4897);
nand U4993 (N_4993,N_4867,N_4886);
and U4994 (N_4994,N_4895,N_4871);
xor U4995 (N_4995,N_4920,N_4816);
and U4996 (N_4996,N_4930,N_4849);
nand U4997 (N_4997,N_4805,N_4848);
nand U4998 (N_4998,N_4909,N_4823);
nand U4999 (N_4999,N_4942,N_4903);
xor U5000 (N_5000,N_4877,N_4803);
xnor U5001 (N_5001,N_4928,N_4944);
and U5002 (N_5002,N_4856,N_4880);
nand U5003 (N_5003,N_4869,N_4830);
nor U5004 (N_5004,N_4934,N_4884);
and U5005 (N_5005,N_4925,N_4932);
xor U5006 (N_5006,N_4821,N_4874);
nor U5007 (N_5007,N_4841,N_4898);
nand U5008 (N_5008,N_4891,N_4845);
nor U5009 (N_5009,N_4817,N_4808);
xnor U5010 (N_5010,N_4943,N_4829);
and U5011 (N_5011,N_4837,N_4865);
and U5012 (N_5012,N_4904,N_4850);
and U5013 (N_5013,N_4926,N_4833);
xor U5014 (N_5014,N_4834,N_4892);
nor U5015 (N_5015,N_4931,N_4902);
nor U5016 (N_5016,N_4831,N_4887);
xnor U5017 (N_5017,N_4818,N_4846);
nand U5018 (N_5018,N_4810,N_4882);
nor U5019 (N_5019,N_4859,N_4916);
and U5020 (N_5020,N_4809,N_4870);
or U5021 (N_5021,N_4927,N_4854);
nor U5022 (N_5022,N_4873,N_4855);
nand U5023 (N_5023,N_4863,N_4945);
or U5024 (N_5024,N_4935,N_4879);
or U5025 (N_5025,N_4912,N_4815);
or U5026 (N_5026,N_4856,N_4849);
xor U5027 (N_5027,N_4885,N_4853);
xor U5028 (N_5028,N_4861,N_4894);
or U5029 (N_5029,N_4892,N_4862);
nor U5030 (N_5030,N_4923,N_4861);
or U5031 (N_5031,N_4843,N_4814);
or U5032 (N_5032,N_4862,N_4871);
or U5033 (N_5033,N_4827,N_4857);
nor U5034 (N_5034,N_4861,N_4818);
and U5035 (N_5035,N_4878,N_4840);
or U5036 (N_5036,N_4855,N_4865);
or U5037 (N_5037,N_4948,N_4843);
and U5038 (N_5038,N_4812,N_4855);
nor U5039 (N_5039,N_4848,N_4906);
or U5040 (N_5040,N_4905,N_4805);
nand U5041 (N_5041,N_4900,N_4937);
or U5042 (N_5042,N_4946,N_4808);
or U5043 (N_5043,N_4812,N_4926);
nand U5044 (N_5044,N_4906,N_4819);
xnor U5045 (N_5045,N_4841,N_4877);
nand U5046 (N_5046,N_4931,N_4849);
xnor U5047 (N_5047,N_4907,N_4828);
nor U5048 (N_5048,N_4800,N_4913);
nand U5049 (N_5049,N_4909,N_4879);
xor U5050 (N_5050,N_4885,N_4910);
nor U5051 (N_5051,N_4812,N_4899);
and U5052 (N_5052,N_4868,N_4917);
and U5053 (N_5053,N_4812,N_4846);
xor U5054 (N_5054,N_4899,N_4831);
and U5055 (N_5055,N_4922,N_4867);
nand U5056 (N_5056,N_4831,N_4856);
nor U5057 (N_5057,N_4900,N_4809);
nand U5058 (N_5058,N_4836,N_4911);
nor U5059 (N_5059,N_4814,N_4857);
or U5060 (N_5060,N_4913,N_4899);
and U5061 (N_5061,N_4856,N_4804);
nor U5062 (N_5062,N_4893,N_4944);
nand U5063 (N_5063,N_4944,N_4947);
nor U5064 (N_5064,N_4875,N_4832);
nand U5065 (N_5065,N_4843,N_4934);
and U5066 (N_5066,N_4945,N_4914);
nand U5067 (N_5067,N_4859,N_4863);
xor U5068 (N_5068,N_4867,N_4843);
and U5069 (N_5069,N_4870,N_4927);
nor U5070 (N_5070,N_4883,N_4931);
nor U5071 (N_5071,N_4918,N_4929);
nor U5072 (N_5072,N_4831,N_4881);
and U5073 (N_5073,N_4824,N_4841);
xnor U5074 (N_5074,N_4889,N_4911);
or U5075 (N_5075,N_4863,N_4872);
or U5076 (N_5076,N_4848,N_4926);
or U5077 (N_5077,N_4854,N_4807);
and U5078 (N_5078,N_4916,N_4925);
or U5079 (N_5079,N_4843,N_4863);
xor U5080 (N_5080,N_4926,N_4818);
xnor U5081 (N_5081,N_4879,N_4887);
xor U5082 (N_5082,N_4829,N_4807);
or U5083 (N_5083,N_4872,N_4911);
xor U5084 (N_5084,N_4897,N_4855);
nand U5085 (N_5085,N_4803,N_4943);
and U5086 (N_5086,N_4863,N_4821);
xor U5087 (N_5087,N_4884,N_4820);
nor U5088 (N_5088,N_4885,N_4846);
or U5089 (N_5089,N_4899,N_4858);
nor U5090 (N_5090,N_4876,N_4877);
or U5091 (N_5091,N_4847,N_4800);
xor U5092 (N_5092,N_4819,N_4829);
or U5093 (N_5093,N_4808,N_4935);
nor U5094 (N_5094,N_4879,N_4922);
nand U5095 (N_5095,N_4858,N_4812);
nand U5096 (N_5096,N_4837,N_4943);
or U5097 (N_5097,N_4818,N_4877);
nand U5098 (N_5098,N_4930,N_4847);
nor U5099 (N_5099,N_4922,N_4882);
nand U5100 (N_5100,N_5086,N_5056);
xnor U5101 (N_5101,N_5016,N_5051);
or U5102 (N_5102,N_5006,N_5059);
or U5103 (N_5103,N_5005,N_5065);
or U5104 (N_5104,N_4960,N_5035);
nor U5105 (N_5105,N_5004,N_4984);
nand U5106 (N_5106,N_5045,N_5095);
or U5107 (N_5107,N_5013,N_5094);
nand U5108 (N_5108,N_5057,N_5055);
nor U5109 (N_5109,N_4953,N_4966);
nand U5110 (N_5110,N_4969,N_5096);
xor U5111 (N_5111,N_4983,N_5073);
or U5112 (N_5112,N_5042,N_4979);
nor U5113 (N_5113,N_5080,N_4997);
or U5114 (N_5114,N_4961,N_5010);
nand U5115 (N_5115,N_5058,N_4955);
or U5116 (N_5116,N_5034,N_4971);
and U5117 (N_5117,N_5038,N_5040);
or U5118 (N_5118,N_4991,N_5017);
nand U5119 (N_5119,N_5097,N_5037);
nor U5120 (N_5120,N_4957,N_4964);
nor U5121 (N_5121,N_4959,N_5020);
nand U5122 (N_5122,N_4995,N_5021);
and U5123 (N_5123,N_4951,N_4965);
and U5124 (N_5124,N_5069,N_5041);
or U5125 (N_5125,N_4980,N_4950);
nand U5126 (N_5126,N_4999,N_5075);
xnor U5127 (N_5127,N_4974,N_4994);
xor U5128 (N_5128,N_5018,N_5044);
nor U5129 (N_5129,N_5079,N_4977);
or U5130 (N_5130,N_5071,N_4956);
or U5131 (N_5131,N_5066,N_5036);
or U5132 (N_5132,N_4981,N_4958);
nand U5133 (N_5133,N_4982,N_5008);
nor U5134 (N_5134,N_5091,N_5027);
nand U5135 (N_5135,N_5030,N_4973);
nand U5136 (N_5136,N_5072,N_5046);
nand U5137 (N_5137,N_5026,N_4978);
nor U5138 (N_5138,N_5023,N_5039);
xnor U5139 (N_5139,N_5099,N_5062);
and U5140 (N_5140,N_5019,N_5049);
or U5141 (N_5141,N_4975,N_5084);
nand U5142 (N_5142,N_4963,N_5054);
and U5143 (N_5143,N_5064,N_5015);
nand U5144 (N_5144,N_5050,N_4972);
nor U5145 (N_5145,N_5002,N_4992);
or U5146 (N_5146,N_5060,N_4962);
or U5147 (N_5147,N_5028,N_4993);
and U5148 (N_5148,N_5012,N_5003);
and U5149 (N_5149,N_5067,N_4970);
nand U5150 (N_5150,N_5009,N_5048);
nor U5151 (N_5151,N_5078,N_4985);
xnor U5152 (N_5152,N_5074,N_4967);
nor U5153 (N_5153,N_4952,N_5025);
or U5154 (N_5154,N_5082,N_5088);
nand U5155 (N_5155,N_4989,N_4986);
or U5156 (N_5156,N_5047,N_5001);
nand U5157 (N_5157,N_5032,N_4954);
or U5158 (N_5158,N_5083,N_4998);
xor U5159 (N_5159,N_4990,N_4987);
and U5160 (N_5160,N_5076,N_4996);
or U5161 (N_5161,N_5022,N_5007);
xor U5162 (N_5162,N_5024,N_5029);
and U5163 (N_5163,N_5052,N_5093);
xor U5164 (N_5164,N_4988,N_5081);
or U5165 (N_5165,N_5089,N_5090);
nor U5166 (N_5166,N_5061,N_5068);
nand U5167 (N_5167,N_4976,N_5098);
nand U5168 (N_5168,N_5070,N_5077);
xor U5169 (N_5169,N_5031,N_5011);
nor U5170 (N_5170,N_5063,N_5092);
or U5171 (N_5171,N_4968,N_5000);
and U5172 (N_5172,N_5033,N_5053);
nor U5173 (N_5173,N_5085,N_5014);
nor U5174 (N_5174,N_5043,N_5087);
and U5175 (N_5175,N_5069,N_5084);
and U5176 (N_5176,N_5068,N_5058);
nand U5177 (N_5177,N_5086,N_4972);
xor U5178 (N_5178,N_4960,N_5046);
and U5179 (N_5179,N_4976,N_5061);
and U5180 (N_5180,N_5069,N_5062);
or U5181 (N_5181,N_5019,N_4973);
xor U5182 (N_5182,N_5086,N_4952);
nor U5183 (N_5183,N_5011,N_4982);
nor U5184 (N_5184,N_5013,N_5095);
or U5185 (N_5185,N_4962,N_4951);
xor U5186 (N_5186,N_5040,N_5092);
xnor U5187 (N_5187,N_4973,N_5056);
and U5188 (N_5188,N_4982,N_4972);
nor U5189 (N_5189,N_4969,N_5098);
nand U5190 (N_5190,N_4985,N_5095);
or U5191 (N_5191,N_4967,N_5053);
or U5192 (N_5192,N_4964,N_4971);
or U5193 (N_5193,N_5021,N_4988);
and U5194 (N_5194,N_4990,N_5050);
or U5195 (N_5195,N_5084,N_4998);
or U5196 (N_5196,N_5091,N_5053);
nor U5197 (N_5197,N_5032,N_4985);
nand U5198 (N_5198,N_5081,N_4951);
and U5199 (N_5199,N_5035,N_5052);
nor U5200 (N_5200,N_5038,N_4967);
nor U5201 (N_5201,N_5060,N_4998);
or U5202 (N_5202,N_4994,N_4997);
and U5203 (N_5203,N_5026,N_5067);
nand U5204 (N_5204,N_4953,N_4957);
and U5205 (N_5205,N_5059,N_4989);
and U5206 (N_5206,N_4950,N_4963);
or U5207 (N_5207,N_5057,N_4994);
nand U5208 (N_5208,N_5034,N_4964);
nor U5209 (N_5209,N_5077,N_5029);
nor U5210 (N_5210,N_4965,N_5004);
and U5211 (N_5211,N_5030,N_5099);
or U5212 (N_5212,N_4983,N_5099);
xor U5213 (N_5213,N_4968,N_5047);
or U5214 (N_5214,N_4967,N_4988);
and U5215 (N_5215,N_5076,N_4977);
nand U5216 (N_5216,N_5034,N_5048);
xor U5217 (N_5217,N_4996,N_5055);
nand U5218 (N_5218,N_4982,N_5025);
nor U5219 (N_5219,N_4994,N_4985);
nand U5220 (N_5220,N_4985,N_5074);
and U5221 (N_5221,N_5067,N_5093);
xor U5222 (N_5222,N_4991,N_5029);
or U5223 (N_5223,N_5051,N_5083);
nand U5224 (N_5224,N_4954,N_4963);
nand U5225 (N_5225,N_5006,N_4978);
nand U5226 (N_5226,N_4987,N_5011);
or U5227 (N_5227,N_5094,N_4996);
and U5228 (N_5228,N_5070,N_5023);
nand U5229 (N_5229,N_5023,N_5017);
nand U5230 (N_5230,N_5084,N_5093);
xnor U5231 (N_5231,N_5040,N_4970);
nand U5232 (N_5232,N_5092,N_4977);
nand U5233 (N_5233,N_4982,N_5015);
or U5234 (N_5234,N_4998,N_5053);
nand U5235 (N_5235,N_5059,N_5051);
nand U5236 (N_5236,N_5096,N_4970);
nand U5237 (N_5237,N_5047,N_5021);
nand U5238 (N_5238,N_5064,N_4991);
or U5239 (N_5239,N_4962,N_5072);
xnor U5240 (N_5240,N_5024,N_5016);
nand U5241 (N_5241,N_5008,N_5038);
nand U5242 (N_5242,N_4954,N_5004);
nand U5243 (N_5243,N_4980,N_5066);
and U5244 (N_5244,N_5091,N_5028);
nor U5245 (N_5245,N_5036,N_5093);
or U5246 (N_5246,N_5056,N_5068);
or U5247 (N_5247,N_5095,N_4994);
nand U5248 (N_5248,N_5075,N_4997);
and U5249 (N_5249,N_5010,N_5095);
or U5250 (N_5250,N_5199,N_5230);
or U5251 (N_5251,N_5248,N_5167);
and U5252 (N_5252,N_5165,N_5177);
nand U5253 (N_5253,N_5220,N_5228);
xor U5254 (N_5254,N_5202,N_5178);
nor U5255 (N_5255,N_5210,N_5129);
nor U5256 (N_5256,N_5219,N_5120);
nor U5257 (N_5257,N_5234,N_5192);
nor U5258 (N_5258,N_5214,N_5191);
or U5259 (N_5259,N_5243,N_5138);
xnor U5260 (N_5260,N_5190,N_5217);
or U5261 (N_5261,N_5204,N_5241);
nor U5262 (N_5262,N_5141,N_5121);
and U5263 (N_5263,N_5145,N_5186);
nor U5264 (N_5264,N_5171,N_5126);
nor U5265 (N_5265,N_5139,N_5207);
xnor U5266 (N_5266,N_5169,N_5215);
nand U5267 (N_5267,N_5123,N_5162);
nand U5268 (N_5268,N_5246,N_5156);
nor U5269 (N_5269,N_5137,N_5163);
and U5270 (N_5270,N_5119,N_5221);
nand U5271 (N_5271,N_5107,N_5249);
nor U5272 (N_5272,N_5102,N_5236);
or U5273 (N_5273,N_5122,N_5218);
or U5274 (N_5274,N_5226,N_5200);
nand U5275 (N_5275,N_5131,N_5238);
or U5276 (N_5276,N_5194,N_5147);
xor U5277 (N_5277,N_5112,N_5232);
xor U5278 (N_5278,N_5117,N_5113);
xnor U5279 (N_5279,N_5143,N_5213);
and U5280 (N_5280,N_5240,N_5108);
and U5281 (N_5281,N_5168,N_5231);
xnor U5282 (N_5282,N_5203,N_5109);
xnor U5283 (N_5283,N_5195,N_5105);
nand U5284 (N_5284,N_5198,N_5106);
and U5285 (N_5285,N_5212,N_5227);
xor U5286 (N_5286,N_5128,N_5244);
nor U5287 (N_5287,N_5125,N_5136);
and U5288 (N_5288,N_5134,N_5208);
nand U5289 (N_5289,N_5114,N_5205);
nand U5290 (N_5290,N_5151,N_5211);
and U5291 (N_5291,N_5115,N_5144);
and U5292 (N_5292,N_5116,N_5157);
nor U5293 (N_5293,N_5140,N_5223);
or U5294 (N_5294,N_5142,N_5100);
nor U5295 (N_5295,N_5153,N_5242);
or U5296 (N_5296,N_5216,N_5181);
xnor U5297 (N_5297,N_5237,N_5224);
or U5298 (N_5298,N_5187,N_5146);
nor U5299 (N_5299,N_5164,N_5103);
or U5300 (N_5300,N_5135,N_5201);
xor U5301 (N_5301,N_5189,N_5247);
xor U5302 (N_5302,N_5174,N_5170);
nor U5303 (N_5303,N_5118,N_5111);
or U5304 (N_5304,N_5233,N_5179);
nand U5305 (N_5305,N_5229,N_5188);
xor U5306 (N_5306,N_5196,N_5183);
nand U5307 (N_5307,N_5175,N_5124);
xnor U5308 (N_5308,N_5206,N_5127);
or U5309 (N_5309,N_5197,N_5176);
and U5310 (N_5310,N_5209,N_5158);
and U5311 (N_5311,N_5245,N_5155);
nand U5312 (N_5312,N_5235,N_5225);
or U5313 (N_5313,N_5185,N_5184);
and U5314 (N_5314,N_5166,N_5182);
xnor U5315 (N_5315,N_5161,N_5110);
xor U5316 (N_5316,N_5132,N_5222);
or U5317 (N_5317,N_5180,N_5130);
nor U5318 (N_5318,N_5148,N_5133);
and U5319 (N_5319,N_5159,N_5160);
nor U5320 (N_5320,N_5104,N_5172);
nand U5321 (N_5321,N_5154,N_5101);
xnor U5322 (N_5322,N_5150,N_5152);
xor U5323 (N_5323,N_5193,N_5149);
nand U5324 (N_5324,N_5173,N_5239);
xnor U5325 (N_5325,N_5222,N_5106);
or U5326 (N_5326,N_5241,N_5145);
nor U5327 (N_5327,N_5176,N_5120);
or U5328 (N_5328,N_5101,N_5147);
nand U5329 (N_5329,N_5106,N_5160);
nor U5330 (N_5330,N_5205,N_5230);
nand U5331 (N_5331,N_5206,N_5108);
nor U5332 (N_5332,N_5128,N_5249);
xnor U5333 (N_5333,N_5241,N_5222);
and U5334 (N_5334,N_5181,N_5137);
and U5335 (N_5335,N_5128,N_5223);
nand U5336 (N_5336,N_5211,N_5179);
or U5337 (N_5337,N_5103,N_5232);
or U5338 (N_5338,N_5247,N_5246);
and U5339 (N_5339,N_5193,N_5248);
nand U5340 (N_5340,N_5228,N_5148);
xnor U5341 (N_5341,N_5171,N_5215);
xor U5342 (N_5342,N_5107,N_5168);
nand U5343 (N_5343,N_5224,N_5159);
nor U5344 (N_5344,N_5171,N_5188);
and U5345 (N_5345,N_5233,N_5160);
nand U5346 (N_5346,N_5195,N_5202);
or U5347 (N_5347,N_5186,N_5146);
xor U5348 (N_5348,N_5205,N_5240);
or U5349 (N_5349,N_5236,N_5242);
nor U5350 (N_5350,N_5169,N_5147);
xor U5351 (N_5351,N_5102,N_5241);
nor U5352 (N_5352,N_5161,N_5230);
or U5353 (N_5353,N_5195,N_5203);
or U5354 (N_5354,N_5142,N_5174);
and U5355 (N_5355,N_5135,N_5158);
nand U5356 (N_5356,N_5105,N_5160);
and U5357 (N_5357,N_5217,N_5144);
nor U5358 (N_5358,N_5245,N_5174);
and U5359 (N_5359,N_5189,N_5235);
xnor U5360 (N_5360,N_5118,N_5103);
nor U5361 (N_5361,N_5206,N_5220);
and U5362 (N_5362,N_5235,N_5160);
or U5363 (N_5363,N_5145,N_5174);
and U5364 (N_5364,N_5127,N_5208);
and U5365 (N_5365,N_5108,N_5189);
xnor U5366 (N_5366,N_5176,N_5219);
xor U5367 (N_5367,N_5232,N_5189);
xor U5368 (N_5368,N_5163,N_5219);
nor U5369 (N_5369,N_5125,N_5230);
nor U5370 (N_5370,N_5106,N_5191);
and U5371 (N_5371,N_5128,N_5168);
xnor U5372 (N_5372,N_5148,N_5176);
nand U5373 (N_5373,N_5160,N_5200);
nor U5374 (N_5374,N_5240,N_5128);
xnor U5375 (N_5375,N_5224,N_5148);
and U5376 (N_5376,N_5169,N_5110);
nand U5377 (N_5377,N_5105,N_5135);
and U5378 (N_5378,N_5108,N_5113);
xnor U5379 (N_5379,N_5135,N_5165);
nor U5380 (N_5380,N_5132,N_5197);
and U5381 (N_5381,N_5100,N_5166);
nand U5382 (N_5382,N_5176,N_5195);
and U5383 (N_5383,N_5115,N_5246);
nor U5384 (N_5384,N_5106,N_5248);
nand U5385 (N_5385,N_5228,N_5105);
nand U5386 (N_5386,N_5132,N_5224);
nand U5387 (N_5387,N_5223,N_5202);
nand U5388 (N_5388,N_5194,N_5159);
and U5389 (N_5389,N_5106,N_5204);
xor U5390 (N_5390,N_5221,N_5105);
xor U5391 (N_5391,N_5184,N_5161);
nand U5392 (N_5392,N_5227,N_5161);
or U5393 (N_5393,N_5112,N_5101);
nor U5394 (N_5394,N_5196,N_5112);
nand U5395 (N_5395,N_5102,N_5211);
nor U5396 (N_5396,N_5154,N_5193);
nand U5397 (N_5397,N_5204,N_5188);
xor U5398 (N_5398,N_5190,N_5141);
and U5399 (N_5399,N_5178,N_5183);
nor U5400 (N_5400,N_5368,N_5311);
nor U5401 (N_5401,N_5346,N_5379);
nor U5402 (N_5402,N_5323,N_5293);
nor U5403 (N_5403,N_5253,N_5394);
or U5404 (N_5404,N_5329,N_5334);
nand U5405 (N_5405,N_5288,N_5302);
nand U5406 (N_5406,N_5287,N_5292);
nor U5407 (N_5407,N_5355,N_5380);
and U5408 (N_5408,N_5252,N_5307);
and U5409 (N_5409,N_5377,N_5277);
xor U5410 (N_5410,N_5396,N_5331);
and U5411 (N_5411,N_5382,N_5359);
xnor U5412 (N_5412,N_5298,N_5306);
and U5413 (N_5413,N_5308,N_5260);
xor U5414 (N_5414,N_5319,N_5291);
and U5415 (N_5415,N_5270,N_5317);
nand U5416 (N_5416,N_5274,N_5272);
nor U5417 (N_5417,N_5374,N_5336);
xnor U5418 (N_5418,N_5387,N_5314);
nor U5419 (N_5419,N_5313,N_5367);
or U5420 (N_5420,N_5285,N_5344);
and U5421 (N_5421,N_5339,N_5326);
and U5422 (N_5422,N_5266,N_5262);
xor U5423 (N_5423,N_5385,N_5320);
nor U5424 (N_5424,N_5349,N_5263);
nor U5425 (N_5425,N_5257,N_5353);
nor U5426 (N_5426,N_5254,N_5269);
or U5427 (N_5427,N_5347,N_5351);
or U5428 (N_5428,N_5304,N_5310);
nand U5429 (N_5429,N_5350,N_5341);
or U5430 (N_5430,N_5395,N_5279);
nand U5431 (N_5431,N_5392,N_5381);
nor U5432 (N_5432,N_5390,N_5259);
xnor U5433 (N_5433,N_5267,N_5316);
nor U5434 (N_5434,N_5386,N_5264);
nand U5435 (N_5435,N_5305,N_5335);
xor U5436 (N_5436,N_5332,N_5297);
nand U5437 (N_5437,N_5278,N_5399);
and U5438 (N_5438,N_5373,N_5398);
or U5439 (N_5439,N_5333,N_5256);
or U5440 (N_5440,N_5251,N_5384);
and U5441 (N_5441,N_5343,N_5275);
nor U5442 (N_5442,N_5363,N_5301);
and U5443 (N_5443,N_5327,N_5337);
and U5444 (N_5444,N_5325,N_5276);
nand U5445 (N_5445,N_5318,N_5361);
and U5446 (N_5446,N_5356,N_5295);
nor U5447 (N_5447,N_5255,N_5338);
or U5448 (N_5448,N_5354,N_5383);
and U5449 (N_5449,N_5360,N_5324);
nand U5450 (N_5450,N_5328,N_5300);
xor U5451 (N_5451,N_5261,N_5294);
nand U5452 (N_5452,N_5364,N_5258);
nor U5453 (N_5453,N_5345,N_5342);
or U5454 (N_5454,N_5369,N_5282);
nand U5455 (N_5455,N_5370,N_5340);
or U5456 (N_5456,N_5366,N_5352);
xnor U5457 (N_5457,N_5286,N_5271);
xnor U5458 (N_5458,N_5388,N_5322);
xor U5459 (N_5459,N_5281,N_5296);
nand U5460 (N_5460,N_5362,N_5393);
nor U5461 (N_5461,N_5315,N_5365);
nand U5462 (N_5462,N_5273,N_5250);
xor U5463 (N_5463,N_5376,N_5397);
and U5464 (N_5464,N_5321,N_5309);
or U5465 (N_5465,N_5303,N_5289);
nor U5466 (N_5466,N_5358,N_5312);
xor U5467 (N_5467,N_5284,N_5372);
nor U5468 (N_5468,N_5389,N_5290);
nor U5469 (N_5469,N_5268,N_5357);
nand U5470 (N_5470,N_5283,N_5299);
xnor U5471 (N_5471,N_5348,N_5280);
nand U5472 (N_5472,N_5371,N_5265);
and U5473 (N_5473,N_5375,N_5391);
nand U5474 (N_5474,N_5378,N_5330);
nand U5475 (N_5475,N_5275,N_5261);
and U5476 (N_5476,N_5293,N_5388);
nand U5477 (N_5477,N_5274,N_5336);
xor U5478 (N_5478,N_5388,N_5267);
xor U5479 (N_5479,N_5307,N_5271);
nor U5480 (N_5480,N_5343,N_5269);
nand U5481 (N_5481,N_5304,N_5377);
xnor U5482 (N_5482,N_5323,N_5346);
xor U5483 (N_5483,N_5264,N_5314);
nand U5484 (N_5484,N_5385,N_5278);
nor U5485 (N_5485,N_5333,N_5299);
or U5486 (N_5486,N_5365,N_5333);
nor U5487 (N_5487,N_5358,N_5317);
and U5488 (N_5488,N_5311,N_5290);
xnor U5489 (N_5489,N_5308,N_5338);
nor U5490 (N_5490,N_5389,N_5343);
nand U5491 (N_5491,N_5313,N_5349);
and U5492 (N_5492,N_5389,N_5284);
nor U5493 (N_5493,N_5268,N_5366);
or U5494 (N_5494,N_5336,N_5348);
or U5495 (N_5495,N_5394,N_5334);
or U5496 (N_5496,N_5304,N_5339);
nor U5497 (N_5497,N_5379,N_5323);
nor U5498 (N_5498,N_5257,N_5390);
nor U5499 (N_5499,N_5353,N_5332);
nor U5500 (N_5500,N_5377,N_5278);
or U5501 (N_5501,N_5369,N_5328);
nand U5502 (N_5502,N_5279,N_5274);
xor U5503 (N_5503,N_5297,N_5330);
and U5504 (N_5504,N_5349,N_5256);
nand U5505 (N_5505,N_5342,N_5371);
nor U5506 (N_5506,N_5368,N_5343);
xnor U5507 (N_5507,N_5309,N_5329);
nor U5508 (N_5508,N_5376,N_5283);
nand U5509 (N_5509,N_5266,N_5349);
and U5510 (N_5510,N_5375,N_5300);
xor U5511 (N_5511,N_5266,N_5319);
nand U5512 (N_5512,N_5296,N_5377);
and U5513 (N_5513,N_5330,N_5261);
nor U5514 (N_5514,N_5295,N_5326);
xnor U5515 (N_5515,N_5357,N_5313);
nand U5516 (N_5516,N_5341,N_5264);
xnor U5517 (N_5517,N_5287,N_5324);
xor U5518 (N_5518,N_5338,N_5318);
or U5519 (N_5519,N_5397,N_5321);
and U5520 (N_5520,N_5335,N_5313);
or U5521 (N_5521,N_5305,N_5276);
xnor U5522 (N_5522,N_5295,N_5388);
xor U5523 (N_5523,N_5252,N_5305);
nand U5524 (N_5524,N_5399,N_5264);
and U5525 (N_5525,N_5264,N_5321);
nor U5526 (N_5526,N_5344,N_5364);
and U5527 (N_5527,N_5332,N_5291);
nand U5528 (N_5528,N_5290,N_5368);
and U5529 (N_5529,N_5375,N_5255);
or U5530 (N_5530,N_5294,N_5370);
or U5531 (N_5531,N_5334,N_5348);
nor U5532 (N_5532,N_5309,N_5393);
xor U5533 (N_5533,N_5386,N_5351);
xor U5534 (N_5534,N_5291,N_5327);
or U5535 (N_5535,N_5311,N_5273);
nand U5536 (N_5536,N_5381,N_5274);
or U5537 (N_5537,N_5378,N_5352);
nand U5538 (N_5538,N_5268,N_5261);
xnor U5539 (N_5539,N_5329,N_5312);
nor U5540 (N_5540,N_5344,N_5257);
nor U5541 (N_5541,N_5298,N_5283);
xnor U5542 (N_5542,N_5326,N_5366);
nor U5543 (N_5543,N_5361,N_5367);
nand U5544 (N_5544,N_5346,N_5304);
and U5545 (N_5545,N_5365,N_5287);
xnor U5546 (N_5546,N_5298,N_5337);
or U5547 (N_5547,N_5268,N_5358);
or U5548 (N_5548,N_5347,N_5381);
xor U5549 (N_5549,N_5359,N_5365);
xor U5550 (N_5550,N_5404,N_5437);
or U5551 (N_5551,N_5426,N_5467);
xnor U5552 (N_5552,N_5420,N_5504);
and U5553 (N_5553,N_5535,N_5466);
or U5554 (N_5554,N_5516,N_5548);
or U5555 (N_5555,N_5501,N_5459);
xnor U5556 (N_5556,N_5545,N_5472);
or U5557 (N_5557,N_5497,N_5529);
nor U5558 (N_5558,N_5452,N_5489);
nand U5559 (N_5559,N_5433,N_5511);
nor U5560 (N_5560,N_5430,N_5498);
or U5561 (N_5561,N_5485,N_5520);
nand U5562 (N_5562,N_5454,N_5522);
xnor U5563 (N_5563,N_5468,N_5428);
and U5564 (N_5564,N_5491,N_5479);
nor U5565 (N_5565,N_5542,N_5407);
nand U5566 (N_5566,N_5425,N_5546);
or U5567 (N_5567,N_5465,N_5443);
or U5568 (N_5568,N_5400,N_5444);
nor U5569 (N_5569,N_5534,N_5533);
xor U5570 (N_5570,N_5528,N_5402);
nor U5571 (N_5571,N_5471,N_5507);
or U5572 (N_5572,N_5494,N_5499);
nor U5573 (N_5573,N_5447,N_5457);
and U5574 (N_5574,N_5495,N_5416);
xor U5575 (N_5575,N_5417,N_5469);
or U5576 (N_5576,N_5502,N_5448);
nor U5577 (N_5577,N_5441,N_5487);
xor U5578 (N_5578,N_5475,N_5438);
or U5579 (N_5579,N_5531,N_5427);
xnor U5580 (N_5580,N_5532,N_5521);
and U5581 (N_5581,N_5523,N_5509);
nor U5582 (N_5582,N_5496,N_5414);
nand U5583 (N_5583,N_5429,N_5519);
or U5584 (N_5584,N_5483,N_5524);
and U5585 (N_5585,N_5537,N_5474);
xnor U5586 (N_5586,N_5462,N_5405);
nand U5587 (N_5587,N_5412,N_5431);
or U5588 (N_5588,N_5484,N_5526);
and U5589 (N_5589,N_5423,N_5421);
and U5590 (N_5590,N_5541,N_5451);
xnor U5591 (N_5591,N_5492,N_5403);
and U5592 (N_5592,N_5445,N_5488);
nor U5593 (N_5593,N_5482,N_5538);
nand U5594 (N_5594,N_5406,N_5470);
nor U5595 (N_5595,N_5476,N_5508);
xor U5596 (N_5596,N_5439,N_5486);
nand U5597 (N_5597,N_5456,N_5446);
nand U5598 (N_5598,N_5422,N_5413);
xnor U5599 (N_5599,N_5503,N_5539);
or U5600 (N_5600,N_5549,N_5518);
nand U5601 (N_5601,N_5408,N_5432);
or U5602 (N_5602,N_5514,N_5510);
nor U5603 (N_5603,N_5540,N_5424);
nand U5604 (N_5604,N_5460,N_5506);
nand U5605 (N_5605,N_5464,N_5473);
and U5606 (N_5606,N_5415,N_5442);
nand U5607 (N_5607,N_5513,N_5458);
and U5608 (N_5608,N_5536,N_5453);
and U5609 (N_5609,N_5434,N_5478);
xor U5610 (N_5610,N_5547,N_5517);
xor U5611 (N_5611,N_5461,N_5512);
and U5612 (N_5612,N_5505,N_5500);
xnor U5613 (N_5613,N_5449,N_5410);
nand U5614 (N_5614,N_5418,N_5440);
xor U5615 (N_5615,N_5435,N_5477);
nand U5616 (N_5616,N_5419,N_5527);
nor U5617 (N_5617,N_5515,N_5525);
and U5618 (N_5618,N_5490,N_5530);
xor U5619 (N_5619,N_5480,N_5450);
or U5620 (N_5620,N_5463,N_5455);
or U5621 (N_5621,N_5411,N_5543);
xor U5622 (N_5622,N_5481,N_5544);
xor U5623 (N_5623,N_5401,N_5436);
or U5624 (N_5624,N_5409,N_5493);
xor U5625 (N_5625,N_5456,N_5401);
nor U5626 (N_5626,N_5515,N_5530);
nor U5627 (N_5627,N_5511,N_5542);
nor U5628 (N_5628,N_5407,N_5549);
or U5629 (N_5629,N_5476,N_5547);
xor U5630 (N_5630,N_5433,N_5481);
nor U5631 (N_5631,N_5473,N_5516);
and U5632 (N_5632,N_5438,N_5504);
xor U5633 (N_5633,N_5528,N_5467);
nor U5634 (N_5634,N_5511,N_5515);
nor U5635 (N_5635,N_5492,N_5462);
xor U5636 (N_5636,N_5508,N_5415);
and U5637 (N_5637,N_5545,N_5435);
or U5638 (N_5638,N_5446,N_5452);
xor U5639 (N_5639,N_5523,N_5451);
nor U5640 (N_5640,N_5465,N_5474);
and U5641 (N_5641,N_5460,N_5547);
xnor U5642 (N_5642,N_5518,N_5418);
or U5643 (N_5643,N_5425,N_5404);
or U5644 (N_5644,N_5525,N_5491);
and U5645 (N_5645,N_5403,N_5439);
xnor U5646 (N_5646,N_5421,N_5407);
xnor U5647 (N_5647,N_5494,N_5501);
or U5648 (N_5648,N_5543,N_5478);
and U5649 (N_5649,N_5432,N_5519);
or U5650 (N_5650,N_5433,N_5464);
and U5651 (N_5651,N_5514,N_5453);
and U5652 (N_5652,N_5545,N_5429);
and U5653 (N_5653,N_5484,N_5543);
nor U5654 (N_5654,N_5542,N_5494);
xnor U5655 (N_5655,N_5456,N_5437);
xnor U5656 (N_5656,N_5432,N_5424);
xor U5657 (N_5657,N_5432,N_5401);
and U5658 (N_5658,N_5412,N_5488);
nor U5659 (N_5659,N_5454,N_5466);
and U5660 (N_5660,N_5467,N_5465);
or U5661 (N_5661,N_5412,N_5497);
or U5662 (N_5662,N_5488,N_5476);
nor U5663 (N_5663,N_5442,N_5486);
and U5664 (N_5664,N_5467,N_5418);
and U5665 (N_5665,N_5410,N_5408);
or U5666 (N_5666,N_5465,N_5491);
xor U5667 (N_5667,N_5527,N_5416);
nor U5668 (N_5668,N_5480,N_5506);
nand U5669 (N_5669,N_5498,N_5544);
xor U5670 (N_5670,N_5434,N_5465);
and U5671 (N_5671,N_5531,N_5441);
xor U5672 (N_5672,N_5456,N_5420);
and U5673 (N_5673,N_5512,N_5513);
xnor U5674 (N_5674,N_5517,N_5518);
or U5675 (N_5675,N_5510,N_5520);
nor U5676 (N_5676,N_5502,N_5514);
and U5677 (N_5677,N_5528,N_5469);
nor U5678 (N_5678,N_5531,N_5435);
xor U5679 (N_5679,N_5432,N_5465);
nor U5680 (N_5680,N_5511,N_5532);
xnor U5681 (N_5681,N_5540,N_5486);
and U5682 (N_5682,N_5463,N_5412);
nor U5683 (N_5683,N_5529,N_5487);
or U5684 (N_5684,N_5460,N_5514);
and U5685 (N_5685,N_5402,N_5420);
nand U5686 (N_5686,N_5471,N_5539);
or U5687 (N_5687,N_5537,N_5455);
xnor U5688 (N_5688,N_5401,N_5511);
nor U5689 (N_5689,N_5447,N_5408);
nand U5690 (N_5690,N_5528,N_5511);
or U5691 (N_5691,N_5402,N_5453);
or U5692 (N_5692,N_5489,N_5532);
nor U5693 (N_5693,N_5542,N_5505);
or U5694 (N_5694,N_5493,N_5426);
nand U5695 (N_5695,N_5445,N_5401);
nor U5696 (N_5696,N_5423,N_5533);
and U5697 (N_5697,N_5486,N_5458);
nand U5698 (N_5698,N_5443,N_5512);
nand U5699 (N_5699,N_5495,N_5423);
nor U5700 (N_5700,N_5636,N_5557);
nor U5701 (N_5701,N_5654,N_5653);
or U5702 (N_5702,N_5590,N_5660);
nor U5703 (N_5703,N_5553,N_5638);
and U5704 (N_5704,N_5678,N_5652);
xor U5705 (N_5705,N_5642,N_5657);
and U5706 (N_5706,N_5576,N_5601);
nor U5707 (N_5707,N_5610,N_5697);
or U5708 (N_5708,N_5551,N_5552);
nor U5709 (N_5709,N_5687,N_5569);
and U5710 (N_5710,N_5618,N_5677);
and U5711 (N_5711,N_5635,N_5641);
nand U5712 (N_5712,N_5662,N_5570);
nand U5713 (N_5713,N_5615,N_5628);
xor U5714 (N_5714,N_5632,N_5575);
and U5715 (N_5715,N_5682,N_5579);
nor U5716 (N_5716,N_5693,N_5679);
nor U5717 (N_5717,N_5622,N_5661);
nand U5718 (N_5718,N_5656,N_5559);
nand U5719 (N_5719,N_5604,N_5668);
or U5720 (N_5720,N_5694,N_5597);
or U5721 (N_5721,N_5586,N_5587);
nor U5722 (N_5722,N_5568,N_5621);
nor U5723 (N_5723,N_5633,N_5592);
nor U5724 (N_5724,N_5648,N_5550);
nand U5725 (N_5725,N_5627,N_5696);
or U5726 (N_5726,N_5602,N_5616);
xor U5727 (N_5727,N_5598,N_5573);
nor U5728 (N_5728,N_5629,N_5680);
nor U5729 (N_5729,N_5623,N_5688);
or U5730 (N_5730,N_5686,N_5650);
nand U5731 (N_5731,N_5625,N_5617);
or U5732 (N_5732,N_5663,N_5584);
or U5733 (N_5733,N_5673,N_5565);
nor U5734 (N_5734,N_5619,N_5631);
and U5735 (N_5735,N_5643,N_5611);
nor U5736 (N_5736,N_5594,N_5560);
and U5737 (N_5737,N_5646,N_5585);
and U5738 (N_5738,N_5609,N_5591);
nand U5739 (N_5739,N_5644,N_5578);
nor U5740 (N_5740,N_5556,N_5670);
nor U5741 (N_5741,N_5608,N_5667);
nand U5742 (N_5742,N_5689,N_5666);
xnor U5743 (N_5743,N_5658,N_5567);
and U5744 (N_5744,N_5675,N_5589);
or U5745 (N_5745,N_5674,N_5593);
or U5746 (N_5746,N_5685,N_5669);
and U5747 (N_5747,N_5620,N_5683);
nand U5748 (N_5748,N_5690,N_5665);
nor U5749 (N_5749,N_5574,N_5672);
or U5750 (N_5750,N_5613,N_5558);
xnor U5751 (N_5751,N_5564,N_5637);
nand U5752 (N_5752,N_5595,N_5695);
and U5753 (N_5753,N_5692,N_5624);
xor U5754 (N_5754,N_5659,N_5582);
or U5755 (N_5755,N_5651,N_5698);
xor U5756 (N_5756,N_5634,N_5612);
or U5757 (N_5757,N_5681,N_5607);
and U5758 (N_5758,N_5647,N_5649);
nor U5759 (N_5759,N_5596,N_5655);
nor U5760 (N_5760,N_5561,N_5566);
nor U5761 (N_5761,N_5645,N_5699);
nand U5762 (N_5762,N_5664,N_5554);
nor U5763 (N_5763,N_5555,N_5684);
and U5764 (N_5764,N_5577,N_5572);
xor U5765 (N_5765,N_5583,N_5563);
nor U5766 (N_5766,N_5614,N_5600);
nand U5767 (N_5767,N_5605,N_5562);
and U5768 (N_5768,N_5606,N_5630);
nand U5769 (N_5769,N_5599,N_5626);
and U5770 (N_5770,N_5580,N_5603);
and U5771 (N_5771,N_5588,N_5640);
nand U5772 (N_5772,N_5581,N_5676);
and U5773 (N_5773,N_5691,N_5671);
nand U5774 (N_5774,N_5571,N_5639);
nand U5775 (N_5775,N_5570,N_5601);
nand U5776 (N_5776,N_5608,N_5575);
nand U5777 (N_5777,N_5670,N_5631);
and U5778 (N_5778,N_5669,N_5640);
nand U5779 (N_5779,N_5618,N_5631);
and U5780 (N_5780,N_5683,N_5578);
or U5781 (N_5781,N_5611,N_5638);
or U5782 (N_5782,N_5654,N_5648);
and U5783 (N_5783,N_5602,N_5686);
xor U5784 (N_5784,N_5586,N_5602);
nor U5785 (N_5785,N_5550,N_5586);
nand U5786 (N_5786,N_5573,N_5672);
nor U5787 (N_5787,N_5633,N_5656);
or U5788 (N_5788,N_5619,N_5642);
and U5789 (N_5789,N_5657,N_5676);
nand U5790 (N_5790,N_5622,N_5569);
and U5791 (N_5791,N_5675,N_5593);
or U5792 (N_5792,N_5680,N_5635);
and U5793 (N_5793,N_5557,N_5574);
xnor U5794 (N_5794,N_5604,N_5588);
xnor U5795 (N_5795,N_5583,N_5635);
nor U5796 (N_5796,N_5628,N_5683);
and U5797 (N_5797,N_5622,N_5552);
and U5798 (N_5798,N_5564,N_5597);
nand U5799 (N_5799,N_5604,N_5597);
or U5800 (N_5800,N_5610,N_5696);
nand U5801 (N_5801,N_5699,N_5618);
nand U5802 (N_5802,N_5632,N_5576);
nor U5803 (N_5803,N_5603,N_5578);
xnor U5804 (N_5804,N_5568,N_5684);
nand U5805 (N_5805,N_5614,N_5635);
xnor U5806 (N_5806,N_5597,N_5689);
nor U5807 (N_5807,N_5648,N_5697);
and U5808 (N_5808,N_5617,N_5634);
xor U5809 (N_5809,N_5654,N_5638);
nor U5810 (N_5810,N_5570,N_5602);
nand U5811 (N_5811,N_5659,N_5591);
and U5812 (N_5812,N_5698,N_5674);
and U5813 (N_5813,N_5660,N_5605);
xnor U5814 (N_5814,N_5577,N_5555);
xor U5815 (N_5815,N_5679,N_5647);
or U5816 (N_5816,N_5620,N_5557);
or U5817 (N_5817,N_5553,N_5609);
nand U5818 (N_5818,N_5635,N_5593);
nor U5819 (N_5819,N_5684,N_5575);
nand U5820 (N_5820,N_5610,N_5588);
nand U5821 (N_5821,N_5672,N_5591);
or U5822 (N_5822,N_5691,N_5656);
nor U5823 (N_5823,N_5648,N_5568);
xnor U5824 (N_5824,N_5584,N_5695);
or U5825 (N_5825,N_5693,N_5572);
xor U5826 (N_5826,N_5611,N_5655);
nand U5827 (N_5827,N_5673,N_5613);
nand U5828 (N_5828,N_5601,N_5692);
xor U5829 (N_5829,N_5689,N_5684);
xnor U5830 (N_5830,N_5594,N_5587);
nor U5831 (N_5831,N_5659,N_5697);
nor U5832 (N_5832,N_5587,N_5563);
nor U5833 (N_5833,N_5581,N_5592);
or U5834 (N_5834,N_5633,N_5631);
or U5835 (N_5835,N_5622,N_5685);
or U5836 (N_5836,N_5556,N_5684);
or U5837 (N_5837,N_5670,N_5635);
or U5838 (N_5838,N_5672,N_5637);
xnor U5839 (N_5839,N_5673,N_5559);
xor U5840 (N_5840,N_5569,N_5570);
nand U5841 (N_5841,N_5567,N_5629);
nor U5842 (N_5842,N_5586,N_5679);
xnor U5843 (N_5843,N_5611,N_5690);
or U5844 (N_5844,N_5561,N_5638);
nor U5845 (N_5845,N_5569,N_5579);
or U5846 (N_5846,N_5605,N_5559);
nand U5847 (N_5847,N_5576,N_5667);
nor U5848 (N_5848,N_5661,N_5677);
and U5849 (N_5849,N_5625,N_5635);
nand U5850 (N_5850,N_5795,N_5786);
nor U5851 (N_5851,N_5802,N_5775);
nor U5852 (N_5852,N_5796,N_5709);
or U5853 (N_5853,N_5793,N_5732);
xor U5854 (N_5854,N_5720,N_5794);
and U5855 (N_5855,N_5797,N_5784);
xor U5856 (N_5856,N_5764,N_5754);
and U5857 (N_5857,N_5808,N_5715);
and U5858 (N_5858,N_5774,N_5813);
and U5859 (N_5859,N_5789,N_5783);
or U5860 (N_5860,N_5822,N_5842);
xnor U5861 (N_5861,N_5701,N_5736);
xnor U5862 (N_5862,N_5766,N_5829);
nor U5863 (N_5863,N_5758,N_5848);
nor U5864 (N_5864,N_5717,N_5777);
and U5865 (N_5865,N_5751,N_5835);
xnor U5866 (N_5866,N_5748,N_5757);
xnor U5867 (N_5867,N_5846,N_5725);
nand U5868 (N_5868,N_5716,N_5756);
nor U5869 (N_5869,N_5713,N_5750);
and U5870 (N_5870,N_5727,N_5812);
and U5871 (N_5871,N_5839,N_5710);
or U5872 (N_5872,N_5801,N_5838);
nand U5873 (N_5873,N_5847,N_5707);
nor U5874 (N_5874,N_5824,N_5714);
nor U5875 (N_5875,N_5738,N_5849);
or U5876 (N_5876,N_5830,N_5826);
nand U5877 (N_5877,N_5763,N_5765);
or U5878 (N_5878,N_5724,N_5825);
and U5879 (N_5879,N_5792,N_5810);
or U5880 (N_5880,N_5843,N_5739);
nor U5881 (N_5881,N_5749,N_5760);
xor U5882 (N_5882,N_5700,N_5799);
nand U5883 (N_5883,N_5819,N_5704);
nand U5884 (N_5884,N_5840,N_5805);
or U5885 (N_5885,N_5818,N_5809);
nor U5886 (N_5886,N_5800,N_5778);
nand U5887 (N_5887,N_5817,N_5771);
nand U5888 (N_5888,N_5806,N_5844);
nor U5889 (N_5889,N_5723,N_5726);
or U5890 (N_5890,N_5761,N_5769);
and U5891 (N_5891,N_5820,N_5711);
nand U5892 (N_5892,N_5781,N_5816);
nor U5893 (N_5893,N_5823,N_5737);
and U5894 (N_5894,N_5755,N_5752);
nand U5895 (N_5895,N_5811,N_5705);
xnor U5896 (N_5896,N_5743,N_5744);
nand U5897 (N_5897,N_5828,N_5773);
nor U5898 (N_5898,N_5719,N_5815);
or U5899 (N_5899,N_5814,N_5706);
nor U5900 (N_5900,N_5722,N_5772);
xnor U5901 (N_5901,N_5746,N_5788);
or U5902 (N_5902,N_5735,N_5845);
nand U5903 (N_5903,N_5834,N_5770);
nor U5904 (N_5904,N_5729,N_5827);
nor U5905 (N_5905,N_5745,N_5741);
nor U5906 (N_5906,N_5836,N_5831);
and U5907 (N_5907,N_5821,N_5731);
xnor U5908 (N_5908,N_5742,N_5804);
or U5909 (N_5909,N_5782,N_5733);
and U5910 (N_5910,N_5798,N_5747);
nor U5911 (N_5911,N_5734,N_5702);
nand U5912 (N_5912,N_5728,N_5785);
nor U5913 (N_5913,N_5779,N_5759);
xnor U5914 (N_5914,N_5776,N_5833);
and U5915 (N_5915,N_5708,N_5841);
nand U5916 (N_5916,N_5837,N_5740);
and U5917 (N_5917,N_5832,N_5807);
and U5918 (N_5918,N_5703,N_5787);
xnor U5919 (N_5919,N_5767,N_5730);
xor U5920 (N_5920,N_5712,N_5803);
nor U5921 (N_5921,N_5780,N_5753);
or U5922 (N_5922,N_5721,N_5762);
nor U5923 (N_5923,N_5790,N_5768);
nand U5924 (N_5924,N_5718,N_5791);
or U5925 (N_5925,N_5725,N_5712);
or U5926 (N_5926,N_5819,N_5787);
xor U5927 (N_5927,N_5813,N_5843);
and U5928 (N_5928,N_5736,N_5792);
nor U5929 (N_5929,N_5773,N_5710);
and U5930 (N_5930,N_5830,N_5772);
nor U5931 (N_5931,N_5831,N_5813);
nor U5932 (N_5932,N_5802,N_5844);
nor U5933 (N_5933,N_5802,N_5744);
nand U5934 (N_5934,N_5787,N_5815);
or U5935 (N_5935,N_5769,N_5798);
and U5936 (N_5936,N_5786,N_5805);
and U5937 (N_5937,N_5767,N_5775);
or U5938 (N_5938,N_5849,N_5823);
and U5939 (N_5939,N_5732,N_5780);
nor U5940 (N_5940,N_5832,N_5703);
or U5941 (N_5941,N_5732,N_5798);
and U5942 (N_5942,N_5843,N_5832);
and U5943 (N_5943,N_5764,N_5839);
and U5944 (N_5944,N_5740,N_5847);
nor U5945 (N_5945,N_5722,N_5794);
nor U5946 (N_5946,N_5743,N_5722);
and U5947 (N_5947,N_5782,N_5813);
or U5948 (N_5948,N_5808,N_5701);
xnor U5949 (N_5949,N_5835,N_5747);
nand U5950 (N_5950,N_5731,N_5712);
xnor U5951 (N_5951,N_5737,N_5785);
xnor U5952 (N_5952,N_5840,N_5770);
xnor U5953 (N_5953,N_5700,N_5788);
or U5954 (N_5954,N_5777,N_5739);
xor U5955 (N_5955,N_5716,N_5844);
xnor U5956 (N_5956,N_5804,N_5832);
nor U5957 (N_5957,N_5820,N_5745);
xor U5958 (N_5958,N_5765,N_5736);
nand U5959 (N_5959,N_5729,N_5821);
nand U5960 (N_5960,N_5848,N_5739);
and U5961 (N_5961,N_5817,N_5810);
nand U5962 (N_5962,N_5783,N_5753);
nand U5963 (N_5963,N_5818,N_5787);
xor U5964 (N_5964,N_5742,N_5710);
or U5965 (N_5965,N_5767,N_5707);
or U5966 (N_5966,N_5827,N_5785);
xnor U5967 (N_5967,N_5729,N_5791);
xnor U5968 (N_5968,N_5807,N_5721);
xor U5969 (N_5969,N_5745,N_5797);
and U5970 (N_5970,N_5804,N_5727);
xor U5971 (N_5971,N_5839,N_5797);
xnor U5972 (N_5972,N_5764,N_5834);
or U5973 (N_5973,N_5702,N_5755);
and U5974 (N_5974,N_5701,N_5700);
nor U5975 (N_5975,N_5771,N_5730);
nand U5976 (N_5976,N_5809,N_5839);
xor U5977 (N_5977,N_5714,N_5845);
or U5978 (N_5978,N_5724,N_5843);
or U5979 (N_5979,N_5792,N_5725);
nand U5980 (N_5980,N_5789,N_5829);
nor U5981 (N_5981,N_5802,N_5752);
or U5982 (N_5982,N_5723,N_5776);
xor U5983 (N_5983,N_5750,N_5806);
and U5984 (N_5984,N_5841,N_5838);
nand U5985 (N_5985,N_5824,N_5704);
xnor U5986 (N_5986,N_5770,N_5743);
nor U5987 (N_5987,N_5711,N_5771);
or U5988 (N_5988,N_5700,N_5704);
and U5989 (N_5989,N_5717,N_5723);
xnor U5990 (N_5990,N_5707,N_5722);
or U5991 (N_5991,N_5716,N_5730);
xnor U5992 (N_5992,N_5738,N_5811);
or U5993 (N_5993,N_5838,N_5842);
xor U5994 (N_5994,N_5722,N_5773);
xnor U5995 (N_5995,N_5805,N_5740);
or U5996 (N_5996,N_5839,N_5834);
nor U5997 (N_5997,N_5711,N_5751);
and U5998 (N_5998,N_5802,N_5812);
or U5999 (N_5999,N_5733,N_5771);
xnor U6000 (N_6000,N_5892,N_5987);
nand U6001 (N_6001,N_5881,N_5990);
or U6002 (N_6002,N_5933,N_5994);
and U6003 (N_6003,N_5925,N_5909);
xor U6004 (N_6004,N_5947,N_5949);
nor U6005 (N_6005,N_5857,N_5867);
nand U6006 (N_6006,N_5924,N_5906);
nand U6007 (N_6007,N_5991,N_5997);
nand U6008 (N_6008,N_5939,N_5916);
nor U6009 (N_6009,N_5913,N_5862);
nor U6010 (N_6010,N_5959,N_5888);
and U6011 (N_6011,N_5960,N_5945);
xor U6012 (N_6012,N_5989,N_5957);
nand U6013 (N_6013,N_5988,N_5978);
nand U6014 (N_6014,N_5850,N_5899);
nand U6015 (N_6015,N_5917,N_5943);
xnor U6016 (N_6016,N_5999,N_5941);
and U6017 (N_6017,N_5889,N_5920);
nor U6018 (N_6018,N_5908,N_5953);
nor U6019 (N_6019,N_5869,N_5885);
or U6020 (N_6020,N_5944,N_5969);
xor U6021 (N_6021,N_5878,N_5884);
and U6022 (N_6022,N_5858,N_5864);
nand U6023 (N_6023,N_5948,N_5852);
or U6024 (N_6024,N_5859,N_5874);
or U6025 (N_6025,N_5901,N_5897);
or U6026 (N_6026,N_5971,N_5940);
nand U6027 (N_6027,N_5932,N_5926);
nor U6028 (N_6028,N_5863,N_5895);
or U6029 (N_6029,N_5860,N_5914);
nand U6030 (N_6030,N_5883,N_5894);
nand U6031 (N_6031,N_5915,N_5993);
xnor U6032 (N_6032,N_5873,N_5865);
nand U6033 (N_6033,N_5985,N_5992);
nand U6034 (N_6034,N_5936,N_5856);
and U6035 (N_6035,N_5928,N_5977);
nand U6036 (N_6036,N_5972,N_5952);
nand U6037 (N_6037,N_5902,N_5967);
nor U6038 (N_6038,N_5882,N_5911);
nor U6039 (N_6039,N_5872,N_5886);
xnor U6040 (N_6040,N_5890,N_5996);
nand U6041 (N_6041,N_5958,N_5927);
xor U6042 (N_6042,N_5934,N_5950);
nor U6043 (N_6043,N_5923,N_5891);
nor U6044 (N_6044,N_5907,N_5931);
or U6045 (N_6045,N_5898,N_5968);
xnor U6046 (N_6046,N_5937,N_5903);
and U6047 (N_6047,N_5866,N_5922);
nand U6048 (N_6048,N_5976,N_5868);
nand U6049 (N_6049,N_5956,N_5893);
nand U6050 (N_6050,N_5983,N_5929);
and U6051 (N_6051,N_5887,N_5981);
xnor U6052 (N_6052,N_5975,N_5984);
xor U6053 (N_6053,N_5973,N_5855);
and U6054 (N_6054,N_5905,N_5918);
or U6055 (N_6055,N_5870,N_5963);
and U6056 (N_6056,N_5982,N_5912);
or U6057 (N_6057,N_5904,N_5979);
nand U6058 (N_6058,N_5946,N_5964);
xor U6059 (N_6059,N_5938,N_5930);
xor U6060 (N_6060,N_5951,N_5965);
and U6061 (N_6061,N_5910,N_5877);
nand U6062 (N_6062,N_5961,N_5876);
nand U6063 (N_6063,N_5995,N_5970);
xnor U6064 (N_6064,N_5998,N_5966);
xnor U6065 (N_6065,N_5879,N_5935);
or U6066 (N_6066,N_5880,N_5875);
nand U6067 (N_6067,N_5871,N_5955);
and U6068 (N_6068,N_5974,N_5854);
or U6069 (N_6069,N_5954,N_5861);
and U6070 (N_6070,N_5962,N_5851);
xor U6071 (N_6071,N_5980,N_5942);
or U6072 (N_6072,N_5919,N_5900);
and U6073 (N_6073,N_5853,N_5896);
or U6074 (N_6074,N_5986,N_5921);
and U6075 (N_6075,N_5931,N_5990);
nor U6076 (N_6076,N_5862,N_5893);
or U6077 (N_6077,N_5961,N_5858);
nand U6078 (N_6078,N_5880,N_5965);
and U6079 (N_6079,N_5862,N_5880);
nor U6080 (N_6080,N_5932,N_5912);
nand U6081 (N_6081,N_5927,N_5899);
nor U6082 (N_6082,N_5906,N_5971);
nand U6083 (N_6083,N_5857,N_5918);
xor U6084 (N_6084,N_5850,N_5966);
nand U6085 (N_6085,N_5957,N_5978);
or U6086 (N_6086,N_5933,N_5957);
and U6087 (N_6087,N_5946,N_5910);
or U6088 (N_6088,N_5925,N_5991);
nand U6089 (N_6089,N_5972,N_5947);
xnor U6090 (N_6090,N_5968,N_5970);
xor U6091 (N_6091,N_5901,N_5965);
and U6092 (N_6092,N_5999,N_5934);
and U6093 (N_6093,N_5992,N_5954);
or U6094 (N_6094,N_5873,N_5850);
nor U6095 (N_6095,N_5894,N_5870);
xor U6096 (N_6096,N_5922,N_5980);
nand U6097 (N_6097,N_5994,N_5873);
nor U6098 (N_6098,N_5921,N_5974);
xor U6099 (N_6099,N_5926,N_5952);
nand U6100 (N_6100,N_5970,N_5864);
and U6101 (N_6101,N_5894,N_5991);
xnor U6102 (N_6102,N_5895,N_5931);
and U6103 (N_6103,N_5855,N_5859);
or U6104 (N_6104,N_5874,N_5922);
or U6105 (N_6105,N_5979,N_5877);
and U6106 (N_6106,N_5882,N_5868);
xor U6107 (N_6107,N_5896,N_5902);
or U6108 (N_6108,N_5861,N_5995);
nor U6109 (N_6109,N_5903,N_5923);
and U6110 (N_6110,N_5940,N_5977);
or U6111 (N_6111,N_5913,N_5907);
and U6112 (N_6112,N_5915,N_5987);
and U6113 (N_6113,N_5929,N_5955);
nand U6114 (N_6114,N_5943,N_5905);
nand U6115 (N_6115,N_5998,N_5983);
nor U6116 (N_6116,N_5855,N_5942);
nand U6117 (N_6117,N_5930,N_5908);
nor U6118 (N_6118,N_5892,N_5881);
and U6119 (N_6119,N_5885,N_5933);
or U6120 (N_6120,N_5880,N_5926);
nand U6121 (N_6121,N_5858,N_5991);
nand U6122 (N_6122,N_5869,N_5992);
xor U6123 (N_6123,N_5945,N_5922);
or U6124 (N_6124,N_5892,N_5967);
or U6125 (N_6125,N_5999,N_5985);
or U6126 (N_6126,N_5862,N_5860);
xor U6127 (N_6127,N_5952,N_5852);
nand U6128 (N_6128,N_5871,N_5927);
nand U6129 (N_6129,N_5920,N_5942);
nand U6130 (N_6130,N_5974,N_5892);
xnor U6131 (N_6131,N_5898,N_5953);
nand U6132 (N_6132,N_5960,N_5924);
nor U6133 (N_6133,N_5912,N_5968);
nor U6134 (N_6134,N_5908,N_5967);
xnor U6135 (N_6135,N_5854,N_5860);
nand U6136 (N_6136,N_5913,N_5864);
nor U6137 (N_6137,N_5864,N_5917);
nand U6138 (N_6138,N_5981,N_5858);
nor U6139 (N_6139,N_5959,N_5997);
xor U6140 (N_6140,N_5908,N_5992);
or U6141 (N_6141,N_5960,N_5886);
xor U6142 (N_6142,N_5983,N_5910);
nor U6143 (N_6143,N_5968,N_5977);
nand U6144 (N_6144,N_5938,N_5934);
nand U6145 (N_6145,N_5997,N_5998);
xnor U6146 (N_6146,N_5885,N_5916);
nand U6147 (N_6147,N_5894,N_5971);
or U6148 (N_6148,N_5987,N_5981);
nand U6149 (N_6149,N_5906,N_5957);
xor U6150 (N_6150,N_6055,N_6032);
xor U6151 (N_6151,N_6129,N_6079);
nor U6152 (N_6152,N_6010,N_6034);
and U6153 (N_6153,N_6005,N_6103);
xnor U6154 (N_6154,N_6043,N_6053);
nand U6155 (N_6155,N_6081,N_6122);
nand U6156 (N_6156,N_6110,N_6117);
nor U6157 (N_6157,N_6024,N_6148);
and U6158 (N_6158,N_6126,N_6069);
xnor U6159 (N_6159,N_6134,N_6080);
or U6160 (N_6160,N_6112,N_6023);
nor U6161 (N_6161,N_6101,N_6042);
and U6162 (N_6162,N_6144,N_6044);
xnor U6163 (N_6163,N_6035,N_6124);
xor U6164 (N_6164,N_6012,N_6123);
or U6165 (N_6165,N_6064,N_6006);
nand U6166 (N_6166,N_6095,N_6108);
xnor U6167 (N_6167,N_6128,N_6036);
nor U6168 (N_6168,N_6030,N_6118);
nor U6169 (N_6169,N_6149,N_6120);
nor U6170 (N_6170,N_6115,N_6119);
or U6171 (N_6171,N_6106,N_6013);
or U6172 (N_6172,N_6008,N_6105);
or U6173 (N_6173,N_6033,N_6072);
and U6174 (N_6174,N_6050,N_6138);
nor U6175 (N_6175,N_6029,N_6109);
and U6176 (N_6176,N_6021,N_6140);
nor U6177 (N_6177,N_6074,N_6048);
nand U6178 (N_6178,N_6039,N_6022);
nor U6179 (N_6179,N_6056,N_6054);
nand U6180 (N_6180,N_6058,N_6094);
or U6181 (N_6181,N_6096,N_6070);
or U6182 (N_6182,N_6015,N_6028);
nand U6183 (N_6183,N_6073,N_6037);
nor U6184 (N_6184,N_6063,N_6040);
xor U6185 (N_6185,N_6003,N_6000);
nor U6186 (N_6186,N_6045,N_6086);
nor U6187 (N_6187,N_6143,N_6136);
nand U6188 (N_6188,N_6062,N_6049);
or U6189 (N_6189,N_6065,N_6099);
xor U6190 (N_6190,N_6046,N_6009);
xnor U6191 (N_6191,N_6145,N_6084);
nor U6192 (N_6192,N_6061,N_6025);
nor U6193 (N_6193,N_6016,N_6077);
and U6194 (N_6194,N_6098,N_6047);
and U6195 (N_6195,N_6087,N_6026);
nor U6196 (N_6196,N_6071,N_6057);
nor U6197 (N_6197,N_6097,N_6102);
or U6198 (N_6198,N_6116,N_6066);
or U6199 (N_6199,N_6017,N_6137);
nand U6200 (N_6200,N_6002,N_6011);
and U6201 (N_6201,N_6127,N_6004);
or U6202 (N_6202,N_6104,N_6083);
and U6203 (N_6203,N_6132,N_6113);
xnor U6204 (N_6204,N_6082,N_6092);
and U6205 (N_6205,N_6111,N_6060);
or U6206 (N_6206,N_6051,N_6089);
xor U6207 (N_6207,N_6019,N_6125);
xnor U6208 (N_6208,N_6052,N_6068);
xnor U6209 (N_6209,N_6031,N_6014);
or U6210 (N_6210,N_6135,N_6146);
nand U6211 (N_6211,N_6141,N_6001);
and U6212 (N_6212,N_6067,N_6121);
nor U6213 (N_6213,N_6093,N_6090);
or U6214 (N_6214,N_6059,N_6088);
nand U6215 (N_6215,N_6027,N_6100);
nand U6216 (N_6216,N_6147,N_6133);
xnor U6217 (N_6217,N_6018,N_6076);
nand U6218 (N_6218,N_6114,N_6139);
nand U6219 (N_6219,N_6091,N_6007);
nand U6220 (N_6220,N_6130,N_6041);
nor U6221 (N_6221,N_6107,N_6142);
or U6222 (N_6222,N_6131,N_6020);
and U6223 (N_6223,N_6085,N_6075);
nor U6224 (N_6224,N_6038,N_6078);
nand U6225 (N_6225,N_6099,N_6108);
and U6226 (N_6226,N_6025,N_6024);
or U6227 (N_6227,N_6010,N_6147);
nor U6228 (N_6228,N_6097,N_6063);
or U6229 (N_6229,N_6000,N_6122);
nor U6230 (N_6230,N_6051,N_6137);
nor U6231 (N_6231,N_6141,N_6103);
xnor U6232 (N_6232,N_6143,N_6067);
xor U6233 (N_6233,N_6047,N_6010);
and U6234 (N_6234,N_6010,N_6141);
or U6235 (N_6235,N_6023,N_6019);
nand U6236 (N_6236,N_6080,N_6016);
xor U6237 (N_6237,N_6013,N_6018);
or U6238 (N_6238,N_6141,N_6052);
or U6239 (N_6239,N_6128,N_6122);
nand U6240 (N_6240,N_6040,N_6120);
nor U6241 (N_6241,N_6022,N_6044);
and U6242 (N_6242,N_6052,N_6071);
xor U6243 (N_6243,N_6096,N_6136);
and U6244 (N_6244,N_6094,N_6102);
or U6245 (N_6245,N_6046,N_6127);
or U6246 (N_6246,N_6086,N_6102);
nor U6247 (N_6247,N_6006,N_6025);
nor U6248 (N_6248,N_6043,N_6071);
nor U6249 (N_6249,N_6005,N_6000);
and U6250 (N_6250,N_6144,N_6061);
or U6251 (N_6251,N_6083,N_6085);
or U6252 (N_6252,N_6075,N_6128);
nand U6253 (N_6253,N_6040,N_6015);
xor U6254 (N_6254,N_6049,N_6000);
and U6255 (N_6255,N_6023,N_6024);
nand U6256 (N_6256,N_6080,N_6086);
or U6257 (N_6257,N_6078,N_6027);
and U6258 (N_6258,N_6075,N_6054);
nand U6259 (N_6259,N_6038,N_6111);
nor U6260 (N_6260,N_6057,N_6019);
xnor U6261 (N_6261,N_6005,N_6134);
nor U6262 (N_6262,N_6003,N_6025);
nor U6263 (N_6263,N_6122,N_6019);
or U6264 (N_6264,N_6036,N_6101);
or U6265 (N_6265,N_6134,N_6065);
and U6266 (N_6266,N_6042,N_6028);
nor U6267 (N_6267,N_6048,N_6085);
or U6268 (N_6268,N_6058,N_6054);
xor U6269 (N_6269,N_6033,N_6053);
and U6270 (N_6270,N_6113,N_6021);
nand U6271 (N_6271,N_6110,N_6020);
xnor U6272 (N_6272,N_6147,N_6111);
nor U6273 (N_6273,N_6099,N_6135);
nand U6274 (N_6274,N_6021,N_6071);
xnor U6275 (N_6275,N_6128,N_6031);
nand U6276 (N_6276,N_6063,N_6071);
nor U6277 (N_6277,N_6081,N_6057);
or U6278 (N_6278,N_6027,N_6131);
nand U6279 (N_6279,N_6050,N_6076);
nand U6280 (N_6280,N_6077,N_6109);
or U6281 (N_6281,N_6103,N_6004);
and U6282 (N_6282,N_6045,N_6016);
xor U6283 (N_6283,N_6049,N_6015);
nor U6284 (N_6284,N_6068,N_6040);
nand U6285 (N_6285,N_6106,N_6029);
nor U6286 (N_6286,N_6108,N_6141);
nor U6287 (N_6287,N_6127,N_6141);
or U6288 (N_6288,N_6077,N_6115);
or U6289 (N_6289,N_6018,N_6075);
nand U6290 (N_6290,N_6093,N_6131);
nor U6291 (N_6291,N_6081,N_6096);
or U6292 (N_6292,N_6138,N_6066);
or U6293 (N_6293,N_6029,N_6141);
or U6294 (N_6294,N_6039,N_6002);
nor U6295 (N_6295,N_6050,N_6022);
nand U6296 (N_6296,N_6027,N_6112);
xor U6297 (N_6297,N_6001,N_6089);
nor U6298 (N_6298,N_6147,N_6039);
xnor U6299 (N_6299,N_6089,N_6015);
nor U6300 (N_6300,N_6269,N_6195);
and U6301 (N_6301,N_6287,N_6290);
and U6302 (N_6302,N_6256,N_6291);
xnor U6303 (N_6303,N_6243,N_6220);
or U6304 (N_6304,N_6258,N_6216);
xnor U6305 (N_6305,N_6214,N_6155);
or U6306 (N_6306,N_6280,N_6190);
nor U6307 (N_6307,N_6180,N_6191);
or U6308 (N_6308,N_6179,N_6233);
nand U6309 (N_6309,N_6197,N_6242);
or U6310 (N_6310,N_6150,N_6182);
nor U6311 (N_6311,N_6249,N_6209);
nor U6312 (N_6312,N_6297,N_6298);
nand U6313 (N_6313,N_6273,N_6227);
nor U6314 (N_6314,N_6270,N_6176);
xnor U6315 (N_6315,N_6283,N_6282);
and U6316 (N_6316,N_6255,N_6274);
nor U6317 (N_6317,N_6163,N_6203);
nor U6318 (N_6318,N_6223,N_6293);
and U6319 (N_6319,N_6228,N_6276);
xor U6320 (N_6320,N_6252,N_6251);
xnor U6321 (N_6321,N_6254,N_6212);
nor U6322 (N_6322,N_6188,N_6263);
nand U6323 (N_6323,N_6198,N_6286);
nand U6324 (N_6324,N_6204,N_6164);
nor U6325 (N_6325,N_6238,N_6262);
xnor U6326 (N_6326,N_6161,N_6217);
or U6327 (N_6327,N_6194,N_6207);
xor U6328 (N_6328,N_6272,N_6205);
nand U6329 (N_6329,N_6157,N_6247);
or U6330 (N_6330,N_6152,N_6178);
and U6331 (N_6331,N_6211,N_6261);
or U6332 (N_6332,N_6170,N_6237);
nor U6333 (N_6333,N_6232,N_6193);
and U6334 (N_6334,N_6200,N_6235);
nand U6335 (N_6335,N_6271,N_6196);
xor U6336 (N_6336,N_6202,N_6264);
nor U6337 (N_6337,N_6166,N_6218);
or U6338 (N_6338,N_6186,N_6168);
or U6339 (N_6339,N_6185,N_6184);
nor U6340 (N_6340,N_6277,N_6284);
or U6341 (N_6341,N_6279,N_6244);
and U6342 (N_6342,N_6172,N_6208);
xor U6343 (N_6343,N_6219,N_6158);
and U6344 (N_6344,N_6201,N_6224);
nand U6345 (N_6345,N_6175,N_6257);
and U6346 (N_6346,N_6295,N_6173);
or U6347 (N_6347,N_6153,N_6292);
and U6348 (N_6348,N_6151,N_6296);
nand U6349 (N_6349,N_6281,N_6192);
or U6350 (N_6350,N_6222,N_6167);
or U6351 (N_6351,N_6240,N_6288);
nand U6352 (N_6352,N_6248,N_6189);
nand U6353 (N_6353,N_6159,N_6169);
nor U6354 (N_6354,N_6187,N_6285);
or U6355 (N_6355,N_6250,N_6253);
and U6356 (N_6356,N_6230,N_6162);
xnor U6357 (N_6357,N_6265,N_6289);
nand U6358 (N_6358,N_6210,N_6206);
nor U6359 (N_6359,N_6259,N_6181);
xnor U6360 (N_6360,N_6165,N_6267);
or U6361 (N_6361,N_6229,N_6177);
xnor U6362 (N_6362,N_6226,N_6299);
and U6363 (N_6363,N_6239,N_6183);
xnor U6364 (N_6364,N_6213,N_6278);
nand U6365 (N_6365,N_6245,N_6294);
nor U6366 (N_6366,N_6246,N_6215);
nor U6367 (N_6367,N_6231,N_6221);
nand U6368 (N_6368,N_6156,N_6174);
nor U6369 (N_6369,N_6268,N_6241);
nor U6370 (N_6370,N_6154,N_6234);
nand U6371 (N_6371,N_6260,N_6266);
nand U6372 (N_6372,N_6160,N_6199);
nand U6373 (N_6373,N_6236,N_6171);
nor U6374 (N_6374,N_6225,N_6275);
nand U6375 (N_6375,N_6248,N_6154);
or U6376 (N_6376,N_6176,N_6266);
nor U6377 (N_6377,N_6190,N_6249);
or U6378 (N_6378,N_6280,N_6253);
nand U6379 (N_6379,N_6282,N_6164);
xnor U6380 (N_6380,N_6201,N_6280);
xnor U6381 (N_6381,N_6233,N_6202);
and U6382 (N_6382,N_6200,N_6193);
or U6383 (N_6383,N_6254,N_6274);
nand U6384 (N_6384,N_6206,N_6194);
nand U6385 (N_6385,N_6230,N_6152);
or U6386 (N_6386,N_6172,N_6288);
or U6387 (N_6387,N_6198,N_6186);
xor U6388 (N_6388,N_6272,N_6243);
nor U6389 (N_6389,N_6272,N_6203);
nand U6390 (N_6390,N_6165,N_6214);
xor U6391 (N_6391,N_6229,N_6210);
nand U6392 (N_6392,N_6275,N_6171);
nand U6393 (N_6393,N_6156,N_6254);
nand U6394 (N_6394,N_6231,N_6217);
nand U6395 (N_6395,N_6244,N_6232);
nand U6396 (N_6396,N_6167,N_6272);
and U6397 (N_6397,N_6268,N_6192);
nand U6398 (N_6398,N_6205,N_6173);
or U6399 (N_6399,N_6264,N_6259);
nor U6400 (N_6400,N_6286,N_6272);
xor U6401 (N_6401,N_6192,N_6161);
nand U6402 (N_6402,N_6150,N_6197);
or U6403 (N_6403,N_6182,N_6282);
nor U6404 (N_6404,N_6249,N_6246);
nor U6405 (N_6405,N_6209,N_6150);
xor U6406 (N_6406,N_6289,N_6239);
nand U6407 (N_6407,N_6227,N_6290);
nand U6408 (N_6408,N_6204,N_6292);
or U6409 (N_6409,N_6282,N_6195);
xnor U6410 (N_6410,N_6268,N_6281);
and U6411 (N_6411,N_6181,N_6283);
xnor U6412 (N_6412,N_6215,N_6273);
and U6413 (N_6413,N_6223,N_6253);
or U6414 (N_6414,N_6257,N_6212);
or U6415 (N_6415,N_6277,N_6222);
nand U6416 (N_6416,N_6295,N_6298);
nor U6417 (N_6417,N_6190,N_6167);
and U6418 (N_6418,N_6151,N_6183);
nand U6419 (N_6419,N_6170,N_6174);
nand U6420 (N_6420,N_6226,N_6264);
nand U6421 (N_6421,N_6287,N_6255);
nor U6422 (N_6422,N_6245,N_6260);
nor U6423 (N_6423,N_6180,N_6241);
or U6424 (N_6424,N_6262,N_6196);
and U6425 (N_6425,N_6258,N_6269);
xor U6426 (N_6426,N_6262,N_6240);
xnor U6427 (N_6427,N_6161,N_6241);
nand U6428 (N_6428,N_6289,N_6258);
xnor U6429 (N_6429,N_6190,N_6199);
and U6430 (N_6430,N_6269,N_6212);
xnor U6431 (N_6431,N_6265,N_6242);
and U6432 (N_6432,N_6207,N_6195);
and U6433 (N_6433,N_6206,N_6281);
or U6434 (N_6434,N_6207,N_6157);
xor U6435 (N_6435,N_6241,N_6294);
and U6436 (N_6436,N_6191,N_6153);
xor U6437 (N_6437,N_6153,N_6263);
and U6438 (N_6438,N_6278,N_6172);
and U6439 (N_6439,N_6265,N_6280);
or U6440 (N_6440,N_6234,N_6183);
nor U6441 (N_6441,N_6294,N_6198);
or U6442 (N_6442,N_6232,N_6174);
and U6443 (N_6443,N_6243,N_6208);
xnor U6444 (N_6444,N_6220,N_6254);
nor U6445 (N_6445,N_6259,N_6173);
and U6446 (N_6446,N_6289,N_6254);
xnor U6447 (N_6447,N_6276,N_6188);
nand U6448 (N_6448,N_6259,N_6209);
nand U6449 (N_6449,N_6269,N_6275);
or U6450 (N_6450,N_6364,N_6357);
xor U6451 (N_6451,N_6359,N_6316);
xnor U6452 (N_6452,N_6337,N_6446);
nand U6453 (N_6453,N_6375,N_6396);
nand U6454 (N_6454,N_6448,N_6300);
nand U6455 (N_6455,N_6352,N_6336);
xnor U6456 (N_6456,N_6304,N_6413);
and U6457 (N_6457,N_6407,N_6447);
or U6458 (N_6458,N_6314,N_6310);
nor U6459 (N_6459,N_6319,N_6440);
or U6460 (N_6460,N_6422,N_6428);
nand U6461 (N_6461,N_6356,N_6429);
nand U6462 (N_6462,N_6311,N_6346);
nor U6463 (N_6463,N_6355,N_6320);
or U6464 (N_6464,N_6431,N_6303);
nand U6465 (N_6465,N_6317,N_6387);
nor U6466 (N_6466,N_6441,N_6312);
and U6467 (N_6467,N_6394,N_6335);
xnor U6468 (N_6468,N_6326,N_6308);
and U6469 (N_6469,N_6384,N_6372);
xor U6470 (N_6470,N_6349,N_6433);
nor U6471 (N_6471,N_6382,N_6432);
xor U6472 (N_6472,N_6302,N_6445);
or U6473 (N_6473,N_6309,N_6323);
xor U6474 (N_6474,N_6385,N_6362);
or U6475 (N_6475,N_6439,N_6412);
or U6476 (N_6476,N_6415,N_6344);
nand U6477 (N_6477,N_6373,N_6327);
xnor U6478 (N_6478,N_6376,N_6391);
nor U6479 (N_6479,N_6435,N_6401);
nor U6480 (N_6480,N_6353,N_6430);
and U6481 (N_6481,N_6423,N_6426);
or U6482 (N_6482,N_6379,N_6417);
and U6483 (N_6483,N_6399,N_6307);
nand U6484 (N_6484,N_6367,N_6437);
or U6485 (N_6485,N_6334,N_6354);
and U6486 (N_6486,N_6404,N_6390);
nor U6487 (N_6487,N_6351,N_6421);
or U6488 (N_6488,N_6398,N_6322);
and U6489 (N_6489,N_6424,N_6330);
and U6490 (N_6490,N_6315,N_6395);
and U6491 (N_6491,N_6383,N_6389);
nand U6492 (N_6492,N_6414,N_6370);
and U6493 (N_6493,N_6388,N_6408);
and U6494 (N_6494,N_6360,N_6331);
xor U6495 (N_6495,N_6411,N_6416);
and U6496 (N_6496,N_6444,N_6425);
xor U6497 (N_6497,N_6325,N_6368);
nand U6498 (N_6498,N_6403,N_6381);
xnor U6499 (N_6499,N_6329,N_6333);
nor U6500 (N_6500,N_6380,N_6434);
nand U6501 (N_6501,N_6348,N_6363);
nor U6502 (N_6502,N_6341,N_6347);
and U6503 (N_6503,N_6342,N_6321);
or U6504 (N_6504,N_6369,N_6305);
nand U6505 (N_6505,N_6377,N_6343);
nor U6506 (N_6506,N_6436,N_6405);
and U6507 (N_6507,N_6419,N_6442);
or U6508 (N_6508,N_6324,N_6350);
or U6509 (N_6509,N_6371,N_6361);
nand U6510 (N_6510,N_6378,N_6328);
xor U6511 (N_6511,N_6420,N_6345);
xor U6512 (N_6512,N_6427,N_6366);
and U6513 (N_6513,N_6410,N_6438);
and U6514 (N_6514,N_6374,N_6313);
and U6515 (N_6515,N_6449,N_6306);
nand U6516 (N_6516,N_6358,N_6418);
nor U6517 (N_6517,N_6393,N_6400);
xor U6518 (N_6518,N_6392,N_6402);
xnor U6519 (N_6519,N_6318,N_6365);
or U6520 (N_6520,N_6332,N_6339);
xor U6521 (N_6521,N_6340,N_6338);
nand U6522 (N_6522,N_6397,N_6409);
and U6523 (N_6523,N_6301,N_6386);
nor U6524 (N_6524,N_6443,N_6406);
xnor U6525 (N_6525,N_6309,N_6402);
or U6526 (N_6526,N_6368,N_6330);
nor U6527 (N_6527,N_6385,N_6355);
nand U6528 (N_6528,N_6303,N_6386);
or U6529 (N_6529,N_6331,N_6372);
or U6530 (N_6530,N_6352,N_6369);
nand U6531 (N_6531,N_6420,N_6428);
and U6532 (N_6532,N_6401,N_6339);
and U6533 (N_6533,N_6402,N_6333);
or U6534 (N_6534,N_6436,N_6336);
xnor U6535 (N_6535,N_6308,N_6446);
nand U6536 (N_6536,N_6303,N_6418);
xnor U6537 (N_6537,N_6440,N_6394);
xor U6538 (N_6538,N_6312,N_6371);
and U6539 (N_6539,N_6445,N_6400);
or U6540 (N_6540,N_6427,N_6409);
nand U6541 (N_6541,N_6334,N_6335);
nand U6542 (N_6542,N_6384,N_6325);
nor U6543 (N_6543,N_6425,N_6420);
nor U6544 (N_6544,N_6400,N_6357);
xor U6545 (N_6545,N_6371,N_6322);
and U6546 (N_6546,N_6303,N_6426);
nand U6547 (N_6547,N_6416,N_6343);
and U6548 (N_6548,N_6304,N_6429);
nor U6549 (N_6549,N_6328,N_6410);
or U6550 (N_6550,N_6338,N_6343);
or U6551 (N_6551,N_6304,N_6326);
or U6552 (N_6552,N_6323,N_6356);
and U6553 (N_6553,N_6418,N_6441);
or U6554 (N_6554,N_6353,N_6355);
nand U6555 (N_6555,N_6301,N_6378);
or U6556 (N_6556,N_6318,N_6328);
and U6557 (N_6557,N_6419,N_6341);
nand U6558 (N_6558,N_6343,N_6359);
or U6559 (N_6559,N_6300,N_6355);
xnor U6560 (N_6560,N_6323,N_6406);
xnor U6561 (N_6561,N_6401,N_6351);
xnor U6562 (N_6562,N_6311,N_6434);
or U6563 (N_6563,N_6359,N_6376);
and U6564 (N_6564,N_6363,N_6358);
and U6565 (N_6565,N_6349,N_6318);
or U6566 (N_6566,N_6390,N_6329);
and U6567 (N_6567,N_6372,N_6332);
or U6568 (N_6568,N_6417,N_6344);
nor U6569 (N_6569,N_6439,N_6358);
xnor U6570 (N_6570,N_6378,N_6447);
xor U6571 (N_6571,N_6357,N_6430);
nor U6572 (N_6572,N_6387,N_6389);
xnor U6573 (N_6573,N_6347,N_6321);
nor U6574 (N_6574,N_6356,N_6397);
or U6575 (N_6575,N_6412,N_6398);
or U6576 (N_6576,N_6336,N_6329);
nand U6577 (N_6577,N_6409,N_6398);
and U6578 (N_6578,N_6426,N_6428);
xnor U6579 (N_6579,N_6353,N_6334);
and U6580 (N_6580,N_6360,N_6328);
nand U6581 (N_6581,N_6400,N_6378);
nor U6582 (N_6582,N_6415,N_6319);
nand U6583 (N_6583,N_6347,N_6404);
and U6584 (N_6584,N_6361,N_6407);
and U6585 (N_6585,N_6374,N_6353);
or U6586 (N_6586,N_6304,N_6428);
and U6587 (N_6587,N_6369,N_6368);
xor U6588 (N_6588,N_6394,N_6347);
or U6589 (N_6589,N_6338,N_6429);
nand U6590 (N_6590,N_6362,N_6368);
nand U6591 (N_6591,N_6389,N_6424);
nand U6592 (N_6592,N_6336,N_6350);
nor U6593 (N_6593,N_6300,N_6339);
nand U6594 (N_6594,N_6358,N_6409);
xor U6595 (N_6595,N_6400,N_6407);
xor U6596 (N_6596,N_6420,N_6353);
nand U6597 (N_6597,N_6428,N_6323);
xor U6598 (N_6598,N_6394,N_6333);
or U6599 (N_6599,N_6365,N_6417);
nand U6600 (N_6600,N_6522,N_6552);
and U6601 (N_6601,N_6528,N_6495);
or U6602 (N_6602,N_6513,N_6489);
and U6603 (N_6603,N_6558,N_6578);
nand U6604 (N_6604,N_6451,N_6459);
and U6605 (N_6605,N_6565,N_6568);
xnor U6606 (N_6606,N_6564,N_6469);
and U6607 (N_6607,N_6595,N_6493);
and U6608 (N_6608,N_6571,N_6572);
nor U6609 (N_6609,N_6580,N_6547);
or U6610 (N_6610,N_6484,N_6476);
or U6611 (N_6611,N_6553,N_6579);
or U6612 (N_6612,N_6587,N_6458);
and U6613 (N_6613,N_6541,N_6574);
xnor U6614 (N_6614,N_6598,N_6550);
or U6615 (N_6615,N_6457,N_6570);
xnor U6616 (N_6616,N_6583,N_6487);
nand U6617 (N_6617,N_6470,N_6546);
nor U6618 (N_6618,N_6536,N_6539);
nor U6619 (N_6619,N_6505,N_6534);
xor U6620 (N_6620,N_6498,N_6511);
or U6621 (N_6621,N_6485,N_6454);
nand U6622 (N_6622,N_6588,N_6562);
nor U6623 (N_6623,N_6460,N_6504);
or U6624 (N_6624,N_6537,N_6532);
nor U6625 (N_6625,N_6491,N_6518);
or U6626 (N_6626,N_6566,N_6509);
or U6627 (N_6627,N_6549,N_6555);
nand U6628 (N_6628,N_6488,N_6502);
xor U6629 (N_6629,N_6575,N_6545);
nand U6630 (N_6630,N_6452,N_6506);
xor U6631 (N_6631,N_6510,N_6473);
and U6632 (N_6632,N_6573,N_6560);
or U6633 (N_6633,N_6543,N_6557);
and U6634 (N_6634,N_6512,N_6576);
and U6635 (N_6635,N_6586,N_6599);
or U6636 (N_6636,N_6519,N_6517);
and U6637 (N_6637,N_6471,N_6478);
nand U6638 (N_6638,N_6563,N_6523);
xnor U6639 (N_6639,N_6569,N_6464);
xnor U6640 (N_6640,N_6490,N_6590);
and U6641 (N_6641,N_6482,N_6592);
or U6642 (N_6642,N_6492,N_6533);
nor U6643 (N_6643,N_6463,N_6529);
and U6644 (N_6644,N_6597,N_6499);
nand U6645 (N_6645,N_6581,N_6594);
or U6646 (N_6646,N_6479,N_6589);
and U6647 (N_6647,N_6561,N_6465);
nor U6648 (N_6648,N_6593,N_6500);
nand U6649 (N_6649,N_6526,N_6556);
nand U6650 (N_6650,N_6584,N_6535);
nor U6651 (N_6651,N_6466,N_6467);
or U6652 (N_6652,N_6462,N_6475);
or U6653 (N_6653,N_6525,N_6548);
nand U6654 (N_6654,N_6567,N_6520);
nor U6655 (N_6655,N_6521,N_6591);
xnor U6656 (N_6656,N_6540,N_6483);
or U6657 (N_6657,N_6472,N_6474);
or U6658 (N_6658,N_6559,N_6494);
nand U6659 (N_6659,N_6480,N_6514);
or U6660 (N_6660,N_6577,N_6507);
nand U6661 (N_6661,N_6486,N_6453);
and U6662 (N_6662,N_6524,N_6538);
and U6663 (N_6663,N_6531,N_6516);
nand U6664 (N_6664,N_6477,N_6542);
nor U6665 (N_6665,N_6554,N_6544);
nand U6666 (N_6666,N_6497,N_6508);
xnor U6667 (N_6667,N_6530,N_6596);
or U6668 (N_6668,N_6456,N_6501);
xnor U6669 (N_6669,N_6503,N_6461);
or U6670 (N_6670,N_6455,N_6468);
xnor U6671 (N_6671,N_6585,N_6450);
nand U6672 (N_6672,N_6515,N_6527);
nand U6673 (N_6673,N_6582,N_6496);
nand U6674 (N_6674,N_6481,N_6551);
nand U6675 (N_6675,N_6488,N_6581);
or U6676 (N_6676,N_6573,N_6477);
nand U6677 (N_6677,N_6467,N_6510);
nand U6678 (N_6678,N_6473,N_6586);
and U6679 (N_6679,N_6570,N_6476);
nor U6680 (N_6680,N_6461,N_6514);
nor U6681 (N_6681,N_6525,N_6555);
nand U6682 (N_6682,N_6490,N_6579);
and U6683 (N_6683,N_6508,N_6589);
and U6684 (N_6684,N_6525,N_6453);
nand U6685 (N_6685,N_6559,N_6503);
and U6686 (N_6686,N_6476,N_6521);
and U6687 (N_6687,N_6599,N_6563);
and U6688 (N_6688,N_6536,N_6541);
nand U6689 (N_6689,N_6528,N_6564);
xor U6690 (N_6690,N_6595,N_6480);
nand U6691 (N_6691,N_6482,N_6545);
and U6692 (N_6692,N_6513,N_6547);
nor U6693 (N_6693,N_6451,N_6495);
nor U6694 (N_6694,N_6555,N_6529);
xor U6695 (N_6695,N_6590,N_6561);
or U6696 (N_6696,N_6524,N_6471);
or U6697 (N_6697,N_6500,N_6452);
nand U6698 (N_6698,N_6450,N_6528);
nand U6699 (N_6699,N_6509,N_6491);
or U6700 (N_6700,N_6548,N_6460);
or U6701 (N_6701,N_6520,N_6570);
or U6702 (N_6702,N_6513,N_6534);
or U6703 (N_6703,N_6528,N_6545);
xnor U6704 (N_6704,N_6470,N_6538);
and U6705 (N_6705,N_6506,N_6592);
nand U6706 (N_6706,N_6498,N_6517);
and U6707 (N_6707,N_6510,N_6463);
and U6708 (N_6708,N_6587,N_6557);
nand U6709 (N_6709,N_6559,N_6541);
nor U6710 (N_6710,N_6453,N_6455);
nand U6711 (N_6711,N_6519,N_6525);
and U6712 (N_6712,N_6550,N_6470);
and U6713 (N_6713,N_6462,N_6577);
xnor U6714 (N_6714,N_6501,N_6476);
xnor U6715 (N_6715,N_6474,N_6558);
nand U6716 (N_6716,N_6567,N_6457);
or U6717 (N_6717,N_6508,N_6565);
nor U6718 (N_6718,N_6556,N_6552);
nand U6719 (N_6719,N_6541,N_6570);
xnor U6720 (N_6720,N_6487,N_6495);
and U6721 (N_6721,N_6575,N_6542);
nor U6722 (N_6722,N_6567,N_6596);
nand U6723 (N_6723,N_6545,N_6560);
nand U6724 (N_6724,N_6465,N_6531);
nand U6725 (N_6725,N_6567,N_6454);
nor U6726 (N_6726,N_6467,N_6472);
nor U6727 (N_6727,N_6550,N_6552);
or U6728 (N_6728,N_6518,N_6550);
nand U6729 (N_6729,N_6464,N_6473);
nand U6730 (N_6730,N_6456,N_6524);
xor U6731 (N_6731,N_6590,N_6584);
nand U6732 (N_6732,N_6598,N_6599);
and U6733 (N_6733,N_6481,N_6465);
or U6734 (N_6734,N_6499,N_6452);
nand U6735 (N_6735,N_6455,N_6514);
and U6736 (N_6736,N_6511,N_6565);
and U6737 (N_6737,N_6570,N_6511);
or U6738 (N_6738,N_6597,N_6470);
nor U6739 (N_6739,N_6527,N_6465);
and U6740 (N_6740,N_6535,N_6524);
nor U6741 (N_6741,N_6573,N_6599);
or U6742 (N_6742,N_6463,N_6454);
nand U6743 (N_6743,N_6505,N_6478);
nor U6744 (N_6744,N_6463,N_6494);
nor U6745 (N_6745,N_6597,N_6460);
xor U6746 (N_6746,N_6559,N_6490);
nor U6747 (N_6747,N_6534,N_6490);
xor U6748 (N_6748,N_6569,N_6553);
and U6749 (N_6749,N_6593,N_6537);
and U6750 (N_6750,N_6694,N_6688);
nor U6751 (N_6751,N_6678,N_6630);
and U6752 (N_6752,N_6676,N_6671);
xnor U6753 (N_6753,N_6712,N_6628);
or U6754 (N_6754,N_6647,N_6746);
nand U6755 (N_6755,N_6657,N_6714);
xor U6756 (N_6756,N_6677,N_6605);
nand U6757 (N_6757,N_6640,N_6743);
and U6758 (N_6758,N_6728,N_6708);
or U6759 (N_6759,N_6650,N_6709);
xnor U6760 (N_6760,N_6698,N_6655);
or U6761 (N_6761,N_6644,N_6689);
nor U6762 (N_6762,N_6690,N_6725);
xnor U6763 (N_6763,N_6631,N_6603);
and U6764 (N_6764,N_6736,N_6619);
xor U6765 (N_6765,N_6648,N_6740);
and U6766 (N_6766,N_6713,N_6741);
or U6767 (N_6767,N_6719,N_6699);
or U6768 (N_6768,N_6666,N_6695);
nand U6769 (N_6769,N_6724,N_6726);
or U6770 (N_6770,N_6601,N_6645);
and U6771 (N_6771,N_6621,N_6654);
or U6772 (N_6772,N_6748,N_6663);
or U6773 (N_6773,N_6646,N_6623);
nand U6774 (N_6774,N_6737,N_6691);
nand U6775 (N_6775,N_6634,N_6617);
nor U6776 (N_6776,N_6609,N_6668);
nand U6777 (N_6777,N_6638,N_6747);
xnor U6778 (N_6778,N_6735,N_6729);
or U6779 (N_6779,N_6625,N_6607);
nand U6780 (N_6780,N_6706,N_6613);
nor U6781 (N_6781,N_6711,N_6656);
or U6782 (N_6782,N_6652,N_6685);
or U6783 (N_6783,N_6679,N_6680);
nor U6784 (N_6784,N_6608,N_6624);
nand U6785 (N_6785,N_6675,N_6693);
nand U6786 (N_6786,N_6633,N_6701);
nand U6787 (N_6787,N_6684,N_6710);
nor U6788 (N_6788,N_6664,N_6742);
and U6789 (N_6789,N_6641,N_6635);
nor U6790 (N_6790,N_6732,N_6720);
or U6791 (N_6791,N_6683,N_6702);
or U6792 (N_6792,N_6700,N_6727);
nor U6793 (N_6793,N_6600,N_6611);
xnor U6794 (N_6794,N_6620,N_6723);
or U6795 (N_6795,N_6739,N_6749);
and U6796 (N_6796,N_6642,N_6653);
xor U6797 (N_6797,N_6718,N_6697);
xor U6798 (N_6798,N_6661,N_6660);
or U6799 (N_6799,N_6730,N_6681);
and U6800 (N_6800,N_6721,N_6696);
xor U6801 (N_6801,N_6649,N_6662);
or U6802 (N_6802,N_6602,N_6626);
xnor U6803 (N_6803,N_6682,N_6704);
xnor U6804 (N_6804,N_6674,N_6672);
nor U6805 (N_6805,N_6717,N_6636);
or U6806 (N_6806,N_6658,N_6733);
or U6807 (N_6807,N_6618,N_6715);
or U6808 (N_6808,N_6651,N_6637);
nor U6809 (N_6809,N_6615,N_6629);
nand U6810 (N_6810,N_6616,N_6744);
xnor U6811 (N_6811,N_6622,N_6705);
and U6812 (N_6812,N_6731,N_6692);
nand U6813 (N_6813,N_6604,N_6606);
nand U6814 (N_6814,N_6703,N_6632);
xor U6815 (N_6815,N_6716,N_6667);
and U6816 (N_6816,N_6610,N_6627);
xor U6817 (N_6817,N_6665,N_6738);
and U6818 (N_6818,N_6639,N_6722);
and U6819 (N_6819,N_6686,N_6673);
or U6820 (N_6820,N_6612,N_6670);
nor U6821 (N_6821,N_6669,N_6614);
nand U6822 (N_6822,N_6734,N_6659);
nor U6823 (N_6823,N_6745,N_6687);
or U6824 (N_6824,N_6643,N_6707);
xor U6825 (N_6825,N_6713,N_6639);
xnor U6826 (N_6826,N_6694,N_6612);
nand U6827 (N_6827,N_6717,N_6656);
xor U6828 (N_6828,N_6672,N_6618);
nor U6829 (N_6829,N_6693,N_6666);
and U6830 (N_6830,N_6602,N_6686);
or U6831 (N_6831,N_6732,N_6651);
or U6832 (N_6832,N_6740,N_6606);
nand U6833 (N_6833,N_6605,N_6601);
or U6834 (N_6834,N_6727,N_6661);
and U6835 (N_6835,N_6642,N_6621);
and U6836 (N_6836,N_6661,N_6715);
or U6837 (N_6837,N_6616,N_6666);
or U6838 (N_6838,N_6600,N_6732);
or U6839 (N_6839,N_6691,N_6642);
nor U6840 (N_6840,N_6746,N_6664);
nand U6841 (N_6841,N_6613,N_6607);
nand U6842 (N_6842,N_6662,N_6732);
nor U6843 (N_6843,N_6680,N_6669);
or U6844 (N_6844,N_6622,N_6681);
or U6845 (N_6845,N_6647,N_6716);
and U6846 (N_6846,N_6616,N_6718);
nand U6847 (N_6847,N_6643,N_6657);
xor U6848 (N_6848,N_6631,N_6689);
nand U6849 (N_6849,N_6640,N_6657);
xor U6850 (N_6850,N_6720,N_6677);
or U6851 (N_6851,N_6674,N_6604);
or U6852 (N_6852,N_6738,N_6604);
and U6853 (N_6853,N_6618,N_6740);
and U6854 (N_6854,N_6649,N_6686);
xor U6855 (N_6855,N_6630,N_6629);
xnor U6856 (N_6856,N_6732,N_6690);
xnor U6857 (N_6857,N_6658,N_6685);
xor U6858 (N_6858,N_6705,N_6616);
xnor U6859 (N_6859,N_6712,N_6696);
xor U6860 (N_6860,N_6708,N_6731);
xor U6861 (N_6861,N_6633,N_6653);
and U6862 (N_6862,N_6729,N_6744);
and U6863 (N_6863,N_6658,N_6713);
xnor U6864 (N_6864,N_6721,N_6732);
or U6865 (N_6865,N_6613,N_6669);
and U6866 (N_6866,N_6729,N_6738);
and U6867 (N_6867,N_6661,N_6617);
and U6868 (N_6868,N_6635,N_6722);
xnor U6869 (N_6869,N_6743,N_6647);
nor U6870 (N_6870,N_6701,N_6600);
and U6871 (N_6871,N_6693,N_6707);
nand U6872 (N_6872,N_6740,N_6655);
xnor U6873 (N_6873,N_6660,N_6739);
or U6874 (N_6874,N_6713,N_6680);
nand U6875 (N_6875,N_6696,N_6689);
nand U6876 (N_6876,N_6621,N_6680);
or U6877 (N_6877,N_6611,N_6746);
nor U6878 (N_6878,N_6633,N_6686);
xor U6879 (N_6879,N_6638,N_6725);
nand U6880 (N_6880,N_6659,N_6635);
or U6881 (N_6881,N_6613,N_6742);
or U6882 (N_6882,N_6635,N_6618);
nor U6883 (N_6883,N_6694,N_6620);
xnor U6884 (N_6884,N_6679,N_6600);
xor U6885 (N_6885,N_6731,N_6652);
xor U6886 (N_6886,N_6635,N_6612);
xnor U6887 (N_6887,N_6690,N_6606);
and U6888 (N_6888,N_6695,N_6600);
nor U6889 (N_6889,N_6635,N_6637);
nor U6890 (N_6890,N_6711,N_6709);
xnor U6891 (N_6891,N_6635,N_6606);
xor U6892 (N_6892,N_6714,N_6739);
nand U6893 (N_6893,N_6690,N_6722);
or U6894 (N_6894,N_6681,N_6719);
nor U6895 (N_6895,N_6686,N_6669);
nand U6896 (N_6896,N_6730,N_6605);
xnor U6897 (N_6897,N_6672,N_6717);
nand U6898 (N_6898,N_6624,N_6721);
nor U6899 (N_6899,N_6660,N_6695);
nor U6900 (N_6900,N_6869,N_6888);
or U6901 (N_6901,N_6863,N_6791);
xnor U6902 (N_6902,N_6872,N_6873);
nand U6903 (N_6903,N_6759,N_6761);
nor U6904 (N_6904,N_6752,N_6851);
or U6905 (N_6905,N_6821,N_6886);
nor U6906 (N_6906,N_6891,N_6878);
or U6907 (N_6907,N_6839,N_6753);
nand U6908 (N_6908,N_6818,N_6892);
nor U6909 (N_6909,N_6853,N_6864);
nand U6910 (N_6910,N_6882,N_6787);
xnor U6911 (N_6911,N_6796,N_6824);
nand U6912 (N_6912,N_6766,N_6849);
and U6913 (N_6913,N_6778,N_6837);
nor U6914 (N_6914,N_6785,N_6825);
nand U6915 (N_6915,N_6842,N_6780);
nand U6916 (N_6916,N_6768,N_6827);
and U6917 (N_6917,N_6846,N_6843);
or U6918 (N_6918,N_6894,N_6845);
nor U6919 (N_6919,N_6893,N_6760);
and U6920 (N_6920,N_6881,N_6838);
or U6921 (N_6921,N_6798,N_6857);
or U6922 (N_6922,N_6833,N_6831);
or U6923 (N_6923,N_6774,N_6899);
xnor U6924 (N_6924,N_6865,N_6754);
xnor U6925 (N_6925,N_6790,N_6871);
xnor U6926 (N_6926,N_6896,N_6793);
or U6927 (N_6927,N_6850,N_6875);
and U6928 (N_6928,N_6777,N_6832);
xnor U6929 (N_6929,N_6884,N_6814);
and U6930 (N_6930,N_6877,N_6804);
or U6931 (N_6931,N_6799,N_6822);
nand U6932 (N_6932,N_6870,N_6756);
xor U6933 (N_6933,N_6826,N_6762);
nor U6934 (N_6934,N_6813,N_6852);
or U6935 (N_6935,N_6823,N_6794);
and U6936 (N_6936,N_6844,N_6854);
xor U6937 (N_6937,N_6786,N_6895);
and U6938 (N_6938,N_6847,N_6859);
xor U6939 (N_6939,N_6763,N_6784);
nor U6940 (N_6940,N_6885,N_6841);
nand U6941 (N_6941,N_6779,N_6755);
nor U6942 (N_6942,N_6806,N_6856);
nor U6943 (N_6943,N_6792,N_6802);
nand U6944 (N_6944,N_6771,N_6770);
and U6945 (N_6945,N_6834,N_6829);
xor U6946 (N_6946,N_6789,N_6758);
xnor U6947 (N_6947,N_6795,N_6889);
nor U6948 (N_6948,N_6751,N_6887);
or U6949 (N_6949,N_6815,N_6890);
nor U6950 (N_6950,N_6874,N_6876);
and U6951 (N_6951,N_6817,N_6880);
xor U6952 (N_6952,N_6830,N_6782);
and U6953 (N_6953,N_6797,N_6775);
xnor U6954 (N_6954,N_6781,N_6767);
or U6955 (N_6955,N_6883,N_6868);
xnor U6956 (N_6956,N_6765,N_6805);
nor U6957 (N_6957,N_6860,N_6879);
nor U6958 (N_6958,N_6858,N_6840);
nand U6959 (N_6959,N_6750,N_6835);
xor U6960 (N_6960,N_6773,N_6803);
xor U6961 (N_6961,N_6855,N_6867);
nand U6962 (N_6962,N_6776,N_6861);
nand U6963 (N_6963,N_6783,N_6800);
xnor U6964 (N_6964,N_6808,N_6816);
or U6965 (N_6965,N_6769,N_6764);
nand U6966 (N_6966,N_6811,N_6812);
and U6967 (N_6967,N_6819,N_6836);
nor U6968 (N_6968,N_6809,N_6772);
xnor U6969 (N_6969,N_6810,N_6820);
nor U6970 (N_6970,N_6866,N_6788);
and U6971 (N_6971,N_6828,N_6862);
nand U6972 (N_6972,N_6757,N_6897);
xnor U6973 (N_6973,N_6807,N_6898);
nor U6974 (N_6974,N_6848,N_6801);
and U6975 (N_6975,N_6867,N_6865);
nand U6976 (N_6976,N_6888,N_6853);
nand U6977 (N_6977,N_6793,N_6795);
nor U6978 (N_6978,N_6844,N_6795);
xor U6979 (N_6979,N_6842,N_6827);
and U6980 (N_6980,N_6823,N_6866);
xnor U6981 (N_6981,N_6836,N_6760);
xor U6982 (N_6982,N_6805,N_6800);
nor U6983 (N_6983,N_6778,N_6871);
xnor U6984 (N_6984,N_6861,N_6844);
nor U6985 (N_6985,N_6798,N_6784);
or U6986 (N_6986,N_6881,N_6812);
xnor U6987 (N_6987,N_6843,N_6895);
nand U6988 (N_6988,N_6797,N_6807);
or U6989 (N_6989,N_6814,N_6811);
nand U6990 (N_6990,N_6815,N_6831);
and U6991 (N_6991,N_6870,N_6814);
xor U6992 (N_6992,N_6819,N_6830);
or U6993 (N_6993,N_6758,N_6819);
and U6994 (N_6994,N_6806,N_6874);
xnor U6995 (N_6995,N_6804,N_6817);
nand U6996 (N_6996,N_6811,N_6877);
and U6997 (N_6997,N_6825,N_6764);
xnor U6998 (N_6998,N_6833,N_6837);
and U6999 (N_6999,N_6809,N_6808);
and U7000 (N_7000,N_6789,N_6771);
xor U7001 (N_7001,N_6860,N_6817);
nand U7002 (N_7002,N_6855,N_6893);
and U7003 (N_7003,N_6792,N_6878);
nand U7004 (N_7004,N_6750,N_6873);
nor U7005 (N_7005,N_6891,N_6888);
nor U7006 (N_7006,N_6863,N_6800);
xnor U7007 (N_7007,N_6765,N_6788);
xnor U7008 (N_7008,N_6761,N_6760);
xnor U7009 (N_7009,N_6878,N_6896);
nor U7010 (N_7010,N_6855,N_6764);
nor U7011 (N_7011,N_6788,N_6843);
nand U7012 (N_7012,N_6789,N_6813);
and U7013 (N_7013,N_6800,N_6834);
nor U7014 (N_7014,N_6803,N_6870);
nor U7015 (N_7015,N_6853,N_6780);
and U7016 (N_7016,N_6838,N_6821);
and U7017 (N_7017,N_6782,N_6770);
xor U7018 (N_7018,N_6866,N_6770);
xor U7019 (N_7019,N_6876,N_6754);
nor U7020 (N_7020,N_6866,N_6829);
nor U7021 (N_7021,N_6847,N_6765);
nor U7022 (N_7022,N_6865,N_6852);
xnor U7023 (N_7023,N_6829,N_6861);
nand U7024 (N_7024,N_6862,N_6829);
nand U7025 (N_7025,N_6862,N_6780);
nand U7026 (N_7026,N_6892,N_6804);
or U7027 (N_7027,N_6774,N_6825);
nand U7028 (N_7028,N_6756,N_6862);
nand U7029 (N_7029,N_6874,N_6784);
and U7030 (N_7030,N_6865,N_6827);
or U7031 (N_7031,N_6887,N_6782);
nor U7032 (N_7032,N_6846,N_6799);
and U7033 (N_7033,N_6834,N_6767);
and U7034 (N_7034,N_6893,N_6807);
or U7035 (N_7035,N_6881,N_6801);
nor U7036 (N_7036,N_6751,N_6834);
xor U7037 (N_7037,N_6820,N_6896);
xor U7038 (N_7038,N_6827,N_6823);
nor U7039 (N_7039,N_6884,N_6813);
nand U7040 (N_7040,N_6831,N_6810);
or U7041 (N_7041,N_6773,N_6840);
xor U7042 (N_7042,N_6876,N_6818);
and U7043 (N_7043,N_6829,N_6843);
xor U7044 (N_7044,N_6895,N_6804);
xnor U7045 (N_7045,N_6882,N_6836);
or U7046 (N_7046,N_6810,N_6891);
nand U7047 (N_7047,N_6766,N_6861);
nand U7048 (N_7048,N_6862,N_6781);
nor U7049 (N_7049,N_6781,N_6844);
nand U7050 (N_7050,N_7006,N_6983);
or U7051 (N_7051,N_6977,N_6991);
nand U7052 (N_7052,N_7035,N_6944);
nand U7053 (N_7053,N_6941,N_6996);
and U7054 (N_7054,N_6945,N_7027);
and U7055 (N_7055,N_7003,N_6910);
nor U7056 (N_7056,N_6971,N_6904);
or U7057 (N_7057,N_7026,N_7032);
or U7058 (N_7058,N_7012,N_6911);
nand U7059 (N_7059,N_7046,N_6921);
or U7060 (N_7060,N_7014,N_6901);
or U7061 (N_7061,N_6962,N_7048);
nor U7062 (N_7062,N_6913,N_7008);
nor U7063 (N_7063,N_7045,N_7038);
and U7064 (N_7064,N_6943,N_6908);
xnor U7065 (N_7065,N_6909,N_6995);
and U7066 (N_7066,N_6939,N_7023);
and U7067 (N_7067,N_6966,N_6975);
or U7068 (N_7068,N_7028,N_6989);
nor U7069 (N_7069,N_6956,N_6917);
and U7070 (N_7070,N_6927,N_6920);
and U7071 (N_7071,N_6999,N_6988);
nand U7072 (N_7072,N_7037,N_6955);
nor U7073 (N_7073,N_6954,N_6923);
xor U7074 (N_7074,N_6970,N_6990);
nor U7075 (N_7075,N_6969,N_7009);
nand U7076 (N_7076,N_7005,N_7019);
xor U7077 (N_7077,N_6902,N_6986);
nor U7078 (N_7078,N_6932,N_6912);
or U7079 (N_7079,N_6918,N_6919);
nor U7080 (N_7080,N_6992,N_6933);
nand U7081 (N_7081,N_6974,N_6905);
xor U7082 (N_7082,N_6931,N_6997);
xor U7083 (N_7083,N_7041,N_6915);
and U7084 (N_7084,N_6935,N_6994);
and U7085 (N_7085,N_6976,N_7030);
nand U7086 (N_7086,N_6948,N_7001);
and U7087 (N_7087,N_6985,N_6914);
xor U7088 (N_7088,N_7020,N_6965);
nor U7089 (N_7089,N_6967,N_6903);
nand U7090 (N_7090,N_6978,N_6916);
nand U7091 (N_7091,N_7047,N_7024);
nor U7092 (N_7092,N_7021,N_6934);
or U7093 (N_7093,N_7011,N_6957);
nor U7094 (N_7094,N_7049,N_6942);
xor U7095 (N_7095,N_7036,N_6964);
xnor U7096 (N_7096,N_7013,N_6924);
and U7097 (N_7097,N_7034,N_6963);
nand U7098 (N_7098,N_6960,N_6925);
or U7099 (N_7099,N_6984,N_7010);
xor U7100 (N_7100,N_6900,N_6952);
nor U7101 (N_7101,N_6993,N_7022);
xnor U7102 (N_7102,N_6949,N_7017);
nand U7103 (N_7103,N_6946,N_6998);
nand U7104 (N_7104,N_6922,N_6930);
xnor U7105 (N_7105,N_7031,N_6982);
and U7106 (N_7106,N_6929,N_6938);
or U7107 (N_7107,N_7018,N_7040);
xor U7108 (N_7108,N_6959,N_7025);
and U7109 (N_7109,N_7039,N_7007);
nor U7110 (N_7110,N_7000,N_6961);
nand U7111 (N_7111,N_6987,N_6958);
and U7112 (N_7112,N_6981,N_6979);
nor U7113 (N_7113,N_6973,N_7033);
nand U7114 (N_7114,N_7015,N_6980);
nand U7115 (N_7115,N_6951,N_7044);
nand U7116 (N_7116,N_6950,N_7029);
and U7117 (N_7117,N_6926,N_6906);
and U7118 (N_7118,N_6947,N_6940);
nand U7119 (N_7119,N_6972,N_6907);
and U7120 (N_7120,N_7004,N_6968);
xor U7121 (N_7121,N_7016,N_6936);
nand U7122 (N_7122,N_7043,N_7002);
nand U7123 (N_7123,N_6928,N_6937);
nand U7124 (N_7124,N_6953,N_7042);
nor U7125 (N_7125,N_7048,N_7023);
and U7126 (N_7126,N_6965,N_6922);
or U7127 (N_7127,N_7029,N_6983);
and U7128 (N_7128,N_7026,N_6985);
or U7129 (N_7129,N_6970,N_6980);
nand U7130 (N_7130,N_7030,N_7016);
nand U7131 (N_7131,N_7013,N_6981);
nor U7132 (N_7132,N_7018,N_6974);
nand U7133 (N_7133,N_6909,N_6924);
or U7134 (N_7134,N_6931,N_7039);
or U7135 (N_7135,N_6978,N_7043);
nand U7136 (N_7136,N_7019,N_7004);
or U7137 (N_7137,N_6940,N_7034);
xor U7138 (N_7138,N_7027,N_6928);
nor U7139 (N_7139,N_7035,N_7016);
or U7140 (N_7140,N_6993,N_6952);
xnor U7141 (N_7141,N_6945,N_7029);
nand U7142 (N_7142,N_6990,N_6907);
xor U7143 (N_7143,N_6924,N_6955);
nand U7144 (N_7144,N_6926,N_6913);
and U7145 (N_7145,N_7000,N_6997);
xor U7146 (N_7146,N_6998,N_7021);
nand U7147 (N_7147,N_6968,N_6986);
or U7148 (N_7148,N_6984,N_7018);
xor U7149 (N_7149,N_7024,N_6943);
and U7150 (N_7150,N_7001,N_6908);
or U7151 (N_7151,N_6912,N_6988);
and U7152 (N_7152,N_7013,N_6997);
nand U7153 (N_7153,N_6993,N_7016);
and U7154 (N_7154,N_6937,N_6906);
nand U7155 (N_7155,N_6962,N_6917);
xor U7156 (N_7156,N_6987,N_6952);
and U7157 (N_7157,N_6904,N_6972);
nor U7158 (N_7158,N_7007,N_6970);
xor U7159 (N_7159,N_6962,N_6926);
and U7160 (N_7160,N_6957,N_7023);
or U7161 (N_7161,N_7040,N_6967);
and U7162 (N_7162,N_6981,N_7043);
and U7163 (N_7163,N_6931,N_6935);
nand U7164 (N_7164,N_7047,N_6919);
or U7165 (N_7165,N_6964,N_6966);
nand U7166 (N_7166,N_6955,N_6991);
and U7167 (N_7167,N_6977,N_6995);
xor U7168 (N_7168,N_7004,N_6925);
and U7169 (N_7169,N_6902,N_6908);
or U7170 (N_7170,N_7004,N_6988);
nand U7171 (N_7171,N_6923,N_6953);
xnor U7172 (N_7172,N_6998,N_7024);
nor U7173 (N_7173,N_6926,N_7012);
nor U7174 (N_7174,N_6983,N_6978);
or U7175 (N_7175,N_6992,N_6972);
xor U7176 (N_7176,N_6965,N_7010);
nor U7177 (N_7177,N_6944,N_7003);
nor U7178 (N_7178,N_7027,N_6983);
or U7179 (N_7179,N_7048,N_7028);
xor U7180 (N_7180,N_6906,N_7038);
and U7181 (N_7181,N_6985,N_6910);
nand U7182 (N_7182,N_6920,N_6948);
xor U7183 (N_7183,N_7023,N_6906);
and U7184 (N_7184,N_7031,N_7016);
xnor U7185 (N_7185,N_6951,N_6919);
nand U7186 (N_7186,N_6930,N_7044);
or U7187 (N_7187,N_7021,N_6938);
and U7188 (N_7188,N_6947,N_6936);
nor U7189 (N_7189,N_7035,N_7037);
xor U7190 (N_7190,N_6935,N_7030);
nor U7191 (N_7191,N_6941,N_7035);
or U7192 (N_7192,N_7045,N_6948);
xor U7193 (N_7193,N_6928,N_7039);
and U7194 (N_7194,N_6919,N_6907);
nand U7195 (N_7195,N_6962,N_6980);
and U7196 (N_7196,N_6980,N_6932);
and U7197 (N_7197,N_6901,N_6915);
xnor U7198 (N_7198,N_6998,N_7045);
nand U7199 (N_7199,N_7039,N_6942);
nand U7200 (N_7200,N_7070,N_7170);
or U7201 (N_7201,N_7182,N_7116);
nand U7202 (N_7202,N_7159,N_7060);
nand U7203 (N_7203,N_7191,N_7168);
xor U7204 (N_7204,N_7066,N_7096);
nor U7205 (N_7205,N_7197,N_7097);
or U7206 (N_7206,N_7064,N_7076);
nand U7207 (N_7207,N_7089,N_7117);
nor U7208 (N_7208,N_7156,N_7124);
nand U7209 (N_7209,N_7147,N_7186);
or U7210 (N_7210,N_7119,N_7052);
or U7211 (N_7211,N_7100,N_7106);
or U7212 (N_7212,N_7166,N_7071);
nor U7213 (N_7213,N_7139,N_7189);
nor U7214 (N_7214,N_7199,N_7181);
nand U7215 (N_7215,N_7132,N_7144);
and U7216 (N_7216,N_7127,N_7152);
and U7217 (N_7217,N_7148,N_7057);
or U7218 (N_7218,N_7172,N_7056);
or U7219 (N_7219,N_7184,N_7082);
xnor U7220 (N_7220,N_7173,N_7098);
nor U7221 (N_7221,N_7088,N_7169);
nor U7222 (N_7222,N_7180,N_7190);
and U7223 (N_7223,N_7069,N_7142);
nand U7224 (N_7224,N_7151,N_7175);
or U7225 (N_7225,N_7154,N_7095);
nor U7226 (N_7226,N_7185,N_7053);
or U7227 (N_7227,N_7103,N_7080);
nor U7228 (N_7228,N_7062,N_7171);
or U7229 (N_7229,N_7155,N_7178);
nor U7230 (N_7230,N_7113,N_7105);
or U7231 (N_7231,N_7065,N_7091);
or U7232 (N_7232,N_7129,N_7087);
and U7233 (N_7233,N_7051,N_7101);
or U7234 (N_7234,N_7090,N_7196);
xor U7235 (N_7235,N_7143,N_7109);
or U7236 (N_7236,N_7141,N_7108);
nor U7237 (N_7237,N_7121,N_7137);
nand U7238 (N_7238,N_7192,N_7164);
nor U7239 (N_7239,N_7114,N_7162);
nand U7240 (N_7240,N_7187,N_7110);
nand U7241 (N_7241,N_7094,N_7093);
nand U7242 (N_7242,N_7118,N_7149);
or U7243 (N_7243,N_7134,N_7150);
nor U7244 (N_7244,N_7084,N_7138);
nand U7245 (N_7245,N_7059,N_7061);
xnor U7246 (N_7246,N_7183,N_7167);
or U7247 (N_7247,N_7058,N_7067);
xor U7248 (N_7248,N_7068,N_7160);
nand U7249 (N_7249,N_7086,N_7195);
or U7250 (N_7250,N_7165,N_7072);
nor U7251 (N_7251,N_7085,N_7133);
or U7252 (N_7252,N_7081,N_7158);
xor U7253 (N_7253,N_7188,N_7079);
or U7254 (N_7254,N_7115,N_7145);
nor U7255 (N_7255,N_7163,N_7128);
or U7256 (N_7256,N_7077,N_7140);
or U7257 (N_7257,N_7126,N_7107);
or U7258 (N_7258,N_7123,N_7157);
and U7259 (N_7259,N_7111,N_7161);
nor U7260 (N_7260,N_7130,N_7153);
xor U7261 (N_7261,N_7125,N_7146);
nand U7262 (N_7262,N_7078,N_7092);
nand U7263 (N_7263,N_7174,N_7177);
xor U7264 (N_7264,N_7194,N_7193);
and U7265 (N_7265,N_7102,N_7135);
or U7266 (N_7266,N_7055,N_7179);
or U7267 (N_7267,N_7120,N_7136);
or U7268 (N_7268,N_7073,N_7075);
and U7269 (N_7269,N_7112,N_7054);
xnor U7270 (N_7270,N_7074,N_7050);
nand U7271 (N_7271,N_7099,N_7063);
and U7272 (N_7272,N_7122,N_7176);
or U7273 (N_7273,N_7083,N_7104);
nand U7274 (N_7274,N_7131,N_7198);
and U7275 (N_7275,N_7100,N_7165);
and U7276 (N_7276,N_7109,N_7194);
xnor U7277 (N_7277,N_7134,N_7187);
xor U7278 (N_7278,N_7053,N_7154);
xnor U7279 (N_7279,N_7140,N_7084);
or U7280 (N_7280,N_7104,N_7094);
xor U7281 (N_7281,N_7157,N_7180);
xnor U7282 (N_7282,N_7126,N_7087);
and U7283 (N_7283,N_7065,N_7051);
nor U7284 (N_7284,N_7148,N_7072);
and U7285 (N_7285,N_7142,N_7166);
xor U7286 (N_7286,N_7107,N_7078);
and U7287 (N_7287,N_7131,N_7173);
or U7288 (N_7288,N_7091,N_7068);
and U7289 (N_7289,N_7135,N_7069);
and U7290 (N_7290,N_7103,N_7079);
xnor U7291 (N_7291,N_7112,N_7192);
nand U7292 (N_7292,N_7067,N_7110);
and U7293 (N_7293,N_7068,N_7192);
nand U7294 (N_7294,N_7147,N_7199);
and U7295 (N_7295,N_7149,N_7068);
xor U7296 (N_7296,N_7186,N_7089);
and U7297 (N_7297,N_7123,N_7103);
nand U7298 (N_7298,N_7103,N_7161);
nor U7299 (N_7299,N_7075,N_7185);
nand U7300 (N_7300,N_7151,N_7108);
or U7301 (N_7301,N_7177,N_7175);
nor U7302 (N_7302,N_7119,N_7173);
nor U7303 (N_7303,N_7098,N_7053);
xnor U7304 (N_7304,N_7107,N_7108);
and U7305 (N_7305,N_7176,N_7149);
nor U7306 (N_7306,N_7153,N_7068);
and U7307 (N_7307,N_7072,N_7180);
or U7308 (N_7308,N_7071,N_7092);
and U7309 (N_7309,N_7106,N_7151);
nand U7310 (N_7310,N_7161,N_7098);
xnor U7311 (N_7311,N_7054,N_7150);
nor U7312 (N_7312,N_7182,N_7172);
or U7313 (N_7313,N_7061,N_7108);
nand U7314 (N_7314,N_7078,N_7186);
or U7315 (N_7315,N_7136,N_7063);
or U7316 (N_7316,N_7075,N_7107);
and U7317 (N_7317,N_7142,N_7083);
nand U7318 (N_7318,N_7185,N_7116);
nand U7319 (N_7319,N_7166,N_7162);
nand U7320 (N_7320,N_7190,N_7072);
nor U7321 (N_7321,N_7186,N_7080);
or U7322 (N_7322,N_7161,N_7087);
nor U7323 (N_7323,N_7098,N_7174);
or U7324 (N_7324,N_7197,N_7050);
xnor U7325 (N_7325,N_7074,N_7105);
xnor U7326 (N_7326,N_7140,N_7120);
and U7327 (N_7327,N_7099,N_7196);
xnor U7328 (N_7328,N_7116,N_7082);
xor U7329 (N_7329,N_7102,N_7068);
nor U7330 (N_7330,N_7060,N_7122);
and U7331 (N_7331,N_7053,N_7123);
and U7332 (N_7332,N_7067,N_7136);
or U7333 (N_7333,N_7105,N_7199);
nand U7334 (N_7334,N_7194,N_7172);
xor U7335 (N_7335,N_7060,N_7192);
xnor U7336 (N_7336,N_7163,N_7164);
and U7337 (N_7337,N_7142,N_7087);
xnor U7338 (N_7338,N_7178,N_7140);
nand U7339 (N_7339,N_7160,N_7138);
nor U7340 (N_7340,N_7172,N_7074);
nor U7341 (N_7341,N_7133,N_7152);
or U7342 (N_7342,N_7059,N_7145);
xnor U7343 (N_7343,N_7144,N_7168);
nand U7344 (N_7344,N_7143,N_7083);
or U7345 (N_7345,N_7151,N_7058);
and U7346 (N_7346,N_7088,N_7198);
xnor U7347 (N_7347,N_7063,N_7092);
nor U7348 (N_7348,N_7189,N_7146);
nand U7349 (N_7349,N_7082,N_7064);
and U7350 (N_7350,N_7206,N_7246);
or U7351 (N_7351,N_7287,N_7301);
xnor U7352 (N_7352,N_7336,N_7327);
nor U7353 (N_7353,N_7255,N_7340);
nor U7354 (N_7354,N_7207,N_7305);
nor U7355 (N_7355,N_7330,N_7347);
nand U7356 (N_7356,N_7284,N_7236);
xnor U7357 (N_7357,N_7277,N_7319);
nor U7358 (N_7358,N_7219,N_7223);
nand U7359 (N_7359,N_7315,N_7225);
and U7360 (N_7360,N_7292,N_7276);
and U7361 (N_7361,N_7263,N_7211);
and U7362 (N_7362,N_7239,N_7249);
xnor U7363 (N_7363,N_7273,N_7346);
nand U7364 (N_7364,N_7215,N_7325);
xor U7365 (N_7365,N_7266,N_7308);
or U7366 (N_7366,N_7250,N_7238);
and U7367 (N_7367,N_7203,N_7261);
nand U7368 (N_7368,N_7201,N_7312);
nor U7369 (N_7369,N_7326,N_7200);
nor U7370 (N_7370,N_7258,N_7221);
nand U7371 (N_7371,N_7322,N_7316);
xnor U7372 (N_7372,N_7279,N_7232);
nand U7373 (N_7373,N_7264,N_7290);
and U7374 (N_7374,N_7245,N_7256);
or U7375 (N_7375,N_7222,N_7304);
and U7376 (N_7376,N_7293,N_7289);
xnor U7377 (N_7377,N_7220,N_7295);
and U7378 (N_7378,N_7229,N_7237);
xor U7379 (N_7379,N_7260,N_7345);
or U7380 (N_7380,N_7343,N_7265);
or U7381 (N_7381,N_7339,N_7328);
xor U7382 (N_7382,N_7333,N_7297);
xor U7383 (N_7383,N_7280,N_7311);
xor U7384 (N_7384,N_7349,N_7224);
or U7385 (N_7385,N_7252,N_7240);
nor U7386 (N_7386,N_7303,N_7272);
and U7387 (N_7387,N_7248,N_7348);
nor U7388 (N_7388,N_7257,N_7204);
and U7389 (N_7389,N_7213,N_7313);
and U7390 (N_7390,N_7323,N_7334);
nor U7391 (N_7391,N_7228,N_7331);
nand U7392 (N_7392,N_7341,N_7282);
nor U7393 (N_7393,N_7278,N_7259);
and U7394 (N_7394,N_7298,N_7318);
nand U7395 (N_7395,N_7332,N_7244);
xnor U7396 (N_7396,N_7217,N_7226);
and U7397 (N_7397,N_7216,N_7214);
or U7398 (N_7398,N_7314,N_7281);
xor U7399 (N_7399,N_7247,N_7306);
nor U7400 (N_7400,N_7231,N_7253);
nor U7401 (N_7401,N_7242,N_7267);
xor U7402 (N_7402,N_7294,N_7243);
nor U7403 (N_7403,N_7210,N_7235);
xor U7404 (N_7404,N_7274,N_7302);
nor U7405 (N_7405,N_7309,N_7342);
or U7406 (N_7406,N_7310,N_7251);
and U7407 (N_7407,N_7291,N_7254);
and U7408 (N_7408,N_7275,N_7208);
xnor U7409 (N_7409,N_7283,N_7209);
nand U7410 (N_7410,N_7288,N_7285);
nor U7411 (N_7411,N_7218,N_7230);
and U7412 (N_7412,N_7317,N_7286);
nor U7413 (N_7413,N_7205,N_7241);
xnor U7414 (N_7414,N_7268,N_7338);
nor U7415 (N_7415,N_7212,N_7300);
or U7416 (N_7416,N_7329,N_7202);
nor U7417 (N_7417,N_7344,N_7321);
xor U7418 (N_7418,N_7227,N_7324);
nor U7419 (N_7419,N_7307,N_7269);
nand U7420 (N_7420,N_7335,N_7262);
xnor U7421 (N_7421,N_7299,N_7270);
nand U7422 (N_7422,N_7271,N_7337);
and U7423 (N_7423,N_7233,N_7296);
xnor U7424 (N_7424,N_7234,N_7320);
nand U7425 (N_7425,N_7294,N_7317);
nor U7426 (N_7426,N_7343,N_7295);
nor U7427 (N_7427,N_7299,N_7265);
xnor U7428 (N_7428,N_7312,N_7276);
and U7429 (N_7429,N_7260,N_7218);
nand U7430 (N_7430,N_7220,N_7322);
nor U7431 (N_7431,N_7240,N_7345);
and U7432 (N_7432,N_7261,N_7279);
and U7433 (N_7433,N_7290,N_7258);
nor U7434 (N_7434,N_7229,N_7248);
nor U7435 (N_7435,N_7249,N_7200);
nor U7436 (N_7436,N_7249,N_7228);
or U7437 (N_7437,N_7312,N_7323);
or U7438 (N_7438,N_7305,N_7270);
or U7439 (N_7439,N_7234,N_7271);
nand U7440 (N_7440,N_7277,N_7230);
nor U7441 (N_7441,N_7252,N_7248);
and U7442 (N_7442,N_7223,N_7249);
nor U7443 (N_7443,N_7345,N_7257);
or U7444 (N_7444,N_7323,N_7296);
or U7445 (N_7445,N_7307,N_7239);
and U7446 (N_7446,N_7279,N_7275);
nand U7447 (N_7447,N_7235,N_7300);
and U7448 (N_7448,N_7270,N_7240);
or U7449 (N_7449,N_7264,N_7253);
and U7450 (N_7450,N_7304,N_7311);
nand U7451 (N_7451,N_7230,N_7219);
nand U7452 (N_7452,N_7277,N_7297);
or U7453 (N_7453,N_7267,N_7257);
nand U7454 (N_7454,N_7201,N_7299);
xnor U7455 (N_7455,N_7347,N_7340);
nor U7456 (N_7456,N_7347,N_7221);
and U7457 (N_7457,N_7270,N_7282);
nand U7458 (N_7458,N_7295,N_7227);
xor U7459 (N_7459,N_7334,N_7345);
or U7460 (N_7460,N_7200,N_7313);
nand U7461 (N_7461,N_7316,N_7295);
and U7462 (N_7462,N_7348,N_7227);
xor U7463 (N_7463,N_7207,N_7240);
nor U7464 (N_7464,N_7235,N_7261);
nand U7465 (N_7465,N_7333,N_7215);
or U7466 (N_7466,N_7307,N_7302);
or U7467 (N_7467,N_7309,N_7267);
nand U7468 (N_7468,N_7339,N_7218);
and U7469 (N_7469,N_7204,N_7311);
xnor U7470 (N_7470,N_7281,N_7263);
nand U7471 (N_7471,N_7278,N_7214);
or U7472 (N_7472,N_7339,N_7216);
xor U7473 (N_7473,N_7326,N_7279);
and U7474 (N_7474,N_7216,N_7321);
xor U7475 (N_7475,N_7329,N_7309);
nand U7476 (N_7476,N_7316,N_7235);
nand U7477 (N_7477,N_7248,N_7211);
and U7478 (N_7478,N_7279,N_7227);
xor U7479 (N_7479,N_7200,N_7218);
and U7480 (N_7480,N_7311,N_7248);
and U7481 (N_7481,N_7271,N_7270);
and U7482 (N_7482,N_7310,N_7211);
or U7483 (N_7483,N_7290,N_7242);
nor U7484 (N_7484,N_7325,N_7262);
and U7485 (N_7485,N_7252,N_7295);
xnor U7486 (N_7486,N_7234,N_7201);
or U7487 (N_7487,N_7303,N_7321);
xor U7488 (N_7488,N_7255,N_7311);
nor U7489 (N_7489,N_7242,N_7322);
and U7490 (N_7490,N_7211,N_7284);
xor U7491 (N_7491,N_7305,N_7234);
nand U7492 (N_7492,N_7317,N_7333);
nand U7493 (N_7493,N_7342,N_7254);
or U7494 (N_7494,N_7236,N_7318);
or U7495 (N_7495,N_7339,N_7268);
nand U7496 (N_7496,N_7317,N_7298);
xnor U7497 (N_7497,N_7325,N_7257);
nor U7498 (N_7498,N_7267,N_7234);
nand U7499 (N_7499,N_7279,N_7327);
nand U7500 (N_7500,N_7470,N_7459);
nor U7501 (N_7501,N_7353,N_7465);
nand U7502 (N_7502,N_7441,N_7351);
and U7503 (N_7503,N_7363,N_7488);
nand U7504 (N_7504,N_7395,N_7359);
nand U7505 (N_7505,N_7388,N_7498);
nand U7506 (N_7506,N_7385,N_7397);
nor U7507 (N_7507,N_7489,N_7439);
nor U7508 (N_7508,N_7497,N_7361);
nor U7509 (N_7509,N_7383,N_7375);
nand U7510 (N_7510,N_7362,N_7421);
nand U7511 (N_7511,N_7446,N_7356);
or U7512 (N_7512,N_7391,N_7409);
xor U7513 (N_7513,N_7437,N_7453);
nand U7514 (N_7514,N_7467,N_7378);
xor U7515 (N_7515,N_7476,N_7430);
xor U7516 (N_7516,N_7457,N_7433);
and U7517 (N_7517,N_7496,N_7486);
xor U7518 (N_7518,N_7412,N_7364);
xnor U7519 (N_7519,N_7490,N_7404);
nand U7520 (N_7520,N_7456,N_7398);
xnor U7521 (N_7521,N_7352,N_7425);
and U7522 (N_7522,N_7464,N_7394);
and U7523 (N_7523,N_7389,N_7436);
nand U7524 (N_7524,N_7372,N_7402);
and U7525 (N_7525,N_7451,N_7387);
nor U7526 (N_7526,N_7405,N_7367);
or U7527 (N_7527,N_7481,N_7458);
or U7528 (N_7528,N_7358,N_7382);
nor U7529 (N_7529,N_7473,N_7444);
or U7530 (N_7530,N_7392,N_7472);
xnor U7531 (N_7531,N_7354,N_7493);
nand U7532 (N_7532,N_7499,N_7494);
nor U7533 (N_7533,N_7450,N_7460);
nand U7534 (N_7534,N_7483,N_7366);
or U7535 (N_7535,N_7442,N_7475);
nor U7536 (N_7536,N_7379,N_7374);
and U7537 (N_7537,N_7403,N_7380);
nor U7538 (N_7538,N_7357,N_7373);
nand U7539 (N_7539,N_7399,N_7360);
xor U7540 (N_7540,N_7365,N_7484);
or U7541 (N_7541,N_7396,N_7455);
nor U7542 (N_7542,N_7381,N_7393);
nand U7543 (N_7543,N_7447,N_7370);
nor U7544 (N_7544,N_7407,N_7369);
xor U7545 (N_7545,N_7432,N_7478);
xnor U7546 (N_7546,N_7461,N_7415);
nand U7547 (N_7547,N_7435,N_7401);
nor U7548 (N_7548,N_7406,N_7449);
nand U7549 (N_7549,N_7452,N_7418);
nand U7550 (N_7550,N_7386,N_7428);
and U7551 (N_7551,N_7424,N_7376);
nor U7552 (N_7552,N_7384,N_7423);
or U7553 (N_7553,N_7371,N_7474);
xnor U7554 (N_7554,N_7426,N_7411);
and U7555 (N_7555,N_7482,N_7438);
nand U7556 (N_7556,N_7477,N_7480);
and U7557 (N_7557,N_7468,N_7491);
nand U7558 (N_7558,N_7408,N_7390);
nand U7559 (N_7559,N_7434,N_7419);
nor U7560 (N_7560,N_7487,N_7410);
nor U7561 (N_7561,N_7427,N_7417);
or U7562 (N_7562,N_7443,N_7422);
and U7563 (N_7563,N_7355,N_7448);
nor U7564 (N_7564,N_7413,N_7454);
and U7565 (N_7565,N_7416,N_7462);
xor U7566 (N_7566,N_7414,N_7492);
nand U7567 (N_7567,N_7420,N_7429);
or U7568 (N_7568,N_7377,N_7469);
nor U7569 (N_7569,N_7471,N_7440);
or U7570 (N_7570,N_7431,N_7350);
nor U7571 (N_7571,N_7466,N_7479);
and U7572 (N_7572,N_7368,N_7495);
nor U7573 (N_7573,N_7463,N_7445);
nor U7574 (N_7574,N_7400,N_7485);
nand U7575 (N_7575,N_7483,N_7494);
and U7576 (N_7576,N_7460,N_7437);
nand U7577 (N_7577,N_7402,N_7379);
nor U7578 (N_7578,N_7488,N_7357);
nor U7579 (N_7579,N_7350,N_7398);
and U7580 (N_7580,N_7405,N_7446);
or U7581 (N_7581,N_7477,N_7468);
xnor U7582 (N_7582,N_7422,N_7393);
xor U7583 (N_7583,N_7431,N_7379);
and U7584 (N_7584,N_7468,N_7376);
xnor U7585 (N_7585,N_7396,N_7375);
xnor U7586 (N_7586,N_7379,N_7403);
nand U7587 (N_7587,N_7481,N_7426);
xnor U7588 (N_7588,N_7474,N_7356);
nand U7589 (N_7589,N_7369,N_7415);
nor U7590 (N_7590,N_7430,N_7433);
and U7591 (N_7591,N_7493,N_7442);
xor U7592 (N_7592,N_7470,N_7408);
nand U7593 (N_7593,N_7459,N_7422);
or U7594 (N_7594,N_7489,N_7420);
nor U7595 (N_7595,N_7354,N_7361);
nand U7596 (N_7596,N_7373,N_7467);
nand U7597 (N_7597,N_7381,N_7456);
xnor U7598 (N_7598,N_7390,N_7374);
nor U7599 (N_7599,N_7418,N_7421);
or U7600 (N_7600,N_7418,N_7435);
or U7601 (N_7601,N_7388,N_7427);
xnor U7602 (N_7602,N_7412,N_7419);
nand U7603 (N_7603,N_7450,N_7363);
nor U7604 (N_7604,N_7439,N_7469);
nand U7605 (N_7605,N_7451,N_7492);
nand U7606 (N_7606,N_7376,N_7370);
nor U7607 (N_7607,N_7448,N_7456);
xor U7608 (N_7608,N_7382,N_7480);
xnor U7609 (N_7609,N_7361,N_7449);
nor U7610 (N_7610,N_7377,N_7490);
nand U7611 (N_7611,N_7373,N_7380);
and U7612 (N_7612,N_7369,N_7449);
xor U7613 (N_7613,N_7479,N_7434);
and U7614 (N_7614,N_7377,N_7494);
xnor U7615 (N_7615,N_7498,N_7453);
nand U7616 (N_7616,N_7399,N_7410);
xnor U7617 (N_7617,N_7391,N_7414);
nor U7618 (N_7618,N_7404,N_7374);
nand U7619 (N_7619,N_7499,N_7401);
and U7620 (N_7620,N_7363,N_7405);
nor U7621 (N_7621,N_7391,N_7371);
or U7622 (N_7622,N_7374,N_7488);
xnor U7623 (N_7623,N_7403,N_7456);
nor U7624 (N_7624,N_7442,N_7372);
and U7625 (N_7625,N_7426,N_7381);
and U7626 (N_7626,N_7443,N_7406);
nor U7627 (N_7627,N_7351,N_7439);
nor U7628 (N_7628,N_7381,N_7391);
and U7629 (N_7629,N_7390,N_7495);
or U7630 (N_7630,N_7413,N_7435);
or U7631 (N_7631,N_7459,N_7452);
nand U7632 (N_7632,N_7447,N_7401);
xnor U7633 (N_7633,N_7442,N_7476);
xor U7634 (N_7634,N_7350,N_7443);
nand U7635 (N_7635,N_7467,N_7470);
nand U7636 (N_7636,N_7353,N_7406);
xor U7637 (N_7637,N_7402,N_7388);
nand U7638 (N_7638,N_7392,N_7459);
nand U7639 (N_7639,N_7370,N_7363);
and U7640 (N_7640,N_7393,N_7455);
or U7641 (N_7641,N_7496,N_7360);
and U7642 (N_7642,N_7401,N_7393);
nand U7643 (N_7643,N_7363,N_7470);
nand U7644 (N_7644,N_7445,N_7428);
nor U7645 (N_7645,N_7484,N_7392);
or U7646 (N_7646,N_7409,N_7399);
xnor U7647 (N_7647,N_7374,N_7494);
nor U7648 (N_7648,N_7378,N_7460);
or U7649 (N_7649,N_7475,N_7362);
nor U7650 (N_7650,N_7601,N_7620);
and U7651 (N_7651,N_7591,N_7501);
or U7652 (N_7652,N_7535,N_7608);
nand U7653 (N_7653,N_7597,N_7534);
xnor U7654 (N_7654,N_7648,N_7632);
nand U7655 (N_7655,N_7506,N_7546);
and U7656 (N_7656,N_7512,N_7555);
nand U7657 (N_7657,N_7614,N_7611);
nor U7658 (N_7658,N_7631,N_7602);
xor U7659 (N_7659,N_7500,N_7539);
nor U7660 (N_7660,N_7531,N_7638);
nand U7661 (N_7661,N_7626,N_7515);
or U7662 (N_7662,N_7634,N_7503);
nand U7663 (N_7663,N_7587,N_7550);
nor U7664 (N_7664,N_7538,N_7599);
xor U7665 (N_7665,N_7572,N_7507);
or U7666 (N_7666,N_7580,N_7577);
nor U7667 (N_7667,N_7588,N_7551);
or U7668 (N_7668,N_7606,N_7504);
xnor U7669 (N_7669,N_7524,N_7583);
or U7670 (N_7670,N_7543,N_7610);
nand U7671 (N_7671,N_7519,N_7568);
or U7672 (N_7672,N_7645,N_7629);
nor U7673 (N_7673,N_7537,N_7624);
and U7674 (N_7674,N_7574,N_7590);
and U7675 (N_7675,N_7511,N_7604);
and U7676 (N_7676,N_7526,N_7544);
nand U7677 (N_7677,N_7522,N_7529);
xnor U7678 (N_7678,N_7617,N_7554);
and U7679 (N_7679,N_7613,N_7567);
nor U7680 (N_7680,N_7510,N_7532);
nor U7681 (N_7681,N_7513,N_7561);
nand U7682 (N_7682,N_7582,N_7641);
or U7683 (N_7683,N_7558,N_7563);
or U7684 (N_7684,N_7553,N_7576);
and U7685 (N_7685,N_7585,N_7622);
nand U7686 (N_7686,N_7605,N_7592);
and U7687 (N_7687,N_7518,N_7616);
and U7688 (N_7688,N_7649,N_7565);
xnor U7689 (N_7689,N_7578,N_7584);
or U7690 (N_7690,N_7628,N_7566);
nand U7691 (N_7691,N_7644,N_7533);
nor U7692 (N_7692,N_7603,N_7593);
nor U7693 (N_7693,N_7502,N_7530);
xnor U7694 (N_7694,N_7564,N_7623);
nor U7695 (N_7695,N_7545,N_7523);
xor U7696 (N_7696,N_7505,N_7625);
nand U7697 (N_7697,N_7594,N_7619);
or U7698 (N_7698,N_7596,N_7621);
or U7699 (N_7699,N_7536,N_7633);
or U7700 (N_7700,N_7639,N_7547);
xnor U7701 (N_7701,N_7571,N_7548);
or U7702 (N_7702,N_7540,N_7595);
nand U7703 (N_7703,N_7630,N_7559);
nand U7704 (N_7704,N_7586,N_7521);
or U7705 (N_7705,N_7525,N_7579);
xnor U7706 (N_7706,N_7573,N_7570);
nor U7707 (N_7707,N_7643,N_7509);
xor U7708 (N_7708,N_7635,N_7647);
and U7709 (N_7709,N_7642,N_7636);
nor U7710 (N_7710,N_7607,N_7560);
xnor U7711 (N_7711,N_7589,N_7556);
or U7712 (N_7712,N_7562,N_7609);
nand U7713 (N_7713,N_7508,N_7520);
nor U7714 (N_7714,N_7514,N_7517);
nand U7715 (N_7715,N_7615,N_7627);
xnor U7716 (N_7716,N_7581,N_7552);
xnor U7717 (N_7717,N_7637,N_7598);
xnor U7718 (N_7718,N_7612,N_7575);
or U7719 (N_7719,N_7600,N_7542);
nor U7720 (N_7720,N_7557,N_7549);
or U7721 (N_7721,N_7528,N_7640);
nor U7722 (N_7722,N_7541,N_7646);
nand U7723 (N_7723,N_7516,N_7527);
or U7724 (N_7724,N_7569,N_7618);
nor U7725 (N_7725,N_7560,N_7614);
and U7726 (N_7726,N_7625,N_7581);
and U7727 (N_7727,N_7574,N_7609);
or U7728 (N_7728,N_7561,N_7505);
nand U7729 (N_7729,N_7516,N_7500);
and U7730 (N_7730,N_7550,N_7538);
and U7731 (N_7731,N_7566,N_7526);
or U7732 (N_7732,N_7565,N_7563);
nor U7733 (N_7733,N_7572,N_7598);
nor U7734 (N_7734,N_7595,N_7640);
xnor U7735 (N_7735,N_7632,N_7523);
xnor U7736 (N_7736,N_7536,N_7572);
and U7737 (N_7737,N_7586,N_7562);
nand U7738 (N_7738,N_7616,N_7559);
nand U7739 (N_7739,N_7556,N_7535);
nor U7740 (N_7740,N_7626,N_7509);
nand U7741 (N_7741,N_7580,N_7560);
nand U7742 (N_7742,N_7605,N_7563);
or U7743 (N_7743,N_7512,N_7591);
xnor U7744 (N_7744,N_7541,N_7613);
or U7745 (N_7745,N_7585,N_7649);
nand U7746 (N_7746,N_7604,N_7536);
xnor U7747 (N_7747,N_7640,N_7624);
nand U7748 (N_7748,N_7533,N_7572);
or U7749 (N_7749,N_7580,N_7537);
nand U7750 (N_7750,N_7583,N_7594);
xnor U7751 (N_7751,N_7553,N_7535);
nand U7752 (N_7752,N_7646,N_7501);
xnor U7753 (N_7753,N_7600,N_7562);
or U7754 (N_7754,N_7594,N_7579);
and U7755 (N_7755,N_7557,N_7626);
xor U7756 (N_7756,N_7570,N_7506);
and U7757 (N_7757,N_7560,N_7539);
and U7758 (N_7758,N_7505,N_7539);
xor U7759 (N_7759,N_7554,N_7513);
xor U7760 (N_7760,N_7647,N_7519);
nand U7761 (N_7761,N_7524,N_7543);
and U7762 (N_7762,N_7613,N_7555);
xor U7763 (N_7763,N_7516,N_7610);
xor U7764 (N_7764,N_7606,N_7563);
or U7765 (N_7765,N_7535,N_7636);
nor U7766 (N_7766,N_7569,N_7557);
and U7767 (N_7767,N_7624,N_7507);
nor U7768 (N_7768,N_7577,N_7526);
nand U7769 (N_7769,N_7511,N_7603);
xnor U7770 (N_7770,N_7589,N_7527);
or U7771 (N_7771,N_7506,N_7647);
nand U7772 (N_7772,N_7509,N_7592);
and U7773 (N_7773,N_7648,N_7607);
or U7774 (N_7774,N_7586,N_7649);
nor U7775 (N_7775,N_7528,N_7553);
xnor U7776 (N_7776,N_7503,N_7536);
and U7777 (N_7777,N_7590,N_7618);
and U7778 (N_7778,N_7545,N_7520);
xor U7779 (N_7779,N_7604,N_7530);
and U7780 (N_7780,N_7503,N_7584);
nand U7781 (N_7781,N_7559,N_7602);
nand U7782 (N_7782,N_7528,N_7527);
or U7783 (N_7783,N_7538,N_7627);
and U7784 (N_7784,N_7557,N_7521);
or U7785 (N_7785,N_7550,N_7522);
xor U7786 (N_7786,N_7545,N_7586);
xor U7787 (N_7787,N_7615,N_7633);
or U7788 (N_7788,N_7554,N_7614);
and U7789 (N_7789,N_7510,N_7522);
nor U7790 (N_7790,N_7648,N_7605);
nand U7791 (N_7791,N_7633,N_7553);
nand U7792 (N_7792,N_7505,N_7541);
nor U7793 (N_7793,N_7531,N_7522);
nor U7794 (N_7794,N_7580,N_7624);
nand U7795 (N_7795,N_7640,N_7567);
xnor U7796 (N_7796,N_7596,N_7564);
and U7797 (N_7797,N_7557,N_7562);
or U7798 (N_7798,N_7516,N_7624);
xor U7799 (N_7799,N_7647,N_7599);
nand U7800 (N_7800,N_7667,N_7665);
nand U7801 (N_7801,N_7657,N_7677);
nand U7802 (N_7802,N_7662,N_7688);
nand U7803 (N_7803,N_7723,N_7798);
nand U7804 (N_7804,N_7782,N_7661);
nor U7805 (N_7805,N_7757,N_7715);
and U7806 (N_7806,N_7651,N_7762);
nand U7807 (N_7807,N_7748,N_7672);
and U7808 (N_7808,N_7676,N_7689);
and U7809 (N_7809,N_7743,N_7731);
xnor U7810 (N_7810,N_7658,N_7738);
or U7811 (N_7811,N_7663,N_7705);
xnor U7812 (N_7812,N_7684,N_7732);
nand U7813 (N_7813,N_7788,N_7787);
xor U7814 (N_7814,N_7668,N_7783);
nand U7815 (N_7815,N_7746,N_7784);
xor U7816 (N_7816,N_7721,N_7682);
xor U7817 (N_7817,N_7742,N_7741);
or U7818 (N_7818,N_7653,N_7704);
nor U7819 (N_7819,N_7713,N_7719);
nor U7820 (N_7820,N_7708,N_7764);
or U7821 (N_7821,N_7726,N_7656);
and U7822 (N_7822,N_7786,N_7673);
or U7823 (N_7823,N_7794,N_7680);
nand U7824 (N_7824,N_7768,N_7754);
nor U7825 (N_7825,N_7650,N_7694);
or U7826 (N_7826,N_7711,N_7777);
nand U7827 (N_7827,N_7749,N_7717);
nor U7828 (N_7828,N_7730,N_7654);
nand U7829 (N_7829,N_7752,N_7693);
and U7830 (N_7830,N_7755,N_7686);
xor U7831 (N_7831,N_7799,N_7702);
xnor U7832 (N_7832,N_7776,N_7670);
xor U7833 (N_7833,N_7770,N_7735);
and U7834 (N_7834,N_7745,N_7760);
nand U7835 (N_7835,N_7766,N_7712);
nand U7836 (N_7836,N_7685,N_7736);
and U7837 (N_7837,N_7698,N_7771);
nor U7838 (N_7838,N_7758,N_7792);
or U7839 (N_7839,N_7692,N_7791);
nand U7840 (N_7840,N_7793,N_7683);
nand U7841 (N_7841,N_7795,N_7737);
nand U7842 (N_7842,N_7671,N_7778);
nor U7843 (N_7843,N_7718,N_7659);
nor U7844 (N_7844,N_7775,N_7706);
or U7845 (N_7845,N_7709,N_7722);
and U7846 (N_7846,N_7769,N_7780);
nor U7847 (N_7847,N_7740,N_7687);
and U7848 (N_7848,N_7720,N_7725);
and U7849 (N_7849,N_7714,N_7700);
nand U7850 (N_7850,N_7669,N_7747);
or U7851 (N_7851,N_7697,N_7664);
nor U7852 (N_7852,N_7727,N_7790);
nand U7853 (N_7853,N_7674,N_7707);
nor U7854 (N_7854,N_7734,N_7724);
nand U7855 (N_7855,N_7710,N_7681);
nand U7856 (N_7856,N_7774,N_7767);
and U7857 (N_7857,N_7696,N_7675);
and U7858 (N_7858,N_7703,N_7744);
and U7859 (N_7859,N_7701,N_7751);
and U7860 (N_7860,N_7773,N_7765);
and U7861 (N_7861,N_7699,N_7739);
xor U7862 (N_7862,N_7750,N_7781);
and U7863 (N_7863,N_7761,N_7797);
nor U7864 (N_7864,N_7728,N_7678);
nand U7865 (N_7865,N_7716,N_7666);
nor U7866 (N_7866,N_7695,N_7779);
or U7867 (N_7867,N_7660,N_7652);
nor U7868 (N_7868,N_7759,N_7733);
and U7869 (N_7869,N_7679,N_7753);
and U7870 (N_7870,N_7763,N_7691);
nand U7871 (N_7871,N_7729,N_7772);
xnor U7872 (N_7872,N_7756,N_7690);
nand U7873 (N_7873,N_7796,N_7785);
and U7874 (N_7874,N_7655,N_7789);
and U7875 (N_7875,N_7739,N_7692);
or U7876 (N_7876,N_7728,N_7743);
nand U7877 (N_7877,N_7694,N_7652);
xor U7878 (N_7878,N_7793,N_7785);
nor U7879 (N_7879,N_7688,N_7746);
xor U7880 (N_7880,N_7709,N_7797);
and U7881 (N_7881,N_7656,N_7750);
nand U7882 (N_7882,N_7674,N_7752);
nand U7883 (N_7883,N_7688,N_7769);
or U7884 (N_7884,N_7689,N_7702);
nand U7885 (N_7885,N_7656,N_7688);
nor U7886 (N_7886,N_7656,N_7692);
nand U7887 (N_7887,N_7656,N_7681);
and U7888 (N_7888,N_7733,N_7796);
or U7889 (N_7889,N_7715,N_7727);
xnor U7890 (N_7890,N_7695,N_7704);
nand U7891 (N_7891,N_7652,N_7767);
and U7892 (N_7892,N_7669,N_7740);
and U7893 (N_7893,N_7742,N_7690);
nor U7894 (N_7894,N_7673,N_7651);
nand U7895 (N_7895,N_7784,N_7760);
and U7896 (N_7896,N_7770,N_7665);
and U7897 (N_7897,N_7768,N_7782);
nand U7898 (N_7898,N_7777,N_7721);
and U7899 (N_7899,N_7658,N_7668);
nor U7900 (N_7900,N_7729,N_7755);
xor U7901 (N_7901,N_7673,N_7676);
and U7902 (N_7902,N_7658,N_7768);
or U7903 (N_7903,N_7693,N_7695);
or U7904 (N_7904,N_7791,N_7798);
or U7905 (N_7905,N_7750,N_7739);
or U7906 (N_7906,N_7791,N_7661);
and U7907 (N_7907,N_7717,N_7785);
or U7908 (N_7908,N_7742,N_7777);
nor U7909 (N_7909,N_7656,N_7714);
or U7910 (N_7910,N_7731,N_7752);
nand U7911 (N_7911,N_7689,N_7650);
nor U7912 (N_7912,N_7749,N_7703);
or U7913 (N_7913,N_7733,N_7671);
and U7914 (N_7914,N_7689,N_7760);
or U7915 (N_7915,N_7758,N_7749);
or U7916 (N_7916,N_7699,N_7663);
xor U7917 (N_7917,N_7699,N_7697);
nor U7918 (N_7918,N_7673,N_7678);
nand U7919 (N_7919,N_7711,N_7650);
nand U7920 (N_7920,N_7733,N_7725);
nand U7921 (N_7921,N_7727,N_7743);
or U7922 (N_7922,N_7785,N_7764);
nor U7923 (N_7923,N_7765,N_7732);
xnor U7924 (N_7924,N_7776,N_7770);
nor U7925 (N_7925,N_7732,N_7734);
or U7926 (N_7926,N_7745,N_7694);
nand U7927 (N_7927,N_7658,N_7716);
xnor U7928 (N_7928,N_7691,N_7767);
or U7929 (N_7929,N_7759,N_7732);
nor U7930 (N_7930,N_7787,N_7696);
xnor U7931 (N_7931,N_7750,N_7699);
or U7932 (N_7932,N_7715,N_7714);
nand U7933 (N_7933,N_7781,N_7787);
xor U7934 (N_7934,N_7660,N_7771);
xnor U7935 (N_7935,N_7758,N_7701);
or U7936 (N_7936,N_7721,N_7792);
and U7937 (N_7937,N_7781,N_7672);
and U7938 (N_7938,N_7772,N_7756);
xnor U7939 (N_7939,N_7689,N_7723);
and U7940 (N_7940,N_7757,N_7760);
nor U7941 (N_7941,N_7672,N_7738);
nand U7942 (N_7942,N_7668,N_7670);
or U7943 (N_7943,N_7744,N_7720);
nor U7944 (N_7944,N_7734,N_7727);
nand U7945 (N_7945,N_7777,N_7791);
nand U7946 (N_7946,N_7688,N_7654);
xnor U7947 (N_7947,N_7709,N_7680);
or U7948 (N_7948,N_7769,N_7733);
nor U7949 (N_7949,N_7693,N_7749);
or U7950 (N_7950,N_7800,N_7936);
xnor U7951 (N_7951,N_7835,N_7888);
and U7952 (N_7952,N_7899,N_7842);
nand U7953 (N_7953,N_7821,N_7940);
xnor U7954 (N_7954,N_7844,N_7810);
xor U7955 (N_7955,N_7874,N_7884);
xor U7956 (N_7956,N_7906,N_7944);
xor U7957 (N_7957,N_7934,N_7945);
and U7958 (N_7958,N_7860,N_7917);
or U7959 (N_7959,N_7859,N_7925);
xnor U7960 (N_7960,N_7938,N_7869);
nor U7961 (N_7961,N_7892,N_7921);
nand U7962 (N_7962,N_7894,N_7834);
xnor U7963 (N_7963,N_7886,N_7832);
xor U7964 (N_7964,N_7912,N_7863);
or U7965 (N_7965,N_7935,N_7898);
nand U7966 (N_7966,N_7919,N_7825);
nor U7967 (N_7967,N_7871,N_7848);
nor U7968 (N_7968,N_7904,N_7937);
nor U7969 (N_7969,N_7932,N_7883);
nand U7970 (N_7970,N_7850,N_7846);
xnor U7971 (N_7971,N_7916,N_7939);
and U7972 (N_7972,N_7882,N_7830);
nand U7973 (N_7973,N_7890,N_7914);
and U7974 (N_7974,N_7818,N_7897);
or U7975 (N_7975,N_7909,N_7828);
nor U7976 (N_7976,N_7929,N_7852);
nand U7977 (N_7977,N_7827,N_7851);
and U7978 (N_7978,N_7901,N_7891);
nand U7979 (N_7979,N_7805,N_7803);
nand U7980 (N_7980,N_7878,N_7942);
xor U7981 (N_7981,N_7920,N_7812);
or U7982 (N_7982,N_7811,N_7826);
or U7983 (N_7983,N_7872,N_7840);
nand U7984 (N_7984,N_7895,N_7902);
nand U7985 (N_7985,N_7815,N_7866);
and U7986 (N_7986,N_7864,N_7949);
nand U7987 (N_7987,N_7856,N_7802);
or U7988 (N_7988,N_7873,N_7907);
and U7989 (N_7989,N_7865,N_7927);
xnor U7990 (N_7990,N_7928,N_7833);
xnor U7991 (N_7991,N_7903,N_7824);
nand U7992 (N_7992,N_7879,N_7876);
nand U7993 (N_7993,N_7931,N_7819);
and U7994 (N_7994,N_7808,N_7820);
nand U7995 (N_7995,N_7941,N_7806);
nand U7996 (N_7996,N_7923,N_7838);
xnor U7997 (N_7997,N_7926,N_7836);
or U7998 (N_7998,N_7837,N_7885);
nand U7999 (N_7999,N_7809,N_7918);
nor U8000 (N_8000,N_7922,N_7807);
xor U8001 (N_8001,N_7862,N_7847);
nand U8002 (N_8002,N_7858,N_7801);
xor U8003 (N_8003,N_7910,N_7947);
or U8004 (N_8004,N_7853,N_7905);
nand U8005 (N_8005,N_7875,N_7814);
or U8006 (N_8006,N_7889,N_7839);
or U8007 (N_8007,N_7870,N_7816);
nor U8008 (N_8008,N_7893,N_7900);
or U8009 (N_8009,N_7829,N_7887);
or U8010 (N_8010,N_7857,N_7861);
xor U8011 (N_8011,N_7804,N_7867);
nor U8012 (N_8012,N_7855,N_7896);
and U8013 (N_8013,N_7831,N_7911);
nand U8014 (N_8014,N_7880,N_7849);
xnor U8015 (N_8015,N_7930,N_7841);
nand U8016 (N_8016,N_7915,N_7813);
xnor U8017 (N_8017,N_7877,N_7913);
xnor U8018 (N_8018,N_7924,N_7948);
or U8019 (N_8019,N_7908,N_7881);
xnor U8020 (N_8020,N_7845,N_7823);
nor U8021 (N_8021,N_7817,N_7868);
or U8022 (N_8022,N_7822,N_7946);
xnor U8023 (N_8023,N_7854,N_7933);
and U8024 (N_8024,N_7943,N_7843);
xor U8025 (N_8025,N_7810,N_7876);
and U8026 (N_8026,N_7839,N_7836);
nand U8027 (N_8027,N_7918,N_7835);
or U8028 (N_8028,N_7817,N_7911);
nand U8029 (N_8029,N_7806,N_7943);
xor U8030 (N_8030,N_7813,N_7900);
xnor U8031 (N_8031,N_7882,N_7821);
or U8032 (N_8032,N_7865,N_7822);
xnor U8033 (N_8033,N_7847,N_7939);
nand U8034 (N_8034,N_7836,N_7879);
and U8035 (N_8035,N_7851,N_7915);
xor U8036 (N_8036,N_7827,N_7874);
or U8037 (N_8037,N_7934,N_7938);
nand U8038 (N_8038,N_7843,N_7933);
nand U8039 (N_8039,N_7864,N_7906);
xor U8040 (N_8040,N_7945,N_7885);
and U8041 (N_8041,N_7864,N_7885);
nand U8042 (N_8042,N_7846,N_7921);
xnor U8043 (N_8043,N_7896,N_7866);
xnor U8044 (N_8044,N_7814,N_7918);
and U8045 (N_8045,N_7909,N_7944);
nand U8046 (N_8046,N_7907,N_7924);
nor U8047 (N_8047,N_7883,N_7933);
nand U8048 (N_8048,N_7943,N_7909);
xor U8049 (N_8049,N_7823,N_7932);
nand U8050 (N_8050,N_7835,N_7849);
nor U8051 (N_8051,N_7848,N_7918);
and U8052 (N_8052,N_7866,N_7918);
xnor U8053 (N_8053,N_7879,N_7802);
and U8054 (N_8054,N_7943,N_7946);
xnor U8055 (N_8055,N_7915,N_7918);
nand U8056 (N_8056,N_7943,N_7870);
xor U8057 (N_8057,N_7867,N_7924);
xor U8058 (N_8058,N_7915,N_7942);
nand U8059 (N_8059,N_7849,N_7856);
or U8060 (N_8060,N_7904,N_7849);
or U8061 (N_8061,N_7803,N_7896);
xor U8062 (N_8062,N_7817,N_7875);
nand U8063 (N_8063,N_7863,N_7836);
xnor U8064 (N_8064,N_7801,N_7881);
nor U8065 (N_8065,N_7884,N_7860);
xnor U8066 (N_8066,N_7928,N_7859);
nor U8067 (N_8067,N_7810,N_7808);
or U8068 (N_8068,N_7816,N_7927);
or U8069 (N_8069,N_7845,N_7858);
xnor U8070 (N_8070,N_7923,N_7842);
and U8071 (N_8071,N_7859,N_7823);
nand U8072 (N_8072,N_7905,N_7838);
or U8073 (N_8073,N_7876,N_7907);
xor U8074 (N_8074,N_7827,N_7903);
nand U8075 (N_8075,N_7857,N_7881);
xor U8076 (N_8076,N_7905,N_7842);
or U8077 (N_8077,N_7852,N_7849);
xor U8078 (N_8078,N_7936,N_7802);
and U8079 (N_8079,N_7887,N_7923);
nor U8080 (N_8080,N_7854,N_7855);
or U8081 (N_8081,N_7848,N_7894);
nand U8082 (N_8082,N_7885,N_7934);
or U8083 (N_8083,N_7861,N_7930);
xnor U8084 (N_8084,N_7906,N_7867);
nor U8085 (N_8085,N_7823,N_7868);
or U8086 (N_8086,N_7883,N_7800);
nor U8087 (N_8087,N_7803,N_7929);
and U8088 (N_8088,N_7916,N_7808);
or U8089 (N_8089,N_7920,N_7917);
nand U8090 (N_8090,N_7825,N_7945);
nor U8091 (N_8091,N_7832,N_7808);
or U8092 (N_8092,N_7830,N_7941);
nand U8093 (N_8093,N_7893,N_7838);
xor U8094 (N_8094,N_7815,N_7927);
or U8095 (N_8095,N_7917,N_7931);
or U8096 (N_8096,N_7861,N_7910);
and U8097 (N_8097,N_7901,N_7915);
or U8098 (N_8098,N_7817,N_7943);
and U8099 (N_8099,N_7920,N_7824);
or U8100 (N_8100,N_8082,N_8076);
and U8101 (N_8101,N_7987,N_7993);
xor U8102 (N_8102,N_7996,N_8042);
and U8103 (N_8103,N_8047,N_8000);
nand U8104 (N_8104,N_7981,N_7970);
nand U8105 (N_8105,N_8007,N_8087);
nand U8106 (N_8106,N_8041,N_8023);
or U8107 (N_8107,N_8039,N_8090);
or U8108 (N_8108,N_8020,N_8033);
nand U8109 (N_8109,N_8061,N_8073);
and U8110 (N_8110,N_8032,N_7972);
nor U8111 (N_8111,N_7978,N_7951);
nand U8112 (N_8112,N_8084,N_8010);
nor U8113 (N_8113,N_8066,N_8014);
or U8114 (N_8114,N_8045,N_8003);
xor U8115 (N_8115,N_8009,N_7965);
or U8116 (N_8116,N_7984,N_7963);
nand U8117 (N_8117,N_8024,N_8037);
xnor U8118 (N_8118,N_8071,N_8028);
and U8119 (N_8119,N_8006,N_8025);
or U8120 (N_8120,N_8004,N_8067);
xor U8121 (N_8121,N_8064,N_8093);
or U8122 (N_8122,N_8005,N_7953);
and U8123 (N_8123,N_8058,N_8013);
and U8124 (N_8124,N_7994,N_7975);
xnor U8125 (N_8125,N_8051,N_8048);
xor U8126 (N_8126,N_8083,N_7974);
xor U8127 (N_8127,N_7961,N_8079);
nand U8128 (N_8128,N_8026,N_7966);
xnor U8129 (N_8129,N_8008,N_8043);
nand U8130 (N_8130,N_8022,N_8088);
or U8131 (N_8131,N_8085,N_7964);
xnor U8132 (N_8132,N_8056,N_7988);
xnor U8133 (N_8133,N_8086,N_8072);
xor U8134 (N_8134,N_8011,N_8002);
xor U8135 (N_8135,N_8057,N_8049);
nand U8136 (N_8136,N_8052,N_8096);
xor U8137 (N_8137,N_8038,N_7979);
nand U8138 (N_8138,N_8017,N_7985);
nor U8139 (N_8139,N_8089,N_7983);
xor U8140 (N_8140,N_8098,N_7958);
or U8141 (N_8141,N_8044,N_7980);
nor U8142 (N_8142,N_8091,N_8034);
nand U8143 (N_8143,N_8035,N_8075);
or U8144 (N_8144,N_8081,N_8054);
or U8145 (N_8145,N_8092,N_8055);
xnor U8146 (N_8146,N_8036,N_7967);
xnor U8147 (N_8147,N_7956,N_7997);
nand U8148 (N_8148,N_8027,N_8019);
and U8149 (N_8149,N_8040,N_7968);
xor U8150 (N_8150,N_8070,N_7991);
or U8151 (N_8151,N_7986,N_8060);
or U8152 (N_8152,N_7973,N_8050);
nor U8153 (N_8153,N_8031,N_7955);
xor U8154 (N_8154,N_8021,N_7995);
and U8155 (N_8155,N_8097,N_7960);
nor U8156 (N_8156,N_8063,N_8068);
nor U8157 (N_8157,N_8069,N_7954);
nor U8158 (N_8158,N_8012,N_7959);
and U8159 (N_8159,N_8029,N_8062);
or U8160 (N_8160,N_7998,N_8078);
nand U8161 (N_8161,N_7976,N_8080);
nor U8162 (N_8162,N_7989,N_7952);
and U8163 (N_8163,N_8001,N_8015);
or U8164 (N_8164,N_7969,N_8018);
and U8165 (N_8165,N_8065,N_7950);
or U8166 (N_8166,N_7977,N_8053);
and U8167 (N_8167,N_8030,N_7971);
and U8168 (N_8168,N_8094,N_7957);
and U8169 (N_8169,N_7982,N_8074);
and U8170 (N_8170,N_8077,N_7990);
nor U8171 (N_8171,N_8046,N_8095);
xor U8172 (N_8172,N_7962,N_8016);
nor U8173 (N_8173,N_8059,N_7992);
xnor U8174 (N_8174,N_8099,N_7999);
nand U8175 (N_8175,N_8063,N_8044);
or U8176 (N_8176,N_8009,N_8023);
nand U8177 (N_8177,N_8044,N_8027);
and U8178 (N_8178,N_8037,N_7980);
or U8179 (N_8179,N_7987,N_8009);
or U8180 (N_8180,N_7970,N_8049);
nand U8181 (N_8181,N_7955,N_8035);
and U8182 (N_8182,N_8038,N_7963);
nor U8183 (N_8183,N_8067,N_8047);
xnor U8184 (N_8184,N_8071,N_7958);
and U8185 (N_8185,N_8062,N_7973);
xor U8186 (N_8186,N_8039,N_8078);
xor U8187 (N_8187,N_7962,N_7980);
xnor U8188 (N_8188,N_7975,N_7986);
xor U8189 (N_8189,N_8041,N_8097);
and U8190 (N_8190,N_8023,N_8074);
nand U8191 (N_8191,N_8059,N_8074);
and U8192 (N_8192,N_8064,N_7997);
xnor U8193 (N_8193,N_8078,N_7999);
and U8194 (N_8194,N_7987,N_8015);
or U8195 (N_8195,N_7972,N_7958);
or U8196 (N_8196,N_7954,N_7959);
and U8197 (N_8197,N_7988,N_7995);
xnor U8198 (N_8198,N_8086,N_7994);
and U8199 (N_8199,N_8091,N_7996);
xnor U8200 (N_8200,N_8099,N_8008);
nor U8201 (N_8201,N_7962,N_7965);
nand U8202 (N_8202,N_8088,N_8071);
nand U8203 (N_8203,N_7979,N_8001);
and U8204 (N_8204,N_7976,N_7987);
nor U8205 (N_8205,N_8004,N_8089);
or U8206 (N_8206,N_8061,N_8018);
nand U8207 (N_8207,N_8058,N_8076);
and U8208 (N_8208,N_8035,N_7984);
or U8209 (N_8209,N_8053,N_8051);
or U8210 (N_8210,N_7975,N_8079);
xor U8211 (N_8211,N_8035,N_7957);
or U8212 (N_8212,N_8086,N_8068);
or U8213 (N_8213,N_7979,N_8098);
and U8214 (N_8214,N_8090,N_8058);
or U8215 (N_8215,N_8084,N_8058);
nor U8216 (N_8216,N_7954,N_8045);
xor U8217 (N_8217,N_7974,N_8070);
or U8218 (N_8218,N_8064,N_8031);
xnor U8219 (N_8219,N_8012,N_8032);
nand U8220 (N_8220,N_7951,N_8092);
nor U8221 (N_8221,N_7951,N_8039);
or U8222 (N_8222,N_8075,N_8074);
nor U8223 (N_8223,N_8038,N_8008);
nor U8224 (N_8224,N_8046,N_7951);
and U8225 (N_8225,N_8015,N_8082);
xnor U8226 (N_8226,N_8078,N_7955);
nor U8227 (N_8227,N_7960,N_8036);
or U8228 (N_8228,N_8007,N_8001);
xor U8229 (N_8229,N_8083,N_8027);
nor U8230 (N_8230,N_8065,N_8035);
nand U8231 (N_8231,N_8095,N_7979);
or U8232 (N_8232,N_8001,N_7975);
nand U8233 (N_8233,N_7991,N_7992);
or U8234 (N_8234,N_8027,N_8018);
xor U8235 (N_8235,N_8025,N_7955);
xnor U8236 (N_8236,N_7960,N_8022);
xor U8237 (N_8237,N_7961,N_8052);
nand U8238 (N_8238,N_8019,N_8086);
nor U8239 (N_8239,N_8042,N_8032);
or U8240 (N_8240,N_8071,N_8089);
and U8241 (N_8241,N_8049,N_8011);
nand U8242 (N_8242,N_8065,N_8071);
and U8243 (N_8243,N_8077,N_8074);
and U8244 (N_8244,N_8059,N_8021);
xnor U8245 (N_8245,N_7991,N_8003);
or U8246 (N_8246,N_8037,N_7991);
nand U8247 (N_8247,N_7951,N_8093);
and U8248 (N_8248,N_8053,N_8084);
and U8249 (N_8249,N_8048,N_8061);
or U8250 (N_8250,N_8218,N_8105);
or U8251 (N_8251,N_8223,N_8197);
nor U8252 (N_8252,N_8195,N_8226);
or U8253 (N_8253,N_8122,N_8244);
nor U8254 (N_8254,N_8162,N_8170);
nand U8255 (N_8255,N_8235,N_8154);
xor U8256 (N_8256,N_8231,N_8128);
nor U8257 (N_8257,N_8148,N_8115);
nor U8258 (N_8258,N_8176,N_8234);
or U8259 (N_8259,N_8144,N_8224);
nor U8260 (N_8260,N_8174,N_8156);
xnor U8261 (N_8261,N_8168,N_8230);
or U8262 (N_8262,N_8183,N_8125);
xnor U8263 (N_8263,N_8107,N_8113);
xor U8264 (N_8264,N_8219,N_8116);
or U8265 (N_8265,N_8126,N_8221);
xor U8266 (N_8266,N_8157,N_8199);
nor U8267 (N_8267,N_8249,N_8160);
and U8268 (N_8268,N_8150,N_8117);
and U8269 (N_8269,N_8139,N_8134);
nor U8270 (N_8270,N_8102,N_8152);
nor U8271 (N_8271,N_8146,N_8100);
and U8272 (N_8272,N_8165,N_8225);
nor U8273 (N_8273,N_8121,N_8149);
nor U8274 (N_8274,N_8111,N_8194);
xnor U8275 (N_8275,N_8210,N_8246);
or U8276 (N_8276,N_8142,N_8184);
or U8277 (N_8277,N_8215,N_8202);
or U8278 (N_8278,N_8151,N_8187);
xor U8279 (N_8279,N_8217,N_8119);
nor U8280 (N_8280,N_8228,N_8123);
or U8281 (N_8281,N_8133,N_8166);
and U8282 (N_8282,N_8220,N_8233);
or U8283 (N_8283,N_8110,N_8137);
and U8284 (N_8284,N_8211,N_8186);
nor U8285 (N_8285,N_8177,N_8138);
nor U8286 (N_8286,N_8169,N_8193);
nor U8287 (N_8287,N_8114,N_8208);
and U8288 (N_8288,N_8209,N_8131);
or U8289 (N_8289,N_8243,N_8214);
and U8290 (N_8290,N_8229,N_8112);
nand U8291 (N_8291,N_8213,N_8188);
nor U8292 (N_8292,N_8158,N_8207);
and U8293 (N_8293,N_8216,N_8127);
or U8294 (N_8294,N_8201,N_8239);
nand U8295 (N_8295,N_8205,N_8141);
or U8296 (N_8296,N_8104,N_8124);
or U8297 (N_8297,N_8159,N_8140);
xor U8298 (N_8298,N_8192,N_8164);
nand U8299 (N_8299,N_8237,N_8120);
xor U8300 (N_8300,N_8241,N_8108);
and U8301 (N_8301,N_8181,N_8167);
nor U8302 (N_8302,N_8204,N_8143);
nand U8303 (N_8303,N_8175,N_8196);
or U8304 (N_8304,N_8145,N_8171);
and U8305 (N_8305,N_8242,N_8147);
nor U8306 (N_8306,N_8238,N_8222);
or U8307 (N_8307,N_8129,N_8136);
or U8308 (N_8308,N_8198,N_8191);
xnor U8309 (N_8309,N_8173,N_8118);
nor U8310 (N_8310,N_8155,N_8240);
nor U8311 (N_8311,N_8179,N_8203);
xnor U8312 (N_8312,N_8182,N_8206);
nand U8313 (N_8313,N_8190,N_8132);
and U8314 (N_8314,N_8227,N_8106);
or U8315 (N_8315,N_8135,N_8101);
and U8316 (N_8316,N_8180,N_8161);
xnor U8317 (N_8317,N_8247,N_8245);
nor U8318 (N_8318,N_8189,N_8185);
xnor U8319 (N_8319,N_8163,N_8130);
or U8320 (N_8320,N_8200,N_8236);
or U8321 (N_8321,N_8153,N_8178);
and U8322 (N_8322,N_8248,N_8212);
xnor U8323 (N_8323,N_8109,N_8232);
nor U8324 (N_8324,N_8172,N_8103);
or U8325 (N_8325,N_8157,N_8220);
nor U8326 (N_8326,N_8218,N_8109);
xnor U8327 (N_8327,N_8123,N_8151);
nand U8328 (N_8328,N_8136,N_8199);
nor U8329 (N_8329,N_8158,N_8165);
nand U8330 (N_8330,N_8175,N_8188);
xor U8331 (N_8331,N_8103,N_8193);
and U8332 (N_8332,N_8112,N_8185);
nor U8333 (N_8333,N_8120,N_8241);
or U8334 (N_8334,N_8108,N_8159);
nand U8335 (N_8335,N_8192,N_8127);
and U8336 (N_8336,N_8156,N_8175);
and U8337 (N_8337,N_8147,N_8232);
or U8338 (N_8338,N_8140,N_8206);
nor U8339 (N_8339,N_8240,N_8161);
or U8340 (N_8340,N_8176,N_8157);
and U8341 (N_8341,N_8121,N_8215);
and U8342 (N_8342,N_8139,N_8118);
xor U8343 (N_8343,N_8216,N_8192);
and U8344 (N_8344,N_8173,N_8239);
xnor U8345 (N_8345,N_8117,N_8127);
xnor U8346 (N_8346,N_8157,N_8104);
or U8347 (N_8347,N_8151,N_8137);
nand U8348 (N_8348,N_8189,N_8163);
and U8349 (N_8349,N_8239,N_8160);
and U8350 (N_8350,N_8130,N_8182);
or U8351 (N_8351,N_8158,N_8193);
or U8352 (N_8352,N_8193,N_8117);
nand U8353 (N_8353,N_8225,N_8246);
nand U8354 (N_8354,N_8101,N_8208);
or U8355 (N_8355,N_8142,N_8100);
or U8356 (N_8356,N_8206,N_8186);
nand U8357 (N_8357,N_8197,N_8202);
or U8358 (N_8358,N_8157,N_8210);
nand U8359 (N_8359,N_8201,N_8192);
nand U8360 (N_8360,N_8142,N_8103);
or U8361 (N_8361,N_8145,N_8108);
nand U8362 (N_8362,N_8146,N_8195);
nor U8363 (N_8363,N_8228,N_8240);
or U8364 (N_8364,N_8177,N_8222);
nand U8365 (N_8365,N_8111,N_8244);
nand U8366 (N_8366,N_8148,N_8130);
and U8367 (N_8367,N_8195,N_8139);
or U8368 (N_8368,N_8176,N_8105);
or U8369 (N_8369,N_8170,N_8243);
or U8370 (N_8370,N_8194,N_8138);
nand U8371 (N_8371,N_8180,N_8194);
nand U8372 (N_8372,N_8104,N_8211);
nand U8373 (N_8373,N_8219,N_8122);
and U8374 (N_8374,N_8249,N_8163);
nor U8375 (N_8375,N_8108,N_8178);
or U8376 (N_8376,N_8181,N_8186);
and U8377 (N_8377,N_8129,N_8158);
nand U8378 (N_8378,N_8160,N_8181);
nand U8379 (N_8379,N_8183,N_8116);
and U8380 (N_8380,N_8100,N_8138);
xnor U8381 (N_8381,N_8173,N_8174);
nor U8382 (N_8382,N_8207,N_8182);
nor U8383 (N_8383,N_8248,N_8195);
nor U8384 (N_8384,N_8187,N_8232);
xnor U8385 (N_8385,N_8236,N_8230);
xnor U8386 (N_8386,N_8189,N_8161);
nand U8387 (N_8387,N_8130,N_8186);
nand U8388 (N_8388,N_8167,N_8192);
nand U8389 (N_8389,N_8147,N_8231);
nor U8390 (N_8390,N_8182,N_8218);
and U8391 (N_8391,N_8244,N_8245);
xnor U8392 (N_8392,N_8151,N_8240);
xor U8393 (N_8393,N_8195,N_8166);
nor U8394 (N_8394,N_8192,N_8221);
or U8395 (N_8395,N_8106,N_8134);
nand U8396 (N_8396,N_8245,N_8156);
xor U8397 (N_8397,N_8182,N_8149);
xor U8398 (N_8398,N_8201,N_8102);
nor U8399 (N_8399,N_8184,N_8226);
nand U8400 (N_8400,N_8265,N_8329);
nor U8401 (N_8401,N_8309,N_8314);
or U8402 (N_8402,N_8337,N_8272);
nor U8403 (N_8403,N_8321,N_8334);
nand U8404 (N_8404,N_8380,N_8282);
nor U8405 (N_8405,N_8353,N_8378);
nand U8406 (N_8406,N_8311,N_8336);
or U8407 (N_8407,N_8346,N_8290);
nor U8408 (N_8408,N_8362,N_8264);
xor U8409 (N_8409,N_8322,N_8278);
nor U8410 (N_8410,N_8304,N_8384);
or U8411 (N_8411,N_8287,N_8361);
nand U8412 (N_8412,N_8285,N_8303);
or U8413 (N_8413,N_8251,N_8333);
or U8414 (N_8414,N_8307,N_8359);
xor U8415 (N_8415,N_8385,N_8393);
and U8416 (N_8416,N_8369,N_8328);
nor U8417 (N_8417,N_8364,N_8350);
or U8418 (N_8418,N_8312,N_8373);
and U8419 (N_8419,N_8399,N_8374);
and U8420 (N_8420,N_8270,N_8302);
xnor U8421 (N_8421,N_8388,N_8269);
nand U8422 (N_8422,N_8300,N_8366);
nand U8423 (N_8423,N_8263,N_8383);
xor U8424 (N_8424,N_8292,N_8254);
and U8425 (N_8425,N_8339,N_8349);
or U8426 (N_8426,N_8275,N_8252);
and U8427 (N_8427,N_8274,N_8368);
or U8428 (N_8428,N_8267,N_8375);
nand U8429 (N_8429,N_8310,N_8352);
or U8430 (N_8430,N_8331,N_8332);
nor U8431 (N_8431,N_8396,N_8294);
and U8432 (N_8432,N_8382,N_8367);
xor U8433 (N_8433,N_8316,N_8360);
and U8434 (N_8434,N_8296,N_8268);
and U8435 (N_8435,N_8255,N_8342);
xor U8436 (N_8436,N_8376,N_8351);
and U8437 (N_8437,N_8319,N_8327);
xor U8438 (N_8438,N_8293,N_8324);
nand U8439 (N_8439,N_8279,N_8390);
nor U8440 (N_8440,N_8397,N_8276);
nand U8441 (N_8441,N_8363,N_8356);
nor U8442 (N_8442,N_8394,N_8392);
nor U8443 (N_8443,N_8357,N_8259);
nor U8444 (N_8444,N_8283,N_8370);
xor U8445 (N_8445,N_8395,N_8391);
nor U8446 (N_8446,N_8354,N_8387);
and U8447 (N_8447,N_8358,N_8297);
xor U8448 (N_8448,N_8250,N_8260);
or U8449 (N_8449,N_8379,N_8338);
and U8450 (N_8450,N_8389,N_8273);
and U8451 (N_8451,N_8365,N_8281);
xnor U8452 (N_8452,N_8280,N_8271);
xnor U8453 (N_8453,N_8295,N_8348);
or U8454 (N_8454,N_8335,N_8266);
and U8455 (N_8455,N_8257,N_8381);
or U8456 (N_8456,N_8289,N_8330);
nor U8457 (N_8457,N_8261,N_8341);
or U8458 (N_8458,N_8256,N_8325);
or U8459 (N_8459,N_8371,N_8386);
or U8460 (N_8460,N_8323,N_8377);
and U8461 (N_8461,N_8372,N_8288);
xnor U8462 (N_8462,N_8317,N_8315);
and U8463 (N_8463,N_8318,N_8299);
or U8464 (N_8464,N_8301,N_8347);
and U8465 (N_8465,N_8308,N_8306);
or U8466 (N_8466,N_8398,N_8343);
or U8467 (N_8467,N_8344,N_8345);
xnor U8468 (N_8468,N_8320,N_8286);
nand U8469 (N_8469,N_8258,N_8326);
xor U8470 (N_8470,N_8313,N_8305);
xnor U8471 (N_8471,N_8277,N_8340);
xor U8472 (N_8472,N_8298,N_8262);
nand U8473 (N_8473,N_8355,N_8253);
nand U8474 (N_8474,N_8284,N_8291);
nand U8475 (N_8475,N_8280,N_8342);
nor U8476 (N_8476,N_8332,N_8399);
nor U8477 (N_8477,N_8252,N_8276);
nand U8478 (N_8478,N_8253,N_8385);
nor U8479 (N_8479,N_8364,N_8279);
xnor U8480 (N_8480,N_8384,N_8353);
and U8481 (N_8481,N_8277,N_8328);
nor U8482 (N_8482,N_8277,N_8396);
or U8483 (N_8483,N_8326,N_8364);
and U8484 (N_8484,N_8288,N_8362);
xor U8485 (N_8485,N_8307,N_8295);
or U8486 (N_8486,N_8354,N_8386);
or U8487 (N_8487,N_8277,N_8384);
nor U8488 (N_8488,N_8251,N_8399);
and U8489 (N_8489,N_8386,N_8339);
xor U8490 (N_8490,N_8398,N_8324);
nand U8491 (N_8491,N_8303,N_8283);
or U8492 (N_8492,N_8314,N_8336);
nor U8493 (N_8493,N_8253,N_8375);
and U8494 (N_8494,N_8363,N_8347);
nand U8495 (N_8495,N_8306,N_8309);
xnor U8496 (N_8496,N_8311,N_8394);
and U8497 (N_8497,N_8272,N_8315);
nand U8498 (N_8498,N_8339,N_8258);
xor U8499 (N_8499,N_8277,N_8278);
xor U8500 (N_8500,N_8386,N_8291);
nand U8501 (N_8501,N_8278,N_8377);
xnor U8502 (N_8502,N_8390,N_8336);
nor U8503 (N_8503,N_8305,N_8373);
xor U8504 (N_8504,N_8271,N_8389);
xnor U8505 (N_8505,N_8314,N_8399);
xor U8506 (N_8506,N_8347,N_8394);
xnor U8507 (N_8507,N_8273,N_8283);
nor U8508 (N_8508,N_8282,N_8342);
or U8509 (N_8509,N_8271,N_8253);
xnor U8510 (N_8510,N_8326,N_8306);
or U8511 (N_8511,N_8298,N_8278);
or U8512 (N_8512,N_8395,N_8311);
nor U8513 (N_8513,N_8387,N_8383);
nor U8514 (N_8514,N_8347,N_8352);
or U8515 (N_8515,N_8287,N_8346);
or U8516 (N_8516,N_8399,N_8360);
or U8517 (N_8517,N_8273,N_8274);
nor U8518 (N_8518,N_8358,N_8346);
nor U8519 (N_8519,N_8301,N_8395);
xnor U8520 (N_8520,N_8329,N_8356);
nor U8521 (N_8521,N_8250,N_8344);
and U8522 (N_8522,N_8394,N_8302);
nand U8523 (N_8523,N_8390,N_8344);
xor U8524 (N_8524,N_8364,N_8328);
or U8525 (N_8525,N_8367,N_8354);
and U8526 (N_8526,N_8305,N_8395);
nor U8527 (N_8527,N_8314,N_8356);
or U8528 (N_8528,N_8359,N_8308);
or U8529 (N_8529,N_8351,N_8326);
xnor U8530 (N_8530,N_8367,N_8296);
and U8531 (N_8531,N_8345,N_8271);
nor U8532 (N_8532,N_8318,N_8330);
and U8533 (N_8533,N_8301,N_8293);
nor U8534 (N_8534,N_8370,N_8250);
xnor U8535 (N_8535,N_8361,N_8300);
and U8536 (N_8536,N_8329,N_8262);
and U8537 (N_8537,N_8290,N_8298);
nand U8538 (N_8538,N_8259,N_8263);
nor U8539 (N_8539,N_8284,N_8383);
nor U8540 (N_8540,N_8257,N_8251);
and U8541 (N_8541,N_8344,N_8309);
xor U8542 (N_8542,N_8328,N_8291);
or U8543 (N_8543,N_8276,N_8283);
nor U8544 (N_8544,N_8390,N_8305);
and U8545 (N_8545,N_8321,N_8360);
xor U8546 (N_8546,N_8259,N_8273);
nand U8547 (N_8547,N_8255,N_8395);
and U8548 (N_8548,N_8254,N_8363);
xnor U8549 (N_8549,N_8326,N_8280);
and U8550 (N_8550,N_8424,N_8541);
or U8551 (N_8551,N_8509,N_8468);
or U8552 (N_8552,N_8437,N_8442);
or U8553 (N_8553,N_8535,N_8434);
nand U8554 (N_8554,N_8498,N_8533);
nand U8555 (N_8555,N_8433,N_8539);
and U8556 (N_8556,N_8531,N_8499);
nor U8557 (N_8557,N_8475,N_8438);
nand U8558 (N_8558,N_8482,N_8547);
nor U8559 (N_8559,N_8441,N_8430);
nor U8560 (N_8560,N_8529,N_8492);
xnor U8561 (N_8561,N_8478,N_8451);
xor U8562 (N_8562,N_8488,N_8505);
and U8563 (N_8563,N_8528,N_8490);
xnor U8564 (N_8564,N_8472,N_8519);
nor U8565 (N_8565,N_8443,N_8508);
and U8566 (N_8566,N_8516,N_8506);
and U8567 (N_8567,N_8402,N_8401);
xnor U8568 (N_8568,N_8517,N_8409);
nand U8569 (N_8569,N_8400,N_8500);
nor U8570 (N_8570,N_8484,N_8538);
or U8571 (N_8571,N_8406,N_8526);
xor U8572 (N_8572,N_8471,N_8456);
nand U8573 (N_8573,N_8515,N_8514);
nor U8574 (N_8574,N_8404,N_8425);
nor U8575 (N_8575,N_8428,N_8523);
nor U8576 (N_8576,N_8532,N_8534);
nand U8577 (N_8577,N_8522,N_8413);
xnor U8578 (N_8578,N_8540,N_8408);
and U8579 (N_8579,N_8491,N_8545);
nor U8580 (N_8580,N_8421,N_8494);
xnor U8581 (N_8581,N_8414,N_8449);
nor U8582 (N_8582,N_8521,N_8503);
nor U8583 (N_8583,N_8518,N_8524);
or U8584 (N_8584,N_8537,N_8549);
xor U8585 (N_8585,N_8445,N_8483);
nand U8586 (N_8586,N_8410,N_8546);
nand U8587 (N_8587,N_8493,N_8417);
nor U8588 (N_8588,N_8465,N_8467);
nand U8589 (N_8589,N_8530,N_8403);
nand U8590 (N_8590,N_8536,N_8415);
nor U8591 (N_8591,N_8520,N_8527);
and U8592 (N_8592,N_8458,N_8457);
and U8593 (N_8593,N_8446,N_8469);
or U8594 (N_8594,N_8416,N_8480);
nor U8595 (N_8595,N_8474,N_8486);
nand U8596 (N_8596,N_8431,N_8476);
and U8597 (N_8597,N_8423,N_8544);
nor U8598 (N_8598,N_8444,N_8489);
xor U8599 (N_8599,N_8497,N_8427);
or U8600 (N_8600,N_8479,N_8473);
nand U8601 (N_8601,N_8477,N_8429);
nand U8602 (N_8602,N_8510,N_8440);
nor U8603 (N_8603,N_8422,N_8511);
nand U8604 (N_8604,N_8412,N_8407);
and U8605 (N_8605,N_8542,N_8462);
nor U8606 (N_8606,N_8452,N_8466);
nand U8607 (N_8607,N_8455,N_8496);
or U8608 (N_8608,N_8459,N_8495);
xor U8609 (N_8609,N_8481,N_8454);
nand U8610 (N_8610,N_8543,N_8436);
and U8611 (N_8611,N_8435,N_8513);
nor U8612 (N_8612,N_8418,N_8420);
nand U8613 (N_8613,N_8432,N_8463);
and U8614 (N_8614,N_8448,N_8419);
or U8615 (N_8615,N_8450,N_8487);
or U8616 (N_8616,N_8502,N_8426);
and U8617 (N_8617,N_8447,N_8525);
nand U8618 (N_8618,N_8470,N_8460);
or U8619 (N_8619,N_8411,N_8507);
nor U8620 (N_8620,N_8485,N_8464);
or U8621 (N_8621,N_8548,N_8461);
xor U8622 (N_8622,N_8439,N_8405);
xnor U8623 (N_8623,N_8501,N_8512);
xor U8624 (N_8624,N_8453,N_8504);
and U8625 (N_8625,N_8425,N_8408);
and U8626 (N_8626,N_8523,N_8520);
or U8627 (N_8627,N_8478,N_8506);
nand U8628 (N_8628,N_8531,N_8498);
xor U8629 (N_8629,N_8528,N_8456);
and U8630 (N_8630,N_8527,N_8429);
xnor U8631 (N_8631,N_8426,N_8423);
xnor U8632 (N_8632,N_8443,N_8527);
and U8633 (N_8633,N_8402,N_8528);
or U8634 (N_8634,N_8528,N_8514);
nand U8635 (N_8635,N_8449,N_8540);
and U8636 (N_8636,N_8465,N_8478);
xnor U8637 (N_8637,N_8513,N_8527);
nor U8638 (N_8638,N_8462,N_8444);
or U8639 (N_8639,N_8540,N_8495);
xor U8640 (N_8640,N_8479,N_8490);
and U8641 (N_8641,N_8521,N_8416);
and U8642 (N_8642,N_8471,N_8499);
or U8643 (N_8643,N_8446,N_8520);
xor U8644 (N_8644,N_8491,N_8401);
and U8645 (N_8645,N_8546,N_8449);
xor U8646 (N_8646,N_8497,N_8418);
nand U8647 (N_8647,N_8463,N_8443);
xnor U8648 (N_8648,N_8504,N_8545);
nor U8649 (N_8649,N_8419,N_8496);
xnor U8650 (N_8650,N_8456,N_8473);
xor U8651 (N_8651,N_8419,N_8484);
xnor U8652 (N_8652,N_8546,N_8528);
xnor U8653 (N_8653,N_8407,N_8435);
and U8654 (N_8654,N_8423,N_8511);
nand U8655 (N_8655,N_8445,N_8456);
nor U8656 (N_8656,N_8423,N_8532);
xnor U8657 (N_8657,N_8475,N_8514);
nand U8658 (N_8658,N_8490,N_8527);
nand U8659 (N_8659,N_8410,N_8536);
and U8660 (N_8660,N_8511,N_8542);
xor U8661 (N_8661,N_8407,N_8537);
xnor U8662 (N_8662,N_8487,N_8423);
xor U8663 (N_8663,N_8408,N_8415);
nand U8664 (N_8664,N_8402,N_8531);
xnor U8665 (N_8665,N_8529,N_8543);
or U8666 (N_8666,N_8410,N_8506);
xor U8667 (N_8667,N_8401,N_8487);
or U8668 (N_8668,N_8407,N_8423);
xnor U8669 (N_8669,N_8545,N_8524);
nand U8670 (N_8670,N_8516,N_8448);
or U8671 (N_8671,N_8467,N_8531);
nand U8672 (N_8672,N_8411,N_8514);
xor U8673 (N_8673,N_8404,N_8544);
nor U8674 (N_8674,N_8515,N_8511);
and U8675 (N_8675,N_8429,N_8500);
xnor U8676 (N_8676,N_8463,N_8429);
or U8677 (N_8677,N_8478,N_8536);
and U8678 (N_8678,N_8433,N_8435);
nand U8679 (N_8679,N_8523,N_8466);
or U8680 (N_8680,N_8412,N_8534);
nand U8681 (N_8681,N_8440,N_8512);
nand U8682 (N_8682,N_8460,N_8527);
nor U8683 (N_8683,N_8488,N_8514);
nand U8684 (N_8684,N_8523,N_8475);
xnor U8685 (N_8685,N_8489,N_8466);
nor U8686 (N_8686,N_8478,N_8514);
and U8687 (N_8687,N_8501,N_8529);
or U8688 (N_8688,N_8410,N_8518);
nand U8689 (N_8689,N_8534,N_8441);
nor U8690 (N_8690,N_8439,N_8450);
nor U8691 (N_8691,N_8500,N_8446);
nand U8692 (N_8692,N_8446,N_8531);
or U8693 (N_8693,N_8453,N_8419);
and U8694 (N_8694,N_8500,N_8436);
or U8695 (N_8695,N_8479,N_8411);
and U8696 (N_8696,N_8482,N_8415);
or U8697 (N_8697,N_8449,N_8514);
xor U8698 (N_8698,N_8546,N_8428);
or U8699 (N_8699,N_8435,N_8453);
nor U8700 (N_8700,N_8566,N_8613);
nor U8701 (N_8701,N_8685,N_8640);
or U8702 (N_8702,N_8648,N_8610);
xnor U8703 (N_8703,N_8553,N_8568);
or U8704 (N_8704,N_8583,N_8570);
and U8705 (N_8705,N_8683,N_8666);
and U8706 (N_8706,N_8642,N_8647);
or U8707 (N_8707,N_8676,N_8605);
and U8708 (N_8708,N_8636,N_8607);
and U8709 (N_8709,N_8616,N_8585);
xor U8710 (N_8710,N_8580,N_8563);
nand U8711 (N_8711,N_8653,N_8635);
nand U8712 (N_8712,N_8630,N_8632);
and U8713 (N_8713,N_8620,N_8612);
nand U8714 (N_8714,N_8554,N_8697);
nor U8715 (N_8715,N_8550,N_8564);
nor U8716 (N_8716,N_8681,N_8565);
nand U8717 (N_8717,N_8567,N_8619);
nand U8718 (N_8718,N_8624,N_8586);
xnor U8719 (N_8719,N_8675,N_8573);
xnor U8720 (N_8720,N_8638,N_8598);
or U8721 (N_8721,N_8657,N_8695);
nor U8722 (N_8722,N_8599,N_8650);
nand U8723 (N_8723,N_8644,N_8628);
nor U8724 (N_8724,N_8561,N_8654);
or U8725 (N_8725,N_8631,N_8581);
or U8726 (N_8726,N_8688,N_8608);
xnor U8727 (N_8727,N_8668,N_8687);
nor U8728 (N_8728,N_8560,N_8555);
nor U8729 (N_8729,N_8667,N_8686);
or U8730 (N_8730,N_8595,N_8662);
xor U8731 (N_8731,N_8593,N_8627);
and U8732 (N_8732,N_8582,N_8614);
nand U8733 (N_8733,N_8634,N_8584);
and U8734 (N_8734,N_8575,N_8684);
or U8735 (N_8735,N_8626,N_8556);
and U8736 (N_8736,N_8574,N_8692);
xnor U8737 (N_8737,N_8661,N_8682);
and U8738 (N_8738,N_8629,N_8569);
nor U8739 (N_8739,N_8663,N_8588);
nand U8740 (N_8740,N_8698,N_8552);
nor U8741 (N_8741,N_8672,N_8699);
nor U8742 (N_8742,N_8617,N_8558);
nor U8743 (N_8743,N_8594,N_8618);
and U8744 (N_8744,N_8689,N_8591);
xnor U8745 (N_8745,N_8551,N_8645);
nor U8746 (N_8746,N_8633,N_8678);
or U8747 (N_8747,N_8670,N_8589);
or U8748 (N_8748,N_8649,N_8597);
and U8749 (N_8749,N_8673,N_8625);
and U8750 (N_8750,N_8646,N_8578);
or U8751 (N_8751,N_8696,N_8604);
or U8752 (N_8752,N_8623,N_8615);
nor U8753 (N_8753,N_8609,N_8665);
and U8754 (N_8754,N_8611,N_8621);
or U8755 (N_8755,N_8577,N_8557);
xnor U8756 (N_8756,N_8596,N_8590);
and U8757 (N_8757,N_8664,N_8679);
and U8758 (N_8758,N_8656,N_8677);
nand U8759 (N_8759,N_8674,N_8659);
xor U8760 (N_8760,N_8602,N_8652);
xor U8761 (N_8761,N_8592,N_8562);
or U8762 (N_8762,N_8660,N_8694);
or U8763 (N_8763,N_8643,N_8690);
or U8764 (N_8764,N_8579,N_8571);
nand U8765 (N_8765,N_8693,N_8587);
xor U8766 (N_8766,N_8655,N_8622);
nand U8767 (N_8767,N_8600,N_8637);
and U8768 (N_8768,N_8601,N_8691);
and U8769 (N_8769,N_8669,N_8606);
xor U8770 (N_8770,N_8680,N_8658);
xor U8771 (N_8771,N_8572,N_8639);
nand U8772 (N_8772,N_8651,N_8671);
nand U8773 (N_8773,N_8603,N_8559);
or U8774 (N_8774,N_8641,N_8576);
xor U8775 (N_8775,N_8629,N_8578);
and U8776 (N_8776,N_8616,N_8659);
xor U8777 (N_8777,N_8609,N_8571);
and U8778 (N_8778,N_8615,N_8564);
nand U8779 (N_8779,N_8554,N_8550);
and U8780 (N_8780,N_8660,N_8684);
or U8781 (N_8781,N_8568,N_8648);
nor U8782 (N_8782,N_8573,N_8630);
nor U8783 (N_8783,N_8555,N_8591);
nand U8784 (N_8784,N_8619,N_8559);
xor U8785 (N_8785,N_8576,N_8620);
nor U8786 (N_8786,N_8570,N_8591);
nor U8787 (N_8787,N_8653,N_8553);
and U8788 (N_8788,N_8696,N_8557);
or U8789 (N_8789,N_8636,N_8618);
and U8790 (N_8790,N_8671,N_8575);
and U8791 (N_8791,N_8596,N_8678);
nand U8792 (N_8792,N_8682,N_8623);
nor U8793 (N_8793,N_8589,N_8669);
nor U8794 (N_8794,N_8573,N_8624);
nand U8795 (N_8795,N_8568,N_8606);
nand U8796 (N_8796,N_8640,N_8564);
or U8797 (N_8797,N_8559,N_8659);
or U8798 (N_8798,N_8641,N_8683);
nor U8799 (N_8799,N_8625,N_8665);
and U8800 (N_8800,N_8675,N_8567);
xor U8801 (N_8801,N_8671,N_8613);
nor U8802 (N_8802,N_8667,N_8641);
nand U8803 (N_8803,N_8594,N_8652);
xnor U8804 (N_8804,N_8575,N_8570);
nor U8805 (N_8805,N_8611,N_8620);
nand U8806 (N_8806,N_8648,N_8590);
nor U8807 (N_8807,N_8660,N_8690);
or U8808 (N_8808,N_8555,N_8663);
nand U8809 (N_8809,N_8663,N_8566);
nor U8810 (N_8810,N_8675,N_8585);
or U8811 (N_8811,N_8594,N_8623);
or U8812 (N_8812,N_8682,N_8660);
nand U8813 (N_8813,N_8611,N_8675);
and U8814 (N_8814,N_8551,N_8591);
or U8815 (N_8815,N_8621,N_8668);
nor U8816 (N_8816,N_8565,N_8636);
and U8817 (N_8817,N_8633,N_8574);
and U8818 (N_8818,N_8622,N_8621);
nor U8819 (N_8819,N_8688,N_8600);
and U8820 (N_8820,N_8600,N_8555);
nor U8821 (N_8821,N_8611,N_8669);
and U8822 (N_8822,N_8610,N_8623);
or U8823 (N_8823,N_8600,N_8683);
nand U8824 (N_8824,N_8687,N_8622);
nor U8825 (N_8825,N_8690,N_8597);
nor U8826 (N_8826,N_8620,N_8658);
xnor U8827 (N_8827,N_8561,N_8575);
nand U8828 (N_8828,N_8565,N_8627);
or U8829 (N_8829,N_8583,N_8696);
xnor U8830 (N_8830,N_8579,N_8688);
and U8831 (N_8831,N_8560,N_8640);
nand U8832 (N_8832,N_8624,N_8600);
and U8833 (N_8833,N_8603,N_8698);
nor U8834 (N_8834,N_8690,N_8646);
nor U8835 (N_8835,N_8560,N_8566);
and U8836 (N_8836,N_8614,N_8654);
or U8837 (N_8837,N_8666,N_8575);
xnor U8838 (N_8838,N_8657,N_8642);
xor U8839 (N_8839,N_8679,N_8666);
or U8840 (N_8840,N_8598,N_8642);
nor U8841 (N_8841,N_8602,N_8611);
nor U8842 (N_8842,N_8695,N_8643);
or U8843 (N_8843,N_8589,N_8599);
nand U8844 (N_8844,N_8679,N_8552);
and U8845 (N_8845,N_8605,N_8677);
xnor U8846 (N_8846,N_8644,N_8599);
nand U8847 (N_8847,N_8596,N_8563);
nor U8848 (N_8848,N_8620,N_8622);
xor U8849 (N_8849,N_8642,N_8699);
or U8850 (N_8850,N_8807,N_8828);
and U8851 (N_8851,N_8790,N_8832);
or U8852 (N_8852,N_8801,N_8731);
xor U8853 (N_8853,N_8743,N_8838);
nand U8854 (N_8854,N_8730,N_8798);
nand U8855 (N_8855,N_8735,N_8806);
nor U8856 (N_8856,N_8826,N_8765);
and U8857 (N_8857,N_8830,N_8739);
and U8858 (N_8858,N_8726,N_8718);
nor U8859 (N_8859,N_8711,N_8837);
or U8860 (N_8860,N_8729,N_8782);
nand U8861 (N_8861,N_8804,N_8706);
or U8862 (N_8862,N_8833,N_8722);
nand U8863 (N_8863,N_8761,N_8840);
and U8864 (N_8864,N_8766,N_8797);
nand U8865 (N_8865,N_8750,N_8792);
nor U8866 (N_8866,N_8728,N_8768);
xor U8867 (N_8867,N_8709,N_8836);
nand U8868 (N_8868,N_8791,N_8755);
nand U8869 (N_8869,N_8841,N_8716);
nand U8870 (N_8870,N_8816,N_8784);
xor U8871 (N_8871,N_8762,N_8732);
nand U8872 (N_8872,N_8758,N_8700);
or U8873 (N_8873,N_8823,N_8745);
or U8874 (N_8874,N_8736,N_8829);
or U8875 (N_8875,N_8808,N_8834);
xor U8876 (N_8876,N_8819,N_8827);
or U8877 (N_8877,N_8835,N_8824);
and U8878 (N_8878,N_8714,N_8831);
xnor U8879 (N_8879,N_8733,N_8847);
xor U8880 (N_8880,N_8810,N_8770);
and U8881 (N_8881,N_8710,N_8751);
or U8882 (N_8882,N_8719,N_8725);
nand U8883 (N_8883,N_8849,N_8715);
or U8884 (N_8884,N_8809,N_8820);
nor U8885 (N_8885,N_8822,N_8779);
or U8886 (N_8886,N_8724,N_8846);
xor U8887 (N_8887,N_8708,N_8777);
xnor U8888 (N_8888,N_8821,N_8723);
and U8889 (N_8889,N_8813,N_8848);
xnor U8890 (N_8890,N_8760,N_8763);
xnor U8891 (N_8891,N_8844,N_8842);
or U8892 (N_8892,N_8752,N_8778);
or U8893 (N_8893,N_8812,N_8746);
or U8894 (N_8894,N_8774,N_8785);
or U8895 (N_8895,N_8817,N_8757);
nor U8896 (N_8896,N_8843,N_8759);
and U8897 (N_8897,N_8756,N_8717);
nand U8898 (N_8898,N_8720,N_8845);
xnor U8899 (N_8899,N_8707,N_8747);
xnor U8900 (N_8900,N_8769,N_8839);
or U8901 (N_8901,N_8803,N_8818);
nor U8902 (N_8902,N_8721,N_8793);
or U8903 (N_8903,N_8740,N_8795);
and U8904 (N_8904,N_8811,N_8825);
nor U8905 (N_8905,N_8799,N_8794);
or U8906 (N_8906,N_8702,N_8773);
nor U8907 (N_8907,N_8780,N_8767);
nor U8908 (N_8908,N_8805,N_8802);
nor U8909 (N_8909,N_8800,N_8753);
xnor U8910 (N_8910,N_8749,N_8781);
xor U8911 (N_8911,N_8815,N_8787);
xor U8912 (N_8912,N_8772,N_8789);
nand U8913 (N_8913,N_8713,N_8786);
and U8914 (N_8914,N_8703,N_8814);
or U8915 (N_8915,N_8748,N_8754);
and U8916 (N_8916,N_8701,N_8742);
nor U8917 (N_8917,N_8705,N_8775);
and U8918 (N_8918,N_8764,N_8788);
xnor U8919 (N_8919,N_8727,N_8741);
or U8920 (N_8920,N_8776,N_8771);
nor U8921 (N_8921,N_8796,N_8744);
nand U8922 (N_8922,N_8783,N_8734);
nand U8923 (N_8923,N_8738,N_8704);
nor U8924 (N_8924,N_8712,N_8737);
or U8925 (N_8925,N_8769,N_8722);
nor U8926 (N_8926,N_8761,N_8844);
or U8927 (N_8927,N_8731,N_8842);
nand U8928 (N_8928,N_8822,N_8803);
or U8929 (N_8929,N_8761,N_8756);
nor U8930 (N_8930,N_8833,N_8734);
nor U8931 (N_8931,N_8832,N_8730);
or U8932 (N_8932,N_8719,N_8771);
nand U8933 (N_8933,N_8795,N_8702);
and U8934 (N_8934,N_8731,N_8721);
and U8935 (N_8935,N_8716,N_8739);
nor U8936 (N_8936,N_8826,N_8716);
nand U8937 (N_8937,N_8822,N_8817);
xor U8938 (N_8938,N_8762,N_8801);
and U8939 (N_8939,N_8828,N_8754);
nand U8940 (N_8940,N_8794,N_8747);
and U8941 (N_8941,N_8756,N_8727);
nor U8942 (N_8942,N_8755,N_8718);
nand U8943 (N_8943,N_8712,N_8811);
or U8944 (N_8944,N_8828,N_8760);
and U8945 (N_8945,N_8723,N_8848);
nor U8946 (N_8946,N_8766,N_8749);
and U8947 (N_8947,N_8842,N_8726);
nor U8948 (N_8948,N_8733,N_8754);
nor U8949 (N_8949,N_8791,N_8757);
nor U8950 (N_8950,N_8798,N_8845);
nand U8951 (N_8951,N_8845,N_8789);
nor U8952 (N_8952,N_8713,N_8743);
or U8953 (N_8953,N_8791,N_8839);
nand U8954 (N_8954,N_8800,N_8702);
and U8955 (N_8955,N_8755,N_8771);
nor U8956 (N_8956,N_8711,N_8811);
nand U8957 (N_8957,N_8720,N_8780);
nor U8958 (N_8958,N_8769,N_8780);
nand U8959 (N_8959,N_8758,N_8723);
nor U8960 (N_8960,N_8741,N_8746);
or U8961 (N_8961,N_8706,N_8847);
nand U8962 (N_8962,N_8825,N_8833);
nand U8963 (N_8963,N_8722,N_8761);
nor U8964 (N_8964,N_8812,N_8766);
or U8965 (N_8965,N_8755,N_8826);
nor U8966 (N_8966,N_8762,N_8825);
or U8967 (N_8967,N_8766,N_8771);
or U8968 (N_8968,N_8806,N_8767);
xor U8969 (N_8969,N_8810,N_8803);
nor U8970 (N_8970,N_8840,N_8823);
nor U8971 (N_8971,N_8737,N_8796);
nor U8972 (N_8972,N_8759,N_8801);
nor U8973 (N_8973,N_8786,N_8716);
or U8974 (N_8974,N_8749,N_8780);
and U8975 (N_8975,N_8822,N_8829);
or U8976 (N_8976,N_8785,N_8763);
and U8977 (N_8977,N_8840,N_8718);
xnor U8978 (N_8978,N_8761,N_8706);
nand U8979 (N_8979,N_8723,N_8725);
and U8980 (N_8980,N_8707,N_8749);
nand U8981 (N_8981,N_8763,N_8820);
and U8982 (N_8982,N_8739,N_8782);
or U8983 (N_8983,N_8703,N_8783);
xnor U8984 (N_8984,N_8781,N_8839);
nor U8985 (N_8985,N_8836,N_8710);
xnor U8986 (N_8986,N_8832,N_8769);
or U8987 (N_8987,N_8840,N_8781);
and U8988 (N_8988,N_8754,N_8799);
nand U8989 (N_8989,N_8702,N_8701);
or U8990 (N_8990,N_8718,N_8795);
and U8991 (N_8991,N_8753,N_8718);
nand U8992 (N_8992,N_8702,N_8819);
nor U8993 (N_8993,N_8709,N_8788);
or U8994 (N_8994,N_8723,N_8704);
nor U8995 (N_8995,N_8824,N_8749);
and U8996 (N_8996,N_8739,N_8838);
nand U8997 (N_8997,N_8745,N_8768);
xor U8998 (N_8998,N_8718,N_8751);
nor U8999 (N_8999,N_8739,N_8810);
and U9000 (N_9000,N_8989,N_8990);
or U9001 (N_9001,N_8894,N_8995);
or U9002 (N_9002,N_8998,N_8982);
nand U9003 (N_9003,N_8933,N_8916);
xor U9004 (N_9004,N_8915,N_8867);
nand U9005 (N_9005,N_8859,N_8903);
xor U9006 (N_9006,N_8880,N_8968);
nand U9007 (N_9007,N_8925,N_8950);
nand U9008 (N_9008,N_8853,N_8871);
nor U9009 (N_9009,N_8908,N_8890);
xor U9010 (N_9010,N_8961,N_8897);
and U9011 (N_9011,N_8921,N_8924);
nand U9012 (N_9012,N_8955,N_8854);
or U9013 (N_9013,N_8910,N_8954);
or U9014 (N_9014,N_8943,N_8957);
xor U9015 (N_9015,N_8856,N_8860);
or U9016 (N_9016,N_8940,N_8918);
and U9017 (N_9017,N_8988,N_8947);
nor U9018 (N_9018,N_8953,N_8977);
nand U9019 (N_9019,N_8981,N_8979);
and U9020 (N_9020,N_8914,N_8978);
or U9021 (N_9021,N_8929,N_8934);
xnor U9022 (N_9022,N_8904,N_8923);
nand U9023 (N_9023,N_8858,N_8958);
or U9024 (N_9024,N_8949,N_8976);
or U9025 (N_9025,N_8899,N_8987);
and U9026 (N_9026,N_8999,N_8877);
xor U9027 (N_9027,N_8959,N_8872);
nor U9028 (N_9028,N_8851,N_8969);
xor U9029 (N_9029,N_8973,N_8935);
nor U9030 (N_9030,N_8932,N_8876);
xnor U9031 (N_9031,N_8928,N_8997);
and U9032 (N_9032,N_8975,N_8907);
nand U9033 (N_9033,N_8912,N_8937);
xor U9034 (N_9034,N_8956,N_8900);
nand U9035 (N_9035,N_8944,N_8893);
or U9036 (N_9036,N_8986,N_8920);
or U9037 (N_9037,N_8960,N_8855);
or U9038 (N_9038,N_8927,N_8974);
nand U9039 (N_9039,N_8906,N_8895);
and U9040 (N_9040,N_8971,N_8905);
nor U9041 (N_9041,N_8892,N_8902);
and U9042 (N_9042,N_8879,N_8922);
nor U9043 (N_9043,N_8862,N_8983);
or U9044 (N_9044,N_8868,N_8898);
nor U9045 (N_9045,N_8873,N_8883);
or U9046 (N_9046,N_8941,N_8970);
or U9047 (N_9047,N_8948,N_8966);
xor U9048 (N_9048,N_8861,N_8946);
or U9049 (N_9049,N_8913,N_8980);
xnor U9050 (N_9050,N_8984,N_8945);
and U9051 (N_9051,N_8952,N_8889);
or U9052 (N_9052,N_8992,N_8991);
or U9053 (N_9053,N_8887,N_8882);
or U9054 (N_9054,N_8896,N_8850);
nand U9055 (N_9055,N_8996,N_8863);
and U9056 (N_9056,N_8938,N_8936);
nor U9057 (N_9057,N_8886,N_8869);
nor U9058 (N_9058,N_8909,N_8901);
nand U9059 (N_9059,N_8993,N_8931);
or U9060 (N_9060,N_8852,N_8874);
or U9061 (N_9061,N_8875,N_8885);
or U9062 (N_9062,N_8911,N_8870);
or U9063 (N_9063,N_8963,N_8864);
nand U9064 (N_9064,N_8962,N_8857);
nor U9065 (N_9065,N_8866,N_8942);
or U9066 (N_9066,N_8888,N_8881);
nand U9067 (N_9067,N_8917,N_8939);
or U9068 (N_9068,N_8865,N_8967);
nor U9069 (N_9069,N_8972,N_8878);
and U9070 (N_9070,N_8930,N_8994);
or U9071 (N_9071,N_8985,N_8919);
or U9072 (N_9072,N_8951,N_8884);
nand U9073 (N_9073,N_8964,N_8926);
xor U9074 (N_9074,N_8891,N_8965);
xnor U9075 (N_9075,N_8935,N_8944);
or U9076 (N_9076,N_8978,N_8967);
or U9077 (N_9077,N_8893,N_8917);
or U9078 (N_9078,N_8934,N_8854);
nor U9079 (N_9079,N_8973,N_8895);
and U9080 (N_9080,N_8960,N_8911);
nor U9081 (N_9081,N_8896,N_8955);
and U9082 (N_9082,N_8895,N_8972);
or U9083 (N_9083,N_8954,N_8855);
nand U9084 (N_9084,N_8934,N_8997);
nor U9085 (N_9085,N_8874,N_8850);
xor U9086 (N_9086,N_8885,N_8888);
or U9087 (N_9087,N_8875,N_8870);
xor U9088 (N_9088,N_8982,N_8995);
or U9089 (N_9089,N_8905,N_8872);
xor U9090 (N_9090,N_8974,N_8950);
nor U9091 (N_9091,N_8965,N_8872);
nand U9092 (N_9092,N_8851,N_8915);
nand U9093 (N_9093,N_8927,N_8933);
and U9094 (N_9094,N_8944,N_8930);
nor U9095 (N_9095,N_8854,N_8943);
and U9096 (N_9096,N_8983,N_8903);
xnor U9097 (N_9097,N_8966,N_8922);
nor U9098 (N_9098,N_8928,N_8876);
nor U9099 (N_9099,N_8866,N_8893);
nand U9100 (N_9100,N_8908,N_8974);
nor U9101 (N_9101,N_8940,N_8930);
xnor U9102 (N_9102,N_8946,N_8901);
nand U9103 (N_9103,N_8960,N_8889);
and U9104 (N_9104,N_8958,N_8898);
or U9105 (N_9105,N_8929,N_8971);
nor U9106 (N_9106,N_8897,N_8950);
nor U9107 (N_9107,N_8981,N_8909);
nand U9108 (N_9108,N_8890,N_8981);
xor U9109 (N_9109,N_8925,N_8900);
xor U9110 (N_9110,N_8969,N_8901);
nor U9111 (N_9111,N_8873,N_8870);
xor U9112 (N_9112,N_8855,N_8919);
xor U9113 (N_9113,N_8926,N_8865);
and U9114 (N_9114,N_8897,N_8864);
or U9115 (N_9115,N_8911,N_8851);
or U9116 (N_9116,N_8966,N_8967);
xnor U9117 (N_9117,N_8902,N_8855);
nand U9118 (N_9118,N_8858,N_8989);
nand U9119 (N_9119,N_8958,N_8872);
and U9120 (N_9120,N_8931,N_8997);
or U9121 (N_9121,N_8985,N_8852);
xnor U9122 (N_9122,N_8947,N_8990);
and U9123 (N_9123,N_8906,N_8903);
xor U9124 (N_9124,N_8974,N_8889);
or U9125 (N_9125,N_8900,N_8862);
and U9126 (N_9126,N_8896,N_8943);
xnor U9127 (N_9127,N_8996,N_8940);
nand U9128 (N_9128,N_8852,N_8944);
nand U9129 (N_9129,N_8928,N_8924);
or U9130 (N_9130,N_8908,N_8984);
xor U9131 (N_9131,N_8893,N_8994);
nor U9132 (N_9132,N_8915,N_8981);
nand U9133 (N_9133,N_8892,N_8882);
or U9134 (N_9134,N_8939,N_8973);
and U9135 (N_9135,N_8959,N_8919);
xor U9136 (N_9136,N_8985,N_8969);
or U9137 (N_9137,N_8943,N_8906);
and U9138 (N_9138,N_8979,N_8954);
nor U9139 (N_9139,N_8943,N_8935);
xor U9140 (N_9140,N_8867,N_8962);
nand U9141 (N_9141,N_8902,N_8933);
nor U9142 (N_9142,N_8915,N_8927);
nor U9143 (N_9143,N_8953,N_8940);
nand U9144 (N_9144,N_8864,N_8891);
and U9145 (N_9145,N_8925,N_8947);
or U9146 (N_9146,N_8975,N_8912);
and U9147 (N_9147,N_8851,N_8863);
and U9148 (N_9148,N_8892,N_8885);
nand U9149 (N_9149,N_8881,N_8852);
and U9150 (N_9150,N_9006,N_9073);
or U9151 (N_9151,N_9116,N_9135);
nor U9152 (N_9152,N_9145,N_9061);
nor U9153 (N_9153,N_9088,N_9014);
or U9154 (N_9154,N_9031,N_9099);
nand U9155 (N_9155,N_9056,N_9075);
or U9156 (N_9156,N_9009,N_9059);
or U9157 (N_9157,N_9016,N_9032);
nand U9158 (N_9158,N_9047,N_9149);
nor U9159 (N_9159,N_9038,N_9008);
xnor U9160 (N_9160,N_9060,N_9139);
nand U9161 (N_9161,N_9003,N_9045);
xor U9162 (N_9162,N_9072,N_9052);
or U9163 (N_9163,N_9085,N_9122);
and U9164 (N_9164,N_9015,N_9025);
xnor U9165 (N_9165,N_9046,N_9082);
xnor U9166 (N_9166,N_9039,N_9078);
nor U9167 (N_9167,N_9097,N_9128);
nor U9168 (N_9168,N_9040,N_9053);
and U9169 (N_9169,N_9105,N_9034);
and U9170 (N_9170,N_9117,N_9069);
and U9171 (N_9171,N_9017,N_9120);
and U9172 (N_9172,N_9033,N_9143);
nor U9173 (N_9173,N_9104,N_9013);
and U9174 (N_9174,N_9030,N_9130);
and U9175 (N_9175,N_9129,N_9028);
nand U9176 (N_9176,N_9068,N_9044);
nor U9177 (N_9177,N_9111,N_9127);
nor U9178 (N_9178,N_9054,N_9140);
nor U9179 (N_9179,N_9050,N_9065);
nand U9180 (N_9180,N_9010,N_9066);
nor U9181 (N_9181,N_9022,N_9002);
nor U9182 (N_9182,N_9125,N_9123);
nand U9183 (N_9183,N_9110,N_9029);
xor U9184 (N_9184,N_9041,N_9051);
xor U9185 (N_9185,N_9000,N_9036);
nor U9186 (N_9186,N_9064,N_9087);
nor U9187 (N_9187,N_9011,N_9098);
nand U9188 (N_9188,N_9023,N_9035);
or U9189 (N_9189,N_9074,N_9077);
nor U9190 (N_9190,N_9037,N_9113);
and U9191 (N_9191,N_9070,N_9100);
and U9192 (N_9192,N_9118,N_9043);
or U9193 (N_9193,N_9142,N_9109);
and U9194 (N_9194,N_9055,N_9084);
nand U9195 (N_9195,N_9114,N_9094);
and U9196 (N_9196,N_9147,N_9063);
xor U9197 (N_9197,N_9136,N_9108);
xor U9198 (N_9198,N_9057,N_9096);
nand U9199 (N_9199,N_9021,N_9049);
or U9200 (N_9200,N_9090,N_9093);
nor U9201 (N_9201,N_9086,N_9076);
or U9202 (N_9202,N_9062,N_9081);
nor U9203 (N_9203,N_9079,N_9106);
nor U9204 (N_9204,N_9092,N_9048);
nand U9205 (N_9205,N_9134,N_9058);
xor U9206 (N_9206,N_9005,N_9119);
xor U9207 (N_9207,N_9112,N_9124);
or U9208 (N_9208,N_9080,N_9019);
xor U9209 (N_9209,N_9067,N_9137);
or U9210 (N_9210,N_9083,N_9027);
xnor U9211 (N_9211,N_9018,N_9107);
or U9212 (N_9212,N_9146,N_9144);
xor U9213 (N_9213,N_9042,N_9133);
xor U9214 (N_9214,N_9004,N_9121);
xnor U9215 (N_9215,N_9091,N_9141);
and U9216 (N_9216,N_9131,N_9132);
nand U9217 (N_9217,N_9020,N_9026);
or U9218 (N_9218,N_9138,N_9095);
nand U9219 (N_9219,N_9089,N_9102);
or U9220 (N_9220,N_9103,N_9115);
nand U9221 (N_9221,N_9024,N_9001);
and U9222 (N_9222,N_9012,N_9071);
or U9223 (N_9223,N_9101,N_9148);
nor U9224 (N_9224,N_9007,N_9126);
or U9225 (N_9225,N_9033,N_9097);
nor U9226 (N_9226,N_9032,N_9092);
nand U9227 (N_9227,N_9079,N_9124);
nor U9228 (N_9228,N_9116,N_9022);
or U9229 (N_9229,N_9019,N_9051);
or U9230 (N_9230,N_9007,N_9083);
and U9231 (N_9231,N_9011,N_9024);
and U9232 (N_9232,N_9076,N_9040);
and U9233 (N_9233,N_9023,N_9048);
nand U9234 (N_9234,N_9133,N_9136);
nand U9235 (N_9235,N_9020,N_9086);
and U9236 (N_9236,N_9052,N_9149);
or U9237 (N_9237,N_9004,N_9069);
nor U9238 (N_9238,N_9034,N_9118);
nor U9239 (N_9239,N_9036,N_9101);
nor U9240 (N_9240,N_9146,N_9118);
nor U9241 (N_9241,N_9135,N_9063);
nand U9242 (N_9242,N_9028,N_9120);
nor U9243 (N_9243,N_9149,N_9090);
or U9244 (N_9244,N_9122,N_9148);
and U9245 (N_9245,N_9021,N_9035);
nor U9246 (N_9246,N_9075,N_9130);
or U9247 (N_9247,N_9022,N_9038);
nor U9248 (N_9248,N_9137,N_9001);
or U9249 (N_9249,N_9075,N_9093);
nor U9250 (N_9250,N_9075,N_9057);
nand U9251 (N_9251,N_9023,N_9149);
or U9252 (N_9252,N_9060,N_9113);
nor U9253 (N_9253,N_9015,N_9001);
xor U9254 (N_9254,N_9037,N_9021);
nor U9255 (N_9255,N_9103,N_9089);
xnor U9256 (N_9256,N_9027,N_9085);
nand U9257 (N_9257,N_9070,N_9135);
xor U9258 (N_9258,N_9059,N_9085);
nand U9259 (N_9259,N_9146,N_9018);
nor U9260 (N_9260,N_9137,N_9013);
nand U9261 (N_9261,N_9086,N_9035);
and U9262 (N_9262,N_9118,N_9107);
or U9263 (N_9263,N_9065,N_9040);
or U9264 (N_9264,N_9052,N_9023);
nand U9265 (N_9265,N_9096,N_9081);
nand U9266 (N_9266,N_9011,N_9128);
and U9267 (N_9267,N_9003,N_9024);
or U9268 (N_9268,N_9069,N_9077);
nor U9269 (N_9269,N_9029,N_9001);
nor U9270 (N_9270,N_9123,N_9117);
or U9271 (N_9271,N_9096,N_9126);
and U9272 (N_9272,N_9098,N_9001);
xnor U9273 (N_9273,N_9051,N_9038);
xnor U9274 (N_9274,N_9118,N_9033);
nor U9275 (N_9275,N_9102,N_9119);
nor U9276 (N_9276,N_9106,N_9082);
xor U9277 (N_9277,N_9077,N_9065);
nor U9278 (N_9278,N_9123,N_9040);
nor U9279 (N_9279,N_9014,N_9119);
nand U9280 (N_9280,N_9023,N_9065);
and U9281 (N_9281,N_9022,N_9100);
nor U9282 (N_9282,N_9065,N_9048);
xnor U9283 (N_9283,N_9057,N_9042);
or U9284 (N_9284,N_9040,N_9138);
nor U9285 (N_9285,N_9040,N_9104);
and U9286 (N_9286,N_9001,N_9005);
xor U9287 (N_9287,N_9002,N_9118);
nand U9288 (N_9288,N_9132,N_9098);
nand U9289 (N_9289,N_9088,N_9054);
nand U9290 (N_9290,N_9050,N_9143);
xnor U9291 (N_9291,N_9000,N_9001);
nand U9292 (N_9292,N_9052,N_9138);
nand U9293 (N_9293,N_9023,N_9063);
xnor U9294 (N_9294,N_9129,N_9092);
or U9295 (N_9295,N_9114,N_9129);
and U9296 (N_9296,N_9147,N_9036);
xor U9297 (N_9297,N_9013,N_9043);
nand U9298 (N_9298,N_9113,N_9131);
or U9299 (N_9299,N_9001,N_9147);
and U9300 (N_9300,N_9188,N_9213);
and U9301 (N_9301,N_9177,N_9210);
nor U9302 (N_9302,N_9194,N_9268);
nand U9303 (N_9303,N_9150,N_9193);
nor U9304 (N_9304,N_9187,N_9294);
and U9305 (N_9305,N_9215,N_9165);
xor U9306 (N_9306,N_9296,N_9290);
and U9307 (N_9307,N_9250,N_9162);
nand U9308 (N_9308,N_9260,N_9183);
nor U9309 (N_9309,N_9209,N_9234);
nand U9310 (N_9310,N_9259,N_9202);
and U9311 (N_9311,N_9236,N_9151);
nand U9312 (N_9312,N_9153,N_9200);
nor U9313 (N_9313,N_9254,N_9217);
and U9314 (N_9314,N_9228,N_9273);
xor U9315 (N_9315,N_9241,N_9218);
or U9316 (N_9316,N_9174,N_9230);
xnor U9317 (N_9317,N_9163,N_9285);
nor U9318 (N_9318,N_9283,N_9212);
nor U9319 (N_9319,N_9261,N_9155);
and U9320 (N_9320,N_9157,N_9172);
or U9321 (N_9321,N_9189,N_9253);
nand U9322 (N_9322,N_9171,N_9208);
nand U9323 (N_9323,N_9258,N_9286);
or U9324 (N_9324,N_9180,N_9279);
xor U9325 (N_9325,N_9229,N_9179);
nor U9326 (N_9326,N_9225,N_9255);
nor U9327 (N_9327,N_9195,N_9167);
nor U9328 (N_9328,N_9198,N_9292);
nand U9329 (N_9329,N_9265,N_9223);
nor U9330 (N_9330,N_9299,N_9244);
xnor U9331 (N_9331,N_9161,N_9170);
or U9332 (N_9332,N_9262,N_9284);
or U9333 (N_9333,N_9275,N_9192);
nand U9334 (N_9334,N_9204,N_9247);
nor U9335 (N_9335,N_9211,N_9175);
or U9336 (N_9336,N_9152,N_9238);
and U9337 (N_9337,N_9278,N_9249);
nor U9338 (N_9338,N_9199,N_9173);
or U9339 (N_9339,N_9291,N_9186);
nor U9340 (N_9340,N_9272,N_9287);
and U9341 (N_9341,N_9164,N_9266);
xor U9342 (N_9342,N_9282,N_9295);
or U9343 (N_9343,N_9274,N_9156);
or U9344 (N_9344,N_9237,N_9169);
or U9345 (N_9345,N_9160,N_9226);
xnor U9346 (N_9346,N_9159,N_9248);
nor U9347 (N_9347,N_9219,N_9239);
or U9348 (N_9348,N_9191,N_9257);
xor U9349 (N_9349,N_9263,N_9158);
xor U9350 (N_9350,N_9297,N_9256);
xnor U9351 (N_9351,N_9205,N_9288);
xor U9352 (N_9352,N_9197,N_9182);
nor U9353 (N_9353,N_9196,N_9201);
or U9354 (N_9354,N_9251,N_9224);
and U9355 (N_9355,N_9166,N_9206);
nor U9356 (N_9356,N_9168,N_9271);
nor U9357 (N_9357,N_9231,N_9240);
nor U9358 (N_9358,N_9181,N_9176);
xnor U9359 (N_9359,N_9245,N_9233);
nand U9360 (N_9360,N_9185,N_9154);
or U9361 (N_9361,N_9235,N_9214);
and U9362 (N_9362,N_9222,N_9207);
xor U9363 (N_9363,N_9270,N_9277);
nand U9364 (N_9364,N_9298,N_9203);
nand U9365 (N_9365,N_9232,N_9220);
nand U9366 (N_9366,N_9221,N_9242);
or U9367 (N_9367,N_9293,N_9190);
nand U9368 (N_9368,N_9227,N_9281);
and U9369 (N_9369,N_9243,N_9264);
xnor U9370 (N_9370,N_9267,N_9269);
nand U9371 (N_9371,N_9276,N_9246);
nand U9372 (N_9372,N_9289,N_9184);
or U9373 (N_9373,N_9216,N_9280);
nand U9374 (N_9374,N_9252,N_9178);
nor U9375 (N_9375,N_9257,N_9245);
xor U9376 (N_9376,N_9232,N_9283);
nand U9377 (N_9377,N_9197,N_9223);
xnor U9378 (N_9378,N_9165,N_9198);
or U9379 (N_9379,N_9173,N_9156);
and U9380 (N_9380,N_9240,N_9254);
and U9381 (N_9381,N_9171,N_9221);
nand U9382 (N_9382,N_9255,N_9159);
nand U9383 (N_9383,N_9157,N_9185);
nor U9384 (N_9384,N_9181,N_9175);
nand U9385 (N_9385,N_9287,N_9264);
and U9386 (N_9386,N_9215,N_9226);
nand U9387 (N_9387,N_9221,N_9220);
xnor U9388 (N_9388,N_9217,N_9209);
nand U9389 (N_9389,N_9250,N_9215);
nand U9390 (N_9390,N_9173,N_9230);
and U9391 (N_9391,N_9185,N_9293);
nor U9392 (N_9392,N_9295,N_9156);
xor U9393 (N_9393,N_9269,N_9229);
xor U9394 (N_9394,N_9276,N_9188);
and U9395 (N_9395,N_9262,N_9201);
nor U9396 (N_9396,N_9296,N_9228);
xnor U9397 (N_9397,N_9226,N_9271);
nor U9398 (N_9398,N_9269,N_9258);
xor U9399 (N_9399,N_9239,N_9159);
nand U9400 (N_9400,N_9271,N_9159);
nand U9401 (N_9401,N_9291,N_9298);
or U9402 (N_9402,N_9238,N_9154);
xor U9403 (N_9403,N_9256,N_9277);
xor U9404 (N_9404,N_9188,N_9184);
nor U9405 (N_9405,N_9212,N_9273);
and U9406 (N_9406,N_9177,N_9268);
nand U9407 (N_9407,N_9251,N_9284);
xor U9408 (N_9408,N_9184,N_9268);
xnor U9409 (N_9409,N_9224,N_9167);
or U9410 (N_9410,N_9258,N_9249);
or U9411 (N_9411,N_9261,N_9238);
nor U9412 (N_9412,N_9253,N_9249);
nand U9413 (N_9413,N_9224,N_9234);
and U9414 (N_9414,N_9205,N_9177);
nand U9415 (N_9415,N_9168,N_9153);
or U9416 (N_9416,N_9150,N_9167);
and U9417 (N_9417,N_9222,N_9244);
nor U9418 (N_9418,N_9235,N_9240);
nor U9419 (N_9419,N_9297,N_9243);
xnor U9420 (N_9420,N_9260,N_9205);
xor U9421 (N_9421,N_9261,N_9227);
or U9422 (N_9422,N_9179,N_9243);
or U9423 (N_9423,N_9221,N_9293);
nand U9424 (N_9424,N_9253,N_9266);
or U9425 (N_9425,N_9265,N_9234);
xor U9426 (N_9426,N_9227,N_9213);
or U9427 (N_9427,N_9258,N_9247);
nor U9428 (N_9428,N_9290,N_9206);
or U9429 (N_9429,N_9227,N_9161);
nand U9430 (N_9430,N_9167,N_9174);
and U9431 (N_9431,N_9246,N_9189);
nor U9432 (N_9432,N_9288,N_9183);
nand U9433 (N_9433,N_9240,N_9207);
or U9434 (N_9434,N_9232,N_9204);
nand U9435 (N_9435,N_9156,N_9289);
nand U9436 (N_9436,N_9211,N_9195);
xor U9437 (N_9437,N_9168,N_9263);
nor U9438 (N_9438,N_9204,N_9162);
nand U9439 (N_9439,N_9281,N_9245);
nand U9440 (N_9440,N_9156,N_9204);
xnor U9441 (N_9441,N_9210,N_9248);
and U9442 (N_9442,N_9261,N_9187);
xor U9443 (N_9443,N_9242,N_9154);
and U9444 (N_9444,N_9198,N_9218);
nor U9445 (N_9445,N_9182,N_9163);
xor U9446 (N_9446,N_9199,N_9237);
nand U9447 (N_9447,N_9189,N_9192);
nor U9448 (N_9448,N_9254,N_9236);
and U9449 (N_9449,N_9268,N_9298);
nand U9450 (N_9450,N_9381,N_9434);
and U9451 (N_9451,N_9405,N_9309);
and U9452 (N_9452,N_9448,N_9386);
and U9453 (N_9453,N_9356,N_9417);
or U9454 (N_9454,N_9332,N_9312);
nor U9455 (N_9455,N_9326,N_9371);
and U9456 (N_9456,N_9366,N_9330);
and U9457 (N_9457,N_9317,N_9430);
nor U9458 (N_9458,N_9337,N_9398);
nand U9459 (N_9459,N_9435,N_9313);
nand U9460 (N_9460,N_9394,N_9319);
nand U9461 (N_9461,N_9302,N_9431);
nand U9462 (N_9462,N_9401,N_9373);
or U9463 (N_9463,N_9389,N_9377);
xnor U9464 (N_9464,N_9374,N_9304);
and U9465 (N_9465,N_9409,N_9367);
or U9466 (N_9466,N_9387,N_9437);
nor U9467 (N_9467,N_9439,N_9449);
xnor U9468 (N_9468,N_9442,N_9412);
or U9469 (N_9469,N_9445,N_9347);
nand U9470 (N_9470,N_9402,N_9426);
nand U9471 (N_9471,N_9329,N_9429);
and U9472 (N_9472,N_9403,N_9399);
xnor U9473 (N_9473,N_9425,N_9310);
or U9474 (N_9474,N_9404,N_9415);
xor U9475 (N_9475,N_9339,N_9393);
or U9476 (N_9476,N_9358,N_9408);
and U9477 (N_9477,N_9359,N_9352);
and U9478 (N_9478,N_9341,N_9418);
xor U9479 (N_9479,N_9413,N_9363);
or U9480 (N_9480,N_9335,N_9385);
nor U9481 (N_9481,N_9416,N_9443);
xnor U9482 (N_9482,N_9305,N_9349);
xnor U9483 (N_9483,N_9361,N_9414);
nor U9484 (N_9484,N_9348,N_9384);
nor U9485 (N_9485,N_9307,N_9438);
xnor U9486 (N_9486,N_9383,N_9395);
xor U9487 (N_9487,N_9325,N_9355);
or U9488 (N_9488,N_9379,N_9391);
or U9489 (N_9489,N_9362,N_9316);
and U9490 (N_9490,N_9400,N_9397);
or U9491 (N_9491,N_9441,N_9407);
or U9492 (N_9492,N_9370,N_9350);
nor U9493 (N_9493,N_9376,N_9343);
or U9494 (N_9494,N_9372,N_9322);
and U9495 (N_9495,N_9432,N_9396);
xnor U9496 (N_9496,N_9331,N_9336);
nor U9497 (N_9497,N_9423,N_9433);
nor U9498 (N_9498,N_9420,N_9380);
nand U9499 (N_9499,N_9424,N_9300);
nor U9500 (N_9500,N_9388,N_9436);
xnor U9501 (N_9501,N_9345,N_9422);
and U9502 (N_9502,N_9421,N_9406);
and U9503 (N_9503,N_9314,N_9365);
nand U9504 (N_9504,N_9328,N_9357);
xor U9505 (N_9505,N_9323,N_9410);
nand U9506 (N_9506,N_9447,N_9419);
nand U9507 (N_9507,N_9321,N_9303);
nand U9508 (N_9508,N_9444,N_9320);
xor U9509 (N_9509,N_9340,N_9368);
xnor U9510 (N_9510,N_9378,N_9308);
nand U9511 (N_9511,N_9327,N_9428);
nand U9512 (N_9512,N_9324,N_9392);
and U9513 (N_9513,N_9318,N_9346);
nor U9514 (N_9514,N_9382,N_9338);
and U9515 (N_9515,N_9311,N_9334);
and U9516 (N_9516,N_9344,N_9427);
or U9517 (N_9517,N_9375,N_9315);
and U9518 (N_9518,N_9354,N_9333);
nor U9519 (N_9519,N_9411,N_9342);
xnor U9520 (N_9520,N_9390,N_9440);
nor U9521 (N_9521,N_9364,N_9301);
or U9522 (N_9522,N_9306,N_9353);
xor U9523 (N_9523,N_9369,N_9446);
or U9524 (N_9524,N_9360,N_9351);
xnor U9525 (N_9525,N_9399,N_9449);
nand U9526 (N_9526,N_9361,N_9436);
and U9527 (N_9527,N_9366,N_9361);
nor U9528 (N_9528,N_9398,N_9413);
nor U9529 (N_9529,N_9342,N_9369);
xor U9530 (N_9530,N_9362,N_9396);
and U9531 (N_9531,N_9310,N_9388);
nand U9532 (N_9532,N_9429,N_9315);
nor U9533 (N_9533,N_9350,N_9426);
nor U9534 (N_9534,N_9306,N_9402);
nand U9535 (N_9535,N_9421,N_9433);
or U9536 (N_9536,N_9441,N_9355);
xnor U9537 (N_9537,N_9408,N_9370);
xor U9538 (N_9538,N_9324,N_9332);
nand U9539 (N_9539,N_9327,N_9334);
nand U9540 (N_9540,N_9418,N_9382);
nand U9541 (N_9541,N_9327,N_9348);
or U9542 (N_9542,N_9426,N_9435);
and U9543 (N_9543,N_9345,N_9372);
or U9544 (N_9544,N_9436,N_9329);
and U9545 (N_9545,N_9421,N_9302);
and U9546 (N_9546,N_9406,N_9449);
nand U9547 (N_9547,N_9403,N_9435);
nor U9548 (N_9548,N_9393,N_9317);
nor U9549 (N_9549,N_9350,N_9325);
nand U9550 (N_9550,N_9310,N_9363);
and U9551 (N_9551,N_9392,N_9330);
nand U9552 (N_9552,N_9412,N_9374);
and U9553 (N_9553,N_9392,N_9365);
or U9554 (N_9554,N_9428,N_9409);
and U9555 (N_9555,N_9310,N_9417);
xor U9556 (N_9556,N_9358,N_9371);
or U9557 (N_9557,N_9342,N_9410);
and U9558 (N_9558,N_9312,N_9342);
or U9559 (N_9559,N_9437,N_9364);
and U9560 (N_9560,N_9319,N_9360);
nor U9561 (N_9561,N_9363,N_9423);
and U9562 (N_9562,N_9314,N_9435);
nand U9563 (N_9563,N_9441,N_9410);
or U9564 (N_9564,N_9393,N_9341);
xnor U9565 (N_9565,N_9416,N_9364);
or U9566 (N_9566,N_9411,N_9365);
xnor U9567 (N_9567,N_9388,N_9331);
nand U9568 (N_9568,N_9432,N_9347);
nor U9569 (N_9569,N_9332,N_9355);
nor U9570 (N_9570,N_9370,N_9355);
xor U9571 (N_9571,N_9355,N_9395);
and U9572 (N_9572,N_9390,N_9325);
xnor U9573 (N_9573,N_9394,N_9301);
nor U9574 (N_9574,N_9360,N_9392);
or U9575 (N_9575,N_9406,N_9389);
xnor U9576 (N_9576,N_9411,N_9408);
and U9577 (N_9577,N_9337,N_9416);
or U9578 (N_9578,N_9333,N_9347);
and U9579 (N_9579,N_9360,N_9355);
or U9580 (N_9580,N_9379,N_9387);
nor U9581 (N_9581,N_9371,N_9447);
or U9582 (N_9582,N_9343,N_9413);
or U9583 (N_9583,N_9419,N_9358);
and U9584 (N_9584,N_9415,N_9326);
xnor U9585 (N_9585,N_9391,N_9434);
nand U9586 (N_9586,N_9337,N_9339);
or U9587 (N_9587,N_9379,N_9338);
nor U9588 (N_9588,N_9343,N_9358);
nor U9589 (N_9589,N_9337,N_9381);
xor U9590 (N_9590,N_9410,N_9371);
and U9591 (N_9591,N_9443,N_9357);
nand U9592 (N_9592,N_9353,N_9329);
xnor U9593 (N_9593,N_9386,N_9357);
and U9594 (N_9594,N_9412,N_9370);
nand U9595 (N_9595,N_9425,N_9341);
xnor U9596 (N_9596,N_9340,N_9443);
nor U9597 (N_9597,N_9346,N_9419);
and U9598 (N_9598,N_9387,N_9413);
or U9599 (N_9599,N_9398,N_9319);
xor U9600 (N_9600,N_9591,N_9534);
or U9601 (N_9601,N_9458,N_9554);
or U9602 (N_9602,N_9575,N_9578);
or U9603 (N_9603,N_9582,N_9490);
nand U9604 (N_9604,N_9527,N_9595);
nor U9605 (N_9605,N_9480,N_9492);
nand U9606 (N_9606,N_9476,N_9455);
and U9607 (N_9607,N_9486,N_9497);
nand U9608 (N_9608,N_9460,N_9545);
nand U9609 (N_9609,N_9518,N_9589);
or U9610 (N_9610,N_9574,N_9462);
nand U9611 (N_9611,N_9576,N_9596);
xor U9612 (N_9612,N_9503,N_9464);
or U9613 (N_9613,N_9547,N_9572);
xor U9614 (N_9614,N_9590,N_9469);
xor U9615 (N_9615,N_9568,N_9569);
and U9616 (N_9616,N_9548,N_9550);
nor U9617 (N_9617,N_9451,N_9535);
or U9618 (N_9618,N_9481,N_9533);
and U9619 (N_9619,N_9473,N_9511);
nand U9620 (N_9620,N_9453,N_9496);
or U9621 (N_9621,N_9594,N_9501);
or U9622 (N_9622,N_9472,N_9489);
nor U9623 (N_9623,N_9459,N_9468);
nand U9624 (N_9624,N_9514,N_9512);
or U9625 (N_9625,N_9493,N_9463);
nand U9626 (N_9626,N_9456,N_9517);
xor U9627 (N_9627,N_9592,N_9452);
nand U9628 (N_9628,N_9539,N_9524);
or U9629 (N_9629,N_9474,N_9552);
nor U9630 (N_9630,N_9507,N_9537);
xnor U9631 (N_9631,N_9483,N_9586);
nor U9632 (N_9632,N_9454,N_9544);
nand U9633 (N_9633,N_9488,N_9504);
nor U9634 (N_9634,N_9487,N_9502);
nand U9635 (N_9635,N_9556,N_9543);
nor U9636 (N_9636,N_9580,N_9581);
nor U9637 (N_9637,N_9515,N_9553);
nor U9638 (N_9638,N_9494,N_9523);
and U9639 (N_9639,N_9529,N_9526);
and U9640 (N_9640,N_9506,N_9482);
nor U9641 (N_9641,N_9467,N_9465);
nand U9642 (N_9642,N_9479,N_9520);
and U9643 (N_9643,N_9565,N_9519);
xor U9644 (N_9644,N_9560,N_9557);
xnor U9645 (N_9645,N_9531,N_9457);
xnor U9646 (N_9646,N_9563,N_9571);
xnor U9647 (N_9647,N_9521,N_9477);
and U9648 (N_9648,N_9471,N_9567);
or U9649 (N_9649,N_9484,N_9525);
xor U9650 (N_9650,N_9516,N_9593);
xor U9651 (N_9651,N_9499,N_9561);
and U9652 (N_9652,N_9478,N_9584);
and U9653 (N_9653,N_9542,N_9546);
nor U9654 (N_9654,N_9536,N_9588);
nand U9655 (N_9655,N_9562,N_9495);
or U9656 (N_9656,N_9491,N_9530);
or U9657 (N_9657,N_9498,N_9461);
nor U9658 (N_9658,N_9587,N_9538);
xor U9659 (N_9659,N_9558,N_9540);
or U9660 (N_9660,N_9528,N_9551);
and U9661 (N_9661,N_9566,N_9577);
nor U9662 (N_9662,N_9510,N_9598);
xnor U9663 (N_9663,N_9564,N_9466);
nor U9664 (N_9664,N_9541,N_9500);
and U9665 (N_9665,N_9509,N_9597);
or U9666 (N_9666,N_9513,N_9470);
xor U9667 (N_9667,N_9450,N_9505);
and U9668 (N_9668,N_9585,N_9559);
nor U9669 (N_9669,N_9549,N_9570);
and U9670 (N_9670,N_9573,N_9599);
xnor U9671 (N_9671,N_9532,N_9485);
or U9672 (N_9672,N_9508,N_9522);
nor U9673 (N_9673,N_9579,N_9475);
nand U9674 (N_9674,N_9555,N_9583);
nor U9675 (N_9675,N_9476,N_9467);
nor U9676 (N_9676,N_9529,N_9516);
nand U9677 (N_9677,N_9572,N_9487);
and U9678 (N_9678,N_9577,N_9562);
nand U9679 (N_9679,N_9566,N_9476);
or U9680 (N_9680,N_9457,N_9468);
xor U9681 (N_9681,N_9474,N_9503);
xor U9682 (N_9682,N_9511,N_9534);
and U9683 (N_9683,N_9580,N_9487);
and U9684 (N_9684,N_9566,N_9580);
nor U9685 (N_9685,N_9533,N_9452);
and U9686 (N_9686,N_9586,N_9556);
nor U9687 (N_9687,N_9524,N_9577);
or U9688 (N_9688,N_9513,N_9581);
nor U9689 (N_9689,N_9547,N_9508);
xnor U9690 (N_9690,N_9461,N_9575);
nor U9691 (N_9691,N_9561,N_9452);
nand U9692 (N_9692,N_9455,N_9599);
or U9693 (N_9693,N_9546,N_9572);
xnor U9694 (N_9694,N_9538,N_9458);
xor U9695 (N_9695,N_9582,N_9488);
nand U9696 (N_9696,N_9499,N_9560);
xor U9697 (N_9697,N_9551,N_9495);
nand U9698 (N_9698,N_9466,N_9497);
xor U9699 (N_9699,N_9475,N_9559);
or U9700 (N_9700,N_9508,N_9561);
xor U9701 (N_9701,N_9523,N_9491);
or U9702 (N_9702,N_9544,N_9496);
and U9703 (N_9703,N_9540,N_9549);
and U9704 (N_9704,N_9555,N_9537);
nand U9705 (N_9705,N_9479,N_9541);
nor U9706 (N_9706,N_9592,N_9532);
xor U9707 (N_9707,N_9586,N_9577);
or U9708 (N_9708,N_9512,N_9567);
or U9709 (N_9709,N_9469,N_9536);
or U9710 (N_9710,N_9543,N_9567);
xor U9711 (N_9711,N_9574,N_9556);
xor U9712 (N_9712,N_9470,N_9523);
nand U9713 (N_9713,N_9462,N_9577);
nand U9714 (N_9714,N_9583,N_9526);
xnor U9715 (N_9715,N_9586,N_9570);
and U9716 (N_9716,N_9476,N_9483);
xnor U9717 (N_9717,N_9514,N_9471);
nor U9718 (N_9718,N_9506,N_9465);
nand U9719 (N_9719,N_9591,N_9576);
xnor U9720 (N_9720,N_9467,N_9523);
or U9721 (N_9721,N_9459,N_9590);
nor U9722 (N_9722,N_9548,N_9586);
xor U9723 (N_9723,N_9542,N_9530);
or U9724 (N_9724,N_9454,N_9535);
nor U9725 (N_9725,N_9527,N_9495);
and U9726 (N_9726,N_9590,N_9534);
and U9727 (N_9727,N_9559,N_9497);
or U9728 (N_9728,N_9475,N_9539);
nand U9729 (N_9729,N_9543,N_9522);
xnor U9730 (N_9730,N_9511,N_9547);
or U9731 (N_9731,N_9451,N_9455);
nand U9732 (N_9732,N_9573,N_9534);
or U9733 (N_9733,N_9467,N_9595);
nand U9734 (N_9734,N_9490,N_9581);
or U9735 (N_9735,N_9465,N_9567);
and U9736 (N_9736,N_9462,N_9490);
or U9737 (N_9737,N_9499,N_9482);
nand U9738 (N_9738,N_9583,N_9566);
or U9739 (N_9739,N_9525,N_9476);
nand U9740 (N_9740,N_9589,N_9456);
xnor U9741 (N_9741,N_9545,N_9463);
xnor U9742 (N_9742,N_9539,N_9499);
nand U9743 (N_9743,N_9595,N_9506);
xnor U9744 (N_9744,N_9505,N_9500);
and U9745 (N_9745,N_9484,N_9589);
and U9746 (N_9746,N_9552,N_9533);
or U9747 (N_9747,N_9529,N_9592);
nor U9748 (N_9748,N_9460,N_9570);
and U9749 (N_9749,N_9481,N_9512);
or U9750 (N_9750,N_9697,N_9685);
xor U9751 (N_9751,N_9649,N_9735);
and U9752 (N_9752,N_9601,N_9747);
nand U9753 (N_9753,N_9722,N_9602);
nand U9754 (N_9754,N_9698,N_9620);
nor U9755 (N_9755,N_9623,N_9640);
and U9756 (N_9756,N_9712,N_9652);
nand U9757 (N_9757,N_9707,N_9713);
nor U9758 (N_9758,N_9714,N_9689);
nor U9759 (N_9759,N_9608,N_9607);
xnor U9760 (N_9760,N_9727,N_9661);
nor U9761 (N_9761,N_9672,N_9673);
and U9762 (N_9762,N_9663,N_9674);
or U9763 (N_9763,N_9635,N_9637);
nor U9764 (N_9764,N_9739,N_9636);
or U9765 (N_9765,N_9730,N_9613);
nand U9766 (N_9766,N_9702,N_9627);
and U9767 (N_9767,N_9671,N_9703);
or U9768 (N_9768,N_9619,N_9614);
nor U9769 (N_9769,N_9741,N_9655);
xnor U9770 (N_9770,N_9669,N_9633);
xnor U9771 (N_9771,N_9676,N_9654);
nand U9772 (N_9772,N_9686,N_9736);
or U9773 (N_9773,N_9650,N_9610);
xor U9774 (N_9774,N_9677,N_9704);
and U9775 (N_9775,N_9681,N_9630);
and U9776 (N_9776,N_9600,N_9734);
xnor U9777 (N_9777,N_9744,N_9638);
or U9778 (N_9778,N_9748,N_9729);
or U9779 (N_9779,N_9706,N_9675);
and U9780 (N_9780,N_9615,N_9603);
nand U9781 (N_9781,N_9721,N_9631);
nand U9782 (N_9782,N_9643,N_9621);
and U9783 (N_9783,N_9645,N_9738);
xor U9784 (N_9784,N_9626,N_9653);
and U9785 (N_9785,N_9646,N_9670);
and U9786 (N_9786,N_9648,N_9737);
nor U9787 (N_9787,N_9732,N_9746);
nor U9788 (N_9788,N_9667,N_9624);
and U9789 (N_9789,N_9651,N_9700);
and U9790 (N_9790,N_9705,N_9743);
and U9791 (N_9791,N_9668,N_9726);
nand U9792 (N_9792,N_9612,N_9666);
or U9793 (N_9793,N_9695,N_9690);
xor U9794 (N_9794,N_9680,N_9684);
nor U9795 (N_9795,N_9644,N_9609);
and U9796 (N_9796,N_9682,N_9647);
xnor U9797 (N_9797,N_9733,N_9665);
xor U9798 (N_9798,N_9628,N_9659);
nand U9799 (N_9799,N_9618,N_9731);
xor U9800 (N_9800,N_9641,N_9718);
nand U9801 (N_9801,N_9740,N_9694);
or U9802 (N_9802,N_9692,N_9656);
nand U9803 (N_9803,N_9724,N_9723);
nand U9804 (N_9804,N_9605,N_9604);
nand U9805 (N_9805,N_9622,N_9716);
xnor U9806 (N_9806,N_9745,N_9696);
and U9807 (N_9807,N_9639,N_9657);
nand U9808 (N_9808,N_9725,N_9617);
and U9809 (N_9809,N_9611,N_9711);
nand U9810 (N_9810,N_9710,N_9691);
nand U9811 (N_9811,N_9708,N_9720);
nand U9812 (N_9812,N_9717,N_9715);
nand U9813 (N_9813,N_9660,N_9625);
and U9814 (N_9814,N_9642,N_9688);
nand U9815 (N_9815,N_9749,N_9606);
nand U9816 (N_9816,N_9699,N_9632);
xnor U9817 (N_9817,N_9658,N_9719);
and U9818 (N_9818,N_9662,N_9709);
or U9819 (N_9819,N_9683,N_9728);
xor U9820 (N_9820,N_9742,N_9687);
and U9821 (N_9821,N_9679,N_9616);
nor U9822 (N_9822,N_9634,N_9693);
nand U9823 (N_9823,N_9701,N_9664);
nor U9824 (N_9824,N_9629,N_9678);
nor U9825 (N_9825,N_9611,N_9602);
nor U9826 (N_9826,N_9634,N_9671);
nand U9827 (N_9827,N_9649,N_9718);
and U9828 (N_9828,N_9659,N_9609);
or U9829 (N_9829,N_9646,N_9621);
nand U9830 (N_9830,N_9652,N_9651);
or U9831 (N_9831,N_9749,N_9691);
or U9832 (N_9832,N_9642,N_9644);
and U9833 (N_9833,N_9728,N_9643);
and U9834 (N_9834,N_9668,N_9680);
and U9835 (N_9835,N_9687,N_9601);
nor U9836 (N_9836,N_9710,N_9672);
or U9837 (N_9837,N_9671,N_9742);
nor U9838 (N_9838,N_9651,N_9717);
nor U9839 (N_9839,N_9669,N_9606);
xor U9840 (N_9840,N_9624,N_9678);
and U9841 (N_9841,N_9617,N_9656);
or U9842 (N_9842,N_9631,N_9705);
nand U9843 (N_9843,N_9628,N_9642);
xnor U9844 (N_9844,N_9740,N_9678);
nand U9845 (N_9845,N_9636,N_9702);
and U9846 (N_9846,N_9749,N_9655);
xor U9847 (N_9847,N_9725,N_9710);
and U9848 (N_9848,N_9691,N_9604);
and U9849 (N_9849,N_9646,N_9698);
xor U9850 (N_9850,N_9611,N_9621);
nor U9851 (N_9851,N_9737,N_9639);
or U9852 (N_9852,N_9647,N_9676);
or U9853 (N_9853,N_9656,N_9714);
or U9854 (N_9854,N_9675,N_9683);
and U9855 (N_9855,N_9607,N_9742);
nand U9856 (N_9856,N_9637,N_9743);
and U9857 (N_9857,N_9700,N_9632);
and U9858 (N_9858,N_9625,N_9609);
nand U9859 (N_9859,N_9635,N_9688);
or U9860 (N_9860,N_9621,N_9723);
xor U9861 (N_9861,N_9647,N_9686);
xnor U9862 (N_9862,N_9650,N_9742);
and U9863 (N_9863,N_9721,N_9717);
nand U9864 (N_9864,N_9654,N_9732);
nand U9865 (N_9865,N_9617,N_9704);
nand U9866 (N_9866,N_9660,N_9692);
nand U9867 (N_9867,N_9722,N_9676);
xnor U9868 (N_9868,N_9725,N_9748);
xnor U9869 (N_9869,N_9720,N_9722);
or U9870 (N_9870,N_9607,N_9703);
nor U9871 (N_9871,N_9721,N_9673);
and U9872 (N_9872,N_9603,N_9671);
xnor U9873 (N_9873,N_9739,N_9602);
xor U9874 (N_9874,N_9661,N_9742);
nand U9875 (N_9875,N_9659,N_9615);
or U9876 (N_9876,N_9714,N_9624);
xnor U9877 (N_9877,N_9609,N_9661);
or U9878 (N_9878,N_9749,N_9637);
xor U9879 (N_9879,N_9602,N_9632);
or U9880 (N_9880,N_9642,N_9704);
xnor U9881 (N_9881,N_9684,N_9606);
xor U9882 (N_9882,N_9649,N_9616);
nand U9883 (N_9883,N_9699,N_9706);
nor U9884 (N_9884,N_9683,N_9684);
nor U9885 (N_9885,N_9673,N_9748);
xor U9886 (N_9886,N_9645,N_9643);
xnor U9887 (N_9887,N_9723,N_9736);
and U9888 (N_9888,N_9749,N_9664);
and U9889 (N_9889,N_9617,N_9689);
nand U9890 (N_9890,N_9619,N_9682);
xnor U9891 (N_9891,N_9718,N_9726);
and U9892 (N_9892,N_9671,N_9617);
and U9893 (N_9893,N_9726,N_9742);
or U9894 (N_9894,N_9716,N_9673);
and U9895 (N_9895,N_9747,N_9650);
or U9896 (N_9896,N_9709,N_9616);
xor U9897 (N_9897,N_9694,N_9646);
nor U9898 (N_9898,N_9647,N_9657);
or U9899 (N_9899,N_9713,N_9693);
and U9900 (N_9900,N_9895,N_9812);
nor U9901 (N_9901,N_9779,N_9834);
nand U9902 (N_9902,N_9821,N_9766);
nor U9903 (N_9903,N_9769,N_9750);
xnor U9904 (N_9904,N_9878,N_9867);
xor U9905 (N_9905,N_9861,N_9877);
xnor U9906 (N_9906,N_9839,N_9848);
xor U9907 (N_9907,N_9862,N_9856);
nor U9908 (N_9908,N_9751,N_9891);
nor U9909 (N_9909,N_9800,N_9882);
or U9910 (N_9910,N_9775,N_9776);
nor U9911 (N_9911,N_9868,N_9801);
nand U9912 (N_9912,N_9825,N_9765);
nor U9913 (N_9913,N_9803,N_9767);
and U9914 (N_9914,N_9754,N_9889);
nand U9915 (N_9915,N_9756,N_9870);
and U9916 (N_9916,N_9817,N_9860);
xor U9917 (N_9917,N_9838,N_9781);
nand U9918 (N_9918,N_9855,N_9790);
nand U9919 (N_9919,N_9771,N_9850);
nor U9920 (N_9920,N_9824,N_9816);
nand U9921 (N_9921,N_9752,N_9755);
or U9922 (N_9922,N_9846,N_9871);
or U9923 (N_9923,N_9898,N_9854);
nor U9924 (N_9924,N_9884,N_9805);
or U9925 (N_9925,N_9883,N_9893);
xnor U9926 (N_9926,N_9836,N_9807);
nand U9927 (N_9927,N_9797,N_9793);
xor U9928 (N_9928,N_9822,N_9837);
xor U9929 (N_9929,N_9813,N_9880);
or U9930 (N_9930,N_9815,N_9760);
or U9931 (N_9931,N_9886,N_9758);
xor U9932 (N_9932,N_9874,N_9772);
nand U9933 (N_9933,N_9842,N_9892);
and U9934 (N_9934,N_9780,N_9827);
xor U9935 (N_9935,N_9764,N_9896);
xor U9936 (N_9936,N_9851,N_9863);
xor U9937 (N_9937,N_9762,N_9757);
or U9938 (N_9938,N_9872,N_9873);
nor U9939 (N_9939,N_9844,N_9823);
nor U9940 (N_9940,N_9876,N_9890);
nand U9941 (N_9941,N_9770,N_9864);
and U9942 (N_9942,N_9833,N_9782);
and U9943 (N_9943,N_9768,N_9879);
nor U9944 (N_9944,N_9753,N_9840);
xor U9945 (N_9945,N_9829,N_9852);
and U9946 (N_9946,N_9792,N_9875);
nor U9947 (N_9947,N_9784,N_9853);
xnor U9948 (N_9948,N_9798,N_9847);
or U9949 (N_9949,N_9778,N_9849);
nand U9950 (N_9950,N_9789,N_9897);
or U9951 (N_9951,N_9881,N_9819);
and U9952 (N_9952,N_9811,N_9899);
xor U9953 (N_9953,N_9808,N_9828);
nand U9954 (N_9954,N_9796,N_9759);
and U9955 (N_9955,N_9831,N_9859);
xnor U9956 (N_9956,N_9869,N_9787);
xor U9957 (N_9957,N_9809,N_9810);
or U9958 (N_9958,N_9761,N_9857);
and U9959 (N_9959,N_9818,N_9806);
nand U9960 (N_9960,N_9885,N_9788);
or U9961 (N_9961,N_9777,N_9865);
xnor U9962 (N_9962,N_9887,N_9785);
nand U9963 (N_9963,N_9799,N_9894);
and U9964 (N_9964,N_9843,N_9888);
and U9965 (N_9965,N_9794,N_9835);
nand U9966 (N_9966,N_9783,N_9804);
xor U9967 (N_9967,N_9858,N_9832);
nand U9968 (N_9968,N_9866,N_9841);
and U9969 (N_9969,N_9795,N_9786);
xor U9970 (N_9970,N_9763,N_9820);
or U9971 (N_9971,N_9791,N_9814);
nand U9972 (N_9972,N_9830,N_9845);
nor U9973 (N_9973,N_9826,N_9773);
or U9974 (N_9974,N_9802,N_9774);
nand U9975 (N_9975,N_9753,N_9854);
and U9976 (N_9976,N_9839,N_9834);
xnor U9977 (N_9977,N_9763,N_9823);
nor U9978 (N_9978,N_9797,N_9786);
or U9979 (N_9979,N_9784,N_9760);
and U9980 (N_9980,N_9762,N_9840);
or U9981 (N_9981,N_9872,N_9759);
nand U9982 (N_9982,N_9892,N_9845);
or U9983 (N_9983,N_9874,N_9832);
xnor U9984 (N_9984,N_9868,N_9796);
or U9985 (N_9985,N_9887,N_9830);
or U9986 (N_9986,N_9753,N_9893);
and U9987 (N_9987,N_9833,N_9811);
and U9988 (N_9988,N_9791,N_9857);
nand U9989 (N_9989,N_9808,N_9754);
xor U9990 (N_9990,N_9878,N_9781);
or U9991 (N_9991,N_9750,N_9751);
and U9992 (N_9992,N_9883,N_9837);
nor U9993 (N_9993,N_9886,N_9782);
or U9994 (N_9994,N_9861,N_9896);
nand U9995 (N_9995,N_9752,N_9816);
nand U9996 (N_9996,N_9837,N_9799);
xnor U9997 (N_9997,N_9867,N_9841);
xnor U9998 (N_9998,N_9862,N_9883);
xor U9999 (N_9999,N_9751,N_9818);
nand U10000 (N_10000,N_9859,N_9777);
and U10001 (N_10001,N_9761,N_9786);
nor U10002 (N_10002,N_9805,N_9794);
or U10003 (N_10003,N_9874,N_9885);
or U10004 (N_10004,N_9846,N_9781);
or U10005 (N_10005,N_9770,N_9797);
nor U10006 (N_10006,N_9832,N_9885);
and U10007 (N_10007,N_9878,N_9827);
nor U10008 (N_10008,N_9804,N_9780);
or U10009 (N_10009,N_9874,N_9755);
nor U10010 (N_10010,N_9792,N_9783);
or U10011 (N_10011,N_9875,N_9811);
nor U10012 (N_10012,N_9881,N_9761);
nor U10013 (N_10013,N_9850,N_9862);
nand U10014 (N_10014,N_9753,N_9778);
nand U10015 (N_10015,N_9826,N_9753);
nor U10016 (N_10016,N_9896,N_9815);
or U10017 (N_10017,N_9897,N_9794);
or U10018 (N_10018,N_9873,N_9802);
nand U10019 (N_10019,N_9843,N_9882);
nor U10020 (N_10020,N_9844,N_9875);
or U10021 (N_10021,N_9849,N_9781);
and U10022 (N_10022,N_9852,N_9830);
nand U10023 (N_10023,N_9804,N_9825);
nand U10024 (N_10024,N_9809,N_9818);
nand U10025 (N_10025,N_9816,N_9803);
and U10026 (N_10026,N_9791,N_9888);
xor U10027 (N_10027,N_9789,N_9762);
or U10028 (N_10028,N_9755,N_9778);
nor U10029 (N_10029,N_9887,N_9814);
or U10030 (N_10030,N_9792,N_9898);
xnor U10031 (N_10031,N_9765,N_9808);
or U10032 (N_10032,N_9881,N_9776);
or U10033 (N_10033,N_9752,N_9819);
nand U10034 (N_10034,N_9782,N_9885);
or U10035 (N_10035,N_9823,N_9802);
or U10036 (N_10036,N_9818,N_9834);
nand U10037 (N_10037,N_9853,N_9876);
nor U10038 (N_10038,N_9820,N_9782);
and U10039 (N_10039,N_9815,N_9822);
and U10040 (N_10040,N_9827,N_9898);
or U10041 (N_10041,N_9769,N_9822);
nor U10042 (N_10042,N_9816,N_9865);
nand U10043 (N_10043,N_9775,N_9756);
nor U10044 (N_10044,N_9832,N_9774);
nand U10045 (N_10045,N_9870,N_9834);
and U10046 (N_10046,N_9875,N_9860);
nand U10047 (N_10047,N_9834,N_9829);
and U10048 (N_10048,N_9760,N_9890);
or U10049 (N_10049,N_9796,N_9814);
xor U10050 (N_10050,N_9988,N_9906);
nand U10051 (N_10051,N_9979,N_9995);
nor U10052 (N_10052,N_10015,N_9966);
or U10053 (N_10053,N_10008,N_10011);
and U10054 (N_10054,N_10002,N_10012);
and U10055 (N_10055,N_10020,N_9918);
or U10056 (N_10056,N_9944,N_9964);
and U10057 (N_10057,N_10004,N_10049);
nor U10058 (N_10058,N_9977,N_10007);
nor U10059 (N_10059,N_9990,N_9986);
or U10060 (N_10060,N_9978,N_9915);
xnor U10061 (N_10061,N_10036,N_10040);
or U10062 (N_10062,N_9965,N_9958);
nand U10063 (N_10063,N_9972,N_10047);
or U10064 (N_10064,N_10043,N_9985);
or U10065 (N_10065,N_9920,N_10024);
nor U10066 (N_10066,N_10019,N_10029);
nand U10067 (N_10067,N_10038,N_9928);
or U10068 (N_10068,N_9922,N_9974);
or U10069 (N_10069,N_9931,N_10045);
nor U10070 (N_10070,N_9905,N_9923);
xor U10071 (N_10071,N_9942,N_10013);
or U10072 (N_10072,N_9952,N_9962);
nand U10073 (N_10073,N_9936,N_10027);
and U10074 (N_10074,N_9956,N_10026);
and U10075 (N_10075,N_9925,N_9902);
xnor U10076 (N_10076,N_9901,N_9954);
and U10077 (N_10077,N_9938,N_10010);
xor U10078 (N_10078,N_9950,N_9941);
and U10079 (N_10079,N_9933,N_9983);
nor U10080 (N_10080,N_10034,N_10022);
xnor U10081 (N_10081,N_10006,N_9907);
or U10082 (N_10082,N_9921,N_10044);
nor U10083 (N_10083,N_9980,N_9917);
or U10084 (N_10084,N_9968,N_9969);
nor U10085 (N_10085,N_9908,N_10017);
or U10086 (N_10086,N_10035,N_9912);
xor U10087 (N_10087,N_9989,N_10028);
and U10088 (N_10088,N_10001,N_9900);
nand U10089 (N_10089,N_9994,N_9926);
and U10090 (N_10090,N_10030,N_10041);
or U10091 (N_10091,N_10009,N_9982);
xor U10092 (N_10092,N_10031,N_10014);
and U10093 (N_10093,N_9996,N_9935);
nand U10094 (N_10094,N_9963,N_9949);
or U10095 (N_10095,N_9997,N_9932);
and U10096 (N_10096,N_9904,N_9913);
xor U10097 (N_10097,N_9959,N_9984);
xor U10098 (N_10098,N_9970,N_9946);
or U10099 (N_10099,N_9957,N_9903);
nand U10100 (N_10100,N_9945,N_9991);
or U10101 (N_10101,N_9909,N_9910);
nand U10102 (N_10102,N_9971,N_10003);
or U10103 (N_10103,N_9927,N_10042);
nor U10104 (N_10104,N_9929,N_9948);
xnor U10105 (N_10105,N_9975,N_9999);
xor U10106 (N_10106,N_9916,N_9981);
nor U10107 (N_10107,N_9939,N_10033);
and U10108 (N_10108,N_10018,N_10039);
and U10109 (N_10109,N_10021,N_9919);
nor U10110 (N_10110,N_9924,N_10000);
and U10111 (N_10111,N_9961,N_9943);
xnor U10112 (N_10112,N_9953,N_9947);
or U10113 (N_10113,N_10046,N_9951);
nand U10114 (N_10114,N_9934,N_10048);
nor U10115 (N_10115,N_9967,N_9993);
or U10116 (N_10116,N_9930,N_10032);
xnor U10117 (N_10117,N_9955,N_9911);
and U10118 (N_10118,N_10037,N_10025);
or U10119 (N_10119,N_9937,N_9940);
nor U10120 (N_10120,N_10016,N_9987);
and U10121 (N_10121,N_10005,N_9998);
and U10122 (N_10122,N_10023,N_9976);
nand U10123 (N_10123,N_9914,N_9992);
nor U10124 (N_10124,N_9973,N_9960);
xor U10125 (N_10125,N_9975,N_9956);
and U10126 (N_10126,N_10017,N_10029);
xor U10127 (N_10127,N_10032,N_9923);
xnor U10128 (N_10128,N_9945,N_9950);
nand U10129 (N_10129,N_10003,N_9910);
nand U10130 (N_10130,N_10042,N_9941);
nor U10131 (N_10131,N_10001,N_10042);
xor U10132 (N_10132,N_9962,N_9943);
nor U10133 (N_10133,N_10030,N_9980);
or U10134 (N_10134,N_9964,N_9958);
and U10135 (N_10135,N_10040,N_9983);
nor U10136 (N_10136,N_10048,N_9945);
xnor U10137 (N_10137,N_9936,N_9920);
nor U10138 (N_10138,N_9991,N_9916);
nand U10139 (N_10139,N_9965,N_10010);
xnor U10140 (N_10140,N_10014,N_9957);
nand U10141 (N_10141,N_9992,N_9993);
nand U10142 (N_10142,N_10028,N_9991);
or U10143 (N_10143,N_9971,N_9969);
nor U10144 (N_10144,N_10015,N_9934);
or U10145 (N_10145,N_9905,N_10015);
and U10146 (N_10146,N_9906,N_9901);
nor U10147 (N_10147,N_10015,N_9925);
xnor U10148 (N_10148,N_9952,N_9955);
nand U10149 (N_10149,N_10039,N_9968);
or U10150 (N_10150,N_9971,N_9981);
or U10151 (N_10151,N_9976,N_9981);
nand U10152 (N_10152,N_9988,N_9973);
and U10153 (N_10153,N_10026,N_9933);
xnor U10154 (N_10154,N_9960,N_10012);
and U10155 (N_10155,N_9978,N_10031);
and U10156 (N_10156,N_9948,N_10026);
nor U10157 (N_10157,N_9994,N_9924);
or U10158 (N_10158,N_9941,N_9977);
nor U10159 (N_10159,N_9929,N_10046);
or U10160 (N_10160,N_9958,N_10025);
and U10161 (N_10161,N_10022,N_9947);
nor U10162 (N_10162,N_9993,N_9976);
or U10163 (N_10163,N_9946,N_9935);
nor U10164 (N_10164,N_9985,N_10029);
or U10165 (N_10165,N_10007,N_10024);
or U10166 (N_10166,N_10031,N_10025);
xor U10167 (N_10167,N_10022,N_9949);
xnor U10168 (N_10168,N_10008,N_10042);
and U10169 (N_10169,N_9977,N_9921);
nor U10170 (N_10170,N_10023,N_9903);
or U10171 (N_10171,N_9918,N_9911);
nor U10172 (N_10172,N_10047,N_10032);
nand U10173 (N_10173,N_10008,N_9956);
and U10174 (N_10174,N_9991,N_9998);
or U10175 (N_10175,N_9984,N_9956);
and U10176 (N_10176,N_9962,N_9997);
nor U10177 (N_10177,N_10033,N_9918);
or U10178 (N_10178,N_10004,N_10029);
or U10179 (N_10179,N_9916,N_9928);
xnor U10180 (N_10180,N_10010,N_9926);
xnor U10181 (N_10181,N_9970,N_10005);
nand U10182 (N_10182,N_9976,N_9925);
and U10183 (N_10183,N_10025,N_10034);
or U10184 (N_10184,N_9970,N_10014);
xnor U10185 (N_10185,N_9919,N_10026);
nand U10186 (N_10186,N_9942,N_10044);
or U10187 (N_10187,N_10017,N_9998);
nor U10188 (N_10188,N_9932,N_9983);
nand U10189 (N_10189,N_9935,N_9962);
xor U10190 (N_10190,N_9956,N_10037);
or U10191 (N_10191,N_9913,N_10038);
xor U10192 (N_10192,N_9945,N_9979);
or U10193 (N_10193,N_9908,N_9975);
nor U10194 (N_10194,N_9921,N_9978);
nor U10195 (N_10195,N_10010,N_10017);
nand U10196 (N_10196,N_9982,N_9927);
nor U10197 (N_10197,N_9978,N_9970);
or U10198 (N_10198,N_10042,N_9984);
and U10199 (N_10199,N_9904,N_10031);
xnor U10200 (N_10200,N_10100,N_10121);
nor U10201 (N_10201,N_10151,N_10184);
xnor U10202 (N_10202,N_10185,N_10109);
and U10203 (N_10203,N_10131,N_10124);
nand U10204 (N_10204,N_10147,N_10191);
nand U10205 (N_10205,N_10066,N_10138);
and U10206 (N_10206,N_10143,N_10178);
nor U10207 (N_10207,N_10080,N_10064);
nor U10208 (N_10208,N_10194,N_10058);
or U10209 (N_10209,N_10174,N_10125);
or U10210 (N_10210,N_10189,N_10160);
nand U10211 (N_10211,N_10126,N_10148);
nor U10212 (N_10212,N_10144,N_10141);
nand U10213 (N_10213,N_10094,N_10116);
xor U10214 (N_10214,N_10068,N_10118);
xnor U10215 (N_10215,N_10106,N_10092);
or U10216 (N_10216,N_10107,N_10072);
or U10217 (N_10217,N_10054,N_10156);
and U10218 (N_10218,N_10087,N_10059);
nand U10219 (N_10219,N_10095,N_10098);
xnor U10220 (N_10220,N_10182,N_10154);
nand U10221 (N_10221,N_10103,N_10134);
or U10222 (N_10222,N_10056,N_10067);
and U10223 (N_10223,N_10161,N_10078);
nor U10224 (N_10224,N_10181,N_10173);
nor U10225 (N_10225,N_10165,N_10104);
xor U10226 (N_10226,N_10129,N_10153);
nand U10227 (N_10227,N_10128,N_10123);
xor U10228 (N_10228,N_10051,N_10079);
nand U10229 (N_10229,N_10145,N_10112);
nand U10230 (N_10230,N_10069,N_10164);
nor U10231 (N_10231,N_10115,N_10071);
and U10232 (N_10232,N_10130,N_10120);
or U10233 (N_10233,N_10169,N_10146);
xor U10234 (N_10234,N_10097,N_10090);
and U10235 (N_10235,N_10060,N_10177);
nor U10236 (N_10236,N_10190,N_10099);
nor U10237 (N_10237,N_10152,N_10162);
nor U10238 (N_10238,N_10199,N_10150);
xor U10239 (N_10239,N_10168,N_10083);
and U10240 (N_10240,N_10180,N_10075);
xor U10241 (N_10241,N_10166,N_10110);
xor U10242 (N_10242,N_10157,N_10187);
and U10243 (N_10243,N_10186,N_10073);
xnor U10244 (N_10244,N_10111,N_10093);
nor U10245 (N_10245,N_10061,N_10088);
and U10246 (N_10246,N_10065,N_10175);
and U10247 (N_10247,N_10133,N_10053);
xor U10248 (N_10248,N_10163,N_10122);
xnor U10249 (N_10249,N_10076,N_10135);
and U10250 (N_10250,N_10070,N_10091);
nor U10251 (N_10251,N_10149,N_10082);
or U10252 (N_10252,N_10055,N_10119);
nor U10253 (N_10253,N_10179,N_10081);
and U10254 (N_10254,N_10195,N_10062);
nor U10255 (N_10255,N_10137,N_10050);
nor U10256 (N_10256,N_10084,N_10183);
and U10257 (N_10257,N_10127,N_10167);
nor U10258 (N_10258,N_10114,N_10057);
or U10259 (N_10259,N_10136,N_10155);
or U10260 (N_10260,N_10101,N_10117);
or U10261 (N_10261,N_10196,N_10142);
nand U10262 (N_10262,N_10139,N_10198);
and U10263 (N_10263,N_10170,N_10132);
xor U10264 (N_10264,N_10108,N_10159);
nand U10265 (N_10265,N_10089,N_10188);
nand U10266 (N_10266,N_10172,N_10140);
nor U10267 (N_10267,N_10052,N_10096);
and U10268 (N_10268,N_10176,N_10158);
xnor U10269 (N_10269,N_10171,N_10063);
nor U10270 (N_10270,N_10077,N_10105);
or U10271 (N_10271,N_10086,N_10192);
nor U10272 (N_10272,N_10113,N_10193);
nor U10273 (N_10273,N_10197,N_10085);
xnor U10274 (N_10274,N_10074,N_10102);
nand U10275 (N_10275,N_10179,N_10067);
or U10276 (N_10276,N_10142,N_10186);
nor U10277 (N_10277,N_10130,N_10160);
xnor U10278 (N_10278,N_10100,N_10067);
xnor U10279 (N_10279,N_10176,N_10153);
and U10280 (N_10280,N_10110,N_10140);
xnor U10281 (N_10281,N_10161,N_10143);
nor U10282 (N_10282,N_10115,N_10166);
nand U10283 (N_10283,N_10122,N_10181);
or U10284 (N_10284,N_10082,N_10105);
and U10285 (N_10285,N_10105,N_10094);
xnor U10286 (N_10286,N_10116,N_10105);
or U10287 (N_10287,N_10178,N_10122);
nor U10288 (N_10288,N_10122,N_10130);
or U10289 (N_10289,N_10053,N_10161);
nand U10290 (N_10290,N_10057,N_10161);
or U10291 (N_10291,N_10155,N_10156);
or U10292 (N_10292,N_10086,N_10050);
nand U10293 (N_10293,N_10097,N_10056);
nor U10294 (N_10294,N_10051,N_10183);
nand U10295 (N_10295,N_10166,N_10190);
nand U10296 (N_10296,N_10050,N_10134);
and U10297 (N_10297,N_10191,N_10060);
and U10298 (N_10298,N_10050,N_10084);
and U10299 (N_10299,N_10127,N_10130);
or U10300 (N_10300,N_10148,N_10121);
xnor U10301 (N_10301,N_10140,N_10114);
nand U10302 (N_10302,N_10095,N_10072);
xnor U10303 (N_10303,N_10166,N_10095);
or U10304 (N_10304,N_10178,N_10088);
and U10305 (N_10305,N_10110,N_10133);
xor U10306 (N_10306,N_10135,N_10170);
or U10307 (N_10307,N_10177,N_10189);
xor U10308 (N_10308,N_10051,N_10060);
xnor U10309 (N_10309,N_10062,N_10051);
nor U10310 (N_10310,N_10132,N_10190);
and U10311 (N_10311,N_10097,N_10185);
nand U10312 (N_10312,N_10158,N_10081);
or U10313 (N_10313,N_10068,N_10133);
and U10314 (N_10314,N_10189,N_10057);
nor U10315 (N_10315,N_10103,N_10112);
nor U10316 (N_10316,N_10105,N_10184);
nand U10317 (N_10317,N_10058,N_10190);
nor U10318 (N_10318,N_10075,N_10149);
and U10319 (N_10319,N_10169,N_10197);
and U10320 (N_10320,N_10186,N_10156);
nand U10321 (N_10321,N_10175,N_10155);
nor U10322 (N_10322,N_10064,N_10156);
nor U10323 (N_10323,N_10197,N_10140);
nand U10324 (N_10324,N_10159,N_10107);
and U10325 (N_10325,N_10164,N_10161);
nor U10326 (N_10326,N_10141,N_10125);
xor U10327 (N_10327,N_10144,N_10054);
nand U10328 (N_10328,N_10150,N_10156);
or U10329 (N_10329,N_10051,N_10182);
or U10330 (N_10330,N_10177,N_10159);
xnor U10331 (N_10331,N_10083,N_10106);
or U10332 (N_10332,N_10147,N_10188);
xnor U10333 (N_10333,N_10102,N_10137);
or U10334 (N_10334,N_10127,N_10181);
and U10335 (N_10335,N_10131,N_10113);
nor U10336 (N_10336,N_10187,N_10184);
nand U10337 (N_10337,N_10092,N_10199);
xor U10338 (N_10338,N_10198,N_10067);
nand U10339 (N_10339,N_10153,N_10065);
nand U10340 (N_10340,N_10183,N_10077);
and U10341 (N_10341,N_10182,N_10140);
or U10342 (N_10342,N_10111,N_10149);
nand U10343 (N_10343,N_10103,N_10147);
xnor U10344 (N_10344,N_10175,N_10052);
nor U10345 (N_10345,N_10077,N_10094);
nand U10346 (N_10346,N_10128,N_10196);
nor U10347 (N_10347,N_10118,N_10054);
xnor U10348 (N_10348,N_10154,N_10125);
nand U10349 (N_10349,N_10169,N_10085);
nand U10350 (N_10350,N_10268,N_10239);
nor U10351 (N_10351,N_10275,N_10228);
nand U10352 (N_10352,N_10322,N_10257);
nand U10353 (N_10353,N_10314,N_10280);
xor U10354 (N_10354,N_10238,N_10214);
and U10355 (N_10355,N_10250,N_10285);
xor U10356 (N_10356,N_10277,N_10294);
nand U10357 (N_10357,N_10346,N_10241);
xor U10358 (N_10358,N_10324,N_10215);
or U10359 (N_10359,N_10335,N_10200);
or U10360 (N_10360,N_10244,N_10343);
and U10361 (N_10361,N_10245,N_10348);
or U10362 (N_10362,N_10295,N_10311);
or U10363 (N_10363,N_10332,N_10273);
or U10364 (N_10364,N_10223,N_10262);
nand U10365 (N_10365,N_10229,N_10253);
xor U10366 (N_10366,N_10220,N_10282);
or U10367 (N_10367,N_10234,N_10306);
xnor U10368 (N_10368,N_10303,N_10263);
or U10369 (N_10369,N_10318,N_10347);
or U10370 (N_10370,N_10261,N_10204);
nand U10371 (N_10371,N_10249,N_10259);
nor U10372 (N_10372,N_10312,N_10291);
and U10373 (N_10373,N_10248,N_10337);
nor U10374 (N_10374,N_10345,N_10320);
xnor U10375 (N_10375,N_10321,N_10325);
nand U10376 (N_10376,N_10300,N_10287);
xnor U10377 (N_10377,N_10236,N_10283);
and U10378 (N_10378,N_10286,N_10316);
nand U10379 (N_10379,N_10213,N_10319);
or U10380 (N_10380,N_10210,N_10328);
nand U10381 (N_10381,N_10330,N_10237);
or U10382 (N_10382,N_10267,N_10327);
xnor U10383 (N_10383,N_10260,N_10240);
nor U10384 (N_10384,N_10258,N_10281);
xnor U10385 (N_10385,N_10265,N_10225);
or U10386 (N_10386,N_10323,N_10329);
xnor U10387 (N_10387,N_10206,N_10218);
or U10388 (N_10388,N_10235,N_10227);
and U10389 (N_10389,N_10222,N_10270);
xor U10390 (N_10390,N_10342,N_10310);
xor U10391 (N_10391,N_10256,N_10271);
nor U10392 (N_10392,N_10207,N_10252);
nor U10393 (N_10393,N_10221,N_10301);
nand U10394 (N_10394,N_10336,N_10243);
or U10395 (N_10395,N_10224,N_10203);
nand U10396 (N_10396,N_10296,N_10212);
nor U10397 (N_10397,N_10217,N_10293);
and U10398 (N_10398,N_10209,N_10231);
nand U10399 (N_10399,N_10326,N_10278);
and U10400 (N_10400,N_10341,N_10247);
nand U10401 (N_10401,N_10233,N_10304);
or U10402 (N_10402,N_10242,N_10315);
xor U10403 (N_10403,N_10255,N_10266);
and U10404 (N_10404,N_10202,N_10289);
nor U10405 (N_10405,N_10308,N_10246);
nand U10406 (N_10406,N_10313,N_10264);
and U10407 (N_10407,N_10302,N_10299);
xor U10408 (N_10408,N_10338,N_10344);
and U10409 (N_10409,N_10333,N_10290);
and U10410 (N_10410,N_10205,N_10309);
nand U10411 (N_10411,N_10208,N_10216);
and U10412 (N_10412,N_10305,N_10272);
xor U10413 (N_10413,N_10279,N_10339);
and U10414 (N_10414,N_10232,N_10349);
nand U10415 (N_10415,N_10211,N_10331);
nand U10416 (N_10416,N_10307,N_10298);
nor U10417 (N_10417,N_10226,N_10317);
or U10418 (N_10418,N_10276,N_10230);
xor U10419 (N_10419,N_10251,N_10254);
nor U10420 (N_10420,N_10201,N_10297);
nand U10421 (N_10421,N_10334,N_10292);
nand U10422 (N_10422,N_10274,N_10284);
nor U10423 (N_10423,N_10288,N_10219);
xnor U10424 (N_10424,N_10340,N_10269);
and U10425 (N_10425,N_10238,N_10322);
nand U10426 (N_10426,N_10216,N_10342);
and U10427 (N_10427,N_10301,N_10342);
nor U10428 (N_10428,N_10223,N_10311);
xor U10429 (N_10429,N_10304,N_10321);
xor U10430 (N_10430,N_10277,N_10310);
or U10431 (N_10431,N_10226,N_10230);
nand U10432 (N_10432,N_10327,N_10237);
nor U10433 (N_10433,N_10316,N_10339);
and U10434 (N_10434,N_10252,N_10240);
nand U10435 (N_10435,N_10260,N_10330);
nand U10436 (N_10436,N_10214,N_10315);
nand U10437 (N_10437,N_10260,N_10288);
nor U10438 (N_10438,N_10326,N_10294);
and U10439 (N_10439,N_10340,N_10255);
xor U10440 (N_10440,N_10231,N_10274);
nor U10441 (N_10441,N_10225,N_10319);
xor U10442 (N_10442,N_10222,N_10300);
and U10443 (N_10443,N_10238,N_10309);
nor U10444 (N_10444,N_10288,N_10209);
xnor U10445 (N_10445,N_10340,N_10226);
nor U10446 (N_10446,N_10304,N_10329);
or U10447 (N_10447,N_10253,N_10217);
xnor U10448 (N_10448,N_10295,N_10205);
and U10449 (N_10449,N_10268,N_10232);
nand U10450 (N_10450,N_10266,N_10260);
nor U10451 (N_10451,N_10213,N_10339);
nor U10452 (N_10452,N_10317,N_10274);
nor U10453 (N_10453,N_10311,N_10342);
and U10454 (N_10454,N_10294,N_10214);
nand U10455 (N_10455,N_10242,N_10297);
nor U10456 (N_10456,N_10336,N_10220);
xor U10457 (N_10457,N_10337,N_10241);
nand U10458 (N_10458,N_10340,N_10201);
and U10459 (N_10459,N_10200,N_10305);
and U10460 (N_10460,N_10261,N_10298);
xnor U10461 (N_10461,N_10295,N_10243);
nor U10462 (N_10462,N_10225,N_10336);
xor U10463 (N_10463,N_10322,N_10229);
nor U10464 (N_10464,N_10274,N_10289);
or U10465 (N_10465,N_10300,N_10211);
xnor U10466 (N_10466,N_10323,N_10233);
nor U10467 (N_10467,N_10242,N_10244);
nand U10468 (N_10468,N_10203,N_10303);
or U10469 (N_10469,N_10295,N_10240);
nor U10470 (N_10470,N_10233,N_10246);
nor U10471 (N_10471,N_10318,N_10208);
or U10472 (N_10472,N_10304,N_10310);
nand U10473 (N_10473,N_10271,N_10200);
nand U10474 (N_10474,N_10295,N_10239);
or U10475 (N_10475,N_10320,N_10241);
or U10476 (N_10476,N_10343,N_10336);
nand U10477 (N_10477,N_10333,N_10279);
and U10478 (N_10478,N_10277,N_10286);
and U10479 (N_10479,N_10284,N_10249);
xor U10480 (N_10480,N_10231,N_10263);
nor U10481 (N_10481,N_10315,N_10206);
nand U10482 (N_10482,N_10336,N_10234);
or U10483 (N_10483,N_10258,N_10223);
or U10484 (N_10484,N_10262,N_10259);
nor U10485 (N_10485,N_10337,N_10234);
or U10486 (N_10486,N_10271,N_10238);
nor U10487 (N_10487,N_10323,N_10237);
or U10488 (N_10488,N_10201,N_10305);
nand U10489 (N_10489,N_10221,N_10283);
xnor U10490 (N_10490,N_10346,N_10221);
and U10491 (N_10491,N_10348,N_10337);
xnor U10492 (N_10492,N_10218,N_10302);
xor U10493 (N_10493,N_10225,N_10312);
or U10494 (N_10494,N_10215,N_10211);
nand U10495 (N_10495,N_10345,N_10270);
nor U10496 (N_10496,N_10269,N_10244);
nand U10497 (N_10497,N_10320,N_10224);
xnor U10498 (N_10498,N_10275,N_10278);
nand U10499 (N_10499,N_10258,N_10205);
and U10500 (N_10500,N_10410,N_10457);
nor U10501 (N_10501,N_10478,N_10374);
nand U10502 (N_10502,N_10433,N_10469);
xnor U10503 (N_10503,N_10389,N_10357);
nor U10504 (N_10504,N_10371,N_10424);
nand U10505 (N_10505,N_10475,N_10422);
nor U10506 (N_10506,N_10489,N_10460);
or U10507 (N_10507,N_10391,N_10495);
or U10508 (N_10508,N_10430,N_10380);
nor U10509 (N_10509,N_10484,N_10413);
or U10510 (N_10510,N_10477,N_10452);
and U10511 (N_10511,N_10474,N_10471);
nor U10512 (N_10512,N_10427,N_10496);
and U10513 (N_10513,N_10438,N_10385);
or U10514 (N_10514,N_10400,N_10355);
and U10515 (N_10515,N_10388,N_10499);
nor U10516 (N_10516,N_10454,N_10370);
nor U10517 (N_10517,N_10434,N_10364);
xnor U10518 (N_10518,N_10441,N_10416);
xnor U10519 (N_10519,N_10498,N_10401);
xor U10520 (N_10520,N_10456,N_10415);
nand U10521 (N_10521,N_10414,N_10491);
nor U10522 (N_10522,N_10365,N_10418);
nand U10523 (N_10523,N_10356,N_10480);
xnor U10524 (N_10524,N_10436,N_10445);
xnor U10525 (N_10525,N_10350,N_10404);
and U10526 (N_10526,N_10351,N_10394);
nor U10527 (N_10527,N_10403,N_10483);
xnor U10528 (N_10528,N_10492,N_10367);
nand U10529 (N_10529,N_10450,N_10486);
xor U10530 (N_10530,N_10381,N_10379);
nor U10531 (N_10531,N_10466,N_10488);
or U10532 (N_10532,N_10493,N_10361);
nor U10533 (N_10533,N_10359,N_10444);
nor U10534 (N_10534,N_10352,N_10412);
or U10535 (N_10535,N_10390,N_10497);
nand U10536 (N_10536,N_10353,N_10462);
nor U10537 (N_10537,N_10479,N_10428);
or U10538 (N_10538,N_10458,N_10420);
and U10539 (N_10539,N_10485,N_10396);
nand U10540 (N_10540,N_10375,N_10369);
nand U10541 (N_10541,N_10448,N_10494);
xor U10542 (N_10542,N_10395,N_10378);
nand U10543 (N_10543,N_10406,N_10425);
nor U10544 (N_10544,N_10363,N_10408);
or U10545 (N_10545,N_10443,N_10451);
xor U10546 (N_10546,N_10397,N_10482);
nand U10547 (N_10547,N_10393,N_10473);
and U10548 (N_10548,N_10437,N_10481);
nor U10549 (N_10549,N_10362,N_10377);
xor U10550 (N_10550,N_10463,N_10358);
or U10551 (N_10551,N_10382,N_10368);
or U10552 (N_10552,N_10487,N_10398);
and U10553 (N_10553,N_10384,N_10464);
xor U10554 (N_10554,N_10439,N_10372);
xnor U10555 (N_10555,N_10455,N_10373);
nand U10556 (N_10556,N_10468,N_10490);
nand U10557 (N_10557,N_10360,N_10442);
xnor U10558 (N_10558,N_10465,N_10467);
or U10559 (N_10559,N_10402,N_10446);
or U10560 (N_10560,N_10447,N_10399);
nand U10561 (N_10561,N_10407,N_10417);
xnor U10562 (N_10562,N_10431,N_10409);
and U10563 (N_10563,N_10426,N_10440);
nand U10564 (N_10564,N_10383,N_10449);
nand U10565 (N_10565,N_10432,N_10429);
or U10566 (N_10566,N_10419,N_10461);
and U10567 (N_10567,N_10411,N_10453);
nand U10568 (N_10568,N_10421,N_10354);
nand U10569 (N_10569,N_10405,N_10459);
or U10570 (N_10570,N_10387,N_10366);
nand U10571 (N_10571,N_10472,N_10470);
and U10572 (N_10572,N_10476,N_10386);
xor U10573 (N_10573,N_10376,N_10392);
nand U10574 (N_10574,N_10423,N_10435);
or U10575 (N_10575,N_10375,N_10496);
nand U10576 (N_10576,N_10451,N_10402);
or U10577 (N_10577,N_10412,N_10449);
or U10578 (N_10578,N_10398,N_10400);
xor U10579 (N_10579,N_10395,N_10363);
nor U10580 (N_10580,N_10432,N_10416);
or U10581 (N_10581,N_10427,N_10460);
xor U10582 (N_10582,N_10450,N_10439);
nand U10583 (N_10583,N_10473,N_10355);
nand U10584 (N_10584,N_10405,N_10411);
or U10585 (N_10585,N_10440,N_10439);
nor U10586 (N_10586,N_10487,N_10382);
xnor U10587 (N_10587,N_10444,N_10353);
nor U10588 (N_10588,N_10404,N_10400);
or U10589 (N_10589,N_10440,N_10467);
nor U10590 (N_10590,N_10385,N_10448);
and U10591 (N_10591,N_10434,N_10359);
nor U10592 (N_10592,N_10446,N_10371);
or U10593 (N_10593,N_10443,N_10420);
nand U10594 (N_10594,N_10429,N_10440);
or U10595 (N_10595,N_10380,N_10415);
or U10596 (N_10596,N_10427,N_10364);
nand U10597 (N_10597,N_10493,N_10407);
nand U10598 (N_10598,N_10458,N_10398);
nand U10599 (N_10599,N_10393,N_10383);
nor U10600 (N_10600,N_10452,N_10406);
and U10601 (N_10601,N_10358,N_10434);
nor U10602 (N_10602,N_10482,N_10471);
xnor U10603 (N_10603,N_10373,N_10399);
nand U10604 (N_10604,N_10442,N_10383);
xor U10605 (N_10605,N_10471,N_10441);
and U10606 (N_10606,N_10395,N_10495);
or U10607 (N_10607,N_10353,N_10455);
nand U10608 (N_10608,N_10439,N_10446);
nor U10609 (N_10609,N_10393,N_10456);
xnor U10610 (N_10610,N_10477,N_10398);
nor U10611 (N_10611,N_10403,N_10484);
and U10612 (N_10612,N_10450,N_10407);
and U10613 (N_10613,N_10472,N_10490);
or U10614 (N_10614,N_10373,N_10469);
or U10615 (N_10615,N_10362,N_10451);
and U10616 (N_10616,N_10369,N_10431);
and U10617 (N_10617,N_10443,N_10378);
and U10618 (N_10618,N_10399,N_10415);
nand U10619 (N_10619,N_10355,N_10374);
or U10620 (N_10620,N_10427,N_10386);
nor U10621 (N_10621,N_10461,N_10456);
xnor U10622 (N_10622,N_10428,N_10366);
nand U10623 (N_10623,N_10457,N_10402);
nand U10624 (N_10624,N_10369,N_10385);
nand U10625 (N_10625,N_10427,N_10365);
or U10626 (N_10626,N_10468,N_10493);
or U10627 (N_10627,N_10366,N_10417);
xor U10628 (N_10628,N_10450,N_10408);
and U10629 (N_10629,N_10499,N_10356);
nor U10630 (N_10630,N_10409,N_10378);
and U10631 (N_10631,N_10385,N_10456);
nand U10632 (N_10632,N_10401,N_10461);
and U10633 (N_10633,N_10372,N_10481);
xnor U10634 (N_10634,N_10427,N_10355);
or U10635 (N_10635,N_10358,N_10354);
or U10636 (N_10636,N_10442,N_10389);
nor U10637 (N_10637,N_10407,N_10359);
and U10638 (N_10638,N_10438,N_10410);
and U10639 (N_10639,N_10387,N_10425);
nand U10640 (N_10640,N_10410,N_10375);
or U10641 (N_10641,N_10489,N_10430);
and U10642 (N_10642,N_10400,N_10408);
nand U10643 (N_10643,N_10372,N_10476);
or U10644 (N_10644,N_10434,N_10437);
and U10645 (N_10645,N_10408,N_10425);
nand U10646 (N_10646,N_10488,N_10433);
nor U10647 (N_10647,N_10493,N_10362);
nand U10648 (N_10648,N_10453,N_10402);
xor U10649 (N_10649,N_10499,N_10395);
or U10650 (N_10650,N_10562,N_10592);
xnor U10651 (N_10651,N_10524,N_10531);
or U10652 (N_10652,N_10512,N_10510);
nand U10653 (N_10653,N_10617,N_10576);
and U10654 (N_10654,N_10616,N_10641);
xor U10655 (N_10655,N_10530,N_10571);
or U10656 (N_10656,N_10543,N_10581);
and U10657 (N_10657,N_10528,N_10522);
and U10658 (N_10658,N_10534,N_10552);
xnor U10659 (N_10659,N_10504,N_10535);
or U10660 (N_10660,N_10648,N_10575);
nor U10661 (N_10661,N_10558,N_10551);
or U10662 (N_10662,N_10642,N_10604);
or U10663 (N_10663,N_10521,N_10589);
nor U10664 (N_10664,N_10501,N_10614);
nand U10665 (N_10665,N_10538,N_10596);
nor U10666 (N_10666,N_10502,N_10585);
nand U10667 (N_10667,N_10608,N_10578);
xor U10668 (N_10668,N_10569,N_10630);
and U10669 (N_10669,N_10579,N_10621);
xor U10670 (N_10670,N_10564,N_10507);
nor U10671 (N_10671,N_10628,N_10577);
nand U10672 (N_10672,N_10505,N_10520);
nor U10673 (N_10673,N_10537,N_10540);
and U10674 (N_10674,N_10627,N_10629);
nor U10675 (N_10675,N_10563,N_10623);
and U10676 (N_10676,N_10635,N_10620);
xor U10677 (N_10677,N_10601,N_10539);
xor U10678 (N_10678,N_10503,N_10515);
nor U10679 (N_10679,N_10559,N_10605);
xnor U10680 (N_10680,N_10568,N_10548);
and U10681 (N_10681,N_10631,N_10519);
nor U10682 (N_10682,N_10595,N_10560);
and U10683 (N_10683,N_10602,N_10598);
and U10684 (N_10684,N_10517,N_10610);
xor U10685 (N_10685,N_10647,N_10638);
and U10686 (N_10686,N_10553,N_10567);
nand U10687 (N_10687,N_10636,N_10586);
and U10688 (N_10688,N_10509,N_10584);
and U10689 (N_10689,N_10500,N_10550);
nor U10690 (N_10690,N_10634,N_10541);
and U10691 (N_10691,N_10587,N_10525);
nor U10692 (N_10692,N_10542,N_10644);
xor U10693 (N_10693,N_10640,N_10612);
or U10694 (N_10694,N_10639,N_10611);
and U10695 (N_10695,N_10637,N_10583);
xor U10696 (N_10696,N_10624,N_10588);
nor U10697 (N_10697,N_10643,N_10622);
nor U10698 (N_10698,N_10600,N_10556);
xor U10699 (N_10699,N_10554,N_10603);
nor U10700 (N_10700,N_10544,N_10619);
nor U10701 (N_10701,N_10555,N_10508);
nand U10702 (N_10702,N_10590,N_10607);
and U10703 (N_10703,N_10593,N_10633);
nand U10704 (N_10704,N_10613,N_10580);
or U10705 (N_10705,N_10599,N_10632);
nand U10706 (N_10706,N_10557,N_10591);
and U10707 (N_10707,N_10526,N_10561);
xnor U10708 (N_10708,N_10511,N_10609);
or U10709 (N_10709,N_10516,N_10527);
xnor U10710 (N_10710,N_10594,N_10582);
nor U10711 (N_10711,N_10514,N_10572);
xor U10712 (N_10712,N_10549,N_10615);
nand U10713 (N_10713,N_10649,N_10570);
nand U10714 (N_10714,N_10606,N_10536);
and U10715 (N_10715,N_10529,N_10597);
nand U10716 (N_10716,N_10626,N_10625);
and U10717 (N_10717,N_10513,N_10566);
and U10718 (N_10718,N_10546,N_10523);
xor U10719 (N_10719,N_10573,N_10574);
nor U10720 (N_10720,N_10518,N_10547);
xnor U10721 (N_10721,N_10646,N_10645);
or U10722 (N_10722,N_10532,N_10545);
or U10723 (N_10723,N_10618,N_10565);
xor U10724 (N_10724,N_10533,N_10506);
xnor U10725 (N_10725,N_10574,N_10566);
or U10726 (N_10726,N_10573,N_10604);
nand U10727 (N_10727,N_10622,N_10570);
xnor U10728 (N_10728,N_10607,N_10625);
or U10729 (N_10729,N_10546,N_10579);
nor U10730 (N_10730,N_10564,N_10524);
and U10731 (N_10731,N_10607,N_10605);
or U10732 (N_10732,N_10524,N_10566);
nor U10733 (N_10733,N_10615,N_10603);
or U10734 (N_10734,N_10601,N_10577);
and U10735 (N_10735,N_10615,N_10624);
and U10736 (N_10736,N_10526,N_10538);
xor U10737 (N_10737,N_10613,N_10567);
xor U10738 (N_10738,N_10538,N_10601);
nor U10739 (N_10739,N_10581,N_10620);
or U10740 (N_10740,N_10584,N_10538);
nor U10741 (N_10741,N_10536,N_10619);
nor U10742 (N_10742,N_10562,N_10637);
nor U10743 (N_10743,N_10636,N_10513);
nor U10744 (N_10744,N_10610,N_10531);
and U10745 (N_10745,N_10619,N_10588);
and U10746 (N_10746,N_10622,N_10541);
or U10747 (N_10747,N_10582,N_10573);
or U10748 (N_10748,N_10514,N_10573);
xor U10749 (N_10749,N_10504,N_10597);
or U10750 (N_10750,N_10590,N_10576);
and U10751 (N_10751,N_10530,N_10534);
nor U10752 (N_10752,N_10564,N_10515);
xor U10753 (N_10753,N_10552,N_10575);
xnor U10754 (N_10754,N_10536,N_10639);
or U10755 (N_10755,N_10528,N_10554);
and U10756 (N_10756,N_10522,N_10569);
and U10757 (N_10757,N_10533,N_10646);
and U10758 (N_10758,N_10543,N_10523);
nor U10759 (N_10759,N_10540,N_10614);
nor U10760 (N_10760,N_10517,N_10566);
nor U10761 (N_10761,N_10599,N_10544);
nand U10762 (N_10762,N_10599,N_10524);
and U10763 (N_10763,N_10603,N_10584);
and U10764 (N_10764,N_10522,N_10558);
and U10765 (N_10765,N_10645,N_10614);
or U10766 (N_10766,N_10581,N_10523);
or U10767 (N_10767,N_10506,N_10596);
and U10768 (N_10768,N_10649,N_10621);
or U10769 (N_10769,N_10596,N_10598);
or U10770 (N_10770,N_10589,N_10586);
or U10771 (N_10771,N_10639,N_10510);
xnor U10772 (N_10772,N_10590,N_10612);
nor U10773 (N_10773,N_10567,N_10618);
and U10774 (N_10774,N_10507,N_10565);
nor U10775 (N_10775,N_10616,N_10532);
nand U10776 (N_10776,N_10549,N_10501);
nor U10777 (N_10777,N_10631,N_10523);
nor U10778 (N_10778,N_10542,N_10595);
and U10779 (N_10779,N_10535,N_10618);
or U10780 (N_10780,N_10511,N_10535);
and U10781 (N_10781,N_10614,N_10571);
nand U10782 (N_10782,N_10636,N_10570);
nor U10783 (N_10783,N_10587,N_10643);
nand U10784 (N_10784,N_10529,N_10610);
or U10785 (N_10785,N_10510,N_10506);
xnor U10786 (N_10786,N_10558,N_10588);
or U10787 (N_10787,N_10570,N_10563);
or U10788 (N_10788,N_10577,N_10512);
or U10789 (N_10789,N_10590,N_10609);
nor U10790 (N_10790,N_10581,N_10536);
nand U10791 (N_10791,N_10614,N_10589);
nand U10792 (N_10792,N_10537,N_10538);
xnor U10793 (N_10793,N_10619,N_10577);
nor U10794 (N_10794,N_10622,N_10604);
or U10795 (N_10795,N_10565,N_10581);
or U10796 (N_10796,N_10629,N_10631);
xnor U10797 (N_10797,N_10641,N_10532);
xor U10798 (N_10798,N_10608,N_10603);
and U10799 (N_10799,N_10569,N_10632);
nand U10800 (N_10800,N_10788,N_10782);
xor U10801 (N_10801,N_10726,N_10785);
nor U10802 (N_10802,N_10719,N_10706);
or U10803 (N_10803,N_10797,N_10714);
nor U10804 (N_10804,N_10681,N_10739);
nor U10805 (N_10805,N_10684,N_10723);
nand U10806 (N_10806,N_10731,N_10754);
xor U10807 (N_10807,N_10769,N_10690);
xor U10808 (N_10808,N_10734,N_10671);
xnor U10809 (N_10809,N_10677,N_10795);
nor U10810 (N_10810,N_10673,N_10652);
nor U10811 (N_10811,N_10781,N_10751);
and U10812 (N_10812,N_10697,N_10799);
nand U10813 (N_10813,N_10704,N_10787);
or U10814 (N_10814,N_10722,N_10696);
nor U10815 (N_10815,N_10727,N_10748);
and U10816 (N_10816,N_10746,N_10667);
xnor U10817 (N_10817,N_10679,N_10772);
nor U10818 (N_10818,N_10777,N_10728);
nor U10819 (N_10819,N_10662,N_10653);
nor U10820 (N_10820,N_10709,N_10670);
xnor U10821 (N_10821,N_10655,N_10718);
nor U10822 (N_10822,N_10651,N_10688);
nand U10823 (N_10823,N_10759,N_10675);
xor U10824 (N_10824,N_10692,N_10796);
nor U10825 (N_10825,N_10745,N_10778);
and U10826 (N_10826,N_10793,N_10654);
nor U10827 (N_10827,N_10701,N_10721);
xor U10828 (N_10828,N_10730,N_10678);
nand U10829 (N_10829,N_10665,N_10767);
nor U10830 (N_10830,N_10775,N_10773);
nor U10831 (N_10831,N_10694,N_10798);
or U10832 (N_10832,N_10676,N_10747);
nand U10833 (N_10833,N_10691,N_10669);
xnor U10834 (N_10834,N_10792,N_10659);
and U10835 (N_10835,N_10741,N_10715);
xnor U10836 (N_10836,N_10786,N_10699);
nor U10837 (N_10837,N_10693,N_10686);
or U10838 (N_10838,N_10749,N_10758);
xor U10839 (N_10839,N_10780,N_10784);
and U10840 (N_10840,N_10668,N_10650);
or U10841 (N_10841,N_10711,N_10702);
xor U10842 (N_10842,N_10687,N_10683);
or U10843 (N_10843,N_10695,N_10768);
and U10844 (N_10844,N_10707,N_10740);
nand U10845 (N_10845,N_10717,N_10744);
nand U10846 (N_10846,N_10752,N_10766);
nand U10847 (N_10847,N_10700,N_10674);
xnor U10848 (N_10848,N_10765,N_10771);
or U10849 (N_10849,N_10672,N_10661);
or U10850 (N_10850,N_10725,N_10762);
nand U10851 (N_10851,N_10664,N_10733);
xnor U10852 (N_10852,N_10720,N_10710);
xor U10853 (N_10853,N_10729,N_10764);
xor U10854 (N_10854,N_10724,N_10750);
or U10855 (N_10855,N_10660,N_10737);
and U10856 (N_10856,N_10713,N_10755);
nand U10857 (N_10857,N_10656,N_10680);
and U10858 (N_10858,N_10761,N_10658);
or U10859 (N_10859,N_10689,N_10703);
or U10860 (N_10860,N_10770,N_10753);
nor U10861 (N_10861,N_10682,N_10663);
xor U10862 (N_10862,N_10698,N_10666);
or U10863 (N_10863,N_10738,N_10705);
and U10864 (N_10864,N_10779,N_10790);
nand U10865 (N_10865,N_10794,N_10763);
nor U10866 (N_10866,N_10685,N_10735);
nor U10867 (N_10867,N_10743,N_10776);
xor U10868 (N_10868,N_10732,N_10791);
nor U10869 (N_10869,N_10789,N_10657);
nor U10870 (N_10870,N_10760,N_10736);
xor U10871 (N_10871,N_10712,N_10742);
and U10872 (N_10872,N_10757,N_10716);
xnor U10873 (N_10873,N_10756,N_10708);
nand U10874 (N_10874,N_10783,N_10774);
or U10875 (N_10875,N_10717,N_10686);
and U10876 (N_10876,N_10671,N_10792);
nand U10877 (N_10877,N_10787,N_10707);
xnor U10878 (N_10878,N_10669,N_10671);
nand U10879 (N_10879,N_10713,N_10785);
nand U10880 (N_10880,N_10669,N_10677);
nand U10881 (N_10881,N_10659,N_10743);
and U10882 (N_10882,N_10764,N_10704);
nor U10883 (N_10883,N_10697,N_10746);
nand U10884 (N_10884,N_10684,N_10699);
nor U10885 (N_10885,N_10667,N_10781);
nand U10886 (N_10886,N_10680,N_10788);
xnor U10887 (N_10887,N_10773,N_10744);
nor U10888 (N_10888,N_10664,N_10690);
nor U10889 (N_10889,N_10766,N_10727);
nand U10890 (N_10890,N_10662,N_10707);
nor U10891 (N_10891,N_10687,N_10758);
nor U10892 (N_10892,N_10664,N_10717);
and U10893 (N_10893,N_10690,N_10798);
and U10894 (N_10894,N_10756,N_10742);
or U10895 (N_10895,N_10704,N_10783);
and U10896 (N_10896,N_10682,N_10777);
and U10897 (N_10897,N_10661,N_10711);
nand U10898 (N_10898,N_10696,N_10770);
and U10899 (N_10899,N_10684,N_10720);
xor U10900 (N_10900,N_10741,N_10723);
nand U10901 (N_10901,N_10755,N_10674);
and U10902 (N_10902,N_10691,N_10676);
xor U10903 (N_10903,N_10748,N_10765);
and U10904 (N_10904,N_10757,N_10737);
nor U10905 (N_10905,N_10661,N_10752);
nor U10906 (N_10906,N_10714,N_10721);
or U10907 (N_10907,N_10684,N_10724);
nand U10908 (N_10908,N_10680,N_10781);
xor U10909 (N_10909,N_10667,N_10759);
or U10910 (N_10910,N_10727,N_10656);
or U10911 (N_10911,N_10770,N_10663);
and U10912 (N_10912,N_10787,N_10771);
nor U10913 (N_10913,N_10759,N_10702);
and U10914 (N_10914,N_10708,N_10762);
xnor U10915 (N_10915,N_10673,N_10747);
nand U10916 (N_10916,N_10684,N_10753);
nor U10917 (N_10917,N_10709,N_10731);
nor U10918 (N_10918,N_10695,N_10659);
nor U10919 (N_10919,N_10799,N_10795);
nor U10920 (N_10920,N_10653,N_10709);
nor U10921 (N_10921,N_10730,N_10702);
and U10922 (N_10922,N_10774,N_10710);
and U10923 (N_10923,N_10672,N_10740);
nor U10924 (N_10924,N_10798,N_10779);
xnor U10925 (N_10925,N_10775,N_10743);
or U10926 (N_10926,N_10777,N_10672);
or U10927 (N_10927,N_10711,N_10750);
or U10928 (N_10928,N_10757,N_10678);
or U10929 (N_10929,N_10693,N_10714);
xnor U10930 (N_10930,N_10749,N_10792);
and U10931 (N_10931,N_10667,N_10670);
nand U10932 (N_10932,N_10774,N_10677);
nor U10933 (N_10933,N_10662,N_10766);
nor U10934 (N_10934,N_10720,N_10688);
and U10935 (N_10935,N_10653,N_10727);
or U10936 (N_10936,N_10750,N_10656);
xor U10937 (N_10937,N_10757,N_10706);
xor U10938 (N_10938,N_10781,N_10653);
nand U10939 (N_10939,N_10752,N_10723);
nor U10940 (N_10940,N_10674,N_10753);
nor U10941 (N_10941,N_10670,N_10671);
nand U10942 (N_10942,N_10730,N_10733);
nor U10943 (N_10943,N_10688,N_10725);
nor U10944 (N_10944,N_10662,N_10747);
nor U10945 (N_10945,N_10687,N_10689);
or U10946 (N_10946,N_10690,N_10670);
nand U10947 (N_10947,N_10733,N_10739);
nor U10948 (N_10948,N_10700,N_10696);
xor U10949 (N_10949,N_10789,N_10723);
or U10950 (N_10950,N_10812,N_10873);
xor U10951 (N_10951,N_10814,N_10853);
or U10952 (N_10952,N_10922,N_10809);
nor U10953 (N_10953,N_10858,N_10813);
or U10954 (N_10954,N_10846,N_10928);
or U10955 (N_10955,N_10883,N_10816);
and U10956 (N_10956,N_10937,N_10841);
or U10957 (N_10957,N_10878,N_10810);
and U10958 (N_10958,N_10882,N_10819);
xor U10959 (N_10959,N_10909,N_10925);
or U10960 (N_10960,N_10916,N_10921);
and U10961 (N_10961,N_10894,N_10806);
nand U10962 (N_10962,N_10835,N_10838);
xor U10963 (N_10963,N_10875,N_10861);
or U10964 (N_10964,N_10919,N_10911);
or U10965 (N_10965,N_10817,N_10939);
xor U10966 (N_10966,N_10926,N_10895);
or U10967 (N_10967,N_10856,N_10826);
nand U10968 (N_10968,N_10855,N_10889);
and U10969 (N_10969,N_10900,N_10907);
and U10970 (N_10970,N_10868,N_10822);
nor U10971 (N_10971,N_10910,N_10897);
nand U10972 (N_10972,N_10876,N_10941);
nor U10973 (N_10973,N_10857,N_10888);
and U10974 (N_10974,N_10940,N_10832);
nand U10975 (N_10975,N_10818,N_10831);
nor U10976 (N_10976,N_10871,N_10912);
xnor U10977 (N_10977,N_10845,N_10935);
or U10978 (N_10978,N_10839,N_10947);
nand U10979 (N_10979,N_10801,N_10945);
nand U10980 (N_10980,N_10828,N_10825);
nand U10981 (N_10981,N_10887,N_10823);
xnor U10982 (N_10982,N_10820,N_10864);
or U10983 (N_10983,N_10836,N_10896);
nor U10984 (N_10984,N_10901,N_10829);
nand U10985 (N_10985,N_10803,N_10874);
or U10986 (N_10986,N_10872,N_10918);
and U10987 (N_10987,N_10860,N_10890);
nor U10988 (N_10988,N_10924,N_10892);
nor U10989 (N_10989,N_10811,N_10824);
or U10990 (N_10990,N_10904,N_10930);
xor U10991 (N_10991,N_10908,N_10844);
xnor U10992 (N_10992,N_10893,N_10923);
nor U10993 (N_10993,N_10833,N_10946);
xnor U10994 (N_10994,N_10936,N_10842);
nor U10995 (N_10995,N_10932,N_10867);
and U10996 (N_10996,N_10942,N_10931);
and U10997 (N_10997,N_10902,N_10886);
or U10998 (N_10998,N_10881,N_10847);
or U10999 (N_10999,N_10849,N_10929);
and U11000 (N_11000,N_10879,N_10915);
nor U11001 (N_11001,N_10884,N_10821);
nand U11002 (N_11002,N_10903,N_10899);
nor U11003 (N_11003,N_10808,N_10948);
xor U11004 (N_11004,N_10834,N_10891);
xor U11005 (N_11005,N_10859,N_10848);
and U11006 (N_11006,N_10898,N_10913);
nand U11007 (N_11007,N_10800,N_10862);
nor U11008 (N_11008,N_10854,N_10933);
or U11009 (N_11009,N_10949,N_10850);
and U11010 (N_11010,N_10837,N_10804);
nor U11011 (N_11011,N_10863,N_10843);
xnor U11012 (N_11012,N_10830,N_10805);
nor U11013 (N_11013,N_10827,N_10866);
or U11014 (N_11014,N_10840,N_10905);
and U11015 (N_11015,N_10944,N_10920);
and U11016 (N_11016,N_10943,N_10927);
nor U11017 (N_11017,N_10938,N_10877);
or U11018 (N_11018,N_10807,N_10914);
or U11019 (N_11019,N_10802,N_10880);
or U11020 (N_11020,N_10852,N_10870);
and U11021 (N_11021,N_10934,N_10851);
nand U11022 (N_11022,N_10917,N_10869);
or U11023 (N_11023,N_10815,N_10906);
nand U11024 (N_11024,N_10865,N_10885);
xor U11025 (N_11025,N_10827,N_10863);
nand U11026 (N_11026,N_10933,N_10863);
nor U11027 (N_11027,N_10919,N_10868);
nor U11028 (N_11028,N_10917,N_10897);
or U11029 (N_11029,N_10801,N_10891);
xor U11030 (N_11030,N_10861,N_10923);
and U11031 (N_11031,N_10861,N_10805);
and U11032 (N_11032,N_10813,N_10888);
or U11033 (N_11033,N_10846,N_10911);
nand U11034 (N_11034,N_10949,N_10840);
and U11035 (N_11035,N_10808,N_10824);
nor U11036 (N_11036,N_10907,N_10883);
xnor U11037 (N_11037,N_10887,N_10911);
and U11038 (N_11038,N_10849,N_10894);
or U11039 (N_11039,N_10838,N_10919);
and U11040 (N_11040,N_10804,N_10840);
nor U11041 (N_11041,N_10823,N_10902);
nand U11042 (N_11042,N_10830,N_10856);
nand U11043 (N_11043,N_10927,N_10886);
nand U11044 (N_11044,N_10818,N_10907);
nand U11045 (N_11045,N_10801,N_10835);
xnor U11046 (N_11046,N_10871,N_10850);
xor U11047 (N_11047,N_10914,N_10916);
xor U11048 (N_11048,N_10946,N_10939);
nand U11049 (N_11049,N_10877,N_10835);
xor U11050 (N_11050,N_10887,N_10855);
or U11051 (N_11051,N_10911,N_10855);
nor U11052 (N_11052,N_10842,N_10929);
nor U11053 (N_11053,N_10821,N_10831);
or U11054 (N_11054,N_10942,N_10800);
and U11055 (N_11055,N_10862,N_10893);
xnor U11056 (N_11056,N_10920,N_10872);
and U11057 (N_11057,N_10804,N_10943);
or U11058 (N_11058,N_10940,N_10886);
or U11059 (N_11059,N_10888,N_10918);
or U11060 (N_11060,N_10880,N_10817);
xnor U11061 (N_11061,N_10901,N_10858);
or U11062 (N_11062,N_10894,N_10933);
and U11063 (N_11063,N_10812,N_10813);
or U11064 (N_11064,N_10935,N_10907);
xor U11065 (N_11065,N_10833,N_10871);
nand U11066 (N_11066,N_10886,N_10900);
xnor U11067 (N_11067,N_10941,N_10868);
nor U11068 (N_11068,N_10867,N_10849);
nand U11069 (N_11069,N_10843,N_10816);
nand U11070 (N_11070,N_10876,N_10940);
and U11071 (N_11071,N_10939,N_10839);
nor U11072 (N_11072,N_10844,N_10925);
or U11073 (N_11073,N_10827,N_10819);
and U11074 (N_11074,N_10897,N_10847);
nand U11075 (N_11075,N_10923,N_10858);
nor U11076 (N_11076,N_10809,N_10948);
and U11077 (N_11077,N_10904,N_10880);
or U11078 (N_11078,N_10917,N_10880);
and U11079 (N_11079,N_10910,N_10874);
nand U11080 (N_11080,N_10942,N_10892);
xnor U11081 (N_11081,N_10854,N_10930);
or U11082 (N_11082,N_10896,N_10898);
nor U11083 (N_11083,N_10905,N_10909);
nor U11084 (N_11084,N_10897,N_10836);
xnor U11085 (N_11085,N_10802,N_10940);
and U11086 (N_11086,N_10946,N_10885);
or U11087 (N_11087,N_10900,N_10821);
xnor U11088 (N_11088,N_10854,N_10828);
nand U11089 (N_11089,N_10918,N_10805);
and U11090 (N_11090,N_10838,N_10908);
or U11091 (N_11091,N_10805,N_10934);
and U11092 (N_11092,N_10843,N_10947);
and U11093 (N_11093,N_10868,N_10818);
nand U11094 (N_11094,N_10803,N_10860);
or U11095 (N_11095,N_10834,N_10860);
nor U11096 (N_11096,N_10829,N_10915);
and U11097 (N_11097,N_10828,N_10860);
and U11098 (N_11098,N_10849,N_10930);
xnor U11099 (N_11099,N_10800,N_10910);
or U11100 (N_11100,N_11008,N_10980);
or U11101 (N_11101,N_11017,N_10983);
nand U11102 (N_11102,N_10981,N_11095);
or U11103 (N_11103,N_10955,N_11078);
nand U11104 (N_11104,N_11092,N_10970);
and U11105 (N_11105,N_11079,N_11099);
xor U11106 (N_11106,N_10951,N_11048);
nor U11107 (N_11107,N_11031,N_10958);
and U11108 (N_11108,N_11065,N_11086);
xor U11109 (N_11109,N_11050,N_10986);
xnor U11110 (N_11110,N_11093,N_10995);
xor U11111 (N_11111,N_11064,N_11037);
and U11112 (N_11112,N_11038,N_10984);
nor U11113 (N_11113,N_10996,N_11066);
nor U11114 (N_11114,N_11090,N_11007);
xnor U11115 (N_11115,N_11083,N_10953);
nand U11116 (N_11116,N_11002,N_10999);
nor U11117 (N_11117,N_11094,N_10972);
xnor U11118 (N_11118,N_11000,N_11057);
or U11119 (N_11119,N_11039,N_11036);
nor U11120 (N_11120,N_11005,N_11076);
xor U11121 (N_11121,N_11033,N_11070);
or U11122 (N_11122,N_11084,N_11015);
or U11123 (N_11123,N_11098,N_11096);
or U11124 (N_11124,N_11047,N_11034);
nor U11125 (N_11125,N_11089,N_11013);
or U11126 (N_11126,N_10962,N_11012);
nand U11127 (N_11127,N_11055,N_10964);
or U11128 (N_11128,N_11091,N_11026);
nor U11129 (N_11129,N_11056,N_10991);
xor U11130 (N_11130,N_10998,N_11080);
nor U11131 (N_11131,N_11063,N_11069);
nand U11132 (N_11132,N_10974,N_10976);
and U11133 (N_11133,N_11027,N_10989);
xor U11134 (N_11134,N_11004,N_11029);
and U11135 (N_11135,N_10982,N_11028);
or U11136 (N_11136,N_11088,N_10971);
or U11137 (N_11137,N_10977,N_10963);
and U11138 (N_11138,N_11082,N_11087);
nand U11139 (N_11139,N_10969,N_11071);
or U11140 (N_11140,N_10952,N_11073);
nand U11141 (N_11141,N_10990,N_11022);
nand U11142 (N_11142,N_11009,N_10975);
or U11143 (N_11143,N_11045,N_11040);
and U11144 (N_11144,N_11051,N_10957);
and U11145 (N_11145,N_11003,N_11041);
or U11146 (N_11146,N_11016,N_11077);
nor U11147 (N_11147,N_10979,N_11081);
and U11148 (N_11148,N_11074,N_10960);
nor U11149 (N_11149,N_11030,N_10954);
nand U11150 (N_11150,N_11018,N_11001);
nor U11151 (N_11151,N_11023,N_11006);
xnor U11152 (N_11152,N_10950,N_11019);
nand U11153 (N_11153,N_11072,N_10956);
nand U11154 (N_11154,N_11059,N_11058);
xor U11155 (N_11155,N_11046,N_11085);
or U11156 (N_11156,N_11052,N_11067);
nor U11157 (N_11157,N_10997,N_10961);
nand U11158 (N_11158,N_11032,N_11062);
nor U11159 (N_11159,N_11014,N_10987);
nand U11160 (N_11160,N_10966,N_10978);
and U11161 (N_11161,N_11025,N_10967);
nor U11162 (N_11162,N_10959,N_11061);
or U11163 (N_11163,N_11049,N_11020);
nand U11164 (N_11164,N_11042,N_10985);
xor U11165 (N_11165,N_11075,N_11035);
and U11166 (N_11166,N_10992,N_11097);
xor U11167 (N_11167,N_11011,N_10994);
nand U11168 (N_11168,N_10988,N_11024);
and U11169 (N_11169,N_11043,N_11044);
and U11170 (N_11170,N_10973,N_11068);
or U11171 (N_11171,N_10968,N_11053);
nand U11172 (N_11172,N_10965,N_11060);
xor U11173 (N_11173,N_11054,N_10993);
and U11174 (N_11174,N_11010,N_11021);
nand U11175 (N_11175,N_11001,N_10973);
nand U11176 (N_11176,N_11050,N_10958);
or U11177 (N_11177,N_11067,N_10966);
nand U11178 (N_11178,N_11012,N_10985);
nor U11179 (N_11179,N_11021,N_11040);
or U11180 (N_11180,N_11095,N_10957);
xor U11181 (N_11181,N_11078,N_11058);
or U11182 (N_11182,N_11014,N_11005);
nor U11183 (N_11183,N_10984,N_11097);
nand U11184 (N_11184,N_10989,N_11041);
nor U11185 (N_11185,N_11084,N_11016);
nand U11186 (N_11186,N_11042,N_10963);
and U11187 (N_11187,N_10954,N_10995);
nor U11188 (N_11188,N_10999,N_11058);
nand U11189 (N_11189,N_11071,N_11027);
nand U11190 (N_11190,N_11007,N_10985);
nand U11191 (N_11191,N_10987,N_11022);
nor U11192 (N_11192,N_11082,N_10987);
xor U11193 (N_11193,N_11091,N_10983);
and U11194 (N_11194,N_10970,N_11010);
nand U11195 (N_11195,N_11012,N_11090);
nand U11196 (N_11196,N_11024,N_10963);
and U11197 (N_11197,N_11066,N_11021);
nand U11198 (N_11198,N_10981,N_11016);
nand U11199 (N_11199,N_11001,N_10961);
nand U11200 (N_11200,N_10962,N_11021);
or U11201 (N_11201,N_11076,N_11058);
xor U11202 (N_11202,N_10988,N_11034);
and U11203 (N_11203,N_11045,N_10977);
and U11204 (N_11204,N_10999,N_10985);
xnor U11205 (N_11205,N_10998,N_10970);
nand U11206 (N_11206,N_11019,N_11013);
xnor U11207 (N_11207,N_11017,N_10985);
xnor U11208 (N_11208,N_11012,N_11074);
nand U11209 (N_11209,N_11011,N_11054);
and U11210 (N_11210,N_10965,N_10979);
xnor U11211 (N_11211,N_11084,N_10996);
nor U11212 (N_11212,N_10992,N_11055);
and U11213 (N_11213,N_11090,N_10991);
and U11214 (N_11214,N_11070,N_11017);
or U11215 (N_11215,N_11092,N_10977);
and U11216 (N_11216,N_11076,N_11002);
nor U11217 (N_11217,N_11071,N_10981);
and U11218 (N_11218,N_11051,N_11017);
or U11219 (N_11219,N_11066,N_11070);
and U11220 (N_11220,N_11025,N_10961);
xor U11221 (N_11221,N_11099,N_10986);
nand U11222 (N_11222,N_11004,N_11096);
and U11223 (N_11223,N_10992,N_10955);
and U11224 (N_11224,N_11055,N_10977);
nor U11225 (N_11225,N_10974,N_10953);
or U11226 (N_11226,N_11096,N_11068);
xnor U11227 (N_11227,N_10959,N_11024);
and U11228 (N_11228,N_11051,N_11035);
xor U11229 (N_11229,N_10958,N_11090);
xor U11230 (N_11230,N_11082,N_11034);
or U11231 (N_11231,N_10976,N_10993);
and U11232 (N_11232,N_11057,N_11046);
xnor U11233 (N_11233,N_11066,N_10984);
xor U11234 (N_11234,N_10972,N_10987);
or U11235 (N_11235,N_10966,N_10972);
nand U11236 (N_11236,N_11025,N_10971);
nor U11237 (N_11237,N_11078,N_10991);
xnor U11238 (N_11238,N_11004,N_11032);
nand U11239 (N_11239,N_11084,N_11048);
or U11240 (N_11240,N_11065,N_10952);
or U11241 (N_11241,N_11023,N_11085);
and U11242 (N_11242,N_10965,N_10988);
xnor U11243 (N_11243,N_11005,N_10980);
xor U11244 (N_11244,N_11060,N_11075);
nor U11245 (N_11245,N_11030,N_11093);
xnor U11246 (N_11246,N_10962,N_11053);
and U11247 (N_11247,N_10954,N_11049);
or U11248 (N_11248,N_11017,N_11068);
and U11249 (N_11249,N_11019,N_11029);
nand U11250 (N_11250,N_11184,N_11205);
nand U11251 (N_11251,N_11164,N_11115);
nor U11252 (N_11252,N_11178,N_11224);
xnor U11253 (N_11253,N_11128,N_11218);
and U11254 (N_11254,N_11185,N_11211);
nand U11255 (N_11255,N_11221,N_11122);
nor U11256 (N_11256,N_11134,N_11138);
and U11257 (N_11257,N_11137,N_11192);
nor U11258 (N_11258,N_11239,N_11194);
nand U11259 (N_11259,N_11208,N_11103);
nor U11260 (N_11260,N_11153,N_11156);
and U11261 (N_11261,N_11206,N_11231);
xor U11262 (N_11262,N_11140,N_11180);
or U11263 (N_11263,N_11223,N_11233);
xor U11264 (N_11264,N_11100,N_11112);
nor U11265 (N_11265,N_11190,N_11227);
xnor U11266 (N_11266,N_11222,N_11121);
xor U11267 (N_11267,N_11157,N_11209);
nand U11268 (N_11268,N_11161,N_11191);
nor U11269 (N_11269,N_11104,N_11226);
and U11270 (N_11270,N_11126,N_11127);
nor U11271 (N_11271,N_11173,N_11110);
nand U11272 (N_11272,N_11242,N_11154);
and U11273 (N_11273,N_11160,N_11247);
xnor U11274 (N_11274,N_11167,N_11169);
xnor U11275 (N_11275,N_11136,N_11113);
nor U11276 (N_11276,N_11129,N_11123);
nand U11277 (N_11277,N_11159,N_11105);
nor U11278 (N_11278,N_11111,N_11106);
xor U11279 (N_11279,N_11132,N_11204);
or U11280 (N_11280,N_11149,N_11193);
or U11281 (N_11281,N_11116,N_11172);
nand U11282 (N_11282,N_11246,N_11143);
nand U11283 (N_11283,N_11133,N_11142);
xor U11284 (N_11284,N_11183,N_11232);
or U11285 (N_11285,N_11155,N_11171);
nor U11286 (N_11286,N_11238,N_11158);
xor U11287 (N_11287,N_11118,N_11109);
nand U11288 (N_11288,N_11125,N_11139);
and U11289 (N_11289,N_11197,N_11230);
and U11290 (N_11290,N_11186,N_11243);
or U11291 (N_11291,N_11141,N_11174);
nor U11292 (N_11292,N_11188,N_11235);
and U11293 (N_11293,N_11214,N_11176);
nand U11294 (N_11294,N_11225,N_11145);
nand U11295 (N_11295,N_11151,N_11236);
nor U11296 (N_11296,N_11212,N_11229);
xor U11297 (N_11297,N_11177,N_11166);
or U11298 (N_11298,N_11234,N_11107);
or U11299 (N_11299,N_11102,N_11150);
or U11300 (N_11300,N_11203,N_11195);
xor U11301 (N_11301,N_11120,N_11200);
nand U11302 (N_11302,N_11130,N_11170);
nand U11303 (N_11303,N_11119,N_11148);
nor U11304 (N_11304,N_11237,N_11135);
xnor U11305 (N_11305,N_11245,N_11131);
xnor U11306 (N_11306,N_11201,N_11249);
xor U11307 (N_11307,N_11114,N_11202);
or U11308 (N_11308,N_11241,N_11163);
nor U11309 (N_11309,N_11179,N_11228);
nand U11310 (N_11310,N_11210,N_11187);
nand U11311 (N_11311,N_11216,N_11144);
xor U11312 (N_11312,N_11199,N_11219);
and U11313 (N_11313,N_11215,N_11101);
and U11314 (N_11314,N_11146,N_11244);
and U11315 (N_11315,N_11124,N_11207);
nand U11316 (N_11316,N_11162,N_11168);
or U11317 (N_11317,N_11248,N_11182);
xor U11318 (N_11318,N_11165,N_11152);
and U11319 (N_11319,N_11117,N_11175);
nand U11320 (N_11320,N_11181,N_11189);
and U11321 (N_11321,N_11217,N_11147);
or U11322 (N_11322,N_11196,N_11240);
nor U11323 (N_11323,N_11198,N_11213);
and U11324 (N_11324,N_11108,N_11220);
or U11325 (N_11325,N_11211,N_11108);
xor U11326 (N_11326,N_11107,N_11157);
nand U11327 (N_11327,N_11235,N_11122);
nand U11328 (N_11328,N_11191,N_11130);
and U11329 (N_11329,N_11119,N_11226);
or U11330 (N_11330,N_11148,N_11205);
nor U11331 (N_11331,N_11190,N_11216);
nand U11332 (N_11332,N_11196,N_11204);
nor U11333 (N_11333,N_11202,N_11132);
or U11334 (N_11334,N_11152,N_11217);
xnor U11335 (N_11335,N_11103,N_11188);
nand U11336 (N_11336,N_11240,N_11126);
or U11337 (N_11337,N_11120,N_11215);
or U11338 (N_11338,N_11116,N_11139);
nand U11339 (N_11339,N_11123,N_11109);
or U11340 (N_11340,N_11114,N_11184);
or U11341 (N_11341,N_11157,N_11184);
nor U11342 (N_11342,N_11139,N_11195);
or U11343 (N_11343,N_11204,N_11160);
nor U11344 (N_11344,N_11215,N_11168);
xnor U11345 (N_11345,N_11127,N_11141);
xor U11346 (N_11346,N_11160,N_11249);
xor U11347 (N_11347,N_11228,N_11192);
or U11348 (N_11348,N_11131,N_11203);
nand U11349 (N_11349,N_11232,N_11143);
or U11350 (N_11350,N_11155,N_11128);
xnor U11351 (N_11351,N_11178,N_11200);
or U11352 (N_11352,N_11205,N_11223);
nand U11353 (N_11353,N_11203,N_11128);
xnor U11354 (N_11354,N_11193,N_11151);
nand U11355 (N_11355,N_11177,N_11109);
nor U11356 (N_11356,N_11127,N_11164);
xnor U11357 (N_11357,N_11183,N_11151);
xor U11358 (N_11358,N_11109,N_11234);
or U11359 (N_11359,N_11146,N_11172);
xnor U11360 (N_11360,N_11126,N_11244);
nand U11361 (N_11361,N_11207,N_11154);
nor U11362 (N_11362,N_11193,N_11186);
or U11363 (N_11363,N_11120,N_11165);
xnor U11364 (N_11364,N_11141,N_11180);
xnor U11365 (N_11365,N_11246,N_11131);
nand U11366 (N_11366,N_11198,N_11117);
nand U11367 (N_11367,N_11169,N_11194);
nor U11368 (N_11368,N_11102,N_11179);
xor U11369 (N_11369,N_11245,N_11170);
nand U11370 (N_11370,N_11141,N_11246);
and U11371 (N_11371,N_11110,N_11185);
or U11372 (N_11372,N_11135,N_11165);
nand U11373 (N_11373,N_11241,N_11154);
nor U11374 (N_11374,N_11192,N_11102);
and U11375 (N_11375,N_11215,N_11103);
or U11376 (N_11376,N_11201,N_11238);
nor U11377 (N_11377,N_11144,N_11224);
or U11378 (N_11378,N_11172,N_11225);
nor U11379 (N_11379,N_11110,N_11171);
xnor U11380 (N_11380,N_11232,N_11170);
xnor U11381 (N_11381,N_11187,N_11149);
and U11382 (N_11382,N_11232,N_11198);
xor U11383 (N_11383,N_11107,N_11207);
nand U11384 (N_11384,N_11238,N_11189);
nor U11385 (N_11385,N_11184,N_11247);
xnor U11386 (N_11386,N_11126,N_11202);
nand U11387 (N_11387,N_11142,N_11171);
nand U11388 (N_11388,N_11190,N_11122);
nor U11389 (N_11389,N_11190,N_11185);
nor U11390 (N_11390,N_11135,N_11126);
xnor U11391 (N_11391,N_11197,N_11121);
nor U11392 (N_11392,N_11193,N_11117);
nand U11393 (N_11393,N_11193,N_11158);
xor U11394 (N_11394,N_11159,N_11114);
or U11395 (N_11395,N_11173,N_11175);
nor U11396 (N_11396,N_11159,N_11153);
nand U11397 (N_11397,N_11101,N_11198);
nand U11398 (N_11398,N_11155,N_11185);
or U11399 (N_11399,N_11109,N_11199);
nor U11400 (N_11400,N_11274,N_11321);
nor U11401 (N_11401,N_11341,N_11368);
nor U11402 (N_11402,N_11392,N_11384);
or U11403 (N_11403,N_11332,N_11294);
nand U11404 (N_11404,N_11299,N_11293);
nor U11405 (N_11405,N_11334,N_11287);
nor U11406 (N_11406,N_11371,N_11336);
nand U11407 (N_11407,N_11300,N_11338);
or U11408 (N_11408,N_11390,N_11272);
nand U11409 (N_11409,N_11314,N_11342);
nor U11410 (N_11410,N_11258,N_11256);
nand U11411 (N_11411,N_11333,N_11298);
or U11412 (N_11412,N_11335,N_11350);
nor U11413 (N_11413,N_11264,N_11296);
or U11414 (N_11414,N_11365,N_11345);
nor U11415 (N_11415,N_11376,N_11303);
nor U11416 (N_11416,N_11363,N_11399);
nand U11417 (N_11417,N_11250,N_11267);
nand U11418 (N_11418,N_11395,N_11396);
and U11419 (N_11419,N_11362,N_11385);
xor U11420 (N_11420,N_11337,N_11319);
and U11421 (N_11421,N_11369,N_11254);
or U11422 (N_11422,N_11343,N_11347);
nand U11423 (N_11423,N_11277,N_11356);
nand U11424 (N_11424,N_11367,N_11340);
nor U11425 (N_11425,N_11318,N_11391);
and U11426 (N_11426,N_11304,N_11358);
nand U11427 (N_11427,N_11360,N_11324);
nor U11428 (N_11428,N_11279,N_11278);
or U11429 (N_11429,N_11305,N_11315);
and U11430 (N_11430,N_11292,N_11285);
nand U11431 (N_11431,N_11309,N_11325);
xnor U11432 (N_11432,N_11301,N_11364);
and U11433 (N_11433,N_11381,N_11323);
or U11434 (N_11434,N_11374,N_11355);
nor U11435 (N_11435,N_11313,N_11387);
or U11436 (N_11436,N_11377,N_11255);
or U11437 (N_11437,N_11295,N_11394);
xnor U11438 (N_11438,N_11386,N_11382);
or U11439 (N_11439,N_11339,N_11306);
and U11440 (N_11440,N_11253,N_11393);
and U11441 (N_11441,N_11378,N_11346);
xnor U11442 (N_11442,N_11327,N_11366);
nand U11443 (N_11443,N_11262,N_11265);
nor U11444 (N_11444,N_11260,N_11283);
or U11445 (N_11445,N_11273,N_11308);
nor U11446 (N_11446,N_11257,N_11251);
xor U11447 (N_11447,N_11344,N_11316);
or U11448 (N_11448,N_11348,N_11261);
nand U11449 (N_11449,N_11259,N_11388);
nand U11450 (N_11450,N_11320,N_11361);
and U11451 (N_11451,N_11397,N_11290);
nand U11452 (N_11452,N_11379,N_11311);
and U11453 (N_11453,N_11322,N_11282);
xor U11454 (N_11454,N_11326,N_11329);
or U11455 (N_11455,N_11281,N_11349);
nand U11456 (N_11456,N_11352,N_11271);
nand U11457 (N_11457,N_11270,N_11289);
or U11458 (N_11458,N_11312,N_11330);
and U11459 (N_11459,N_11380,N_11269);
and U11460 (N_11460,N_11307,N_11353);
and U11461 (N_11461,N_11328,N_11372);
xor U11462 (N_11462,N_11302,N_11383);
xor U11463 (N_11463,N_11354,N_11389);
or U11464 (N_11464,N_11359,N_11331);
nor U11465 (N_11465,N_11373,N_11284);
nand U11466 (N_11466,N_11375,N_11275);
xnor U11467 (N_11467,N_11297,N_11263);
xnor U11468 (N_11468,N_11266,N_11398);
nor U11469 (N_11469,N_11276,N_11280);
or U11470 (N_11470,N_11252,N_11310);
and U11471 (N_11471,N_11286,N_11291);
and U11472 (N_11472,N_11357,N_11351);
or U11473 (N_11473,N_11317,N_11288);
nor U11474 (N_11474,N_11268,N_11370);
nand U11475 (N_11475,N_11349,N_11390);
xor U11476 (N_11476,N_11284,N_11304);
or U11477 (N_11477,N_11345,N_11261);
xor U11478 (N_11478,N_11313,N_11341);
nor U11479 (N_11479,N_11285,N_11311);
and U11480 (N_11480,N_11336,N_11385);
nor U11481 (N_11481,N_11258,N_11307);
and U11482 (N_11482,N_11279,N_11363);
xnor U11483 (N_11483,N_11274,N_11303);
nand U11484 (N_11484,N_11337,N_11321);
and U11485 (N_11485,N_11349,N_11361);
and U11486 (N_11486,N_11304,N_11300);
nor U11487 (N_11487,N_11301,N_11381);
nand U11488 (N_11488,N_11339,N_11266);
and U11489 (N_11489,N_11330,N_11393);
or U11490 (N_11490,N_11258,N_11344);
and U11491 (N_11491,N_11354,N_11359);
nand U11492 (N_11492,N_11341,N_11289);
and U11493 (N_11493,N_11362,N_11272);
nand U11494 (N_11494,N_11280,N_11326);
nor U11495 (N_11495,N_11341,N_11252);
xor U11496 (N_11496,N_11334,N_11293);
nand U11497 (N_11497,N_11324,N_11293);
nand U11498 (N_11498,N_11299,N_11345);
nand U11499 (N_11499,N_11398,N_11260);
xnor U11500 (N_11500,N_11265,N_11274);
and U11501 (N_11501,N_11337,N_11379);
xnor U11502 (N_11502,N_11272,N_11254);
nand U11503 (N_11503,N_11276,N_11395);
xor U11504 (N_11504,N_11266,N_11285);
xor U11505 (N_11505,N_11351,N_11268);
nor U11506 (N_11506,N_11284,N_11288);
and U11507 (N_11507,N_11383,N_11387);
or U11508 (N_11508,N_11371,N_11350);
nor U11509 (N_11509,N_11280,N_11263);
nand U11510 (N_11510,N_11334,N_11273);
xnor U11511 (N_11511,N_11298,N_11284);
nand U11512 (N_11512,N_11287,N_11302);
nor U11513 (N_11513,N_11322,N_11355);
xnor U11514 (N_11514,N_11373,N_11341);
or U11515 (N_11515,N_11302,N_11367);
xnor U11516 (N_11516,N_11379,N_11302);
nor U11517 (N_11517,N_11369,N_11376);
xnor U11518 (N_11518,N_11257,N_11379);
xnor U11519 (N_11519,N_11340,N_11318);
nor U11520 (N_11520,N_11272,N_11377);
nor U11521 (N_11521,N_11394,N_11323);
or U11522 (N_11522,N_11288,N_11289);
xnor U11523 (N_11523,N_11266,N_11384);
or U11524 (N_11524,N_11362,N_11315);
xor U11525 (N_11525,N_11364,N_11259);
or U11526 (N_11526,N_11389,N_11367);
nor U11527 (N_11527,N_11250,N_11354);
nand U11528 (N_11528,N_11378,N_11259);
nor U11529 (N_11529,N_11345,N_11366);
xnor U11530 (N_11530,N_11271,N_11378);
nor U11531 (N_11531,N_11251,N_11342);
nand U11532 (N_11532,N_11259,N_11275);
nor U11533 (N_11533,N_11261,N_11385);
nand U11534 (N_11534,N_11317,N_11303);
xnor U11535 (N_11535,N_11361,N_11287);
and U11536 (N_11536,N_11346,N_11343);
nor U11537 (N_11537,N_11319,N_11307);
xnor U11538 (N_11538,N_11344,N_11353);
nor U11539 (N_11539,N_11295,N_11250);
or U11540 (N_11540,N_11288,N_11279);
xor U11541 (N_11541,N_11255,N_11300);
xor U11542 (N_11542,N_11389,N_11295);
nor U11543 (N_11543,N_11313,N_11311);
xor U11544 (N_11544,N_11283,N_11288);
nand U11545 (N_11545,N_11296,N_11390);
xor U11546 (N_11546,N_11313,N_11296);
xnor U11547 (N_11547,N_11372,N_11363);
or U11548 (N_11548,N_11371,N_11344);
xnor U11549 (N_11549,N_11362,N_11254);
nand U11550 (N_11550,N_11449,N_11539);
xnor U11551 (N_11551,N_11455,N_11542);
and U11552 (N_11552,N_11425,N_11530);
or U11553 (N_11553,N_11412,N_11423);
nand U11554 (N_11554,N_11446,N_11524);
and U11555 (N_11555,N_11513,N_11491);
xnor U11556 (N_11556,N_11473,N_11430);
or U11557 (N_11557,N_11439,N_11436);
xor U11558 (N_11558,N_11408,N_11471);
xnor U11559 (N_11559,N_11548,N_11431);
xor U11560 (N_11560,N_11472,N_11438);
nand U11561 (N_11561,N_11515,N_11478);
xnor U11562 (N_11562,N_11461,N_11497);
nor U11563 (N_11563,N_11443,N_11484);
or U11564 (N_11564,N_11428,N_11459);
and U11565 (N_11565,N_11482,N_11535);
or U11566 (N_11566,N_11502,N_11448);
xnor U11567 (N_11567,N_11467,N_11532);
nand U11568 (N_11568,N_11549,N_11493);
and U11569 (N_11569,N_11462,N_11418);
and U11570 (N_11570,N_11410,N_11518);
or U11571 (N_11571,N_11538,N_11437);
and U11572 (N_11572,N_11528,N_11480);
nand U11573 (N_11573,N_11463,N_11419);
nand U11574 (N_11574,N_11504,N_11498);
nor U11575 (N_11575,N_11426,N_11469);
and U11576 (N_11576,N_11522,N_11416);
or U11577 (N_11577,N_11490,N_11440);
nand U11578 (N_11578,N_11406,N_11475);
nand U11579 (N_11579,N_11488,N_11505);
and U11580 (N_11580,N_11421,N_11402);
nor U11581 (N_11581,N_11424,N_11514);
nand U11582 (N_11582,N_11435,N_11525);
nor U11583 (N_11583,N_11442,N_11457);
xor U11584 (N_11584,N_11464,N_11546);
or U11585 (N_11585,N_11527,N_11523);
nor U11586 (N_11586,N_11520,N_11453);
and U11587 (N_11587,N_11451,N_11534);
or U11588 (N_11588,N_11486,N_11517);
or U11589 (N_11589,N_11470,N_11545);
nand U11590 (N_11590,N_11407,N_11444);
nand U11591 (N_11591,N_11541,N_11432);
and U11592 (N_11592,N_11506,N_11509);
nor U11593 (N_11593,N_11401,N_11417);
xnor U11594 (N_11594,N_11413,N_11479);
nand U11595 (N_11595,N_11405,N_11445);
and U11596 (N_11596,N_11516,N_11489);
and U11597 (N_11597,N_11429,N_11433);
or U11598 (N_11598,N_11533,N_11537);
nor U11599 (N_11599,N_11529,N_11414);
or U11600 (N_11600,N_11508,N_11420);
xnor U11601 (N_11601,N_11492,N_11536);
or U11602 (N_11602,N_11531,N_11411);
nor U11603 (N_11603,N_11543,N_11465);
xnor U11604 (N_11604,N_11526,N_11450);
xnor U11605 (N_11605,N_11409,N_11476);
nand U11606 (N_11606,N_11521,N_11499);
nor U11607 (N_11607,N_11422,N_11500);
nor U11608 (N_11608,N_11547,N_11454);
nor U11609 (N_11609,N_11481,N_11511);
nor U11610 (N_11610,N_11483,N_11400);
xnor U11611 (N_11611,N_11495,N_11404);
nor U11612 (N_11612,N_11519,N_11544);
nand U11613 (N_11613,N_11427,N_11456);
nor U11614 (N_11614,N_11415,N_11452);
or U11615 (N_11615,N_11512,N_11468);
and U11616 (N_11616,N_11496,N_11501);
nor U11617 (N_11617,N_11460,N_11434);
and U11618 (N_11618,N_11466,N_11494);
xnor U11619 (N_11619,N_11487,N_11477);
xor U11620 (N_11620,N_11474,N_11540);
nor U11621 (N_11621,N_11441,N_11458);
nor U11622 (N_11622,N_11485,N_11403);
nor U11623 (N_11623,N_11510,N_11503);
nand U11624 (N_11624,N_11447,N_11507);
nand U11625 (N_11625,N_11524,N_11530);
nand U11626 (N_11626,N_11490,N_11491);
nor U11627 (N_11627,N_11531,N_11427);
xnor U11628 (N_11628,N_11432,N_11495);
xnor U11629 (N_11629,N_11412,N_11503);
and U11630 (N_11630,N_11468,N_11459);
xnor U11631 (N_11631,N_11483,N_11515);
or U11632 (N_11632,N_11514,N_11468);
nand U11633 (N_11633,N_11440,N_11503);
xnor U11634 (N_11634,N_11417,N_11457);
or U11635 (N_11635,N_11420,N_11483);
and U11636 (N_11636,N_11516,N_11409);
nor U11637 (N_11637,N_11471,N_11482);
and U11638 (N_11638,N_11485,N_11413);
and U11639 (N_11639,N_11468,N_11520);
and U11640 (N_11640,N_11502,N_11412);
or U11641 (N_11641,N_11520,N_11459);
nand U11642 (N_11642,N_11419,N_11405);
xnor U11643 (N_11643,N_11544,N_11548);
nor U11644 (N_11644,N_11491,N_11530);
or U11645 (N_11645,N_11463,N_11532);
or U11646 (N_11646,N_11514,N_11459);
and U11647 (N_11647,N_11508,N_11438);
and U11648 (N_11648,N_11467,N_11444);
and U11649 (N_11649,N_11429,N_11426);
nor U11650 (N_11650,N_11475,N_11492);
nand U11651 (N_11651,N_11432,N_11526);
and U11652 (N_11652,N_11511,N_11544);
or U11653 (N_11653,N_11413,N_11527);
nor U11654 (N_11654,N_11447,N_11400);
xnor U11655 (N_11655,N_11517,N_11419);
and U11656 (N_11656,N_11529,N_11436);
nand U11657 (N_11657,N_11521,N_11450);
nand U11658 (N_11658,N_11484,N_11462);
or U11659 (N_11659,N_11538,N_11507);
nor U11660 (N_11660,N_11425,N_11487);
or U11661 (N_11661,N_11483,N_11536);
nand U11662 (N_11662,N_11502,N_11543);
or U11663 (N_11663,N_11543,N_11487);
xnor U11664 (N_11664,N_11548,N_11405);
and U11665 (N_11665,N_11501,N_11490);
nor U11666 (N_11666,N_11469,N_11406);
or U11667 (N_11667,N_11405,N_11426);
nand U11668 (N_11668,N_11464,N_11414);
xor U11669 (N_11669,N_11447,N_11459);
nand U11670 (N_11670,N_11458,N_11497);
and U11671 (N_11671,N_11441,N_11451);
nor U11672 (N_11672,N_11480,N_11458);
or U11673 (N_11673,N_11411,N_11477);
nand U11674 (N_11674,N_11487,N_11535);
and U11675 (N_11675,N_11503,N_11420);
nand U11676 (N_11676,N_11416,N_11449);
nor U11677 (N_11677,N_11492,N_11472);
nor U11678 (N_11678,N_11535,N_11541);
xor U11679 (N_11679,N_11429,N_11404);
nand U11680 (N_11680,N_11517,N_11412);
xnor U11681 (N_11681,N_11526,N_11504);
xnor U11682 (N_11682,N_11529,N_11511);
and U11683 (N_11683,N_11442,N_11496);
and U11684 (N_11684,N_11503,N_11511);
nand U11685 (N_11685,N_11447,N_11421);
xor U11686 (N_11686,N_11536,N_11528);
nand U11687 (N_11687,N_11498,N_11438);
nand U11688 (N_11688,N_11515,N_11497);
or U11689 (N_11689,N_11548,N_11538);
or U11690 (N_11690,N_11514,N_11538);
nand U11691 (N_11691,N_11408,N_11421);
nor U11692 (N_11692,N_11411,N_11503);
xor U11693 (N_11693,N_11448,N_11435);
nor U11694 (N_11694,N_11479,N_11546);
xor U11695 (N_11695,N_11507,N_11521);
nand U11696 (N_11696,N_11434,N_11435);
nor U11697 (N_11697,N_11528,N_11456);
nor U11698 (N_11698,N_11472,N_11545);
nor U11699 (N_11699,N_11413,N_11469);
and U11700 (N_11700,N_11620,N_11635);
or U11701 (N_11701,N_11673,N_11699);
xor U11702 (N_11702,N_11562,N_11601);
xor U11703 (N_11703,N_11643,N_11588);
nor U11704 (N_11704,N_11616,N_11647);
or U11705 (N_11705,N_11671,N_11644);
and U11706 (N_11706,N_11609,N_11606);
nor U11707 (N_11707,N_11667,N_11555);
and U11708 (N_11708,N_11633,N_11629);
xnor U11709 (N_11709,N_11589,N_11657);
xnor U11710 (N_11710,N_11557,N_11655);
and U11711 (N_11711,N_11551,N_11582);
and U11712 (N_11712,N_11651,N_11691);
nor U11713 (N_11713,N_11613,N_11670);
nand U11714 (N_11714,N_11672,N_11685);
and U11715 (N_11715,N_11576,N_11554);
and U11716 (N_11716,N_11624,N_11563);
or U11717 (N_11717,N_11638,N_11631);
or U11718 (N_11718,N_11634,N_11607);
or U11719 (N_11719,N_11664,N_11580);
nor U11720 (N_11720,N_11566,N_11642);
nand U11721 (N_11721,N_11608,N_11679);
nor U11722 (N_11722,N_11641,N_11560);
and U11723 (N_11723,N_11577,N_11684);
nor U11724 (N_11724,N_11586,N_11660);
xnor U11725 (N_11725,N_11668,N_11661);
or U11726 (N_11726,N_11570,N_11688);
or U11727 (N_11727,N_11597,N_11678);
xnor U11728 (N_11728,N_11675,N_11689);
or U11729 (N_11729,N_11697,N_11579);
nand U11730 (N_11730,N_11604,N_11677);
xor U11731 (N_11731,N_11578,N_11599);
and U11732 (N_11732,N_11662,N_11611);
nor U11733 (N_11733,N_11571,N_11621);
and U11734 (N_11734,N_11594,N_11610);
nand U11735 (N_11735,N_11619,N_11612);
and U11736 (N_11736,N_11694,N_11686);
nor U11737 (N_11737,N_11569,N_11598);
nand U11738 (N_11738,N_11639,N_11654);
nand U11739 (N_11739,N_11592,N_11663);
nand U11740 (N_11740,N_11623,N_11565);
xor U11741 (N_11741,N_11605,N_11676);
xnor U11742 (N_11742,N_11567,N_11614);
nor U11743 (N_11743,N_11618,N_11627);
nor U11744 (N_11744,N_11559,N_11674);
nor U11745 (N_11745,N_11682,N_11665);
nand U11746 (N_11746,N_11575,N_11652);
xor U11747 (N_11747,N_11659,N_11587);
xor U11748 (N_11748,N_11585,N_11593);
xnor U11749 (N_11749,N_11602,N_11572);
xor U11750 (N_11750,N_11574,N_11692);
or U11751 (N_11751,N_11637,N_11687);
or U11752 (N_11752,N_11581,N_11656);
nor U11753 (N_11753,N_11658,N_11553);
or U11754 (N_11754,N_11630,N_11622);
xnor U11755 (N_11755,N_11632,N_11653);
xor U11756 (N_11756,N_11646,N_11583);
nor U11757 (N_11757,N_11556,N_11615);
nor U11758 (N_11758,N_11669,N_11695);
and U11759 (N_11759,N_11693,N_11573);
nor U11760 (N_11760,N_11595,N_11564);
or U11761 (N_11761,N_11625,N_11690);
nor U11762 (N_11762,N_11552,N_11666);
nand U11763 (N_11763,N_11626,N_11648);
or U11764 (N_11764,N_11683,N_11617);
nor U11765 (N_11765,N_11600,N_11603);
nand U11766 (N_11766,N_11628,N_11558);
nand U11767 (N_11767,N_11568,N_11640);
nand U11768 (N_11768,N_11584,N_11650);
and U11769 (N_11769,N_11636,N_11681);
nand U11770 (N_11770,N_11698,N_11645);
or U11771 (N_11771,N_11591,N_11696);
xor U11772 (N_11772,N_11590,N_11561);
nand U11773 (N_11773,N_11649,N_11550);
nor U11774 (N_11774,N_11596,N_11680);
nand U11775 (N_11775,N_11605,N_11699);
nand U11776 (N_11776,N_11683,N_11663);
and U11777 (N_11777,N_11654,N_11695);
nor U11778 (N_11778,N_11608,N_11577);
nor U11779 (N_11779,N_11558,N_11636);
nand U11780 (N_11780,N_11692,N_11602);
nor U11781 (N_11781,N_11589,N_11570);
and U11782 (N_11782,N_11594,N_11631);
xnor U11783 (N_11783,N_11569,N_11556);
nor U11784 (N_11784,N_11694,N_11550);
or U11785 (N_11785,N_11669,N_11614);
nand U11786 (N_11786,N_11672,N_11598);
nor U11787 (N_11787,N_11620,N_11693);
nand U11788 (N_11788,N_11655,N_11619);
or U11789 (N_11789,N_11621,N_11589);
nor U11790 (N_11790,N_11671,N_11589);
nand U11791 (N_11791,N_11599,N_11640);
nor U11792 (N_11792,N_11671,N_11639);
and U11793 (N_11793,N_11631,N_11588);
and U11794 (N_11794,N_11662,N_11694);
nand U11795 (N_11795,N_11569,N_11633);
and U11796 (N_11796,N_11600,N_11662);
nand U11797 (N_11797,N_11585,N_11570);
xnor U11798 (N_11798,N_11560,N_11691);
nor U11799 (N_11799,N_11650,N_11647);
and U11800 (N_11800,N_11606,N_11631);
and U11801 (N_11801,N_11641,N_11585);
and U11802 (N_11802,N_11556,N_11632);
nor U11803 (N_11803,N_11645,N_11625);
nand U11804 (N_11804,N_11652,N_11569);
and U11805 (N_11805,N_11669,N_11577);
xnor U11806 (N_11806,N_11555,N_11646);
or U11807 (N_11807,N_11551,N_11597);
nor U11808 (N_11808,N_11551,N_11642);
and U11809 (N_11809,N_11626,N_11571);
nand U11810 (N_11810,N_11573,N_11624);
nor U11811 (N_11811,N_11578,N_11638);
nand U11812 (N_11812,N_11587,N_11644);
and U11813 (N_11813,N_11558,N_11691);
and U11814 (N_11814,N_11574,N_11698);
and U11815 (N_11815,N_11566,N_11585);
or U11816 (N_11816,N_11595,N_11644);
or U11817 (N_11817,N_11591,N_11669);
and U11818 (N_11818,N_11631,N_11667);
xnor U11819 (N_11819,N_11603,N_11586);
xor U11820 (N_11820,N_11679,N_11650);
or U11821 (N_11821,N_11554,N_11615);
xor U11822 (N_11822,N_11594,N_11628);
or U11823 (N_11823,N_11578,N_11637);
or U11824 (N_11824,N_11631,N_11562);
xnor U11825 (N_11825,N_11571,N_11608);
or U11826 (N_11826,N_11619,N_11653);
or U11827 (N_11827,N_11679,N_11586);
nand U11828 (N_11828,N_11688,N_11626);
or U11829 (N_11829,N_11653,N_11687);
nand U11830 (N_11830,N_11630,N_11559);
and U11831 (N_11831,N_11581,N_11552);
nand U11832 (N_11832,N_11682,N_11616);
nand U11833 (N_11833,N_11671,N_11585);
and U11834 (N_11834,N_11686,N_11565);
and U11835 (N_11835,N_11692,N_11667);
xor U11836 (N_11836,N_11648,N_11632);
and U11837 (N_11837,N_11635,N_11610);
and U11838 (N_11838,N_11666,N_11676);
and U11839 (N_11839,N_11587,N_11641);
or U11840 (N_11840,N_11647,N_11681);
nand U11841 (N_11841,N_11640,N_11686);
nor U11842 (N_11842,N_11642,N_11698);
nor U11843 (N_11843,N_11698,N_11685);
or U11844 (N_11844,N_11566,N_11601);
xnor U11845 (N_11845,N_11599,N_11572);
and U11846 (N_11846,N_11651,N_11600);
nand U11847 (N_11847,N_11687,N_11613);
nand U11848 (N_11848,N_11616,N_11665);
and U11849 (N_11849,N_11565,N_11690);
and U11850 (N_11850,N_11806,N_11826);
xor U11851 (N_11851,N_11727,N_11704);
xnor U11852 (N_11852,N_11825,N_11717);
and U11853 (N_11853,N_11810,N_11820);
nand U11854 (N_11854,N_11788,N_11744);
or U11855 (N_11855,N_11742,N_11736);
and U11856 (N_11856,N_11740,N_11776);
or U11857 (N_11857,N_11721,N_11706);
or U11858 (N_11858,N_11731,N_11802);
nor U11859 (N_11859,N_11803,N_11770);
nor U11860 (N_11860,N_11800,N_11749);
xnor U11861 (N_11861,N_11720,N_11796);
and U11862 (N_11862,N_11743,N_11758);
and U11863 (N_11863,N_11842,N_11748);
nand U11864 (N_11864,N_11794,N_11759);
xnor U11865 (N_11865,N_11738,N_11797);
and U11866 (N_11866,N_11832,N_11712);
and U11867 (N_11867,N_11775,N_11734);
or U11868 (N_11868,N_11715,N_11762);
xor U11869 (N_11869,N_11739,N_11790);
nor U11870 (N_11870,N_11745,N_11822);
nor U11871 (N_11871,N_11707,N_11829);
or U11872 (N_11872,N_11763,N_11753);
nand U11873 (N_11873,N_11793,N_11837);
xor U11874 (N_11874,N_11840,N_11845);
and U11875 (N_11875,N_11761,N_11816);
xor U11876 (N_11876,N_11783,N_11769);
nand U11877 (N_11877,N_11710,N_11771);
nand U11878 (N_11878,N_11765,N_11801);
xor U11879 (N_11879,N_11785,N_11756);
xnor U11880 (N_11880,N_11755,N_11773);
nand U11881 (N_11881,N_11823,N_11701);
and U11882 (N_11882,N_11804,N_11713);
xor U11883 (N_11883,N_11780,N_11774);
and U11884 (N_11884,N_11846,N_11752);
nor U11885 (N_11885,N_11784,N_11722);
or U11886 (N_11886,N_11830,N_11786);
nand U11887 (N_11887,N_11798,N_11792);
and U11888 (N_11888,N_11705,N_11811);
and U11889 (N_11889,N_11828,N_11714);
xnor U11890 (N_11890,N_11813,N_11844);
nor U11891 (N_11891,N_11737,N_11835);
xor U11892 (N_11892,N_11724,N_11709);
or U11893 (N_11893,N_11728,N_11849);
or U11894 (N_11894,N_11781,N_11700);
and U11895 (N_11895,N_11815,N_11841);
xor U11896 (N_11896,N_11809,N_11789);
or U11897 (N_11897,N_11750,N_11827);
or U11898 (N_11898,N_11807,N_11795);
xor U11899 (N_11899,N_11725,N_11791);
xor U11900 (N_11900,N_11726,N_11768);
xor U11901 (N_11901,N_11767,N_11777);
xnor U11902 (N_11902,N_11836,N_11735);
or U11903 (N_11903,N_11812,N_11843);
or U11904 (N_11904,N_11732,N_11847);
or U11905 (N_11905,N_11787,N_11834);
or U11906 (N_11906,N_11754,N_11711);
nand U11907 (N_11907,N_11838,N_11833);
nor U11908 (N_11908,N_11760,N_11772);
and U11909 (N_11909,N_11818,N_11824);
xor U11910 (N_11910,N_11799,N_11821);
or U11911 (N_11911,N_11831,N_11733);
or U11912 (N_11912,N_11702,N_11741);
nor U11913 (N_11913,N_11766,N_11764);
and U11914 (N_11914,N_11757,N_11805);
xnor U11915 (N_11915,N_11778,N_11808);
nor U11916 (N_11916,N_11814,N_11817);
xnor U11917 (N_11917,N_11839,N_11723);
nor U11918 (N_11918,N_11716,N_11719);
or U11919 (N_11919,N_11729,N_11819);
xor U11920 (N_11920,N_11751,N_11782);
nand U11921 (N_11921,N_11746,N_11708);
nor U11922 (N_11922,N_11718,N_11730);
nand U11923 (N_11923,N_11747,N_11703);
nand U11924 (N_11924,N_11779,N_11848);
nor U11925 (N_11925,N_11824,N_11804);
or U11926 (N_11926,N_11766,N_11806);
or U11927 (N_11927,N_11778,N_11752);
and U11928 (N_11928,N_11755,N_11712);
xor U11929 (N_11929,N_11815,N_11791);
nand U11930 (N_11930,N_11727,N_11847);
and U11931 (N_11931,N_11801,N_11834);
nand U11932 (N_11932,N_11708,N_11754);
nand U11933 (N_11933,N_11745,N_11709);
xor U11934 (N_11934,N_11778,N_11842);
and U11935 (N_11935,N_11758,N_11735);
or U11936 (N_11936,N_11843,N_11754);
nor U11937 (N_11937,N_11762,N_11760);
and U11938 (N_11938,N_11788,N_11808);
nand U11939 (N_11939,N_11848,N_11837);
nor U11940 (N_11940,N_11789,N_11715);
nor U11941 (N_11941,N_11782,N_11753);
nand U11942 (N_11942,N_11840,N_11702);
nand U11943 (N_11943,N_11751,N_11784);
nor U11944 (N_11944,N_11728,N_11745);
xnor U11945 (N_11945,N_11754,N_11758);
nand U11946 (N_11946,N_11788,N_11840);
xor U11947 (N_11947,N_11723,N_11709);
and U11948 (N_11948,N_11755,N_11746);
nand U11949 (N_11949,N_11758,N_11777);
or U11950 (N_11950,N_11768,N_11794);
xor U11951 (N_11951,N_11788,N_11773);
nor U11952 (N_11952,N_11702,N_11831);
nand U11953 (N_11953,N_11796,N_11815);
xor U11954 (N_11954,N_11796,N_11755);
or U11955 (N_11955,N_11794,N_11750);
nor U11956 (N_11956,N_11815,N_11788);
nor U11957 (N_11957,N_11719,N_11838);
nor U11958 (N_11958,N_11779,N_11814);
xor U11959 (N_11959,N_11743,N_11748);
and U11960 (N_11960,N_11735,N_11825);
and U11961 (N_11961,N_11826,N_11748);
or U11962 (N_11962,N_11799,N_11823);
or U11963 (N_11963,N_11807,N_11801);
nand U11964 (N_11964,N_11835,N_11709);
nand U11965 (N_11965,N_11823,N_11840);
and U11966 (N_11966,N_11702,N_11726);
nand U11967 (N_11967,N_11762,N_11714);
nand U11968 (N_11968,N_11716,N_11730);
nor U11969 (N_11969,N_11769,N_11829);
xor U11970 (N_11970,N_11761,N_11841);
nor U11971 (N_11971,N_11720,N_11799);
xor U11972 (N_11972,N_11845,N_11712);
xnor U11973 (N_11973,N_11790,N_11741);
or U11974 (N_11974,N_11839,N_11747);
or U11975 (N_11975,N_11812,N_11718);
xor U11976 (N_11976,N_11748,N_11754);
or U11977 (N_11977,N_11792,N_11700);
and U11978 (N_11978,N_11752,N_11780);
nor U11979 (N_11979,N_11800,N_11798);
and U11980 (N_11980,N_11806,N_11734);
and U11981 (N_11981,N_11794,N_11722);
or U11982 (N_11982,N_11785,N_11804);
nor U11983 (N_11983,N_11795,N_11758);
or U11984 (N_11984,N_11756,N_11791);
nand U11985 (N_11985,N_11839,N_11718);
and U11986 (N_11986,N_11821,N_11815);
nand U11987 (N_11987,N_11749,N_11713);
or U11988 (N_11988,N_11788,N_11791);
or U11989 (N_11989,N_11767,N_11727);
nand U11990 (N_11990,N_11778,N_11785);
and U11991 (N_11991,N_11728,N_11712);
nand U11992 (N_11992,N_11829,N_11754);
xnor U11993 (N_11993,N_11822,N_11778);
nor U11994 (N_11994,N_11801,N_11821);
nor U11995 (N_11995,N_11849,N_11706);
nor U11996 (N_11996,N_11780,N_11849);
nor U11997 (N_11997,N_11848,N_11827);
and U11998 (N_11998,N_11833,N_11845);
and U11999 (N_11999,N_11731,N_11837);
xnor U12000 (N_12000,N_11863,N_11986);
nand U12001 (N_12001,N_11942,N_11894);
nand U12002 (N_12002,N_11901,N_11977);
nor U12003 (N_12003,N_11889,N_11955);
or U12004 (N_12004,N_11897,N_11946);
xor U12005 (N_12005,N_11898,N_11918);
xor U12006 (N_12006,N_11872,N_11912);
nand U12007 (N_12007,N_11945,N_11974);
nor U12008 (N_12008,N_11926,N_11919);
xnor U12009 (N_12009,N_11993,N_11956);
nor U12010 (N_12010,N_11948,N_11911);
or U12011 (N_12011,N_11879,N_11874);
nor U12012 (N_12012,N_11936,N_11856);
or U12013 (N_12013,N_11937,N_11921);
or U12014 (N_12014,N_11997,N_11966);
xnor U12015 (N_12015,N_11870,N_11975);
xnor U12016 (N_12016,N_11891,N_11862);
nand U12017 (N_12017,N_11989,N_11866);
nor U12018 (N_12018,N_11960,N_11953);
xnor U12019 (N_12019,N_11859,N_11983);
nor U12020 (N_12020,N_11885,N_11924);
xor U12021 (N_12021,N_11853,N_11904);
nand U12022 (N_12022,N_11857,N_11871);
xor U12023 (N_12023,N_11878,N_11938);
nand U12024 (N_12024,N_11935,N_11855);
xor U12025 (N_12025,N_11860,N_11922);
xor U12026 (N_12026,N_11959,N_11934);
xnor U12027 (N_12027,N_11888,N_11962);
nor U12028 (N_12028,N_11927,N_11958);
nand U12029 (N_12029,N_11909,N_11964);
nor U12030 (N_12030,N_11972,N_11940);
nor U12031 (N_12031,N_11923,N_11906);
nand U12032 (N_12032,N_11984,N_11982);
nand U12033 (N_12033,N_11925,N_11932);
and U12034 (N_12034,N_11903,N_11852);
xnor U12035 (N_12035,N_11887,N_11886);
nand U12036 (N_12036,N_11913,N_11917);
nand U12037 (N_12037,N_11890,N_11861);
and U12038 (N_12038,N_11883,N_11979);
nand U12039 (N_12039,N_11876,N_11865);
nand U12040 (N_12040,N_11928,N_11971);
or U12041 (N_12041,N_11929,N_11965);
xor U12042 (N_12042,N_11882,N_11949);
and U12043 (N_12043,N_11910,N_11947);
nor U12044 (N_12044,N_11933,N_11952);
nand U12045 (N_12045,N_11994,N_11873);
or U12046 (N_12046,N_11985,N_11884);
nand U12047 (N_12047,N_11920,N_11976);
xnor U12048 (N_12048,N_11988,N_11943);
xnor U12049 (N_12049,N_11895,N_11969);
or U12050 (N_12050,N_11892,N_11967);
nor U12051 (N_12051,N_11858,N_11868);
or U12052 (N_12052,N_11899,N_11854);
or U12053 (N_12053,N_11893,N_11954);
nand U12054 (N_12054,N_11902,N_11914);
xor U12055 (N_12055,N_11850,N_11941);
nand U12056 (N_12056,N_11981,N_11999);
xor U12057 (N_12057,N_11970,N_11875);
nor U12058 (N_12058,N_11867,N_11930);
and U12059 (N_12059,N_11896,N_11944);
nand U12060 (N_12060,N_11869,N_11957);
nor U12061 (N_12061,N_11864,N_11915);
or U12062 (N_12062,N_11939,N_11992);
nor U12063 (N_12063,N_11991,N_11905);
or U12064 (N_12064,N_11978,N_11881);
nor U12065 (N_12065,N_11907,N_11968);
xor U12066 (N_12066,N_11987,N_11998);
or U12067 (N_12067,N_11908,N_11990);
and U12068 (N_12068,N_11996,N_11916);
and U12069 (N_12069,N_11931,N_11950);
xnor U12070 (N_12070,N_11851,N_11900);
and U12071 (N_12071,N_11961,N_11963);
xor U12072 (N_12072,N_11951,N_11880);
xnor U12073 (N_12073,N_11973,N_11980);
nor U12074 (N_12074,N_11877,N_11995);
nand U12075 (N_12075,N_11905,N_11888);
xnor U12076 (N_12076,N_11877,N_11859);
and U12077 (N_12077,N_11883,N_11918);
nor U12078 (N_12078,N_11992,N_11983);
xnor U12079 (N_12079,N_11886,N_11980);
nor U12080 (N_12080,N_11949,N_11980);
nor U12081 (N_12081,N_11877,N_11899);
nand U12082 (N_12082,N_11930,N_11927);
nand U12083 (N_12083,N_11895,N_11941);
or U12084 (N_12084,N_11895,N_11960);
nand U12085 (N_12085,N_11894,N_11921);
xor U12086 (N_12086,N_11992,N_11855);
and U12087 (N_12087,N_11975,N_11997);
or U12088 (N_12088,N_11971,N_11896);
nor U12089 (N_12089,N_11941,N_11966);
nor U12090 (N_12090,N_11910,N_11915);
and U12091 (N_12091,N_11866,N_11964);
and U12092 (N_12092,N_11978,N_11987);
or U12093 (N_12093,N_11953,N_11927);
xnor U12094 (N_12094,N_11875,N_11879);
nand U12095 (N_12095,N_11948,N_11906);
or U12096 (N_12096,N_11871,N_11946);
nand U12097 (N_12097,N_11935,N_11875);
xnor U12098 (N_12098,N_11979,N_11998);
or U12099 (N_12099,N_11981,N_11878);
nor U12100 (N_12100,N_11854,N_11878);
and U12101 (N_12101,N_11987,N_11964);
nor U12102 (N_12102,N_11881,N_11935);
or U12103 (N_12103,N_11909,N_11941);
or U12104 (N_12104,N_11921,N_11880);
xnor U12105 (N_12105,N_11868,N_11986);
or U12106 (N_12106,N_11995,N_11911);
or U12107 (N_12107,N_11985,N_11921);
xor U12108 (N_12108,N_11937,N_11880);
or U12109 (N_12109,N_11957,N_11871);
nor U12110 (N_12110,N_11898,N_11891);
nor U12111 (N_12111,N_11965,N_11952);
or U12112 (N_12112,N_11938,N_11999);
and U12113 (N_12113,N_11963,N_11889);
xor U12114 (N_12114,N_11866,N_11962);
and U12115 (N_12115,N_11948,N_11908);
and U12116 (N_12116,N_11857,N_11984);
and U12117 (N_12117,N_11921,N_11964);
and U12118 (N_12118,N_11919,N_11998);
nor U12119 (N_12119,N_11993,N_11970);
or U12120 (N_12120,N_11869,N_11905);
and U12121 (N_12121,N_11975,N_11965);
nor U12122 (N_12122,N_11988,N_11999);
and U12123 (N_12123,N_11932,N_11869);
and U12124 (N_12124,N_11922,N_11969);
nand U12125 (N_12125,N_11984,N_11852);
nand U12126 (N_12126,N_11887,N_11863);
nor U12127 (N_12127,N_11895,N_11905);
nor U12128 (N_12128,N_11940,N_11903);
or U12129 (N_12129,N_11861,N_11922);
and U12130 (N_12130,N_11920,N_11926);
or U12131 (N_12131,N_11854,N_11903);
nor U12132 (N_12132,N_11862,N_11890);
nor U12133 (N_12133,N_11931,N_11895);
or U12134 (N_12134,N_11891,N_11911);
nand U12135 (N_12135,N_11953,N_11978);
nand U12136 (N_12136,N_11852,N_11906);
nor U12137 (N_12137,N_11879,N_11951);
or U12138 (N_12138,N_11913,N_11956);
xor U12139 (N_12139,N_11960,N_11916);
nand U12140 (N_12140,N_11900,N_11909);
nand U12141 (N_12141,N_11857,N_11917);
or U12142 (N_12142,N_11975,N_11874);
and U12143 (N_12143,N_11913,N_11910);
and U12144 (N_12144,N_11925,N_11942);
nand U12145 (N_12145,N_11978,N_11920);
xor U12146 (N_12146,N_11916,N_11934);
or U12147 (N_12147,N_11948,N_11973);
nor U12148 (N_12148,N_11988,N_11870);
xnor U12149 (N_12149,N_11892,N_11909);
and U12150 (N_12150,N_12125,N_12043);
and U12151 (N_12151,N_12136,N_12000);
or U12152 (N_12152,N_12098,N_12116);
nand U12153 (N_12153,N_12040,N_12135);
or U12154 (N_12154,N_12063,N_12102);
or U12155 (N_12155,N_12038,N_12120);
nand U12156 (N_12156,N_12097,N_12047);
nand U12157 (N_12157,N_12096,N_12101);
and U12158 (N_12158,N_12094,N_12024);
xor U12159 (N_12159,N_12025,N_12100);
xnor U12160 (N_12160,N_12133,N_12075);
nor U12161 (N_12161,N_12067,N_12039);
xnor U12162 (N_12162,N_12031,N_12140);
nand U12163 (N_12163,N_12126,N_12121);
and U12164 (N_12164,N_12078,N_12138);
or U12165 (N_12165,N_12144,N_12026);
and U12166 (N_12166,N_12130,N_12048);
nand U12167 (N_12167,N_12035,N_12089);
nor U12168 (N_12168,N_12110,N_12131);
and U12169 (N_12169,N_12014,N_12060);
or U12170 (N_12170,N_12112,N_12088);
nand U12171 (N_12171,N_12147,N_12134);
nor U12172 (N_12172,N_12149,N_12127);
nor U12173 (N_12173,N_12137,N_12082);
and U12174 (N_12174,N_12142,N_12080);
xnor U12175 (N_12175,N_12056,N_12030);
nor U12176 (N_12176,N_12010,N_12001);
and U12177 (N_12177,N_12020,N_12057);
xor U12178 (N_12178,N_12052,N_12033);
or U12179 (N_12179,N_12087,N_12103);
and U12180 (N_12180,N_12058,N_12036);
nand U12181 (N_12181,N_12064,N_12093);
and U12182 (N_12182,N_12049,N_12046);
xor U12183 (N_12183,N_12041,N_12105);
xor U12184 (N_12184,N_12005,N_12143);
or U12185 (N_12185,N_12028,N_12129);
nand U12186 (N_12186,N_12077,N_12109);
xnor U12187 (N_12187,N_12104,N_12084);
nand U12188 (N_12188,N_12081,N_12118);
xor U12189 (N_12189,N_12122,N_12062);
nor U12190 (N_12190,N_12090,N_12059);
and U12191 (N_12191,N_12021,N_12074);
or U12192 (N_12192,N_12011,N_12017);
and U12193 (N_12193,N_12092,N_12108);
nand U12194 (N_12194,N_12085,N_12071);
or U12195 (N_12195,N_12006,N_12032);
or U12196 (N_12196,N_12128,N_12076);
nor U12197 (N_12197,N_12013,N_12061);
nand U12198 (N_12198,N_12065,N_12073);
nand U12199 (N_12199,N_12007,N_12027);
xor U12200 (N_12200,N_12012,N_12051);
nor U12201 (N_12201,N_12015,N_12066);
nand U12202 (N_12202,N_12083,N_12044);
and U12203 (N_12203,N_12114,N_12139);
xor U12204 (N_12204,N_12069,N_12123);
nor U12205 (N_12205,N_12008,N_12050);
nand U12206 (N_12206,N_12106,N_12117);
and U12207 (N_12207,N_12068,N_12003);
and U12208 (N_12208,N_12042,N_12009);
and U12209 (N_12209,N_12086,N_12099);
nand U12210 (N_12210,N_12079,N_12019);
xnor U12211 (N_12211,N_12115,N_12141);
xor U12212 (N_12212,N_12004,N_12029);
xnor U12213 (N_12213,N_12072,N_12016);
nor U12214 (N_12214,N_12119,N_12002);
and U12215 (N_12215,N_12018,N_12148);
nand U12216 (N_12216,N_12055,N_12070);
or U12217 (N_12217,N_12145,N_12023);
and U12218 (N_12218,N_12091,N_12034);
xnor U12219 (N_12219,N_12054,N_12095);
nand U12220 (N_12220,N_12045,N_12037);
or U12221 (N_12221,N_12111,N_12053);
and U12222 (N_12222,N_12022,N_12132);
or U12223 (N_12223,N_12146,N_12113);
xnor U12224 (N_12224,N_12124,N_12107);
xor U12225 (N_12225,N_12146,N_12032);
nor U12226 (N_12226,N_12134,N_12069);
nor U12227 (N_12227,N_12145,N_12092);
xor U12228 (N_12228,N_12065,N_12071);
xor U12229 (N_12229,N_12118,N_12067);
and U12230 (N_12230,N_12008,N_12033);
nand U12231 (N_12231,N_12131,N_12148);
and U12232 (N_12232,N_12087,N_12124);
nor U12233 (N_12233,N_12072,N_12012);
xnor U12234 (N_12234,N_12061,N_12014);
and U12235 (N_12235,N_12032,N_12026);
and U12236 (N_12236,N_12131,N_12058);
xnor U12237 (N_12237,N_12058,N_12031);
nor U12238 (N_12238,N_12032,N_12015);
nor U12239 (N_12239,N_12065,N_12137);
nand U12240 (N_12240,N_12002,N_12126);
nor U12241 (N_12241,N_12046,N_12030);
and U12242 (N_12242,N_12026,N_12056);
nor U12243 (N_12243,N_12149,N_12007);
or U12244 (N_12244,N_12014,N_12077);
or U12245 (N_12245,N_12046,N_12047);
or U12246 (N_12246,N_12129,N_12146);
and U12247 (N_12247,N_12114,N_12015);
nand U12248 (N_12248,N_12101,N_12007);
and U12249 (N_12249,N_12033,N_12127);
xor U12250 (N_12250,N_12006,N_12146);
nor U12251 (N_12251,N_12081,N_12093);
nor U12252 (N_12252,N_12087,N_12077);
or U12253 (N_12253,N_12013,N_12131);
xor U12254 (N_12254,N_12062,N_12119);
or U12255 (N_12255,N_12075,N_12076);
nand U12256 (N_12256,N_12085,N_12059);
nand U12257 (N_12257,N_12082,N_12036);
xor U12258 (N_12258,N_12114,N_12007);
nor U12259 (N_12259,N_12069,N_12130);
and U12260 (N_12260,N_12045,N_12047);
and U12261 (N_12261,N_12005,N_12070);
xnor U12262 (N_12262,N_12008,N_12046);
and U12263 (N_12263,N_12038,N_12006);
nor U12264 (N_12264,N_12075,N_12069);
nor U12265 (N_12265,N_12036,N_12056);
xor U12266 (N_12266,N_12139,N_12131);
or U12267 (N_12267,N_12027,N_12092);
or U12268 (N_12268,N_12038,N_12121);
nor U12269 (N_12269,N_12066,N_12080);
nand U12270 (N_12270,N_12122,N_12093);
and U12271 (N_12271,N_12033,N_12086);
xnor U12272 (N_12272,N_12066,N_12148);
nand U12273 (N_12273,N_12027,N_12104);
nand U12274 (N_12274,N_12010,N_12138);
or U12275 (N_12275,N_12146,N_12132);
and U12276 (N_12276,N_12070,N_12058);
or U12277 (N_12277,N_12042,N_12143);
xor U12278 (N_12278,N_12139,N_12100);
or U12279 (N_12279,N_12100,N_12070);
nand U12280 (N_12280,N_12026,N_12022);
xnor U12281 (N_12281,N_12136,N_12106);
and U12282 (N_12282,N_12081,N_12139);
nor U12283 (N_12283,N_12137,N_12138);
nand U12284 (N_12284,N_12124,N_12045);
nand U12285 (N_12285,N_12088,N_12107);
nand U12286 (N_12286,N_12056,N_12137);
or U12287 (N_12287,N_12128,N_12060);
nand U12288 (N_12288,N_12130,N_12013);
nand U12289 (N_12289,N_12053,N_12117);
xor U12290 (N_12290,N_12017,N_12094);
or U12291 (N_12291,N_12006,N_12103);
or U12292 (N_12292,N_12062,N_12096);
nand U12293 (N_12293,N_12013,N_12049);
or U12294 (N_12294,N_12096,N_12014);
xnor U12295 (N_12295,N_12010,N_12140);
xnor U12296 (N_12296,N_12034,N_12107);
xnor U12297 (N_12297,N_12147,N_12094);
nand U12298 (N_12298,N_12054,N_12131);
nand U12299 (N_12299,N_12020,N_12063);
xnor U12300 (N_12300,N_12257,N_12196);
or U12301 (N_12301,N_12245,N_12298);
nor U12302 (N_12302,N_12268,N_12240);
or U12303 (N_12303,N_12182,N_12188);
xnor U12304 (N_12304,N_12152,N_12189);
nand U12305 (N_12305,N_12265,N_12237);
and U12306 (N_12306,N_12234,N_12204);
and U12307 (N_12307,N_12158,N_12186);
and U12308 (N_12308,N_12166,N_12230);
xnor U12309 (N_12309,N_12161,N_12267);
nor U12310 (N_12310,N_12259,N_12222);
xor U12311 (N_12311,N_12178,N_12205);
xnor U12312 (N_12312,N_12180,N_12275);
and U12313 (N_12313,N_12209,N_12197);
and U12314 (N_12314,N_12170,N_12253);
and U12315 (N_12315,N_12194,N_12242);
and U12316 (N_12316,N_12271,N_12216);
nor U12317 (N_12317,N_12262,N_12248);
and U12318 (N_12318,N_12278,N_12235);
xnor U12319 (N_12319,N_12206,N_12174);
or U12320 (N_12320,N_12281,N_12159);
or U12321 (N_12321,N_12241,N_12173);
or U12322 (N_12322,N_12282,N_12263);
or U12323 (N_12323,N_12215,N_12277);
or U12324 (N_12324,N_12199,N_12162);
nand U12325 (N_12325,N_12295,N_12157);
and U12326 (N_12326,N_12255,N_12283);
nand U12327 (N_12327,N_12276,N_12214);
nor U12328 (N_12328,N_12231,N_12184);
nand U12329 (N_12329,N_12286,N_12198);
or U12330 (N_12330,N_12250,N_12254);
nand U12331 (N_12331,N_12249,N_12287);
nor U12332 (N_12332,N_12229,N_12191);
or U12333 (N_12333,N_12238,N_12181);
or U12334 (N_12334,N_12280,N_12270);
nand U12335 (N_12335,N_12273,N_12172);
and U12336 (N_12336,N_12227,N_12296);
nor U12337 (N_12337,N_12176,N_12261);
nor U12338 (N_12338,N_12165,N_12274);
nor U12339 (N_12339,N_12290,N_12297);
nand U12340 (N_12340,N_12244,N_12200);
and U12341 (N_12341,N_12272,N_12247);
xnor U12342 (N_12342,N_12156,N_12167);
nand U12343 (N_12343,N_12284,N_12177);
nor U12344 (N_12344,N_12236,N_12285);
nor U12345 (N_12345,N_12169,N_12201);
nor U12346 (N_12346,N_12258,N_12226);
or U12347 (N_12347,N_12223,N_12232);
or U12348 (N_12348,N_12155,N_12211);
or U12349 (N_12349,N_12264,N_12171);
or U12350 (N_12350,N_12202,N_12299);
or U12351 (N_12351,N_12218,N_12224);
nor U12352 (N_12352,N_12168,N_12210);
and U12353 (N_12353,N_12239,N_12203);
and U12354 (N_12354,N_12221,N_12294);
xnor U12355 (N_12355,N_12183,N_12150);
nand U12356 (N_12356,N_12251,N_12233);
xnor U12357 (N_12357,N_12193,N_12192);
nor U12358 (N_12358,N_12208,N_12293);
nor U12359 (N_12359,N_12164,N_12269);
and U12360 (N_12360,N_12190,N_12187);
and U12361 (N_12361,N_12217,N_12179);
nand U12362 (N_12362,N_12151,N_12260);
nor U12363 (N_12363,N_12288,N_12212);
nor U12364 (N_12364,N_12163,N_12289);
or U12365 (N_12365,N_12252,N_12153);
nor U12366 (N_12366,N_12279,N_12291);
nor U12367 (N_12367,N_12207,N_12160);
or U12368 (N_12368,N_12185,N_12154);
or U12369 (N_12369,N_12246,N_12220);
and U12370 (N_12370,N_12219,N_12266);
xnor U12371 (N_12371,N_12195,N_12243);
and U12372 (N_12372,N_12225,N_12228);
or U12373 (N_12373,N_12213,N_12256);
or U12374 (N_12374,N_12175,N_12292);
nor U12375 (N_12375,N_12267,N_12201);
nor U12376 (N_12376,N_12268,N_12228);
xor U12377 (N_12377,N_12204,N_12172);
or U12378 (N_12378,N_12201,N_12184);
and U12379 (N_12379,N_12218,N_12193);
nor U12380 (N_12380,N_12214,N_12215);
nand U12381 (N_12381,N_12218,N_12196);
or U12382 (N_12382,N_12201,N_12160);
xnor U12383 (N_12383,N_12203,N_12165);
nand U12384 (N_12384,N_12179,N_12151);
and U12385 (N_12385,N_12228,N_12266);
nand U12386 (N_12386,N_12246,N_12163);
nor U12387 (N_12387,N_12295,N_12234);
and U12388 (N_12388,N_12175,N_12239);
nand U12389 (N_12389,N_12230,N_12213);
or U12390 (N_12390,N_12205,N_12176);
nand U12391 (N_12391,N_12251,N_12279);
xnor U12392 (N_12392,N_12229,N_12299);
xnor U12393 (N_12393,N_12184,N_12217);
and U12394 (N_12394,N_12220,N_12244);
or U12395 (N_12395,N_12255,N_12223);
nor U12396 (N_12396,N_12272,N_12210);
and U12397 (N_12397,N_12267,N_12217);
nor U12398 (N_12398,N_12209,N_12279);
xnor U12399 (N_12399,N_12231,N_12269);
or U12400 (N_12400,N_12168,N_12251);
and U12401 (N_12401,N_12291,N_12170);
or U12402 (N_12402,N_12167,N_12224);
nor U12403 (N_12403,N_12219,N_12190);
xor U12404 (N_12404,N_12250,N_12187);
xnor U12405 (N_12405,N_12223,N_12241);
or U12406 (N_12406,N_12269,N_12289);
nor U12407 (N_12407,N_12233,N_12189);
xor U12408 (N_12408,N_12170,N_12177);
nand U12409 (N_12409,N_12227,N_12249);
and U12410 (N_12410,N_12279,N_12282);
nand U12411 (N_12411,N_12151,N_12186);
and U12412 (N_12412,N_12201,N_12245);
nand U12413 (N_12413,N_12166,N_12172);
or U12414 (N_12414,N_12262,N_12192);
nor U12415 (N_12415,N_12218,N_12150);
or U12416 (N_12416,N_12182,N_12254);
and U12417 (N_12417,N_12281,N_12237);
nor U12418 (N_12418,N_12174,N_12261);
nor U12419 (N_12419,N_12292,N_12156);
nand U12420 (N_12420,N_12260,N_12168);
xor U12421 (N_12421,N_12180,N_12257);
and U12422 (N_12422,N_12186,N_12189);
and U12423 (N_12423,N_12298,N_12250);
or U12424 (N_12424,N_12163,N_12250);
xor U12425 (N_12425,N_12182,N_12248);
xor U12426 (N_12426,N_12292,N_12189);
xor U12427 (N_12427,N_12254,N_12237);
nor U12428 (N_12428,N_12166,N_12164);
xor U12429 (N_12429,N_12153,N_12255);
nand U12430 (N_12430,N_12266,N_12202);
nor U12431 (N_12431,N_12170,N_12195);
nand U12432 (N_12432,N_12256,N_12221);
nand U12433 (N_12433,N_12259,N_12162);
or U12434 (N_12434,N_12205,N_12280);
or U12435 (N_12435,N_12169,N_12217);
nand U12436 (N_12436,N_12295,N_12261);
or U12437 (N_12437,N_12173,N_12232);
xor U12438 (N_12438,N_12190,N_12162);
or U12439 (N_12439,N_12169,N_12203);
or U12440 (N_12440,N_12160,N_12229);
nor U12441 (N_12441,N_12287,N_12214);
xor U12442 (N_12442,N_12259,N_12193);
xor U12443 (N_12443,N_12209,N_12227);
or U12444 (N_12444,N_12268,N_12242);
nand U12445 (N_12445,N_12280,N_12175);
or U12446 (N_12446,N_12152,N_12222);
or U12447 (N_12447,N_12269,N_12251);
or U12448 (N_12448,N_12159,N_12202);
nand U12449 (N_12449,N_12291,N_12268);
xnor U12450 (N_12450,N_12364,N_12333);
and U12451 (N_12451,N_12353,N_12428);
or U12452 (N_12452,N_12416,N_12404);
nor U12453 (N_12453,N_12396,N_12310);
nor U12454 (N_12454,N_12447,N_12394);
or U12455 (N_12455,N_12331,N_12444);
or U12456 (N_12456,N_12442,N_12322);
nand U12457 (N_12457,N_12448,N_12405);
xnor U12458 (N_12458,N_12374,N_12362);
nor U12459 (N_12459,N_12412,N_12318);
nand U12460 (N_12460,N_12383,N_12425);
nor U12461 (N_12461,N_12367,N_12373);
xor U12462 (N_12462,N_12351,N_12363);
nand U12463 (N_12463,N_12323,N_12431);
xor U12464 (N_12464,N_12346,N_12314);
nor U12465 (N_12465,N_12382,N_12427);
or U12466 (N_12466,N_12319,N_12342);
or U12467 (N_12467,N_12399,N_12417);
xor U12468 (N_12468,N_12301,N_12419);
and U12469 (N_12469,N_12380,N_12391);
and U12470 (N_12470,N_12359,N_12326);
or U12471 (N_12471,N_12377,N_12343);
xor U12472 (N_12472,N_12408,N_12354);
or U12473 (N_12473,N_12386,N_12324);
nand U12474 (N_12474,N_12340,N_12316);
xor U12475 (N_12475,N_12423,N_12437);
nand U12476 (N_12476,N_12446,N_12360);
xnor U12477 (N_12477,N_12349,N_12372);
xnor U12478 (N_12478,N_12411,N_12376);
xor U12479 (N_12479,N_12369,N_12356);
and U12480 (N_12480,N_12317,N_12371);
nor U12481 (N_12481,N_12312,N_12433);
nand U12482 (N_12482,N_12387,N_12361);
and U12483 (N_12483,N_12426,N_12395);
nand U12484 (N_12484,N_12375,N_12401);
nor U12485 (N_12485,N_12339,N_12300);
xnor U12486 (N_12486,N_12332,N_12379);
nor U12487 (N_12487,N_12422,N_12303);
nor U12488 (N_12488,N_12305,N_12306);
and U12489 (N_12489,N_12440,N_12388);
xnor U12490 (N_12490,N_12410,N_12304);
xor U12491 (N_12491,N_12415,N_12420);
nand U12492 (N_12492,N_12355,N_12325);
nor U12493 (N_12493,N_12350,N_12403);
or U12494 (N_12494,N_12368,N_12344);
or U12495 (N_12495,N_12439,N_12414);
nand U12496 (N_12496,N_12429,N_12315);
nand U12497 (N_12497,N_12432,N_12358);
nor U12498 (N_12498,N_12413,N_12424);
and U12499 (N_12499,N_12441,N_12378);
or U12500 (N_12500,N_12370,N_12334);
nor U12501 (N_12501,N_12313,N_12435);
nand U12502 (N_12502,N_12328,N_12335);
nand U12503 (N_12503,N_12345,N_12308);
nor U12504 (N_12504,N_12418,N_12320);
nor U12505 (N_12505,N_12327,N_12337);
xor U12506 (N_12506,N_12436,N_12357);
and U12507 (N_12507,N_12393,N_12397);
and U12508 (N_12508,N_12309,N_12398);
or U12509 (N_12509,N_12341,N_12347);
nor U12510 (N_12510,N_12385,N_12321);
and U12511 (N_12511,N_12443,N_12302);
xor U12512 (N_12512,N_12389,N_12330);
xor U12513 (N_12513,N_12402,N_12348);
and U12514 (N_12514,N_12445,N_12366);
or U12515 (N_12515,N_12400,N_12421);
nand U12516 (N_12516,N_12390,N_12430);
and U12517 (N_12517,N_12384,N_12352);
and U12518 (N_12518,N_12434,N_12409);
nor U12519 (N_12519,N_12449,N_12311);
or U12520 (N_12520,N_12406,N_12381);
xor U12521 (N_12521,N_12438,N_12336);
xor U12522 (N_12522,N_12392,N_12365);
xnor U12523 (N_12523,N_12338,N_12307);
nand U12524 (N_12524,N_12407,N_12329);
and U12525 (N_12525,N_12326,N_12330);
nor U12526 (N_12526,N_12387,N_12355);
nand U12527 (N_12527,N_12423,N_12435);
nand U12528 (N_12528,N_12327,N_12446);
and U12529 (N_12529,N_12345,N_12340);
nor U12530 (N_12530,N_12374,N_12371);
nor U12531 (N_12531,N_12307,N_12406);
nor U12532 (N_12532,N_12447,N_12423);
nor U12533 (N_12533,N_12338,N_12334);
nand U12534 (N_12534,N_12372,N_12420);
or U12535 (N_12535,N_12442,N_12311);
xnor U12536 (N_12536,N_12449,N_12316);
nor U12537 (N_12537,N_12419,N_12438);
or U12538 (N_12538,N_12387,N_12329);
nand U12539 (N_12539,N_12427,N_12301);
or U12540 (N_12540,N_12440,N_12355);
or U12541 (N_12541,N_12330,N_12409);
or U12542 (N_12542,N_12304,N_12343);
nand U12543 (N_12543,N_12304,N_12440);
nand U12544 (N_12544,N_12384,N_12439);
xor U12545 (N_12545,N_12336,N_12370);
nand U12546 (N_12546,N_12310,N_12317);
and U12547 (N_12547,N_12388,N_12433);
and U12548 (N_12548,N_12329,N_12312);
xor U12549 (N_12549,N_12442,N_12434);
and U12550 (N_12550,N_12400,N_12325);
nand U12551 (N_12551,N_12414,N_12373);
nor U12552 (N_12552,N_12357,N_12344);
or U12553 (N_12553,N_12319,N_12315);
or U12554 (N_12554,N_12343,N_12400);
xnor U12555 (N_12555,N_12323,N_12385);
nor U12556 (N_12556,N_12359,N_12310);
xor U12557 (N_12557,N_12377,N_12329);
xor U12558 (N_12558,N_12396,N_12425);
nor U12559 (N_12559,N_12311,N_12440);
and U12560 (N_12560,N_12432,N_12363);
or U12561 (N_12561,N_12386,N_12346);
nand U12562 (N_12562,N_12359,N_12402);
and U12563 (N_12563,N_12322,N_12361);
nor U12564 (N_12564,N_12329,N_12402);
nand U12565 (N_12565,N_12317,N_12338);
nand U12566 (N_12566,N_12383,N_12419);
nand U12567 (N_12567,N_12411,N_12335);
or U12568 (N_12568,N_12423,N_12446);
or U12569 (N_12569,N_12380,N_12355);
or U12570 (N_12570,N_12378,N_12401);
xnor U12571 (N_12571,N_12323,N_12313);
nand U12572 (N_12572,N_12327,N_12430);
or U12573 (N_12573,N_12354,N_12413);
and U12574 (N_12574,N_12393,N_12418);
nand U12575 (N_12575,N_12413,N_12318);
and U12576 (N_12576,N_12354,N_12389);
and U12577 (N_12577,N_12399,N_12434);
and U12578 (N_12578,N_12326,N_12334);
or U12579 (N_12579,N_12368,N_12392);
or U12580 (N_12580,N_12339,N_12383);
or U12581 (N_12581,N_12433,N_12358);
xnor U12582 (N_12582,N_12304,N_12394);
or U12583 (N_12583,N_12390,N_12303);
xor U12584 (N_12584,N_12378,N_12382);
or U12585 (N_12585,N_12444,N_12364);
nor U12586 (N_12586,N_12438,N_12335);
nand U12587 (N_12587,N_12313,N_12386);
nor U12588 (N_12588,N_12341,N_12447);
and U12589 (N_12589,N_12317,N_12308);
nor U12590 (N_12590,N_12300,N_12317);
xor U12591 (N_12591,N_12324,N_12408);
xor U12592 (N_12592,N_12433,N_12323);
and U12593 (N_12593,N_12362,N_12308);
or U12594 (N_12594,N_12406,N_12398);
and U12595 (N_12595,N_12444,N_12429);
nor U12596 (N_12596,N_12308,N_12445);
nor U12597 (N_12597,N_12413,N_12439);
nand U12598 (N_12598,N_12344,N_12309);
and U12599 (N_12599,N_12310,N_12430);
and U12600 (N_12600,N_12490,N_12549);
nor U12601 (N_12601,N_12530,N_12588);
nor U12602 (N_12602,N_12590,N_12454);
or U12603 (N_12603,N_12467,N_12583);
and U12604 (N_12604,N_12565,N_12513);
nand U12605 (N_12605,N_12533,N_12573);
and U12606 (N_12606,N_12586,N_12546);
xnor U12607 (N_12607,N_12507,N_12478);
and U12608 (N_12608,N_12482,N_12452);
xor U12609 (N_12609,N_12472,N_12563);
nand U12610 (N_12610,N_12574,N_12518);
or U12611 (N_12611,N_12468,N_12493);
and U12612 (N_12612,N_12496,N_12509);
nand U12613 (N_12613,N_12551,N_12593);
nand U12614 (N_12614,N_12587,N_12508);
nand U12615 (N_12615,N_12471,N_12599);
xor U12616 (N_12616,N_12477,N_12528);
xnor U12617 (N_12617,N_12475,N_12538);
nor U12618 (N_12618,N_12495,N_12519);
xor U12619 (N_12619,N_12480,N_12502);
nand U12620 (N_12620,N_12512,N_12517);
and U12621 (N_12621,N_12531,N_12559);
or U12622 (N_12622,N_12506,N_12459);
nor U12623 (N_12623,N_12575,N_12570);
nand U12624 (N_12624,N_12564,N_12532);
nor U12625 (N_12625,N_12579,N_12536);
xor U12626 (N_12626,N_12543,N_12534);
or U12627 (N_12627,N_12545,N_12527);
nand U12628 (N_12628,N_12469,N_12541);
xnor U12629 (N_12629,N_12465,N_12484);
xnor U12630 (N_12630,N_12515,N_12470);
or U12631 (N_12631,N_12466,N_12558);
nor U12632 (N_12632,N_12486,N_12456);
and U12633 (N_12633,N_12571,N_12594);
nor U12634 (N_12634,N_12492,N_12562);
nand U12635 (N_12635,N_12491,N_12554);
or U12636 (N_12636,N_12503,N_12557);
xnor U12637 (N_12637,N_12514,N_12487);
nand U12638 (N_12638,N_12483,N_12568);
nor U12639 (N_12639,N_12516,N_12537);
xor U12640 (N_12640,N_12455,N_12540);
nor U12641 (N_12641,N_12520,N_12453);
and U12642 (N_12642,N_12505,N_12524);
nor U12643 (N_12643,N_12462,N_12589);
xnor U12644 (N_12644,N_12548,N_12510);
xor U12645 (N_12645,N_12458,N_12522);
nand U12646 (N_12646,N_12498,N_12535);
or U12647 (N_12647,N_12578,N_12576);
or U12648 (N_12648,N_12485,N_12463);
nor U12649 (N_12649,N_12474,N_12553);
and U12650 (N_12650,N_12569,N_12499);
and U12651 (N_12651,N_12596,N_12523);
nand U12652 (N_12652,N_12566,N_12504);
nand U12653 (N_12653,N_12521,N_12460);
or U12654 (N_12654,N_12451,N_12584);
or U12655 (N_12655,N_12497,N_12598);
or U12656 (N_12656,N_12539,N_12556);
xor U12657 (N_12657,N_12547,N_12597);
or U12658 (N_12658,N_12581,N_12529);
nand U12659 (N_12659,N_12560,N_12595);
or U12660 (N_12660,N_12525,N_12591);
nor U12661 (N_12661,N_12582,N_12567);
or U12662 (N_12662,N_12473,N_12457);
nor U12663 (N_12663,N_12464,N_12511);
nand U12664 (N_12664,N_12481,N_12585);
nand U12665 (N_12665,N_12592,N_12550);
nand U12666 (N_12666,N_12476,N_12577);
and U12667 (N_12667,N_12494,N_12572);
nor U12668 (N_12668,N_12544,N_12552);
and U12669 (N_12669,N_12561,N_12488);
nand U12670 (N_12670,N_12479,N_12450);
nand U12671 (N_12671,N_12542,N_12580);
nand U12672 (N_12672,N_12555,N_12526);
nor U12673 (N_12673,N_12461,N_12501);
nor U12674 (N_12674,N_12489,N_12500);
or U12675 (N_12675,N_12450,N_12546);
or U12676 (N_12676,N_12570,N_12453);
and U12677 (N_12677,N_12593,N_12544);
xnor U12678 (N_12678,N_12563,N_12525);
or U12679 (N_12679,N_12464,N_12539);
xor U12680 (N_12680,N_12452,N_12479);
or U12681 (N_12681,N_12563,N_12505);
xnor U12682 (N_12682,N_12537,N_12475);
nand U12683 (N_12683,N_12469,N_12546);
nand U12684 (N_12684,N_12535,N_12551);
and U12685 (N_12685,N_12511,N_12548);
xor U12686 (N_12686,N_12520,N_12535);
nand U12687 (N_12687,N_12462,N_12511);
or U12688 (N_12688,N_12556,N_12586);
or U12689 (N_12689,N_12468,N_12471);
nand U12690 (N_12690,N_12533,N_12575);
or U12691 (N_12691,N_12503,N_12504);
nand U12692 (N_12692,N_12489,N_12521);
xnor U12693 (N_12693,N_12473,N_12471);
nor U12694 (N_12694,N_12544,N_12459);
and U12695 (N_12695,N_12459,N_12532);
and U12696 (N_12696,N_12552,N_12531);
xnor U12697 (N_12697,N_12568,N_12492);
xor U12698 (N_12698,N_12491,N_12548);
nor U12699 (N_12699,N_12472,N_12564);
or U12700 (N_12700,N_12552,N_12546);
xor U12701 (N_12701,N_12550,N_12533);
nor U12702 (N_12702,N_12462,N_12561);
xor U12703 (N_12703,N_12498,N_12450);
or U12704 (N_12704,N_12488,N_12493);
nor U12705 (N_12705,N_12479,N_12499);
or U12706 (N_12706,N_12588,N_12597);
or U12707 (N_12707,N_12532,N_12494);
nor U12708 (N_12708,N_12475,N_12550);
nor U12709 (N_12709,N_12471,N_12485);
xor U12710 (N_12710,N_12477,N_12582);
or U12711 (N_12711,N_12599,N_12575);
nor U12712 (N_12712,N_12570,N_12520);
and U12713 (N_12713,N_12460,N_12565);
nand U12714 (N_12714,N_12598,N_12533);
or U12715 (N_12715,N_12526,N_12530);
or U12716 (N_12716,N_12531,N_12483);
nand U12717 (N_12717,N_12543,N_12524);
nand U12718 (N_12718,N_12572,N_12585);
nand U12719 (N_12719,N_12483,N_12498);
nand U12720 (N_12720,N_12584,N_12564);
or U12721 (N_12721,N_12516,N_12508);
nor U12722 (N_12722,N_12480,N_12594);
or U12723 (N_12723,N_12451,N_12481);
nand U12724 (N_12724,N_12536,N_12508);
nand U12725 (N_12725,N_12517,N_12555);
nor U12726 (N_12726,N_12464,N_12570);
xor U12727 (N_12727,N_12517,N_12456);
and U12728 (N_12728,N_12497,N_12552);
or U12729 (N_12729,N_12589,N_12582);
xor U12730 (N_12730,N_12571,N_12451);
nor U12731 (N_12731,N_12518,N_12527);
or U12732 (N_12732,N_12546,N_12453);
and U12733 (N_12733,N_12456,N_12577);
and U12734 (N_12734,N_12466,N_12496);
or U12735 (N_12735,N_12593,N_12453);
or U12736 (N_12736,N_12560,N_12593);
and U12737 (N_12737,N_12474,N_12536);
nor U12738 (N_12738,N_12538,N_12565);
or U12739 (N_12739,N_12549,N_12539);
nand U12740 (N_12740,N_12598,N_12557);
or U12741 (N_12741,N_12545,N_12520);
nor U12742 (N_12742,N_12468,N_12512);
nand U12743 (N_12743,N_12571,N_12578);
nor U12744 (N_12744,N_12522,N_12461);
or U12745 (N_12745,N_12566,N_12547);
nor U12746 (N_12746,N_12505,N_12480);
nand U12747 (N_12747,N_12453,N_12541);
or U12748 (N_12748,N_12592,N_12464);
or U12749 (N_12749,N_12535,N_12481);
and U12750 (N_12750,N_12651,N_12614);
nand U12751 (N_12751,N_12600,N_12626);
nor U12752 (N_12752,N_12641,N_12678);
and U12753 (N_12753,N_12701,N_12681);
nand U12754 (N_12754,N_12686,N_12741);
and U12755 (N_12755,N_12687,N_12718);
and U12756 (N_12756,N_12663,N_12668);
nor U12757 (N_12757,N_12624,N_12609);
or U12758 (N_12758,N_12698,N_12731);
nand U12759 (N_12759,N_12722,N_12732);
and U12760 (N_12760,N_12610,N_12738);
nor U12761 (N_12761,N_12720,N_12700);
and U12762 (N_12762,N_12690,N_12608);
nand U12763 (N_12763,N_12664,N_12615);
nand U12764 (N_12764,N_12719,N_12693);
nand U12765 (N_12765,N_12637,N_12653);
and U12766 (N_12766,N_12642,N_12748);
xnor U12767 (N_12767,N_12747,N_12714);
nor U12768 (N_12768,N_12625,N_12733);
or U12769 (N_12769,N_12697,N_12666);
nand U12770 (N_12770,N_12650,N_12679);
or U12771 (N_12771,N_12671,N_12665);
nor U12772 (N_12772,N_12640,N_12737);
nor U12773 (N_12773,N_12727,N_12716);
nor U12774 (N_12774,N_12601,N_12611);
nand U12775 (N_12775,N_12672,N_12736);
and U12776 (N_12776,N_12675,N_12696);
nor U12777 (N_12777,N_12724,N_12646);
nor U12778 (N_12778,N_12649,N_12746);
nor U12779 (N_12779,N_12629,N_12618);
or U12780 (N_12780,N_12702,N_12677);
and U12781 (N_12781,N_12710,N_12689);
or U12782 (N_12782,N_12743,N_12669);
nand U12783 (N_12783,N_12656,N_12706);
nand U12784 (N_12784,N_12670,N_12606);
or U12785 (N_12785,N_12632,N_12667);
xor U12786 (N_12786,N_12729,N_12734);
and U12787 (N_12787,N_12692,N_12707);
xor U12788 (N_12788,N_12717,N_12728);
and U12789 (N_12789,N_12683,N_12634);
nand U12790 (N_12790,N_12682,N_12648);
or U12791 (N_12791,N_12631,N_12703);
nor U12792 (N_12792,N_12725,N_12705);
or U12793 (N_12793,N_12605,N_12622);
and U12794 (N_12794,N_12709,N_12712);
nand U12795 (N_12795,N_12699,N_12645);
xor U12796 (N_12796,N_12744,N_12691);
nor U12797 (N_12797,N_12704,N_12654);
xnor U12798 (N_12798,N_12643,N_12715);
nand U12799 (N_12799,N_12620,N_12658);
or U12800 (N_12800,N_12708,N_12730);
or U12801 (N_12801,N_12613,N_12742);
or U12802 (N_12802,N_12635,N_12657);
nor U12803 (N_12803,N_12673,N_12740);
xor U12804 (N_12804,N_12726,N_12662);
and U12805 (N_12805,N_12694,N_12711);
nor U12806 (N_12806,N_12603,N_12655);
or U12807 (N_12807,N_12749,N_12627);
nand U12808 (N_12808,N_12723,N_12688);
nor U12809 (N_12809,N_12684,N_12607);
or U12810 (N_12810,N_12713,N_12604);
nand U12811 (N_12811,N_12638,N_12633);
xor U12812 (N_12812,N_12636,N_12695);
or U12813 (N_12813,N_12674,N_12647);
nand U12814 (N_12814,N_12660,N_12652);
and U12815 (N_12815,N_12745,N_12621);
or U12816 (N_12816,N_12602,N_12680);
and U12817 (N_12817,N_12676,N_12612);
or U12818 (N_12818,N_12628,N_12659);
or U12819 (N_12819,N_12644,N_12721);
nand U12820 (N_12820,N_12623,N_12616);
and U12821 (N_12821,N_12630,N_12661);
and U12822 (N_12822,N_12619,N_12639);
xor U12823 (N_12823,N_12617,N_12685);
xor U12824 (N_12824,N_12735,N_12739);
nor U12825 (N_12825,N_12668,N_12644);
nor U12826 (N_12826,N_12664,N_12629);
nand U12827 (N_12827,N_12706,N_12712);
nand U12828 (N_12828,N_12651,N_12654);
nor U12829 (N_12829,N_12655,N_12719);
nand U12830 (N_12830,N_12630,N_12604);
or U12831 (N_12831,N_12683,N_12653);
nand U12832 (N_12832,N_12734,N_12741);
nor U12833 (N_12833,N_12714,N_12657);
or U12834 (N_12834,N_12688,N_12629);
and U12835 (N_12835,N_12699,N_12716);
or U12836 (N_12836,N_12606,N_12609);
xnor U12837 (N_12837,N_12687,N_12631);
nor U12838 (N_12838,N_12657,N_12666);
nand U12839 (N_12839,N_12704,N_12720);
or U12840 (N_12840,N_12652,N_12703);
xnor U12841 (N_12841,N_12604,N_12727);
nand U12842 (N_12842,N_12678,N_12723);
nor U12843 (N_12843,N_12637,N_12729);
nor U12844 (N_12844,N_12629,N_12748);
nand U12845 (N_12845,N_12695,N_12647);
and U12846 (N_12846,N_12629,N_12609);
nand U12847 (N_12847,N_12600,N_12732);
or U12848 (N_12848,N_12719,N_12695);
and U12849 (N_12849,N_12664,N_12705);
xnor U12850 (N_12850,N_12707,N_12629);
nor U12851 (N_12851,N_12748,N_12728);
xor U12852 (N_12852,N_12722,N_12644);
nor U12853 (N_12853,N_12704,N_12743);
nand U12854 (N_12854,N_12664,N_12741);
nor U12855 (N_12855,N_12682,N_12675);
nor U12856 (N_12856,N_12724,N_12613);
and U12857 (N_12857,N_12679,N_12725);
nand U12858 (N_12858,N_12607,N_12644);
nor U12859 (N_12859,N_12697,N_12707);
and U12860 (N_12860,N_12678,N_12727);
nand U12861 (N_12861,N_12618,N_12660);
or U12862 (N_12862,N_12697,N_12619);
nand U12863 (N_12863,N_12615,N_12688);
xnor U12864 (N_12864,N_12631,N_12629);
xnor U12865 (N_12865,N_12647,N_12663);
nor U12866 (N_12866,N_12612,N_12640);
nand U12867 (N_12867,N_12655,N_12666);
or U12868 (N_12868,N_12719,N_12706);
nand U12869 (N_12869,N_12691,N_12683);
nand U12870 (N_12870,N_12619,N_12721);
and U12871 (N_12871,N_12616,N_12685);
and U12872 (N_12872,N_12658,N_12661);
or U12873 (N_12873,N_12614,N_12649);
nand U12874 (N_12874,N_12665,N_12716);
or U12875 (N_12875,N_12669,N_12657);
nor U12876 (N_12876,N_12645,N_12625);
nor U12877 (N_12877,N_12738,N_12732);
xor U12878 (N_12878,N_12746,N_12659);
xor U12879 (N_12879,N_12680,N_12729);
xnor U12880 (N_12880,N_12687,N_12640);
nor U12881 (N_12881,N_12712,N_12654);
and U12882 (N_12882,N_12745,N_12626);
and U12883 (N_12883,N_12700,N_12703);
xnor U12884 (N_12884,N_12703,N_12725);
nand U12885 (N_12885,N_12613,N_12643);
xor U12886 (N_12886,N_12718,N_12626);
nand U12887 (N_12887,N_12685,N_12703);
xor U12888 (N_12888,N_12631,N_12654);
nor U12889 (N_12889,N_12660,N_12713);
xnor U12890 (N_12890,N_12748,N_12700);
and U12891 (N_12891,N_12636,N_12728);
and U12892 (N_12892,N_12625,N_12726);
xnor U12893 (N_12893,N_12698,N_12632);
or U12894 (N_12894,N_12700,N_12744);
or U12895 (N_12895,N_12742,N_12655);
nor U12896 (N_12896,N_12743,N_12637);
nor U12897 (N_12897,N_12729,N_12737);
nand U12898 (N_12898,N_12644,N_12684);
and U12899 (N_12899,N_12637,N_12718);
xor U12900 (N_12900,N_12752,N_12849);
nor U12901 (N_12901,N_12855,N_12838);
nor U12902 (N_12902,N_12879,N_12872);
nand U12903 (N_12903,N_12788,N_12794);
nor U12904 (N_12904,N_12889,N_12813);
nand U12905 (N_12905,N_12759,N_12899);
xor U12906 (N_12906,N_12777,N_12831);
xnor U12907 (N_12907,N_12754,N_12875);
nor U12908 (N_12908,N_12793,N_12874);
nand U12909 (N_12909,N_12764,N_12823);
nor U12910 (N_12910,N_12857,N_12871);
and U12911 (N_12911,N_12837,N_12828);
and U12912 (N_12912,N_12807,N_12882);
or U12913 (N_12913,N_12842,N_12783);
nand U12914 (N_12914,N_12843,N_12888);
nand U12915 (N_12915,N_12845,N_12775);
or U12916 (N_12916,N_12852,N_12760);
xor U12917 (N_12917,N_12817,N_12799);
and U12918 (N_12918,N_12846,N_12892);
and U12919 (N_12919,N_12771,N_12804);
nand U12920 (N_12920,N_12755,N_12766);
nor U12921 (N_12921,N_12770,N_12840);
or U12922 (N_12922,N_12769,N_12854);
nand U12923 (N_12923,N_12792,N_12824);
xor U12924 (N_12924,N_12853,N_12781);
and U12925 (N_12925,N_12765,N_12819);
nand U12926 (N_12926,N_12833,N_12774);
and U12927 (N_12927,N_12863,N_12779);
nor U12928 (N_12928,N_12885,N_12841);
nand U12929 (N_12929,N_12773,N_12812);
nand U12930 (N_12930,N_12876,N_12758);
nor U12931 (N_12931,N_12822,N_12891);
nor U12932 (N_12932,N_12866,N_12784);
xor U12933 (N_12933,N_12862,N_12851);
xor U12934 (N_12934,N_12751,N_12801);
nand U12935 (N_12935,N_12815,N_12830);
and U12936 (N_12936,N_12761,N_12878);
xnor U12937 (N_12937,N_12894,N_12798);
nor U12938 (N_12938,N_12893,N_12811);
nor U12939 (N_12939,N_12767,N_12895);
nand U12940 (N_12940,N_12836,N_12847);
nor U12941 (N_12941,N_12825,N_12756);
or U12942 (N_12942,N_12797,N_12826);
xor U12943 (N_12943,N_12776,N_12860);
and U12944 (N_12944,N_12757,N_12821);
and U12945 (N_12945,N_12805,N_12835);
xor U12946 (N_12946,N_12818,N_12896);
nand U12947 (N_12947,N_12834,N_12763);
xor U12948 (N_12948,N_12787,N_12865);
nand U12949 (N_12949,N_12810,N_12806);
nand U12950 (N_12950,N_12795,N_12869);
or U12951 (N_12951,N_12802,N_12832);
and U12952 (N_12952,N_12861,N_12864);
nand U12953 (N_12953,N_12753,N_12844);
nor U12954 (N_12954,N_12814,N_12803);
xnor U12955 (N_12955,N_12850,N_12877);
xnor U12956 (N_12956,N_12897,N_12829);
or U12957 (N_12957,N_12800,N_12782);
nand U12958 (N_12958,N_12886,N_12808);
or U12959 (N_12959,N_12750,N_12791);
xor U12960 (N_12960,N_12898,N_12839);
nor U12961 (N_12961,N_12789,N_12827);
and U12962 (N_12962,N_12816,N_12867);
nand U12963 (N_12963,N_12762,N_12848);
nand U12964 (N_12964,N_12887,N_12778);
or U12965 (N_12965,N_12880,N_12884);
nand U12966 (N_12966,N_12768,N_12881);
nand U12967 (N_12967,N_12786,N_12883);
xnor U12968 (N_12968,N_12859,N_12772);
and U12969 (N_12969,N_12890,N_12785);
and U12970 (N_12970,N_12870,N_12856);
xnor U12971 (N_12971,N_12809,N_12780);
nand U12972 (N_12972,N_12820,N_12796);
or U12973 (N_12973,N_12868,N_12873);
or U12974 (N_12974,N_12790,N_12858);
xnor U12975 (N_12975,N_12781,N_12879);
and U12976 (N_12976,N_12761,N_12791);
xor U12977 (N_12977,N_12805,N_12847);
xnor U12978 (N_12978,N_12894,N_12828);
nand U12979 (N_12979,N_12885,N_12751);
xor U12980 (N_12980,N_12858,N_12880);
xor U12981 (N_12981,N_12863,N_12833);
nand U12982 (N_12982,N_12856,N_12750);
and U12983 (N_12983,N_12888,N_12831);
nand U12984 (N_12984,N_12889,N_12839);
and U12985 (N_12985,N_12810,N_12754);
xor U12986 (N_12986,N_12789,N_12791);
and U12987 (N_12987,N_12820,N_12765);
nand U12988 (N_12988,N_12759,N_12847);
or U12989 (N_12989,N_12779,N_12844);
nand U12990 (N_12990,N_12817,N_12829);
nor U12991 (N_12991,N_12812,N_12844);
or U12992 (N_12992,N_12787,N_12780);
xor U12993 (N_12993,N_12869,N_12870);
or U12994 (N_12994,N_12788,N_12829);
and U12995 (N_12995,N_12795,N_12803);
xor U12996 (N_12996,N_12855,N_12863);
nand U12997 (N_12997,N_12826,N_12819);
nand U12998 (N_12998,N_12827,N_12791);
xnor U12999 (N_12999,N_12874,N_12813);
nand U13000 (N_13000,N_12792,N_12814);
xor U13001 (N_13001,N_12855,N_12798);
nand U13002 (N_13002,N_12887,N_12867);
and U13003 (N_13003,N_12870,N_12783);
or U13004 (N_13004,N_12761,N_12866);
nor U13005 (N_13005,N_12876,N_12873);
nand U13006 (N_13006,N_12860,N_12893);
or U13007 (N_13007,N_12845,N_12832);
and U13008 (N_13008,N_12869,N_12863);
nand U13009 (N_13009,N_12763,N_12851);
nand U13010 (N_13010,N_12779,N_12751);
nor U13011 (N_13011,N_12831,N_12790);
xnor U13012 (N_13012,N_12796,N_12804);
nor U13013 (N_13013,N_12782,N_12855);
xor U13014 (N_13014,N_12772,N_12865);
nor U13015 (N_13015,N_12890,N_12789);
or U13016 (N_13016,N_12798,N_12763);
nand U13017 (N_13017,N_12761,N_12788);
or U13018 (N_13018,N_12792,N_12806);
nand U13019 (N_13019,N_12856,N_12763);
and U13020 (N_13020,N_12865,N_12806);
xor U13021 (N_13021,N_12807,N_12795);
nand U13022 (N_13022,N_12784,N_12877);
xnor U13023 (N_13023,N_12816,N_12829);
nand U13024 (N_13024,N_12841,N_12803);
or U13025 (N_13025,N_12787,N_12818);
or U13026 (N_13026,N_12892,N_12859);
xor U13027 (N_13027,N_12847,N_12866);
or U13028 (N_13028,N_12810,N_12751);
nand U13029 (N_13029,N_12793,N_12870);
or U13030 (N_13030,N_12760,N_12835);
xnor U13031 (N_13031,N_12760,N_12891);
nor U13032 (N_13032,N_12817,N_12830);
xnor U13033 (N_13033,N_12842,N_12790);
nand U13034 (N_13034,N_12775,N_12817);
nor U13035 (N_13035,N_12824,N_12799);
nand U13036 (N_13036,N_12898,N_12855);
xnor U13037 (N_13037,N_12809,N_12755);
nand U13038 (N_13038,N_12869,N_12785);
or U13039 (N_13039,N_12855,N_12752);
and U13040 (N_13040,N_12763,N_12760);
xnor U13041 (N_13041,N_12829,N_12753);
xor U13042 (N_13042,N_12896,N_12893);
or U13043 (N_13043,N_12780,N_12864);
or U13044 (N_13044,N_12847,N_12799);
or U13045 (N_13045,N_12838,N_12845);
nor U13046 (N_13046,N_12875,N_12815);
xnor U13047 (N_13047,N_12881,N_12889);
xor U13048 (N_13048,N_12760,N_12880);
nor U13049 (N_13049,N_12799,N_12831);
nor U13050 (N_13050,N_13041,N_13046);
xor U13051 (N_13051,N_12902,N_13028);
xnor U13052 (N_13052,N_13044,N_12919);
and U13053 (N_13053,N_12959,N_13007);
xor U13054 (N_13054,N_12917,N_12952);
or U13055 (N_13055,N_12996,N_13021);
nand U13056 (N_13056,N_12965,N_13033);
xnor U13057 (N_13057,N_13038,N_13029);
nor U13058 (N_13058,N_12903,N_13030);
nor U13059 (N_13059,N_12920,N_12934);
nor U13060 (N_13060,N_13001,N_12945);
xor U13061 (N_13061,N_13003,N_12936);
and U13062 (N_13062,N_12933,N_12915);
and U13063 (N_13063,N_13039,N_12947);
or U13064 (N_13064,N_12982,N_13002);
nor U13065 (N_13065,N_12943,N_12979);
nand U13066 (N_13066,N_12997,N_13031);
and U13067 (N_13067,N_12985,N_13006);
nand U13068 (N_13068,N_12928,N_13022);
xor U13069 (N_13069,N_13043,N_12984);
xnor U13070 (N_13070,N_13012,N_12932);
or U13071 (N_13071,N_13035,N_12904);
and U13072 (N_13072,N_13015,N_12922);
nand U13073 (N_13073,N_13017,N_12901);
and U13074 (N_13074,N_12916,N_12925);
and U13075 (N_13075,N_12998,N_12910);
xor U13076 (N_13076,N_12908,N_12968);
and U13077 (N_13077,N_12948,N_13014);
xor U13078 (N_13078,N_12963,N_12973);
or U13079 (N_13079,N_12927,N_12909);
xor U13080 (N_13080,N_13024,N_12921);
nor U13081 (N_13081,N_12977,N_12969);
nor U13082 (N_13082,N_12992,N_12914);
nor U13083 (N_13083,N_13013,N_13008);
nor U13084 (N_13084,N_12995,N_12980);
nand U13085 (N_13085,N_12930,N_12967);
nand U13086 (N_13086,N_13020,N_13040);
and U13087 (N_13087,N_12949,N_12993);
or U13088 (N_13088,N_12962,N_12974);
and U13089 (N_13089,N_12960,N_12940);
nand U13090 (N_13090,N_13049,N_12913);
nand U13091 (N_13091,N_13000,N_13025);
xnor U13092 (N_13092,N_12924,N_12971);
nand U13093 (N_13093,N_13036,N_13042);
xnor U13094 (N_13094,N_12983,N_12907);
xor U13095 (N_13095,N_13047,N_12944);
and U13096 (N_13096,N_13034,N_12938);
nand U13097 (N_13097,N_12961,N_12956);
xnor U13098 (N_13098,N_13009,N_12990);
xnor U13099 (N_13099,N_12978,N_13019);
or U13100 (N_13100,N_12951,N_12900);
nand U13101 (N_13101,N_13037,N_12941);
nand U13102 (N_13102,N_12970,N_12999);
nand U13103 (N_13103,N_12929,N_12926);
xor U13104 (N_13104,N_12955,N_13016);
and U13105 (N_13105,N_12964,N_12911);
nand U13106 (N_13106,N_12937,N_13032);
nor U13107 (N_13107,N_13026,N_13018);
nor U13108 (N_13108,N_12975,N_12958);
and U13109 (N_13109,N_12939,N_12946);
xnor U13110 (N_13110,N_12953,N_12981);
nand U13111 (N_13111,N_13045,N_12906);
or U13112 (N_13112,N_12954,N_12923);
or U13113 (N_13113,N_12987,N_13023);
xnor U13114 (N_13114,N_12966,N_12976);
xor U13115 (N_13115,N_12912,N_12950);
nor U13116 (N_13116,N_12972,N_12957);
nand U13117 (N_13117,N_13011,N_12994);
xor U13118 (N_13118,N_12942,N_12988);
or U13119 (N_13119,N_12991,N_12918);
xor U13120 (N_13120,N_12931,N_13004);
nand U13121 (N_13121,N_12989,N_13027);
nand U13122 (N_13122,N_12905,N_12986);
xor U13123 (N_13123,N_13048,N_12935);
nor U13124 (N_13124,N_13005,N_13010);
xor U13125 (N_13125,N_12911,N_12930);
xor U13126 (N_13126,N_12965,N_12991);
or U13127 (N_13127,N_12904,N_12945);
nor U13128 (N_13128,N_13007,N_13024);
and U13129 (N_13129,N_12979,N_12957);
xnor U13130 (N_13130,N_12985,N_12987);
nand U13131 (N_13131,N_12934,N_13027);
or U13132 (N_13132,N_12923,N_13011);
or U13133 (N_13133,N_13015,N_13019);
and U13134 (N_13134,N_13014,N_12976);
xnor U13135 (N_13135,N_12909,N_13034);
and U13136 (N_13136,N_13007,N_12942);
nor U13137 (N_13137,N_12930,N_13003);
and U13138 (N_13138,N_13027,N_12947);
nand U13139 (N_13139,N_12914,N_13012);
xor U13140 (N_13140,N_12959,N_12958);
nand U13141 (N_13141,N_12993,N_13035);
xnor U13142 (N_13142,N_12995,N_13043);
or U13143 (N_13143,N_12938,N_13008);
and U13144 (N_13144,N_13012,N_13014);
or U13145 (N_13145,N_12980,N_12988);
nor U13146 (N_13146,N_13009,N_13044);
and U13147 (N_13147,N_12940,N_12923);
nand U13148 (N_13148,N_12969,N_13033);
xor U13149 (N_13149,N_12975,N_13004);
nor U13150 (N_13150,N_12904,N_12998);
nand U13151 (N_13151,N_12972,N_13034);
nor U13152 (N_13152,N_13024,N_12901);
nor U13153 (N_13153,N_12943,N_12928);
and U13154 (N_13154,N_13032,N_12974);
nand U13155 (N_13155,N_12953,N_12915);
and U13156 (N_13156,N_13006,N_12960);
or U13157 (N_13157,N_13048,N_13030);
nand U13158 (N_13158,N_12988,N_12957);
xor U13159 (N_13159,N_13030,N_13031);
xnor U13160 (N_13160,N_13006,N_13015);
nand U13161 (N_13161,N_12932,N_12994);
nand U13162 (N_13162,N_13010,N_12989);
and U13163 (N_13163,N_13005,N_12984);
and U13164 (N_13164,N_12956,N_13019);
xor U13165 (N_13165,N_12945,N_13045);
nand U13166 (N_13166,N_13023,N_12969);
or U13167 (N_13167,N_12956,N_12930);
nand U13168 (N_13168,N_12913,N_13028);
nand U13169 (N_13169,N_12926,N_12912);
or U13170 (N_13170,N_13016,N_12999);
or U13171 (N_13171,N_12996,N_13018);
nand U13172 (N_13172,N_12999,N_13018);
or U13173 (N_13173,N_12996,N_13012);
nor U13174 (N_13174,N_13046,N_12980);
nand U13175 (N_13175,N_12994,N_12937);
nor U13176 (N_13176,N_12950,N_13025);
nor U13177 (N_13177,N_12968,N_13010);
xor U13178 (N_13178,N_12919,N_13010);
and U13179 (N_13179,N_13046,N_12922);
or U13180 (N_13180,N_12964,N_12949);
and U13181 (N_13181,N_13044,N_13018);
or U13182 (N_13182,N_13013,N_12942);
nor U13183 (N_13183,N_12937,N_12950);
and U13184 (N_13184,N_12971,N_13011);
xnor U13185 (N_13185,N_12963,N_13024);
or U13186 (N_13186,N_12985,N_13029);
nand U13187 (N_13187,N_12925,N_13018);
and U13188 (N_13188,N_12906,N_12941);
nor U13189 (N_13189,N_12998,N_12905);
nand U13190 (N_13190,N_12989,N_12948);
nand U13191 (N_13191,N_13030,N_12980);
and U13192 (N_13192,N_12903,N_12996);
nand U13193 (N_13193,N_12928,N_13012);
nor U13194 (N_13194,N_12939,N_13047);
and U13195 (N_13195,N_12999,N_13024);
nand U13196 (N_13196,N_12994,N_12969);
nand U13197 (N_13197,N_12916,N_12922);
nand U13198 (N_13198,N_12967,N_12981);
nand U13199 (N_13199,N_12934,N_13028);
and U13200 (N_13200,N_13153,N_13096);
xor U13201 (N_13201,N_13099,N_13148);
xnor U13202 (N_13202,N_13063,N_13141);
nor U13203 (N_13203,N_13056,N_13081);
nor U13204 (N_13204,N_13164,N_13117);
or U13205 (N_13205,N_13109,N_13107);
nor U13206 (N_13206,N_13089,N_13119);
nor U13207 (N_13207,N_13080,N_13131);
xnor U13208 (N_13208,N_13095,N_13177);
and U13209 (N_13209,N_13124,N_13171);
nand U13210 (N_13210,N_13083,N_13086);
or U13211 (N_13211,N_13197,N_13151);
or U13212 (N_13212,N_13174,N_13175);
nand U13213 (N_13213,N_13192,N_13051);
or U13214 (N_13214,N_13184,N_13157);
xor U13215 (N_13215,N_13140,N_13193);
nand U13216 (N_13216,N_13071,N_13159);
xor U13217 (N_13217,N_13058,N_13191);
nand U13218 (N_13218,N_13134,N_13070);
nor U13219 (N_13219,N_13093,N_13129);
or U13220 (N_13220,N_13092,N_13108);
or U13221 (N_13221,N_13150,N_13160);
nand U13222 (N_13222,N_13116,N_13061);
nor U13223 (N_13223,N_13106,N_13054);
nand U13224 (N_13224,N_13183,N_13069);
nand U13225 (N_13225,N_13082,N_13180);
nand U13226 (N_13226,N_13172,N_13123);
or U13227 (N_13227,N_13078,N_13102);
or U13228 (N_13228,N_13179,N_13156);
nor U13229 (N_13229,N_13166,N_13052);
or U13230 (N_13230,N_13103,N_13186);
nor U13231 (N_13231,N_13143,N_13162);
nor U13232 (N_13232,N_13077,N_13145);
and U13233 (N_13233,N_13087,N_13152);
nand U13234 (N_13234,N_13115,N_13199);
xnor U13235 (N_13235,N_13084,N_13062);
nor U13236 (N_13236,N_13074,N_13176);
and U13237 (N_13237,N_13125,N_13079);
xor U13238 (N_13238,N_13154,N_13101);
nor U13239 (N_13239,N_13068,N_13196);
xor U13240 (N_13240,N_13060,N_13163);
nor U13241 (N_13241,N_13149,N_13121);
and U13242 (N_13242,N_13178,N_13118);
or U13243 (N_13243,N_13059,N_13127);
nor U13244 (N_13244,N_13188,N_13100);
or U13245 (N_13245,N_13050,N_13146);
or U13246 (N_13246,N_13073,N_13128);
xnor U13247 (N_13247,N_13057,N_13189);
nor U13248 (N_13248,N_13190,N_13168);
or U13249 (N_13249,N_13198,N_13185);
nor U13250 (N_13250,N_13097,N_13122);
nand U13251 (N_13251,N_13133,N_13169);
nor U13252 (N_13252,N_13142,N_13147);
or U13253 (N_13253,N_13161,N_13085);
xor U13254 (N_13254,N_13098,N_13053);
and U13255 (N_13255,N_13111,N_13072);
xor U13256 (N_13256,N_13165,N_13167);
xor U13257 (N_13257,N_13130,N_13076);
or U13258 (N_13258,N_13170,N_13126);
nand U13259 (N_13259,N_13067,N_13112);
xnor U13260 (N_13260,N_13158,N_13105);
nand U13261 (N_13261,N_13137,N_13094);
nor U13262 (N_13262,N_13055,N_13135);
or U13263 (N_13263,N_13136,N_13066);
xor U13264 (N_13264,N_13187,N_13088);
nor U13265 (N_13265,N_13173,N_13155);
or U13266 (N_13266,N_13064,N_13132);
xor U13267 (N_13267,N_13195,N_13113);
and U13268 (N_13268,N_13120,N_13194);
xor U13269 (N_13269,N_13075,N_13181);
and U13270 (N_13270,N_13139,N_13138);
nor U13271 (N_13271,N_13090,N_13110);
and U13272 (N_13272,N_13104,N_13144);
nor U13273 (N_13273,N_13065,N_13091);
xnor U13274 (N_13274,N_13114,N_13182);
nor U13275 (N_13275,N_13143,N_13130);
and U13276 (N_13276,N_13114,N_13147);
or U13277 (N_13277,N_13111,N_13162);
xor U13278 (N_13278,N_13199,N_13062);
and U13279 (N_13279,N_13190,N_13179);
nand U13280 (N_13280,N_13195,N_13188);
or U13281 (N_13281,N_13153,N_13144);
or U13282 (N_13282,N_13065,N_13113);
and U13283 (N_13283,N_13170,N_13143);
nand U13284 (N_13284,N_13138,N_13061);
and U13285 (N_13285,N_13183,N_13087);
and U13286 (N_13286,N_13180,N_13133);
and U13287 (N_13287,N_13112,N_13084);
nor U13288 (N_13288,N_13108,N_13174);
nand U13289 (N_13289,N_13072,N_13196);
or U13290 (N_13290,N_13172,N_13148);
xnor U13291 (N_13291,N_13093,N_13100);
nand U13292 (N_13292,N_13190,N_13196);
and U13293 (N_13293,N_13174,N_13173);
and U13294 (N_13294,N_13089,N_13110);
or U13295 (N_13295,N_13133,N_13065);
xor U13296 (N_13296,N_13187,N_13116);
nand U13297 (N_13297,N_13176,N_13077);
nand U13298 (N_13298,N_13087,N_13158);
xor U13299 (N_13299,N_13167,N_13151);
nand U13300 (N_13300,N_13107,N_13128);
and U13301 (N_13301,N_13081,N_13125);
nand U13302 (N_13302,N_13157,N_13179);
nor U13303 (N_13303,N_13058,N_13069);
and U13304 (N_13304,N_13197,N_13053);
and U13305 (N_13305,N_13093,N_13124);
or U13306 (N_13306,N_13195,N_13154);
or U13307 (N_13307,N_13161,N_13147);
or U13308 (N_13308,N_13154,N_13078);
nor U13309 (N_13309,N_13124,N_13098);
nand U13310 (N_13310,N_13178,N_13198);
or U13311 (N_13311,N_13159,N_13055);
or U13312 (N_13312,N_13134,N_13068);
nand U13313 (N_13313,N_13055,N_13161);
nand U13314 (N_13314,N_13130,N_13074);
nor U13315 (N_13315,N_13058,N_13169);
or U13316 (N_13316,N_13177,N_13168);
nor U13317 (N_13317,N_13108,N_13180);
nor U13318 (N_13318,N_13091,N_13188);
nand U13319 (N_13319,N_13142,N_13103);
and U13320 (N_13320,N_13108,N_13065);
nor U13321 (N_13321,N_13138,N_13164);
nand U13322 (N_13322,N_13098,N_13086);
nand U13323 (N_13323,N_13094,N_13098);
xnor U13324 (N_13324,N_13152,N_13150);
or U13325 (N_13325,N_13097,N_13157);
or U13326 (N_13326,N_13151,N_13053);
or U13327 (N_13327,N_13067,N_13103);
nor U13328 (N_13328,N_13190,N_13063);
nand U13329 (N_13329,N_13088,N_13069);
nand U13330 (N_13330,N_13128,N_13079);
nand U13331 (N_13331,N_13191,N_13074);
or U13332 (N_13332,N_13100,N_13129);
and U13333 (N_13333,N_13081,N_13180);
xor U13334 (N_13334,N_13078,N_13187);
or U13335 (N_13335,N_13174,N_13086);
and U13336 (N_13336,N_13195,N_13132);
nand U13337 (N_13337,N_13053,N_13071);
xnor U13338 (N_13338,N_13164,N_13110);
xor U13339 (N_13339,N_13108,N_13133);
nand U13340 (N_13340,N_13076,N_13191);
xor U13341 (N_13341,N_13124,N_13103);
nor U13342 (N_13342,N_13123,N_13076);
or U13343 (N_13343,N_13193,N_13177);
nor U13344 (N_13344,N_13164,N_13120);
nand U13345 (N_13345,N_13087,N_13080);
or U13346 (N_13346,N_13157,N_13158);
and U13347 (N_13347,N_13137,N_13102);
nor U13348 (N_13348,N_13073,N_13170);
xnor U13349 (N_13349,N_13188,N_13124);
nand U13350 (N_13350,N_13285,N_13338);
xor U13351 (N_13351,N_13204,N_13302);
or U13352 (N_13352,N_13321,N_13274);
and U13353 (N_13353,N_13300,N_13288);
nor U13354 (N_13354,N_13268,N_13296);
nand U13355 (N_13355,N_13335,N_13346);
or U13356 (N_13356,N_13243,N_13254);
and U13357 (N_13357,N_13250,N_13205);
nand U13358 (N_13358,N_13322,N_13290);
nand U13359 (N_13359,N_13269,N_13291);
or U13360 (N_13360,N_13241,N_13212);
and U13361 (N_13361,N_13245,N_13294);
and U13362 (N_13362,N_13329,N_13292);
nor U13363 (N_13363,N_13202,N_13343);
and U13364 (N_13364,N_13234,N_13267);
and U13365 (N_13365,N_13320,N_13281);
nor U13366 (N_13366,N_13217,N_13242);
xor U13367 (N_13367,N_13210,N_13272);
nor U13368 (N_13368,N_13298,N_13216);
xor U13369 (N_13369,N_13283,N_13264);
xor U13370 (N_13370,N_13276,N_13328);
xnor U13371 (N_13371,N_13271,N_13253);
or U13372 (N_13372,N_13209,N_13327);
or U13373 (N_13373,N_13293,N_13229);
xnor U13374 (N_13374,N_13223,N_13227);
or U13375 (N_13375,N_13230,N_13336);
nor U13376 (N_13376,N_13219,N_13330);
xnor U13377 (N_13377,N_13236,N_13248);
and U13378 (N_13378,N_13282,N_13333);
or U13379 (N_13379,N_13239,N_13326);
or U13380 (N_13380,N_13307,N_13317);
nand U13381 (N_13381,N_13309,N_13306);
nor U13382 (N_13382,N_13332,N_13228);
and U13383 (N_13383,N_13237,N_13313);
nand U13384 (N_13384,N_13339,N_13257);
nand U13385 (N_13385,N_13232,N_13265);
nor U13386 (N_13386,N_13235,N_13231);
nand U13387 (N_13387,N_13258,N_13214);
nor U13388 (N_13388,N_13225,N_13246);
xnor U13389 (N_13389,N_13251,N_13284);
or U13390 (N_13390,N_13348,N_13287);
xor U13391 (N_13391,N_13266,N_13295);
xnor U13392 (N_13392,N_13224,N_13261);
nor U13393 (N_13393,N_13203,N_13319);
nor U13394 (N_13394,N_13303,N_13263);
and U13395 (N_13395,N_13256,N_13344);
nor U13396 (N_13396,N_13218,N_13340);
and U13397 (N_13397,N_13222,N_13308);
nor U13398 (N_13398,N_13315,N_13255);
nand U13399 (N_13399,N_13200,N_13349);
or U13400 (N_13400,N_13277,N_13238);
or U13401 (N_13401,N_13312,N_13305);
and U13402 (N_13402,N_13337,N_13334);
xnor U13403 (N_13403,N_13259,N_13342);
or U13404 (N_13404,N_13310,N_13299);
or U13405 (N_13405,N_13341,N_13221);
nor U13406 (N_13406,N_13220,N_13247);
xor U13407 (N_13407,N_13297,N_13301);
xnor U13408 (N_13408,N_13304,N_13260);
or U13409 (N_13409,N_13275,N_13273);
or U13410 (N_13410,N_13279,N_13215);
or U13411 (N_13411,N_13249,N_13201);
and U13412 (N_13412,N_13345,N_13280);
or U13413 (N_13413,N_13318,N_13325);
nor U13414 (N_13414,N_13252,N_13211);
or U13415 (N_13415,N_13208,N_13226);
and U13416 (N_13416,N_13316,N_13207);
or U13417 (N_13417,N_13323,N_13262);
xnor U13418 (N_13418,N_13311,N_13213);
xor U13419 (N_13419,N_13289,N_13278);
nor U13420 (N_13420,N_13324,N_13286);
nor U13421 (N_13421,N_13233,N_13270);
or U13422 (N_13422,N_13314,N_13331);
or U13423 (N_13423,N_13240,N_13206);
or U13424 (N_13424,N_13244,N_13347);
xor U13425 (N_13425,N_13213,N_13286);
or U13426 (N_13426,N_13222,N_13256);
or U13427 (N_13427,N_13304,N_13320);
nand U13428 (N_13428,N_13348,N_13238);
and U13429 (N_13429,N_13298,N_13231);
xnor U13430 (N_13430,N_13248,N_13270);
nand U13431 (N_13431,N_13215,N_13209);
nor U13432 (N_13432,N_13249,N_13203);
xnor U13433 (N_13433,N_13291,N_13236);
or U13434 (N_13434,N_13340,N_13303);
nor U13435 (N_13435,N_13338,N_13202);
or U13436 (N_13436,N_13279,N_13326);
and U13437 (N_13437,N_13208,N_13270);
nor U13438 (N_13438,N_13232,N_13335);
nand U13439 (N_13439,N_13286,N_13279);
nand U13440 (N_13440,N_13333,N_13322);
xor U13441 (N_13441,N_13244,N_13295);
xnor U13442 (N_13442,N_13229,N_13245);
and U13443 (N_13443,N_13237,N_13314);
nor U13444 (N_13444,N_13257,N_13248);
or U13445 (N_13445,N_13338,N_13316);
nand U13446 (N_13446,N_13227,N_13319);
xnor U13447 (N_13447,N_13340,N_13294);
and U13448 (N_13448,N_13212,N_13225);
or U13449 (N_13449,N_13207,N_13321);
and U13450 (N_13450,N_13293,N_13247);
xnor U13451 (N_13451,N_13253,N_13303);
nor U13452 (N_13452,N_13290,N_13205);
nand U13453 (N_13453,N_13235,N_13283);
nor U13454 (N_13454,N_13217,N_13237);
and U13455 (N_13455,N_13240,N_13233);
or U13456 (N_13456,N_13228,N_13280);
nor U13457 (N_13457,N_13340,N_13258);
nor U13458 (N_13458,N_13233,N_13321);
and U13459 (N_13459,N_13328,N_13325);
and U13460 (N_13460,N_13200,N_13255);
nand U13461 (N_13461,N_13234,N_13291);
nor U13462 (N_13462,N_13347,N_13217);
nand U13463 (N_13463,N_13253,N_13285);
xor U13464 (N_13464,N_13243,N_13329);
nand U13465 (N_13465,N_13202,N_13262);
nor U13466 (N_13466,N_13348,N_13295);
nand U13467 (N_13467,N_13305,N_13284);
or U13468 (N_13468,N_13230,N_13330);
or U13469 (N_13469,N_13275,N_13345);
xnor U13470 (N_13470,N_13287,N_13336);
or U13471 (N_13471,N_13291,N_13286);
or U13472 (N_13472,N_13346,N_13289);
nor U13473 (N_13473,N_13261,N_13344);
xor U13474 (N_13474,N_13204,N_13321);
xnor U13475 (N_13475,N_13211,N_13258);
nor U13476 (N_13476,N_13300,N_13234);
and U13477 (N_13477,N_13265,N_13229);
or U13478 (N_13478,N_13315,N_13205);
xnor U13479 (N_13479,N_13259,N_13324);
xor U13480 (N_13480,N_13304,N_13321);
and U13481 (N_13481,N_13285,N_13274);
xor U13482 (N_13482,N_13284,N_13334);
xnor U13483 (N_13483,N_13301,N_13210);
and U13484 (N_13484,N_13305,N_13277);
nor U13485 (N_13485,N_13287,N_13321);
xor U13486 (N_13486,N_13260,N_13220);
or U13487 (N_13487,N_13222,N_13202);
nor U13488 (N_13488,N_13320,N_13212);
nand U13489 (N_13489,N_13202,N_13251);
and U13490 (N_13490,N_13281,N_13276);
nand U13491 (N_13491,N_13261,N_13296);
or U13492 (N_13492,N_13346,N_13251);
nor U13493 (N_13493,N_13262,N_13259);
and U13494 (N_13494,N_13281,N_13331);
and U13495 (N_13495,N_13201,N_13344);
nor U13496 (N_13496,N_13203,N_13221);
xor U13497 (N_13497,N_13347,N_13210);
xnor U13498 (N_13498,N_13321,N_13246);
or U13499 (N_13499,N_13225,N_13264);
or U13500 (N_13500,N_13394,N_13399);
nor U13501 (N_13501,N_13383,N_13499);
nor U13502 (N_13502,N_13435,N_13434);
nor U13503 (N_13503,N_13440,N_13482);
nand U13504 (N_13504,N_13371,N_13448);
nand U13505 (N_13505,N_13454,N_13474);
xor U13506 (N_13506,N_13403,N_13477);
xor U13507 (N_13507,N_13445,N_13398);
nand U13508 (N_13508,N_13414,N_13361);
nor U13509 (N_13509,N_13393,N_13369);
xnor U13510 (N_13510,N_13379,N_13408);
and U13511 (N_13511,N_13473,N_13405);
nand U13512 (N_13512,N_13424,N_13491);
nand U13513 (N_13513,N_13367,N_13498);
and U13514 (N_13514,N_13433,N_13382);
and U13515 (N_13515,N_13372,N_13460);
nand U13516 (N_13516,N_13356,N_13436);
nand U13517 (N_13517,N_13396,N_13485);
or U13518 (N_13518,N_13457,N_13364);
nand U13519 (N_13519,N_13497,N_13442);
xor U13520 (N_13520,N_13409,N_13432);
and U13521 (N_13521,N_13384,N_13450);
xor U13522 (N_13522,N_13446,N_13401);
xnor U13523 (N_13523,N_13428,N_13465);
nand U13524 (N_13524,N_13378,N_13480);
nor U13525 (N_13525,N_13471,N_13486);
nand U13526 (N_13526,N_13483,N_13468);
and U13527 (N_13527,N_13478,N_13487);
and U13528 (N_13528,N_13415,N_13387);
xor U13529 (N_13529,N_13492,N_13366);
or U13530 (N_13530,N_13417,N_13449);
nand U13531 (N_13531,N_13464,N_13430);
or U13532 (N_13532,N_13385,N_13395);
nor U13533 (N_13533,N_13466,N_13370);
nand U13534 (N_13534,N_13444,N_13397);
nand U13535 (N_13535,N_13493,N_13388);
nor U13536 (N_13536,N_13475,N_13459);
nor U13537 (N_13537,N_13462,N_13476);
nand U13538 (N_13538,N_13443,N_13365);
xnor U13539 (N_13539,N_13423,N_13437);
nand U13540 (N_13540,N_13429,N_13377);
nand U13541 (N_13541,N_13494,N_13421);
nand U13542 (N_13542,N_13407,N_13376);
nor U13543 (N_13543,N_13455,N_13422);
and U13544 (N_13544,N_13375,N_13431);
nand U13545 (N_13545,N_13351,N_13456);
or U13546 (N_13546,N_13495,N_13380);
and U13547 (N_13547,N_13390,N_13439);
nor U13548 (N_13548,N_13363,N_13452);
and U13549 (N_13549,N_13425,N_13353);
xnor U13550 (N_13550,N_13426,N_13420);
or U13551 (N_13551,N_13496,N_13402);
nand U13552 (N_13552,N_13481,N_13386);
or U13553 (N_13553,N_13427,N_13451);
xnor U13554 (N_13554,N_13463,N_13411);
nand U13555 (N_13555,N_13469,N_13490);
and U13556 (N_13556,N_13410,N_13381);
and U13557 (N_13557,N_13412,N_13453);
nand U13558 (N_13558,N_13357,N_13389);
nor U13559 (N_13559,N_13489,N_13484);
or U13560 (N_13560,N_13461,N_13373);
xor U13561 (N_13561,N_13362,N_13447);
xnor U13562 (N_13562,N_13488,N_13358);
and U13563 (N_13563,N_13419,N_13374);
xor U13564 (N_13564,N_13416,N_13352);
or U13565 (N_13565,N_13360,N_13354);
and U13566 (N_13566,N_13350,N_13413);
and U13567 (N_13567,N_13467,N_13470);
nand U13568 (N_13568,N_13472,N_13355);
nand U13569 (N_13569,N_13368,N_13392);
and U13570 (N_13570,N_13404,N_13441);
xnor U13571 (N_13571,N_13400,N_13438);
xor U13572 (N_13572,N_13418,N_13406);
nor U13573 (N_13573,N_13391,N_13458);
nand U13574 (N_13574,N_13479,N_13359);
nand U13575 (N_13575,N_13449,N_13446);
nor U13576 (N_13576,N_13446,N_13437);
and U13577 (N_13577,N_13365,N_13469);
nand U13578 (N_13578,N_13395,N_13498);
nand U13579 (N_13579,N_13434,N_13477);
nor U13580 (N_13580,N_13464,N_13392);
or U13581 (N_13581,N_13413,N_13443);
and U13582 (N_13582,N_13399,N_13483);
nand U13583 (N_13583,N_13421,N_13415);
nand U13584 (N_13584,N_13479,N_13466);
nor U13585 (N_13585,N_13388,N_13444);
xnor U13586 (N_13586,N_13361,N_13471);
xor U13587 (N_13587,N_13419,N_13402);
xnor U13588 (N_13588,N_13480,N_13414);
nand U13589 (N_13589,N_13494,N_13427);
nand U13590 (N_13590,N_13351,N_13404);
nor U13591 (N_13591,N_13393,N_13431);
or U13592 (N_13592,N_13353,N_13486);
nor U13593 (N_13593,N_13429,N_13419);
and U13594 (N_13594,N_13412,N_13371);
nor U13595 (N_13595,N_13379,N_13460);
nor U13596 (N_13596,N_13481,N_13374);
nand U13597 (N_13597,N_13483,N_13370);
xor U13598 (N_13598,N_13374,N_13429);
and U13599 (N_13599,N_13375,N_13405);
nor U13600 (N_13600,N_13495,N_13454);
nand U13601 (N_13601,N_13350,N_13471);
and U13602 (N_13602,N_13459,N_13462);
nor U13603 (N_13603,N_13455,N_13437);
nand U13604 (N_13604,N_13471,N_13417);
and U13605 (N_13605,N_13457,N_13465);
xnor U13606 (N_13606,N_13368,N_13487);
or U13607 (N_13607,N_13407,N_13383);
and U13608 (N_13608,N_13456,N_13410);
and U13609 (N_13609,N_13386,N_13358);
and U13610 (N_13610,N_13414,N_13440);
nor U13611 (N_13611,N_13365,N_13453);
nand U13612 (N_13612,N_13364,N_13460);
nand U13613 (N_13613,N_13439,N_13473);
nand U13614 (N_13614,N_13431,N_13443);
nand U13615 (N_13615,N_13466,N_13357);
or U13616 (N_13616,N_13462,N_13475);
nand U13617 (N_13617,N_13463,N_13409);
nand U13618 (N_13618,N_13418,N_13427);
xor U13619 (N_13619,N_13354,N_13497);
nand U13620 (N_13620,N_13355,N_13403);
nor U13621 (N_13621,N_13471,N_13377);
or U13622 (N_13622,N_13383,N_13472);
and U13623 (N_13623,N_13421,N_13404);
nand U13624 (N_13624,N_13384,N_13406);
nand U13625 (N_13625,N_13422,N_13353);
or U13626 (N_13626,N_13478,N_13476);
nand U13627 (N_13627,N_13483,N_13476);
or U13628 (N_13628,N_13488,N_13439);
nand U13629 (N_13629,N_13432,N_13357);
nor U13630 (N_13630,N_13357,N_13361);
nand U13631 (N_13631,N_13434,N_13353);
or U13632 (N_13632,N_13378,N_13463);
nand U13633 (N_13633,N_13361,N_13401);
nor U13634 (N_13634,N_13373,N_13372);
nand U13635 (N_13635,N_13479,N_13454);
and U13636 (N_13636,N_13432,N_13480);
xnor U13637 (N_13637,N_13434,N_13433);
xor U13638 (N_13638,N_13404,N_13481);
xnor U13639 (N_13639,N_13378,N_13474);
and U13640 (N_13640,N_13476,N_13453);
and U13641 (N_13641,N_13413,N_13465);
nor U13642 (N_13642,N_13467,N_13350);
and U13643 (N_13643,N_13356,N_13471);
xor U13644 (N_13644,N_13367,N_13450);
or U13645 (N_13645,N_13454,N_13434);
and U13646 (N_13646,N_13393,N_13491);
nor U13647 (N_13647,N_13441,N_13434);
nor U13648 (N_13648,N_13361,N_13442);
or U13649 (N_13649,N_13416,N_13423);
and U13650 (N_13650,N_13524,N_13571);
and U13651 (N_13651,N_13602,N_13625);
xor U13652 (N_13652,N_13509,N_13558);
xnor U13653 (N_13653,N_13636,N_13544);
xnor U13654 (N_13654,N_13582,N_13628);
nor U13655 (N_13655,N_13517,N_13549);
nor U13656 (N_13656,N_13633,N_13634);
nor U13657 (N_13657,N_13592,N_13501);
nor U13658 (N_13658,N_13564,N_13624);
and U13659 (N_13659,N_13503,N_13646);
and U13660 (N_13660,N_13559,N_13539);
and U13661 (N_13661,N_13529,N_13561);
nand U13662 (N_13662,N_13505,N_13599);
xnor U13663 (N_13663,N_13565,N_13572);
xor U13664 (N_13664,N_13626,N_13570);
nand U13665 (N_13665,N_13545,N_13635);
nand U13666 (N_13666,N_13641,N_13631);
or U13667 (N_13667,N_13598,N_13504);
nand U13668 (N_13668,N_13629,N_13613);
and U13669 (N_13669,N_13638,N_13563);
and U13670 (N_13670,N_13640,N_13531);
xnor U13671 (N_13671,N_13536,N_13630);
nand U13672 (N_13672,N_13502,N_13575);
or U13673 (N_13673,N_13555,N_13609);
nor U13674 (N_13674,N_13579,N_13557);
nand U13675 (N_13675,N_13615,N_13585);
or U13676 (N_13676,N_13548,N_13623);
and U13677 (N_13677,N_13526,N_13577);
xor U13678 (N_13678,N_13586,N_13632);
xor U13679 (N_13679,N_13590,N_13589);
nor U13680 (N_13680,N_13600,N_13617);
nor U13681 (N_13681,N_13540,N_13645);
or U13682 (N_13682,N_13533,N_13606);
nand U13683 (N_13683,N_13596,N_13560);
and U13684 (N_13684,N_13593,N_13546);
and U13685 (N_13685,N_13607,N_13622);
nor U13686 (N_13686,N_13610,N_13552);
nor U13687 (N_13687,N_13566,N_13541);
nand U13688 (N_13688,N_13512,N_13511);
and U13689 (N_13689,N_13520,N_13538);
xnor U13690 (N_13690,N_13614,N_13543);
or U13691 (N_13691,N_13581,N_13611);
nand U13692 (N_13692,N_13618,N_13527);
nand U13693 (N_13693,N_13621,N_13525);
nor U13694 (N_13694,N_13574,N_13508);
and U13695 (N_13695,N_13594,N_13601);
nor U13696 (N_13696,N_13608,N_13643);
nor U13697 (N_13697,N_13583,N_13516);
and U13698 (N_13698,N_13642,N_13530);
xnor U13699 (N_13699,N_13522,N_13547);
nor U13700 (N_13700,N_13507,N_13604);
xnor U13701 (N_13701,N_13584,N_13556);
nand U13702 (N_13702,N_13528,N_13612);
nand U13703 (N_13703,N_13569,N_13587);
xnor U13704 (N_13704,N_13513,N_13554);
nor U13705 (N_13705,N_13537,N_13580);
xnor U13706 (N_13706,N_13567,N_13644);
or U13707 (N_13707,N_13616,N_13510);
xor U13708 (N_13708,N_13519,N_13553);
nand U13709 (N_13709,N_13627,N_13573);
and U13710 (N_13710,N_13649,N_13576);
or U13711 (N_13711,N_13532,N_13620);
nand U13712 (N_13712,N_13500,N_13550);
or U13713 (N_13713,N_13637,N_13605);
and U13714 (N_13714,N_13514,N_13595);
and U13715 (N_13715,N_13603,N_13597);
and U13716 (N_13716,N_13523,N_13648);
nand U13717 (N_13717,N_13562,N_13551);
xnor U13718 (N_13718,N_13591,N_13518);
nand U13719 (N_13719,N_13515,N_13535);
nor U13720 (N_13720,N_13647,N_13639);
or U13721 (N_13721,N_13578,N_13588);
or U13722 (N_13722,N_13568,N_13619);
and U13723 (N_13723,N_13534,N_13542);
and U13724 (N_13724,N_13521,N_13506);
nor U13725 (N_13725,N_13564,N_13618);
and U13726 (N_13726,N_13617,N_13621);
or U13727 (N_13727,N_13524,N_13598);
and U13728 (N_13728,N_13590,N_13546);
and U13729 (N_13729,N_13622,N_13610);
or U13730 (N_13730,N_13642,N_13630);
and U13731 (N_13731,N_13594,N_13583);
nor U13732 (N_13732,N_13513,N_13546);
nor U13733 (N_13733,N_13522,N_13534);
and U13734 (N_13734,N_13518,N_13615);
or U13735 (N_13735,N_13551,N_13554);
or U13736 (N_13736,N_13588,N_13602);
xnor U13737 (N_13737,N_13611,N_13536);
nand U13738 (N_13738,N_13533,N_13512);
nor U13739 (N_13739,N_13638,N_13615);
nor U13740 (N_13740,N_13590,N_13632);
nand U13741 (N_13741,N_13534,N_13509);
xor U13742 (N_13742,N_13525,N_13597);
xnor U13743 (N_13743,N_13589,N_13503);
xor U13744 (N_13744,N_13550,N_13624);
or U13745 (N_13745,N_13536,N_13623);
nor U13746 (N_13746,N_13500,N_13640);
nand U13747 (N_13747,N_13523,N_13515);
xnor U13748 (N_13748,N_13516,N_13578);
and U13749 (N_13749,N_13530,N_13600);
or U13750 (N_13750,N_13513,N_13638);
xor U13751 (N_13751,N_13608,N_13551);
or U13752 (N_13752,N_13616,N_13583);
and U13753 (N_13753,N_13531,N_13536);
xnor U13754 (N_13754,N_13533,N_13570);
or U13755 (N_13755,N_13588,N_13508);
nor U13756 (N_13756,N_13637,N_13526);
nor U13757 (N_13757,N_13617,N_13583);
nand U13758 (N_13758,N_13507,N_13611);
nor U13759 (N_13759,N_13509,N_13500);
nor U13760 (N_13760,N_13620,N_13512);
and U13761 (N_13761,N_13587,N_13635);
or U13762 (N_13762,N_13546,N_13553);
and U13763 (N_13763,N_13514,N_13644);
xor U13764 (N_13764,N_13518,N_13647);
or U13765 (N_13765,N_13648,N_13506);
or U13766 (N_13766,N_13503,N_13541);
xnor U13767 (N_13767,N_13629,N_13530);
xor U13768 (N_13768,N_13543,N_13572);
and U13769 (N_13769,N_13616,N_13542);
nor U13770 (N_13770,N_13519,N_13611);
nand U13771 (N_13771,N_13567,N_13611);
or U13772 (N_13772,N_13643,N_13504);
xnor U13773 (N_13773,N_13591,N_13605);
xnor U13774 (N_13774,N_13510,N_13636);
xor U13775 (N_13775,N_13588,N_13561);
nor U13776 (N_13776,N_13616,N_13540);
nor U13777 (N_13777,N_13520,N_13580);
nor U13778 (N_13778,N_13523,N_13542);
xnor U13779 (N_13779,N_13617,N_13633);
nor U13780 (N_13780,N_13588,N_13642);
nor U13781 (N_13781,N_13502,N_13580);
nand U13782 (N_13782,N_13556,N_13583);
and U13783 (N_13783,N_13631,N_13519);
nand U13784 (N_13784,N_13509,N_13613);
nand U13785 (N_13785,N_13550,N_13508);
nand U13786 (N_13786,N_13507,N_13591);
nor U13787 (N_13787,N_13541,N_13523);
and U13788 (N_13788,N_13549,N_13624);
nor U13789 (N_13789,N_13588,N_13514);
xor U13790 (N_13790,N_13563,N_13511);
nor U13791 (N_13791,N_13501,N_13524);
or U13792 (N_13792,N_13559,N_13557);
and U13793 (N_13793,N_13537,N_13543);
nor U13794 (N_13794,N_13634,N_13564);
and U13795 (N_13795,N_13553,N_13505);
and U13796 (N_13796,N_13584,N_13579);
and U13797 (N_13797,N_13635,N_13574);
and U13798 (N_13798,N_13540,N_13537);
nor U13799 (N_13799,N_13530,N_13606);
nand U13800 (N_13800,N_13736,N_13769);
or U13801 (N_13801,N_13666,N_13791);
nand U13802 (N_13802,N_13688,N_13659);
or U13803 (N_13803,N_13777,N_13762);
and U13804 (N_13804,N_13674,N_13765);
xnor U13805 (N_13805,N_13658,N_13778);
or U13806 (N_13806,N_13718,N_13707);
nand U13807 (N_13807,N_13668,N_13684);
xor U13808 (N_13808,N_13759,N_13673);
nand U13809 (N_13809,N_13716,N_13671);
nand U13810 (N_13810,N_13774,N_13746);
nor U13811 (N_13811,N_13715,N_13680);
or U13812 (N_13812,N_13723,N_13689);
xor U13813 (N_13813,N_13705,N_13734);
or U13814 (N_13814,N_13748,N_13683);
and U13815 (N_13815,N_13799,N_13768);
nor U13816 (N_13816,N_13726,N_13754);
or U13817 (N_13817,N_13795,N_13706);
or U13818 (N_13818,N_13787,N_13784);
nor U13819 (N_13819,N_13770,N_13731);
nand U13820 (N_13820,N_13662,N_13792);
xnor U13821 (N_13821,N_13693,N_13697);
nor U13822 (N_13822,N_13737,N_13696);
xor U13823 (N_13823,N_13656,N_13650);
nand U13824 (N_13824,N_13758,N_13665);
and U13825 (N_13825,N_13661,N_13744);
nor U13826 (N_13826,N_13789,N_13740);
or U13827 (N_13827,N_13678,N_13719);
xor U13828 (N_13828,N_13767,N_13763);
nor U13829 (N_13829,N_13670,N_13663);
and U13830 (N_13830,N_13729,N_13738);
xor U13831 (N_13831,N_13781,N_13692);
xnor U13832 (N_13832,N_13750,N_13788);
or U13833 (N_13833,N_13793,N_13798);
nand U13834 (N_13834,N_13681,N_13755);
and U13835 (N_13835,N_13752,N_13717);
xor U13836 (N_13836,N_13790,N_13794);
nand U13837 (N_13837,N_13771,N_13780);
nand U13838 (N_13838,N_13653,N_13669);
or U13839 (N_13839,N_13710,N_13725);
xnor U13840 (N_13840,N_13772,N_13700);
and U13841 (N_13841,N_13728,N_13651);
nand U13842 (N_13842,N_13757,N_13749);
nor U13843 (N_13843,N_13751,N_13753);
nor U13844 (N_13844,N_13694,N_13775);
nor U13845 (N_13845,N_13733,N_13779);
nor U13846 (N_13846,N_13785,N_13732);
xnor U13847 (N_13847,N_13672,N_13766);
nor U13848 (N_13848,N_13742,N_13730);
nand U13849 (N_13849,N_13695,N_13704);
and U13850 (N_13850,N_13677,N_13796);
xor U13851 (N_13851,N_13735,N_13664);
nor U13852 (N_13852,N_13682,N_13676);
xor U13853 (N_13853,N_13782,N_13727);
xnor U13854 (N_13854,N_13714,N_13739);
xor U13855 (N_13855,N_13776,N_13722);
xor U13856 (N_13856,N_13724,N_13760);
or U13857 (N_13857,N_13721,N_13657);
nand U13858 (N_13858,N_13698,N_13745);
or U13859 (N_13859,N_13720,N_13786);
or U13860 (N_13860,N_13667,N_13687);
nand U13861 (N_13861,N_13783,N_13761);
xnor U13862 (N_13862,N_13711,N_13699);
xnor U13863 (N_13863,N_13690,N_13660);
nor U13864 (N_13864,N_13654,N_13709);
nor U13865 (N_13865,N_13713,N_13652);
or U13866 (N_13866,N_13701,N_13686);
and U13867 (N_13867,N_13691,N_13685);
xnor U13868 (N_13868,N_13743,N_13708);
nand U13869 (N_13869,N_13797,N_13764);
nand U13870 (N_13870,N_13741,N_13747);
nor U13871 (N_13871,N_13675,N_13773);
and U13872 (N_13872,N_13655,N_13756);
and U13873 (N_13873,N_13712,N_13679);
and U13874 (N_13874,N_13702,N_13703);
nand U13875 (N_13875,N_13664,N_13799);
nand U13876 (N_13876,N_13669,N_13777);
or U13877 (N_13877,N_13767,N_13691);
and U13878 (N_13878,N_13757,N_13673);
and U13879 (N_13879,N_13788,N_13768);
nor U13880 (N_13880,N_13737,N_13668);
nand U13881 (N_13881,N_13695,N_13783);
nand U13882 (N_13882,N_13755,N_13794);
nor U13883 (N_13883,N_13691,N_13701);
and U13884 (N_13884,N_13701,N_13651);
nand U13885 (N_13885,N_13706,N_13772);
nor U13886 (N_13886,N_13680,N_13665);
nand U13887 (N_13887,N_13683,N_13776);
or U13888 (N_13888,N_13762,N_13688);
or U13889 (N_13889,N_13788,N_13753);
nand U13890 (N_13890,N_13719,N_13736);
nor U13891 (N_13891,N_13785,N_13728);
nand U13892 (N_13892,N_13781,N_13754);
and U13893 (N_13893,N_13732,N_13761);
or U13894 (N_13894,N_13755,N_13739);
or U13895 (N_13895,N_13703,N_13784);
nor U13896 (N_13896,N_13768,N_13785);
xor U13897 (N_13897,N_13669,N_13789);
nor U13898 (N_13898,N_13738,N_13766);
xnor U13899 (N_13899,N_13681,N_13784);
and U13900 (N_13900,N_13650,N_13704);
nor U13901 (N_13901,N_13776,N_13762);
nor U13902 (N_13902,N_13795,N_13694);
and U13903 (N_13903,N_13755,N_13706);
nand U13904 (N_13904,N_13795,N_13719);
and U13905 (N_13905,N_13670,N_13682);
or U13906 (N_13906,N_13732,N_13779);
nand U13907 (N_13907,N_13781,N_13695);
xor U13908 (N_13908,N_13695,N_13701);
nand U13909 (N_13909,N_13673,N_13748);
and U13910 (N_13910,N_13666,N_13785);
nand U13911 (N_13911,N_13729,N_13658);
and U13912 (N_13912,N_13795,N_13744);
xor U13913 (N_13913,N_13777,N_13708);
nor U13914 (N_13914,N_13718,N_13747);
xnor U13915 (N_13915,N_13734,N_13733);
xnor U13916 (N_13916,N_13677,N_13692);
and U13917 (N_13917,N_13695,N_13759);
or U13918 (N_13918,N_13676,N_13707);
nor U13919 (N_13919,N_13760,N_13716);
xnor U13920 (N_13920,N_13655,N_13657);
and U13921 (N_13921,N_13716,N_13762);
or U13922 (N_13922,N_13707,N_13692);
xor U13923 (N_13923,N_13752,N_13784);
and U13924 (N_13924,N_13785,N_13718);
nor U13925 (N_13925,N_13674,N_13711);
and U13926 (N_13926,N_13769,N_13709);
nand U13927 (N_13927,N_13708,N_13787);
xor U13928 (N_13928,N_13695,N_13752);
or U13929 (N_13929,N_13758,N_13781);
nand U13930 (N_13930,N_13760,N_13759);
nand U13931 (N_13931,N_13651,N_13774);
and U13932 (N_13932,N_13652,N_13663);
and U13933 (N_13933,N_13714,N_13794);
nand U13934 (N_13934,N_13662,N_13698);
or U13935 (N_13935,N_13779,N_13746);
xnor U13936 (N_13936,N_13697,N_13679);
xnor U13937 (N_13937,N_13752,N_13786);
and U13938 (N_13938,N_13686,N_13784);
nand U13939 (N_13939,N_13722,N_13731);
and U13940 (N_13940,N_13761,N_13753);
nor U13941 (N_13941,N_13789,N_13655);
or U13942 (N_13942,N_13715,N_13768);
nor U13943 (N_13943,N_13685,N_13739);
or U13944 (N_13944,N_13741,N_13664);
or U13945 (N_13945,N_13739,N_13733);
nand U13946 (N_13946,N_13672,N_13695);
or U13947 (N_13947,N_13766,N_13754);
and U13948 (N_13948,N_13665,N_13692);
or U13949 (N_13949,N_13745,N_13794);
and U13950 (N_13950,N_13888,N_13927);
and U13951 (N_13951,N_13934,N_13866);
nor U13952 (N_13952,N_13814,N_13838);
or U13953 (N_13953,N_13919,N_13902);
nand U13954 (N_13954,N_13860,N_13899);
and U13955 (N_13955,N_13900,N_13808);
or U13956 (N_13956,N_13874,N_13868);
nand U13957 (N_13957,N_13831,N_13824);
or U13958 (N_13958,N_13800,N_13908);
and U13959 (N_13959,N_13869,N_13842);
nor U13960 (N_13960,N_13820,N_13804);
or U13961 (N_13961,N_13819,N_13871);
and U13962 (N_13962,N_13889,N_13851);
nor U13963 (N_13963,N_13859,N_13893);
or U13964 (N_13964,N_13840,N_13827);
or U13965 (N_13965,N_13911,N_13920);
and U13966 (N_13966,N_13822,N_13855);
nand U13967 (N_13967,N_13903,N_13914);
or U13968 (N_13968,N_13816,N_13890);
nor U13969 (N_13969,N_13844,N_13873);
nand U13970 (N_13970,N_13846,N_13940);
or U13971 (N_13971,N_13882,N_13916);
xor U13972 (N_13972,N_13850,N_13917);
nor U13973 (N_13973,N_13807,N_13885);
or U13974 (N_13974,N_13837,N_13865);
and U13975 (N_13975,N_13937,N_13939);
nor U13976 (N_13976,N_13817,N_13830);
and U13977 (N_13977,N_13936,N_13884);
nor U13978 (N_13978,N_13922,N_13905);
nor U13979 (N_13979,N_13848,N_13943);
and U13980 (N_13980,N_13834,N_13941);
xor U13981 (N_13981,N_13921,N_13935);
and U13982 (N_13982,N_13826,N_13867);
and U13983 (N_13983,N_13926,N_13811);
xor U13984 (N_13984,N_13862,N_13913);
nand U13985 (N_13985,N_13895,N_13938);
nand U13986 (N_13986,N_13815,N_13947);
nand U13987 (N_13987,N_13856,N_13877);
nor U13988 (N_13988,N_13883,N_13946);
xnor U13989 (N_13989,N_13847,N_13894);
xor U13990 (N_13990,N_13887,N_13929);
xnor U13991 (N_13991,N_13909,N_13853);
nand U13992 (N_13992,N_13880,N_13898);
nor U13993 (N_13993,N_13876,N_13861);
xnor U13994 (N_13994,N_13949,N_13944);
or U13995 (N_13995,N_13803,N_13915);
xor U13996 (N_13996,N_13864,N_13836);
nand U13997 (N_13997,N_13818,N_13825);
xor U13998 (N_13998,N_13806,N_13863);
nand U13999 (N_13999,N_13904,N_13881);
or U14000 (N_14000,N_13802,N_13924);
or U14001 (N_14001,N_13854,N_13896);
or U14002 (N_14002,N_13948,N_13892);
xor U14003 (N_14003,N_13910,N_13886);
and U14004 (N_14004,N_13810,N_13945);
nand U14005 (N_14005,N_13832,N_13933);
and U14006 (N_14006,N_13858,N_13843);
nor U14007 (N_14007,N_13809,N_13907);
nor U14008 (N_14008,N_13812,N_13849);
nand U14009 (N_14009,N_13813,N_13823);
or U14010 (N_14010,N_13912,N_13932);
or U14011 (N_14011,N_13828,N_13857);
and U14012 (N_14012,N_13801,N_13897);
nor U14013 (N_14013,N_13852,N_13870);
and U14014 (N_14014,N_13872,N_13805);
and U14015 (N_14015,N_13906,N_13925);
and U14016 (N_14016,N_13835,N_13829);
nand U14017 (N_14017,N_13821,N_13918);
nor U14018 (N_14018,N_13878,N_13879);
and U14019 (N_14019,N_13875,N_13930);
and U14020 (N_14020,N_13928,N_13923);
or U14021 (N_14021,N_13901,N_13931);
nor U14022 (N_14022,N_13891,N_13845);
xor U14023 (N_14023,N_13833,N_13942);
nor U14024 (N_14024,N_13839,N_13841);
xnor U14025 (N_14025,N_13922,N_13874);
nand U14026 (N_14026,N_13891,N_13934);
nor U14027 (N_14027,N_13873,N_13890);
nand U14028 (N_14028,N_13946,N_13895);
and U14029 (N_14029,N_13911,N_13875);
xnor U14030 (N_14030,N_13890,N_13844);
nor U14031 (N_14031,N_13833,N_13924);
or U14032 (N_14032,N_13895,N_13948);
nor U14033 (N_14033,N_13813,N_13825);
or U14034 (N_14034,N_13942,N_13845);
nor U14035 (N_14035,N_13842,N_13819);
and U14036 (N_14036,N_13885,N_13924);
nor U14037 (N_14037,N_13931,N_13899);
nor U14038 (N_14038,N_13800,N_13846);
xnor U14039 (N_14039,N_13937,N_13887);
xor U14040 (N_14040,N_13907,N_13860);
and U14041 (N_14041,N_13942,N_13830);
xnor U14042 (N_14042,N_13934,N_13878);
nor U14043 (N_14043,N_13863,N_13937);
xnor U14044 (N_14044,N_13923,N_13947);
and U14045 (N_14045,N_13822,N_13947);
nand U14046 (N_14046,N_13806,N_13886);
and U14047 (N_14047,N_13839,N_13810);
xor U14048 (N_14048,N_13839,N_13924);
xnor U14049 (N_14049,N_13893,N_13862);
and U14050 (N_14050,N_13842,N_13888);
xnor U14051 (N_14051,N_13846,N_13883);
and U14052 (N_14052,N_13881,N_13852);
nand U14053 (N_14053,N_13823,N_13844);
xnor U14054 (N_14054,N_13817,N_13848);
and U14055 (N_14055,N_13881,N_13937);
nor U14056 (N_14056,N_13899,N_13826);
or U14057 (N_14057,N_13824,N_13933);
nand U14058 (N_14058,N_13828,N_13916);
xor U14059 (N_14059,N_13884,N_13893);
xnor U14060 (N_14060,N_13906,N_13935);
nand U14061 (N_14061,N_13805,N_13836);
nand U14062 (N_14062,N_13844,N_13891);
and U14063 (N_14063,N_13806,N_13802);
nor U14064 (N_14064,N_13929,N_13922);
nor U14065 (N_14065,N_13873,N_13939);
xnor U14066 (N_14066,N_13868,N_13876);
or U14067 (N_14067,N_13937,N_13921);
and U14068 (N_14068,N_13835,N_13892);
or U14069 (N_14069,N_13921,N_13890);
xor U14070 (N_14070,N_13917,N_13886);
or U14071 (N_14071,N_13920,N_13838);
and U14072 (N_14072,N_13899,N_13872);
and U14073 (N_14073,N_13863,N_13849);
nor U14074 (N_14074,N_13826,N_13862);
xor U14075 (N_14075,N_13885,N_13880);
nor U14076 (N_14076,N_13805,N_13884);
nand U14077 (N_14077,N_13910,N_13877);
nor U14078 (N_14078,N_13938,N_13832);
and U14079 (N_14079,N_13841,N_13937);
xnor U14080 (N_14080,N_13934,N_13893);
and U14081 (N_14081,N_13948,N_13840);
or U14082 (N_14082,N_13888,N_13914);
and U14083 (N_14083,N_13878,N_13827);
or U14084 (N_14084,N_13939,N_13902);
nand U14085 (N_14085,N_13909,N_13947);
and U14086 (N_14086,N_13805,N_13849);
nand U14087 (N_14087,N_13826,N_13855);
xnor U14088 (N_14088,N_13875,N_13917);
xnor U14089 (N_14089,N_13874,N_13946);
xor U14090 (N_14090,N_13918,N_13942);
nor U14091 (N_14091,N_13843,N_13921);
and U14092 (N_14092,N_13873,N_13935);
or U14093 (N_14093,N_13908,N_13896);
nor U14094 (N_14094,N_13898,N_13896);
and U14095 (N_14095,N_13843,N_13851);
or U14096 (N_14096,N_13904,N_13802);
nand U14097 (N_14097,N_13947,N_13868);
nor U14098 (N_14098,N_13823,N_13920);
or U14099 (N_14099,N_13817,N_13809);
xnor U14100 (N_14100,N_14079,N_14049);
and U14101 (N_14101,N_14000,N_14094);
nor U14102 (N_14102,N_14088,N_13962);
or U14103 (N_14103,N_13956,N_13999);
nand U14104 (N_14104,N_14005,N_14096);
nor U14105 (N_14105,N_13958,N_13952);
xor U14106 (N_14106,N_14001,N_14076);
or U14107 (N_14107,N_14039,N_14030);
or U14108 (N_14108,N_14099,N_13995);
nor U14109 (N_14109,N_14020,N_13992);
and U14110 (N_14110,N_14085,N_14002);
or U14111 (N_14111,N_13964,N_13959);
nor U14112 (N_14112,N_13996,N_14078);
or U14113 (N_14113,N_14023,N_13981);
xor U14114 (N_14114,N_14042,N_14071);
nor U14115 (N_14115,N_14058,N_14051);
and U14116 (N_14116,N_14047,N_14087);
nand U14117 (N_14117,N_14065,N_14014);
xor U14118 (N_14118,N_13961,N_13977);
xnor U14119 (N_14119,N_14070,N_13954);
or U14120 (N_14120,N_13986,N_14041);
nor U14121 (N_14121,N_14026,N_14009);
nand U14122 (N_14122,N_13991,N_14040);
nor U14123 (N_14123,N_14043,N_14074);
nor U14124 (N_14124,N_13980,N_14003);
and U14125 (N_14125,N_13976,N_13965);
xnor U14126 (N_14126,N_14095,N_14077);
and U14127 (N_14127,N_13984,N_14055);
nand U14128 (N_14128,N_14013,N_14044);
xnor U14129 (N_14129,N_14081,N_14015);
nand U14130 (N_14130,N_14091,N_13970);
nor U14131 (N_14131,N_14057,N_14056);
xor U14132 (N_14132,N_13955,N_14048);
nor U14133 (N_14133,N_14016,N_13966);
nand U14134 (N_14134,N_14032,N_14033);
nand U14135 (N_14135,N_14021,N_14037);
nor U14136 (N_14136,N_14069,N_13971);
nand U14137 (N_14137,N_13979,N_13974);
nor U14138 (N_14138,N_14008,N_13983);
xnor U14139 (N_14139,N_14063,N_14004);
and U14140 (N_14140,N_14034,N_13951);
and U14141 (N_14141,N_14007,N_13993);
nor U14142 (N_14142,N_14067,N_13957);
xnor U14143 (N_14143,N_14053,N_14019);
or U14144 (N_14144,N_13975,N_14031);
xnor U14145 (N_14145,N_14086,N_14006);
xor U14146 (N_14146,N_13969,N_14027);
nor U14147 (N_14147,N_14097,N_13963);
nand U14148 (N_14148,N_14024,N_14092);
xnor U14149 (N_14149,N_14098,N_13987);
and U14150 (N_14150,N_14045,N_14012);
and U14151 (N_14151,N_14036,N_13950);
xnor U14152 (N_14152,N_13960,N_14018);
and U14153 (N_14153,N_14068,N_13978);
and U14154 (N_14154,N_13998,N_14073);
and U14155 (N_14155,N_14054,N_14050);
xnor U14156 (N_14156,N_14062,N_13994);
and U14157 (N_14157,N_14022,N_14075);
xnor U14158 (N_14158,N_13982,N_14061);
nor U14159 (N_14159,N_14066,N_14072);
xor U14160 (N_14160,N_14017,N_14035);
and U14161 (N_14161,N_13997,N_13990);
or U14162 (N_14162,N_14025,N_14083);
xor U14163 (N_14163,N_13953,N_13988);
nor U14164 (N_14164,N_14010,N_13967);
xor U14165 (N_14165,N_14059,N_13989);
or U14166 (N_14166,N_14038,N_14064);
and U14167 (N_14167,N_13972,N_14080);
nand U14168 (N_14168,N_14052,N_14082);
nand U14169 (N_14169,N_14028,N_14089);
or U14170 (N_14170,N_13968,N_14090);
or U14171 (N_14171,N_13973,N_14093);
and U14172 (N_14172,N_14011,N_14029);
xor U14173 (N_14173,N_14084,N_13985);
xor U14174 (N_14174,N_14046,N_14060);
nor U14175 (N_14175,N_14072,N_13989);
and U14176 (N_14176,N_14075,N_14066);
xor U14177 (N_14177,N_14042,N_14077);
nor U14178 (N_14178,N_14055,N_14019);
and U14179 (N_14179,N_14087,N_14075);
or U14180 (N_14180,N_14058,N_14068);
xnor U14181 (N_14181,N_14055,N_14046);
or U14182 (N_14182,N_14091,N_13974);
nand U14183 (N_14183,N_14009,N_13976);
or U14184 (N_14184,N_14005,N_14015);
or U14185 (N_14185,N_14089,N_13990);
or U14186 (N_14186,N_13978,N_14094);
nor U14187 (N_14187,N_14085,N_13973);
and U14188 (N_14188,N_13967,N_13973);
nor U14189 (N_14189,N_13956,N_14027);
nor U14190 (N_14190,N_14005,N_13962);
nor U14191 (N_14191,N_14064,N_14042);
xnor U14192 (N_14192,N_14058,N_13981);
or U14193 (N_14193,N_14042,N_14047);
xor U14194 (N_14194,N_13994,N_13962);
and U14195 (N_14195,N_14006,N_14098);
or U14196 (N_14196,N_14096,N_14030);
xor U14197 (N_14197,N_14042,N_14091);
and U14198 (N_14198,N_14096,N_13952);
or U14199 (N_14199,N_14031,N_13971);
nand U14200 (N_14200,N_14036,N_13962);
or U14201 (N_14201,N_14055,N_13992);
xor U14202 (N_14202,N_14051,N_14092);
nand U14203 (N_14203,N_14074,N_14081);
nor U14204 (N_14204,N_14082,N_14038);
nor U14205 (N_14205,N_14023,N_13979);
nor U14206 (N_14206,N_14046,N_14020);
and U14207 (N_14207,N_14085,N_13968);
or U14208 (N_14208,N_14054,N_14064);
or U14209 (N_14209,N_14074,N_14002);
or U14210 (N_14210,N_13971,N_13972);
xnor U14211 (N_14211,N_14094,N_14037);
nand U14212 (N_14212,N_14069,N_14016);
nor U14213 (N_14213,N_14077,N_14096);
or U14214 (N_14214,N_13981,N_14036);
and U14215 (N_14215,N_13979,N_13960);
or U14216 (N_14216,N_13961,N_13981);
and U14217 (N_14217,N_14003,N_13961);
nand U14218 (N_14218,N_13981,N_13986);
and U14219 (N_14219,N_14053,N_14000);
and U14220 (N_14220,N_13970,N_14079);
or U14221 (N_14221,N_14029,N_14018);
and U14222 (N_14222,N_14031,N_13955);
nand U14223 (N_14223,N_14035,N_14052);
nand U14224 (N_14224,N_14081,N_14065);
xor U14225 (N_14225,N_13984,N_13990);
nand U14226 (N_14226,N_13992,N_13991);
nand U14227 (N_14227,N_14059,N_13972);
and U14228 (N_14228,N_14070,N_14099);
and U14229 (N_14229,N_14007,N_14058);
xnor U14230 (N_14230,N_14080,N_13971);
xnor U14231 (N_14231,N_14054,N_13984);
or U14232 (N_14232,N_14030,N_14086);
nor U14233 (N_14233,N_13981,N_14089);
nand U14234 (N_14234,N_14004,N_13957);
and U14235 (N_14235,N_14083,N_13995);
nand U14236 (N_14236,N_14063,N_14046);
or U14237 (N_14237,N_13999,N_14096);
xor U14238 (N_14238,N_14033,N_13953);
and U14239 (N_14239,N_13996,N_14010);
nor U14240 (N_14240,N_14001,N_13965);
nor U14241 (N_14241,N_14044,N_14042);
and U14242 (N_14242,N_14040,N_14014);
or U14243 (N_14243,N_14071,N_14015);
nor U14244 (N_14244,N_14094,N_14008);
or U14245 (N_14245,N_13988,N_14076);
xor U14246 (N_14246,N_14057,N_14073);
or U14247 (N_14247,N_14065,N_14021);
nand U14248 (N_14248,N_14027,N_14036);
nand U14249 (N_14249,N_14069,N_14061);
nor U14250 (N_14250,N_14190,N_14143);
nand U14251 (N_14251,N_14142,N_14213);
nor U14252 (N_14252,N_14202,N_14185);
xnor U14253 (N_14253,N_14123,N_14187);
and U14254 (N_14254,N_14179,N_14219);
nand U14255 (N_14255,N_14113,N_14188);
and U14256 (N_14256,N_14216,N_14114);
nand U14257 (N_14257,N_14173,N_14122);
and U14258 (N_14258,N_14116,N_14151);
nor U14259 (N_14259,N_14101,N_14126);
xor U14260 (N_14260,N_14248,N_14249);
or U14261 (N_14261,N_14139,N_14140);
and U14262 (N_14262,N_14183,N_14106);
nand U14263 (N_14263,N_14132,N_14224);
and U14264 (N_14264,N_14209,N_14242);
and U14265 (N_14265,N_14233,N_14110);
xnor U14266 (N_14266,N_14189,N_14170);
or U14267 (N_14267,N_14223,N_14230);
nor U14268 (N_14268,N_14150,N_14119);
nor U14269 (N_14269,N_14239,N_14196);
and U14270 (N_14270,N_14246,N_14131);
and U14271 (N_14271,N_14177,N_14217);
nor U14272 (N_14272,N_14228,N_14163);
nand U14273 (N_14273,N_14135,N_14166);
nor U14274 (N_14274,N_14200,N_14164);
or U14275 (N_14275,N_14149,N_14171);
xor U14276 (N_14276,N_14137,N_14180);
and U14277 (N_14277,N_14229,N_14227);
nor U14278 (N_14278,N_14192,N_14201);
nand U14279 (N_14279,N_14136,N_14148);
nor U14280 (N_14280,N_14232,N_14161);
xnor U14281 (N_14281,N_14117,N_14193);
nor U14282 (N_14282,N_14167,N_14152);
xor U14283 (N_14283,N_14146,N_14147);
or U14284 (N_14284,N_14247,N_14208);
nand U14285 (N_14285,N_14220,N_14211);
or U14286 (N_14286,N_14194,N_14218);
nor U14287 (N_14287,N_14172,N_14100);
and U14288 (N_14288,N_14118,N_14207);
nand U14289 (N_14289,N_14231,N_14221);
xnor U14290 (N_14290,N_14153,N_14212);
and U14291 (N_14291,N_14127,N_14160);
nand U14292 (N_14292,N_14204,N_14130);
and U14293 (N_14293,N_14214,N_14103);
and U14294 (N_14294,N_14120,N_14156);
xor U14295 (N_14295,N_14141,N_14109);
xnor U14296 (N_14296,N_14111,N_14115);
nand U14297 (N_14297,N_14206,N_14125);
nand U14298 (N_14298,N_14154,N_14236);
nand U14299 (N_14299,N_14107,N_14159);
and U14300 (N_14300,N_14128,N_14168);
xor U14301 (N_14301,N_14176,N_14195);
nand U14302 (N_14302,N_14145,N_14121);
nor U14303 (N_14303,N_14178,N_14197);
or U14304 (N_14304,N_14157,N_14198);
nand U14305 (N_14305,N_14240,N_14174);
nand U14306 (N_14306,N_14238,N_14225);
or U14307 (N_14307,N_14134,N_14138);
nand U14308 (N_14308,N_14226,N_14133);
nand U14309 (N_14309,N_14144,N_14124);
or U14310 (N_14310,N_14102,N_14182);
nor U14311 (N_14311,N_14245,N_14205);
nor U14312 (N_14312,N_14129,N_14186);
or U14313 (N_14313,N_14210,N_14155);
nand U14314 (N_14314,N_14169,N_14165);
nand U14315 (N_14315,N_14108,N_14203);
and U14316 (N_14316,N_14243,N_14215);
and U14317 (N_14317,N_14105,N_14244);
nor U14318 (N_14318,N_14235,N_14112);
or U14319 (N_14319,N_14104,N_14158);
nor U14320 (N_14320,N_14237,N_14162);
nand U14321 (N_14321,N_14222,N_14184);
nand U14322 (N_14322,N_14241,N_14234);
xnor U14323 (N_14323,N_14199,N_14175);
or U14324 (N_14324,N_14191,N_14181);
xor U14325 (N_14325,N_14153,N_14120);
nor U14326 (N_14326,N_14130,N_14124);
or U14327 (N_14327,N_14103,N_14129);
and U14328 (N_14328,N_14151,N_14173);
and U14329 (N_14329,N_14162,N_14127);
or U14330 (N_14330,N_14136,N_14179);
xnor U14331 (N_14331,N_14171,N_14236);
nor U14332 (N_14332,N_14105,N_14190);
nand U14333 (N_14333,N_14124,N_14231);
nor U14334 (N_14334,N_14195,N_14166);
nand U14335 (N_14335,N_14178,N_14148);
nor U14336 (N_14336,N_14120,N_14222);
xnor U14337 (N_14337,N_14113,N_14184);
or U14338 (N_14338,N_14219,N_14145);
nor U14339 (N_14339,N_14181,N_14132);
nand U14340 (N_14340,N_14242,N_14178);
and U14341 (N_14341,N_14234,N_14215);
xor U14342 (N_14342,N_14238,N_14105);
xor U14343 (N_14343,N_14202,N_14159);
nor U14344 (N_14344,N_14228,N_14159);
and U14345 (N_14345,N_14103,N_14141);
xnor U14346 (N_14346,N_14162,N_14221);
xnor U14347 (N_14347,N_14159,N_14155);
nor U14348 (N_14348,N_14121,N_14146);
nand U14349 (N_14349,N_14211,N_14152);
and U14350 (N_14350,N_14199,N_14240);
or U14351 (N_14351,N_14113,N_14148);
xnor U14352 (N_14352,N_14106,N_14118);
xor U14353 (N_14353,N_14123,N_14244);
nand U14354 (N_14354,N_14148,N_14226);
nand U14355 (N_14355,N_14183,N_14178);
xnor U14356 (N_14356,N_14191,N_14109);
nand U14357 (N_14357,N_14105,N_14207);
xor U14358 (N_14358,N_14105,N_14189);
xnor U14359 (N_14359,N_14186,N_14221);
nor U14360 (N_14360,N_14196,N_14119);
and U14361 (N_14361,N_14145,N_14147);
nand U14362 (N_14362,N_14216,N_14153);
or U14363 (N_14363,N_14203,N_14163);
xor U14364 (N_14364,N_14207,N_14126);
nor U14365 (N_14365,N_14216,N_14145);
nand U14366 (N_14366,N_14199,N_14109);
or U14367 (N_14367,N_14204,N_14197);
and U14368 (N_14368,N_14138,N_14201);
xor U14369 (N_14369,N_14139,N_14213);
nor U14370 (N_14370,N_14137,N_14242);
or U14371 (N_14371,N_14143,N_14179);
xnor U14372 (N_14372,N_14149,N_14222);
and U14373 (N_14373,N_14198,N_14185);
xnor U14374 (N_14374,N_14170,N_14241);
or U14375 (N_14375,N_14195,N_14217);
nor U14376 (N_14376,N_14221,N_14102);
nand U14377 (N_14377,N_14133,N_14189);
and U14378 (N_14378,N_14112,N_14247);
or U14379 (N_14379,N_14175,N_14150);
and U14380 (N_14380,N_14107,N_14155);
nand U14381 (N_14381,N_14175,N_14232);
and U14382 (N_14382,N_14170,N_14175);
nor U14383 (N_14383,N_14244,N_14145);
nand U14384 (N_14384,N_14126,N_14229);
nor U14385 (N_14385,N_14189,N_14123);
xnor U14386 (N_14386,N_14115,N_14133);
xor U14387 (N_14387,N_14186,N_14231);
nor U14388 (N_14388,N_14139,N_14234);
and U14389 (N_14389,N_14240,N_14145);
nor U14390 (N_14390,N_14241,N_14199);
and U14391 (N_14391,N_14192,N_14228);
and U14392 (N_14392,N_14237,N_14165);
xor U14393 (N_14393,N_14190,N_14240);
and U14394 (N_14394,N_14231,N_14246);
or U14395 (N_14395,N_14215,N_14163);
and U14396 (N_14396,N_14133,N_14158);
nand U14397 (N_14397,N_14139,N_14222);
or U14398 (N_14398,N_14108,N_14182);
or U14399 (N_14399,N_14199,N_14168);
or U14400 (N_14400,N_14279,N_14358);
nor U14401 (N_14401,N_14381,N_14389);
and U14402 (N_14402,N_14298,N_14321);
or U14403 (N_14403,N_14386,N_14259);
or U14404 (N_14404,N_14383,N_14351);
nand U14405 (N_14405,N_14343,N_14364);
xor U14406 (N_14406,N_14257,N_14376);
nor U14407 (N_14407,N_14337,N_14303);
and U14408 (N_14408,N_14283,N_14355);
or U14409 (N_14409,N_14282,N_14286);
or U14410 (N_14410,N_14330,N_14378);
xor U14411 (N_14411,N_14338,N_14258);
nor U14412 (N_14412,N_14326,N_14306);
nand U14413 (N_14413,N_14371,N_14276);
nor U14414 (N_14414,N_14393,N_14366);
and U14415 (N_14415,N_14333,N_14292);
or U14416 (N_14416,N_14301,N_14290);
nand U14417 (N_14417,N_14356,N_14325);
or U14418 (N_14418,N_14250,N_14294);
or U14419 (N_14419,N_14287,N_14275);
and U14420 (N_14420,N_14300,N_14308);
or U14421 (N_14421,N_14387,N_14353);
xnor U14422 (N_14422,N_14305,N_14352);
nor U14423 (N_14423,N_14254,N_14372);
nand U14424 (N_14424,N_14314,N_14361);
and U14425 (N_14425,N_14293,N_14379);
or U14426 (N_14426,N_14331,N_14296);
nand U14427 (N_14427,N_14342,N_14396);
and U14428 (N_14428,N_14281,N_14318);
xnor U14429 (N_14429,N_14375,N_14272);
and U14430 (N_14430,N_14322,N_14374);
and U14431 (N_14431,N_14288,N_14302);
xnor U14432 (N_14432,N_14265,N_14362);
or U14433 (N_14433,N_14398,N_14267);
and U14434 (N_14434,N_14368,N_14345);
xor U14435 (N_14435,N_14385,N_14336);
nor U14436 (N_14436,N_14285,N_14307);
or U14437 (N_14437,N_14394,N_14274);
nand U14438 (N_14438,N_14297,N_14332);
and U14439 (N_14439,N_14320,N_14367);
xnor U14440 (N_14440,N_14316,N_14319);
nor U14441 (N_14441,N_14348,N_14255);
xor U14442 (N_14442,N_14392,N_14399);
nand U14443 (N_14443,N_14365,N_14390);
nor U14444 (N_14444,N_14280,N_14289);
nor U14445 (N_14445,N_14324,N_14339);
and U14446 (N_14446,N_14271,N_14388);
and U14447 (N_14447,N_14373,N_14309);
xnor U14448 (N_14448,N_14347,N_14377);
and U14449 (N_14449,N_14317,N_14312);
or U14450 (N_14450,N_14261,N_14369);
nand U14451 (N_14451,N_14344,N_14329);
and U14452 (N_14452,N_14323,N_14341);
nand U14453 (N_14453,N_14384,N_14310);
and U14454 (N_14454,N_14335,N_14295);
or U14455 (N_14455,N_14270,N_14252);
xor U14456 (N_14456,N_14260,N_14382);
xnor U14457 (N_14457,N_14397,N_14346);
xor U14458 (N_14458,N_14313,N_14349);
or U14459 (N_14459,N_14395,N_14284);
or U14460 (N_14460,N_14256,N_14278);
xor U14461 (N_14461,N_14315,N_14263);
xor U14462 (N_14462,N_14299,N_14291);
nor U14463 (N_14463,N_14334,N_14370);
nor U14464 (N_14464,N_14273,N_14251);
xor U14465 (N_14465,N_14359,N_14311);
nand U14466 (N_14466,N_14327,N_14264);
nand U14467 (N_14467,N_14363,N_14268);
and U14468 (N_14468,N_14277,N_14350);
nor U14469 (N_14469,N_14269,N_14266);
nor U14470 (N_14470,N_14253,N_14340);
and U14471 (N_14471,N_14262,N_14357);
nor U14472 (N_14472,N_14360,N_14328);
and U14473 (N_14473,N_14380,N_14391);
or U14474 (N_14474,N_14354,N_14304);
or U14475 (N_14475,N_14388,N_14327);
xnor U14476 (N_14476,N_14326,N_14286);
xor U14477 (N_14477,N_14343,N_14274);
and U14478 (N_14478,N_14340,N_14272);
nand U14479 (N_14479,N_14377,N_14282);
nor U14480 (N_14480,N_14331,N_14347);
nor U14481 (N_14481,N_14305,N_14387);
or U14482 (N_14482,N_14272,N_14262);
nor U14483 (N_14483,N_14319,N_14332);
or U14484 (N_14484,N_14303,N_14361);
nor U14485 (N_14485,N_14369,N_14266);
and U14486 (N_14486,N_14376,N_14252);
nand U14487 (N_14487,N_14350,N_14357);
or U14488 (N_14488,N_14260,N_14275);
xor U14489 (N_14489,N_14393,N_14257);
nor U14490 (N_14490,N_14290,N_14288);
and U14491 (N_14491,N_14304,N_14361);
and U14492 (N_14492,N_14360,N_14317);
nor U14493 (N_14493,N_14289,N_14388);
nor U14494 (N_14494,N_14356,N_14282);
nor U14495 (N_14495,N_14322,N_14270);
or U14496 (N_14496,N_14332,N_14314);
and U14497 (N_14497,N_14377,N_14322);
xnor U14498 (N_14498,N_14251,N_14263);
or U14499 (N_14499,N_14259,N_14276);
nor U14500 (N_14500,N_14268,N_14317);
nand U14501 (N_14501,N_14295,N_14366);
and U14502 (N_14502,N_14371,N_14357);
nor U14503 (N_14503,N_14256,N_14344);
or U14504 (N_14504,N_14303,N_14326);
xor U14505 (N_14505,N_14344,N_14335);
and U14506 (N_14506,N_14342,N_14301);
and U14507 (N_14507,N_14335,N_14338);
nor U14508 (N_14508,N_14393,N_14357);
and U14509 (N_14509,N_14397,N_14252);
or U14510 (N_14510,N_14261,N_14356);
nor U14511 (N_14511,N_14333,N_14267);
nand U14512 (N_14512,N_14380,N_14331);
or U14513 (N_14513,N_14297,N_14394);
nor U14514 (N_14514,N_14399,N_14263);
or U14515 (N_14515,N_14285,N_14296);
nor U14516 (N_14516,N_14386,N_14397);
nor U14517 (N_14517,N_14354,N_14381);
nor U14518 (N_14518,N_14379,N_14281);
nor U14519 (N_14519,N_14372,N_14335);
and U14520 (N_14520,N_14344,N_14353);
nand U14521 (N_14521,N_14323,N_14321);
or U14522 (N_14522,N_14339,N_14307);
nand U14523 (N_14523,N_14260,N_14351);
and U14524 (N_14524,N_14379,N_14310);
or U14525 (N_14525,N_14330,N_14371);
xor U14526 (N_14526,N_14399,N_14295);
and U14527 (N_14527,N_14390,N_14251);
and U14528 (N_14528,N_14255,N_14395);
and U14529 (N_14529,N_14269,N_14334);
and U14530 (N_14530,N_14359,N_14253);
and U14531 (N_14531,N_14375,N_14253);
and U14532 (N_14532,N_14381,N_14254);
nor U14533 (N_14533,N_14345,N_14317);
or U14534 (N_14534,N_14339,N_14361);
or U14535 (N_14535,N_14376,N_14365);
nor U14536 (N_14536,N_14274,N_14258);
xor U14537 (N_14537,N_14385,N_14395);
xor U14538 (N_14538,N_14383,N_14339);
nand U14539 (N_14539,N_14393,N_14296);
nor U14540 (N_14540,N_14299,N_14337);
or U14541 (N_14541,N_14324,N_14333);
nor U14542 (N_14542,N_14309,N_14396);
and U14543 (N_14543,N_14392,N_14253);
and U14544 (N_14544,N_14290,N_14356);
xor U14545 (N_14545,N_14279,N_14312);
nand U14546 (N_14546,N_14357,N_14380);
nand U14547 (N_14547,N_14293,N_14389);
xnor U14548 (N_14548,N_14342,N_14365);
and U14549 (N_14549,N_14364,N_14270);
nand U14550 (N_14550,N_14432,N_14538);
xor U14551 (N_14551,N_14503,N_14478);
or U14552 (N_14552,N_14507,N_14518);
and U14553 (N_14553,N_14421,N_14455);
nor U14554 (N_14554,N_14469,N_14470);
nor U14555 (N_14555,N_14522,N_14464);
nand U14556 (N_14556,N_14403,N_14449);
or U14557 (N_14557,N_14439,N_14480);
or U14558 (N_14558,N_14490,N_14400);
or U14559 (N_14559,N_14409,N_14498);
xnor U14560 (N_14560,N_14420,N_14505);
xnor U14561 (N_14561,N_14476,N_14483);
xnor U14562 (N_14562,N_14487,N_14404);
nor U14563 (N_14563,N_14504,N_14419);
xor U14564 (N_14564,N_14506,N_14516);
xor U14565 (N_14565,N_14405,N_14456);
xnor U14566 (N_14566,N_14494,N_14486);
nand U14567 (N_14567,N_14466,N_14406);
xnor U14568 (N_14568,N_14446,N_14477);
nand U14569 (N_14569,N_14465,N_14441);
or U14570 (N_14570,N_14544,N_14495);
or U14571 (N_14571,N_14435,N_14491);
xor U14572 (N_14572,N_14443,N_14467);
xnor U14573 (N_14573,N_14452,N_14461);
xnor U14574 (N_14574,N_14541,N_14423);
or U14575 (N_14575,N_14457,N_14526);
nor U14576 (N_14576,N_14524,N_14549);
xor U14577 (N_14577,N_14489,N_14417);
and U14578 (N_14578,N_14523,N_14407);
or U14579 (N_14579,N_14459,N_14448);
xnor U14580 (N_14580,N_14427,N_14513);
nand U14581 (N_14581,N_14434,N_14528);
and U14582 (N_14582,N_14473,N_14540);
nand U14583 (N_14583,N_14532,N_14501);
or U14584 (N_14584,N_14496,N_14547);
and U14585 (N_14585,N_14521,N_14440);
or U14586 (N_14586,N_14537,N_14502);
nor U14587 (N_14587,N_14431,N_14430);
or U14588 (N_14588,N_14482,N_14509);
nor U14589 (N_14589,N_14408,N_14425);
or U14590 (N_14590,N_14429,N_14493);
or U14591 (N_14591,N_14462,N_14536);
nand U14592 (N_14592,N_14539,N_14481);
or U14593 (N_14593,N_14492,N_14415);
and U14594 (N_14594,N_14548,N_14530);
nor U14595 (N_14595,N_14525,N_14531);
nor U14596 (N_14596,N_14412,N_14460);
or U14597 (N_14597,N_14414,N_14511);
nor U14598 (N_14598,N_14436,N_14508);
xnor U14599 (N_14599,N_14454,N_14422);
nor U14600 (N_14600,N_14401,N_14426);
or U14601 (N_14601,N_14515,N_14533);
nor U14602 (N_14602,N_14438,N_14542);
nand U14603 (N_14603,N_14444,N_14411);
and U14604 (N_14604,N_14445,N_14517);
xor U14605 (N_14605,N_14519,N_14485);
and U14606 (N_14606,N_14497,N_14453);
nand U14607 (N_14607,N_14442,N_14418);
or U14608 (N_14608,N_14514,N_14433);
nor U14609 (N_14609,N_14472,N_14499);
or U14610 (N_14610,N_14545,N_14468);
and U14611 (N_14611,N_14451,N_14529);
xnor U14612 (N_14612,N_14512,N_14484);
xnor U14613 (N_14613,N_14413,N_14475);
and U14614 (N_14614,N_14424,N_14535);
nor U14615 (N_14615,N_14428,N_14520);
or U14616 (N_14616,N_14410,N_14534);
xnor U14617 (N_14617,N_14458,N_14543);
nand U14618 (N_14618,N_14474,N_14402);
or U14619 (N_14619,N_14479,N_14471);
and U14620 (N_14620,N_14527,N_14447);
and U14621 (N_14621,N_14488,N_14450);
nor U14622 (N_14622,N_14416,N_14463);
nand U14623 (N_14623,N_14500,N_14510);
or U14624 (N_14624,N_14546,N_14437);
nor U14625 (N_14625,N_14480,N_14545);
or U14626 (N_14626,N_14533,N_14471);
and U14627 (N_14627,N_14479,N_14505);
nor U14628 (N_14628,N_14454,N_14448);
nand U14629 (N_14629,N_14414,N_14491);
and U14630 (N_14630,N_14420,N_14500);
and U14631 (N_14631,N_14489,N_14438);
nor U14632 (N_14632,N_14505,N_14489);
nor U14633 (N_14633,N_14410,N_14436);
nor U14634 (N_14634,N_14507,N_14449);
xor U14635 (N_14635,N_14465,N_14530);
xnor U14636 (N_14636,N_14492,N_14413);
nor U14637 (N_14637,N_14460,N_14474);
nor U14638 (N_14638,N_14459,N_14530);
xnor U14639 (N_14639,N_14537,N_14513);
xnor U14640 (N_14640,N_14485,N_14408);
nor U14641 (N_14641,N_14503,N_14477);
nand U14642 (N_14642,N_14474,N_14546);
nand U14643 (N_14643,N_14458,N_14438);
and U14644 (N_14644,N_14451,N_14424);
or U14645 (N_14645,N_14483,N_14446);
nor U14646 (N_14646,N_14425,N_14412);
nor U14647 (N_14647,N_14524,N_14445);
nand U14648 (N_14648,N_14468,N_14509);
or U14649 (N_14649,N_14414,N_14541);
and U14650 (N_14650,N_14516,N_14436);
xor U14651 (N_14651,N_14452,N_14495);
and U14652 (N_14652,N_14413,N_14470);
and U14653 (N_14653,N_14487,N_14419);
nand U14654 (N_14654,N_14463,N_14459);
and U14655 (N_14655,N_14539,N_14471);
nor U14656 (N_14656,N_14518,N_14445);
or U14657 (N_14657,N_14447,N_14529);
or U14658 (N_14658,N_14527,N_14466);
or U14659 (N_14659,N_14454,N_14524);
nand U14660 (N_14660,N_14504,N_14414);
nand U14661 (N_14661,N_14458,N_14539);
nand U14662 (N_14662,N_14484,N_14518);
and U14663 (N_14663,N_14539,N_14478);
nand U14664 (N_14664,N_14539,N_14483);
nand U14665 (N_14665,N_14470,N_14497);
nor U14666 (N_14666,N_14473,N_14498);
or U14667 (N_14667,N_14482,N_14490);
or U14668 (N_14668,N_14447,N_14523);
xnor U14669 (N_14669,N_14410,N_14536);
or U14670 (N_14670,N_14448,N_14522);
xnor U14671 (N_14671,N_14540,N_14472);
or U14672 (N_14672,N_14430,N_14422);
xnor U14673 (N_14673,N_14494,N_14529);
nand U14674 (N_14674,N_14474,N_14417);
nor U14675 (N_14675,N_14450,N_14547);
nand U14676 (N_14676,N_14513,N_14441);
nor U14677 (N_14677,N_14495,N_14406);
or U14678 (N_14678,N_14526,N_14416);
or U14679 (N_14679,N_14534,N_14435);
nand U14680 (N_14680,N_14521,N_14482);
nand U14681 (N_14681,N_14436,N_14491);
nand U14682 (N_14682,N_14452,N_14440);
or U14683 (N_14683,N_14498,N_14491);
nand U14684 (N_14684,N_14406,N_14544);
nor U14685 (N_14685,N_14507,N_14519);
nor U14686 (N_14686,N_14406,N_14509);
nand U14687 (N_14687,N_14528,N_14511);
nor U14688 (N_14688,N_14408,N_14445);
nor U14689 (N_14689,N_14417,N_14521);
nor U14690 (N_14690,N_14519,N_14547);
and U14691 (N_14691,N_14474,N_14504);
and U14692 (N_14692,N_14541,N_14433);
nand U14693 (N_14693,N_14431,N_14408);
or U14694 (N_14694,N_14498,N_14469);
and U14695 (N_14695,N_14491,N_14489);
xnor U14696 (N_14696,N_14537,N_14517);
nor U14697 (N_14697,N_14459,N_14432);
and U14698 (N_14698,N_14464,N_14443);
nand U14699 (N_14699,N_14480,N_14468);
and U14700 (N_14700,N_14571,N_14605);
nand U14701 (N_14701,N_14699,N_14603);
and U14702 (N_14702,N_14596,N_14607);
nand U14703 (N_14703,N_14556,N_14568);
nor U14704 (N_14704,N_14643,N_14640);
xor U14705 (N_14705,N_14561,N_14698);
nor U14706 (N_14706,N_14560,N_14609);
or U14707 (N_14707,N_14633,N_14625);
or U14708 (N_14708,N_14618,N_14581);
nand U14709 (N_14709,N_14668,N_14653);
or U14710 (N_14710,N_14595,N_14578);
or U14711 (N_14711,N_14644,N_14648);
nand U14712 (N_14712,N_14647,N_14606);
and U14713 (N_14713,N_14635,N_14665);
xor U14714 (N_14714,N_14599,N_14654);
nor U14715 (N_14715,N_14646,N_14630);
xnor U14716 (N_14716,N_14558,N_14637);
xnor U14717 (N_14717,N_14604,N_14569);
or U14718 (N_14718,N_14610,N_14592);
nand U14719 (N_14719,N_14674,N_14615);
nand U14720 (N_14720,N_14664,N_14591);
xnor U14721 (N_14721,N_14667,N_14628);
nand U14722 (N_14722,N_14572,N_14690);
xnor U14723 (N_14723,N_14634,N_14680);
nor U14724 (N_14724,N_14621,N_14689);
or U14725 (N_14725,N_14682,N_14657);
or U14726 (N_14726,N_14641,N_14565);
xnor U14727 (N_14727,N_14554,N_14583);
xor U14728 (N_14728,N_14669,N_14666);
nor U14729 (N_14729,N_14602,N_14656);
or U14730 (N_14730,N_14652,N_14584);
xor U14731 (N_14731,N_14691,N_14608);
nand U14732 (N_14732,N_14624,N_14622);
xnor U14733 (N_14733,N_14629,N_14623);
nor U14734 (N_14734,N_14676,N_14645);
nand U14735 (N_14735,N_14582,N_14631);
or U14736 (N_14736,N_14553,N_14580);
xor U14737 (N_14737,N_14579,N_14686);
nor U14738 (N_14738,N_14589,N_14679);
xnor U14739 (N_14739,N_14632,N_14642);
or U14740 (N_14740,N_14574,N_14566);
xor U14741 (N_14741,N_14673,N_14614);
xor U14742 (N_14742,N_14658,N_14672);
nor U14743 (N_14743,N_14626,N_14585);
xnor U14744 (N_14744,N_14586,N_14587);
xor U14745 (N_14745,N_14611,N_14601);
or U14746 (N_14746,N_14678,N_14697);
nand U14747 (N_14747,N_14681,N_14597);
nor U14748 (N_14748,N_14564,N_14557);
xor U14749 (N_14749,N_14627,N_14651);
nand U14750 (N_14750,N_14692,N_14675);
or U14751 (N_14751,N_14567,N_14638);
nor U14752 (N_14752,N_14590,N_14685);
nand U14753 (N_14753,N_14573,N_14693);
or U14754 (N_14754,N_14684,N_14695);
and U14755 (N_14755,N_14688,N_14552);
or U14756 (N_14756,N_14570,N_14649);
nand U14757 (N_14757,N_14677,N_14594);
or U14758 (N_14758,N_14696,N_14694);
or U14759 (N_14759,N_14598,N_14575);
nand U14760 (N_14760,N_14639,N_14612);
and U14761 (N_14761,N_14661,N_14636);
nand U14762 (N_14762,N_14559,N_14550);
xnor U14763 (N_14763,N_14670,N_14662);
nor U14764 (N_14764,N_14576,N_14663);
or U14765 (N_14765,N_14588,N_14650);
xor U14766 (N_14766,N_14659,N_14616);
nor U14767 (N_14767,N_14551,N_14655);
xnor U14768 (N_14768,N_14660,N_14683);
and U14769 (N_14769,N_14600,N_14563);
nor U14770 (N_14770,N_14613,N_14577);
or U14771 (N_14771,N_14619,N_14593);
nand U14772 (N_14772,N_14617,N_14620);
and U14773 (N_14773,N_14671,N_14555);
or U14774 (N_14774,N_14562,N_14687);
nor U14775 (N_14775,N_14654,N_14660);
nor U14776 (N_14776,N_14692,N_14624);
or U14777 (N_14777,N_14669,N_14611);
nand U14778 (N_14778,N_14590,N_14665);
or U14779 (N_14779,N_14619,N_14687);
or U14780 (N_14780,N_14698,N_14670);
nor U14781 (N_14781,N_14563,N_14644);
nand U14782 (N_14782,N_14577,N_14606);
or U14783 (N_14783,N_14646,N_14672);
nand U14784 (N_14784,N_14637,N_14554);
and U14785 (N_14785,N_14604,N_14687);
and U14786 (N_14786,N_14580,N_14646);
nand U14787 (N_14787,N_14623,N_14683);
nor U14788 (N_14788,N_14606,N_14601);
or U14789 (N_14789,N_14656,N_14556);
or U14790 (N_14790,N_14658,N_14576);
nor U14791 (N_14791,N_14637,N_14569);
nor U14792 (N_14792,N_14569,N_14652);
xor U14793 (N_14793,N_14592,N_14611);
xnor U14794 (N_14794,N_14556,N_14695);
xor U14795 (N_14795,N_14672,N_14679);
xnor U14796 (N_14796,N_14566,N_14587);
nor U14797 (N_14797,N_14619,N_14648);
and U14798 (N_14798,N_14622,N_14652);
nor U14799 (N_14799,N_14603,N_14686);
xor U14800 (N_14800,N_14698,N_14634);
or U14801 (N_14801,N_14563,N_14590);
and U14802 (N_14802,N_14600,N_14676);
xnor U14803 (N_14803,N_14592,N_14585);
and U14804 (N_14804,N_14581,N_14554);
nor U14805 (N_14805,N_14569,N_14621);
or U14806 (N_14806,N_14697,N_14691);
xor U14807 (N_14807,N_14564,N_14692);
xnor U14808 (N_14808,N_14650,N_14602);
nand U14809 (N_14809,N_14631,N_14565);
and U14810 (N_14810,N_14691,N_14666);
or U14811 (N_14811,N_14592,N_14640);
nand U14812 (N_14812,N_14605,N_14615);
and U14813 (N_14813,N_14652,N_14673);
nor U14814 (N_14814,N_14586,N_14678);
or U14815 (N_14815,N_14621,N_14615);
nor U14816 (N_14816,N_14602,N_14555);
nand U14817 (N_14817,N_14690,N_14566);
and U14818 (N_14818,N_14644,N_14673);
or U14819 (N_14819,N_14619,N_14686);
nand U14820 (N_14820,N_14655,N_14649);
xor U14821 (N_14821,N_14561,N_14571);
xor U14822 (N_14822,N_14686,N_14574);
nand U14823 (N_14823,N_14613,N_14630);
nand U14824 (N_14824,N_14570,N_14600);
nand U14825 (N_14825,N_14662,N_14584);
and U14826 (N_14826,N_14613,N_14698);
nor U14827 (N_14827,N_14579,N_14565);
nor U14828 (N_14828,N_14699,N_14645);
or U14829 (N_14829,N_14667,N_14555);
and U14830 (N_14830,N_14646,N_14582);
or U14831 (N_14831,N_14653,N_14664);
and U14832 (N_14832,N_14611,N_14589);
xnor U14833 (N_14833,N_14558,N_14652);
xor U14834 (N_14834,N_14610,N_14673);
nand U14835 (N_14835,N_14661,N_14617);
nor U14836 (N_14836,N_14685,N_14667);
xnor U14837 (N_14837,N_14627,N_14665);
or U14838 (N_14838,N_14569,N_14602);
xnor U14839 (N_14839,N_14556,N_14564);
nand U14840 (N_14840,N_14683,N_14599);
nor U14841 (N_14841,N_14597,N_14645);
nor U14842 (N_14842,N_14693,N_14561);
nor U14843 (N_14843,N_14552,N_14663);
xor U14844 (N_14844,N_14613,N_14597);
nand U14845 (N_14845,N_14647,N_14631);
xnor U14846 (N_14846,N_14673,N_14667);
or U14847 (N_14847,N_14579,N_14566);
or U14848 (N_14848,N_14637,N_14563);
nand U14849 (N_14849,N_14678,N_14683);
nand U14850 (N_14850,N_14755,N_14711);
or U14851 (N_14851,N_14709,N_14716);
and U14852 (N_14852,N_14790,N_14802);
nand U14853 (N_14853,N_14777,N_14704);
nor U14854 (N_14854,N_14813,N_14756);
or U14855 (N_14855,N_14706,N_14730);
and U14856 (N_14856,N_14783,N_14771);
or U14857 (N_14857,N_14788,N_14846);
nor U14858 (N_14858,N_14710,N_14837);
and U14859 (N_14859,N_14816,N_14735);
or U14860 (N_14860,N_14833,N_14829);
and U14861 (N_14861,N_14726,N_14824);
or U14862 (N_14862,N_14724,N_14725);
xnor U14863 (N_14863,N_14809,N_14845);
and U14864 (N_14864,N_14791,N_14843);
nand U14865 (N_14865,N_14848,N_14807);
nor U14866 (N_14866,N_14737,N_14733);
or U14867 (N_14867,N_14789,N_14750);
nand U14868 (N_14868,N_14826,N_14804);
and U14869 (N_14869,N_14743,N_14740);
nand U14870 (N_14870,N_14715,N_14774);
xnor U14871 (N_14871,N_14708,N_14701);
and U14872 (N_14872,N_14792,N_14717);
nand U14873 (N_14873,N_14799,N_14723);
nor U14874 (N_14874,N_14794,N_14759);
nor U14875 (N_14875,N_14738,N_14842);
nand U14876 (N_14876,N_14747,N_14830);
nand U14877 (N_14877,N_14705,N_14836);
xnor U14878 (N_14878,N_14764,N_14754);
xor U14879 (N_14879,N_14834,N_14731);
nor U14880 (N_14880,N_14827,N_14782);
nor U14881 (N_14881,N_14838,N_14806);
or U14882 (N_14882,N_14812,N_14766);
nor U14883 (N_14883,N_14796,N_14840);
nand U14884 (N_14884,N_14748,N_14803);
and U14885 (N_14885,N_14793,N_14815);
xor U14886 (N_14886,N_14784,N_14721);
xor U14887 (N_14887,N_14780,N_14787);
and U14888 (N_14888,N_14847,N_14811);
nand U14889 (N_14889,N_14767,N_14739);
and U14890 (N_14890,N_14772,N_14700);
or U14891 (N_14891,N_14720,N_14745);
or U14892 (N_14892,N_14768,N_14746);
or U14893 (N_14893,N_14734,N_14757);
or U14894 (N_14894,N_14763,N_14817);
nand U14895 (N_14895,N_14823,N_14729);
and U14896 (N_14896,N_14736,N_14810);
or U14897 (N_14897,N_14832,N_14814);
nand U14898 (N_14898,N_14801,N_14714);
and U14899 (N_14899,N_14785,N_14831);
xor U14900 (N_14900,N_14707,N_14722);
nor U14901 (N_14901,N_14713,N_14775);
nand U14902 (N_14902,N_14835,N_14800);
nand U14903 (N_14903,N_14744,N_14822);
xor U14904 (N_14904,N_14718,N_14778);
and U14905 (N_14905,N_14727,N_14769);
and U14906 (N_14906,N_14765,N_14805);
and U14907 (N_14907,N_14741,N_14712);
or U14908 (N_14908,N_14761,N_14770);
nand U14909 (N_14909,N_14844,N_14742);
nand U14910 (N_14910,N_14808,N_14732);
and U14911 (N_14911,N_14751,N_14821);
and U14912 (N_14912,N_14752,N_14839);
nand U14913 (N_14913,N_14818,N_14749);
nor U14914 (N_14914,N_14702,N_14825);
and U14915 (N_14915,N_14828,N_14798);
or U14916 (N_14916,N_14786,N_14820);
and U14917 (N_14917,N_14849,N_14797);
xnor U14918 (N_14918,N_14781,N_14773);
xnor U14919 (N_14919,N_14753,N_14703);
xor U14920 (N_14920,N_14762,N_14779);
xnor U14921 (N_14921,N_14760,N_14719);
nor U14922 (N_14922,N_14795,N_14776);
nand U14923 (N_14923,N_14758,N_14841);
and U14924 (N_14924,N_14728,N_14819);
nor U14925 (N_14925,N_14710,N_14827);
or U14926 (N_14926,N_14757,N_14741);
nor U14927 (N_14927,N_14836,N_14834);
nor U14928 (N_14928,N_14776,N_14705);
and U14929 (N_14929,N_14820,N_14798);
or U14930 (N_14930,N_14716,N_14824);
and U14931 (N_14931,N_14777,N_14831);
or U14932 (N_14932,N_14764,N_14745);
xnor U14933 (N_14933,N_14707,N_14710);
or U14934 (N_14934,N_14823,N_14811);
xor U14935 (N_14935,N_14730,N_14714);
and U14936 (N_14936,N_14797,N_14807);
nor U14937 (N_14937,N_14707,N_14816);
and U14938 (N_14938,N_14839,N_14791);
xor U14939 (N_14939,N_14738,N_14748);
or U14940 (N_14940,N_14715,N_14710);
nand U14941 (N_14941,N_14810,N_14717);
xor U14942 (N_14942,N_14847,N_14755);
or U14943 (N_14943,N_14797,N_14821);
xor U14944 (N_14944,N_14755,N_14831);
xnor U14945 (N_14945,N_14723,N_14735);
nor U14946 (N_14946,N_14714,N_14716);
nor U14947 (N_14947,N_14797,N_14711);
nand U14948 (N_14948,N_14710,N_14774);
nand U14949 (N_14949,N_14742,N_14779);
and U14950 (N_14950,N_14778,N_14731);
xnor U14951 (N_14951,N_14722,N_14751);
xor U14952 (N_14952,N_14808,N_14812);
nor U14953 (N_14953,N_14834,N_14712);
nor U14954 (N_14954,N_14741,N_14754);
nand U14955 (N_14955,N_14739,N_14723);
xor U14956 (N_14956,N_14730,N_14838);
nand U14957 (N_14957,N_14750,N_14847);
or U14958 (N_14958,N_14773,N_14759);
and U14959 (N_14959,N_14716,N_14728);
or U14960 (N_14960,N_14735,N_14756);
nand U14961 (N_14961,N_14752,N_14843);
or U14962 (N_14962,N_14728,N_14706);
and U14963 (N_14963,N_14844,N_14756);
or U14964 (N_14964,N_14717,N_14843);
xor U14965 (N_14965,N_14715,N_14806);
xor U14966 (N_14966,N_14849,N_14794);
or U14967 (N_14967,N_14721,N_14716);
nor U14968 (N_14968,N_14823,N_14798);
nor U14969 (N_14969,N_14703,N_14748);
and U14970 (N_14970,N_14751,N_14767);
or U14971 (N_14971,N_14849,N_14782);
nor U14972 (N_14972,N_14718,N_14711);
or U14973 (N_14973,N_14710,N_14753);
xnor U14974 (N_14974,N_14714,N_14773);
xor U14975 (N_14975,N_14796,N_14845);
nor U14976 (N_14976,N_14715,N_14777);
and U14977 (N_14977,N_14834,N_14718);
nand U14978 (N_14978,N_14780,N_14722);
and U14979 (N_14979,N_14710,N_14731);
xor U14980 (N_14980,N_14751,N_14719);
or U14981 (N_14981,N_14774,N_14760);
xor U14982 (N_14982,N_14835,N_14830);
nand U14983 (N_14983,N_14784,N_14846);
and U14984 (N_14984,N_14727,N_14829);
nand U14985 (N_14985,N_14831,N_14774);
or U14986 (N_14986,N_14784,N_14761);
nor U14987 (N_14987,N_14701,N_14776);
xnor U14988 (N_14988,N_14821,N_14710);
or U14989 (N_14989,N_14843,N_14811);
and U14990 (N_14990,N_14726,N_14794);
nand U14991 (N_14991,N_14814,N_14737);
nand U14992 (N_14992,N_14811,N_14819);
nor U14993 (N_14993,N_14716,N_14777);
xnor U14994 (N_14994,N_14763,N_14748);
nand U14995 (N_14995,N_14817,N_14754);
and U14996 (N_14996,N_14792,N_14805);
xnor U14997 (N_14997,N_14798,N_14728);
or U14998 (N_14998,N_14823,N_14713);
nand U14999 (N_14999,N_14813,N_14703);
nor UO_0 (O_0,N_14869,N_14929);
nand UO_1 (O_1,N_14912,N_14985);
or UO_2 (O_2,N_14925,N_14961);
nor UO_3 (O_3,N_14955,N_14997);
or UO_4 (O_4,N_14851,N_14906);
xor UO_5 (O_5,N_14882,N_14922);
nor UO_6 (O_6,N_14893,N_14910);
nand UO_7 (O_7,N_14953,N_14965);
xnor UO_8 (O_8,N_14939,N_14887);
and UO_9 (O_9,N_14948,N_14870);
xnor UO_10 (O_10,N_14987,N_14917);
nor UO_11 (O_11,N_14931,N_14940);
and UO_12 (O_12,N_14962,N_14899);
xor UO_13 (O_13,N_14990,N_14976);
or UO_14 (O_14,N_14889,N_14991);
or UO_15 (O_15,N_14969,N_14850);
and UO_16 (O_16,N_14919,N_14937);
or UO_17 (O_17,N_14968,N_14949);
and UO_18 (O_18,N_14879,N_14943);
and UO_19 (O_19,N_14909,N_14905);
xor UO_20 (O_20,N_14945,N_14902);
nand UO_21 (O_21,N_14914,N_14880);
and UO_22 (O_22,N_14983,N_14868);
and UO_23 (O_23,N_14999,N_14863);
nand UO_24 (O_24,N_14954,N_14957);
and UO_25 (O_25,N_14876,N_14977);
nor UO_26 (O_26,N_14970,N_14856);
or UO_27 (O_27,N_14926,N_14938);
nand UO_28 (O_28,N_14988,N_14854);
nand UO_29 (O_29,N_14871,N_14892);
xnor UO_30 (O_30,N_14900,N_14908);
nor UO_31 (O_31,N_14951,N_14916);
nor UO_32 (O_32,N_14875,N_14979);
or UO_33 (O_33,N_14975,N_14858);
nand UO_34 (O_34,N_14982,N_14867);
xor UO_35 (O_35,N_14959,N_14878);
nand UO_36 (O_36,N_14932,N_14896);
and UO_37 (O_37,N_14915,N_14927);
and UO_38 (O_38,N_14862,N_14956);
nand UO_39 (O_39,N_14860,N_14861);
and UO_40 (O_40,N_14884,N_14903);
nand UO_41 (O_41,N_14980,N_14964);
xor UO_42 (O_42,N_14942,N_14859);
nand UO_43 (O_43,N_14907,N_14958);
xor UO_44 (O_44,N_14874,N_14857);
nand UO_45 (O_45,N_14911,N_14890);
xnor UO_46 (O_46,N_14974,N_14895);
nand UO_47 (O_47,N_14978,N_14885);
and UO_48 (O_48,N_14941,N_14888);
nand UO_49 (O_49,N_14981,N_14947);
xnor UO_50 (O_50,N_14992,N_14986);
nand UO_51 (O_51,N_14883,N_14973);
and UO_52 (O_52,N_14994,N_14898);
or UO_53 (O_53,N_14936,N_14989);
nor UO_54 (O_54,N_14891,N_14894);
nand UO_55 (O_55,N_14934,N_14877);
and UO_56 (O_56,N_14855,N_14852);
or UO_57 (O_57,N_14853,N_14864);
nand UO_58 (O_58,N_14966,N_14967);
nand UO_59 (O_59,N_14972,N_14935);
nand UO_60 (O_60,N_14993,N_14995);
or UO_61 (O_61,N_14918,N_14901);
nor UO_62 (O_62,N_14950,N_14971);
nor UO_63 (O_63,N_14881,N_14933);
and UO_64 (O_64,N_14998,N_14873);
and UO_65 (O_65,N_14924,N_14930);
xnor UO_66 (O_66,N_14920,N_14996);
and UO_67 (O_67,N_14952,N_14960);
and UO_68 (O_68,N_14866,N_14904);
and UO_69 (O_69,N_14865,N_14913);
and UO_70 (O_70,N_14928,N_14963);
nand UO_71 (O_71,N_14921,N_14897);
nand UO_72 (O_72,N_14886,N_14944);
and UO_73 (O_73,N_14872,N_14923);
xor UO_74 (O_74,N_14946,N_14984);
nand UO_75 (O_75,N_14931,N_14988);
nor UO_76 (O_76,N_14887,N_14892);
nand UO_77 (O_77,N_14873,N_14910);
or UO_78 (O_78,N_14869,N_14906);
nand UO_79 (O_79,N_14961,N_14878);
and UO_80 (O_80,N_14940,N_14894);
or UO_81 (O_81,N_14960,N_14908);
and UO_82 (O_82,N_14984,N_14961);
nor UO_83 (O_83,N_14983,N_14972);
nand UO_84 (O_84,N_14963,N_14940);
or UO_85 (O_85,N_14913,N_14961);
or UO_86 (O_86,N_14995,N_14921);
and UO_87 (O_87,N_14886,N_14870);
nand UO_88 (O_88,N_14918,N_14948);
and UO_89 (O_89,N_14897,N_14862);
nor UO_90 (O_90,N_14903,N_14969);
nand UO_91 (O_91,N_14982,N_14906);
nand UO_92 (O_92,N_14897,N_14983);
nor UO_93 (O_93,N_14967,N_14935);
nor UO_94 (O_94,N_14942,N_14879);
nor UO_95 (O_95,N_14851,N_14913);
nor UO_96 (O_96,N_14855,N_14908);
nor UO_97 (O_97,N_14964,N_14995);
nand UO_98 (O_98,N_14907,N_14972);
and UO_99 (O_99,N_14868,N_14870);
nand UO_100 (O_100,N_14852,N_14909);
nand UO_101 (O_101,N_14928,N_14926);
xor UO_102 (O_102,N_14948,N_14882);
nand UO_103 (O_103,N_14903,N_14906);
or UO_104 (O_104,N_14882,N_14903);
nand UO_105 (O_105,N_14903,N_14995);
xor UO_106 (O_106,N_14947,N_14878);
nand UO_107 (O_107,N_14860,N_14871);
nand UO_108 (O_108,N_14905,N_14916);
nand UO_109 (O_109,N_14867,N_14977);
nor UO_110 (O_110,N_14862,N_14977);
nor UO_111 (O_111,N_14922,N_14935);
nor UO_112 (O_112,N_14946,N_14855);
and UO_113 (O_113,N_14995,N_14878);
or UO_114 (O_114,N_14863,N_14910);
nor UO_115 (O_115,N_14978,N_14956);
or UO_116 (O_116,N_14961,N_14896);
or UO_117 (O_117,N_14961,N_14900);
nand UO_118 (O_118,N_14893,N_14972);
xor UO_119 (O_119,N_14942,N_14893);
or UO_120 (O_120,N_14979,N_14990);
xor UO_121 (O_121,N_14952,N_14890);
xor UO_122 (O_122,N_14912,N_14966);
and UO_123 (O_123,N_14866,N_14886);
or UO_124 (O_124,N_14929,N_14952);
and UO_125 (O_125,N_14949,N_14853);
xnor UO_126 (O_126,N_14886,N_14941);
or UO_127 (O_127,N_14953,N_14876);
and UO_128 (O_128,N_14920,N_14936);
nand UO_129 (O_129,N_14955,N_14910);
nor UO_130 (O_130,N_14879,N_14885);
nor UO_131 (O_131,N_14951,N_14939);
and UO_132 (O_132,N_14950,N_14875);
or UO_133 (O_133,N_14866,N_14874);
xor UO_134 (O_134,N_14897,N_14959);
nand UO_135 (O_135,N_14894,N_14961);
or UO_136 (O_136,N_14893,N_14990);
nor UO_137 (O_137,N_14938,N_14984);
xnor UO_138 (O_138,N_14976,N_14926);
xor UO_139 (O_139,N_14934,N_14913);
nand UO_140 (O_140,N_14969,N_14869);
and UO_141 (O_141,N_14898,N_14978);
xnor UO_142 (O_142,N_14889,N_14947);
nor UO_143 (O_143,N_14878,N_14953);
xor UO_144 (O_144,N_14964,N_14918);
or UO_145 (O_145,N_14956,N_14894);
nand UO_146 (O_146,N_14945,N_14946);
nor UO_147 (O_147,N_14861,N_14994);
nor UO_148 (O_148,N_14976,N_14935);
xnor UO_149 (O_149,N_14958,N_14979);
nor UO_150 (O_150,N_14908,N_14954);
nand UO_151 (O_151,N_14913,N_14864);
xnor UO_152 (O_152,N_14933,N_14948);
nor UO_153 (O_153,N_14895,N_14920);
nor UO_154 (O_154,N_14926,N_14882);
or UO_155 (O_155,N_14951,N_14925);
and UO_156 (O_156,N_14971,N_14872);
xor UO_157 (O_157,N_14887,N_14969);
and UO_158 (O_158,N_14955,N_14948);
nand UO_159 (O_159,N_14908,N_14901);
nor UO_160 (O_160,N_14886,N_14900);
nand UO_161 (O_161,N_14989,N_14913);
nand UO_162 (O_162,N_14859,N_14923);
nor UO_163 (O_163,N_14965,N_14882);
xnor UO_164 (O_164,N_14999,N_14876);
or UO_165 (O_165,N_14898,N_14857);
or UO_166 (O_166,N_14934,N_14942);
nand UO_167 (O_167,N_14854,N_14884);
or UO_168 (O_168,N_14932,N_14945);
and UO_169 (O_169,N_14922,N_14916);
nand UO_170 (O_170,N_14939,N_14999);
xor UO_171 (O_171,N_14974,N_14882);
and UO_172 (O_172,N_14871,N_14955);
and UO_173 (O_173,N_14909,N_14860);
nand UO_174 (O_174,N_14959,N_14908);
and UO_175 (O_175,N_14870,N_14874);
nand UO_176 (O_176,N_14979,N_14884);
xnor UO_177 (O_177,N_14980,N_14859);
xnor UO_178 (O_178,N_14979,N_14942);
xnor UO_179 (O_179,N_14984,N_14915);
nor UO_180 (O_180,N_14959,N_14998);
or UO_181 (O_181,N_14899,N_14991);
and UO_182 (O_182,N_14935,N_14957);
nand UO_183 (O_183,N_14881,N_14915);
or UO_184 (O_184,N_14888,N_14950);
or UO_185 (O_185,N_14863,N_14902);
nor UO_186 (O_186,N_14997,N_14977);
or UO_187 (O_187,N_14860,N_14930);
xor UO_188 (O_188,N_14882,N_14864);
nor UO_189 (O_189,N_14885,N_14984);
xnor UO_190 (O_190,N_14914,N_14994);
and UO_191 (O_191,N_14857,N_14967);
xnor UO_192 (O_192,N_14930,N_14925);
and UO_193 (O_193,N_14932,N_14863);
xor UO_194 (O_194,N_14911,N_14936);
and UO_195 (O_195,N_14982,N_14952);
nand UO_196 (O_196,N_14916,N_14987);
xnor UO_197 (O_197,N_14995,N_14897);
or UO_198 (O_198,N_14873,N_14969);
xor UO_199 (O_199,N_14966,N_14904);
and UO_200 (O_200,N_14868,N_14873);
nor UO_201 (O_201,N_14870,N_14904);
nand UO_202 (O_202,N_14918,N_14859);
xnor UO_203 (O_203,N_14999,N_14972);
and UO_204 (O_204,N_14882,N_14968);
nor UO_205 (O_205,N_14999,N_14953);
and UO_206 (O_206,N_14869,N_14945);
or UO_207 (O_207,N_14859,N_14959);
or UO_208 (O_208,N_14936,N_14951);
nor UO_209 (O_209,N_14898,N_14860);
nand UO_210 (O_210,N_14938,N_14865);
or UO_211 (O_211,N_14913,N_14899);
or UO_212 (O_212,N_14967,N_14958);
or UO_213 (O_213,N_14917,N_14991);
xor UO_214 (O_214,N_14930,N_14978);
nand UO_215 (O_215,N_14962,N_14926);
and UO_216 (O_216,N_14931,N_14976);
xnor UO_217 (O_217,N_14994,N_14964);
and UO_218 (O_218,N_14947,N_14965);
nand UO_219 (O_219,N_14897,N_14987);
nor UO_220 (O_220,N_14963,N_14995);
nor UO_221 (O_221,N_14895,N_14980);
nand UO_222 (O_222,N_14961,N_14980);
xnor UO_223 (O_223,N_14902,N_14955);
or UO_224 (O_224,N_14885,N_14882);
and UO_225 (O_225,N_14977,N_14866);
nor UO_226 (O_226,N_14927,N_14890);
and UO_227 (O_227,N_14877,N_14931);
xnor UO_228 (O_228,N_14966,N_14985);
and UO_229 (O_229,N_14935,N_14855);
xor UO_230 (O_230,N_14997,N_14887);
or UO_231 (O_231,N_14913,N_14892);
and UO_232 (O_232,N_14980,N_14887);
nand UO_233 (O_233,N_14902,N_14908);
or UO_234 (O_234,N_14998,N_14922);
xor UO_235 (O_235,N_14873,N_14883);
nand UO_236 (O_236,N_14922,N_14860);
or UO_237 (O_237,N_14905,N_14927);
nand UO_238 (O_238,N_14895,N_14898);
nand UO_239 (O_239,N_14976,N_14995);
xnor UO_240 (O_240,N_14922,N_14927);
nand UO_241 (O_241,N_14961,N_14928);
nor UO_242 (O_242,N_14858,N_14875);
or UO_243 (O_243,N_14864,N_14859);
and UO_244 (O_244,N_14902,N_14986);
nand UO_245 (O_245,N_14929,N_14973);
nor UO_246 (O_246,N_14948,N_14860);
and UO_247 (O_247,N_14961,N_14869);
or UO_248 (O_248,N_14910,N_14853);
nor UO_249 (O_249,N_14867,N_14956);
xnor UO_250 (O_250,N_14989,N_14979);
or UO_251 (O_251,N_14976,N_14971);
or UO_252 (O_252,N_14904,N_14913);
xor UO_253 (O_253,N_14950,N_14942);
xnor UO_254 (O_254,N_14866,N_14927);
nand UO_255 (O_255,N_14941,N_14952);
xnor UO_256 (O_256,N_14894,N_14887);
nand UO_257 (O_257,N_14971,N_14866);
xor UO_258 (O_258,N_14979,N_14951);
xor UO_259 (O_259,N_14988,N_14933);
nor UO_260 (O_260,N_14977,N_14883);
nor UO_261 (O_261,N_14915,N_14951);
nor UO_262 (O_262,N_14987,N_14928);
xor UO_263 (O_263,N_14906,N_14899);
and UO_264 (O_264,N_14924,N_14929);
xor UO_265 (O_265,N_14922,N_14951);
and UO_266 (O_266,N_14877,N_14969);
xor UO_267 (O_267,N_14877,N_14869);
xnor UO_268 (O_268,N_14970,N_14946);
nand UO_269 (O_269,N_14957,N_14984);
nand UO_270 (O_270,N_14906,N_14908);
xnor UO_271 (O_271,N_14988,N_14957);
nand UO_272 (O_272,N_14923,N_14868);
and UO_273 (O_273,N_14852,N_14928);
xor UO_274 (O_274,N_14945,N_14989);
nor UO_275 (O_275,N_14950,N_14880);
xor UO_276 (O_276,N_14886,N_14854);
nand UO_277 (O_277,N_14990,N_14942);
nor UO_278 (O_278,N_14911,N_14986);
nand UO_279 (O_279,N_14945,N_14915);
nand UO_280 (O_280,N_14988,N_14940);
xor UO_281 (O_281,N_14859,N_14919);
and UO_282 (O_282,N_14926,N_14934);
and UO_283 (O_283,N_14857,N_14969);
and UO_284 (O_284,N_14949,N_14892);
and UO_285 (O_285,N_14908,N_14858);
nor UO_286 (O_286,N_14954,N_14850);
xnor UO_287 (O_287,N_14905,N_14947);
nand UO_288 (O_288,N_14986,N_14883);
nand UO_289 (O_289,N_14956,N_14857);
and UO_290 (O_290,N_14965,N_14961);
and UO_291 (O_291,N_14957,N_14982);
nand UO_292 (O_292,N_14885,N_14977);
nor UO_293 (O_293,N_14945,N_14883);
nand UO_294 (O_294,N_14925,N_14919);
or UO_295 (O_295,N_14932,N_14858);
and UO_296 (O_296,N_14885,N_14914);
xor UO_297 (O_297,N_14984,N_14951);
nand UO_298 (O_298,N_14879,N_14915);
xor UO_299 (O_299,N_14859,N_14978);
xnor UO_300 (O_300,N_14982,N_14903);
nand UO_301 (O_301,N_14930,N_14996);
nor UO_302 (O_302,N_14959,N_14852);
and UO_303 (O_303,N_14987,N_14941);
nand UO_304 (O_304,N_14874,N_14917);
and UO_305 (O_305,N_14939,N_14987);
and UO_306 (O_306,N_14896,N_14897);
nand UO_307 (O_307,N_14968,N_14855);
xnor UO_308 (O_308,N_14896,N_14871);
or UO_309 (O_309,N_14960,N_14965);
nor UO_310 (O_310,N_14970,N_14933);
or UO_311 (O_311,N_14917,N_14907);
or UO_312 (O_312,N_14909,N_14929);
or UO_313 (O_313,N_14858,N_14931);
and UO_314 (O_314,N_14920,N_14908);
nor UO_315 (O_315,N_14895,N_14853);
nor UO_316 (O_316,N_14895,N_14937);
nand UO_317 (O_317,N_14987,N_14860);
xor UO_318 (O_318,N_14927,N_14884);
xor UO_319 (O_319,N_14979,N_14902);
and UO_320 (O_320,N_14907,N_14895);
nand UO_321 (O_321,N_14960,N_14999);
nand UO_322 (O_322,N_14904,N_14890);
nand UO_323 (O_323,N_14910,N_14871);
nor UO_324 (O_324,N_14979,N_14856);
and UO_325 (O_325,N_14886,N_14968);
or UO_326 (O_326,N_14875,N_14933);
and UO_327 (O_327,N_14902,N_14997);
and UO_328 (O_328,N_14897,N_14927);
or UO_329 (O_329,N_14993,N_14877);
and UO_330 (O_330,N_14927,N_14857);
or UO_331 (O_331,N_14981,N_14990);
nand UO_332 (O_332,N_14952,N_14851);
xor UO_333 (O_333,N_14915,N_14985);
or UO_334 (O_334,N_14906,N_14966);
nand UO_335 (O_335,N_14890,N_14866);
nor UO_336 (O_336,N_14949,N_14980);
xnor UO_337 (O_337,N_14970,N_14901);
xnor UO_338 (O_338,N_14905,N_14878);
xnor UO_339 (O_339,N_14855,N_14980);
or UO_340 (O_340,N_14917,N_14936);
nor UO_341 (O_341,N_14974,N_14918);
xnor UO_342 (O_342,N_14996,N_14850);
and UO_343 (O_343,N_14910,N_14902);
or UO_344 (O_344,N_14871,N_14943);
nor UO_345 (O_345,N_14997,N_14850);
and UO_346 (O_346,N_14998,N_14966);
nor UO_347 (O_347,N_14935,N_14958);
or UO_348 (O_348,N_14982,N_14917);
nor UO_349 (O_349,N_14946,N_14980);
and UO_350 (O_350,N_14902,N_14881);
nor UO_351 (O_351,N_14878,N_14999);
nor UO_352 (O_352,N_14998,N_14917);
nor UO_353 (O_353,N_14885,N_14940);
and UO_354 (O_354,N_14979,N_14967);
or UO_355 (O_355,N_14921,N_14982);
and UO_356 (O_356,N_14855,N_14970);
or UO_357 (O_357,N_14878,N_14850);
and UO_358 (O_358,N_14900,N_14872);
nor UO_359 (O_359,N_14948,N_14876);
nor UO_360 (O_360,N_14958,N_14994);
nand UO_361 (O_361,N_14910,N_14896);
xnor UO_362 (O_362,N_14930,N_14934);
nor UO_363 (O_363,N_14914,N_14981);
and UO_364 (O_364,N_14918,N_14851);
xor UO_365 (O_365,N_14962,N_14880);
or UO_366 (O_366,N_14859,N_14975);
nor UO_367 (O_367,N_14933,N_14931);
nand UO_368 (O_368,N_14861,N_14960);
xnor UO_369 (O_369,N_14887,N_14877);
xor UO_370 (O_370,N_14995,N_14885);
and UO_371 (O_371,N_14934,N_14904);
and UO_372 (O_372,N_14915,N_14919);
nor UO_373 (O_373,N_14911,N_14963);
or UO_374 (O_374,N_14996,N_14882);
xor UO_375 (O_375,N_14982,N_14931);
or UO_376 (O_376,N_14933,N_14919);
xor UO_377 (O_377,N_14883,N_14937);
xnor UO_378 (O_378,N_14946,N_14903);
and UO_379 (O_379,N_14983,N_14992);
nor UO_380 (O_380,N_14955,N_14974);
nor UO_381 (O_381,N_14943,N_14863);
xor UO_382 (O_382,N_14949,N_14864);
and UO_383 (O_383,N_14925,N_14960);
xor UO_384 (O_384,N_14974,N_14980);
nor UO_385 (O_385,N_14937,N_14968);
xor UO_386 (O_386,N_14889,N_14968);
and UO_387 (O_387,N_14939,N_14963);
nand UO_388 (O_388,N_14979,N_14850);
or UO_389 (O_389,N_14948,N_14914);
or UO_390 (O_390,N_14978,N_14974);
and UO_391 (O_391,N_14927,N_14924);
xor UO_392 (O_392,N_14868,N_14901);
or UO_393 (O_393,N_14948,N_14941);
nor UO_394 (O_394,N_14875,N_14925);
nand UO_395 (O_395,N_14895,N_14938);
or UO_396 (O_396,N_14989,N_14867);
nand UO_397 (O_397,N_14895,N_14923);
nand UO_398 (O_398,N_14868,N_14896);
nand UO_399 (O_399,N_14898,N_14977);
xnor UO_400 (O_400,N_14897,N_14871);
nor UO_401 (O_401,N_14999,N_14992);
or UO_402 (O_402,N_14914,N_14954);
xor UO_403 (O_403,N_14961,N_14861);
or UO_404 (O_404,N_14867,N_14889);
xnor UO_405 (O_405,N_14878,N_14889);
and UO_406 (O_406,N_14947,N_14977);
nand UO_407 (O_407,N_14918,N_14984);
nor UO_408 (O_408,N_14979,N_14853);
nor UO_409 (O_409,N_14887,N_14941);
or UO_410 (O_410,N_14856,N_14932);
or UO_411 (O_411,N_14911,N_14994);
nand UO_412 (O_412,N_14998,N_14947);
nor UO_413 (O_413,N_14981,N_14903);
xor UO_414 (O_414,N_14921,N_14972);
and UO_415 (O_415,N_14851,N_14938);
nand UO_416 (O_416,N_14853,N_14926);
or UO_417 (O_417,N_14982,N_14891);
nor UO_418 (O_418,N_14894,N_14853);
nor UO_419 (O_419,N_14902,N_14977);
nor UO_420 (O_420,N_14905,N_14854);
or UO_421 (O_421,N_14949,N_14925);
and UO_422 (O_422,N_14920,N_14930);
and UO_423 (O_423,N_14973,N_14903);
xor UO_424 (O_424,N_14927,N_14981);
and UO_425 (O_425,N_14877,N_14868);
xnor UO_426 (O_426,N_14988,N_14946);
or UO_427 (O_427,N_14981,N_14888);
xor UO_428 (O_428,N_14860,N_14911);
nand UO_429 (O_429,N_14871,N_14909);
nand UO_430 (O_430,N_14866,N_14928);
and UO_431 (O_431,N_14972,N_14932);
xnor UO_432 (O_432,N_14864,N_14989);
nand UO_433 (O_433,N_14952,N_14964);
nor UO_434 (O_434,N_14995,N_14916);
or UO_435 (O_435,N_14991,N_14874);
or UO_436 (O_436,N_14939,N_14903);
nand UO_437 (O_437,N_14889,N_14880);
nand UO_438 (O_438,N_14925,N_14993);
nand UO_439 (O_439,N_14982,N_14936);
nor UO_440 (O_440,N_14946,N_14862);
and UO_441 (O_441,N_14866,N_14896);
nor UO_442 (O_442,N_14900,N_14871);
nor UO_443 (O_443,N_14900,N_14929);
xor UO_444 (O_444,N_14906,N_14897);
and UO_445 (O_445,N_14989,N_14917);
nor UO_446 (O_446,N_14905,N_14855);
and UO_447 (O_447,N_14962,N_14855);
and UO_448 (O_448,N_14921,N_14960);
xnor UO_449 (O_449,N_14857,N_14859);
xor UO_450 (O_450,N_14953,N_14962);
xor UO_451 (O_451,N_14989,N_14855);
nand UO_452 (O_452,N_14964,N_14992);
nand UO_453 (O_453,N_14958,N_14897);
or UO_454 (O_454,N_14941,N_14883);
xor UO_455 (O_455,N_14964,N_14979);
nor UO_456 (O_456,N_14979,N_14888);
or UO_457 (O_457,N_14902,N_14983);
xnor UO_458 (O_458,N_14889,N_14939);
xor UO_459 (O_459,N_14914,N_14979);
xor UO_460 (O_460,N_14866,N_14962);
and UO_461 (O_461,N_14899,N_14971);
and UO_462 (O_462,N_14881,N_14894);
or UO_463 (O_463,N_14917,N_14859);
and UO_464 (O_464,N_14931,N_14942);
xor UO_465 (O_465,N_14984,N_14953);
xnor UO_466 (O_466,N_14923,N_14993);
nor UO_467 (O_467,N_14927,N_14993);
or UO_468 (O_468,N_14948,N_14887);
or UO_469 (O_469,N_14919,N_14875);
xor UO_470 (O_470,N_14968,N_14978);
or UO_471 (O_471,N_14909,N_14882);
xor UO_472 (O_472,N_14854,N_14903);
nand UO_473 (O_473,N_14936,N_14870);
or UO_474 (O_474,N_14852,N_14995);
or UO_475 (O_475,N_14960,N_14852);
xnor UO_476 (O_476,N_14976,N_14966);
nand UO_477 (O_477,N_14994,N_14941);
nand UO_478 (O_478,N_14938,N_14977);
nor UO_479 (O_479,N_14942,N_14907);
nor UO_480 (O_480,N_14889,N_14887);
xor UO_481 (O_481,N_14948,N_14852);
nor UO_482 (O_482,N_14987,N_14970);
nor UO_483 (O_483,N_14971,N_14860);
nor UO_484 (O_484,N_14891,N_14858);
xnor UO_485 (O_485,N_14967,N_14867);
nor UO_486 (O_486,N_14909,N_14916);
and UO_487 (O_487,N_14918,N_14853);
xnor UO_488 (O_488,N_14948,N_14877);
xnor UO_489 (O_489,N_14993,N_14915);
nor UO_490 (O_490,N_14936,N_14855);
or UO_491 (O_491,N_14958,N_14964);
or UO_492 (O_492,N_14904,N_14960);
nor UO_493 (O_493,N_14958,N_14968);
or UO_494 (O_494,N_14865,N_14881);
nand UO_495 (O_495,N_14917,N_14927);
or UO_496 (O_496,N_14998,N_14860);
nor UO_497 (O_497,N_14908,N_14860);
xor UO_498 (O_498,N_14883,N_14895);
xnor UO_499 (O_499,N_14920,N_14890);
xor UO_500 (O_500,N_14968,N_14908);
xnor UO_501 (O_501,N_14940,N_14967);
or UO_502 (O_502,N_14879,N_14993);
xor UO_503 (O_503,N_14980,N_14948);
nor UO_504 (O_504,N_14901,N_14993);
or UO_505 (O_505,N_14934,N_14983);
nand UO_506 (O_506,N_14912,N_14883);
nor UO_507 (O_507,N_14982,N_14873);
or UO_508 (O_508,N_14988,N_14935);
nand UO_509 (O_509,N_14910,N_14890);
and UO_510 (O_510,N_14855,N_14863);
and UO_511 (O_511,N_14879,N_14910);
nor UO_512 (O_512,N_14979,N_14971);
nand UO_513 (O_513,N_14870,N_14896);
and UO_514 (O_514,N_14861,N_14932);
or UO_515 (O_515,N_14898,N_14972);
and UO_516 (O_516,N_14874,N_14983);
and UO_517 (O_517,N_14900,N_14956);
xnor UO_518 (O_518,N_14943,N_14963);
nand UO_519 (O_519,N_14863,N_14961);
nand UO_520 (O_520,N_14872,N_14917);
or UO_521 (O_521,N_14885,N_14930);
and UO_522 (O_522,N_14931,N_14917);
xor UO_523 (O_523,N_14992,N_14862);
xor UO_524 (O_524,N_14928,N_14911);
and UO_525 (O_525,N_14922,N_14924);
nor UO_526 (O_526,N_14872,N_14952);
and UO_527 (O_527,N_14929,N_14964);
nor UO_528 (O_528,N_14967,N_14938);
xnor UO_529 (O_529,N_14876,N_14879);
xnor UO_530 (O_530,N_14945,N_14909);
and UO_531 (O_531,N_14985,N_14968);
or UO_532 (O_532,N_14856,N_14919);
nor UO_533 (O_533,N_14907,N_14871);
nor UO_534 (O_534,N_14929,N_14991);
xor UO_535 (O_535,N_14981,N_14896);
nand UO_536 (O_536,N_14993,N_14898);
or UO_537 (O_537,N_14854,N_14852);
xnor UO_538 (O_538,N_14958,N_14873);
nor UO_539 (O_539,N_14973,N_14922);
nor UO_540 (O_540,N_14955,N_14968);
nand UO_541 (O_541,N_14873,N_14890);
and UO_542 (O_542,N_14876,N_14874);
and UO_543 (O_543,N_14883,N_14851);
nor UO_544 (O_544,N_14974,N_14969);
nor UO_545 (O_545,N_14957,N_14975);
nor UO_546 (O_546,N_14874,N_14889);
and UO_547 (O_547,N_14993,N_14911);
nand UO_548 (O_548,N_14902,N_14854);
nand UO_549 (O_549,N_14876,N_14980);
nor UO_550 (O_550,N_14979,N_14999);
and UO_551 (O_551,N_14977,N_14952);
nand UO_552 (O_552,N_14978,N_14961);
nor UO_553 (O_553,N_14961,N_14967);
xnor UO_554 (O_554,N_14935,N_14966);
nor UO_555 (O_555,N_14970,N_14910);
xor UO_556 (O_556,N_14993,N_14990);
and UO_557 (O_557,N_14943,N_14993);
xor UO_558 (O_558,N_14938,N_14896);
and UO_559 (O_559,N_14861,N_14967);
and UO_560 (O_560,N_14962,N_14869);
and UO_561 (O_561,N_14871,N_14928);
nor UO_562 (O_562,N_14965,N_14969);
xor UO_563 (O_563,N_14927,N_14902);
xnor UO_564 (O_564,N_14958,N_14880);
and UO_565 (O_565,N_14887,N_14949);
xor UO_566 (O_566,N_14948,N_14858);
nor UO_567 (O_567,N_14950,N_14951);
or UO_568 (O_568,N_14969,N_14911);
nor UO_569 (O_569,N_14983,N_14943);
xnor UO_570 (O_570,N_14993,N_14969);
and UO_571 (O_571,N_14958,N_14932);
nor UO_572 (O_572,N_14948,N_14957);
xnor UO_573 (O_573,N_14878,N_14898);
nor UO_574 (O_574,N_14850,N_14854);
xor UO_575 (O_575,N_14874,N_14949);
nor UO_576 (O_576,N_14899,N_14977);
or UO_577 (O_577,N_14963,N_14962);
nand UO_578 (O_578,N_14950,N_14876);
and UO_579 (O_579,N_14991,N_14878);
xnor UO_580 (O_580,N_14977,N_14980);
xor UO_581 (O_581,N_14928,N_14941);
nor UO_582 (O_582,N_14859,N_14882);
or UO_583 (O_583,N_14901,N_14942);
nand UO_584 (O_584,N_14869,N_14863);
and UO_585 (O_585,N_14969,N_14870);
nor UO_586 (O_586,N_14885,N_14935);
nor UO_587 (O_587,N_14922,N_14906);
xor UO_588 (O_588,N_14895,N_14918);
and UO_589 (O_589,N_14934,N_14966);
nand UO_590 (O_590,N_14863,N_14927);
nand UO_591 (O_591,N_14938,N_14992);
or UO_592 (O_592,N_14979,N_14868);
nor UO_593 (O_593,N_14880,N_14953);
nor UO_594 (O_594,N_14983,N_14930);
xnor UO_595 (O_595,N_14918,N_14917);
xnor UO_596 (O_596,N_14945,N_14884);
xor UO_597 (O_597,N_14909,N_14985);
xnor UO_598 (O_598,N_14960,N_14995);
and UO_599 (O_599,N_14934,N_14920);
or UO_600 (O_600,N_14905,N_14874);
xnor UO_601 (O_601,N_14943,N_14937);
nand UO_602 (O_602,N_14873,N_14904);
xnor UO_603 (O_603,N_14884,N_14880);
nor UO_604 (O_604,N_14894,N_14856);
xnor UO_605 (O_605,N_14955,N_14934);
and UO_606 (O_606,N_14898,N_14909);
and UO_607 (O_607,N_14896,N_14952);
nor UO_608 (O_608,N_14923,N_14857);
nand UO_609 (O_609,N_14978,N_14854);
or UO_610 (O_610,N_14998,N_14957);
or UO_611 (O_611,N_14998,N_14983);
nand UO_612 (O_612,N_14927,N_14935);
nand UO_613 (O_613,N_14882,N_14978);
xor UO_614 (O_614,N_14918,N_14899);
or UO_615 (O_615,N_14951,N_14991);
nor UO_616 (O_616,N_14851,N_14977);
nand UO_617 (O_617,N_14978,N_14936);
or UO_618 (O_618,N_14867,N_14937);
nor UO_619 (O_619,N_14924,N_14925);
or UO_620 (O_620,N_14987,N_14862);
nand UO_621 (O_621,N_14896,N_14895);
nor UO_622 (O_622,N_14968,N_14967);
xnor UO_623 (O_623,N_14993,N_14910);
and UO_624 (O_624,N_14852,N_14983);
and UO_625 (O_625,N_14926,N_14929);
and UO_626 (O_626,N_14978,N_14860);
and UO_627 (O_627,N_14997,N_14876);
xor UO_628 (O_628,N_14968,N_14903);
and UO_629 (O_629,N_14944,N_14906);
nor UO_630 (O_630,N_14946,N_14934);
and UO_631 (O_631,N_14852,N_14898);
and UO_632 (O_632,N_14976,N_14887);
and UO_633 (O_633,N_14929,N_14911);
or UO_634 (O_634,N_14934,N_14990);
and UO_635 (O_635,N_14964,N_14970);
and UO_636 (O_636,N_14871,N_14980);
or UO_637 (O_637,N_14910,N_14998);
xor UO_638 (O_638,N_14983,N_14971);
xor UO_639 (O_639,N_14922,N_14937);
nand UO_640 (O_640,N_14971,N_14955);
or UO_641 (O_641,N_14908,N_14956);
or UO_642 (O_642,N_14958,N_14867);
or UO_643 (O_643,N_14860,N_14924);
nand UO_644 (O_644,N_14934,N_14915);
nand UO_645 (O_645,N_14986,N_14898);
nor UO_646 (O_646,N_14910,N_14997);
nor UO_647 (O_647,N_14885,N_14864);
nand UO_648 (O_648,N_14988,N_14996);
nand UO_649 (O_649,N_14970,N_14912);
nand UO_650 (O_650,N_14854,N_14857);
or UO_651 (O_651,N_14998,N_14851);
and UO_652 (O_652,N_14928,N_14959);
or UO_653 (O_653,N_14911,N_14957);
or UO_654 (O_654,N_14884,N_14948);
xnor UO_655 (O_655,N_14958,N_14940);
nor UO_656 (O_656,N_14965,N_14938);
and UO_657 (O_657,N_14933,N_14911);
and UO_658 (O_658,N_14911,N_14858);
and UO_659 (O_659,N_14895,N_14902);
nand UO_660 (O_660,N_14922,N_14928);
and UO_661 (O_661,N_14903,N_14961);
and UO_662 (O_662,N_14977,N_14964);
and UO_663 (O_663,N_14858,N_14909);
and UO_664 (O_664,N_14879,N_14946);
nor UO_665 (O_665,N_14976,N_14912);
or UO_666 (O_666,N_14930,N_14958);
and UO_667 (O_667,N_14890,N_14968);
nor UO_668 (O_668,N_14902,N_14937);
nor UO_669 (O_669,N_14962,N_14927);
xnor UO_670 (O_670,N_14858,N_14967);
nand UO_671 (O_671,N_14957,N_14869);
or UO_672 (O_672,N_14861,N_14983);
nand UO_673 (O_673,N_14925,N_14890);
or UO_674 (O_674,N_14985,N_14956);
nor UO_675 (O_675,N_14926,N_14915);
nand UO_676 (O_676,N_14957,N_14868);
and UO_677 (O_677,N_14941,N_14864);
or UO_678 (O_678,N_14982,N_14915);
nor UO_679 (O_679,N_14912,N_14986);
nor UO_680 (O_680,N_14980,N_14947);
and UO_681 (O_681,N_14921,N_14987);
and UO_682 (O_682,N_14922,N_14864);
nor UO_683 (O_683,N_14923,N_14883);
nor UO_684 (O_684,N_14868,N_14903);
nor UO_685 (O_685,N_14870,N_14851);
xor UO_686 (O_686,N_14995,N_14891);
nand UO_687 (O_687,N_14928,N_14909);
or UO_688 (O_688,N_14925,N_14907);
xor UO_689 (O_689,N_14962,N_14959);
or UO_690 (O_690,N_14903,N_14897);
xnor UO_691 (O_691,N_14864,N_14943);
nor UO_692 (O_692,N_14925,N_14893);
xnor UO_693 (O_693,N_14859,N_14960);
and UO_694 (O_694,N_14869,N_14925);
xor UO_695 (O_695,N_14889,N_14890);
nor UO_696 (O_696,N_14856,N_14928);
nand UO_697 (O_697,N_14909,N_14925);
nand UO_698 (O_698,N_14883,N_14954);
nand UO_699 (O_699,N_14898,N_14889);
or UO_700 (O_700,N_14897,N_14980);
nand UO_701 (O_701,N_14933,N_14963);
nor UO_702 (O_702,N_14855,N_14892);
or UO_703 (O_703,N_14955,N_14993);
or UO_704 (O_704,N_14992,N_14903);
and UO_705 (O_705,N_14876,N_14913);
or UO_706 (O_706,N_14914,N_14894);
or UO_707 (O_707,N_14932,N_14923);
or UO_708 (O_708,N_14865,N_14900);
nor UO_709 (O_709,N_14920,N_14891);
nand UO_710 (O_710,N_14939,N_14906);
and UO_711 (O_711,N_14873,N_14985);
nor UO_712 (O_712,N_14978,N_14946);
xor UO_713 (O_713,N_14926,N_14880);
nor UO_714 (O_714,N_14976,N_14991);
nand UO_715 (O_715,N_14866,N_14956);
nand UO_716 (O_716,N_14961,N_14875);
xnor UO_717 (O_717,N_14973,N_14924);
and UO_718 (O_718,N_14942,N_14920);
xor UO_719 (O_719,N_14975,N_14909);
or UO_720 (O_720,N_14857,N_14938);
or UO_721 (O_721,N_14871,N_14930);
or UO_722 (O_722,N_14996,N_14895);
nand UO_723 (O_723,N_14916,N_14880);
and UO_724 (O_724,N_14918,N_14992);
or UO_725 (O_725,N_14967,N_14866);
and UO_726 (O_726,N_14879,N_14986);
xnor UO_727 (O_727,N_14940,N_14948);
nand UO_728 (O_728,N_14894,N_14959);
xor UO_729 (O_729,N_14890,N_14991);
or UO_730 (O_730,N_14902,N_14982);
xor UO_731 (O_731,N_14991,N_14999);
or UO_732 (O_732,N_14925,N_14998);
and UO_733 (O_733,N_14911,N_14942);
xor UO_734 (O_734,N_14882,N_14898);
nand UO_735 (O_735,N_14963,N_14885);
nor UO_736 (O_736,N_14971,N_14895);
xnor UO_737 (O_737,N_14904,N_14953);
xnor UO_738 (O_738,N_14862,N_14900);
and UO_739 (O_739,N_14872,N_14901);
or UO_740 (O_740,N_14910,N_14943);
and UO_741 (O_741,N_14872,N_14860);
nand UO_742 (O_742,N_14978,N_14928);
nor UO_743 (O_743,N_14852,N_14989);
nor UO_744 (O_744,N_14940,N_14989);
and UO_745 (O_745,N_14965,N_14878);
nand UO_746 (O_746,N_14881,N_14924);
or UO_747 (O_747,N_14862,N_14981);
or UO_748 (O_748,N_14906,N_14855);
nor UO_749 (O_749,N_14872,N_14965);
nor UO_750 (O_750,N_14982,N_14855);
xor UO_751 (O_751,N_14921,N_14947);
nor UO_752 (O_752,N_14925,N_14857);
nand UO_753 (O_753,N_14982,N_14962);
and UO_754 (O_754,N_14952,N_14869);
xor UO_755 (O_755,N_14853,N_14933);
xor UO_756 (O_756,N_14865,N_14917);
nand UO_757 (O_757,N_14963,N_14915);
and UO_758 (O_758,N_14987,N_14891);
and UO_759 (O_759,N_14857,N_14886);
or UO_760 (O_760,N_14943,N_14927);
and UO_761 (O_761,N_14851,N_14854);
nor UO_762 (O_762,N_14882,N_14954);
nor UO_763 (O_763,N_14964,N_14942);
nor UO_764 (O_764,N_14874,N_14922);
or UO_765 (O_765,N_14973,N_14958);
xor UO_766 (O_766,N_14953,N_14955);
nand UO_767 (O_767,N_14856,N_14931);
and UO_768 (O_768,N_14944,N_14930);
nor UO_769 (O_769,N_14858,N_14958);
nand UO_770 (O_770,N_14986,N_14919);
nand UO_771 (O_771,N_14878,N_14969);
nand UO_772 (O_772,N_14999,N_14922);
and UO_773 (O_773,N_14850,N_14945);
and UO_774 (O_774,N_14949,N_14947);
and UO_775 (O_775,N_14989,N_14924);
and UO_776 (O_776,N_14951,N_14945);
and UO_777 (O_777,N_14999,N_14852);
xnor UO_778 (O_778,N_14882,N_14963);
or UO_779 (O_779,N_14977,N_14905);
or UO_780 (O_780,N_14943,N_14953);
or UO_781 (O_781,N_14857,N_14961);
nor UO_782 (O_782,N_14983,N_14914);
xor UO_783 (O_783,N_14859,N_14966);
and UO_784 (O_784,N_14869,N_14993);
or UO_785 (O_785,N_14923,N_14891);
nand UO_786 (O_786,N_14952,N_14937);
nor UO_787 (O_787,N_14866,N_14938);
nand UO_788 (O_788,N_14945,N_14987);
nand UO_789 (O_789,N_14892,N_14984);
and UO_790 (O_790,N_14994,N_14895);
nand UO_791 (O_791,N_14933,N_14923);
or UO_792 (O_792,N_14927,N_14959);
nand UO_793 (O_793,N_14867,N_14948);
nor UO_794 (O_794,N_14965,N_14920);
nand UO_795 (O_795,N_14950,N_14991);
nand UO_796 (O_796,N_14981,N_14929);
or UO_797 (O_797,N_14981,N_14850);
nand UO_798 (O_798,N_14969,N_14858);
or UO_799 (O_799,N_14977,N_14979);
nor UO_800 (O_800,N_14999,N_14968);
or UO_801 (O_801,N_14933,N_14934);
or UO_802 (O_802,N_14943,N_14930);
and UO_803 (O_803,N_14994,N_14892);
and UO_804 (O_804,N_14858,N_14889);
xor UO_805 (O_805,N_14961,N_14948);
nor UO_806 (O_806,N_14902,N_14975);
xor UO_807 (O_807,N_14937,N_14855);
xor UO_808 (O_808,N_14939,N_14990);
nand UO_809 (O_809,N_14910,N_14895);
xnor UO_810 (O_810,N_14869,N_14960);
nor UO_811 (O_811,N_14996,N_14914);
and UO_812 (O_812,N_14950,N_14934);
and UO_813 (O_813,N_14932,N_14994);
nor UO_814 (O_814,N_14993,N_14858);
nand UO_815 (O_815,N_14977,N_14932);
xor UO_816 (O_816,N_14951,N_14964);
nor UO_817 (O_817,N_14857,N_14939);
or UO_818 (O_818,N_14981,N_14919);
or UO_819 (O_819,N_14974,N_14888);
and UO_820 (O_820,N_14945,N_14975);
and UO_821 (O_821,N_14932,N_14876);
or UO_822 (O_822,N_14978,N_14907);
xor UO_823 (O_823,N_14964,N_14999);
and UO_824 (O_824,N_14925,N_14990);
and UO_825 (O_825,N_14912,N_14909);
or UO_826 (O_826,N_14904,N_14859);
and UO_827 (O_827,N_14962,N_14854);
nand UO_828 (O_828,N_14941,N_14897);
nor UO_829 (O_829,N_14875,N_14871);
xnor UO_830 (O_830,N_14965,N_14931);
nor UO_831 (O_831,N_14991,N_14980);
or UO_832 (O_832,N_14927,N_14860);
xnor UO_833 (O_833,N_14947,N_14873);
nor UO_834 (O_834,N_14946,N_14886);
xor UO_835 (O_835,N_14982,N_14940);
and UO_836 (O_836,N_14983,N_14988);
nand UO_837 (O_837,N_14971,N_14923);
nor UO_838 (O_838,N_14994,N_14878);
xor UO_839 (O_839,N_14933,N_14962);
xnor UO_840 (O_840,N_14885,N_14877);
nand UO_841 (O_841,N_14918,N_14931);
xnor UO_842 (O_842,N_14962,N_14922);
or UO_843 (O_843,N_14901,N_14912);
xor UO_844 (O_844,N_14987,N_14947);
xnor UO_845 (O_845,N_14900,N_14958);
xnor UO_846 (O_846,N_14969,N_14853);
or UO_847 (O_847,N_14853,N_14932);
nand UO_848 (O_848,N_14927,N_14871);
or UO_849 (O_849,N_14854,N_14895);
or UO_850 (O_850,N_14876,N_14862);
or UO_851 (O_851,N_14854,N_14938);
nand UO_852 (O_852,N_14920,N_14949);
and UO_853 (O_853,N_14853,N_14850);
xnor UO_854 (O_854,N_14977,N_14896);
nor UO_855 (O_855,N_14931,N_14981);
xnor UO_856 (O_856,N_14981,N_14978);
nand UO_857 (O_857,N_14887,N_14851);
nand UO_858 (O_858,N_14981,N_14952);
nor UO_859 (O_859,N_14957,N_14932);
or UO_860 (O_860,N_14963,N_14901);
xor UO_861 (O_861,N_14882,N_14969);
nor UO_862 (O_862,N_14933,N_14884);
and UO_863 (O_863,N_14951,N_14865);
and UO_864 (O_864,N_14900,N_14955);
nor UO_865 (O_865,N_14940,N_14986);
xor UO_866 (O_866,N_14943,N_14990);
and UO_867 (O_867,N_14941,N_14898);
nor UO_868 (O_868,N_14981,N_14993);
and UO_869 (O_869,N_14879,N_14898);
nor UO_870 (O_870,N_14959,N_14889);
xnor UO_871 (O_871,N_14917,N_14903);
xor UO_872 (O_872,N_14916,N_14924);
or UO_873 (O_873,N_14943,N_14914);
nand UO_874 (O_874,N_14986,N_14884);
or UO_875 (O_875,N_14939,N_14856);
and UO_876 (O_876,N_14948,N_14979);
nor UO_877 (O_877,N_14929,N_14934);
and UO_878 (O_878,N_14931,N_14857);
xnor UO_879 (O_879,N_14985,N_14975);
xor UO_880 (O_880,N_14886,N_14985);
nand UO_881 (O_881,N_14994,N_14946);
nand UO_882 (O_882,N_14865,N_14895);
nor UO_883 (O_883,N_14924,N_14955);
nand UO_884 (O_884,N_14977,N_14993);
nand UO_885 (O_885,N_14866,N_14987);
nand UO_886 (O_886,N_14987,N_14900);
nor UO_887 (O_887,N_14948,N_14910);
nor UO_888 (O_888,N_14931,N_14897);
or UO_889 (O_889,N_14975,N_14952);
nor UO_890 (O_890,N_14917,N_14861);
and UO_891 (O_891,N_14875,N_14877);
and UO_892 (O_892,N_14997,N_14892);
or UO_893 (O_893,N_14931,N_14970);
nand UO_894 (O_894,N_14909,N_14938);
nand UO_895 (O_895,N_14873,N_14889);
nand UO_896 (O_896,N_14990,N_14860);
nand UO_897 (O_897,N_14892,N_14854);
and UO_898 (O_898,N_14955,N_14863);
nor UO_899 (O_899,N_14984,N_14919);
xnor UO_900 (O_900,N_14999,N_14990);
and UO_901 (O_901,N_14873,N_14885);
and UO_902 (O_902,N_14998,N_14907);
nand UO_903 (O_903,N_14883,N_14959);
xor UO_904 (O_904,N_14981,N_14923);
and UO_905 (O_905,N_14887,N_14861);
nand UO_906 (O_906,N_14950,N_14861);
nor UO_907 (O_907,N_14918,N_14976);
xor UO_908 (O_908,N_14891,N_14906);
nand UO_909 (O_909,N_14922,N_14963);
or UO_910 (O_910,N_14895,N_14928);
xor UO_911 (O_911,N_14938,N_14928);
xor UO_912 (O_912,N_14977,N_14929);
nand UO_913 (O_913,N_14899,N_14943);
and UO_914 (O_914,N_14958,N_14992);
xor UO_915 (O_915,N_14963,N_14998);
nor UO_916 (O_916,N_14948,N_14857);
xnor UO_917 (O_917,N_14978,N_14896);
or UO_918 (O_918,N_14994,N_14854);
xor UO_919 (O_919,N_14997,N_14901);
or UO_920 (O_920,N_14861,N_14958);
and UO_921 (O_921,N_14884,N_14917);
xnor UO_922 (O_922,N_14978,N_14983);
nand UO_923 (O_923,N_14910,N_14931);
xnor UO_924 (O_924,N_14850,N_14923);
xor UO_925 (O_925,N_14990,N_14904);
nor UO_926 (O_926,N_14899,N_14942);
nor UO_927 (O_927,N_14999,N_14860);
and UO_928 (O_928,N_14853,N_14883);
or UO_929 (O_929,N_14867,N_14919);
nor UO_930 (O_930,N_14859,N_14866);
or UO_931 (O_931,N_14855,N_14896);
nand UO_932 (O_932,N_14923,N_14982);
or UO_933 (O_933,N_14917,N_14876);
and UO_934 (O_934,N_14932,N_14894);
xnor UO_935 (O_935,N_14870,N_14998);
xor UO_936 (O_936,N_14936,N_14987);
nor UO_937 (O_937,N_14866,N_14879);
and UO_938 (O_938,N_14857,N_14896);
nor UO_939 (O_939,N_14985,N_14944);
nor UO_940 (O_940,N_14948,N_14951);
nor UO_941 (O_941,N_14972,N_14930);
nand UO_942 (O_942,N_14950,N_14972);
nor UO_943 (O_943,N_14884,N_14874);
xor UO_944 (O_944,N_14850,N_14903);
or UO_945 (O_945,N_14857,N_14975);
nand UO_946 (O_946,N_14886,N_14893);
or UO_947 (O_947,N_14936,N_14902);
nand UO_948 (O_948,N_14962,N_14957);
nand UO_949 (O_949,N_14960,N_14955);
xnor UO_950 (O_950,N_14903,N_14918);
and UO_951 (O_951,N_14963,N_14886);
and UO_952 (O_952,N_14958,N_14961);
xnor UO_953 (O_953,N_14955,N_14986);
xor UO_954 (O_954,N_14863,N_14953);
xor UO_955 (O_955,N_14950,N_14872);
nand UO_956 (O_956,N_14945,N_14944);
xnor UO_957 (O_957,N_14905,N_14912);
or UO_958 (O_958,N_14969,N_14988);
nand UO_959 (O_959,N_14936,N_14958);
and UO_960 (O_960,N_14993,N_14932);
nor UO_961 (O_961,N_14956,N_14938);
or UO_962 (O_962,N_14955,N_14926);
nand UO_963 (O_963,N_14869,N_14988);
and UO_964 (O_964,N_14860,N_14875);
and UO_965 (O_965,N_14888,N_14944);
nor UO_966 (O_966,N_14965,N_14913);
xnor UO_967 (O_967,N_14876,N_14872);
nand UO_968 (O_968,N_14991,N_14971);
nand UO_969 (O_969,N_14955,N_14894);
nor UO_970 (O_970,N_14958,N_14983);
xnor UO_971 (O_971,N_14854,N_14991);
xnor UO_972 (O_972,N_14932,N_14961);
xor UO_973 (O_973,N_14919,N_14885);
xnor UO_974 (O_974,N_14964,N_14907);
and UO_975 (O_975,N_14922,N_14907);
nor UO_976 (O_976,N_14989,N_14953);
nand UO_977 (O_977,N_14886,N_14973);
or UO_978 (O_978,N_14913,N_14901);
or UO_979 (O_979,N_14956,N_14914);
xnor UO_980 (O_980,N_14876,N_14952);
xnor UO_981 (O_981,N_14987,N_14935);
and UO_982 (O_982,N_14955,N_14914);
xnor UO_983 (O_983,N_14876,N_14912);
nand UO_984 (O_984,N_14963,N_14949);
and UO_985 (O_985,N_14881,N_14942);
and UO_986 (O_986,N_14937,N_14935);
nor UO_987 (O_987,N_14978,N_14970);
and UO_988 (O_988,N_14944,N_14884);
nand UO_989 (O_989,N_14959,N_14922);
and UO_990 (O_990,N_14860,N_14995);
and UO_991 (O_991,N_14976,N_14980);
nand UO_992 (O_992,N_14934,N_14952);
and UO_993 (O_993,N_14908,N_14887);
nand UO_994 (O_994,N_14903,N_14865);
nor UO_995 (O_995,N_14900,N_14962);
nand UO_996 (O_996,N_14975,N_14976);
and UO_997 (O_997,N_14894,N_14882);
nor UO_998 (O_998,N_14924,N_14936);
or UO_999 (O_999,N_14929,N_14992);
nand UO_1000 (O_1000,N_14972,N_14870);
and UO_1001 (O_1001,N_14935,N_14951);
nor UO_1002 (O_1002,N_14959,N_14896);
nand UO_1003 (O_1003,N_14868,N_14871);
and UO_1004 (O_1004,N_14959,N_14875);
or UO_1005 (O_1005,N_14851,N_14940);
nand UO_1006 (O_1006,N_14884,N_14864);
nand UO_1007 (O_1007,N_14955,N_14940);
and UO_1008 (O_1008,N_14946,N_14920);
and UO_1009 (O_1009,N_14969,N_14940);
xnor UO_1010 (O_1010,N_14868,N_14866);
nand UO_1011 (O_1011,N_14877,N_14895);
nor UO_1012 (O_1012,N_14867,N_14916);
nor UO_1013 (O_1013,N_14960,N_14938);
or UO_1014 (O_1014,N_14953,N_14850);
nor UO_1015 (O_1015,N_14910,N_14989);
nor UO_1016 (O_1016,N_14907,N_14877);
or UO_1017 (O_1017,N_14992,N_14913);
xor UO_1018 (O_1018,N_14950,N_14862);
nand UO_1019 (O_1019,N_14865,N_14902);
nand UO_1020 (O_1020,N_14913,N_14897);
nand UO_1021 (O_1021,N_14871,N_14913);
and UO_1022 (O_1022,N_14997,N_14987);
nor UO_1023 (O_1023,N_14979,N_14881);
and UO_1024 (O_1024,N_14974,N_14853);
nand UO_1025 (O_1025,N_14962,N_14863);
nand UO_1026 (O_1026,N_14896,N_14926);
nand UO_1027 (O_1027,N_14931,N_14854);
or UO_1028 (O_1028,N_14953,N_14886);
nor UO_1029 (O_1029,N_14924,N_14877);
or UO_1030 (O_1030,N_14916,N_14856);
and UO_1031 (O_1031,N_14986,N_14984);
and UO_1032 (O_1032,N_14928,N_14913);
nor UO_1033 (O_1033,N_14994,N_14949);
nand UO_1034 (O_1034,N_14876,N_14854);
or UO_1035 (O_1035,N_14888,N_14947);
nor UO_1036 (O_1036,N_14944,N_14940);
xnor UO_1037 (O_1037,N_14911,N_14947);
xnor UO_1038 (O_1038,N_14872,N_14939);
nor UO_1039 (O_1039,N_14972,N_14883);
nor UO_1040 (O_1040,N_14956,N_14925);
or UO_1041 (O_1041,N_14853,N_14914);
nor UO_1042 (O_1042,N_14892,N_14907);
or UO_1043 (O_1043,N_14870,N_14924);
and UO_1044 (O_1044,N_14852,N_14971);
nor UO_1045 (O_1045,N_14924,N_14898);
nor UO_1046 (O_1046,N_14979,N_14855);
and UO_1047 (O_1047,N_14959,N_14911);
and UO_1048 (O_1048,N_14904,N_14897);
nor UO_1049 (O_1049,N_14911,N_14941);
xor UO_1050 (O_1050,N_14948,N_14935);
and UO_1051 (O_1051,N_14864,N_14978);
or UO_1052 (O_1052,N_14909,N_14892);
and UO_1053 (O_1053,N_14869,N_14938);
nor UO_1054 (O_1054,N_14945,N_14859);
xnor UO_1055 (O_1055,N_14934,N_14956);
xor UO_1056 (O_1056,N_14942,N_14862);
and UO_1057 (O_1057,N_14893,N_14887);
or UO_1058 (O_1058,N_14915,N_14898);
and UO_1059 (O_1059,N_14880,N_14954);
and UO_1060 (O_1060,N_14996,N_14867);
xnor UO_1061 (O_1061,N_14958,N_14944);
nand UO_1062 (O_1062,N_14862,N_14867);
or UO_1063 (O_1063,N_14924,N_14918);
and UO_1064 (O_1064,N_14887,N_14989);
or UO_1065 (O_1065,N_14989,N_14985);
or UO_1066 (O_1066,N_14867,N_14978);
nand UO_1067 (O_1067,N_14871,N_14953);
or UO_1068 (O_1068,N_14974,N_14851);
nand UO_1069 (O_1069,N_14921,N_14992);
and UO_1070 (O_1070,N_14949,N_14865);
nand UO_1071 (O_1071,N_14901,N_14914);
nor UO_1072 (O_1072,N_14965,N_14948);
nor UO_1073 (O_1073,N_14876,N_14995);
nor UO_1074 (O_1074,N_14935,N_14975);
and UO_1075 (O_1075,N_14966,N_14919);
nor UO_1076 (O_1076,N_14871,N_14886);
nor UO_1077 (O_1077,N_14912,N_14891);
or UO_1078 (O_1078,N_14957,N_14952);
or UO_1079 (O_1079,N_14892,N_14919);
nor UO_1080 (O_1080,N_14903,N_14975);
or UO_1081 (O_1081,N_14919,N_14909);
nor UO_1082 (O_1082,N_14961,N_14943);
nand UO_1083 (O_1083,N_14935,N_14979);
and UO_1084 (O_1084,N_14923,N_14917);
or UO_1085 (O_1085,N_14855,N_14974);
or UO_1086 (O_1086,N_14925,N_14879);
nand UO_1087 (O_1087,N_14998,N_14937);
nor UO_1088 (O_1088,N_14908,N_14994);
and UO_1089 (O_1089,N_14899,N_14917);
nor UO_1090 (O_1090,N_14915,N_14920);
xnor UO_1091 (O_1091,N_14938,N_14958);
nor UO_1092 (O_1092,N_14921,N_14970);
nor UO_1093 (O_1093,N_14875,N_14885);
or UO_1094 (O_1094,N_14884,N_14887);
nand UO_1095 (O_1095,N_14972,N_14994);
and UO_1096 (O_1096,N_14963,N_14862);
or UO_1097 (O_1097,N_14973,N_14993);
nor UO_1098 (O_1098,N_14955,N_14927);
and UO_1099 (O_1099,N_14923,N_14920);
and UO_1100 (O_1100,N_14908,N_14991);
or UO_1101 (O_1101,N_14940,N_14925);
and UO_1102 (O_1102,N_14930,N_14995);
nor UO_1103 (O_1103,N_14871,N_14861);
nor UO_1104 (O_1104,N_14896,N_14968);
nand UO_1105 (O_1105,N_14959,N_14979);
nand UO_1106 (O_1106,N_14891,N_14935);
nand UO_1107 (O_1107,N_14934,N_14862);
nor UO_1108 (O_1108,N_14979,N_14928);
nand UO_1109 (O_1109,N_14976,N_14865);
nand UO_1110 (O_1110,N_14949,N_14902);
xnor UO_1111 (O_1111,N_14985,N_14933);
and UO_1112 (O_1112,N_14883,N_14928);
or UO_1113 (O_1113,N_14906,N_14988);
or UO_1114 (O_1114,N_14917,N_14895);
nor UO_1115 (O_1115,N_14925,N_14991);
nand UO_1116 (O_1116,N_14883,N_14870);
nor UO_1117 (O_1117,N_14913,N_14908);
and UO_1118 (O_1118,N_14898,N_14961);
xor UO_1119 (O_1119,N_14863,N_14888);
or UO_1120 (O_1120,N_14974,N_14961);
and UO_1121 (O_1121,N_14965,N_14955);
and UO_1122 (O_1122,N_14933,N_14900);
xnor UO_1123 (O_1123,N_14915,N_14900);
nor UO_1124 (O_1124,N_14979,N_14900);
or UO_1125 (O_1125,N_14968,N_14980);
nand UO_1126 (O_1126,N_14943,N_14965);
and UO_1127 (O_1127,N_14877,N_14978);
nand UO_1128 (O_1128,N_14987,N_14990);
or UO_1129 (O_1129,N_14887,N_14968);
and UO_1130 (O_1130,N_14996,N_14945);
or UO_1131 (O_1131,N_14935,N_14915);
or UO_1132 (O_1132,N_14900,N_14853);
or UO_1133 (O_1133,N_14996,N_14908);
nand UO_1134 (O_1134,N_14856,N_14941);
xnor UO_1135 (O_1135,N_14861,N_14999);
and UO_1136 (O_1136,N_14866,N_14997);
and UO_1137 (O_1137,N_14950,N_14923);
nand UO_1138 (O_1138,N_14946,N_14853);
nor UO_1139 (O_1139,N_14971,N_14975);
and UO_1140 (O_1140,N_14854,N_14986);
xor UO_1141 (O_1141,N_14947,N_14978);
nor UO_1142 (O_1142,N_14956,N_14880);
xnor UO_1143 (O_1143,N_14873,N_14946);
and UO_1144 (O_1144,N_14914,N_14920);
nor UO_1145 (O_1145,N_14854,N_14946);
nor UO_1146 (O_1146,N_14928,N_14896);
or UO_1147 (O_1147,N_14992,N_14969);
and UO_1148 (O_1148,N_14966,N_14930);
nand UO_1149 (O_1149,N_14882,N_14895);
or UO_1150 (O_1150,N_14954,N_14889);
nand UO_1151 (O_1151,N_14877,N_14945);
xnor UO_1152 (O_1152,N_14915,N_14897);
nand UO_1153 (O_1153,N_14901,N_14996);
nand UO_1154 (O_1154,N_14974,N_14979);
nor UO_1155 (O_1155,N_14947,N_14869);
xnor UO_1156 (O_1156,N_14898,N_14948);
xnor UO_1157 (O_1157,N_14949,N_14850);
nor UO_1158 (O_1158,N_14929,N_14887);
xnor UO_1159 (O_1159,N_14878,N_14930);
xor UO_1160 (O_1160,N_14872,N_14941);
and UO_1161 (O_1161,N_14986,N_14983);
nor UO_1162 (O_1162,N_14938,N_14902);
xnor UO_1163 (O_1163,N_14891,N_14966);
and UO_1164 (O_1164,N_14990,N_14950);
nor UO_1165 (O_1165,N_14975,N_14996);
xnor UO_1166 (O_1166,N_14933,N_14986);
or UO_1167 (O_1167,N_14967,N_14914);
and UO_1168 (O_1168,N_14873,N_14859);
nor UO_1169 (O_1169,N_14952,N_14927);
xnor UO_1170 (O_1170,N_14874,N_14986);
nand UO_1171 (O_1171,N_14997,N_14858);
xnor UO_1172 (O_1172,N_14884,N_14899);
nand UO_1173 (O_1173,N_14866,N_14871);
nor UO_1174 (O_1174,N_14992,N_14931);
nand UO_1175 (O_1175,N_14977,N_14940);
nand UO_1176 (O_1176,N_14894,N_14883);
xnor UO_1177 (O_1177,N_14913,N_14980);
and UO_1178 (O_1178,N_14855,N_14889);
xor UO_1179 (O_1179,N_14852,N_14890);
nand UO_1180 (O_1180,N_14995,N_14958);
nor UO_1181 (O_1181,N_14862,N_14856);
nor UO_1182 (O_1182,N_14905,N_14994);
or UO_1183 (O_1183,N_14929,N_14994);
xor UO_1184 (O_1184,N_14964,N_14987);
xnor UO_1185 (O_1185,N_14980,N_14877);
nor UO_1186 (O_1186,N_14853,N_14865);
or UO_1187 (O_1187,N_14984,N_14875);
and UO_1188 (O_1188,N_14860,N_14874);
or UO_1189 (O_1189,N_14990,N_14894);
or UO_1190 (O_1190,N_14955,N_14954);
nor UO_1191 (O_1191,N_14914,N_14966);
nand UO_1192 (O_1192,N_14860,N_14894);
xnor UO_1193 (O_1193,N_14975,N_14862);
nand UO_1194 (O_1194,N_14996,N_14943);
and UO_1195 (O_1195,N_14896,N_14999);
nand UO_1196 (O_1196,N_14907,N_14893);
or UO_1197 (O_1197,N_14932,N_14852);
nand UO_1198 (O_1198,N_14863,N_14934);
and UO_1199 (O_1199,N_14930,N_14965);
nand UO_1200 (O_1200,N_14857,N_14947);
or UO_1201 (O_1201,N_14863,N_14924);
or UO_1202 (O_1202,N_14966,N_14858);
nor UO_1203 (O_1203,N_14975,N_14995);
nand UO_1204 (O_1204,N_14931,N_14996);
or UO_1205 (O_1205,N_14888,N_14990);
nand UO_1206 (O_1206,N_14951,N_14955);
and UO_1207 (O_1207,N_14855,N_14971);
nor UO_1208 (O_1208,N_14863,N_14973);
xor UO_1209 (O_1209,N_14867,N_14984);
or UO_1210 (O_1210,N_14965,N_14988);
or UO_1211 (O_1211,N_14946,N_14957);
nand UO_1212 (O_1212,N_14953,N_14901);
and UO_1213 (O_1213,N_14996,N_14852);
nor UO_1214 (O_1214,N_14870,N_14992);
xor UO_1215 (O_1215,N_14872,N_14884);
and UO_1216 (O_1216,N_14932,N_14867);
nor UO_1217 (O_1217,N_14914,N_14980);
or UO_1218 (O_1218,N_14937,N_14932);
and UO_1219 (O_1219,N_14850,N_14858);
xor UO_1220 (O_1220,N_14934,N_14936);
xnor UO_1221 (O_1221,N_14865,N_14922);
or UO_1222 (O_1222,N_14961,N_14872);
or UO_1223 (O_1223,N_14933,N_14904);
and UO_1224 (O_1224,N_14987,N_14961);
nor UO_1225 (O_1225,N_14894,N_14921);
and UO_1226 (O_1226,N_14965,N_14884);
and UO_1227 (O_1227,N_14956,N_14881);
xnor UO_1228 (O_1228,N_14916,N_14942);
nand UO_1229 (O_1229,N_14916,N_14897);
nand UO_1230 (O_1230,N_14893,N_14881);
nor UO_1231 (O_1231,N_14858,N_14886);
nor UO_1232 (O_1232,N_14951,N_14908);
xnor UO_1233 (O_1233,N_14962,N_14996);
xnor UO_1234 (O_1234,N_14897,N_14981);
nor UO_1235 (O_1235,N_14957,N_14892);
and UO_1236 (O_1236,N_14926,N_14945);
and UO_1237 (O_1237,N_14967,N_14951);
or UO_1238 (O_1238,N_14890,N_14938);
xnor UO_1239 (O_1239,N_14899,N_14896);
xor UO_1240 (O_1240,N_14905,N_14887);
nor UO_1241 (O_1241,N_14975,N_14876);
nor UO_1242 (O_1242,N_14992,N_14998);
and UO_1243 (O_1243,N_14870,N_14859);
nor UO_1244 (O_1244,N_14921,N_14985);
or UO_1245 (O_1245,N_14945,N_14910);
nand UO_1246 (O_1246,N_14889,N_14961);
and UO_1247 (O_1247,N_14984,N_14882);
nor UO_1248 (O_1248,N_14882,N_14872);
nand UO_1249 (O_1249,N_14946,N_14960);
nor UO_1250 (O_1250,N_14956,N_14947);
and UO_1251 (O_1251,N_14895,N_14945);
xnor UO_1252 (O_1252,N_14969,N_14863);
or UO_1253 (O_1253,N_14988,N_14917);
nand UO_1254 (O_1254,N_14921,N_14867);
xor UO_1255 (O_1255,N_14921,N_14997);
xor UO_1256 (O_1256,N_14859,N_14922);
nor UO_1257 (O_1257,N_14994,N_14871);
nor UO_1258 (O_1258,N_14965,N_14871);
and UO_1259 (O_1259,N_14932,N_14964);
xor UO_1260 (O_1260,N_14909,N_14997);
and UO_1261 (O_1261,N_14995,N_14969);
nand UO_1262 (O_1262,N_14996,N_14889);
nand UO_1263 (O_1263,N_14961,N_14887);
nor UO_1264 (O_1264,N_14954,N_14913);
nand UO_1265 (O_1265,N_14992,N_14922);
nor UO_1266 (O_1266,N_14866,N_14957);
nor UO_1267 (O_1267,N_14920,N_14916);
and UO_1268 (O_1268,N_14895,N_14879);
nor UO_1269 (O_1269,N_14873,N_14864);
nor UO_1270 (O_1270,N_14910,N_14904);
and UO_1271 (O_1271,N_14997,N_14884);
xor UO_1272 (O_1272,N_14956,N_14982);
and UO_1273 (O_1273,N_14894,N_14984);
nand UO_1274 (O_1274,N_14909,N_14865);
and UO_1275 (O_1275,N_14919,N_14870);
nor UO_1276 (O_1276,N_14868,N_14913);
xnor UO_1277 (O_1277,N_14981,N_14964);
nand UO_1278 (O_1278,N_14953,N_14921);
or UO_1279 (O_1279,N_14972,N_14875);
xor UO_1280 (O_1280,N_14883,N_14891);
xor UO_1281 (O_1281,N_14930,N_14935);
xnor UO_1282 (O_1282,N_14911,N_14913);
xnor UO_1283 (O_1283,N_14961,N_14868);
xor UO_1284 (O_1284,N_14925,N_14901);
and UO_1285 (O_1285,N_14982,N_14986);
or UO_1286 (O_1286,N_14919,N_14992);
nor UO_1287 (O_1287,N_14953,N_14919);
or UO_1288 (O_1288,N_14873,N_14879);
or UO_1289 (O_1289,N_14900,N_14944);
xor UO_1290 (O_1290,N_14976,N_14968);
nand UO_1291 (O_1291,N_14974,N_14857);
or UO_1292 (O_1292,N_14955,N_14918);
nand UO_1293 (O_1293,N_14992,N_14892);
or UO_1294 (O_1294,N_14856,N_14883);
nand UO_1295 (O_1295,N_14984,N_14993);
or UO_1296 (O_1296,N_14892,N_14942);
nand UO_1297 (O_1297,N_14891,N_14953);
xnor UO_1298 (O_1298,N_14959,N_14850);
or UO_1299 (O_1299,N_14897,N_14854);
or UO_1300 (O_1300,N_14986,N_14957);
and UO_1301 (O_1301,N_14922,N_14964);
nor UO_1302 (O_1302,N_14970,N_14890);
or UO_1303 (O_1303,N_14977,N_14872);
xnor UO_1304 (O_1304,N_14921,N_14860);
and UO_1305 (O_1305,N_14889,N_14920);
xnor UO_1306 (O_1306,N_14921,N_14954);
xor UO_1307 (O_1307,N_14910,N_14976);
and UO_1308 (O_1308,N_14928,N_14865);
and UO_1309 (O_1309,N_14970,N_14966);
and UO_1310 (O_1310,N_14992,N_14975);
nand UO_1311 (O_1311,N_14910,N_14911);
and UO_1312 (O_1312,N_14935,N_14955);
or UO_1313 (O_1313,N_14942,N_14861);
nand UO_1314 (O_1314,N_14906,N_14857);
nor UO_1315 (O_1315,N_14898,N_14979);
and UO_1316 (O_1316,N_14968,N_14995);
xnor UO_1317 (O_1317,N_14982,N_14948);
nor UO_1318 (O_1318,N_14885,N_14857);
nor UO_1319 (O_1319,N_14916,N_14955);
and UO_1320 (O_1320,N_14937,N_14851);
nand UO_1321 (O_1321,N_14933,N_14885);
xnor UO_1322 (O_1322,N_14921,N_14889);
nand UO_1323 (O_1323,N_14966,N_14931);
nor UO_1324 (O_1324,N_14994,N_14875);
nor UO_1325 (O_1325,N_14971,N_14882);
xor UO_1326 (O_1326,N_14920,N_14924);
nor UO_1327 (O_1327,N_14931,N_14950);
xnor UO_1328 (O_1328,N_14942,N_14915);
nor UO_1329 (O_1329,N_14996,N_14947);
xor UO_1330 (O_1330,N_14970,N_14939);
nor UO_1331 (O_1331,N_14864,N_14871);
and UO_1332 (O_1332,N_14930,N_14959);
nand UO_1333 (O_1333,N_14967,N_14957);
nand UO_1334 (O_1334,N_14881,N_14953);
xor UO_1335 (O_1335,N_14901,N_14950);
nor UO_1336 (O_1336,N_14857,N_14954);
xor UO_1337 (O_1337,N_14891,N_14910);
and UO_1338 (O_1338,N_14852,N_14934);
and UO_1339 (O_1339,N_14946,N_14888);
and UO_1340 (O_1340,N_14959,N_14861);
and UO_1341 (O_1341,N_14869,N_14903);
and UO_1342 (O_1342,N_14921,N_14879);
nor UO_1343 (O_1343,N_14865,N_14851);
xor UO_1344 (O_1344,N_14977,N_14870);
and UO_1345 (O_1345,N_14933,N_14896);
or UO_1346 (O_1346,N_14886,N_14852);
or UO_1347 (O_1347,N_14933,N_14984);
nand UO_1348 (O_1348,N_14978,N_14888);
or UO_1349 (O_1349,N_14963,N_14996);
nand UO_1350 (O_1350,N_14892,N_14884);
nand UO_1351 (O_1351,N_14934,N_14986);
xor UO_1352 (O_1352,N_14996,N_14872);
nor UO_1353 (O_1353,N_14915,N_14909);
nor UO_1354 (O_1354,N_14900,N_14990);
nand UO_1355 (O_1355,N_14937,N_14988);
nor UO_1356 (O_1356,N_14899,N_14877);
and UO_1357 (O_1357,N_14971,N_14953);
and UO_1358 (O_1358,N_14967,N_14992);
nand UO_1359 (O_1359,N_14871,N_14912);
nor UO_1360 (O_1360,N_14859,N_14865);
xor UO_1361 (O_1361,N_14893,N_14997);
nor UO_1362 (O_1362,N_14851,N_14900);
xnor UO_1363 (O_1363,N_14963,N_14930);
xor UO_1364 (O_1364,N_14861,N_14901);
nand UO_1365 (O_1365,N_14852,N_14880);
or UO_1366 (O_1366,N_14973,N_14965);
xnor UO_1367 (O_1367,N_14905,N_14851);
or UO_1368 (O_1368,N_14896,N_14997);
nand UO_1369 (O_1369,N_14868,N_14972);
nor UO_1370 (O_1370,N_14946,N_14938);
xor UO_1371 (O_1371,N_14990,N_14963);
or UO_1372 (O_1372,N_14932,N_14929);
or UO_1373 (O_1373,N_14980,N_14989);
nand UO_1374 (O_1374,N_14928,N_14996);
xnor UO_1375 (O_1375,N_14966,N_14892);
or UO_1376 (O_1376,N_14860,N_14936);
or UO_1377 (O_1377,N_14897,N_14986);
xor UO_1378 (O_1378,N_14920,N_14888);
nand UO_1379 (O_1379,N_14923,N_14861);
nand UO_1380 (O_1380,N_14945,N_14928);
or UO_1381 (O_1381,N_14861,N_14876);
or UO_1382 (O_1382,N_14893,N_14922);
nor UO_1383 (O_1383,N_14914,N_14992);
or UO_1384 (O_1384,N_14882,N_14919);
or UO_1385 (O_1385,N_14915,N_14974);
or UO_1386 (O_1386,N_14928,N_14864);
nand UO_1387 (O_1387,N_14911,N_14974);
nand UO_1388 (O_1388,N_14883,N_14898);
or UO_1389 (O_1389,N_14882,N_14877);
xor UO_1390 (O_1390,N_14930,N_14939);
and UO_1391 (O_1391,N_14974,N_14907);
and UO_1392 (O_1392,N_14977,N_14860);
xor UO_1393 (O_1393,N_14870,N_14965);
and UO_1394 (O_1394,N_14907,N_14929);
and UO_1395 (O_1395,N_14990,N_14945);
and UO_1396 (O_1396,N_14875,N_14976);
and UO_1397 (O_1397,N_14913,N_14973);
and UO_1398 (O_1398,N_14896,N_14925);
nor UO_1399 (O_1399,N_14850,N_14925);
nand UO_1400 (O_1400,N_14945,N_14979);
xor UO_1401 (O_1401,N_14866,N_14954);
nand UO_1402 (O_1402,N_14908,N_14981);
or UO_1403 (O_1403,N_14992,N_14855);
nor UO_1404 (O_1404,N_14933,N_14872);
nand UO_1405 (O_1405,N_14963,N_14964);
and UO_1406 (O_1406,N_14959,N_14945);
nand UO_1407 (O_1407,N_14863,N_14862);
and UO_1408 (O_1408,N_14870,N_14971);
nor UO_1409 (O_1409,N_14968,N_14942);
nor UO_1410 (O_1410,N_14925,N_14903);
and UO_1411 (O_1411,N_14926,N_14997);
xor UO_1412 (O_1412,N_14957,N_14942);
and UO_1413 (O_1413,N_14860,N_14903);
xnor UO_1414 (O_1414,N_14987,N_14890);
xnor UO_1415 (O_1415,N_14886,N_14918);
nand UO_1416 (O_1416,N_14917,N_14922);
or UO_1417 (O_1417,N_14891,N_14855);
nor UO_1418 (O_1418,N_14875,N_14884);
nand UO_1419 (O_1419,N_14974,N_14914);
or UO_1420 (O_1420,N_14893,N_14905);
nand UO_1421 (O_1421,N_14921,N_14942);
xor UO_1422 (O_1422,N_14990,N_14985);
nand UO_1423 (O_1423,N_14896,N_14904);
and UO_1424 (O_1424,N_14952,N_14938);
nor UO_1425 (O_1425,N_14916,N_14964);
and UO_1426 (O_1426,N_14868,N_14953);
and UO_1427 (O_1427,N_14938,N_14893);
or UO_1428 (O_1428,N_14855,N_14879);
and UO_1429 (O_1429,N_14856,N_14994);
nor UO_1430 (O_1430,N_14990,N_14949);
or UO_1431 (O_1431,N_14991,N_14983);
or UO_1432 (O_1432,N_14853,N_14955);
nor UO_1433 (O_1433,N_14974,N_14868);
and UO_1434 (O_1434,N_14963,N_14880);
nor UO_1435 (O_1435,N_14934,N_14897);
nor UO_1436 (O_1436,N_14983,N_14881);
xnor UO_1437 (O_1437,N_14981,N_14909);
nand UO_1438 (O_1438,N_14985,N_14888);
xor UO_1439 (O_1439,N_14979,N_14878);
and UO_1440 (O_1440,N_14990,N_14889);
xor UO_1441 (O_1441,N_14901,N_14926);
or UO_1442 (O_1442,N_14902,N_14969);
xnor UO_1443 (O_1443,N_14880,N_14910);
nand UO_1444 (O_1444,N_14927,N_14987);
and UO_1445 (O_1445,N_14937,N_14891);
and UO_1446 (O_1446,N_14865,N_14897);
nor UO_1447 (O_1447,N_14850,N_14867);
nand UO_1448 (O_1448,N_14850,N_14915);
xor UO_1449 (O_1449,N_14984,N_14893);
xor UO_1450 (O_1450,N_14972,N_14911);
and UO_1451 (O_1451,N_14855,N_14925);
nand UO_1452 (O_1452,N_14993,N_14881);
nand UO_1453 (O_1453,N_14870,N_14905);
nor UO_1454 (O_1454,N_14873,N_14983);
xor UO_1455 (O_1455,N_14956,N_14919);
or UO_1456 (O_1456,N_14903,N_14983);
or UO_1457 (O_1457,N_14853,N_14930);
nor UO_1458 (O_1458,N_14862,N_14936);
xor UO_1459 (O_1459,N_14859,N_14878);
xor UO_1460 (O_1460,N_14947,N_14875);
nor UO_1461 (O_1461,N_14938,N_14914);
and UO_1462 (O_1462,N_14899,N_14975);
nand UO_1463 (O_1463,N_14966,N_14873);
xor UO_1464 (O_1464,N_14957,N_14886);
nand UO_1465 (O_1465,N_14927,N_14983);
nor UO_1466 (O_1466,N_14944,N_14890);
nand UO_1467 (O_1467,N_14889,N_14978);
nor UO_1468 (O_1468,N_14874,N_14978);
nor UO_1469 (O_1469,N_14878,N_14906);
and UO_1470 (O_1470,N_14877,N_14960);
nor UO_1471 (O_1471,N_14988,N_14975);
nor UO_1472 (O_1472,N_14902,N_14852);
xnor UO_1473 (O_1473,N_14989,N_14984);
nor UO_1474 (O_1474,N_14853,N_14957);
or UO_1475 (O_1475,N_14920,N_14945);
xnor UO_1476 (O_1476,N_14940,N_14980);
nor UO_1477 (O_1477,N_14944,N_14943);
nand UO_1478 (O_1478,N_14862,N_14861);
nor UO_1479 (O_1479,N_14863,N_14877);
nor UO_1480 (O_1480,N_14913,N_14856);
or UO_1481 (O_1481,N_14898,N_14990);
or UO_1482 (O_1482,N_14856,N_14907);
and UO_1483 (O_1483,N_14968,N_14975);
xnor UO_1484 (O_1484,N_14902,N_14904);
or UO_1485 (O_1485,N_14909,N_14993);
or UO_1486 (O_1486,N_14924,N_14984);
xnor UO_1487 (O_1487,N_14948,N_14953);
xor UO_1488 (O_1488,N_14984,N_14967);
and UO_1489 (O_1489,N_14997,N_14944);
or UO_1490 (O_1490,N_14963,N_14993);
nand UO_1491 (O_1491,N_14969,N_14894);
or UO_1492 (O_1492,N_14973,N_14946);
and UO_1493 (O_1493,N_14973,N_14926);
nor UO_1494 (O_1494,N_14993,N_14912);
nand UO_1495 (O_1495,N_14909,N_14947);
nor UO_1496 (O_1496,N_14981,N_14868);
xnor UO_1497 (O_1497,N_14934,N_14878);
nor UO_1498 (O_1498,N_14868,N_14986);
nor UO_1499 (O_1499,N_14941,N_14884);
and UO_1500 (O_1500,N_14890,N_14967);
or UO_1501 (O_1501,N_14939,N_14904);
nor UO_1502 (O_1502,N_14933,N_14876);
xnor UO_1503 (O_1503,N_14902,N_14970);
and UO_1504 (O_1504,N_14871,N_14858);
and UO_1505 (O_1505,N_14867,N_14863);
nand UO_1506 (O_1506,N_14868,N_14933);
or UO_1507 (O_1507,N_14990,N_14913);
and UO_1508 (O_1508,N_14912,N_14860);
and UO_1509 (O_1509,N_14902,N_14965);
nand UO_1510 (O_1510,N_14941,N_14940);
nand UO_1511 (O_1511,N_14988,N_14961);
or UO_1512 (O_1512,N_14982,N_14851);
xnor UO_1513 (O_1513,N_14889,N_14899);
and UO_1514 (O_1514,N_14945,N_14972);
or UO_1515 (O_1515,N_14930,N_14977);
xor UO_1516 (O_1516,N_14928,N_14952);
or UO_1517 (O_1517,N_14995,N_14979);
nand UO_1518 (O_1518,N_14930,N_14929);
nor UO_1519 (O_1519,N_14894,N_14982);
xor UO_1520 (O_1520,N_14891,N_14964);
and UO_1521 (O_1521,N_14865,N_14878);
and UO_1522 (O_1522,N_14991,N_14880);
or UO_1523 (O_1523,N_14962,N_14897);
xnor UO_1524 (O_1524,N_14903,N_14891);
xnor UO_1525 (O_1525,N_14960,N_14862);
xor UO_1526 (O_1526,N_14958,N_14918);
nor UO_1527 (O_1527,N_14922,N_14953);
xnor UO_1528 (O_1528,N_14948,N_14909);
or UO_1529 (O_1529,N_14926,N_14866);
xor UO_1530 (O_1530,N_14881,N_14869);
nand UO_1531 (O_1531,N_14853,N_14972);
nor UO_1532 (O_1532,N_14919,N_14979);
or UO_1533 (O_1533,N_14920,N_14951);
nor UO_1534 (O_1534,N_14878,N_14913);
nand UO_1535 (O_1535,N_14969,N_14923);
nand UO_1536 (O_1536,N_14991,N_14920);
nand UO_1537 (O_1537,N_14984,N_14978);
nand UO_1538 (O_1538,N_14998,N_14953);
or UO_1539 (O_1539,N_14953,N_14931);
nor UO_1540 (O_1540,N_14995,N_14928);
and UO_1541 (O_1541,N_14971,N_14868);
or UO_1542 (O_1542,N_14926,N_14993);
nor UO_1543 (O_1543,N_14853,N_14984);
and UO_1544 (O_1544,N_14961,N_14999);
and UO_1545 (O_1545,N_14992,N_14896);
xnor UO_1546 (O_1546,N_14976,N_14982);
nand UO_1547 (O_1547,N_14950,N_14912);
nand UO_1548 (O_1548,N_14987,N_14974);
xnor UO_1549 (O_1549,N_14941,N_14906);
and UO_1550 (O_1550,N_14851,N_14951);
and UO_1551 (O_1551,N_14941,N_14855);
nor UO_1552 (O_1552,N_14949,N_14906);
nand UO_1553 (O_1553,N_14943,N_14851);
nor UO_1554 (O_1554,N_14866,N_14919);
or UO_1555 (O_1555,N_14859,N_14883);
nand UO_1556 (O_1556,N_14859,N_14973);
or UO_1557 (O_1557,N_14942,N_14882);
and UO_1558 (O_1558,N_14942,N_14909);
xor UO_1559 (O_1559,N_14896,N_14886);
or UO_1560 (O_1560,N_14949,N_14860);
nand UO_1561 (O_1561,N_14943,N_14866);
nor UO_1562 (O_1562,N_14926,N_14979);
xor UO_1563 (O_1563,N_14856,N_14955);
and UO_1564 (O_1564,N_14925,N_14953);
nand UO_1565 (O_1565,N_14890,N_14948);
xnor UO_1566 (O_1566,N_14989,N_14850);
or UO_1567 (O_1567,N_14872,N_14909);
nor UO_1568 (O_1568,N_14936,N_14965);
nor UO_1569 (O_1569,N_14935,N_14850);
and UO_1570 (O_1570,N_14986,N_14852);
or UO_1571 (O_1571,N_14939,N_14892);
nor UO_1572 (O_1572,N_14859,N_14863);
nor UO_1573 (O_1573,N_14894,N_14979);
nor UO_1574 (O_1574,N_14945,N_14934);
nand UO_1575 (O_1575,N_14946,N_14895);
nand UO_1576 (O_1576,N_14956,N_14943);
and UO_1577 (O_1577,N_14989,N_14905);
or UO_1578 (O_1578,N_14936,N_14942);
nor UO_1579 (O_1579,N_14943,N_14934);
or UO_1580 (O_1580,N_14871,N_14958);
xor UO_1581 (O_1581,N_14942,N_14993);
nand UO_1582 (O_1582,N_14899,N_14983);
xor UO_1583 (O_1583,N_14973,N_14936);
nand UO_1584 (O_1584,N_14964,N_14930);
xor UO_1585 (O_1585,N_14896,N_14939);
nor UO_1586 (O_1586,N_14858,N_14955);
or UO_1587 (O_1587,N_14850,N_14866);
nor UO_1588 (O_1588,N_14901,N_14898);
xor UO_1589 (O_1589,N_14951,N_14877);
and UO_1590 (O_1590,N_14889,N_14877);
and UO_1591 (O_1591,N_14942,N_14896);
nor UO_1592 (O_1592,N_14950,N_14855);
or UO_1593 (O_1593,N_14955,N_14872);
nor UO_1594 (O_1594,N_14985,N_14877);
nor UO_1595 (O_1595,N_14874,N_14908);
and UO_1596 (O_1596,N_14907,N_14966);
nand UO_1597 (O_1597,N_14932,N_14882);
or UO_1598 (O_1598,N_14990,N_14928);
nor UO_1599 (O_1599,N_14927,N_14934);
xnor UO_1600 (O_1600,N_14905,N_14895);
nor UO_1601 (O_1601,N_14883,N_14908);
or UO_1602 (O_1602,N_14868,N_14938);
nand UO_1603 (O_1603,N_14949,N_14950);
nor UO_1604 (O_1604,N_14885,N_14869);
nand UO_1605 (O_1605,N_14940,N_14895);
and UO_1606 (O_1606,N_14864,N_14857);
or UO_1607 (O_1607,N_14867,N_14925);
nand UO_1608 (O_1608,N_14887,N_14880);
and UO_1609 (O_1609,N_14941,N_14939);
nand UO_1610 (O_1610,N_14868,N_14917);
nor UO_1611 (O_1611,N_14982,N_14924);
and UO_1612 (O_1612,N_14964,N_14861);
or UO_1613 (O_1613,N_14952,N_14893);
nand UO_1614 (O_1614,N_14919,N_14862);
or UO_1615 (O_1615,N_14896,N_14945);
nand UO_1616 (O_1616,N_14921,N_14916);
nor UO_1617 (O_1617,N_14901,N_14994);
and UO_1618 (O_1618,N_14998,N_14934);
or UO_1619 (O_1619,N_14919,N_14923);
nor UO_1620 (O_1620,N_14946,N_14926);
nor UO_1621 (O_1621,N_14908,N_14905);
nand UO_1622 (O_1622,N_14999,N_14912);
xnor UO_1623 (O_1623,N_14963,N_14856);
nand UO_1624 (O_1624,N_14970,N_14979);
xnor UO_1625 (O_1625,N_14969,N_14895);
and UO_1626 (O_1626,N_14870,N_14916);
nand UO_1627 (O_1627,N_14855,N_14945);
and UO_1628 (O_1628,N_14997,N_14959);
nand UO_1629 (O_1629,N_14988,N_14870);
and UO_1630 (O_1630,N_14866,N_14918);
or UO_1631 (O_1631,N_14918,N_14882);
nand UO_1632 (O_1632,N_14907,N_14873);
nand UO_1633 (O_1633,N_14863,N_14992);
nand UO_1634 (O_1634,N_14945,N_14868);
nand UO_1635 (O_1635,N_14927,N_14907);
nor UO_1636 (O_1636,N_14994,N_14907);
and UO_1637 (O_1637,N_14972,N_14894);
xnor UO_1638 (O_1638,N_14968,N_14904);
nand UO_1639 (O_1639,N_14930,N_14954);
nand UO_1640 (O_1640,N_14980,N_14992);
or UO_1641 (O_1641,N_14859,N_14916);
or UO_1642 (O_1642,N_14962,N_14950);
nor UO_1643 (O_1643,N_14942,N_14958);
or UO_1644 (O_1644,N_14975,N_14974);
nor UO_1645 (O_1645,N_14990,N_14936);
and UO_1646 (O_1646,N_14964,N_14961);
nor UO_1647 (O_1647,N_14922,N_14858);
nor UO_1648 (O_1648,N_14938,N_14873);
xnor UO_1649 (O_1649,N_14964,N_14950);
nand UO_1650 (O_1650,N_14990,N_14946);
nor UO_1651 (O_1651,N_14929,N_14953);
and UO_1652 (O_1652,N_14897,N_14891);
and UO_1653 (O_1653,N_14967,N_14982);
nor UO_1654 (O_1654,N_14866,N_14939);
and UO_1655 (O_1655,N_14855,N_14913);
xor UO_1656 (O_1656,N_14976,N_14870);
and UO_1657 (O_1657,N_14908,N_14890);
or UO_1658 (O_1658,N_14851,N_14858);
or UO_1659 (O_1659,N_14876,N_14973);
nand UO_1660 (O_1660,N_14979,N_14899);
xor UO_1661 (O_1661,N_14913,N_14854);
or UO_1662 (O_1662,N_14967,N_14903);
nand UO_1663 (O_1663,N_14970,N_14936);
nand UO_1664 (O_1664,N_14943,N_14889);
xor UO_1665 (O_1665,N_14959,N_14947);
and UO_1666 (O_1666,N_14852,N_14892);
xnor UO_1667 (O_1667,N_14965,N_14989);
and UO_1668 (O_1668,N_14879,N_14883);
or UO_1669 (O_1669,N_14987,N_14932);
xnor UO_1670 (O_1670,N_14865,N_14873);
nand UO_1671 (O_1671,N_14933,N_14937);
or UO_1672 (O_1672,N_14949,N_14903);
or UO_1673 (O_1673,N_14913,N_14950);
xnor UO_1674 (O_1674,N_14912,N_14945);
or UO_1675 (O_1675,N_14904,N_14999);
xor UO_1676 (O_1676,N_14996,N_14926);
and UO_1677 (O_1677,N_14919,N_14980);
nor UO_1678 (O_1678,N_14852,N_14940);
nand UO_1679 (O_1679,N_14991,N_14978);
xnor UO_1680 (O_1680,N_14949,N_14930);
xnor UO_1681 (O_1681,N_14897,N_14870);
or UO_1682 (O_1682,N_14910,N_14914);
nand UO_1683 (O_1683,N_14964,N_14852);
and UO_1684 (O_1684,N_14964,N_14917);
xor UO_1685 (O_1685,N_14913,N_14887);
xor UO_1686 (O_1686,N_14967,N_14936);
nand UO_1687 (O_1687,N_14935,N_14938);
xor UO_1688 (O_1688,N_14874,N_14897);
nand UO_1689 (O_1689,N_14941,N_14881);
and UO_1690 (O_1690,N_14903,N_14892);
or UO_1691 (O_1691,N_14901,N_14882);
nand UO_1692 (O_1692,N_14996,N_14857);
nor UO_1693 (O_1693,N_14959,N_14920);
xnor UO_1694 (O_1694,N_14933,N_14989);
xnor UO_1695 (O_1695,N_14950,N_14918);
and UO_1696 (O_1696,N_14945,N_14911);
nor UO_1697 (O_1697,N_14935,N_14895);
nand UO_1698 (O_1698,N_14952,N_14883);
nor UO_1699 (O_1699,N_14909,N_14930);
nor UO_1700 (O_1700,N_14859,N_14970);
nand UO_1701 (O_1701,N_14938,N_14957);
nand UO_1702 (O_1702,N_14908,N_14999);
and UO_1703 (O_1703,N_14948,N_14973);
xor UO_1704 (O_1704,N_14955,N_14908);
nor UO_1705 (O_1705,N_14934,N_14912);
or UO_1706 (O_1706,N_14945,N_14994);
xnor UO_1707 (O_1707,N_14942,N_14871);
or UO_1708 (O_1708,N_14929,N_14901);
nand UO_1709 (O_1709,N_14995,N_14910);
nand UO_1710 (O_1710,N_14944,N_14920);
nand UO_1711 (O_1711,N_14869,N_14992);
xor UO_1712 (O_1712,N_14924,N_14928);
or UO_1713 (O_1713,N_14992,N_14910);
nor UO_1714 (O_1714,N_14976,N_14873);
nand UO_1715 (O_1715,N_14945,N_14907);
nor UO_1716 (O_1716,N_14968,N_14983);
nor UO_1717 (O_1717,N_14952,N_14874);
nand UO_1718 (O_1718,N_14852,N_14962);
nand UO_1719 (O_1719,N_14929,N_14922);
nor UO_1720 (O_1720,N_14940,N_14900);
nor UO_1721 (O_1721,N_14954,N_14951);
or UO_1722 (O_1722,N_14994,N_14863);
nand UO_1723 (O_1723,N_14964,N_14873);
and UO_1724 (O_1724,N_14965,N_14924);
nor UO_1725 (O_1725,N_14967,N_14944);
xor UO_1726 (O_1726,N_14999,N_14998);
or UO_1727 (O_1727,N_14855,N_14972);
nand UO_1728 (O_1728,N_14889,N_14974);
or UO_1729 (O_1729,N_14916,N_14893);
nor UO_1730 (O_1730,N_14881,N_14991);
or UO_1731 (O_1731,N_14891,N_14888);
xnor UO_1732 (O_1732,N_14935,N_14974);
and UO_1733 (O_1733,N_14947,N_14917);
nor UO_1734 (O_1734,N_14939,N_14878);
nor UO_1735 (O_1735,N_14992,N_14951);
nor UO_1736 (O_1736,N_14886,N_14895);
xnor UO_1737 (O_1737,N_14858,N_14953);
nand UO_1738 (O_1738,N_14924,N_14855);
nand UO_1739 (O_1739,N_14872,N_14912);
xnor UO_1740 (O_1740,N_14943,N_14971);
xor UO_1741 (O_1741,N_14896,N_14948);
xnor UO_1742 (O_1742,N_14924,N_14991);
or UO_1743 (O_1743,N_14909,N_14886);
xnor UO_1744 (O_1744,N_14863,N_14871);
xor UO_1745 (O_1745,N_14927,N_14978);
nand UO_1746 (O_1746,N_14943,N_14978);
and UO_1747 (O_1747,N_14859,N_14926);
nand UO_1748 (O_1748,N_14932,N_14924);
nand UO_1749 (O_1749,N_14941,N_14982);
nand UO_1750 (O_1750,N_14904,N_14945);
and UO_1751 (O_1751,N_14882,N_14944);
nor UO_1752 (O_1752,N_14984,N_14910);
or UO_1753 (O_1753,N_14913,N_14858);
xnor UO_1754 (O_1754,N_14976,N_14853);
xnor UO_1755 (O_1755,N_14895,N_14892);
nor UO_1756 (O_1756,N_14914,N_14852);
and UO_1757 (O_1757,N_14968,N_14912);
nand UO_1758 (O_1758,N_14963,N_14999);
nor UO_1759 (O_1759,N_14924,N_14993);
nand UO_1760 (O_1760,N_14939,N_14867);
xnor UO_1761 (O_1761,N_14938,N_14939);
xnor UO_1762 (O_1762,N_14895,N_14903);
or UO_1763 (O_1763,N_14894,N_14954);
and UO_1764 (O_1764,N_14913,N_14924);
or UO_1765 (O_1765,N_14977,N_14890);
or UO_1766 (O_1766,N_14897,N_14900);
nand UO_1767 (O_1767,N_14997,N_14904);
xor UO_1768 (O_1768,N_14990,N_14974);
xnor UO_1769 (O_1769,N_14928,N_14955);
xor UO_1770 (O_1770,N_14936,N_14986);
nand UO_1771 (O_1771,N_14956,N_14915);
and UO_1772 (O_1772,N_14898,N_14984);
nor UO_1773 (O_1773,N_14864,N_14976);
and UO_1774 (O_1774,N_14926,N_14992);
and UO_1775 (O_1775,N_14940,N_14945);
or UO_1776 (O_1776,N_14962,N_14851);
nand UO_1777 (O_1777,N_14920,N_14998);
xnor UO_1778 (O_1778,N_14931,N_14955);
or UO_1779 (O_1779,N_14878,N_14998);
or UO_1780 (O_1780,N_14963,N_14934);
xnor UO_1781 (O_1781,N_14875,N_14943);
xnor UO_1782 (O_1782,N_14873,N_14928);
or UO_1783 (O_1783,N_14890,N_14894);
xor UO_1784 (O_1784,N_14976,N_14947);
and UO_1785 (O_1785,N_14900,N_14984);
and UO_1786 (O_1786,N_14866,N_14968);
nor UO_1787 (O_1787,N_14946,N_14975);
xor UO_1788 (O_1788,N_14995,N_14855);
xor UO_1789 (O_1789,N_14996,N_14933);
nor UO_1790 (O_1790,N_14909,N_14963);
xor UO_1791 (O_1791,N_14979,N_14940);
nor UO_1792 (O_1792,N_14969,N_14999);
or UO_1793 (O_1793,N_14866,N_14878);
or UO_1794 (O_1794,N_14968,N_14916);
nor UO_1795 (O_1795,N_14920,N_14881);
xnor UO_1796 (O_1796,N_14988,N_14905);
and UO_1797 (O_1797,N_14972,N_14951);
nor UO_1798 (O_1798,N_14950,N_14927);
xnor UO_1799 (O_1799,N_14916,N_14993);
xnor UO_1800 (O_1800,N_14897,N_14997);
xor UO_1801 (O_1801,N_14859,N_14907);
nand UO_1802 (O_1802,N_14971,N_14920);
and UO_1803 (O_1803,N_14880,N_14974);
nor UO_1804 (O_1804,N_14930,N_14868);
or UO_1805 (O_1805,N_14959,N_14876);
nor UO_1806 (O_1806,N_14948,N_14866);
xnor UO_1807 (O_1807,N_14917,N_14948);
nor UO_1808 (O_1808,N_14904,N_14956);
xor UO_1809 (O_1809,N_14919,N_14880);
xnor UO_1810 (O_1810,N_14934,N_14881);
nand UO_1811 (O_1811,N_14872,N_14964);
nor UO_1812 (O_1812,N_14904,N_14855);
nor UO_1813 (O_1813,N_14946,N_14864);
xor UO_1814 (O_1814,N_14889,N_14885);
nor UO_1815 (O_1815,N_14893,N_14939);
and UO_1816 (O_1816,N_14876,N_14996);
nor UO_1817 (O_1817,N_14945,N_14942);
or UO_1818 (O_1818,N_14898,N_14885);
and UO_1819 (O_1819,N_14904,N_14863);
or UO_1820 (O_1820,N_14993,N_14996);
nand UO_1821 (O_1821,N_14852,N_14927);
xnor UO_1822 (O_1822,N_14992,N_14940);
xor UO_1823 (O_1823,N_14866,N_14915);
nand UO_1824 (O_1824,N_14997,N_14947);
or UO_1825 (O_1825,N_14958,N_14917);
nor UO_1826 (O_1826,N_14977,N_14920);
nand UO_1827 (O_1827,N_14869,N_14979);
and UO_1828 (O_1828,N_14980,N_14941);
or UO_1829 (O_1829,N_14935,N_14962);
xor UO_1830 (O_1830,N_14874,N_14982);
nand UO_1831 (O_1831,N_14976,N_14961);
nand UO_1832 (O_1832,N_14953,N_14898);
or UO_1833 (O_1833,N_14920,N_14882);
nand UO_1834 (O_1834,N_14871,N_14915);
or UO_1835 (O_1835,N_14997,N_14863);
xnor UO_1836 (O_1836,N_14918,N_14919);
nor UO_1837 (O_1837,N_14855,N_14967);
nand UO_1838 (O_1838,N_14852,N_14863);
and UO_1839 (O_1839,N_14865,N_14908);
nand UO_1840 (O_1840,N_14879,N_14903);
nor UO_1841 (O_1841,N_14889,N_14969);
nand UO_1842 (O_1842,N_14924,N_14921);
or UO_1843 (O_1843,N_14992,N_14860);
nand UO_1844 (O_1844,N_14924,N_14995);
xnor UO_1845 (O_1845,N_14906,N_14919);
and UO_1846 (O_1846,N_14967,N_14931);
and UO_1847 (O_1847,N_14930,N_14902);
xnor UO_1848 (O_1848,N_14935,N_14881);
and UO_1849 (O_1849,N_14915,N_14864);
or UO_1850 (O_1850,N_14959,N_14860);
nor UO_1851 (O_1851,N_14879,N_14947);
nand UO_1852 (O_1852,N_14854,N_14887);
nand UO_1853 (O_1853,N_14916,N_14868);
or UO_1854 (O_1854,N_14921,N_14854);
xor UO_1855 (O_1855,N_14928,N_14997);
and UO_1856 (O_1856,N_14937,N_14920);
nor UO_1857 (O_1857,N_14974,N_14856);
nor UO_1858 (O_1858,N_14900,N_14992);
or UO_1859 (O_1859,N_14907,N_14955);
and UO_1860 (O_1860,N_14894,N_14975);
or UO_1861 (O_1861,N_14959,N_14985);
or UO_1862 (O_1862,N_14936,N_14923);
nor UO_1863 (O_1863,N_14949,N_14876);
or UO_1864 (O_1864,N_14874,N_14980);
nand UO_1865 (O_1865,N_14855,N_14881);
and UO_1866 (O_1866,N_14925,N_14887);
xor UO_1867 (O_1867,N_14993,N_14991);
xor UO_1868 (O_1868,N_14891,N_14929);
nor UO_1869 (O_1869,N_14852,N_14987);
and UO_1870 (O_1870,N_14978,N_14855);
nor UO_1871 (O_1871,N_14988,N_14909);
nor UO_1872 (O_1872,N_14990,N_14989);
xor UO_1873 (O_1873,N_14972,N_14974);
or UO_1874 (O_1874,N_14890,N_14912);
or UO_1875 (O_1875,N_14968,N_14925);
or UO_1876 (O_1876,N_14966,N_14910);
nand UO_1877 (O_1877,N_14976,N_14868);
nor UO_1878 (O_1878,N_14918,N_14996);
and UO_1879 (O_1879,N_14944,N_14876);
and UO_1880 (O_1880,N_14973,N_14933);
or UO_1881 (O_1881,N_14996,N_14925);
and UO_1882 (O_1882,N_14940,N_14997);
nor UO_1883 (O_1883,N_14989,N_14914);
nor UO_1884 (O_1884,N_14875,N_14908);
xor UO_1885 (O_1885,N_14852,N_14938);
and UO_1886 (O_1886,N_14973,N_14908);
and UO_1887 (O_1887,N_14854,N_14930);
xnor UO_1888 (O_1888,N_14965,N_14987);
or UO_1889 (O_1889,N_14995,N_14926);
or UO_1890 (O_1890,N_14875,N_14966);
nand UO_1891 (O_1891,N_14910,N_14889);
xnor UO_1892 (O_1892,N_14875,N_14863);
or UO_1893 (O_1893,N_14977,N_14991);
xnor UO_1894 (O_1894,N_14878,N_14854);
xnor UO_1895 (O_1895,N_14996,N_14938);
nor UO_1896 (O_1896,N_14989,N_14946);
or UO_1897 (O_1897,N_14989,N_14997);
and UO_1898 (O_1898,N_14886,N_14914);
nand UO_1899 (O_1899,N_14997,N_14908);
nor UO_1900 (O_1900,N_14883,N_14926);
nand UO_1901 (O_1901,N_14948,N_14991);
nand UO_1902 (O_1902,N_14959,N_14917);
or UO_1903 (O_1903,N_14902,N_14929);
nand UO_1904 (O_1904,N_14973,N_14864);
or UO_1905 (O_1905,N_14852,N_14973);
nor UO_1906 (O_1906,N_14870,N_14999);
xnor UO_1907 (O_1907,N_14886,N_14856);
and UO_1908 (O_1908,N_14867,N_14983);
xnor UO_1909 (O_1909,N_14926,N_14862);
nor UO_1910 (O_1910,N_14887,N_14933);
xnor UO_1911 (O_1911,N_14987,N_14940);
or UO_1912 (O_1912,N_14936,N_14882);
nand UO_1913 (O_1913,N_14925,N_14933);
or UO_1914 (O_1914,N_14895,N_14949);
and UO_1915 (O_1915,N_14869,N_14964);
xor UO_1916 (O_1916,N_14952,N_14924);
xor UO_1917 (O_1917,N_14951,N_14895);
nand UO_1918 (O_1918,N_14933,N_14920);
nor UO_1919 (O_1919,N_14877,N_14941);
or UO_1920 (O_1920,N_14852,N_14970);
and UO_1921 (O_1921,N_14959,N_14866);
xnor UO_1922 (O_1922,N_14947,N_14970);
nor UO_1923 (O_1923,N_14908,N_14967);
nand UO_1924 (O_1924,N_14973,N_14928);
or UO_1925 (O_1925,N_14926,N_14912);
xnor UO_1926 (O_1926,N_14993,N_14945);
and UO_1927 (O_1927,N_14882,N_14891);
nand UO_1928 (O_1928,N_14970,N_14930);
and UO_1929 (O_1929,N_14967,N_14871);
nor UO_1930 (O_1930,N_14867,N_14891);
or UO_1931 (O_1931,N_14877,N_14991);
nand UO_1932 (O_1932,N_14906,N_14979);
xor UO_1933 (O_1933,N_14971,N_14935);
nor UO_1934 (O_1934,N_14885,N_14896);
nand UO_1935 (O_1935,N_14872,N_14892);
and UO_1936 (O_1936,N_14919,N_14976);
or UO_1937 (O_1937,N_14851,N_14864);
nor UO_1938 (O_1938,N_14950,N_14870);
or UO_1939 (O_1939,N_14951,N_14850);
nor UO_1940 (O_1940,N_14859,N_14929);
nand UO_1941 (O_1941,N_14944,N_14862);
nor UO_1942 (O_1942,N_14931,N_14932);
and UO_1943 (O_1943,N_14996,N_14973);
nand UO_1944 (O_1944,N_14958,N_14988);
and UO_1945 (O_1945,N_14980,N_14951);
xnor UO_1946 (O_1946,N_14869,N_14920);
nand UO_1947 (O_1947,N_14964,N_14853);
nor UO_1948 (O_1948,N_14915,N_14913);
or UO_1949 (O_1949,N_14910,N_14996);
nor UO_1950 (O_1950,N_14994,N_14886);
and UO_1951 (O_1951,N_14999,N_14877);
xnor UO_1952 (O_1952,N_14959,N_14977);
nand UO_1953 (O_1953,N_14864,N_14904);
and UO_1954 (O_1954,N_14894,N_14998);
xor UO_1955 (O_1955,N_14871,N_14979);
xor UO_1956 (O_1956,N_14965,N_14949);
or UO_1957 (O_1957,N_14900,N_14996);
or UO_1958 (O_1958,N_14925,N_14868);
nand UO_1959 (O_1959,N_14962,N_14924);
xnor UO_1960 (O_1960,N_14973,N_14867);
xnor UO_1961 (O_1961,N_14865,N_14906);
and UO_1962 (O_1962,N_14994,N_14880);
or UO_1963 (O_1963,N_14908,N_14881);
xor UO_1964 (O_1964,N_14986,N_14962);
or UO_1965 (O_1965,N_14966,N_14933);
xnor UO_1966 (O_1966,N_14987,N_14898);
nand UO_1967 (O_1967,N_14945,N_14854);
or UO_1968 (O_1968,N_14935,N_14961);
nand UO_1969 (O_1969,N_14903,N_14872);
xnor UO_1970 (O_1970,N_14929,N_14993);
xnor UO_1971 (O_1971,N_14877,N_14920);
and UO_1972 (O_1972,N_14939,N_14981);
and UO_1973 (O_1973,N_14888,N_14999);
and UO_1974 (O_1974,N_14969,N_14933);
nor UO_1975 (O_1975,N_14997,N_14906);
nand UO_1976 (O_1976,N_14853,N_14998);
nand UO_1977 (O_1977,N_14929,N_14855);
xor UO_1978 (O_1978,N_14881,N_14985);
or UO_1979 (O_1979,N_14951,N_14926);
and UO_1980 (O_1980,N_14874,N_14881);
xnor UO_1981 (O_1981,N_14891,N_14884);
nand UO_1982 (O_1982,N_14983,N_14947);
nand UO_1983 (O_1983,N_14925,N_14948);
or UO_1984 (O_1984,N_14865,N_14973);
nor UO_1985 (O_1985,N_14933,N_14871);
nand UO_1986 (O_1986,N_14953,N_14970);
xnor UO_1987 (O_1987,N_14964,N_14954);
or UO_1988 (O_1988,N_14867,N_14991);
and UO_1989 (O_1989,N_14942,N_14866);
and UO_1990 (O_1990,N_14913,N_14953);
nand UO_1991 (O_1991,N_14893,N_14961);
and UO_1992 (O_1992,N_14966,N_14980);
xnor UO_1993 (O_1993,N_14992,N_14916);
xor UO_1994 (O_1994,N_14933,N_14983);
nor UO_1995 (O_1995,N_14963,N_14907);
xor UO_1996 (O_1996,N_14929,N_14987);
xor UO_1997 (O_1997,N_14981,N_14891);
nor UO_1998 (O_1998,N_14877,N_14954);
nor UO_1999 (O_1999,N_14870,N_14850);
endmodule