module basic_500_3000_500_30_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_84,In_367);
and U1 (N_1,In_377,In_359);
nor U2 (N_2,In_81,In_270);
nor U3 (N_3,In_424,In_383);
nor U4 (N_4,In_39,In_147);
nor U5 (N_5,In_490,In_326);
nand U6 (N_6,In_24,In_355);
nand U7 (N_7,In_465,In_25);
nor U8 (N_8,In_427,In_276);
and U9 (N_9,In_64,In_480);
nand U10 (N_10,In_152,In_482);
and U11 (N_11,In_341,In_145);
and U12 (N_12,In_325,In_305);
nor U13 (N_13,In_259,In_193);
nor U14 (N_14,In_393,In_99);
nor U15 (N_15,In_257,In_202);
nor U16 (N_16,In_345,In_352);
or U17 (N_17,In_183,In_18);
nor U18 (N_18,In_115,In_440);
nand U19 (N_19,In_336,In_309);
nand U20 (N_20,In_229,In_131);
or U21 (N_21,In_250,In_220);
or U22 (N_22,In_174,In_179);
or U23 (N_23,In_41,In_280);
nand U24 (N_24,In_247,In_211);
nor U25 (N_25,In_304,In_2);
and U26 (N_26,In_258,In_187);
or U27 (N_27,In_101,In_429);
or U28 (N_28,In_37,In_76);
or U29 (N_29,In_201,In_374);
nand U30 (N_30,In_303,In_119);
nand U31 (N_31,In_172,In_290);
nand U32 (N_32,In_88,In_185);
xnor U33 (N_33,In_168,In_292);
nor U34 (N_34,In_379,In_239);
and U35 (N_35,In_112,In_46);
xor U36 (N_36,In_8,In_364);
or U37 (N_37,In_333,In_230);
xor U38 (N_38,In_446,In_478);
and U39 (N_39,In_488,In_432);
and U40 (N_40,In_436,In_36);
or U41 (N_41,In_10,In_254);
or U42 (N_42,In_418,In_205);
or U43 (N_43,In_256,In_159);
or U44 (N_44,In_176,In_396);
or U45 (N_45,In_195,In_394);
xor U46 (N_46,In_49,In_302);
xor U47 (N_47,In_189,In_380);
and U48 (N_48,In_126,In_332);
and U49 (N_49,In_154,In_27);
xnor U50 (N_50,In_12,In_426);
nor U51 (N_51,In_19,In_80);
nor U52 (N_52,In_70,In_151);
nand U53 (N_53,In_32,In_44);
nand U54 (N_54,In_261,In_219);
nor U55 (N_55,In_221,In_362);
nand U56 (N_56,In_338,In_199);
xor U57 (N_57,In_372,In_373);
xor U58 (N_58,In_417,In_416);
nand U59 (N_59,In_233,In_390);
xnor U60 (N_60,In_387,In_375);
and U61 (N_61,In_59,In_441);
nor U62 (N_62,In_58,In_82);
nand U63 (N_63,In_241,In_384);
or U64 (N_64,In_125,In_100);
xor U65 (N_65,In_334,In_213);
nand U66 (N_66,In_356,In_231);
xor U67 (N_67,In_102,In_210);
or U68 (N_68,In_28,In_425);
or U69 (N_69,In_204,In_78);
xor U70 (N_70,In_354,In_408);
nand U71 (N_71,In_170,In_473);
or U72 (N_72,In_83,In_472);
or U73 (N_73,In_128,In_243);
nand U74 (N_74,In_263,In_272);
and U75 (N_75,In_327,In_53);
and U76 (N_76,In_21,In_225);
xor U77 (N_77,In_497,In_422);
xnor U78 (N_78,In_1,In_16);
nand U79 (N_79,In_207,In_435);
nand U80 (N_80,In_411,In_349);
nand U81 (N_81,In_124,In_66);
nand U82 (N_82,In_34,In_97);
nand U83 (N_83,In_85,In_454);
or U84 (N_84,In_395,In_378);
and U85 (N_85,In_5,In_200);
nand U86 (N_86,In_388,In_42);
nand U87 (N_87,In_52,In_47);
or U88 (N_88,In_463,In_437);
nand U89 (N_89,In_228,In_319);
or U90 (N_90,In_314,In_245);
nor U91 (N_91,In_363,In_468);
nand U92 (N_92,In_48,In_289);
xnor U93 (N_93,In_281,In_191);
nor U94 (N_94,In_246,In_320);
nand U95 (N_95,In_452,In_471);
nand U96 (N_96,In_121,In_392);
or U97 (N_97,In_20,In_316);
xor U98 (N_98,In_123,In_38);
and U99 (N_99,In_114,In_353);
or U100 (N_100,N_30,N_42);
xor U101 (N_101,In_188,In_376);
nor U102 (N_102,In_265,N_86);
xnor U103 (N_103,N_85,In_266);
nand U104 (N_104,N_61,In_344);
and U105 (N_105,N_68,In_167);
nand U106 (N_106,In_160,In_237);
nand U107 (N_107,In_89,In_90);
and U108 (N_108,In_50,In_491);
xor U109 (N_109,N_84,In_14);
nor U110 (N_110,In_158,In_461);
xor U111 (N_111,In_318,N_83);
nand U112 (N_112,In_448,In_430);
nor U113 (N_113,In_389,In_391);
nor U114 (N_114,In_234,In_442);
and U115 (N_115,N_44,In_120);
nor U116 (N_116,In_456,In_148);
or U117 (N_117,In_339,N_89);
and U118 (N_118,In_227,In_475);
and U119 (N_119,In_129,In_369);
or U120 (N_120,In_209,In_87);
nor U121 (N_121,N_21,In_94);
and U122 (N_122,In_98,In_68);
nand U123 (N_123,In_141,N_48);
nand U124 (N_124,In_322,In_255);
nor U125 (N_125,N_97,In_153);
nand U126 (N_126,In_409,In_342);
or U127 (N_127,N_77,N_60);
or U128 (N_128,N_92,In_324);
nand U129 (N_129,N_47,In_118);
nor U130 (N_130,N_35,In_312);
and U131 (N_131,In_136,In_69);
nor U132 (N_132,In_65,In_335);
or U133 (N_133,In_150,In_43);
xnor U134 (N_134,In_370,In_190);
or U135 (N_135,N_13,In_365);
and U136 (N_136,In_177,N_9);
nand U137 (N_137,In_445,N_96);
nor U138 (N_138,In_130,In_11);
nand U139 (N_139,In_343,In_400);
or U140 (N_140,In_328,N_70);
and U141 (N_141,In_157,In_419);
or U142 (N_142,N_11,In_61);
or U143 (N_143,In_346,In_13);
and U144 (N_144,In_348,In_110);
and U145 (N_145,In_453,In_212);
or U146 (N_146,In_23,In_404);
or U147 (N_147,In_171,In_3);
nand U148 (N_148,In_73,N_53);
nor U149 (N_149,In_6,N_8);
and U150 (N_150,N_43,In_311);
and U151 (N_151,In_279,In_351);
or U152 (N_152,N_52,In_51);
nor U153 (N_153,In_186,In_358);
nor U154 (N_154,In_248,In_499);
or U155 (N_155,In_40,In_460);
and U156 (N_156,N_17,In_149);
xnor U157 (N_157,N_32,In_0);
or U158 (N_158,In_242,In_477);
or U159 (N_159,In_226,In_218);
or U160 (N_160,N_55,In_108);
or U161 (N_161,In_414,N_78);
xor U162 (N_162,In_371,In_252);
or U163 (N_163,In_412,In_135);
nand U164 (N_164,In_466,In_79);
xor U165 (N_165,N_36,N_62);
and U166 (N_166,N_28,In_143);
nand U167 (N_167,In_262,In_476);
nor U168 (N_168,In_405,N_23);
xnor U169 (N_169,N_4,In_340);
nand U170 (N_170,In_274,In_268);
xnor U171 (N_171,In_295,In_33);
or U172 (N_172,In_57,In_317);
nand U173 (N_173,In_26,In_144);
xnor U174 (N_174,In_264,In_223);
xnor U175 (N_175,In_249,N_29);
nor U176 (N_176,In_155,In_483);
nand U177 (N_177,N_74,N_25);
or U178 (N_178,In_103,In_301);
nor U179 (N_179,In_308,N_63);
xnor U180 (N_180,N_0,In_30);
nor U181 (N_181,In_55,In_63);
and U182 (N_182,In_447,N_19);
or U183 (N_183,In_307,In_107);
xnor U184 (N_184,In_166,In_253);
and U185 (N_185,In_206,N_75);
nor U186 (N_186,N_49,In_493);
or U187 (N_187,N_15,N_20);
and U188 (N_188,In_434,In_357);
nand U189 (N_189,In_116,N_45);
or U190 (N_190,In_175,In_71);
nor U191 (N_191,In_180,In_485);
or U192 (N_192,In_306,N_57);
nand U193 (N_193,In_407,N_46);
xor U194 (N_194,In_169,In_277);
and U195 (N_195,In_457,N_67);
nand U196 (N_196,N_40,N_72);
xor U197 (N_197,In_122,In_4);
or U198 (N_198,N_88,In_215);
xnor U199 (N_199,N_38,In_496);
xor U200 (N_200,In_439,N_37);
and U201 (N_201,N_34,In_288);
nand U202 (N_202,In_208,N_100);
or U203 (N_203,N_176,N_95);
xor U204 (N_204,N_180,N_39);
xor U205 (N_205,In_132,N_113);
xnor U206 (N_206,In_31,In_35);
nor U207 (N_207,N_26,N_64);
nand U208 (N_208,N_87,N_181);
nand U209 (N_209,N_142,N_58);
nor U210 (N_210,N_59,In_109);
and U211 (N_211,N_71,In_7);
nor U212 (N_212,N_5,N_3);
xor U213 (N_213,In_299,N_151);
nand U214 (N_214,N_119,In_184);
xnor U215 (N_215,N_162,N_65);
nor U216 (N_216,N_2,In_410);
nor U217 (N_217,N_106,N_114);
xnor U218 (N_218,In_117,N_1);
xor U219 (N_219,In_397,N_121);
nor U220 (N_220,N_51,In_293);
nor U221 (N_221,N_50,N_16);
nand U222 (N_222,In_401,N_82);
or U223 (N_223,N_110,In_399);
or U224 (N_224,In_294,In_382);
or U225 (N_225,In_214,N_167);
nand U226 (N_226,In_240,N_197);
or U227 (N_227,In_481,N_138);
xnor U228 (N_228,In_474,In_321);
nor U229 (N_229,N_183,N_182);
and U230 (N_230,In_469,In_95);
or U231 (N_231,N_193,N_12);
or U232 (N_232,In_423,In_282);
xnor U233 (N_233,In_106,N_185);
nor U234 (N_234,In_450,In_287);
nand U235 (N_235,In_224,In_331);
xnor U236 (N_236,In_194,N_169);
xor U237 (N_237,In_164,In_310);
nor U238 (N_238,N_22,In_222);
nand U239 (N_239,In_91,N_168);
nand U240 (N_240,N_134,In_298);
nor U241 (N_241,In_96,N_157);
nor U242 (N_242,N_128,In_139);
nor U243 (N_243,In_415,In_217);
nand U244 (N_244,N_69,In_406);
nor U245 (N_245,N_148,N_108);
xor U246 (N_246,N_120,N_131);
nor U247 (N_247,N_54,N_135);
nand U248 (N_248,In_300,In_462);
and U249 (N_249,In_385,N_79);
and U250 (N_250,In_438,N_187);
and U251 (N_251,In_350,In_347);
and U252 (N_252,In_484,In_402);
nor U253 (N_253,In_464,In_486);
nor U254 (N_254,N_179,In_232);
or U255 (N_255,In_146,In_467);
nand U256 (N_256,In_420,N_190);
xor U257 (N_257,N_150,N_170);
or U258 (N_258,N_166,In_444);
xor U259 (N_259,In_75,In_421);
or U260 (N_260,N_126,N_104);
nor U261 (N_261,In_92,In_271);
or U262 (N_262,In_15,N_125);
nand U263 (N_263,In_86,In_9);
and U264 (N_264,N_24,N_124);
and U265 (N_265,N_115,In_291);
nand U266 (N_266,In_386,N_172);
and U267 (N_267,N_143,In_360);
xor U268 (N_268,In_113,In_297);
xnor U269 (N_269,In_162,N_99);
nor U270 (N_270,In_313,In_330);
and U271 (N_271,In_329,In_45);
nand U272 (N_272,In_156,In_29);
and U273 (N_273,In_56,N_158);
nor U274 (N_274,In_337,N_139);
xor U275 (N_275,In_451,In_93);
nand U276 (N_276,In_197,In_428);
nor U277 (N_277,In_494,N_80);
nor U278 (N_278,In_251,N_111);
and U279 (N_279,N_198,In_489);
nor U280 (N_280,N_152,In_296);
nand U281 (N_281,N_33,N_154);
and U282 (N_282,In_181,N_14);
or U283 (N_283,N_199,In_244);
nor U284 (N_284,N_27,In_449);
nand U285 (N_285,N_116,N_159);
xnor U286 (N_286,In_192,In_161);
nor U287 (N_287,N_98,N_173);
nor U288 (N_288,N_186,In_498);
xnor U289 (N_289,In_142,N_164);
xor U290 (N_290,N_129,N_31);
nor U291 (N_291,In_140,N_188);
xnor U292 (N_292,In_163,N_178);
or U293 (N_293,N_189,In_238);
or U294 (N_294,N_160,In_470);
nor U295 (N_295,In_17,In_105);
xor U296 (N_296,N_191,N_165);
or U297 (N_297,In_137,In_286);
nor U298 (N_298,N_91,In_198);
nand U299 (N_299,N_118,N_132);
nor U300 (N_300,N_201,N_205);
nand U301 (N_301,N_6,N_297);
or U302 (N_302,In_196,N_93);
nor U303 (N_303,In_134,N_221);
and U304 (N_304,N_281,In_495);
nand U305 (N_305,In_111,In_492);
or U306 (N_306,N_252,In_74);
nor U307 (N_307,In_273,N_231);
and U308 (N_308,N_253,N_7);
and U309 (N_309,N_271,In_487);
or U310 (N_310,N_163,N_296);
nand U311 (N_311,N_226,N_267);
xnor U312 (N_312,N_174,N_216);
or U313 (N_313,N_256,N_222);
xor U314 (N_314,In_67,N_250);
nand U315 (N_315,N_141,N_171);
and U316 (N_316,In_323,N_268);
nor U317 (N_317,N_280,In_62);
xnor U318 (N_318,In_284,N_155);
and U319 (N_319,N_261,N_215);
or U320 (N_320,N_229,N_290);
or U321 (N_321,N_230,N_282);
nand U322 (N_322,In_54,N_260);
nor U323 (N_323,N_293,N_249);
and U324 (N_324,In_403,In_22);
nand U325 (N_325,In_283,N_140);
nand U326 (N_326,N_184,In_138);
nand U327 (N_327,N_90,N_10);
and U328 (N_328,N_262,N_136);
or U329 (N_329,In_315,N_177);
xor U330 (N_330,N_240,N_130);
nand U331 (N_331,In_72,N_291);
and U332 (N_332,N_105,N_257);
or U333 (N_333,In_366,N_245);
or U334 (N_334,N_127,N_73);
and U335 (N_335,N_202,N_219);
and U336 (N_336,N_234,In_236);
xnor U337 (N_337,N_287,N_208);
or U338 (N_338,N_41,N_195);
xnor U339 (N_339,N_273,N_224);
xnor U340 (N_340,In_459,N_103);
nand U341 (N_341,In_235,In_285);
or U342 (N_342,N_145,N_233);
or U343 (N_343,N_235,N_192);
nor U344 (N_344,N_212,N_292);
or U345 (N_345,N_238,N_269);
nor U346 (N_346,N_223,N_289);
nand U347 (N_347,N_76,N_241);
nand U348 (N_348,N_200,N_206);
xor U349 (N_349,N_214,N_258);
xnor U350 (N_350,N_112,N_210);
nand U351 (N_351,N_217,N_255);
nor U352 (N_352,N_213,N_101);
nand U353 (N_353,In_398,In_413);
or U354 (N_354,N_94,In_260);
or U355 (N_355,N_144,N_275);
xor U356 (N_356,N_56,N_227);
nand U357 (N_357,N_264,N_203);
and U358 (N_358,In_178,N_149);
xnor U359 (N_359,N_66,N_107);
xnor U360 (N_360,N_243,N_156);
nand U361 (N_361,In_165,N_299);
xnor U362 (N_362,N_146,N_220);
nor U363 (N_363,In_275,N_246);
and U364 (N_364,N_218,N_286);
and U365 (N_365,N_247,In_455);
nand U366 (N_366,In_104,N_196);
nand U367 (N_367,N_265,N_161);
and U368 (N_368,N_123,N_109);
nand U369 (N_369,N_263,N_254);
nand U370 (N_370,N_137,In_458);
or U371 (N_371,N_266,N_133);
nand U372 (N_372,In_203,N_279);
and U373 (N_373,N_18,N_284);
nor U374 (N_374,In_269,N_207);
xor U375 (N_375,In_431,N_147);
and U376 (N_376,N_194,N_272);
nand U377 (N_377,In_433,N_276);
xnor U378 (N_378,N_175,N_211);
nor U379 (N_379,N_236,N_122);
or U380 (N_380,In_77,In_361);
and U381 (N_381,N_228,N_298);
and U382 (N_382,In_216,In_443);
and U383 (N_383,N_232,In_267);
xnor U384 (N_384,N_270,N_295);
or U385 (N_385,In_479,In_182);
nand U386 (N_386,N_283,N_244);
nand U387 (N_387,In_127,N_274);
xor U388 (N_388,N_294,In_173);
and U389 (N_389,N_277,N_248);
nand U390 (N_390,N_285,N_259);
or U391 (N_391,N_239,N_278);
xnor U392 (N_392,N_204,In_368);
nand U393 (N_393,N_251,N_225);
nand U394 (N_394,N_102,In_278);
and U395 (N_395,N_81,N_288);
nor U396 (N_396,N_153,In_60);
nand U397 (N_397,In_133,N_117);
nand U398 (N_398,In_381,N_242);
xor U399 (N_399,N_209,N_237);
and U400 (N_400,N_328,N_347);
and U401 (N_401,N_360,N_337);
or U402 (N_402,N_317,N_389);
or U403 (N_403,N_398,N_370);
nor U404 (N_404,N_330,N_373);
xnor U405 (N_405,N_312,N_362);
xnor U406 (N_406,N_352,N_380);
nor U407 (N_407,N_315,N_381);
xnor U408 (N_408,N_343,N_369);
nand U409 (N_409,N_364,N_319);
or U410 (N_410,N_372,N_320);
xor U411 (N_411,N_358,N_376);
xnor U412 (N_412,N_354,N_357);
nand U413 (N_413,N_333,N_327);
nor U414 (N_414,N_386,N_396);
nand U415 (N_415,N_385,N_378);
xor U416 (N_416,N_325,N_321);
nor U417 (N_417,N_371,N_301);
nand U418 (N_418,N_390,N_311);
nand U419 (N_419,N_375,N_365);
and U420 (N_420,N_305,N_382);
or U421 (N_421,N_367,N_310);
nor U422 (N_422,N_314,N_383);
and U423 (N_423,N_306,N_329);
and U424 (N_424,N_338,N_350);
nand U425 (N_425,N_302,N_339);
nand U426 (N_426,N_309,N_303);
and U427 (N_427,N_391,N_341);
nor U428 (N_428,N_334,N_313);
nand U429 (N_429,N_395,N_349);
xnor U430 (N_430,N_392,N_366);
and U431 (N_431,N_387,N_353);
and U432 (N_432,N_324,N_331);
xor U433 (N_433,N_332,N_316);
nand U434 (N_434,N_368,N_336);
nand U435 (N_435,N_394,N_326);
xnor U436 (N_436,N_384,N_318);
nor U437 (N_437,N_359,N_342);
or U438 (N_438,N_377,N_399);
nand U439 (N_439,N_308,N_322);
and U440 (N_440,N_344,N_355);
and U441 (N_441,N_351,N_323);
and U442 (N_442,N_361,N_388);
and U443 (N_443,N_340,N_345);
xor U444 (N_444,N_356,N_304);
nor U445 (N_445,N_348,N_346);
xnor U446 (N_446,N_379,N_307);
or U447 (N_447,N_393,N_397);
xor U448 (N_448,N_300,N_335);
xor U449 (N_449,N_363,N_374);
xor U450 (N_450,N_323,N_366);
xor U451 (N_451,N_335,N_318);
or U452 (N_452,N_330,N_393);
nand U453 (N_453,N_345,N_323);
and U454 (N_454,N_373,N_387);
nand U455 (N_455,N_319,N_361);
nand U456 (N_456,N_309,N_393);
xor U457 (N_457,N_336,N_313);
nand U458 (N_458,N_396,N_363);
or U459 (N_459,N_372,N_334);
and U460 (N_460,N_365,N_337);
nand U461 (N_461,N_323,N_308);
nand U462 (N_462,N_395,N_341);
xnor U463 (N_463,N_389,N_377);
nor U464 (N_464,N_310,N_369);
xor U465 (N_465,N_369,N_335);
nor U466 (N_466,N_372,N_330);
xnor U467 (N_467,N_313,N_357);
or U468 (N_468,N_334,N_353);
xnor U469 (N_469,N_369,N_349);
and U470 (N_470,N_353,N_314);
and U471 (N_471,N_316,N_330);
nand U472 (N_472,N_341,N_348);
and U473 (N_473,N_308,N_398);
or U474 (N_474,N_317,N_356);
nor U475 (N_475,N_359,N_367);
and U476 (N_476,N_344,N_378);
nand U477 (N_477,N_378,N_398);
xnor U478 (N_478,N_349,N_311);
or U479 (N_479,N_370,N_339);
nand U480 (N_480,N_354,N_394);
xor U481 (N_481,N_370,N_367);
or U482 (N_482,N_339,N_327);
or U483 (N_483,N_358,N_345);
nand U484 (N_484,N_311,N_368);
nand U485 (N_485,N_345,N_364);
xor U486 (N_486,N_322,N_359);
xnor U487 (N_487,N_383,N_348);
xor U488 (N_488,N_389,N_361);
nand U489 (N_489,N_317,N_328);
and U490 (N_490,N_381,N_331);
nand U491 (N_491,N_335,N_366);
nand U492 (N_492,N_341,N_379);
nand U493 (N_493,N_330,N_364);
and U494 (N_494,N_353,N_331);
and U495 (N_495,N_365,N_359);
or U496 (N_496,N_342,N_387);
xor U497 (N_497,N_362,N_323);
nand U498 (N_498,N_345,N_361);
xor U499 (N_499,N_385,N_339);
and U500 (N_500,N_443,N_458);
and U501 (N_501,N_431,N_407);
and U502 (N_502,N_499,N_481);
nand U503 (N_503,N_484,N_416);
or U504 (N_504,N_418,N_408);
nor U505 (N_505,N_467,N_457);
or U506 (N_506,N_483,N_441);
nand U507 (N_507,N_406,N_417);
nor U508 (N_508,N_438,N_450);
nand U509 (N_509,N_427,N_412);
nor U510 (N_510,N_428,N_455);
or U511 (N_511,N_469,N_452);
or U512 (N_512,N_449,N_444);
or U513 (N_513,N_492,N_451);
xnor U514 (N_514,N_471,N_479);
xor U515 (N_515,N_464,N_490);
or U516 (N_516,N_422,N_410);
and U517 (N_517,N_421,N_403);
xnor U518 (N_518,N_402,N_404);
nand U519 (N_519,N_419,N_468);
nor U520 (N_520,N_447,N_437);
or U521 (N_521,N_440,N_480);
xor U522 (N_522,N_489,N_497);
and U523 (N_523,N_439,N_475);
and U524 (N_524,N_436,N_462);
nand U525 (N_525,N_442,N_487);
and U526 (N_526,N_446,N_456);
xor U527 (N_527,N_477,N_461);
xor U528 (N_528,N_429,N_423);
nand U529 (N_529,N_434,N_494);
nand U530 (N_530,N_453,N_420);
or U531 (N_531,N_478,N_454);
or U532 (N_532,N_413,N_482);
nor U533 (N_533,N_465,N_460);
nand U534 (N_534,N_495,N_485);
nand U535 (N_535,N_470,N_445);
or U536 (N_536,N_424,N_498);
nor U537 (N_537,N_491,N_493);
or U538 (N_538,N_432,N_430);
and U539 (N_539,N_488,N_466);
nor U540 (N_540,N_459,N_463);
nand U541 (N_541,N_426,N_411);
nand U542 (N_542,N_472,N_433);
or U543 (N_543,N_425,N_474);
xor U544 (N_544,N_435,N_405);
xnor U545 (N_545,N_486,N_476);
nand U546 (N_546,N_401,N_448);
and U547 (N_547,N_409,N_414);
or U548 (N_548,N_496,N_400);
and U549 (N_549,N_415,N_473);
and U550 (N_550,N_472,N_499);
and U551 (N_551,N_450,N_429);
xor U552 (N_552,N_449,N_484);
nand U553 (N_553,N_463,N_404);
and U554 (N_554,N_486,N_416);
and U555 (N_555,N_470,N_486);
nand U556 (N_556,N_473,N_413);
nor U557 (N_557,N_478,N_468);
or U558 (N_558,N_456,N_415);
and U559 (N_559,N_420,N_466);
nor U560 (N_560,N_409,N_455);
xnor U561 (N_561,N_489,N_464);
or U562 (N_562,N_484,N_476);
xnor U563 (N_563,N_453,N_479);
xor U564 (N_564,N_441,N_408);
xor U565 (N_565,N_497,N_435);
and U566 (N_566,N_479,N_431);
nand U567 (N_567,N_448,N_418);
or U568 (N_568,N_418,N_447);
nor U569 (N_569,N_434,N_419);
xor U570 (N_570,N_414,N_468);
nor U571 (N_571,N_491,N_421);
and U572 (N_572,N_416,N_456);
and U573 (N_573,N_488,N_421);
nand U574 (N_574,N_458,N_497);
or U575 (N_575,N_424,N_446);
or U576 (N_576,N_498,N_472);
xnor U577 (N_577,N_425,N_463);
nor U578 (N_578,N_453,N_429);
or U579 (N_579,N_471,N_436);
or U580 (N_580,N_415,N_480);
and U581 (N_581,N_451,N_493);
xnor U582 (N_582,N_421,N_408);
nand U583 (N_583,N_498,N_444);
xor U584 (N_584,N_466,N_472);
xnor U585 (N_585,N_485,N_475);
or U586 (N_586,N_495,N_447);
xnor U587 (N_587,N_449,N_456);
or U588 (N_588,N_424,N_493);
and U589 (N_589,N_404,N_410);
and U590 (N_590,N_499,N_419);
nand U591 (N_591,N_490,N_491);
nor U592 (N_592,N_416,N_442);
and U593 (N_593,N_417,N_489);
and U594 (N_594,N_491,N_419);
xnor U595 (N_595,N_462,N_430);
nor U596 (N_596,N_469,N_432);
xor U597 (N_597,N_456,N_459);
nand U598 (N_598,N_496,N_452);
xor U599 (N_599,N_402,N_419);
or U600 (N_600,N_518,N_507);
nor U601 (N_601,N_595,N_590);
or U602 (N_602,N_549,N_597);
nor U603 (N_603,N_556,N_505);
nand U604 (N_604,N_523,N_516);
or U605 (N_605,N_574,N_593);
nor U606 (N_606,N_509,N_573);
and U607 (N_607,N_572,N_565);
xnor U608 (N_608,N_592,N_510);
or U609 (N_609,N_538,N_577);
and U610 (N_610,N_513,N_534);
xnor U611 (N_611,N_563,N_506);
nor U612 (N_612,N_599,N_596);
or U613 (N_613,N_508,N_528);
or U614 (N_614,N_570,N_526);
xnor U615 (N_615,N_554,N_552);
xor U616 (N_616,N_575,N_529);
xor U617 (N_617,N_560,N_582);
nor U618 (N_618,N_502,N_540);
xnor U619 (N_619,N_581,N_594);
or U620 (N_620,N_588,N_525);
nand U621 (N_621,N_561,N_569);
and U622 (N_622,N_559,N_520);
nand U623 (N_623,N_591,N_521);
nor U624 (N_624,N_579,N_546);
nor U625 (N_625,N_585,N_576);
nand U626 (N_626,N_543,N_503);
xor U627 (N_627,N_571,N_598);
nand U628 (N_628,N_515,N_524);
nor U629 (N_629,N_553,N_533);
or U630 (N_630,N_541,N_547);
and U631 (N_631,N_500,N_539);
nand U632 (N_632,N_544,N_578);
xor U633 (N_633,N_562,N_545);
and U634 (N_634,N_512,N_551);
xor U635 (N_635,N_511,N_504);
xnor U636 (N_636,N_517,N_589);
and U637 (N_637,N_550,N_536);
xnor U638 (N_638,N_557,N_566);
and U639 (N_639,N_537,N_586);
nand U640 (N_640,N_584,N_568);
nand U641 (N_641,N_583,N_514);
xnor U642 (N_642,N_535,N_501);
or U643 (N_643,N_522,N_587);
or U644 (N_644,N_542,N_531);
and U645 (N_645,N_564,N_527);
or U646 (N_646,N_580,N_555);
nor U647 (N_647,N_530,N_567);
xnor U648 (N_648,N_532,N_558);
nand U649 (N_649,N_519,N_548);
and U650 (N_650,N_579,N_501);
and U651 (N_651,N_501,N_572);
nor U652 (N_652,N_533,N_547);
nor U653 (N_653,N_513,N_535);
xnor U654 (N_654,N_573,N_520);
nor U655 (N_655,N_583,N_599);
nor U656 (N_656,N_562,N_569);
nor U657 (N_657,N_570,N_548);
xor U658 (N_658,N_591,N_541);
xor U659 (N_659,N_584,N_575);
nand U660 (N_660,N_501,N_551);
and U661 (N_661,N_535,N_534);
and U662 (N_662,N_570,N_595);
xnor U663 (N_663,N_581,N_558);
nand U664 (N_664,N_524,N_555);
and U665 (N_665,N_551,N_549);
and U666 (N_666,N_581,N_572);
nand U667 (N_667,N_585,N_581);
xnor U668 (N_668,N_539,N_504);
or U669 (N_669,N_564,N_556);
and U670 (N_670,N_594,N_564);
and U671 (N_671,N_566,N_552);
xor U672 (N_672,N_580,N_567);
nand U673 (N_673,N_597,N_538);
nor U674 (N_674,N_596,N_595);
nor U675 (N_675,N_585,N_579);
xnor U676 (N_676,N_563,N_556);
and U677 (N_677,N_589,N_504);
nand U678 (N_678,N_537,N_561);
xor U679 (N_679,N_570,N_533);
and U680 (N_680,N_588,N_576);
or U681 (N_681,N_572,N_512);
nand U682 (N_682,N_529,N_560);
or U683 (N_683,N_583,N_586);
nor U684 (N_684,N_520,N_574);
or U685 (N_685,N_552,N_519);
xnor U686 (N_686,N_512,N_527);
or U687 (N_687,N_594,N_598);
and U688 (N_688,N_553,N_525);
xor U689 (N_689,N_539,N_587);
nand U690 (N_690,N_576,N_551);
or U691 (N_691,N_556,N_555);
or U692 (N_692,N_587,N_544);
nand U693 (N_693,N_517,N_524);
xnor U694 (N_694,N_539,N_564);
nor U695 (N_695,N_588,N_531);
or U696 (N_696,N_506,N_558);
nand U697 (N_697,N_574,N_566);
and U698 (N_698,N_501,N_521);
nor U699 (N_699,N_517,N_510);
nor U700 (N_700,N_641,N_618);
or U701 (N_701,N_679,N_695);
nor U702 (N_702,N_616,N_648);
nand U703 (N_703,N_667,N_622);
nor U704 (N_704,N_659,N_694);
xnor U705 (N_705,N_675,N_661);
nor U706 (N_706,N_631,N_685);
and U707 (N_707,N_691,N_642);
xor U708 (N_708,N_672,N_693);
nor U709 (N_709,N_686,N_624);
and U710 (N_710,N_643,N_684);
nor U711 (N_711,N_670,N_692);
xor U712 (N_712,N_646,N_668);
and U713 (N_713,N_683,N_634);
nand U714 (N_714,N_656,N_620);
and U715 (N_715,N_637,N_651);
or U716 (N_716,N_665,N_664);
nand U717 (N_717,N_608,N_617);
xnor U718 (N_718,N_638,N_688);
nand U719 (N_719,N_611,N_629);
xor U720 (N_720,N_639,N_699);
nand U721 (N_721,N_663,N_644);
nor U722 (N_722,N_690,N_615);
or U723 (N_723,N_653,N_625);
nor U724 (N_724,N_601,N_673);
xnor U725 (N_725,N_689,N_635);
or U726 (N_726,N_650,N_636);
nor U727 (N_727,N_671,N_662);
or U728 (N_728,N_605,N_619);
nor U729 (N_729,N_640,N_697);
and U730 (N_730,N_654,N_678);
nor U731 (N_731,N_682,N_655);
nor U732 (N_732,N_657,N_687);
xor U733 (N_733,N_649,N_676);
xnor U734 (N_734,N_647,N_645);
nor U735 (N_735,N_604,N_652);
or U736 (N_736,N_600,N_626);
nor U737 (N_737,N_609,N_606);
or U738 (N_738,N_627,N_632);
and U739 (N_739,N_660,N_612);
or U740 (N_740,N_698,N_680);
nor U741 (N_741,N_633,N_674);
nor U742 (N_742,N_610,N_614);
nand U743 (N_743,N_681,N_630);
and U744 (N_744,N_658,N_696);
nor U745 (N_745,N_677,N_623);
and U746 (N_746,N_628,N_669);
xnor U747 (N_747,N_613,N_621);
or U748 (N_748,N_602,N_666);
nor U749 (N_749,N_603,N_607);
nand U750 (N_750,N_686,N_622);
xnor U751 (N_751,N_683,N_663);
nor U752 (N_752,N_686,N_690);
xnor U753 (N_753,N_612,N_667);
nand U754 (N_754,N_661,N_631);
nor U755 (N_755,N_694,N_650);
xnor U756 (N_756,N_668,N_647);
nand U757 (N_757,N_655,N_612);
and U758 (N_758,N_615,N_624);
xor U759 (N_759,N_643,N_671);
nor U760 (N_760,N_663,N_678);
nor U761 (N_761,N_612,N_666);
nor U762 (N_762,N_615,N_619);
xnor U763 (N_763,N_684,N_644);
nand U764 (N_764,N_611,N_676);
nor U765 (N_765,N_644,N_612);
nand U766 (N_766,N_689,N_622);
xor U767 (N_767,N_692,N_634);
nor U768 (N_768,N_687,N_619);
nand U769 (N_769,N_608,N_671);
or U770 (N_770,N_655,N_644);
nand U771 (N_771,N_628,N_688);
nand U772 (N_772,N_691,N_685);
nand U773 (N_773,N_623,N_695);
or U774 (N_774,N_681,N_679);
or U775 (N_775,N_645,N_602);
nand U776 (N_776,N_676,N_682);
nand U777 (N_777,N_627,N_609);
or U778 (N_778,N_627,N_637);
and U779 (N_779,N_609,N_684);
xnor U780 (N_780,N_699,N_618);
and U781 (N_781,N_666,N_689);
and U782 (N_782,N_640,N_699);
and U783 (N_783,N_678,N_670);
or U784 (N_784,N_676,N_610);
and U785 (N_785,N_619,N_608);
xnor U786 (N_786,N_642,N_619);
or U787 (N_787,N_624,N_676);
nand U788 (N_788,N_646,N_621);
xnor U789 (N_789,N_610,N_617);
xnor U790 (N_790,N_648,N_632);
and U791 (N_791,N_697,N_679);
xor U792 (N_792,N_636,N_631);
xor U793 (N_793,N_682,N_646);
nor U794 (N_794,N_677,N_603);
and U795 (N_795,N_677,N_602);
nor U796 (N_796,N_695,N_609);
nand U797 (N_797,N_633,N_699);
xnor U798 (N_798,N_610,N_615);
nand U799 (N_799,N_631,N_675);
nor U800 (N_800,N_704,N_786);
nor U801 (N_801,N_708,N_778);
and U802 (N_802,N_772,N_753);
xnor U803 (N_803,N_707,N_732);
and U804 (N_804,N_751,N_792);
or U805 (N_805,N_701,N_748);
and U806 (N_806,N_794,N_713);
or U807 (N_807,N_767,N_779);
nand U808 (N_808,N_775,N_745);
or U809 (N_809,N_782,N_752);
nand U810 (N_810,N_718,N_796);
or U811 (N_811,N_787,N_731);
or U812 (N_812,N_784,N_720);
nand U813 (N_813,N_733,N_738);
or U814 (N_814,N_770,N_724);
xor U815 (N_815,N_771,N_714);
nor U816 (N_816,N_760,N_765);
and U817 (N_817,N_777,N_766);
or U818 (N_818,N_776,N_715);
nor U819 (N_819,N_774,N_737);
nor U820 (N_820,N_783,N_739);
or U821 (N_821,N_759,N_710);
nand U822 (N_822,N_726,N_756);
nand U823 (N_823,N_735,N_788);
and U824 (N_824,N_761,N_736);
or U825 (N_825,N_702,N_746);
nand U826 (N_826,N_795,N_762);
and U827 (N_827,N_790,N_727);
nand U828 (N_828,N_769,N_755);
nor U829 (N_829,N_763,N_744);
nand U830 (N_830,N_729,N_734);
or U831 (N_831,N_722,N_728);
and U832 (N_832,N_781,N_716);
xnor U833 (N_833,N_742,N_711);
nor U834 (N_834,N_703,N_798);
or U835 (N_835,N_709,N_749);
nor U836 (N_836,N_785,N_780);
xor U837 (N_837,N_754,N_725);
or U838 (N_838,N_719,N_797);
and U839 (N_839,N_706,N_750);
and U840 (N_840,N_721,N_712);
xor U841 (N_841,N_730,N_700);
nor U842 (N_842,N_705,N_757);
nor U843 (N_843,N_741,N_789);
and U844 (N_844,N_791,N_717);
nand U845 (N_845,N_758,N_799);
xor U846 (N_846,N_747,N_743);
and U847 (N_847,N_723,N_773);
and U848 (N_848,N_764,N_793);
or U849 (N_849,N_740,N_768);
nor U850 (N_850,N_727,N_789);
or U851 (N_851,N_737,N_729);
and U852 (N_852,N_786,N_755);
or U853 (N_853,N_705,N_762);
nand U854 (N_854,N_722,N_711);
or U855 (N_855,N_795,N_728);
or U856 (N_856,N_706,N_772);
and U857 (N_857,N_776,N_771);
xnor U858 (N_858,N_784,N_799);
and U859 (N_859,N_704,N_767);
nand U860 (N_860,N_782,N_742);
xnor U861 (N_861,N_795,N_785);
nor U862 (N_862,N_719,N_757);
and U863 (N_863,N_709,N_702);
nand U864 (N_864,N_762,N_707);
nor U865 (N_865,N_722,N_778);
nor U866 (N_866,N_753,N_754);
nand U867 (N_867,N_735,N_737);
xor U868 (N_868,N_734,N_778);
nand U869 (N_869,N_734,N_775);
nand U870 (N_870,N_753,N_703);
nand U871 (N_871,N_751,N_724);
or U872 (N_872,N_759,N_767);
nand U873 (N_873,N_797,N_760);
nand U874 (N_874,N_785,N_763);
and U875 (N_875,N_789,N_709);
and U876 (N_876,N_703,N_759);
and U877 (N_877,N_747,N_741);
xnor U878 (N_878,N_797,N_795);
or U879 (N_879,N_754,N_751);
xor U880 (N_880,N_782,N_709);
xnor U881 (N_881,N_748,N_760);
nor U882 (N_882,N_736,N_735);
xor U883 (N_883,N_715,N_765);
nand U884 (N_884,N_704,N_760);
and U885 (N_885,N_769,N_745);
and U886 (N_886,N_766,N_726);
or U887 (N_887,N_776,N_753);
or U888 (N_888,N_799,N_786);
and U889 (N_889,N_719,N_764);
xor U890 (N_890,N_761,N_740);
nor U891 (N_891,N_778,N_703);
nand U892 (N_892,N_705,N_728);
and U893 (N_893,N_728,N_771);
or U894 (N_894,N_752,N_718);
nor U895 (N_895,N_737,N_734);
nand U896 (N_896,N_774,N_707);
and U897 (N_897,N_788,N_768);
nor U898 (N_898,N_726,N_744);
nor U899 (N_899,N_738,N_799);
and U900 (N_900,N_836,N_810);
nor U901 (N_901,N_868,N_817);
and U902 (N_902,N_846,N_897);
xor U903 (N_903,N_893,N_872);
or U904 (N_904,N_889,N_804);
nand U905 (N_905,N_860,N_814);
nor U906 (N_906,N_813,N_838);
nor U907 (N_907,N_892,N_848);
nand U908 (N_908,N_826,N_878);
or U909 (N_909,N_876,N_847);
xnor U910 (N_910,N_886,N_831);
or U911 (N_911,N_870,N_822);
nor U912 (N_912,N_856,N_873);
nand U913 (N_913,N_806,N_891);
nor U914 (N_914,N_815,N_898);
nand U915 (N_915,N_839,N_803);
and U916 (N_916,N_830,N_842);
nand U917 (N_917,N_874,N_829);
nand U918 (N_918,N_855,N_851);
nand U919 (N_919,N_835,N_864);
nor U920 (N_920,N_899,N_884);
nand U921 (N_921,N_877,N_800);
and U922 (N_922,N_869,N_820);
nor U923 (N_923,N_849,N_885);
nor U924 (N_924,N_834,N_894);
xnor U925 (N_925,N_823,N_871);
nand U926 (N_926,N_812,N_828);
and U927 (N_927,N_883,N_845);
nand U928 (N_928,N_890,N_808);
and U929 (N_929,N_887,N_867);
nor U930 (N_930,N_895,N_840);
nor U931 (N_931,N_816,N_854);
nor U932 (N_932,N_888,N_841);
or U933 (N_933,N_821,N_850);
nand U934 (N_934,N_832,N_866);
and U935 (N_935,N_809,N_827);
or U936 (N_936,N_852,N_862);
and U937 (N_937,N_875,N_853);
nor U938 (N_938,N_818,N_805);
and U939 (N_939,N_819,N_858);
nand U940 (N_940,N_861,N_825);
nand U941 (N_941,N_880,N_896);
and U942 (N_942,N_879,N_837);
or U943 (N_943,N_844,N_811);
and U944 (N_944,N_857,N_881);
or U945 (N_945,N_807,N_802);
nand U946 (N_946,N_843,N_865);
or U947 (N_947,N_859,N_801);
and U948 (N_948,N_824,N_882);
nor U949 (N_949,N_863,N_833);
nand U950 (N_950,N_891,N_818);
or U951 (N_951,N_855,N_854);
or U952 (N_952,N_886,N_888);
nor U953 (N_953,N_810,N_816);
nand U954 (N_954,N_807,N_880);
or U955 (N_955,N_849,N_899);
or U956 (N_956,N_871,N_852);
nor U957 (N_957,N_842,N_880);
nand U958 (N_958,N_865,N_814);
xnor U959 (N_959,N_823,N_805);
and U960 (N_960,N_836,N_870);
nand U961 (N_961,N_869,N_857);
xor U962 (N_962,N_861,N_820);
nand U963 (N_963,N_864,N_899);
nor U964 (N_964,N_864,N_813);
nor U965 (N_965,N_810,N_807);
or U966 (N_966,N_884,N_863);
and U967 (N_967,N_817,N_844);
xor U968 (N_968,N_819,N_872);
or U969 (N_969,N_803,N_870);
xnor U970 (N_970,N_853,N_851);
nor U971 (N_971,N_893,N_847);
nand U972 (N_972,N_860,N_852);
nor U973 (N_973,N_850,N_830);
and U974 (N_974,N_832,N_899);
nand U975 (N_975,N_851,N_802);
and U976 (N_976,N_841,N_820);
nand U977 (N_977,N_877,N_868);
nor U978 (N_978,N_899,N_860);
xnor U979 (N_979,N_891,N_808);
nand U980 (N_980,N_893,N_899);
nand U981 (N_981,N_827,N_807);
xor U982 (N_982,N_810,N_898);
nand U983 (N_983,N_893,N_862);
xnor U984 (N_984,N_823,N_846);
nand U985 (N_985,N_878,N_815);
or U986 (N_986,N_833,N_868);
or U987 (N_987,N_817,N_864);
nor U988 (N_988,N_819,N_862);
or U989 (N_989,N_838,N_854);
nand U990 (N_990,N_824,N_810);
nor U991 (N_991,N_848,N_865);
or U992 (N_992,N_885,N_882);
nor U993 (N_993,N_823,N_847);
and U994 (N_994,N_836,N_843);
xnor U995 (N_995,N_812,N_863);
nor U996 (N_996,N_890,N_803);
xor U997 (N_997,N_896,N_832);
nor U998 (N_998,N_890,N_834);
and U999 (N_999,N_819,N_877);
or U1000 (N_1000,N_969,N_953);
nand U1001 (N_1001,N_911,N_941);
or U1002 (N_1002,N_934,N_976);
nand U1003 (N_1003,N_931,N_928);
nand U1004 (N_1004,N_906,N_973);
nor U1005 (N_1005,N_919,N_990);
and U1006 (N_1006,N_966,N_908);
xnor U1007 (N_1007,N_910,N_992);
nand U1008 (N_1008,N_999,N_943);
or U1009 (N_1009,N_907,N_950);
or U1010 (N_1010,N_937,N_935);
and U1011 (N_1011,N_972,N_940);
or U1012 (N_1012,N_900,N_955);
nor U1013 (N_1013,N_995,N_989);
xor U1014 (N_1014,N_970,N_982);
xnor U1015 (N_1015,N_916,N_985);
nand U1016 (N_1016,N_909,N_915);
and U1017 (N_1017,N_929,N_933);
or U1018 (N_1018,N_980,N_913);
or U1019 (N_1019,N_939,N_946);
xor U1020 (N_1020,N_926,N_904);
nor U1021 (N_1021,N_967,N_945);
and U1022 (N_1022,N_922,N_984);
and U1023 (N_1023,N_961,N_951);
and U1024 (N_1024,N_905,N_925);
and U1025 (N_1025,N_998,N_981);
and U1026 (N_1026,N_986,N_936);
nor U1027 (N_1027,N_977,N_949);
nor U1028 (N_1028,N_962,N_921);
xnor U1029 (N_1029,N_914,N_930);
or U1030 (N_1030,N_952,N_924);
nand U1031 (N_1031,N_959,N_996);
xnor U1032 (N_1032,N_938,N_957);
nor U1033 (N_1033,N_912,N_956);
and U1034 (N_1034,N_901,N_954);
and U1035 (N_1035,N_960,N_987);
nand U1036 (N_1036,N_979,N_971);
nand U1037 (N_1037,N_920,N_964);
nor U1038 (N_1038,N_963,N_997);
nand U1039 (N_1039,N_923,N_927);
xnor U1040 (N_1040,N_942,N_917);
or U1041 (N_1041,N_918,N_965);
nor U1042 (N_1042,N_994,N_975);
nand U1043 (N_1043,N_944,N_947);
or U1044 (N_1044,N_974,N_958);
nand U1045 (N_1045,N_978,N_932);
or U1046 (N_1046,N_903,N_988);
nor U1047 (N_1047,N_993,N_968);
xnor U1048 (N_1048,N_991,N_948);
nand U1049 (N_1049,N_983,N_902);
and U1050 (N_1050,N_936,N_915);
or U1051 (N_1051,N_994,N_990);
and U1052 (N_1052,N_948,N_981);
nand U1053 (N_1053,N_992,N_907);
nand U1054 (N_1054,N_967,N_906);
and U1055 (N_1055,N_916,N_920);
nand U1056 (N_1056,N_905,N_901);
nor U1057 (N_1057,N_919,N_989);
xor U1058 (N_1058,N_979,N_973);
nand U1059 (N_1059,N_923,N_919);
and U1060 (N_1060,N_927,N_918);
nor U1061 (N_1061,N_985,N_989);
nand U1062 (N_1062,N_970,N_912);
nor U1063 (N_1063,N_962,N_918);
xor U1064 (N_1064,N_986,N_938);
and U1065 (N_1065,N_969,N_921);
or U1066 (N_1066,N_910,N_955);
xnor U1067 (N_1067,N_989,N_925);
nor U1068 (N_1068,N_932,N_979);
nand U1069 (N_1069,N_932,N_965);
and U1070 (N_1070,N_918,N_929);
or U1071 (N_1071,N_979,N_996);
xor U1072 (N_1072,N_964,N_905);
nor U1073 (N_1073,N_920,N_970);
xnor U1074 (N_1074,N_983,N_958);
nand U1075 (N_1075,N_903,N_901);
or U1076 (N_1076,N_911,N_953);
nand U1077 (N_1077,N_919,N_946);
xor U1078 (N_1078,N_950,N_995);
nand U1079 (N_1079,N_977,N_920);
xor U1080 (N_1080,N_904,N_940);
or U1081 (N_1081,N_976,N_926);
and U1082 (N_1082,N_956,N_993);
or U1083 (N_1083,N_906,N_932);
or U1084 (N_1084,N_962,N_983);
nand U1085 (N_1085,N_978,N_901);
nand U1086 (N_1086,N_963,N_913);
nor U1087 (N_1087,N_907,N_919);
xor U1088 (N_1088,N_930,N_981);
nor U1089 (N_1089,N_943,N_924);
xor U1090 (N_1090,N_925,N_929);
or U1091 (N_1091,N_909,N_904);
xor U1092 (N_1092,N_957,N_916);
nand U1093 (N_1093,N_999,N_979);
xor U1094 (N_1094,N_975,N_934);
or U1095 (N_1095,N_989,N_944);
or U1096 (N_1096,N_911,N_943);
xor U1097 (N_1097,N_982,N_943);
nor U1098 (N_1098,N_956,N_940);
nor U1099 (N_1099,N_943,N_989);
nor U1100 (N_1100,N_1036,N_1018);
xnor U1101 (N_1101,N_1047,N_1070);
and U1102 (N_1102,N_1020,N_1056);
and U1103 (N_1103,N_1086,N_1025);
nor U1104 (N_1104,N_1066,N_1048);
nand U1105 (N_1105,N_1096,N_1017);
xnor U1106 (N_1106,N_1095,N_1080);
or U1107 (N_1107,N_1082,N_1008);
xor U1108 (N_1108,N_1021,N_1050);
nor U1109 (N_1109,N_1073,N_1064);
nand U1110 (N_1110,N_1092,N_1007);
or U1111 (N_1111,N_1031,N_1067);
nor U1112 (N_1112,N_1079,N_1012);
nor U1113 (N_1113,N_1040,N_1049);
or U1114 (N_1114,N_1022,N_1076);
and U1115 (N_1115,N_1065,N_1001);
xnor U1116 (N_1116,N_1089,N_1085);
nor U1117 (N_1117,N_1088,N_1027);
nand U1118 (N_1118,N_1039,N_1029);
xnor U1119 (N_1119,N_1074,N_1071);
nand U1120 (N_1120,N_1010,N_1051);
and U1121 (N_1121,N_1077,N_1006);
and U1122 (N_1122,N_1093,N_1043);
or U1123 (N_1123,N_1084,N_1094);
xnor U1124 (N_1124,N_1037,N_1055);
or U1125 (N_1125,N_1013,N_1097);
and U1126 (N_1126,N_1063,N_1091);
and U1127 (N_1127,N_1099,N_1054);
nor U1128 (N_1128,N_1032,N_1053);
xor U1129 (N_1129,N_1016,N_1005);
xor U1130 (N_1130,N_1046,N_1026);
or U1131 (N_1131,N_1098,N_1028);
xor U1132 (N_1132,N_1004,N_1038);
and U1133 (N_1133,N_1041,N_1003);
xor U1134 (N_1134,N_1014,N_1059);
and U1135 (N_1135,N_1015,N_1000);
or U1136 (N_1136,N_1078,N_1062);
nand U1137 (N_1137,N_1011,N_1087);
nand U1138 (N_1138,N_1072,N_1068);
nand U1139 (N_1139,N_1058,N_1023);
and U1140 (N_1140,N_1002,N_1057);
nand U1141 (N_1141,N_1034,N_1033);
xnor U1142 (N_1142,N_1035,N_1081);
or U1143 (N_1143,N_1009,N_1024);
nand U1144 (N_1144,N_1030,N_1060);
and U1145 (N_1145,N_1061,N_1075);
xnor U1146 (N_1146,N_1083,N_1069);
and U1147 (N_1147,N_1045,N_1052);
and U1148 (N_1148,N_1019,N_1090);
nor U1149 (N_1149,N_1044,N_1042);
and U1150 (N_1150,N_1043,N_1031);
xnor U1151 (N_1151,N_1022,N_1078);
and U1152 (N_1152,N_1017,N_1060);
nor U1153 (N_1153,N_1093,N_1032);
nand U1154 (N_1154,N_1075,N_1078);
xor U1155 (N_1155,N_1024,N_1064);
nand U1156 (N_1156,N_1079,N_1011);
xor U1157 (N_1157,N_1075,N_1019);
or U1158 (N_1158,N_1094,N_1019);
nand U1159 (N_1159,N_1020,N_1061);
nor U1160 (N_1160,N_1084,N_1018);
nor U1161 (N_1161,N_1028,N_1047);
nand U1162 (N_1162,N_1014,N_1012);
nand U1163 (N_1163,N_1061,N_1004);
nor U1164 (N_1164,N_1058,N_1033);
or U1165 (N_1165,N_1017,N_1037);
nor U1166 (N_1166,N_1084,N_1088);
nor U1167 (N_1167,N_1098,N_1087);
and U1168 (N_1168,N_1075,N_1090);
or U1169 (N_1169,N_1094,N_1009);
nor U1170 (N_1170,N_1031,N_1056);
and U1171 (N_1171,N_1095,N_1068);
nand U1172 (N_1172,N_1049,N_1071);
nor U1173 (N_1173,N_1057,N_1084);
or U1174 (N_1174,N_1054,N_1019);
or U1175 (N_1175,N_1064,N_1019);
xor U1176 (N_1176,N_1063,N_1023);
xor U1177 (N_1177,N_1070,N_1061);
xor U1178 (N_1178,N_1092,N_1074);
nand U1179 (N_1179,N_1031,N_1091);
or U1180 (N_1180,N_1038,N_1052);
or U1181 (N_1181,N_1086,N_1020);
xnor U1182 (N_1182,N_1009,N_1008);
and U1183 (N_1183,N_1095,N_1091);
nand U1184 (N_1184,N_1051,N_1020);
and U1185 (N_1185,N_1080,N_1074);
nor U1186 (N_1186,N_1050,N_1020);
and U1187 (N_1187,N_1057,N_1050);
xnor U1188 (N_1188,N_1066,N_1077);
xnor U1189 (N_1189,N_1007,N_1083);
xnor U1190 (N_1190,N_1026,N_1022);
and U1191 (N_1191,N_1065,N_1016);
nor U1192 (N_1192,N_1045,N_1011);
xnor U1193 (N_1193,N_1081,N_1080);
or U1194 (N_1194,N_1036,N_1029);
nand U1195 (N_1195,N_1030,N_1004);
nand U1196 (N_1196,N_1037,N_1048);
or U1197 (N_1197,N_1078,N_1010);
nor U1198 (N_1198,N_1078,N_1038);
and U1199 (N_1199,N_1031,N_1062);
xor U1200 (N_1200,N_1184,N_1191);
and U1201 (N_1201,N_1128,N_1105);
nor U1202 (N_1202,N_1193,N_1142);
nor U1203 (N_1203,N_1131,N_1194);
or U1204 (N_1204,N_1107,N_1181);
nand U1205 (N_1205,N_1122,N_1189);
and U1206 (N_1206,N_1129,N_1182);
nand U1207 (N_1207,N_1103,N_1124);
and U1208 (N_1208,N_1106,N_1173);
nand U1209 (N_1209,N_1121,N_1153);
nand U1210 (N_1210,N_1170,N_1137);
nor U1211 (N_1211,N_1147,N_1136);
nor U1212 (N_1212,N_1143,N_1187);
or U1213 (N_1213,N_1169,N_1178);
or U1214 (N_1214,N_1175,N_1157);
or U1215 (N_1215,N_1167,N_1104);
and U1216 (N_1216,N_1149,N_1113);
or U1217 (N_1217,N_1134,N_1130);
and U1218 (N_1218,N_1119,N_1120);
and U1219 (N_1219,N_1159,N_1125);
nor U1220 (N_1220,N_1146,N_1126);
and U1221 (N_1221,N_1199,N_1108);
nand U1222 (N_1222,N_1172,N_1158);
nor U1223 (N_1223,N_1185,N_1198);
xor U1224 (N_1224,N_1141,N_1196);
or U1225 (N_1225,N_1133,N_1112);
and U1226 (N_1226,N_1117,N_1100);
or U1227 (N_1227,N_1180,N_1151);
xnor U1228 (N_1228,N_1171,N_1188);
xor U1229 (N_1229,N_1114,N_1197);
nand U1230 (N_1230,N_1168,N_1186);
xor U1231 (N_1231,N_1195,N_1154);
or U1232 (N_1232,N_1155,N_1140);
or U1233 (N_1233,N_1177,N_1162);
xor U1234 (N_1234,N_1179,N_1138);
nor U1235 (N_1235,N_1161,N_1152);
and U1236 (N_1236,N_1165,N_1109);
or U1237 (N_1237,N_1192,N_1115);
nand U1238 (N_1238,N_1163,N_1102);
nor U1239 (N_1239,N_1148,N_1144);
xnor U1240 (N_1240,N_1111,N_1176);
xor U1241 (N_1241,N_1183,N_1101);
nand U1242 (N_1242,N_1174,N_1116);
and U1243 (N_1243,N_1164,N_1150);
nand U1244 (N_1244,N_1135,N_1166);
nor U1245 (N_1245,N_1145,N_1118);
xnor U1246 (N_1246,N_1123,N_1190);
xnor U1247 (N_1247,N_1127,N_1110);
and U1248 (N_1248,N_1156,N_1132);
nor U1249 (N_1249,N_1139,N_1160);
nand U1250 (N_1250,N_1187,N_1134);
xor U1251 (N_1251,N_1104,N_1160);
or U1252 (N_1252,N_1107,N_1136);
nand U1253 (N_1253,N_1146,N_1186);
xor U1254 (N_1254,N_1141,N_1156);
nand U1255 (N_1255,N_1166,N_1153);
nor U1256 (N_1256,N_1179,N_1137);
and U1257 (N_1257,N_1120,N_1115);
or U1258 (N_1258,N_1120,N_1123);
and U1259 (N_1259,N_1166,N_1177);
and U1260 (N_1260,N_1145,N_1153);
or U1261 (N_1261,N_1122,N_1117);
and U1262 (N_1262,N_1154,N_1156);
or U1263 (N_1263,N_1181,N_1155);
and U1264 (N_1264,N_1126,N_1129);
nor U1265 (N_1265,N_1157,N_1177);
nand U1266 (N_1266,N_1164,N_1107);
and U1267 (N_1267,N_1178,N_1191);
xor U1268 (N_1268,N_1189,N_1138);
or U1269 (N_1269,N_1116,N_1171);
or U1270 (N_1270,N_1140,N_1156);
nor U1271 (N_1271,N_1121,N_1163);
nor U1272 (N_1272,N_1189,N_1165);
xnor U1273 (N_1273,N_1131,N_1178);
nor U1274 (N_1274,N_1155,N_1118);
xnor U1275 (N_1275,N_1188,N_1154);
and U1276 (N_1276,N_1100,N_1185);
and U1277 (N_1277,N_1179,N_1142);
xnor U1278 (N_1278,N_1190,N_1176);
and U1279 (N_1279,N_1161,N_1194);
or U1280 (N_1280,N_1196,N_1113);
nor U1281 (N_1281,N_1173,N_1127);
or U1282 (N_1282,N_1109,N_1151);
xor U1283 (N_1283,N_1101,N_1191);
and U1284 (N_1284,N_1190,N_1198);
xor U1285 (N_1285,N_1154,N_1120);
nor U1286 (N_1286,N_1163,N_1160);
or U1287 (N_1287,N_1134,N_1135);
nand U1288 (N_1288,N_1161,N_1158);
xor U1289 (N_1289,N_1183,N_1137);
nor U1290 (N_1290,N_1119,N_1173);
nand U1291 (N_1291,N_1149,N_1114);
and U1292 (N_1292,N_1172,N_1160);
or U1293 (N_1293,N_1113,N_1173);
xnor U1294 (N_1294,N_1145,N_1132);
xor U1295 (N_1295,N_1188,N_1141);
or U1296 (N_1296,N_1120,N_1138);
nor U1297 (N_1297,N_1188,N_1126);
nand U1298 (N_1298,N_1154,N_1198);
nand U1299 (N_1299,N_1140,N_1160);
or U1300 (N_1300,N_1219,N_1210);
xnor U1301 (N_1301,N_1201,N_1221);
nand U1302 (N_1302,N_1262,N_1297);
or U1303 (N_1303,N_1274,N_1273);
nor U1304 (N_1304,N_1278,N_1254);
and U1305 (N_1305,N_1264,N_1205);
or U1306 (N_1306,N_1250,N_1224);
or U1307 (N_1307,N_1291,N_1207);
or U1308 (N_1308,N_1293,N_1267);
or U1309 (N_1309,N_1257,N_1232);
or U1310 (N_1310,N_1204,N_1225);
nor U1311 (N_1311,N_1288,N_1220);
or U1312 (N_1312,N_1258,N_1261);
and U1313 (N_1313,N_1282,N_1271);
or U1314 (N_1314,N_1223,N_1206);
xnor U1315 (N_1315,N_1246,N_1238);
or U1316 (N_1316,N_1241,N_1272);
nor U1317 (N_1317,N_1268,N_1215);
nor U1318 (N_1318,N_1255,N_1251);
nand U1319 (N_1319,N_1239,N_1285);
xor U1320 (N_1320,N_1235,N_1253);
xor U1321 (N_1321,N_1234,N_1259);
nor U1322 (N_1322,N_1217,N_1281);
nor U1323 (N_1323,N_1203,N_1260);
and U1324 (N_1324,N_1214,N_1296);
or U1325 (N_1325,N_1295,N_1263);
or U1326 (N_1326,N_1245,N_1228);
nor U1327 (N_1327,N_1283,N_1244);
nor U1328 (N_1328,N_1212,N_1277);
and U1329 (N_1329,N_1209,N_1226);
or U1330 (N_1330,N_1287,N_1249);
nand U1331 (N_1331,N_1292,N_1275);
nor U1332 (N_1332,N_1213,N_1240);
nor U1333 (N_1333,N_1243,N_1279);
or U1334 (N_1334,N_1227,N_1231);
or U1335 (N_1335,N_1256,N_1294);
xor U1336 (N_1336,N_1298,N_1270);
or U1337 (N_1337,N_1284,N_1247);
or U1338 (N_1338,N_1202,N_1248);
and U1339 (N_1339,N_1237,N_1286);
xnor U1340 (N_1340,N_1252,N_1242);
nor U1341 (N_1341,N_1216,N_1269);
or U1342 (N_1342,N_1229,N_1290);
or U1343 (N_1343,N_1265,N_1280);
nand U1344 (N_1344,N_1208,N_1299);
and U1345 (N_1345,N_1200,N_1276);
nand U1346 (N_1346,N_1230,N_1233);
xor U1347 (N_1347,N_1289,N_1266);
and U1348 (N_1348,N_1222,N_1211);
xnor U1349 (N_1349,N_1236,N_1218);
nand U1350 (N_1350,N_1269,N_1281);
xnor U1351 (N_1351,N_1256,N_1218);
nor U1352 (N_1352,N_1221,N_1204);
nor U1353 (N_1353,N_1240,N_1284);
xor U1354 (N_1354,N_1236,N_1288);
or U1355 (N_1355,N_1291,N_1280);
xor U1356 (N_1356,N_1205,N_1212);
nand U1357 (N_1357,N_1289,N_1219);
nor U1358 (N_1358,N_1226,N_1275);
or U1359 (N_1359,N_1224,N_1270);
xor U1360 (N_1360,N_1204,N_1202);
xnor U1361 (N_1361,N_1235,N_1291);
and U1362 (N_1362,N_1229,N_1232);
xnor U1363 (N_1363,N_1249,N_1213);
and U1364 (N_1364,N_1272,N_1207);
xnor U1365 (N_1365,N_1253,N_1285);
nor U1366 (N_1366,N_1231,N_1268);
xnor U1367 (N_1367,N_1258,N_1206);
nor U1368 (N_1368,N_1202,N_1262);
or U1369 (N_1369,N_1276,N_1208);
or U1370 (N_1370,N_1210,N_1255);
and U1371 (N_1371,N_1295,N_1254);
nand U1372 (N_1372,N_1207,N_1287);
xor U1373 (N_1373,N_1239,N_1248);
nor U1374 (N_1374,N_1293,N_1296);
nand U1375 (N_1375,N_1266,N_1287);
or U1376 (N_1376,N_1269,N_1233);
nand U1377 (N_1377,N_1245,N_1255);
and U1378 (N_1378,N_1298,N_1206);
xnor U1379 (N_1379,N_1275,N_1248);
and U1380 (N_1380,N_1254,N_1251);
xor U1381 (N_1381,N_1273,N_1271);
xnor U1382 (N_1382,N_1293,N_1220);
nor U1383 (N_1383,N_1269,N_1295);
or U1384 (N_1384,N_1272,N_1203);
nor U1385 (N_1385,N_1206,N_1262);
nor U1386 (N_1386,N_1289,N_1234);
nor U1387 (N_1387,N_1217,N_1278);
nor U1388 (N_1388,N_1287,N_1223);
and U1389 (N_1389,N_1208,N_1204);
nor U1390 (N_1390,N_1259,N_1256);
or U1391 (N_1391,N_1227,N_1219);
xor U1392 (N_1392,N_1256,N_1266);
nand U1393 (N_1393,N_1238,N_1242);
nand U1394 (N_1394,N_1265,N_1230);
xnor U1395 (N_1395,N_1214,N_1202);
nor U1396 (N_1396,N_1273,N_1224);
and U1397 (N_1397,N_1298,N_1223);
and U1398 (N_1398,N_1208,N_1297);
and U1399 (N_1399,N_1267,N_1217);
nand U1400 (N_1400,N_1387,N_1344);
and U1401 (N_1401,N_1301,N_1310);
nand U1402 (N_1402,N_1336,N_1312);
nand U1403 (N_1403,N_1369,N_1314);
and U1404 (N_1404,N_1306,N_1393);
and U1405 (N_1405,N_1321,N_1383);
xnor U1406 (N_1406,N_1315,N_1390);
and U1407 (N_1407,N_1395,N_1368);
xnor U1408 (N_1408,N_1363,N_1349);
or U1409 (N_1409,N_1318,N_1392);
nor U1410 (N_1410,N_1332,N_1367);
or U1411 (N_1411,N_1302,N_1348);
and U1412 (N_1412,N_1355,N_1356);
and U1413 (N_1413,N_1343,N_1325);
or U1414 (N_1414,N_1347,N_1364);
nor U1415 (N_1415,N_1308,N_1326);
nor U1416 (N_1416,N_1388,N_1338);
or U1417 (N_1417,N_1305,N_1328);
and U1418 (N_1418,N_1397,N_1319);
nand U1419 (N_1419,N_1381,N_1375);
and U1420 (N_1420,N_1307,N_1396);
nor U1421 (N_1421,N_1334,N_1330);
and U1422 (N_1422,N_1317,N_1360);
nand U1423 (N_1423,N_1399,N_1351);
xnor U1424 (N_1424,N_1300,N_1359);
xor U1425 (N_1425,N_1385,N_1362);
nand U1426 (N_1426,N_1384,N_1389);
xor U1427 (N_1427,N_1374,N_1398);
or U1428 (N_1428,N_1373,N_1358);
and U1429 (N_1429,N_1333,N_1340);
or U1430 (N_1430,N_1377,N_1323);
and U1431 (N_1431,N_1366,N_1357);
or U1432 (N_1432,N_1391,N_1331);
or U1433 (N_1433,N_1345,N_1311);
xnor U1434 (N_1434,N_1346,N_1341);
xor U1435 (N_1435,N_1322,N_1320);
and U1436 (N_1436,N_1342,N_1379);
xor U1437 (N_1437,N_1339,N_1376);
nand U1438 (N_1438,N_1371,N_1303);
nor U1439 (N_1439,N_1354,N_1353);
nand U1440 (N_1440,N_1372,N_1316);
nor U1441 (N_1441,N_1327,N_1313);
xor U1442 (N_1442,N_1309,N_1335);
and U1443 (N_1443,N_1361,N_1352);
nand U1444 (N_1444,N_1337,N_1386);
or U1445 (N_1445,N_1350,N_1382);
or U1446 (N_1446,N_1380,N_1365);
nor U1447 (N_1447,N_1324,N_1304);
nand U1448 (N_1448,N_1329,N_1378);
nand U1449 (N_1449,N_1370,N_1394);
nand U1450 (N_1450,N_1322,N_1366);
xnor U1451 (N_1451,N_1363,N_1356);
or U1452 (N_1452,N_1312,N_1322);
nand U1453 (N_1453,N_1356,N_1315);
xnor U1454 (N_1454,N_1353,N_1325);
nand U1455 (N_1455,N_1344,N_1351);
or U1456 (N_1456,N_1354,N_1373);
nor U1457 (N_1457,N_1392,N_1326);
nor U1458 (N_1458,N_1348,N_1386);
or U1459 (N_1459,N_1310,N_1374);
xor U1460 (N_1460,N_1374,N_1355);
and U1461 (N_1461,N_1333,N_1337);
and U1462 (N_1462,N_1393,N_1313);
nor U1463 (N_1463,N_1327,N_1322);
and U1464 (N_1464,N_1366,N_1394);
nand U1465 (N_1465,N_1329,N_1374);
xor U1466 (N_1466,N_1358,N_1320);
xor U1467 (N_1467,N_1373,N_1332);
nand U1468 (N_1468,N_1391,N_1388);
xor U1469 (N_1469,N_1352,N_1345);
nand U1470 (N_1470,N_1322,N_1336);
xnor U1471 (N_1471,N_1352,N_1311);
and U1472 (N_1472,N_1371,N_1381);
nand U1473 (N_1473,N_1368,N_1314);
or U1474 (N_1474,N_1397,N_1346);
and U1475 (N_1475,N_1366,N_1302);
xor U1476 (N_1476,N_1319,N_1359);
and U1477 (N_1477,N_1365,N_1304);
or U1478 (N_1478,N_1331,N_1340);
and U1479 (N_1479,N_1354,N_1367);
and U1480 (N_1480,N_1380,N_1312);
and U1481 (N_1481,N_1340,N_1396);
nand U1482 (N_1482,N_1312,N_1342);
xnor U1483 (N_1483,N_1336,N_1367);
nand U1484 (N_1484,N_1346,N_1311);
and U1485 (N_1485,N_1320,N_1363);
nand U1486 (N_1486,N_1341,N_1372);
nor U1487 (N_1487,N_1387,N_1366);
and U1488 (N_1488,N_1387,N_1388);
xnor U1489 (N_1489,N_1365,N_1300);
or U1490 (N_1490,N_1321,N_1324);
or U1491 (N_1491,N_1340,N_1390);
xnor U1492 (N_1492,N_1301,N_1378);
and U1493 (N_1493,N_1352,N_1386);
xnor U1494 (N_1494,N_1363,N_1301);
or U1495 (N_1495,N_1373,N_1313);
or U1496 (N_1496,N_1356,N_1384);
nand U1497 (N_1497,N_1310,N_1314);
nor U1498 (N_1498,N_1308,N_1374);
nand U1499 (N_1499,N_1376,N_1360);
and U1500 (N_1500,N_1426,N_1438);
or U1501 (N_1501,N_1451,N_1432);
nor U1502 (N_1502,N_1462,N_1455);
nor U1503 (N_1503,N_1402,N_1437);
xnor U1504 (N_1504,N_1401,N_1499);
or U1505 (N_1505,N_1420,N_1476);
xnor U1506 (N_1506,N_1453,N_1496);
and U1507 (N_1507,N_1443,N_1404);
xnor U1508 (N_1508,N_1460,N_1471);
nor U1509 (N_1509,N_1465,N_1457);
and U1510 (N_1510,N_1492,N_1434);
or U1511 (N_1511,N_1486,N_1487);
and U1512 (N_1512,N_1405,N_1447);
xor U1513 (N_1513,N_1407,N_1418);
and U1514 (N_1514,N_1424,N_1469);
nand U1515 (N_1515,N_1421,N_1417);
xor U1516 (N_1516,N_1473,N_1400);
nand U1517 (N_1517,N_1456,N_1406);
xnor U1518 (N_1518,N_1411,N_1475);
or U1519 (N_1519,N_1498,N_1454);
xnor U1520 (N_1520,N_1415,N_1441);
nor U1521 (N_1521,N_1495,N_1450);
xnor U1522 (N_1522,N_1408,N_1419);
nor U1523 (N_1523,N_1482,N_1466);
or U1524 (N_1524,N_1461,N_1413);
nor U1525 (N_1525,N_1468,N_1479);
xnor U1526 (N_1526,N_1427,N_1483);
and U1527 (N_1527,N_1409,N_1422);
nor U1528 (N_1528,N_1429,N_1481);
or U1529 (N_1529,N_1464,N_1403);
nand U1530 (N_1530,N_1412,N_1458);
nor U1531 (N_1531,N_1414,N_1459);
and U1532 (N_1532,N_1439,N_1449);
and U1533 (N_1533,N_1440,N_1490);
and U1534 (N_1534,N_1474,N_1425);
nor U1535 (N_1535,N_1431,N_1444);
xor U1536 (N_1536,N_1477,N_1493);
xor U1537 (N_1537,N_1442,N_1430);
and U1538 (N_1538,N_1423,N_1435);
nor U1539 (N_1539,N_1436,N_1448);
or U1540 (N_1540,N_1488,N_1470);
or U1541 (N_1541,N_1472,N_1467);
nor U1542 (N_1542,N_1433,N_1480);
xor U1543 (N_1543,N_1446,N_1478);
xor U1544 (N_1544,N_1489,N_1410);
or U1545 (N_1545,N_1428,N_1494);
nand U1546 (N_1546,N_1463,N_1416);
and U1547 (N_1547,N_1445,N_1497);
or U1548 (N_1548,N_1484,N_1485);
xor U1549 (N_1549,N_1452,N_1491);
xnor U1550 (N_1550,N_1428,N_1409);
xnor U1551 (N_1551,N_1416,N_1426);
or U1552 (N_1552,N_1497,N_1460);
nor U1553 (N_1553,N_1468,N_1488);
nor U1554 (N_1554,N_1495,N_1414);
and U1555 (N_1555,N_1430,N_1450);
nand U1556 (N_1556,N_1410,N_1443);
xor U1557 (N_1557,N_1465,N_1424);
nor U1558 (N_1558,N_1443,N_1482);
xor U1559 (N_1559,N_1424,N_1405);
nand U1560 (N_1560,N_1460,N_1408);
or U1561 (N_1561,N_1409,N_1498);
xnor U1562 (N_1562,N_1427,N_1439);
or U1563 (N_1563,N_1455,N_1449);
nand U1564 (N_1564,N_1488,N_1442);
and U1565 (N_1565,N_1429,N_1453);
nor U1566 (N_1566,N_1425,N_1438);
and U1567 (N_1567,N_1420,N_1419);
xor U1568 (N_1568,N_1444,N_1418);
xnor U1569 (N_1569,N_1413,N_1425);
and U1570 (N_1570,N_1405,N_1427);
nand U1571 (N_1571,N_1411,N_1400);
or U1572 (N_1572,N_1408,N_1424);
nor U1573 (N_1573,N_1469,N_1452);
nand U1574 (N_1574,N_1495,N_1482);
xnor U1575 (N_1575,N_1401,N_1496);
and U1576 (N_1576,N_1454,N_1487);
or U1577 (N_1577,N_1467,N_1454);
nand U1578 (N_1578,N_1405,N_1496);
nand U1579 (N_1579,N_1475,N_1452);
and U1580 (N_1580,N_1461,N_1478);
and U1581 (N_1581,N_1486,N_1443);
or U1582 (N_1582,N_1445,N_1485);
xor U1583 (N_1583,N_1480,N_1449);
and U1584 (N_1584,N_1461,N_1437);
xnor U1585 (N_1585,N_1488,N_1485);
nand U1586 (N_1586,N_1450,N_1465);
and U1587 (N_1587,N_1495,N_1481);
and U1588 (N_1588,N_1416,N_1488);
nand U1589 (N_1589,N_1432,N_1480);
or U1590 (N_1590,N_1477,N_1409);
nand U1591 (N_1591,N_1414,N_1418);
nand U1592 (N_1592,N_1483,N_1479);
nand U1593 (N_1593,N_1425,N_1487);
nand U1594 (N_1594,N_1440,N_1470);
xor U1595 (N_1595,N_1427,N_1417);
nor U1596 (N_1596,N_1415,N_1499);
nand U1597 (N_1597,N_1476,N_1442);
xnor U1598 (N_1598,N_1413,N_1434);
or U1599 (N_1599,N_1417,N_1462);
and U1600 (N_1600,N_1548,N_1582);
and U1601 (N_1601,N_1580,N_1558);
nor U1602 (N_1602,N_1562,N_1519);
and U1603 (N_1603,N_1570,N_1573);
xor U1604 (N_1604,N_1521,N_1599);
nor U1605 (N_1605,N_1546,N_1515);
and U1606 (N_1606,N_1592,N_1528);
nand U1607 (N_1607,N_1527,N_1577);
and U1608 (N_1608,N_1524,N_1538);
xor U1609 (N_1609,N_1550,N_1532);
xnor U1610 (N_1610,N_1554,N_1531);
and U1611 (N_1611,N_1574,N_1537);
nand U1612 (N_1612,N_1503,N_1506);
and U1613 (N_1613,N_1513,N_1545);
xor U1614 (N_1614,N_1584,N_1539);
or U1615 (N_1615,N_1501,N_1526);
nor U1616 (N_1616,N_1543,N_1510);
nor U1617 (N_1617,N_1585,N_1564);
xnor U1618 (N_1618,N_1568,N_1552);
nor U1619 (N_1619,N_1504,N_1575);
and U1620 (N_1620,N_1502,N_1511);
or U1621 (N_1621,N_1572,N_1597);
or U1622 (N_1622,N_1508,N_1598);
nor U1623 (N_1623,N_1540,N_1533);
and U1624 (N_1624,N_1505,N_1518);
nor U1625 (N_1625,N_1516,N_1517);
and U1626 (N_1626,N_1593,N_1587);
and U1627 (N_1627,N_1509,N_1530);
xor U1628 (N_1628,N_1520,N_1522);
xor U1629 (N_1629,N_1547,N_1535);
and U1630 (N_1630,N_1579,N_1595);
xnor U1631 (N_1631,N_1523,N_1559);
xor U1632 (N_1632,N_1553,N_1561);
nor U1633 (N_1633,N_1560,N_1542);
xor U1634 (N_1634,N_1544,N_1514);
and U1635 (N_1635,N_1500,N_1565);
nand U1636 (N_1636,N_1571,N_1594);
and U1637 (N_1637,N_1578,N_1557);
nor U1638 (N_1638,N_1576,N_1529);
nor U1639 (N_1639,N_1507,N_1569);
xnor U1640 (N_1640,N_1536,N_1541);
xor U1641 (N_1641,N_1555,N_1566);
and U1642 (N_1642,N_1588,N_1586);
xnor U1643 (N_1643,N_1534,N_1551);
nor U1644 (N_1644,N_1590,N_1556);
nand U1645 (N_1645,N_1549,N_1563);
xnor U1646 (N_1646,N_1596,N_1589);
nor U1647 (N_1647,N_1581,N_1512);
nor U1648 (N_1648,N_1583,N_1567);
and U1649 (N_1649,N_1525,N_1591);
and U1650 (N_1650,N_1522,N_1574);
and U1651 (N_1651,N_1567,N_1541);
nor U1652 (N_1652,N_1570,N_1566);
nand U1653 (N_1653,N_1591,N_1585);
xnor U1654 (N_1654,N_1500,N_1517);
and U1655 (N_1655,N_1531,N_1569);
and U1656 (N_1656,N_1534,N_1589);
nand U1657 (N_1657,N_1594,N_1592);
nor U1658 (N_1658,N_1579,N_1526);
and U1659 (N_1659,N_1574,N_1552);
or U1660 (N_1660,N_1522,N_1553);
nand U1661 (N_1661,N_1588,N_1555);
xnor U1662 (N_1662,N_1529,N_1538);
and U1663 (N_1663,N_1525,N_1511);
nor U1664 (N_1664,N_1534,N_1573);
xnor U1665 (N_1665,N_1591,N_1548);
nor U1666 (N_1666,N_1588,N_1544);
or U1667 (N_1667,N_1501,N_1511);
nand U1668 (N_1668,N_1579,N_1515);
nand U1669 (N_1669,N_1518,N_1521);
nor U1670 (N_1670,N_1559,N_1514);
nor U1671 (N_1671,N_1551,N_1545);
and U1672 (N_1672,N_1582,N_1512);
nand U1673 (N_1673,N_1541,N_1532);
and U1674 (N_1674,N_1569,N_1580);
nor U1675 (N_1675,N_1524,N_1509);
xor U1676 (N_1676,N_1587,N_1554);
or U1677 (N_1677,N_1510,N_1534);
and U1678 (N_1678,N_1598,N_1542);
nand U1679 (N_1679,N_1565,N_1527);
and U1680 (N_1680,N_1552,N_1579);
or U1681 (N_1681,N_1534,N_1532);
nand U1682 (N_1682,N_1582,N_1531);
or U1683 (N_1683,N_1573,N_1521);
nand U1684 (N_1684,N_1552,N_1523);
xnor U1685 (N_1685,N_1544,N_1584);
and U1686 (N_1686,N_1529,N_1516);
or U1687 (N_1687,N_1575,N_1535);
xor U1688 (N_1688,N_1563,N_1525);
xnor U1689 (N_1689,N_1519,N_1568);
or U1690 (N_1690,N_1512,N_1553);
xor U1691 (N_1691,N_1500,N_1552);
and U1692 (N_1692,N_1573,N_1583);
or U1693 (N_1693,N_1573,N_1512);
and U1694 (N_1694,N_1584,N_1516);
or U1695 (N_1695,N_1536,N_1553);
nor U1696 (N_1696,N_1519,N_1549);
xnor U1697 (N_1697,N_1535,N_1546);
or U1698 (N_1698,N_1584,N_1503);
or U1699 (N_1699,N_1584,N_1568);
xor U1700 (N_1700,N_1652,N_1613);
and U1701 (N_1701,N_1669,N_1698);
nand U1702 (N_1702,N_1655,N_1658);
and U1703 (N_1703,N_1676,N_1693);
or U1704 (N_1704,N_1646,N_1673);
or U1705 (N_1705,N_1665,N_1647);
nor U1706 (N_1706,N_1650,N_1684);
xor U1707 (N_1707,N_1690,N_1680);
nand U1708 (N_1708,N_1668,N_1622);
nor U1709 (N_1709,N_1695,N_1632);
or U1710 (N_1710,N_1606,N_1687);
and U1711 (N_1711,N_1691,N_1615);
or U1712 (N_1712,N_1628,N_1634);
nand U1713 (N_1713,N_1685,N_1608);
or U1714 (N_1714,N_1683,N_1659);
or U1715 (N_1715,N_1619,N_1630);
nor U1716 (N_1716,N_1636,N_1620);
or U1717 (N_1717,N_1642,N_1679);
or U1718 (N_1718,N_1661,N_1645);
and U1719 (N_1719,N_1618,N_1611);
and U1720 (N_1720,N_1648,N_1604);
xnor U1721 (N_1721,N_1631,N_1629);
xor U1722 (N_1722,N_1670,N_1640);
and U1723 (N_1723,N_1688,N_1654);
xor U1724 (N_1724,N_1637,N_1651);
nand U1725 (N_1725,N_1624,N_1660);
xor U1726 (N_1726,N_1667,N_1638);
and U1727 (N_1727,N_1666,N_1635);
xnor U1728 (N_1728,N_1657,N_1681);
and U1729 (N_1729,N_1614,N_1600);
or U1730 (N_1730,N_1610,N_1694);
or U1731 (N_1731,N_1641,N_1675);
and U1732 (N_1732,N_1612,N_1677);
and U1733 (N_1733,N_1663,N_1686);
or U1734 (N_1734,N_1605,N_1692);
xor U1735 (N_1735,N_1601,N_1649);
nor U1736 (N_1736,N_1625,N_1682);
and U1737 (N_1737,N_1602,N_1616);
or U1738 (N_1738,N_1699,N_1627);
xnor U1739 (N_1739,N_1696,N_1656);
or U1740 (N_1740,N_1633,N_1662);
and U1741 (N_1741,N_1603,N_1644);
nor U1742 (N_1742,N_1609,N_1689);
or U1743 (N_1743,N_1672,N_1674);
xor U1744 (N_1744,N_1617,N_1653);
nand U1745 (N_1745,N_1678,N_1697);
nor U1746 (N_1746,N_1621,N_1623);
nand U1747 (N_1747,N_1639,N_1607);
or U1748 (N_1748,N_1626,N_1664);
or U1749 (N_1749,N_1671,N_1643);
nor U1750 (N_1750,N_1619,N_1656);
or U1751 (N_1751,N_1665,N_1642);
nor U1752 (N_1752,N_1669,N_1626);
nand U1753 (N_1753,N_1633,N_1629);
nand U1754 (N_1754,N_1680,N_1602);
and U1755 (N_1755,N_1638,N_1627);
and U1756 (N_1756,N_1616,N_1614);
nor U1757 (N_1757,N_1699,N_1682);
nand U1758 (N_1758,N_1623,N_1679);
and U1759 (N_1759,N_1603,N_1609);
or U1760 (N_1760,N_1688,N_1628);
or U1761 (N_1761,N_1651,N_1665);
xor U1762 (N_1762,N_1688,N_1659);
xnor U1763 (N_1763,N_1637,N_1619);
xnor U1764 (N_1764,N_1607,N_1626);
and U1765 (N_1765,N_1603,N_1669);
xnor U1766 (N_1766,N_1614,N_1675);
xnor U1767 (N_1767,N_1605,N_1689);
xor U1768 (N_1768,N_1640,N_1699);
nand U1769 (N_1769,N_1654,N_1698);
and U1770 (N_1770,N_1656,N_1634);
and U1771 (N_1771,N_1612,N_1688);
nand U1772 (N_1772,N_1640,N_1685);
nand U1773 (N_1773,N_1601,N_1651);
and U1774 (N_1774,N_1658,N_1628);
nor U1775 (N_1775,N_1663,N_1681);
nor U1776 (N_1776,N_1668,N_1631);
and U1777 (N_1777,N_1685,N_1623);
xor U1778 (N_1778,N_1612,N_1698);
and U1779 (N_1779,N_1620,N_1691);
or U1780 (N_1780,N_1622,N_1636);
nor U1781 (N_1781,N_1670,N_1608);
nor U1782 (N_1782,N_1620,N_1675);
xor U1783 (N_1783,N_1649,N_1694);
xnor U1784 (N_1784,N_1683,N_1611);
xnor U1785 (N_1785,N_1641,N_1625);
and U1786 (N_1786,N_1615,N_1680);
or U1787 (N_1787,N_1600,N_1635);
nand U1788 (N_1788,N_1677,N_1639);
or U1789 (N_1789,N_1640,N_1629);
nor U1790 (N_1790,N_1690,N_1617);
nor U1791 (N_1791,N_1619,N_1660);
nand U1792 (N_1792,N_1656,N_1667);
or U1793 (N_1793,N_1606,N_1600);
xor U1794 (N_1794,N_1696,N_1637);
xor U1795 (N_1795,N_1630,N_1673);
nor U1796 (N_1796,N_1687,N_1664);
and U1797 (N_1797,N_1661,N_1633);
xor U1798 (N_1798,N_1675,N_1619);
nor U1799 (N_1799,N_1697,N_1611);
nand U1800 (N_1800,N_1722,N_1746);
nor U1801 (N_1801,N_1756,N_1788);
and U1802 (N_1802,N_1760,N_1739);
nor U1803 (N_1803,N_1759,N_1798);
nor U1804 (N_1804,N_1753,N_1708);
nor U1805 (N_1805,N_1723,N_1742);
and U1806 (N_1806,N_1777,N_1733);
nor U1807 (N_1807,N_1749,N_1772);
or U1808 (N_1808,N_1719,N_1778);
nor U1809 (N_1809,N_1764,N_1736);
xnor U1810 (N_1810,N_1721,N_1737);
or U1811 (N_1811,N_1754,N_1703);
and U1812 (N_1812,N_1751,N_1757);
nor U1813 (N_1813,N_1713,N_1790);
nand U1814 (N_1814,N_1781,N_1726);
nor U1815 (N_1815,N_1735,N_1785);
and U1816 (N_1816,N_1782,N_1720);
xor U1817 (N_1817,N_1741,N_1780);
and U1818 (N_1818,N_1797,N_1786);
nor U1819 (N_1819,N_1792,N_1745);
xnor U1820 (N_1820,N_1765,N_1775);
or U1821 (N_1821,N_1795,N_1715);
or U1822 (N_1822,N_1705,N_1734);
and U1823 (N_1823,N_1784,N_1766);
nand U1824 (N_1824,N_1768,N_1773);
nor U1825 (N_1825,N_1725,N_1750);
nor U1826 (N_1826,N_1793,N_1730);
xnor U1827 (N_1827,N_1783,N_1702);
and U1828 (N_1828,N_1711,N_1796);
nor U1829 (N_1829,N_1774,N_1752);
and U1830 (N_1830,N_1709,N_1763);
xor U1831 (N_1831,N_1769,N_1762);
and U1832 (N_1832,N_1776,N_1710);
and U1833 (N_1833,N_1714,N_1743);
nor U1834 (N_1834,N_1779,N_1718);
nand U1835 (N_1835,N_1727,N_1712);
nand U1836 (N_1836,N_1787,N_1717);
nor U1837 (N_1837,N_1707,N_1731);
nor U1838 (N_1838,N_1706,N_1794);
or U1839 (N_1839,N_1700,N_1758);
xnor U1840 (N_1840,N_1740,N_1744);
nand U1841 (N_1841,N_1728,N_1791);
nand U1842 (N_1842,N_1770,N_1789);
nand U1843 (N_1843,N_1738,N_1701);
and U1844 (N_1844,N_1767,N_1771);
and U1845 (N_1845,N_1761,N_1716);
nor U1846 (N_1846,N_1747,N_1799);
and U1847 (N_1847,N_1704,N_1724);
xnor U1848 (N_1848,N_1748,N_1755);
nand U1849 (N_1849,N_1729,N_1732);
nand U1850 (N_1850,N_1783,N_1741);
nand U1851 (N_1851,N_1732,N_1707);
and U1852 (N_1852,N_1783,N_1780);
nand U1853 (N_1853,N_1716,N_1786);
or U1854 (N_1854,N_1776,N_1735);
nand U1855 (N_1855,N_1719,N_1738);
or U1856 (N_1856,N_1772,N_1777);
nand U1857 (N_1857,N_1715,N_1796);
xnor U1858 (N_1858,N_1711,N_1794);
and U1859 (N_1859,N_1766,N_1713);
nand U1860 (N_1860,N_1768,N_1782);
and U1861 (N_1861,N_1768,N_1746);
nand U1862 (N_1862,N_1771,N_1708);
xnor U1863 (N_1863,N_1750,N_1753);
or U1864 (N_1864,N_1733,N_1789);
nor U1865 (N_1865,N_1762,N_1724);
nor U1866 (N_1866,N_1791,N_1720);
nor U1867 (N_1867,N_1749,N_1745);
xor U1868 (N_1868,N_1798,N_1792);
nor U1869 (N_1869,N_1770,N_1781);
and U1870 (N_1870,N_1716,N_1723);
and U1871 (N_1871,N_1759,N_1743);
xor U1872 (N_1872,N_1765,N_1774);
nor U1873 (N_1873,N_1782,N_1728);
xor U1874 (N_1874,N_1785,N_1769);
xor U1875 (N_1875,N_1724,N_1799);
nand U1876 (N_1876,N_1743,N_1740);
or U1877 (N_1877,N_1704,N_1754);
and U1878 (N_1878,N_1707,N_1706);
nand U1879 (N_1879,N_1726,N_1792);
and U1880 (N_1880,N_1762,N_1754);
xor U1881 (N_1881,N_1731,N_1704);
and U1882 (N_1882,N_1720,N_1716);
and U1883 (N_1883,N_1724,N_1735);
and U1884 (N_1884,N_1721,N_1761);
or U1885 (N_1885,N_1743,N_1798);
xnor U1886 (N_1886,N_1757,N_1756);
nand U1887 (N_1887,N_1775,N_1774);
xor U1888 (N_1888,N_1732,N_1736);
nand U1889 (N_1889,N_1765,N_1762);
nand U1890 (N_1890,N_1772,N_1713);
nor U1891 (N_1891,N_1761,N_1756);
and U1892 (N_1892,N_1758,N_1740);
xor U1893 (N_1893,N_1728,N_1708);
and U1894 (N_1894,N_1719,N_1795);
and U1895 (N_1895,N_1772,N_1752);
and U1896 (N_1896,N_1707,N_1719);
nor U1897 (N_1897,N_1793,N_1742);
nor U1898 (N_1898,N_1719,N_1798);
and U1899 (N_1899,N_1781,N_1794);
nand U1900 (N_1900,N_1838,N_1812);
nand U1901 (N_1901,N_1817,N_1860);
xnor U1902 (N_1902,N_1814,N_1876);
nor U1903 (N_1903,N_1884,N_1865);
xor U1904 (N_1904,N_1843,N_1820);
or U1905 (N_1905,N_1804,N_1867);
xnor U1906 (N_1906,N_1844,N_1894);
and U1907 (N_1907,N_1828,N_1855);
or U1908 (N_1908,N_1866,N_1861);
nand U1909 (N_1909,N_1898,N_1875);
xor U1910 (N_1910,N_1888,N_1889);
nand U1911 (N_1911,N_1895,N_1849);
or U1912 (N_1912,N_1878,N_1822);
and U1913 (N_1913,N_1803,N_1858);
xor U1914 (N_1914,N_1864,N_1829);
xnor U1915 (N_1915,N_1863,N_1852);
or U1916 (N_1916,N_1841,N_1827);
nand U1917 (N_1917,N_1837,N_1887);
nand U1918 (N_1918,N_1802,N_1824);
and U1919 (N_1919,N_1856,N_1857);
nor U1920 (N_1920,N_1809,N_1813);
xnor U1921 (N_1921,N_1868,N_1810);
or U1922 (N_1922,N_1859,N_1872);
nand U1923 (N_1923,N_1883,N_1899);
nor U1924 (N_1924,N_1836,N_1873);
and U1925 (N_1925,N_1818,N_1826);
nor U1926 (N_1926,N_1877,N_1821);
nor U1927 (N_1927,N_1808,N_1886);
xnor U1928 (N_1928,N_1893,N_1806);
nand U1929 (N_1929,N_1891,N_1871);
xor U1930 (N_1930,N_1846,N_1835);
or U1931 (N_1931,N_1879,N_1851);
or U1932 (N_1932,N_1834,N_1854);
or U1933 (N_1933,N_1823,N_1830);
and U1934 (N_1934,N_1832,N_1825);
nand U1935 (N_1935,N_1845,N_1885);
or U1936 (N_1936,N_1840,N_1819);
and U1937 (N_1937,N_1890,N_1897);
nor U1938 (N_1938,N_1811,N_1839);
nor U1939 (N_1939,N_1869,N_1880);
and U1940 (N_1940,N_1831,N_1816);
nand U1941 (N_1941,N_1833,N_1847);
and U1942 (N_1942,N_1850,N_1882);
or U1943 (N_1943,N_1801,N_1842);
xnor U1944 (N_1944,N_1853,N_1862);
nor U1945 (N_1945,N_1815,N_1892);
and U1946 (N_1946,N_1848,N_1896);
or U1947 (N_1947,N_1874,N_1881);
and U1948 (N_1948,N_1807,N_1870);
or U1949 (N_1949,N_1805,N_1800);
or U1950 (N_1950,N_1830,N_1843);
nand U1951 (N_1951,N_1876,N_1823);
and U1952 (N_1952,N_1856,N_1825);
and U1953 (N_1953,N_1819,N_1858);
nor U1954 (N_1954,N_1861,N_1882);
nor U1955 (N_1955,N_1845,N_1897);
xnor U1956 (N_1956,N_1852,N_1872);
nand U1957 (N_1957,N_1888,N_1890);
and U1958 (N_1958,N_1828,N_1806);
nand U1959 (N_1959,N_1890,N_1823);
nand U1960 (N_1960,N_1893,N_1820);
xor U1961 (N_1961,N_1898,N_1866);
nand U1962 (N_1962,N_1852,N_1874);
and U1963 (N_1963,N_1860,N_1874);
nand U1964 (N_1964,N_1813,N_1839);
and U1965 (N_1965,N_1821,N_1889);
nor U1966 (N_1966,N_1808,N_1813);
and U1967 (N_1967,N_1818,N_1882);
nor U1968 (N_1968,N_1893,N_1895);
and U1969 (N_1969,N_1839,N_1826);
xor U1970 (N_1970,N_1822,N_1820);
and U1971 (N_1971,N_1840,N_1848);
and U1972 (N_1972,N_1837,N_1890);
nor U1973 (N_1973,N_1848,N_1841);
xor U1974 (N_1974,N_1843,N_1816);
xnor U1975 (N_1975,N_1861,N_1837);
xor U1976 (N_1976,N_1880,N_1813);
nor U1977 (N_1977,N_1845,N_1879);
nor U1978 (N_1978,N_1855,N_1893);
or U1979 (N_1979,N_1859,N_1863);
nor U1980 (N_1980,N_1863,N_1825);
nor U1981 (N_1981,N_1894,N_1803);
nor U1982 (N_1982,N_1805,N_1888);
and U1983 (N_1983,N_1809,N_1839);
or U1984 (N_1984,N_1810,N_1830);
nand U1985 (N_1985,N_1858,N_1830);
or U1986 (N_1986,N_1834,N_1892);
and U1987 (N_1987,N_1825,N_1803);
and U1988 (N_1988,N_1864,N_1827);
and U1989 (N_1989,N_1821,N_1891);
or U1990 (N_1990,N_1842,N_1807);
or U1991 (N_1991,N_1897,N_1858);
nor U1992 (N_1992,N_1843,N_1879);
and U1993 (N_1993,N_1880,N_1802);
or U1994 (N_1994,N_1895,N_1839);
or U1995 (N_1995,N_1892,N_1817);
nand U1996 (N_1996,N_1808,N_1819);
nand U1997 (N_1997,N_1838,N_1807);
nand U1998 (N_1998,N_1834,N_1829);
and U1999 (N_1999,N_1803,N_1821);
nand U2000 (N_2000,N_1957,N_1970);
nand U2001 (N_2001,N_1959,N_1920);
and U2002 (N_2002,N_1968,N_1911);
or U2003 (N_2003,N_1938,N_1993);
or U2004 (N_2004,N_1994,N_1985);
or U2005 (N_2005,N_1997,N_1978);
xor U2006 (N_2006,N_1928,N_1908);
xor U2007 (N_2007,N_1914,N_1919);
or U2008 (N_2008,N_1945,N_1934);
nand U2009 (N_2009,N_1958,N_1947);
nor U2010 (N_2010,N_1989,N_1998);
or U2011 (N_2011,N_1984,N_1955);
nor U2012 (N_2012,N_1999,N_1922);
nor U2013 (N_2013,N_1943,N_1988);
or U2014 (N_2014,N_1979,N_1940);
xnor U2015 (N_2015,N_1996,N_1921);
or U2016 (N_2016,N_1916,N_1933);
nand U2017 (N_2017,N_1949,N_1965);
xor U2018 (N_2018,N_1924,N_1967);
and U2019 (N_2019,N_1910,N_1926);
nand U2020 (N_2020,N_1953,N_1982);
and U2021 (N_2021,N_1929,N_1927);
nand U2022 (N_2022,N_1952,N_1944);
xor U2023 (N_2023,N_1975,N_1905);
nand U2024 (N_2024,N_1976,N_1939);
nor U2025 (N_2025,N_1981,N_1969);
or U2026 (N_2026,N_1901,N_1960);
nor U2027 (N_2027,N_1980,N_1937);
nor U2028 (N_2028,N_1942,N_1956);
nor U2029 (N_2029,N_1948,N_1932);
nor U2030 (N_2030,N_1931,N_1986);
nor U2031 (N_2031,N_1992,N_1990);
nand U2032 (N_2032,N_1963,N_1917);
and U2033 (N_2033,N_1961,N_1983);
and U2034 (N_2034,N_1936,N_1966);
or U2035 (N_2035,N_1902,N_1918);
and U2036 (N_2036,N_1904,N_1972);
or U2037 (N_2037,N_1935,N_1909);
xnor U2038 (N_2038,N_1946,N_1971);
or U2039 (N_2039,N_1923,N_1900);
nand U2040 (N_2040,N_1930,N_1954);
and U2041 (N_2041,N_1951,N_1964);
nand U2042 (N_2042,N_1913,N_1950);
and U2043 (N_2043,N_1912,N_1907);
or U2044 (N_2044,N_1925,N_1962);
nor U2045 (N_2045,N_1974,N_1915);
nor U2046 (N_2046,N_1995,N_1903);
nor U2047 (N_2047,N_1941,N_1991);
or U2048 (N_2048,N_1987,N_1977);
and U2049 (N_2049,N_1906,N_1973);
or U2050 (N_2050,N_1963,N_1910);
nor U2051 (N_2051,N_1927,N_1922);
and U2052 (N_2052,N_1948,N_1929);
nand U2053 (N_2053,N_1906,N_1986);
nor U2054 (N_2054,N_1926,N_1967);
nor U2055 (N_2055,N_1948,N_1958);
nand U2056 (N_2056,N_1908,N_1917);
and U2057 (N_2057,N_1933,N_1998);
or U2058 (N_2058,N_1916,N_1967);
or U2059 (N_2059,N_1917,N_1968);
nor U2060 (N_2060,N_1981,N_1918);
nand U2061 (N_2061,N_1912,N_1994);
nand U2062 (N_2062,N_1934,N_1969);
and U2063 (N_2063,N_1929,N_1998);
nor U2064 (N_2064,N_1907,N_1917);
and U2065 (N_2065,N_1970,N_1999);
and U2066 (N_2066,N_1940,N_1937);
and U2067 (N_2067,N_1920,N_1958);
or U2068 (N_2068,N_1970,N_1916);
nor U2069 (N_2069,N_1957,N_1916);
or U2070 (N_2070,N_1934,N_1975);
or U2071 (N_2071,N_1961,N_1954);
nand U2072 (N_2072,N_1907,N_1962);
xor U2073 (N_2073,N_1938,N_1987);
or U2074 (N_2074,N_1960,N_1929);
nor U2075 (N_2075,N_1966,N_1984);
xor U2076 (N_2076,N_1955,N_1961);
nor U2077 (N_2077,N_1936,N_1942);
nand U2078 (N_2078,N_1969,N_1974);
nor U2079 (N_2079,N_1900,N_1913);
nand U2080 (N_2080,N_1958,N_1951);
nand U2081 (N_2081,N_1930,N_1959);
nor U2082 (N_2082,N_1969,N_1999);
and U2083 (N_2083,N_1969,N_1910);
xnor U2084 (N_2084,N_1934,N_1996);
xnor U2085 (N_2085,N_1985,N_1934);
or U2086 (N_2086,N_1929,N_1996);
and U2087 (N_2087,N_1957,N_1918);
and U2088 (N_2088,N_1970,N_1982);
and U2089 (N_2089,N_1993,N_1920);
and U2090 (N_2090,N_1958,N_1956);
nand U2091 (N_2091,N_1934,N_1964);
xnor U2092 (N_2092,N_1983,N_1935);
and U2093 (N_2093,N_1924,N_1968);
xnor U2094 (N_2094,N_1962,N_1939);
and U2095 (N_2095,N_1910,N_1906);
and U2096 (N_2096,N_1998,N_1990);
or U2097 (N_2097,N_1931,N_1962);
and U2098 (N_2098,N_1935,N_1930);
or U2099 (N_2099,N_1920,N_1907);
nand U2100 (N_2100,N_2000,N_2009);
nand U2101 (N_2101,N_2039,N_2014);
or U2102 (N_2102,N_2035,N_2092);
nand U2103 (N_2103,N_2001,N_2048);
nor U2104 (N_2104,N_2062,N_2013);
and U2105 (N_2105,N_2073,N_2004);
xor U2106 (N_2106,N_2057,N_2074);
and U2107 (N_2107,N_2064,N_2012);
and U2108 (N_2108,N_2082,N_2026);
and U2109 (N_2109,N_2003,N_2088);
and U2110 (N_2110,N_2091,N_2005);
or U2111 (N_2111,N_2095,N_2090);
xnor U2112 (N_2112,N_2018,N_2032);
and U2113 (N_2113,N_2008,N_2072);
nand U2114 (N_2114,N_2042,N_2036);
or U2115 (N_2115,N_2098,N_2029);
and U2116 (N_2116,N_2099,N_2031);
or U2117 (N_2117,N_2030,N_2034);
nand U2118 (N_2118,N_2015,N_2081);
or U2119 (N_2119,N_2017,N_2068);
nor U2120 (N_2120,N_2071,N_2006);
nand U2121 (N_2121,N_2046,N_2043);
and U2122 (N_2122,N_2045,N_2033);
nor U2123 (N_2123,N_2075,N_2019);
and U2124 (N_2124,N_2002,N_2021);
or U2125 (N_2125,N_2084,N_2060);
nor U2126 (N_2126,N_2067,N_2007);
nand U2127 (N_2127,N_2097,N_2028);
xor U2128 (N_2128,N_2051,N_2023);
nor U2129 (N_2129,N_2038,N_2079);
nor U2130 (N_2130,N_2083,N_2096);
nor U2131 (N_2131,N_2011,N_2055);
nand U2132 (N_2132,N_2027,N_2087);
nand U2133 (N_2133,N_2093,N_2065);
or U2134 (N_2134,N_2010,N_2020);
and U2135 (N_2135,N_2063,N_2049);
and U2136 (N_2136,N_2086,N_2054);
nand U2137 (N_2137,N_2066,N_2070);
or U2138 (N_2138,N_2077,N_2052);
or U2139 (N_2139,N_2040,N_2047);
or U2140 (N_2140,N_2050,N_2058);
xor U2141 (N_2141,N_2085,N_2094);
nor U2142 (N_2142,N_2041,N_2044);
or U2143 (N_2143,N_2024,N_2037);
and U2144 (N_2144,N_2069,N_2056);
or U2145 (N_2145,N_2076,N_2025);
nor U2146 (N_2146,N_2016,N_2061);
nor U2147 (N_2147,N_2089,N_2053);
xnor U2148 (N_2148,N_2078,N_2059);
or U2149 (N_2149,N_2080,N_2022);
nand U2150 (N_2150,N_2072,N_2047);
or U2151 (N_2151,N_2038,N_2043);
or U2152 (N_2152,N_2007,N_2029);
and U2153 (N_2153,N_2098,N_2063);
and U2154 (N_2154,N_2086,N_2029);
nor U2155 (N_2155,N_2018,N_2042);
nand U2156 (N_2156,N_2044,N_2067);
nand U2157 (N_2157,N_2059,N_2049);
and U2158 (N_2158,N_2022,N_2013);
and U2159 (N_2159,N_2092,N_2052);
nor U2160 (N_2160,N_2084,N_2091);
xnor U2161 (N_2161,N_2027,N_2068);
and U2162 (N_2162,N_2036,N_2044);
and U2163 (N_2163,N_2063,N_2004);
or U2164 (N_2164,N_2030,N_2087);
xnor U2165 (N_2165,N_2007,N_2055);
and U2166 (N_2166,N_2073,N_2072);
xnor U2167 (N_2167,N_2074,N_2019);
and U2168 (N_2168,N_2097,N_2025);
nand U2169 (N_2169,N_2078,N_2045);
and U2170 (N_2170,N_2005,N_2055);
nor U2171 (N_2171,N_2006,N_2027);
nor U2172 (N_2172,N_2031,N_2029);
nor U2173 (N_2173,N_2080,N_2060);
nor U2174 (N_2174,N_2086,N_2021);
nor U2175 (N_2175,N_2036,N_2013);
or U2176 (N_2176,N_2022,N_2040);
xor U2177 (N_2177,N_2025,N_2039);
and U2178 (N_2178,N_2073,N_2007);
nand U2179 (N_2179,N_2030,N_2018);
nand U2180 (N_2180,N_2082,N_2066);
or U2181 (N_2181,N_2023,N_2013);
xor U2182 (N_2182,N_2059,N_2065);
or U2183 (N_2183,N_2006,N_2017);
xnor U2184 (N_2184,N_2091,N_2024);
xnor U2185 (N_2185,N_2076,N_2000);
nor U2186 (N_2186,N_2011,N_2032);
xor U2187 (N_2187,N_2003,N_2082);
or U2188 (N_2188,N_2011,N_2064);
and U2189 (N_2189,N_2034,N_2056);
or U2190 (N_2190,N_2083,N_2050);
nor U2191 (N_2191,N_2096,N_2047);
or U2192 (N_2192,N_2082,N_2021);
nor U2193 (N_2193,N_2059,N_2013);
xnor U2194 (N_2194,N_2057,N_2049);
xor U2195 (N_2195,N_2030,N_2099);
nand U2196 (N_2196,N_2064,N_2086);
nor U2197 (N_2197,N_2042,N_2059);
nor U2198 (N_2198,N_2029,N_2073);
nand U2199 (N_2199,N_2026,N_2048);
nor U2200 (N_2200,N_2102,N_2129);
nand U2201 (N_2201,N_2177,N_2192);
or U2202 (N_2202,N_2194,N_2196);
nand U2203 (N_2203,N_2113,N_2156);
nor U2204 (N_2204,N_2173,N_2187);
xor U2205 (N_2205,N_2121,N_2162);
nor U2206 (N_2206,N_2106,N_2182);
or U2207 (N_2207,N_2136,N_2188);
nor U2208 (N_2208,N_2138,N_2189);
nor U2209 (N_2209,N_2146,N_2179);
and U2210 (N_2210,N_2122,N_2174);
nand U2211 (N_2211,N_2114,N_2167);
nor U2212 (N_2212,N_2193,N_2153);
xnor U2213 (N_2213,N_2161,N_2152);
nand U2214 (N_2214,N_2186,N_2105);
nand U2215 (N_2215,N_2150,N_2134);
nor U2216 (N_2216,N_2151,N_2139);
and U2217 (N_2217,N_2184,N_2166);
xor U2218 (N_2218,N_2109,N_2130);
xor U2219 (N_2219,N_2128,N_2171);
xor U2220 (N_2220,N_2175,N_2131);
xor U2221 (N_2221,N_2185,N_2147);
and U2222 (N_2222,N_2180,N_2158);
xor U2223 (N_2223,N_2190,N_2198);
or U2224 (N_2224,N_2104,N_2154);
nand U2225 (N_2225,N_2183,N_2110);
nand U2226 (N_2226,N_2123,N_2197);
nand U2227 (N_2227,N_2126,N_2195);
nor U2228 (N_2228,N_2191,N_2143);
nand U2229 (N_2229,N_2165,N_2135);
nand U2230 (N_2230,N_2145,N_2149);
xor U2231 (N_2231,N_2169,N_2148);
and U2232 (N_2232,N_2100,N_2170);
xnor U2233 (N_2233,N_2116,N_2140);
nand U2234 (N_2234,N_2118,N_2157);
nor U2235 (N_2235,N_2181,N_2112);
nand U2236 (N_2236,N_2137,N_2133);
xor U2237 (N_2237,N_2142,N_2125);
or U2238 (N_2238,N_2103,N_2119);
xnor U2239 (N_2239,N_2155,N_2163);
and U2240 (N_2240,N_2107,N_2168);
xnor U2241 (N_2241,N_2141,N_2124);
and U2242 (N_2242,N_2127,N_2132);
and U2243 (N_2243,N_2115,N_2120);
or U2244 (N_2244,N_2159,N_2172);
and U2245 (N_2245,N_2164,N_2178);
and U2246 (N_2246,N_2199,N_2101);
or U2247 (N_2247,N_2160,N_2176);
and U2248 (N_2248,N_2111,N_2117);
nand U2249 (N_2249,N_2144,N_2108);
or U2250 (N_2250,N_2165,N_2182);
xnor U2251 (N_2251,N_2105,N_2122);
and U2252 (N_2252,N_2111,N_2134);
or U2253 (N_2253,N_2182,N_2147);
nor U2254 (N_2254,N_2192,N_2199);
or U2255 (N_2255,N_2138,N_2114);
xor U2256 (N_2256,N_2130,N_2195);
nor U2257 (N_2257,N_2110,N_2171);
nor U2258 (N_2258,N_2115,N_2134);
nor U2259 (N_2259,N_2145,N_2173);
and U2260 (N_2260,N_2185,N_2196);
nor U2261 (N_2261,N_2176,N_2137);
or U2262 (N_2262,N_2170,N_2169);
or U2263 (N_2263,N_2181,N_2188);
or U2264 (N_2264,N_2155,N_2177);
nand U2265 (N_2265,N_2169,N_2154);
xnor U2266 (N_2266,N_2113,N_2120);
nand U2267 (N_2267,N_2133,N_2176);
nor U2268 (N_2268,N_2158,N_2140);
or U2269 (N_2269,N_2108,N_2135);
nand U2270 (N_2270,N_2115,N_2190);
and U2271 (N_2271,N_2189,N_2120);
nand U2272 (N_2272,N_2104,N_2161);
and U2273 (N_2273,N_2153,N_2171);
nand U2274 (N_2274,N_2101,N_2124);
or U2275 (N_2275,N_2174,N_2154);
nand U2276 (N_2276,N_2146,N_2120);
xnor U2277 (N_2277,N_2160,N_2117);
and U2278 (N_2278,N_2181,N_2178);
and U2279 (N_2279,N_2146,N_2108);
nor U2280 (N_2280,N_2124,N_2148);
xnor U2281 (N_2281,N_2145,N_2153);
nor U2282 (N_2282,N_2159,N_2193);
xnor U2283 (N_2283,N_2188,N_2106);
and U2284 (N_2284,N_2161,N_2135);
nand U2285 (N_2285,N_2143,N_2132);
nor U2286 (N_2286,N_2174,N_2120);
and U2287 (N_2287,N_2161,N_2166);
nand U2288 (N_2288,N_2183,N_2168);
and U2289 (N_2289,N_2104,N_2152);
or U2290 (N_2290,N_2122,N_2171);
or U2291 (N_2291,N_2103,N_2163);
and U2292 (N_2292,N_2116,N_2115);
nor U2293 (N_2293,N_2140,N_2103);
nand U2294 (N_2294,N_2100,N_2150);
nand U2295 (N_2295,N_2194,N_2165);
nor U2296 (N_2296,N_2187,N_2137);
nand U2297 (N_2297,N_2184,N_2140);
and U2298 (N_2298,N_2156,N_2163);
xnor U2299 (N_2299,N_2174,N_2151);
nand U2300 (N_2300,N_2271,N_2226);
or U2301 (N_2301,N_2251,N_2265);
nand U2302 (N_2302,N_2259,N_2255);
and U2303 (N_2303,N_2281,N_2266);
or U2304 (N_2304,N_2244,N_2230);
or U2305 (N_2305,N_2212,N_2290);
or U2306 (N_2306,N_2282,N_2224);
or U2307 (N_2307,N_2291,N_2289);
or U2308 (N_2308,N_2200,N_2228);
xor U2309 (N_2309,N_2277,N_2235);
or U2310 (N_2310,N_2258,N_2202);
nor U2311 (N_2311,N_2227,N_2243);
nand U2312 (N_2312,N_2296,N_2247);
or U2313 (N_2313,N_2254,N_2283);
nand U2314 (N_2314,N_2272,N_2245);
and U2315 (N_2315,N_2279,N_2284);
nor U2316 (N_2316,N_2262,N_2299);
nand U2317 (N_2317,N_2252,N_2246);
nor U2318 (N_2318,N_2203,N_2240);
nand U2319 (N_2319,N_2238,N_2273);
and U2320 (N_2320,N_2237,N_2209);
nand U2321 (N_2321,N_2253,N_2270);
nand U2322 (N_2322,N_2286,N_2293);
nor U2323 (N_2323,N_2207,N_2264);
nor U2324 (N_2324,N_2229,N_2216);
xor U2325 (N_2325,N_2278,N_2219);
or U2326 (N_2326,N_2218,N_2234);
nand U2327 (N_2327,N_2269,N_2233);
and U2328 (N_2328,N_2263,N_2280);
nor U2329 (N_2329,N_2221,N_2231);
nor U2330 (N_2330,N_2204,N_2205);
or U2331 (N_2331,N_2220,N_2292);
nand U2332 (N_2332,N_2294,N_2297);
nor U2333 (N_2333,N_2248,N_2239);
or U2334 (N_2334,N_2225,N_2213);
or U2335 (N_2335,N_2260,N_2256);
nor U2336 (N_2336,N_2275,N_2222);
and U2337 (N_2337,N_2208,N_2274);
xnor U2338 (N_2338,N_2267,N_2236);
or U2339 (N_2339,N_2287,N_2232);
or U2340 (N_2340,N_2268,N_2285);
or U2341 (N_2341,N_2261,N_2250);
or U2342 (N_2342,N_2210,N_2206);
or U2343 (N_2343,N_2201,N_2249);
nor U2344 (N_2344,N_2276,N_2211);
xnor U2345 (N_2345,N_2257,N_2288);
xnor U2346 (N_2346,N_2298,N_2215);
and U2347 (N_2347,N_2214,N_2242);
xor U2348 (N_2348,N_2217,N_2241);
and U2349 (N_2349,N_2295,N_2223);
or U2350 (N_2350,N_2284,N_2278);
nor U2351 (N_2351,N_2230,N_2217);
xor U2352 (N_2352,N_2245,N_2291);
or U2353 (N_2353,N_2281,N_2268);
and U2354 (N_2354,N_2213,N_2207);
or U2355 (N_2355,N_2212,N_2252);
and U2356 (N_2356,N_2267,N_2253);
nand U2357 (N_2357,N_2247,N_2298);
or U2358 (N_2358,N_2286,N_2234);
xor U2359 (N_2359,N_2211,N_2258);
nand U2360 (N_2360,N_2239,N_2219);
nor U2361 (N_2361,N_2289,N_2224);
nor U2362 (N_2362,N_2211,N_2212);
or U2363 (N_2363,N_2297,N_2221);
or U2364 (N_2364,N_2212,N_2289);
nor U2365 (N_2365,N_2267,N_2231);
nor U2366 (N_2366,N_2288,N_2249);
xnor U2367 (N_2367,N_2228,N_2292);
xor U2368 (N_2368,N_2279,N_2267);
and U2369 (N_2369,N_2258,N_2273);
nand U2370 (N_2370,N_2298,N_2235);
nand U2371 (N_2371,N_2251,N_2225);
nand U2372 (N_2372,N_2208,N_2242);
xnor U2373 (N_2373,N_2240,N_2273);
nor U2374 (N_2374,N_2290,N_2279);
xor U2375 (N_2375,N_2290,N_2248);
or U2376 (N_2376,N_2208,N_2291);
xnor U2377 (N_2377,N_2249,N_2257);
or U2378 (N_2378,N_2220,N_2286);
nand U2379 (N_2379,N_2236,N_2245);
or U2380 (N_2380,N_2276,N_2273);
or U2381 (N_2381,N_2248,N_2259);
xor U2382 (N_2382,N_2289,N_2297);
xnor U2383 (N_2383,N_2274,N_2231);
nand U2384 (N_2384,N_2248,N_2271);
xnor U2385 (N_2385,N_2235,N_2210);
xnor U2386 (N_2386,N_2225,N_2276);
xor U2387 (N_2387,N_2240,N_2299);
nand U2388 (N_2388,N_2232,N_2273);
nand U2389 (N_2389,N_2242,N_2274);
nand U2390 (N_2390,N_2295,N_2252);
and U2391 (N_2391,N_2273,N_2212);
or U2392 (N_2392,N_2267,N_2257);
nand U2393 (N_2393,N_2249,N_2269);
and U2394 (N_2394,N_2218,N_2233);
nand U2395 (N_2395,N_2228,N_2235);
nand U2396 (N_2396,N_2215,N_2274);
or U2397 (N_2397,N_2255,N_2223);
xnor U2398 (N_2398,N_2243,N_2200);
xnor U2399 (N_2399,N_2202,N_2265);
nor U2400 (N_2400,N_2370,N_2346);
xor U2401 (N_2401,N_2340,N_2312);
nor U2402 (N_2402,N_2380,N_2399);
nand U2403 (N_2403,N_2342,N_2389);
nand U2404 (N_2404,N_2384,N_2352);
or U2405 (N_2405,N_2390,N_2328);
nor U2406 (N_2406,N_2381,N_2307);
nor U2407 (N_2407,N_2331,N_2333);
nand U2408 (N_2408,N_2336,N_2366);
nand U2409 (N_2409,N_2396,N_2337);
and U2410 (N_2410,N_2383,N_2388);
or U2411 (N_2411,N_2315,N_2357);
nand U2412 (N_2412,N_2364,N_2371);
and U2413 (N_2413,N_2304,N_2311);
or U2414 (N_2414,N_2393,N_2392);
nor U2415 (N_2415,N_2395,N_2375);
and U2416 (N_2416,N_2317,N_2313);
and U2417 (N_2417,N_2361,N_2363);
nor U2418 (N_2418,N_2324,N_2398);
xor U2419 (N_2419,N_2308,N_2314);
xnor U2420 (N_2420,N_2377,N_2385);
xor U2421 (N_2421,N_2330,N_2368);
xnor U2422 (N_2422,N_2347,N_2353);
xor U2423 (N_2423,N_2365,N_2391);
nand U2424 (N_2424,N_2367,N_2306);
nand U2425 (N_2425,N_2303,N_2302);
or U2426 (N_2426,N_2323,N_2316);
or U2427 (N_2427,N_2358,N_2356);
nor U2428 (N_2428,N_2332,N_2397);
and U2429 (N_2429,N_2345,N_2320);
nand U2430 (N_2430,N_2339,N_2355);
or U2431 (N_2431,N_2387,N_2310);
nand U2432 (N_2432,N_2359,N_2372);
or U2433 (N_2433,N_2309,N_2327);
or U2434 (N_2434,N_2301,N_2319);
xnor U2435 (N_2435,N_2349,N_2369);
nand U2436 (N_2436,N_2386,N_2348);
nand U2437 (N_2437,N_2322,N_2379);
nor U2438 (N_2438,N_2334,N_2325);
xnor U2439 (N_2439,N_2338,N_2354);
nand U2440 (N_2440,N_2376,N_2321);
xnor U2441 (N_2441,N_2382,N_2378);
or U2442 (N_2442,N_2344,N_2374);
nand U2443 (N_2443,N_2305,N_2329);
or U2444 (N_2444,N_2300,N_2341);
nand U2445 (N_2445,N_2360,N_2318);
nor U2446 (N_2446,N_2373,N_2394);
xor U2447 (N_2447,N_2326,N_2343);
nand U2448 (N_2448,N_2362,N_2335);
xnor U2449 (N_2449,N_2350,N_2351);
xnor U2450 (N_2450,N_2369,N_2337);
and U2451 (N_2451,N_2358,N_2311);
nand U2452 (N_2452,N_2351,N_2314);
or U2453 (N_2453,N_2344,N_2340);
xnor U2454 (N_2454,N_2336,N_2380);
xor U2455 (N_2455,N_2351,N_2333);
nor U2456 (N_2456,N_2332,N_2321);
xor U2457 (N_2457,N_2397,N_2308);
nand U2458 (N_2458,N_2307,N_2347);
xor U2459 (N_2459,N_2327,N_2384);
nand U2460 (N_2460,N_2300,N_2366);
xor U2461 (N_2461,N_2337,N_2392);
or U2462 (N_2462,N_2381,N_2390);
or U2463 (N_2463,N_2384,N_2374);
nand U2464 (N_2464,N_2397,N_2389);
and U2465 (N_2465,N_2300,N_2359);
nand U2466 (N_2466,N_2328,N_2384);
nor U2467 (N_2467,N_2369,N_2396);
or U2468 (N_2468,N_2302,N_2398);
xor U2469 (N_2469,N_2366,N_2339);
xnor U2470 (N_2470,N_2304,N_2342);
nand U2471 (N_2471,N_2337,N_2367);
and U2472 (N_2472,N_2337,N_2359);
nor U2473 (N_2473,N_2361,N_2336);
and U2474 (N_2474,N_2316,N_2343);
or U2475 (N_2475,N_2332,N_2354);
nand U2476 (N_2476,N_2383,N_2359);
xnor U2477 (N_2477,N_2311,N_2320);
or U2478 (N_2478,N_2354,N_2350);
or U2479 (N_2479,N_2392,N_2362);
nor U2480 (N_2480,N_2305,N_2335);
xor U2481 (N_2481,N_2374,N_2393);
xnor U2482 (N_2482,N_2348,N_2343);
or U2483 (N_2483,N_2353,N_2379);
nand U2484 (N_2484,N_2336,N_2305);
xor U2485 (N_2485,N_2360,N_2389);
xor U2486 (N_2486,N_2374,N_2341);
and U2487 (N_2487,N_2319,N_2347);
or U2488 (N_2488,N_2345,N_2399);
or U2489 (N_2489,N_2393,N_2362);
nand U2490 (N_2490,N_2340,N_2301);
nand U2491 (N_2491,N_2356,N_2391);
and U2492 (N_2492,N_2307,N_2304);
nand U2493 (N_2493,N_2347,N_2339);
nand U2494 (N_2494,N_2358,N_2315);
xor U2495 (N_2495,N_2311,N_2316);
and U2496 (N_2496,N_2388,N_2351);
xor U2497 (N_2497,N_2308,N_2321);
or U2498 (N_2498,N_2330,N_2346);
or U2499 (N_2499,N_2392,N_2339);
nor U2500 (N_2500,N_2458,N_2426);
and U2501 (N_2501,N_2479,N_2484);
or U2502 (N_2502,N_2407,N_2434);
and U2503 (N_2503,N_2419,N_2432);
nand U2504 (N_2504,N_2411,N_2442);
nand U2505 (N_2505,N_2487,N_2404);
xor U2506 (N_2506,N_2460,N_2449);
nor U2507 (N_2507,N_2451,N_2455);
nor U2508 (N_2508,N_2429,N_2463);
nand U2509 (N_2509,N_2415,N_2457);
nor U2510 (N_2510,N_2464,N_2441);
xor U2511 (N_2511,N_2435,N_2436);
or U2512 (N_2512,N_2433,N_2444);
and U2513 (N_2513,N_2405,N_2412);
and U2514 (N_2514,N_2440,N_2480);
xor U2515 (N_2515,N_2478,N_2438);
xor U2516 (N_2516,N_2421,N_2437);
nor U2517 (N_2517,N_2443,N_2494);
or U2518 (N_2518,N_2454,N_2400);
nand U2519 (N_2519,N_2485,N_2450);
nor U2520 (N_2520,N_2486,N_2467);
or U2521 (N_2521,N_2420,N_2496);
and U2522 (N_2522,N_2498,N_2414);
xnor U2523 (N_2523,N_2491,N_2427);
or U2524 (N_2524,N_2459,N_2481);
and U2525 (N_2525,N_2416,N_2413);
nor U2526 (N_2526,N_2406,N_2482);
nand U2527 (N_2527,N_2483,N_2488);
xnor U2528 (N_2528,N_2428,N_2453);
xor U2529 (N_2529,N_2477,N_2476);
and U2530 (N_2530,N_2410,N_2446);
xnor U2531 (N_2531,N_2469,N_2462);
nor U2532 (N_2532,N_2489,N_2445);
and U2533 (N_2533,N_2499,N_2422);
nor U2534 (N_2534,N_2475,N_2465);
and U2535 (N_2535,N_2495,N_2409);
nor U2536 (N_2536,N_2473,N_2490);
or U2537 (N_2537,N_2448,N_2468);
or U2538 (N_2538,N_2403,N_2417);
xnor U2539 (N_2539,N_2466,N_2439);
nand U2540 (N_2540,N_2408,N_2493);
or U2541 (N_2541,N_2447,N_2423);
nor U2542 (N_2542,N_2472,N_2425);
and U2543 (N_2543,N_2492,N_2461);
or U2544 (N_2544,N_2474,N_2452);
or U2545 (N_2545,N_2471,N_2418);
xnor U2546 (N_2546,N_2430,N_2431);
nand U2547 (N_2547,N_2401,N_2402);
nand U2548 (N_2548,N_2470,N_2497);
or U2549 (N_2549,N_2424,N_2456);
xnor U2550 (N_2550,N_2492,N_2463);
nor U2551 (N_2551,N_2468,N_2457);
nand U2552 (N_2552,N_2493,N_2499);
and U2553 (N_2553,N_2450,N_2486);
nand U2554 (N_2554,N_2439,N_2441);
nand U2555 (N_2555,N_2443,N_2481);
and U2556 (N_2556,N_2440,N_2494);
and U2557 (N_2557,N_2433,N_2495);
or U2558 (N_2558,N_2492,N_2443);
nor U2559 (N_2559,N_2411,N_2414);
nand U2560 (N_2560,N_2428,N_2465);
nand U2561 (N_2561,N_2484,N_2458);
and U2562 (N_2562,N_2412,N_2403);
nor U2563 (N_2563,N_2407,N_2483);
or U2564 (N_2564,N_2401,N_2407);
and U2565 (N_2565,N_2471,N_2459);
and U2566 (N_2566,N_2426,N_2463);
nand U2567 (N_2567,N_2494,N_2490);
nand U2568 (N_2568,N_2460,N_2481);
nand U2569 (N_2569,N_2456,N_2425);
xnor U2570 (N_2570,N_2483,N_2474);
and U2571 (N_2571,N_2437,N_2483);
nor U2572 (N_2572,N_2451,N_2402);
nand U2573 (N_2573,N_2408,N_2447);
nor U2574 (N_2574,N_2478,N_2489);
xnor U2575 (N_2575,N_2457,N_2431);
nand U2576 (N_2576,N_2472,N_2470);
and U2577 (N_2577,N_2435,N_2469);
nor U2578 (N_2578,N_2460,N_2443);
and U2579 (N_2579,N_2460,N_2492);
and U2580 (N_2580,N_2417,N_2430);
nand U2581 (N_2581,N_2402,N_2422);
nor U2582 (N_2582,N_2481,N_2420);
or U2583 (N_2583,N_2446,N_2424);
or U2584 (N_2584,N_2452,N_2428);
and U2585 (N_2585,N_2486,N_2485);
or U2586 (N_2586,N_2433,N_2430);
nor U2587 (N_2587,N_2443,N_2418);
and U2588 (N_2588,N_2475,N_2447);
or U2589 (N_2589,N_2463,N_2478);
nor U2590 (N_2590,N_2422,N_2465);
and U2591 (N_2591,N_2486,N_2471);
and U2592 (N_2592,N_2419,N_2438);
and U2593 (N_2593,N_2490,N_2433);
xor U2594 (N_2594,N_2445,N_2466);
nor U2595 (N_2595,N_2464,N_2425);
nand U2596 (N_2596,N_2474,N_2438);
or U2597 (N_2597,N_2425,N_2462);
xnor U2598 (N_2598,N_2425,N_2410);
nand U2599 (N_2599,N_2439,N_2461);
and U2600 (N_2600,N_2507,N_2589);
xor U2601 (N_2601,N_2524,N_2503);
nand U2602 (N_2602,N_2518,N_2555);
nand U2603 (N_2603,N_2558,N_2597);
nor U2604 (N_2604,N_2541,N_2585);
or U2605 (N_2605,N_2530,N_2568);
xor U2606 (N_2606,N_2560,N_2514);
nand U2607 (N_2607,N_2502,N_2557);
or U2608 (N_2608,N_2535,N_2519);
nor U2609 (N_2609,N_2515,N_2588);
or U2610 (N_2610,N_2505,N_2581);
xor U2611 (N_2611,N_2594,N_2550);
nor U2612 (N_2612,N_2595,N_2587);
and U2613 (N_2613,N_2592,N_2582);
nand U2614 (N_2614,N_2596,N_2538);
xnor U2615 (N_2615,N_2561,N_2525);
nor U2616 (N_2616,N_2500,N_2573);
nand U2617 (N_2617,N_2553,N_2556);
or U2618 (N_2618,N_2508,N_2565);
xor U2619 (N_2619,N_2572,N_2574);
or U2620 (N_2620,N_2540,N_2523);
and U2621 (N_2621,N_2569,N_2528);
nor U2622 (N_2622,N_2520,N_2593);
or U2623 (N_2623,N_2577,N_2562);
xnor U2624 (N_2624,N_2575,N_2578);
nand U2625 (N_2625,N_2504,N_2563);
nor U2626 (N_2626,N_2580,N_2571);
xor U2627 (N_2627,N_2510,N_2546);
and U2628 (N_2628,N_2544,N_2533);
xor U2629 (N_2629,N_2517,N_2511);
nand U2630 (N_2630,N_2584,N_2586);
xnor U2631 (N_2631,N_2512,N_2590);
xor U2632 (N_2632,N_2527,N_2516);
xor U2633 (N_2633,N_2531,N_2547);
or U2634 (N_2634,N_2552,N_2551);
nor U2635 (N_2635,N_2522,N_2513);
or U2636 (N_2636,N_2576,N_2549);
nor U2637 (N_2637,N_2566,N_2567);
and U2638 (N_2638,N_2545,N_2598);
nor U2639 (N_2639,N_2559,N_2542);
nor U2640 (N_2640,N_2536,N_2501);
xnor U2641 (N_2641,N_2506,N_2570);
nand U2642 (N_2642,N_2543,N_2532);
xnor U2643 (N_2643,N_2599,N_2554);
and U2644 (N_2644,N_2509,N_2548);
xnor U2645 (N_2645,N_2526,N_2521);
xor U2646 (N_2646,N_2539,N_2579);
and U2647 (N_2647,N_2591,N_2529);
or U2648 (N_2648,N_2564,N_2583);
and U2649 (N_2649,N_2534,N_2537);
xnor U2650 (N_2650,N_2555,N_2599);
nand U2651 (N_2651,N_2507,N_2524);
and U2652 (N_2652,N_2596,N_2593);
or U2653 (N_2653,N_2522,N_2579);
or U2654 (N_2654,N_2537,N_2531);
or U2655 (N_2655,N_2562,N_2512);
xor U2656 (N_2656,N_2527,N_2525);
and U2657 (N_2657,N_2527,N_2582);
or U2658 (N_2658,N_2539,N_2562);
nand U2659 (N_2659,N_2558,N_2574);
xor U2660 (N_2660,N_2529,N_2547);
or U2661 (N_2661,N_2579,N_2572);
nand U2662 (N_2662,N_2599,N_2516);
nand U2663 (N_2663,N_2552,N_2544);
nand U2664 (N_2664,N_2565,N_2583);
and U2665 (N_2665,N_2510,N_2539);
xor U2666 (N_2666,N_2511,N_2554);
xnor U2667 (N_2667,N_2578,N_2509);
and U2668 (N_2668,N_2557,N_2599);
nor U2669 (N_2669,N_2586,N_2599);
xor U2670 (N_2670,N_2527,N_2502);
xor U2671 (N_2671,N_2523,N_2552);
and U2672 (N_2672,N_2586,N_2582);
and U2673 (N_2673,N_2543,N_2597);
and U2674 (N_2674,N_2554,N_2523);
nor U2675 (N_2675,N_2598,N_2523);
or U2676 (N_2676,N_2578,N_2552);
nor U2677 (N_2677,N_2505,N_2525);
nand U2678 (N_2678,N_2588,N_2596);
nor U2679 (N_2679,N_2502,N_2588);
nand U2680 (N_2680,N_2502,N_2563);
xnor U2681 (N_2681,N_2539,N_2538);
or U2682 (N_2682,N_2530,N_2548);
or U2683 (N_2683,N_2580,N_2509);
nand U2684 (N_2684,N_2546,N_2538);
nor U2685 (N_2685,N_2583,N_2555);
xnor U2686 (N_2686,N_2513,N_2510);
and U2687 (N_2687,N_2550,N_2582);
and U2688 (N_2688,N_2594,N_2584);
nand U2689 (N_2689,N_2555,N_2531);
xor U2690 (N_2690,N_2565,N_2535);
nand U2691 (N_2691,N_2572,N_2510);
xnor U2692 (N_2692,N_2508,N_2582);
and U2693 (N_2693,N_2567,N_2592);
nor U2694 (N_2694,N_2580,N_2506);
nand U2695 (N_2695,N_2594,N_2542);
xnor U2696 (N_2696,N_2595,N_2570);
nor U2697 (N_2697,N_2545,N_2591);
xnor U2698 (N_2698,N_2507,N_2575);
nor U2699 (N_2699,N_2559,N_2576);
nor U2700 (N_2700,N_2669,N_2644);
nor U2701 (N_2701,N_2670,N_2681);
or U2702 (N_2702,N_2609,N_2652);
nor U2703 (N_2703,N_2640,N_2699);
nand U2704 (N_2704,N_2665,N_2666);
nand U2705 (N_2705,N_2602,N_2632);
and U2706 (N_2706,N_2680,N_2610);
xnor U2707 (N_2707,N_2635,N_2653);
or U2708 (N_2708,N_2657,N_2673);
xor U2709 (N_2709,N_2676,N_2611);
nand U2710 (N_2710,N_2604,N_2636);
nor U2711 (N_2711,N_2619,N_2674);
nor U2712 (N_2712,N_2698,N_2690);
or U2713 (N_2713,N_2623,N_2683);
and U2714 (N_2714,N_2693,N_2664);
nor U2715 (N_2715,N_2638,N_2615);
nand U2716 (N_2716,N_2684,N_2662);
nand U2717 (N_2717,N_2601,N_2645);
xnor U2718 (N_2718,N_2672,N_2647);
nand U2719 (N_2719,N_2663,N_2634);
or U2720 (N_2720,N_2646,N_2648);
xnor U2721 (N_2721,N_2633,N_2651);
and U2722 (N_2722,N_2618,N_2629);
and U2723 (N_2723,N_2656,N_2671);
xnor U2724 (N_2724,N_2682,N_2622);
and U2725 (N_2725,N_2649,N_2603);
or U2726 (N_2726,N_2675,N_2607);
or U2727 (N_2727,N_2642,N_2668);
and U2728 (N_2728,N_2621,N_2659);
or U2729 (N_2729,N_2612,N_2620);
nor U2730 (N_2730,N_2605,N_2696);
nand U2731 (N_2731,N_2661,N_2626);
and U2732 (N_2732,N_2625,N_2685);
xor U2733 (N_2733,N_2697,N_2658);
nor U2734 (N_2734,N_2654,N_2643);
and U2735 (N_2735,N_2616,N_2677);
nor U2736 (N_2736,N_2655,N_2627);
nor U2737 (N_2737,N_2687,N_2679);
nor U2738 (N_2738,N_2606,N_2691);
or U2739 (N_2739,N_2650,N_2686);
nor U2740 (N_2740,N_2600,N_2639);
xor U2741 (N_2741,N_2667,N_2689);
and U2742 (N_2742,N_2613,N_2692);
and U2743 (N_2743,N_2614,N_2630);
and U2744 (N_2744,N_2695,N_2637);
nor U2745 (N_2745,N_2628,N_2631);
or U2746 (N_2746,N_2688,N_2694);
or U2747 (N_2747,N_2641,N_2624);
and U2748 (N_2748,N_2617,N_2660);
nor U2749 (N_2749,N_2608,N_2678);
nor U2750 (N_2750,N_2667,N_2632);
xnor U2751 (N_2751,N_2625,N_2657);
nor U2752 (N_2752,N_2605,N_2658);
nor U2753 (N_2753,N_2662,N_2620);
nand U2754 (N_2754,N_2619,N_2658);
xnor U2755 (N_2755,N_2653,N_2629);
nor U2756 (N_2756,N_2695,N_2648);
nor U2757 (N_2757,N_2634,N_2654);
or U2758 (N_2758,N_2684,N_2650);
xnor U2759 (N_2759,N_2659,N_2671);
nand U2760 (N_2760,N_2680,N_2673);
xor U2761 (N_2761,N_2691,N_2640);
xor U2762 (N_2762,N_2665,N_2603);
xor U2763 (N_2763,N_2640,N_2608);
xnor U2764 (N_2764,N_2610,N_2627);
or U2765 (N_2765,N_2627,N_2680);
and U2766 (N_2766,N_2638,N_2600);
nand U2767 (N_2767,N_2657,N_2612);
xor U2768 (N_2768,N_2678,N_2639);
and U2769 (N_2769,N_2688,N_2652);
nand U2770 (N_2770,N_2665,N_2659);
and U2771 (N_2771,N_2616,N_2692);
nand U2772 (N_2772,N_2682,N_2600);
xnor U2773 (N_2773,N_2628,N_2642);
nor U2774 (N_2774,N_2605,N_2606);
nor U2775 (N_2775,N_2673,N_2602);
and U2776 (N_2776,N_2669,N_2640);
xor U2777 (N_2777,N_2647,N_2637);
nor U2778 (N_2778,N_2635,N_2647);
xnor U2779 (N_2779,N_2641,N_2633);
xor U2780 (N_2780,N_2688,N_2617);
or U2781 (N_2781,N_2650,N_2609);
nand U2782 (N_2782,N_2615,N_2617);
and U2783 (N_2783,N_2643,N_2640);
nor U2784 (N_2784,N_2690,N_2637);
nand U2785 (N_2785,N_2691,N_2674);
nor U2786 (N_2786,N_2673,N_2660);
and U2787 (N_2787,N_2626,N_2635);
nand U2788 (N_2788,N_2639,N_2693);
nor U2789 (N_2789,N_2619,N_2608);
and U2790 (N_2790,N_2605,N_2698);
nor U2791 (N_2791,N_2686,N_2697);
xor U2792 (N_2792,N_2625,N_2607);
or U2793 (N_2793,N_2611,N_2650);
xor U2794 (N_2794,N_2658,N_2680);
nor U2795 (N_2795,N_2659,N_2607);
nand U2796 (N_2796,N_2635,N_2661);
nand U2797 (N_2797,N_2638,N_2659);
nand U2798 (N_2798,N_2609,N_2690);
xnor U2799 (N_2799,N_2617,N_2657);
nand U2800 (N_2800,N_2772,N_2741);
nand U2801 (N_2801,N_2742,N_2799);
and U2802 (N_2802,N_2703,N_2739);
xnor U2803 (N_2803,N_2736,N_2782);
and U2804 (N_2804,N_2719,N_2740);
and U2805 (N_2805,N_2788,N_2709);
or U2806 (N_2806,N_2781,N_2754);
and U2807 (N_2807,N_2744,N_2718);
nor U2808 (N_2808,N_2777,N_2701);
nor U2809 (N_2809,N_2785,N_2756);
nand U2810 (N_2810,N_2751,N_2729);
nor U2811 (N_2811,N_2796,N_2791);
xnor U2812 (N_2812,N_2766,N_2767);
nand U2813 (N_2813,N_2717,N_2727);
and U2814 (N_2814,N_2708,N_2774);
nor U2815 (N_2815,N_2790,N_2735);
and U2816 (N_2816,N_2761,N_2780);
xnor U2817 (N_2817,N_2792,N_2764);
xor U2818 (N_2818,N_2789,N_2795);
xor U2819 (N_2819,N_2702,N_2787);
xor U2820 (N_2820,N_2720,N_2738);
xnor U2821 (N_2821,N_2752,N_2714);
and U2822 (N_2822,N_2749,N_2730);
nor U2823 (N_2823,N_2723,N_2783);
nand U2824 (N_2824,N_2710,N_2728);
nor U2825 (N_2825,N_2768,N_2784);
or U2826 (N_2826,N_2748,N_2725);
nor U2827 (N_2827,N_2705,N_2737);
and U2828 (N_2828,N_2704,N_2773);
or U2829 (N_2829,N_2707,N_2712);
nand U2830 (N_2830,N_2721,N_2731);
or U2831 (N_2831,N_2778,N_2793);
nand U2832 (N_2832,N_2753,N_2760);
nor U2833 (N_2833,N_2798,N_2716);
xor U2834 (N_2834,N_2779,N_2769);
xnor U2835 (N_2835,N_2762,N_2755);
xor U2836 (N_2836,N_2786,N_2763);
nand U2837 (N_2837,N_2771,N_2757);
nand U2838 (N_2838,N_2794,N_2711);
nand U2839 (N_2839,N_2732,N_2734);
nand U2840 (N_2840,N_2797,N_2765);
xnor U2841 (N_2841,N_2746,N_2713);
xor U2842 (N_2842,N_2733,N_2700);
or U2843 (N_2843,N_2706,N_2722);
nor U2844 (N_2844,N_2726,N_2770);
nand U2845 (N_2845,N_2743,N_2747);
and U2846 (N_2846,N_2715,N_2775);
or U2847 (N_2847,N_2759,N_2750);
or U2848 (N_2848,N_2724,N_2745);
nor U2849 (N_2849,N_2758,N_2776);
nor U2850 (N_2850,N_2717,N_2707);
and U2851 (N_2851,N_2762,N_2757);
nor U2852 (N_2852,N_2714,N_2756);
or U2853 (N_2853,N_2738,N_2767);
and U2854 (N_2854,N_2724,N_2742);
xor U2855 (N_2855,N_2724,N_2761);
nand U2856 (N_2856,N_2786,N_2731);
nor U2857 (N_2857,N_2762,N_2785);
or U2858 (N_2858,N_2732,N_2730);
nand U2859 (N_2859,N_2771,N_2776);
and U2860 (N_2860,N_2700,N_2701);
nand U2861 (N_2861,N_2753,N_2778);
and U2862 (N_2862,N_2708,N_2713);
nand U2863 (N_2863,N_2766,N_2727);
or U2864 (N_2864,N_2762,N_2704);
nor U2865 (N_2865,N_2737,N_2748);
and U2866 (N_2866,N_2701,N_2730);
xnor U2867 (N_2867,N_2782,N_2757);
xnor U2868 (N_2868,N_2707,N_2710);
xor U2869 (N_2869,N_2794,N_2738);
and U2870 (N_2870,N_2734,N_2784);
or U2871 (N_2871,N_2747,N_2764);
and U2872 (N_2872,N_2771,N_2714);
xor U2873 (N_2873,N_2746,N_2769);
nor U2874 (N_2874,N_2716,N_2776);
nor U2875 (N_2875,N_2729,N_2739);
or U2876 (N_2876,N_2705,N_2720);
xor U2877 (N_2877,N_2793,N_2709);
and U2878 (N_2878,N_2746,N_2717);
and U2879 (N_2879,N_2782,N_2774);
xnor U2880 (N_2880,N_2787,N_2741);
nand U2881 (N_2881,N_2798,N_2763);
and U2882 (N_2882,N_2788,N_2713);
xnor U2883 (N_2883,N_2733,N_2716);
xor U2884 (N_2884,N_2769,N_2749);
or U2885 (N_2885,N_2750,N_2712);
xnor U2886 (N_2886,N_2761,N_2751);
xor U2887 (N_2887,N_2743,N_2786);
nand U2888 (N_2888,N_2771,N_2797);
nor U2889 (N_2889,N_2798,N_2718);
nand U2890 (N_2890,N_2789,N_2702);
nor U2891 (N_2891,N_2776,N_2757);
nor U2892 (N_2892,N_2796,N_2715);
and U2893 (N_2893,N_2768,N_2723);
or U2894 (N_2894,N_2758,N_2704);
nor U2895 (N_2895,N_2710,N_2704);
and U2896 (N_2896,N_2748,N_2707);
nor U2897 (N_2897,N_2729,N_2790);
or U2898 (N_2898,N_2716,N_2709);
or U2899 (N_2899,N_2787,N_2735);
xnor U2900 (N_2900,N_2879,N_2809);
or U2901 (N_2901,N_2840,N_2830);
and U2902 (N_2902,N_2864,N_2842);
nand U2903 (N_2903,N_2825,N_2841);
or U2904 (N_2904,N_2800,N_2818);
nor U2905 (N_2905,N_2860,N_2897);
or U2906 (N_2906,N_2857,N_2806);
or U2907 (N_2907,N_2812,N_2894);
nor U2908 (N_2908,N_2861,N_2835);
nor U2909 (N_2909,N_2878,N_2808);
nor U2910 (N_2910,N_2850,N_2834);
xnor U2911 (N_2911,N_2868,N_2844);
or U2912 (N_2912,N_2828,N_2846);
xor U2913 (N_2913,N_2807,N_2851);
nor U2914 (N_2914,N_2875,N_2876);
nand U2915 (N_2915,N_2881,N_2867);
or U2916 (N_2916,N_2896,N_2874);
xnor U2917 (N_2917,N_2827,N_2866);
and U2918 (N_2918,N_2898,N_2892);
nor U2919 (N_2919,N_2805,N_2877);
xnor U2920 (N_2920,N_2816,N_2829);
or U2921 (N_2921,N_2813,N_2859);
and U2922 (N_2922,N_2801,N_2847);
nand U2923 (N_2923,N_2882,N_2855);
nand U2924 (N_2924,N_2802,N_2863);
xnor U2925 (N_2925,N_2887,N_2843);
nand U2926 (N_2926,N_2853,N_2837);
xnor U2927 (N_2927,N_2821,N_2854);
and U2928 (N_2928,N_2889,N_2849);
and U2929 (N_2929,N_2862,N_2852);
nor U2930 (N_2930,N_2858,N_2869);
nand U2931 (N_2931,N_2885,N_2890);
nor U2932 (N_2932,N_2865,N_2833);
xnor U2933 (N_2933,N_2819,N_2826);
xor U2934 (N_2934,N_2880,N_2831);
or U2935 (N_2935,N_2870,N_2820);
or U2936 (N_2936,N_2803,N_2872);
nand U2937 (N_2937,N_2871,N_2836);
xnor U2938 (N_2938,N_2845,N_2848);
nand U2939 (N_2939,N_2815,N_2883);
nand U2940 (N_2940,N_2817,N_2811);
and U2941 (N_2941,N_2873,N_2888);
nor U2942 (N_2942,N_2838,N_2824);
nor U2943 (N_2943,N_2810,N_2891);
nor U2944 (N_2944,N_2804,N_2886);
or U2945 (N_2945,N_2832,N_2823);
or U2946 (N_2946,N_2856,N_2814);
nor U2947 (N_2947,N_2895,N_2822);
xor U2948 (N_2948,N_2899,N_2839);
or U2949 (N_2949,N_2893,N_2884);
xnor U2950 (N_2950,N_2811,N_2841);
nand U2951 (N_2951,N_2879,N_2885);
nand U2952 (N_2952,N_2868,N_2864);
or U2953 (N_2953,N_2802,N_2884);
or U2954 (N_2954,N_2890,N_2813);
xnor U2955 (N_2955,N_2890,N_2875);
nand U2956 (N_2956,N_2886,N_2806);
xnor U2957 (N_2957,N_2800,N_2824);
xor U2958 (N_2958,N_2895,N_2827);
and U2959 (N_2959,N_2878,N_2845);
and U2960 (N_2960,N_2832,N_2811);
or U2961 (N_2961,N_2886,N_2882);
or U2962 (N_2962,N_2843,N_2837);
nor U2963 (N_2963,N_2813,N_2894);
and U2964 (N_2964,N_2849,N_2804);
or U2965 (N_2965,N_2885,N_2827);
nand U2966 (N_2966,N_2860,N_2800);
nor U2967 (N_2967,N_2801,N_2813);
and U2968 (N_2968,N_2836,N_2837);
xor U2969 (N_2969,N_2851,N_2865);
or U2970 (N_2970,N_2861,N_2852);
nor U2971 (N_2971,N_2863,N_2842);
and U2972 (N_2972,N_2862,N_2810);
xnor U2973 (N_2973,N_2827,N_2878);
nand U2974 (N_2974,N_2882,N_2811);
nand U2975 (N_2975,N_2882,N_2877);
and U2976 (N_2976,N_2824,N_2859);
nor U2977 (N_2977,N_2828,N_2837);
or U2978 (N_2978,N_2852,N_2894);
and U2979 (N_2979,N_2811,N_2881);
or U2980 (N_2980,N_2868,N_2805);
or U2981 (N_2981,N_2887,N_2815);
xor U2982 (N_2982,N_2842,N_2849);
and U2983 (N_2983,N_2820,N_2882);
or U2984 (N_2984,N_2839,N_2863);
or U2985 (N_2985,N_2849,N_2877);
nor U2986 (N_2986,N_2834,N_2826);
xnor U2987 (N_2987,N_2848,N_2844);
nand U2988 (N_2988,N_2835,N_2826);
nor U2989 (N_2989,N_2864,N_2897);
and U2990 (N_2990,N_2854,N_2814);
or U2991 (N_2991,N_2806,N_2809);
xor U2992 (N_2992,N_2864,N_2865);
or U2993 (N_2993,N_2864,N_2844);
and U2994 (N_2994,N_2800,N_2803);
xnor U2995 (N_2995,N_2836,N_2816);
nand U2996 (N_2996,N_2891,N_2836);
xor U2997 (N_2997,N_2815,N_2821);
and U2998 (N_2998,N_2891,N_2872);
xnor U2999 (N_2999,N_2828,N_2801);
nor UO_0 (O_0,N_2901,N_2929);
or UO_1 (O_1,N_2970,N_2982);
or UO_2 (O_2,N_2930,N_2903);
or UO_3 (O_3,N_2915,N_2977);
xor UO_4 (O_4,N_2900,N_2980);
nor UO_5 (O_5,N_2908,N_2922);
or UO_6 (O_6,N_2979,N_2939);
nor UO_7 (O_7,N_2952,N_2988);
and UO_8 (O_8,N_2953,N_2945);
nand UO_9 (O_9,N_2917,N_2976);
or UO_10 (O_10,N_2916,N_2919);
nor UO_11 (O_11,N_2950,N_2968);
and UO_12 (O_12,N_2963,N_2960);
or UO_13 (O_13,N_2906,N_2990);
and UO_14 (O_14,N_2937,N_2994);
or UO_15 (O_15,N_2947,N_2924);
or UO_16 (O_16,N_2902,N_2956);
xnor UO_17 (O_17,N_2920,N_2997);
or UO_18 (O_18,N_2983,N_2949);
xor UO_19 (O_19,N_2989,N_2911);
and UO_20 (O_20,N_2992,N_2943);
xor UO_21 (O_21,N_2964,N_2966);
nand UO_22 (O_22,N_2936,N_2923);
nor UO_23 (O_23,N_2985,N_2995);
and UO_24 (O_24,N_2996,N_2907);
nand UO_25 (O_25,N_2972,N_2913);
nor UO_26 (O_26,N_2957,N_2932);
or UO_27 (O_27,N_2986,N_2971);
or UO_28 (O_28,N_2905,N_2933);
nor UO_29 (O_29,N_2991,N_2987);
nand UO_30 (O_30,N_2904,N_2969);
or UO_31 (O_31,N_2993,N_2984);
nand UO_32 (O_32,N_2958,N_2926);
xor UO_33 (O_33,N_2914,N_2981);
or UO_34 (O_34,N_2931,N_2962);
and UO_35 (O_35,N_2918,N_2925);
xor UO_36 (O_36,N_2909,N_2978);
xnor UO_37 (O_37,N_2973,N_2938);
xnor UO_38 (O_38,N_2934,N_2999);
or UO_39 (O_39,N_2944,N_2961);
nor UO_40 (O_40,N_2959,N_2941);
and UO_41 (O_41,N_2954,N_2912);
xor UO_42 (O_42,N_2927,N_2928);
xnor UO_43 (O_43,N_2948,N_2946);
nand UO_44 (O_44,N_2942,N_2921);
nor UO_45 (O_45,N_2974,N_2955);
or UO_46 (O_46,N_2975,N_2967);
or UO_47 (O_47,N_2935,N_2910);
xor UO_48 (O_48,N_2951,N_2998);
nor UO_49 (O_49,N_2940,N_2965);
nand UO_50 (O_50,N_2988,N_2968);
nor UO_51 (O_51,N_2961,N_2919);
and UO_52 (O_52,N_2912,N_2904);
nor UO_53 (O_53,N_2989,N_2979);
xnor UO_54 (O_54,N_2911,N_2914);
and UO_55 (O_55,N_2926,N_2963);
nor UO_56 (O_56,N_2970,N_2934);
nor UO_57 (O_57,N_2946,N_2990);
and UO_58 (O_58,N_2957,N_2907);
and UO_59 (O_59,N_2919,N_2936);
or UO_60 (O_60,N_2979,N_2909);
or UO_61 (O_61,N_2971,N_2951);
nor UO_62 (O_62,N_2942,N_2974);
nand UO_63 (O_63,N_2924,N_2952);
nor UO_64 (O_64,N_2955,N_2981);
xor UO_65 (O_65,N_2937,N_2940);
or UO_66 (O_66,N_2961,N_2939);
nand UO_67 (O_67,N_2954,N_2995);
nand UO_68 (O_68,N_2997,N_2905);
nand UO_69 (O_69,N_2927,N_2993);
nor UO_70 (O_70,N_2915,N_2911);
nor UO_71 (O_71,N_2987,N_2972);
nand UO_72 (O_72,N_2907,N_2915);
and UO_73 (O_73,N_2921,N_2903);
xnor UO_74 (O_74,N_2906,N_2994);
or UO_75 (O_75,N_2995,N_2981);
xor UO_76 (O_76,N_2948,N_2938);
xor UO_77 (O_77,N_2915,N_2925);
nor UO_78 (O_78,N_2916,N_2936);
or UO_79 (O_79,N_2935,N_2945);
xnor UO_80 (O_80,N_2937,N_2991);
and UO_81 (O_81,N_2940,N_2949);
and UO_82 (O_82,N_2976,N_2951);
xnor UO_83 (O_83,N_2949,N_2932);
nor UO_84 (O_84,N_2976,N_2948);
nand UO_85 (O_85,N_2968,N_2939);
xnor UO_86 (O_86,N_2989,N_2941);
nor UO_87 (O_87,N_2978,N_2913);
nor UO_88 (O_88,N_2947,N_2922);
xnor UO_89 (O_89,N_2913,N_2982);
and UO_90 (O_90,N_2909,N_2913);
nor UO_91 (O_91,N_2958,N_2967);
xnor UO_92 (O_92,N_2910,N_2973);
and UO_93 (O_93,N_2915,N_2951);
or UO_94 (O_94,N_2979,N_2941);
nand UO_95 (O_95,N_2956,N_2960);
and UO_96 (O_96,N_2905,N_2906);
nor UO_97 (O_97,N_2954,N_2952);
xnor UO_98 (O_98,N_2953,N_2984);
xor UO_99 (O_99,N_2960,N_2906);
or UO_100 (O_100,N_2963,N_2944);
nand UO_101 (O_101,N_2945,N_2960);
and UO_102 (O_102,N_2938,N_2979);
nand UO_103 (O_103,N_2930,N_2902);
nand UO_104 (O_104,N_2907,N_2930);
nand UO_105 (O_105,N_2980,N_2976);
xor UO_106 (O_106,N_2912,N_2930);
xnor UO_107 (O_107,N_2954,N_2977);
xor UO_108 (O_108,N_2951,N_2987);
or UO_109 (O_109,N_2907,N_2954);
and UO_110 (O_110,N_2940,N_2950);
nand UO_111 (O_111,N_2972,N_2969);
nor UO_112 (O_112,N_2972,N_2959);
xor UO_113 (O_113,N_2979,N_2919);
nand UO_114 (O_114,N_2936,N_2997);
and UO_115 (O_115,N_2916,N_2996);
nor UO_116 (O_116,N_2920,N_2980);
nor UO_117 (O_117,N_2989,N_2964);
xor UO_118 (O_118,N_2904,N_2999);
nor UO_119 (O_119,N_2921,N_2938);
or UO_120 (O_120,N_2971,N_2998);
xor UO_121 (O_121,N_2938,N_2911);
nor UO_122 (O_122,N_2960,N_2938);
nand UO_123 (O_123,N_2988,N_2984);
and UO_124 (O_124,N_2922,N_2959);
xnor UO_125 (O_125,N_2919,N_2951);
nor UO_126 (O_126,N_2910,N_2998);
xor UO_127 (O_127,N_2956,N_2920);
and UO_128 (O_128,N_2962,N_2964);
and UO_129 (O_129,N_2916,N_2912);
nand UO_130 (O_130,N_2937,N_2946);
or UO_131 (O_131,N_2905,N_2955);
and UO_132 (O_132,N_2972,N_2934);
nand UO_133 (O_133,N_2939,N_2957);
nand UO_134 (O_134,N_2954,N_2931);
xor UO_135 (O_135,N_2973,N_2952);
or UO_136 (O_136,N_2905,N_2953);
nor UO_137 (O_137,N_2951,N_2967);
nor UO_138 (O_138,N_2914,N_2909);
xor UO_139 (O_139,N_2956,N_2973);
and UO_140 (O_140,N_2976,N_2966);
or UO_141 (O_141,N_2944,N_2968);
nor UO_142 (O_142,N_2919,N_2928);
and UO_143 (O_143,N_2934,N_2909);
xnor UO_144 (O_144,N_2919,N_2912);
xnor UO_145 (O_145,N_2926,N_2909);
nand UO_146 (O_146,N_2947,N_2979);
and UO_147 (O_147,N_2914,N_2903);
nor UO_148 (O_148,N_2909,N_2975);
and UO_149 (O_149,N_2943,N_2977);
and UO_150 (O_150,N_2946,N_2993);
xnor UO_151 (O_151,N_2998,N_2960);
or UO_152 (O_152,N_2963,N_2920);
nand UO_153 (O_153,N_2979,N_2932);
xor UO_154 (O_154,N_2920,N_2911);
xnor UO_155 (O_155,N_2959,N_2988);
nand UO_156 (O_156,N_2937,N_2919);
and UO_157 (O_157,N_2939,N_2919);
xnor UO_158 (O_158,N_2951,N_2955);
xor UO_159 (O_159,N_2914,N_2975);
nand UO_160 (O_160,N_2962,N_2976);
or UO_161 (O_161,N_2970,N_2902);
nor UO_162 (O_162,N_2978,N_2905);
and UO_163 (O_163,N_2976,N_2963);
nor UO_164 (O_164,N_2905,N_2995);
or UO_165 (O_165,N_2931,N_2941);
nor UO_166 (O_166,N_2997,N_2934);
nand UO_167 (O_167,N_2936,N_2906);
and UO_168 (O_168,N_2973,N_2925);
nand UO_169 (O_169,N_2943,N_2985);
and UO_170 (O_170,N_2981,N_2983);
or UO_171 (O_171,N_2961,N_2960);
and UO_172 (O_172,N_2978,N_2986);
nor UO_173 (O_173,N_2988,N_2992);
or UO_174 (O_174,N_2918,N_2929);
nor UO_175 (O_175,N_2950,N_2917);
or UO_176 (O_176,N_2954,N_2936);
nand UO_177 (O_177,N_2920,N_2957);
and UO_178 (O_178,N_2971,N_2919);
nor UO_179 (O_179,N_2911,N_2993);
xnor UO_180 (O_180,N_2937,N_2902);
or UO_181 (O_181,N_2907,N_2919);
nor UO_182 (O_182,N_2991,N_2965);
or UO_183 (O_183,N_2917,N_2984);
nor UO_184 (O_184,N_2976,N_2974);
xor UO_185 (O_185,N_2957,N_2966);
xnor UO_186 (O_186,N_2987,N_2934);
and UO_187 (O_187,N_2942,N_2995);
or UO_188 (O_188,N_2970,N_2956);
and UO_189 (O_189,N_2905,N_2941);
and UO_190 (O_190,N_2929,N_2998);
nor UO_191 (O_191,N_2927,N_2906);
or UO_192 (O_192,N_2964,N_2913);
and UO_193 (O_193,N_2994,N_2929);
xor UO_194 (O_194,N_2919,N_2922);
nand UO_195 (O_195,N_2922,N_2979);
and UO_196 (O_196,N_2981,N_2952);
xnor UO_197 (O_197,N_2932,N_2947);
xnor UO_198 (O_198,N_2944,N_2919);
nor UO_199 (O_199,N_2927,N_2901);
nor UO_200 (O_200,N_2934,N_2945);
and UO_201 (O_201,N_2917,N_2942);
nand UO_202 (O_202,N_2942,N_2980);
nor UO_203 (O_203,N_2975,N_2978);
xnor UO_204 (O_204,N_2960,N_2902);
and UO_205 (O_205,N_2907,N_2992);
nor UO_206 (O_206,N_2926,N_2947);
and UO_207 (O_207,N_2955,N_2925);
nand UO_208 (O_208,N_2971,N_2903);
nor UO_209 (O_209,N_2906,N_2973);
and UO_210 (O_210,N_2937,N_2969);
nor UO_211 (O_211,N_2986,N_2967);
nand UO_212 (O_212,N_2990,N_2979);
nand UO_213 (O_213,N_2987,N_2942);
nand UO_214 (O_214,N_2983,N_2942);
nor UO_215 (O_215,N_2936,N_2973);
xnor UO_216 (O_216,N_2971,N_2980);
xor UO_217 (O_217,N_2909,N_2942);
and UO_218 (O_218,N_2921,N_2987);
or UO_219 (O_219,N_2996,N_2915);
or UO_220 (O_220,N_2923,N_2922);
nand UO_221 (O_221,N_2965,N_2999);
nor UO_222 (O_222,N_2964,N_2954);
or UO_223 (O_223,N_2982,N_2927);
xor UO_224 (O_224,N_2925,N_2950);
nand UO_225 (O_225,N_2913,N_2902);
and UO_226 (O_226,N_2960,N_2994);
nor UO_227 (O_227,N_2968,N_2916);
nand UO_228 (O_228,N_2945,N_2967);
or UO_229 (O_229,N_2940,N_2938);
nand UO_230 (O_230,N_2950,N_2910);
and UO_231 (O_231,N_2928,N_2993);
nor UO_232 (O_232,N_2994,N_2992);
or UO_233 (O_233,N_2910,N_2997);
and UO_234 (O_234,N_2954,N_2905);
xnor UO_235 (O_235,N_2980,N_2954);
and UO_236 (O_236,N_2936,N_2947);
and UO_237 (O_237,N_2989,N_2924);
or UO_238 (O_238,N_2985,N_2963);
xor UO_239 (O_239,N_2986,N_2954);
and UO_240 (O_240,N_2993,N_2989);
nor UO_241 (O_241,N_2936,N_2903);
xor UO_242 (O_242,N_2946,N_2982);
nor UO_243 (O_243,N_2998,N_2958);
or UO_244 (O_244,N_2912,N_2968);
xor UO_245 (O_245,N_2948,N_2965);
or UO_246 (O_246,N_2923,N_2940);
or UO_247 (O_247,N_2901,N_2962);
or UO_248 (O_248,N_2969,N_2973);
xor UO_249 (O_249,N_2940,N_2971);
nand UO_250 (O_250,N_2904,N_2922);
xor UO_251 (O_251,N_2953,N_2937);
xor UO_252 (O_252,N_2970,N_2917);
xnor UO_253 (O_253,N_2902,N_2910);
nand UO_254 (O_254,N_2975,N_2919);
or UO_255 (O_255,N_2972,N_2976);
nand UO_256 (O_256,N_2937,N_2910);
xnor UO_257 (O_257,N_2971,N_2987);
xor UO_258 (O_258,N_2937,N_2932);
and UO_259 (O_259,N_2953,N_2997);
xor UO_260 (O_260,N_2939,N_2952);
and UO_261 (O_261,N_2958,N_2923);
and UO_262 (O_262,N_2918,N_2940);
nor UO_263 (O_263,N_2918,N_2955);
or UO_264 (O_264,N_2986,N_2970);
nand UO_265 (O_265,N_2984,N_2971);
nor UO_266 (O_266,N_2956,N_2964);
and UO_267 (O_267,N_2944,N_2973);
xor UO_268 (O_268,N_2975,N_2956);
nor UO_269 (O_269,N_2959,N_2955);
nor UO_270 (O_270,N_2980,N_2952);
and UO_271 (O_271,N_2914,N_2949);
or UO_272 (O_272,N_2947,N_2957);
nor UO_273 (O_273,N_2990,N_2999);
xor UO_274 (O_274,N_2920,N_2919);
or UO_275 (O_275,N_2933,N_2912);
and UO_276 (O_276,N_2985,N_2909);
or UO_277 (O_277,N_2993,N_2924);
xor UO_278 (O_278,N_2945,N_2995);
or UO_279 (O_279,N_2929,N_2960);
or UO_280 (O_280,N_2903,N_2979);
and UO_281 (O_281,N_2929,N_2964);
nor UO_282 (O_282,N_2915,N_2998);
nor UO_283 (O_283,N_2938,N_2942);
or UO_284 (O_284,N_2955,N_2910);
xor UO_285 (O_285,N_2992,N_2918);
xor UO_286 (O_286,N_2942,N_2991);
nor UO_287 (O_287,N_2930,N_2957);
or UO_288 (O_288,N_2913,N_2921);
nor UO_289 (O_289,N_2981,N_2997);
or UO_290 (O_290,N_2967,N_2910);
or UO_291 (O_291,N_2958,N_2915);
nand UO_292 (O_292,N_2918,N_2982);
nor UO_293 (O_293,N_2933,N_2975);
nand UO_294 (O_294,N_2999,N_2955);
and UO_295 (O_295,N_2913,N_2916);
or UO_296 (O_296,N_2947,N_2939);
and UO_297 (O_297,N_2999,N_2919);
nand UO_298 (O_298,N_2943,N_2931);
nand UO_299 (O_299,N_2966,N_2981);
nand UO_300 (O_300,N_2906,N_2957);
and UO_301 (O_301,N_2985,N_2955);
xor UO_302 (O_302,N_2987,N_2907);
nand UO_303 (O_303,N_2916,N_2905);
nor UO_304 (O_304,N_2903,N_2961);
nand UO_305 (O_305,N_2917,N_2952);
nor UO_306 (O_306,N_2946,N_2900);
nand UO_307 (O_307,N_2931,N_2947);
nand UO_308 (O_308,N_2922,N_2967);
nor UO_309 (O_309,N_2955,N_2968);
nor UO_310 (O_310,N_2986,N_2931);
nand UO_311 (O_311,N_2914,N_2994);
xnor UO_312 (O_312,N_2958,N_2951);
or UO_313 (O_313,N_2900,N_2988);
nor UO_314 (O_314,N_2961,N_2916);
xor UO_315 (O_315,N_2939,N_2996);
xnor UO_316 (O_316,N_2963,N_2970);
nor UO_317 (O_317,N_2925,N_2946);
nand UO_318 (O_318,N_2912,N_2949);
xnor UO_319 (O_319,N_2922,N_2928);
and UO_320 (O_320,N_2963,N_2916);
xor UO_321 (O_321,N_2962,N_2912);
xnor UO_322 (O_322,N_2913,N_2960);
and UO_323 (O_323,N_2959,N_2913);
nor UO_324 (O_324,N_2980,N_2964);
and UO_325 (O_325,N_2988,N_2972);
nor UO_326 (O_326,N_2943,N_2950);
nand UO_327 (O_327,N_2914,N_2932);
nand UO_328 (O_328,N_2930,N_2975);
xor UO_329 (O_329,N_2964,N_2927);
xor UO_330 (O_330,N_2928,N_2902);
nor UO_331 (O_331,N_2944,N_2987);
or UO_332 (O_332,N_2938,N_2989);
and UO_333 (O_333,N_2973,N_2940);
xnor UO_334 (O_334,N_2928,N_2943);
nor UO_335 (O_335,N_2946,N_2936);
or UO_336 (O_336,N_2998,N_2963);
and UO_337 (O_337,N_2915,N_2968);
nor UO_338 (O_338,N_2941,N_2920);
or UO_339 (O_339,N_2940,N_2960);
and UO_340 (O_340,N_2942,N_2913);
nor UO_341 (O_341,N_2964,N_2930);
nor UO_342 (O_342,N_2959,N_2944);
or UO_343 (O_343,N_2936,N_2979);
and UO_344 (O_344,N_2953,N_2924);
xor UO_345 (O_345,N_2932,N_2910);
or UO_346 (O_346,N_2924,N_2970);
and UO_347 (O_347,N_2971,N_2923);
nor UO_348 (O_348,N_2923,N_2919);
nand UO_349 (O_349,N_2942,N_2997);
and UO_350 (O_350,N_2901,N_2996);
xnor UO_351 (O_351,N_2978,N_2943);
or UO_352 (O_352,N_2910,N_2963);
and UO_353 (O_353,N_2917,N_2998);
nor UO_354 (O_354,N_2984,N_2987);
xnor UO_355 (O_355,N_2947,N_2920);
and UO_356 (O_356,N_2956,N_2935);
and UO_357 (O_357,N_2908,N_2944);
or UO_358 (O_358,N_2954,N_2942);
xnor UO_359 (O_359,N_2978,N_2934);
xnor UO_360 (O_360,N_2992,N_2911);
nor UO_361 (O_361,N_2936,N_2976);
or UO_362 (O_362,N_2946,N_2988);
nor UO_363 (O_363,N_2942,N_2981);
and UO_364 (O_364,N_2955,N_2948);
xor UO_365 (O_365,N_2983,N_2991);
or UO_366 (O_366,N_2961,N_2900);
and UO_367 (O_367,N_2932,N_2989);
nor UO_368 (O_368,N_2919,N_2970);
or UO_369 (O_369,N_2956,N_2916);
xor UO_370 (O_370,N_2993,N_2941);
xnor UO_371 (O_371,N_2941,N_2922);
nand UO_372 (O_372,N_2905,N_2917);
or UO_373 (O_373,N_2992,N_2916);
or UO_374 (O_374,N_2945,N_2991);
xor UO_375 (O_375,N_2928,N_2951);
xnor UO_376 (O_376,N_2952,N_2943);
or UO_377 (O_377,N_2956,N_2953);
nor UO_378 (O_378,N_2937,N_2978);
and UO_379 (O_379,N_2959,N_2957);
or UO_380 (O_380,N_2942,N_2955);
nand UO_381 (O_381,N_2966,N_2947);
xor UO_382 (O_382,N_2994,N_2964);
and UO_383 (O_383,N_2938,N_2909);
and UO_384 (O_384,N_2990,N_2969);
and UO_385 (O_385,N_2990,N_2919);
nand UO_386 (O_386,N_2907,N_2923);
or UO_387 (O_387,N_2936,N_2964);
nand UO_388 (O_388,N_2950,N_2932);
nor UO_389 (O_389,N_2956,N_2986);
and UO_390 (O_390,N_2934,N_2955);
nand UO_391 (O_391,N_2948,N_2998);
nor UO_392 (O_392,N_2969,N_2915);
nand UO_393 (O_393,N_2925,N_2928);
and UO_394 (O_394,N_2935,N_2988);
nand UO_395 (O_395,N_2936,N_2996);
xnor UO_396 (O_396,N_2963,N_2997);
nand UO_397 (O_397,N_2993,N_2918);
or UO_398 (O_398,N_2915,N_2970);
and UO_399 (O_399,N_2903,N_2926);
and UO_400 (O_400,N_2902,N_2901);
nand UO_401 (O_401,N_2997,N_2987);
or UO_402 (O_402,N_2931,N_2926);
nor UO_403 (O_403,N_2979,N_2957);
and UO_404 (O_404,N_2980,N_2989);
nor UO_405 (O_405,N_2943,N_2959);
or UO_406 (O_406,N_2958,N_2936);
or UO_407 (O_407,N_2968,N_2919);
nor UO_408 (O_408,N_2927,N_2912);
and UO_409 (O_409,N_2964,N_2951);
and UO_410 (O_410,N_2914,N_2974);
or UO_411 (O_411,N_2987,N_2950);
or UO_412 (O_412,N_2910,N_2978);
or UO_413 (O_413,N_2965,N_2934);
xnor UO_414 (O_414,N_2996,N_2927);
nand UO_415 (O_415,N_2958,N_2973);
nor UO_416 (O_416,N_2966,N_2997);
and UO_417 (O_417,N_2912,N_2944);
xor UO_418 (O_418,N_2993,N_2934);
or UO_419 (O_419,N_2950,N_2907);
nand UO_420 (O_420,N_2935,N_2933);
and UO_421 (O_421,N_2987,N_2964);
xnor UO_422 (O_422,N_2932,N_2961);
xnor UO_423 (O_423,N_2982,N_2952);
or UO_424 (O_424,N_2910,N_2926);
nor UO_425 (O_425,N_2944,N_2935);
nor UO_426 (O_426,N_2962,N_2987);
nand UO_427 (O_427,N_2917,N_2977);
nand UO_428 (O_428,N_2929,N_2913);
or UO_429 (O_429,N_2932,N_2911);
xor UO_430 (O_430,N_2922,N_2986);
xnor UO_431 (O_431,N_2962,N_2930);
nor UO_432 (O_432,N_2911,N_2908);
nor UO_433 (O_433,N_2982,N_2934);
or UO_434 (O_434,N_2957,N_2956);
xnor UO_435 (O_435,N_2978,N_2924);
and UO_436 (O_436,N_2901,N_2958);
and UO_437 (O_437,N_2961,N_2957);
and UO_438 (O_438,N_2999,N_2973);
nor UO_439 (O_439,N_2914,N_2953);
and UO_440 (O_440,N_2989,N_2978);
xnor UO_441 (O_441,N_2916,N_2946);
nand UO_442 (O_442,N_2980,N_2937);
or UO_443 (O_443,N_2963,N_2937);
xnor UO_444 (O_444,N_2950,N_2911);
nor UO_445 (O_445,N_2961,N_2956);
xnor UO_446 (O_446,N_2930,N_2952);
nand UO_447 (O_447,N_2947,N_2983);
or UO_448 (O_448,N_2992,N_2986);
nor UO_449 (O_449,N_2947,N_2901);
nor UO_450 (O_450,N_2912,N_2969);
xor UO_451 (O_451,N_2911,N_2969);
and UO_452 (O_452,N_2916,N_2909);
nand UO_453 (O_453,N_2926,N_2966);
or UO_454 (O_454,N_2955,N_2961);
xor UO_455 (O_455,N_2973,N_2900);
nor UO_456 (O_456,N_2969,N_2952);
or UO_457 (O_457,N_2979,N_2999);
and UO_458 (O_458,N_2977,N_2930);
nor UO_459 (O_459,N_2996,N_2974);
and UO_460 (O_460,N_2931,N_2983);
and UO_461 (O_461,N_2943,N_2914);
nor UO_462 (O_462,N_2909,N_2924);
nor UO_463 (O_463,N_2978,N_2957);
nand UO_464 (O_464,N_2982,N_2961);
nor UO_465 (O_465,N_2941,N_2945);
and UO_466 (O_466,N_2974,N_2918);
xor UO_467 (O_467,N_2923,N_2937);
nand UO_468 (O_468,N_2939,N_2936);
nor UO_469 (O_469,N_2906,N_2924);
xor UO_470 (O_470,N_2969,N_2982);
or UO_471 (O_471,N_2938,N_2966);
or UO_472 (O_472,N_2983,N_2992);
or UO_473 (O_473,N_2998,N_2930);
or UO_474 (O_474,N_2948,N_2926);
nor UO_475 (O_475,N_2987,N_2935);
nor UO_476 (O_476,N_2974,N_2963);
or UO_477 (O_477,N_2962,N_2908);
xnor UO_478 (O_478,N_2913,N_2930);
nand UO_479 (O_479,N_2957,N_2925);
nor UO_480 (O_480,N_2994,N_2988);
nand UO_481 (O_481,N_2990,N_2986);
or UO_482 (O_482,N_2970,N_2958);
xnor UO_483 (O_483,N_2934,N_2950);
xor UO_484 (O_484,N_2970,N_2925);
nor UO_485 (O_485,N_2974,N_2982);
and UO_486 (O_486,N_2942,N_2931);
and UO_487 (O_487,N_2992,N_2900);
and UO_488 (O_488,N_2995,N_2920);
xor UO_489 (O_489,N_2998,N_2990);
or UO_490 (O_490,N_2907,N_2927);
xnor UO_491 (O_491,N_2905,N_2956);
nor UO_492 (O_492,N_2977,N_2955);
xnor UO_493 (O_493,N_2907,N_2967);
xor UO_494 (O_494,N_2992,N_2902);
xor UO_495 (O_495,N_2964,N_2957);
and UO_496 (O_496,N_2928,N_2980);
and UO_497 (O_497,N_2929,N_2949);
nand UO_498 (O_498,N_2949,N_2922);
nand UO_499 (O_499,N_2952,N_2937);
endmodule