module basic_5000_50000_5000_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_4328,In_1581);
or U1 (N_1,In_2360,In_3389);
nor U2 (N_2,In_3406,In_4225);
and U3 (N_3,In_995,In_4965);
nand U4 (N_4,In_2408,In_4239);
nor U5 (N_5,In_1726,In_802);
nor U6 (N_6,In_360,In_249);
and U7 (N_7,In_3034,In_4297);
and U8 (N_8,In_197,In_3713);
nand U9 (N_9,In_4571,In_4096);
or U10 (N_10,In_104,In_1071);
and U11 (N_11,In_2516,In_34);
nor U12 (N_12,In_1374,In_1175);
or U13 (N_13,In_533,In_2817);
nor U14 (N_14,In_1112,In_471);
nand U15 (N_15,In_3162,In_3345);
or U16 (N_16,In_4625,In_1395);
or U17 (N_17,In_1085,In_3896);
nand U18 (N_18,In_2785,In_729);
nor U19 (N_19,In_2891,In_4268);
or U20 (N_20,In_1222,In_1350);
xor U21 (N_21,In_3718,In_786);
xor U22 (N_22,In_1436,In_4326);
or U23 (N_23,In_309,In_1540);
and U24 (N_24,In_4934,In_89);
xnor U25 (N_25,In_968,In_4336);
nand U26 (N_26,In_3182,In_1714);
xnor U27 (N_27,In_2925,In_3);
or U28 (N_28,In_1722,In_772);
xor U29 (N_29,In_1300,In_956);
nand U30 (N_30,In_2474,In_3376);
nor U31 (N_31,In_4006,In_4659);
xnor U32 (N_32,In_4022,In_390);
or U33 (N_33,In_1546,In_3271);
nand U34 (N_34,In_2828,In_3469);
nor U35 (N_35,In_593,In_2297);
nand U36 (N_36,In_3971,In_1621);
or U37 (N_37,In_1002,In_3094);
xnor U38 (N_38,In_3481,In_2560);
or U39 (N_39,In_1160,In_209);
nor U40 (N_40,In_3688,In_2367);
and U41 (N_41,In_1593,In_3213);
nand U42 (N_42,In_2200,In_3083);
or U43 (N_43,In_2406,In_359);
or U44 (N_44,In_4802,In_2740);
xor U45 (N_45,In_2806,In_2219);
and U46 (N_46,In_4139,In_3489);
nand U47 (N_47,In_2656,In_2136);
or U48 (N_48,In_2050,In_4294);
and U49 (N_49,In_3757,In_326);
nor U50 (N_50,In_3842,In_301);
xor U51 (N_51,In_2939,In_3535);
xnor U52 (N_52,In_32,In_906);
nand U53 (N_53,In_3789,In_3076);
and U54 (N_54,In_1569,In_929);
nand U55 (N_55,In_988,In_1104);
and U56 (N_56,In_520,In_4766);
nand U57 (N_57,In_71,In_3049);
or U58 (N_58,In_4719,In_3772);
and U59 (N_59,In_4843,In_1848);
and U60 (N_60,In_1503,In_3326);
nor U61 (N_61,In_4630,In_3024);
or U62 (N_62,In_4039,In_728);
and U63 (N_63,In_228,In_2549);
and U64 (N_64,In_4542,In_2552);
nor U65 (N_65,In_3092,In_3671);
nor U66 (N_66,In_4455,In_290);
and U67 (N_67,In_4560,In_1629);
or U68 (N_68,In_3091,In_3110);
or U69 (N_69,In_2016,In_3126);
and U70 (N_70,In_4673,In_4536);
nand U71 (N_71,In_3267,In_2147);
and U72 (N_72,In_95,In_4358);
nor U73 (N_73,In_2840,In_756);
xnor U74 (N_74,In_1872,In_1542);
nand U75 (N_75,In_1095,In_3189);
or U76 (N_76,In_2410,In_3235);
nand U77 (N_77,In_1319,In_2600);
nor U78 (N_78,In_834,In_332);
and U79 (N_79,In_3036,In_779);
nand U80 (N_80,In_3550,In_3264);
nand U81 (N_81,In_886,In_4587);
or U82 (N_82,In_3350,In_1885);
nand U83 (N_83,In_1105,In_2567);
nor U84 (N_84,In_3428,In_4230);
xor U85 (N_85,In_4547,In_4482);
nand U86 (N_86,In_1197,In_4024);
or U87 (N_87,In_3392,In_4506);
nand U88 (N_88,In_3624,In_3736);
nand U89 (N_89,In_4304,In_1428);
and U90 (N_90,In_1277,In_3784);
and U91 (N_91,In_2524,In_1834);
nor U92 (N_92,In_1662,In_547);
and U93 (N_93,In_3433,In_3445);
and U94 (N_94,In_3722,In_1548);
nand U95 (N_95,In_4084,In_1194);
xor U96 (N_96,In_626,In_414);
or U97 (N_97,In_1437,In_2454);
nand U98 (N_98,In_665,In_595);
nand U99 (N_99,In_4957,In_438);
nand U100 (N_100,In_3773,In_2696);
or U101 (N_101,In_494,In_3467);
nand U102 (N_102,In_3561,In_640);
nand U103 (N_103,In_1559,In_4056);
nor U104 (N_104,In_3030,In_3287);
nor U105 (N_105,In_4503,In_2232);
and U106 (N_106,In_1142,In_4150);
xnor U107 (N_107,In_231,In_1989);
and U108 (N_108,In_1801,In_199);
nand U109 (N_109,In_4157,In_3988);
nand U110 (N_110,In_4199,In_872);
nand U111 (N_111,In_240,In_2397);
xor U112 (N_112,In_1249,In_2679);
nand U113 (N_113,In_1132,In_2929);
nand U114 (N_114,In_4977,In_3894);
and U115 (N_115,In_939,In_2058);
xnor U116 (N_116,In_3554,In_40);
and U117 (N_117,In_769,In_2803);
and U118 (N_118,In_3727,In_4208);
nand U119 (N_119,In_3976,In_2370);
or U120 (N_120,In_4705,In_3650);
and U121 (N_121,In_3626,In_2513);
xor U122 (N_122,In_4858,In_4606);
nand U123 (N_123,In_4025,In_1878);
nor U124 (N_124,In_2722,In_3869);
nor U125 (N_125,In_2018,In_537);
nor U126 (N_126,In_3037,In_4841);
nand U127 (N_127,In_541,In_554);
or U128 (N_128,In_465,In_3482);
nor U129 (N_129,In_2966,In_1557);
or U130 (N_130,In_4877,In_2731);
and U131 (N_131,In_3021,In_2555);
nand U132 (N_132,In_1740,In_1995);
xnor U133 (N_133,In_1487,In_4395);
and U134 (N_134,In_283,In_3760);
or U135 (N_135,In_4464,In_244);
nand U136 (N_136,In_523,In_1278);
nor U137 (N_137,In_3101,In_3663);
or U138 (N_138,In_1092,In_2546);
xnor U139 (N_139,In_325,In_1576);
or U140 (N_140,In_4295,In_2654);
or U141 (N_141,In_1727,In_2180);
xor U142 (N_142,In_1154,In_2871);
nor U143 (N_143,In_3479,In_1620);
nor U144 (N_144,In_2063,In_1167);
or U145 (N_145,In_4098,In_2564);
xor U146 (N_146,In_2575,In_1490);
or U147 (N_147,In_4551,In_4062);
and U148 (N_148,In_2212,In_3812);
nor U149 (N_149,In_2621,In_121);
nand U150 (N_150,In_1813,In_3129);
nand U151 (N_151,In_4716,In_2206);
or U152 (N_152,In_3953,In_2968);
and U153 (N_153,In_2222,In_4377);
nand U154 (N_154,In_1238,In_3415);
or U155 (N_155,In_4317,In_1803);
and U156 (N_156,In_526,In_2436);
nand U157 (N_157,In_741,In_4829);
nand U158 (N_158,In_2745,In_4605);
or U159 (N_159,In_4773,In_4123);
xor U160 (N_160,In_511,In_2962);
or U161 (N_161,In_2563,In_3690);
xnor U162 (N_162,In_885,In_269);
xor U163 (N_163,In_2375,In_850);
xor U164 (N_164,In_1296,In_4881);
xnor U165 (N_165,In_4701,In_924);
and U166 (N_166,In_621,In_223);
nor U167 (N_167,In_4759,In_696);
nor U168 (N_168,In_4253,In_4921);
or U169 (N_169,In_2257,In_3693);
nand U170 (N_170,In_4930,In_113);
nor U171 (N_171,In_4472,In_67);
and U172 (N_172,In_2495,In_1121);
or U173 (N_173,In_1931,In_4867);
or U174 (N_174,In_2044,In_1728);
nor U175 (N_175,In_2814,In_3141);
or U176 (N_176,In_3446,In_3518);
and U177 (N_177,In_4436,In_3526);
xor U178 (N_178,In_4601,In_3405);
and U179 (N_179,In_2706,In_3174);
or U180 (N_180,In_905,In_1405);
nor U181 (N_181,In_970,In_2580);
xor U182 (N_182,In_3848,In_30);
or U183 (N_183,In_2277,In_3991);
nor U184 (N_184,In_4362,In_3364);
xor U185 (N_185,In_3199,In_74);
and U186 (N_186,In_208,In_4939);
nand U187 (N_187,In_58,In_4623);
nor U188 (N_188,In_2686,In_490);
nand U189 (N_189,In_1688,In_3765);
or U190 (N_190,In_862,In_4220);
xnor U191 (N_191,In_1516,In_3378);
and U192 (N_192,In_2320,In_2490);
nand U193 (N_193,In_4009,In_4197);
nand U194 (N_194,In_726,In_3029);
and U195 (N_195,In_3439,In_1215);
nor U196 (N_196,In_4776,In_766);
or U197 (N_197,In_1709,In_1274);
nor U198 (N_198,In_4189,In_1847);
and U199 (N_199,In_4653,In_702);
nand U200 (N_200,In_2221,In_1207);
nor U201 (N_201,In_4669,In_2841);
nand U202 (N_202,In_1065,In_2215);
nand U203 (N_203,In_923,In_758);
nand U204 (N_204,In_2718,In_708);
nor U205 (N_205,In_77,In_4651);
nand U206 (N_206,In_3994,In_3924);
xnor U207 (N_207,In_1669,In_2444);
and U208 (N_208,In_1473,In_3057);
nand U209 (N_209,In_3438,In_2046);
and U210 (N_210,In_3590,In_1280);
nor U211 (N_211,In_3532,In_4683);
or U212 (N_212,In_2576,In_2970);
and U213 (N_213,In_2682,In_647);
nand U214 (N_214,In_506,In_484);
xor U215 (N_215,In_773,In_4767);
nor U216 (N_216,In_4219,In_2847);
or U217 (N_217,In_791,In_211);
and U218 (N_218,In_3654,In_1515);
xor U219 (N_219,In_765,In_4037);
or U220 (N_220,In_2164,In_200);
nor U221 (N_221,In_3181,In_2298);
and U222 (N_222,In_3601,In_842);
or U223 (N_223,In_1743,In_3011);
or U224 (N_224,In_3062,In_338);
nand U225 (N_225,In_3293,In_1285);
and U226 (N_226,In_4805,In_3973);
nand U227 (N_227,In_1959,In_2496);
nand U228 (N_228,In_2240,In_3735);
xnor U229 (N_229,In_4207,In_4308);
xnor U230 (N_230,In_3102,In_318);
nand U231 (N_231,In_3290,In_3192);
nor U232 (N_232,In_2933,In_4280);
nand U233 (N_233,In_2274,In_3764);
nand U234 (N_234,In_497,In_198);
and U235 (N_235,In_1413,In_3946);
or U236 (N_236,In_2168,In_2752);
xnor U237 (N_237,In_4698,In_4964);
nand U238 (N_238,In_946,In_3336);
xor U239 (N_239,In_3357,In_835);
nor U240 (N_240,In_2315,In_1262);
xor U241 (N_241,In_307,In_2651);
or U242 (N_242,In_2897,In_3571);
xor U243 (N_243,In_2479,In_4912);
or U244 (N_244,In_2793,In_704);
nand U245 (N_245,In_451,In_1140);
nor U246 (N_246,In_568,In_1391);
or U247 (N_247,In_2707,In_3344);
or U248 (N_248,In_342,In_658);
and U249 (N_249,In_3634,In_860);
and U250 (N_250,In_972,In_2505);
and U251 (N_251,In_3979,In_1416);
nand U252 (N_252,In_4201,In_4051);
xor U253 (N_253,In_3952,In_4130);
xor U254 (N_254,In_4909,In_1764);
or U255 (N_255,In_1565,In_263);
nand U256 (N_256,In_1307,In_4764);
and U257 (N_257,In_1076,In_3221);
or U258 (N_258,In_3067,In_4182);
and U259 (N_259,In_1725,In_1054);
nor U260 (N_260,In_2211,In_1499);
and U261 (N_261,In_1116,In_3215);
nand U262 (N_262,In_617,In_587);
xnor U263 (N_263,In_3868,In_757);
and U264 (N_264,In_559,In_3012);
or U265 (N_265,In_4332,In_4307);
xnor U266 (N_266,In_2204,In_3921);
and U267 (N_267,In_2171,In_967);
or U268 (N_268,In_1053,In_3105);
nand U269 (N_269,In_4596,In_1288);
and U270 (N_270,In_2392,In_4520);
nor U271 (N_271,In_3200,In_11);
nor U272 (N_272,In_480,In_2059);
or U273 (N_273,In_4710,In_4413);
nand U274 (N_274,In_420,In_1470);
nand U275 (N_275,In_4165,In_685);
and U276 (N_276,In_2174,In_2019);
or U277 (N_277,In_4272,In_560);
and U278 (N_278,In_2771,In_2708);
xnor U279 (N_279,In_2156,In_543);
nor U280 (N_280,In_2007,In_2636);
or U281 (N_281,In_2339,In_3104);
and U282 (N_282,In_1228,In_1827);
and U283 (N_283,In_3202,In_69);
nand U284 (N_284,In_3609,In_2862);
or U285 (N_285,In_408,In_395);
and U286 (N_286,In_4687,In_1013);
or U287 (N_287,In_3513,In_133);
or U288 (N_288,In_1275,In_399);
nor U289 (N_289,In_590,In_4450);
nor U290 (N_290,In_4576,In_1097);
and U291 (N_291,In_4343,In_8);
or U292 (N_292,In_501,In_57);
or U293 (N_293,In_1911,In_3417);
and U294 (N_294,In_4554,In_402);
nand U295 (N_295,In_1298,In_2231);
or U296 (N_296,In_3472,In_4402);
and U297 (N_297,In_2721,In_4092);
xor U298 (N_298,In_4363,In_4539);
xor U299 (N_299,In_1840,In_3849);
nand U300 (N_300,In_4209,In_798);
nand U301 (N_301,In_3879,In_4963);
or U302 (N_302,In_1073,In_1720);
and U303 (N_303,In_4137,In_1927);
nor U304 (N_304,In_1412,In_4211);
xnor U305 (N_305,In_4176,In_636);
nor U306 (N_306,In_3943,In_4310);
and U307 (N_307,In_1493,In_2661);
nand U308 (N_308,In_4846,In_1291);
nand U309 (N_309,In_4043,In_2511);
nor U310 (N_310,In_2057,In_4848);
and U311 (N_311,In_4240,In_2162);
nor U312 (N_312,In_2714,In_1435);
nor U313 (N_313,In_2312,In_1019);
nand U314 (N_314,In_4751,In_4706);
xor U315 (N_315,In_527,In_1164);
nor U316 (N_316,In_994,In_744);
and U317 (N_317,In_2247,In_2477);
or U318 (N_318,In_2885,In_2758);
nor U319 (N_319,In_750,In_461);
and U320 (N_320,In_2356,In_1538);
nor U321 (N_321,In_205,In_407);
nor U322 (N_322,In_3004,In_1052);
and U323 (N_323,In_838,In_2955);
nor U324 (N_324,In_4899,In_3954);
xor U325 (N_325,In_37,In_4016);
xor U326 (N_326,In_2846,In_1506);
nand U327 (N_327,In_4195,In_1924);
nand U328 (N_328,In_24,In_1525);
nand U329 (N_329,In_3567,In_4515);
or U330 (N_330,In_4597,In_1809);
xor U331 (N_331,In_4237,In_128);
xnor U332 (N_332,In_83,In_1637);
nor U333 (N_333,In_4690,In_1657);
xor U334 (N_334,In_122,In_4271);
nand U335 (N_335,In_837,In_2311);
nand U336 (N_336,In_1083,In_3338);
and U337 (N_337,In_1510,In_118);
xor U338 (N_338,In_59,In_2306);
nand U339 (N_339,In_3209,In_3730);
or U340 (N_340,In_3368,In_3777);
nor U341 (N_341,In_1220,In_1254);
and U342 (N_342,In_4541,In_4958);
xor U343 (N_343,In_1929,In_4465);
and U344 (N_344,In_1876,In_22);
xnor U345 (N_345,In_1336,In_2042);
and U346 (N_346,In_3726,In_170);
nand U347 (N_347,In_813,In_887);
and U348 (N_348,In_3632,In_2591);
xnor U349 (N_349,In_4948,In_2083);
or U350 (N_350,In_3606,In_610);
or U351 (N_351,In_109,In_1068);
or U352 (N_352,In_2643,In_2028);
nand U353 (N_353,In_927,In_1842);
nor U354 (N_354,In_852,In_3099);
nand U355 (N_355,In_3507,In_1987);
and U356 (N_356,In_695,In_4386);
and U357 (N_357,In_571,In_2514);
nand U358 (N_358,In_3116,In_3697);
and U359 (N_359,In_1839,In_3332);
or U360 (N_360,In_4089,In_39);
nand U361 (N_361,In_4447,In_2123);
xor U362 (N_362,In_4346,In_4610);
or U363 (N_363,In_3164,In_462);
nand U364 (N_364,In_3000,In_352);
xnor U365 (N_365,In_893,In_131);
nand U366 (N_366,In_3488,In_220);
xor U367 (N_367,In_4278,In_1912);
and U368 (N_368,In_3574,In_1712);
or U369 (N_369,In_4734,In_3889);
nand U370 (N_370,In_1600,In_320);
and U371 (N_371,In_19,In_528);
nand U372 (N_372,In_2908,In_683);
xor U373 (N_373,In_1494,In_578);
nor U374 (N_374,In_2244,In_3819);
xor U375 (N_375,In_3674,In_164);
or U376 (N_376,In_2744,In_2673);
nor U377 (N_377,In_44,In_2003);
nor U378 (N_378,In_1252,In_2602);
nor U379 (N_379,In_1102,In_3755);
and U380 (N_380,In_3808,In_1508);
and U381 (N_381,In_1123,In_3270);
nor U382 (N_382,In_3802,In_4086);
nor U383 (N_383,In_4354,In_1696);
nand U384 (N_384,In_637,In_4248);
or U385 (N_385,In_277,In_4978);
and U386 (N_386,In_1265,In_4441);
or U387 (N_387,In_4947,In_2622);
and U388 (N_388,In_3804,In_2798);
nor U389 (N_389,In_4969,In_4642);
nor U390 (N_390,In_3843,In_990);
or U391 (N_391,In_2776,In_1545);
xor U392 (N_392,In_472,In_4142);
xor U393 (N_393,In_423,In_2394);
and U394 (N_394,In_2405,In_1359);
and U395 (N_395,In_151,In_4353);
nand U396 (N_396,In_1321,In_4565);
or U397 (N_397,In_1532,In_317);
nand U398 (N_398,In_4911,In_4493);
xor U399 (N_399,In_2617,In_1241);
xnor U400 (N_400,In_2227,In_3448);
nand U401 (N_401,In_964,In_1676);
nor U402 (N_402,In_2012,In_1214);
or U403 (N_403,In_1653,In_2482);
or U404 (N_404,In_3915,In_4648);
xnor U405 (N_405,In_4111,In_4793);
xor U406 (N_406,In_3173,In_219);
and U407 (N_407,In_3006,In_3124);
and U408 (N_408,In_4933,In_2569);
nor U409 (N_409,In_2309,In_689);
or U410 (N_410,In_1426,In_4257);
nand U411 (N_411,In_2005,In_1124);
xor U412 (N_412,In_3087,In_4488);
xor U413 (N_413,In_2074,In_4010);
xnor U414 (N_414,In_1198,In_2048);
or U415 (N_415,In_2431,In_4992);
nor U416 (N_416,In_1820,In_4632);
nand U417 (N_417,In_4847,In_3207);
nor U418 (N_418,In_4997,In_549);
and U419 (N_419,In_1447,In_1287);
nor U420 (N_420,In_794,In_2228);
or U421 (N_421,In_2856,In_4404);
nand U422 (N_422,In_2570,In_2484);
nand U423 (N_423,In_1710,In_1571);
or U424 (N_424,In_2066,In_4399);
nor U425 (N_425,In_1385,In_194);
xor U426 (N_426,In_586,In_4035);
xor U427 (N_427,In_3888,In_4255);
or U428 (N_428,In_4770,In_4518);
or U429 (N_429,In_1836,In_4627);
or U430 (N_430,In_2521,In_4558);
or U431 (N_431,In_1587,In_357);
xnor U432 (N_432,In_3331,In_980);
or U433 (N_433,In_2006,In_2415);
xnor U434 (N_434,In_3038,In_4063);
and U435 (N_435,In_1382,In_3762);
or U436 (N_436,In_2184,In_3410);
and U437 (N_437,In_2254,In_3020);
and U438 (N_438,In_1831,In_2697);
nand U439 (N_439,In_2928,In_1425);
or U440 (N_440,In_2157,In_406);
and U441 (N_441,In_2811,In_2121);
nand U442 (N_442,In_4507,In_1877);
xor U443 (N_443,In_1145,In_2684);
nand U444 (N_444,In_3964,In_1477);
xnor U445 (N_445,In_3680,In_3065);
xor U446 (N_446,In_1509,In_2336);
nor U447 (N_447,In_1458,In_2378);
and U448 (N_448,In_4882,In_314);
nand U449 (N_449,In_2276,In_3635);
nor U450 (N_450,In_2537,In_1675);
nor U451 (N_451,In_188,In_3325);
nor U452 (N_452,In_392,In_4898);
and U453 (N_453,In_4616,In_1816);
nor U454 (N_454,In_1334,In_4820);
nand U455 (N_455,In_4049,In_3531);
or U456 (N_456,In_4186,In_4247);
nand U457 (N_457,In_2813,In_1129);
nor U458 (N_458,In_276,In_3778);
nand U459 (N_459,In_1534,In_187);
nand U460 (N_460,In_4030,In_3462);
and U461 (N_461,In_4607,In_687);
xnor U462 (N_462,In_2509,In_2216);
nor U463 (N_463,In_3534,In_4754);
nand U464 (N_464,In_2690,In_3337);
nor U465 (N_465,In_4755,In_4801);
nand U466 (N_466,In_1967,In_4810);
nor U467 (N_467,In_4187,In_216);
nand U468 (N_468,In_3908,In_975);
and U469 (N_469,In_346,In_1267);
nand U470 (N_470,In_1830,In_62);
or U471 (N_471,In_2723,In_2150);
or U472 (N_472,In_20,In_3905);
nor U473 (N_473,In_2559,In_4298);
or U474 (N_474,In_2238,In_4214);
or U475 (N_475,In_1928,In_3224);
or U476 (N_476,In_75,In_4835);
or U477 (N_477,In_2676,In_1846);
or U478 (N_478,In_3568,In_4168);
nor U479 (N_479,In_3453,In_335);
xor U480 (N_480,In_1772,In_4549);
xor U481 (N_481,In_488,In_4046);
or U482 (N_482,In_907,In_3340);
and U483 (N_483,In_2849,In_902);
nand U484 (N_484,In_3549,In_1161);
nor U485 (N_485,In_265,In_1560);
nand U486 (N_486,In_3045,In_4634);
and U487 (N_487,In_3656,In_2198);
xor U488 (N_488,In_1971,In_1818);
nor U489 (N_489,In_4804,In_4366);
or U490 (N_490,In_1256,In_4420);
xor U491 (N_491,In_442,In_755);
and U492 (N_492,In_4663,In_3125);
or U493 (N_493,In_3519,In_2937);
or U494 (N_494,In_378,In_1103);
nand U495 (N_495,In_98,In_799);
xor U496 (N_496,In_2314,In_3247);
xor U497 (N_497,In_3967,In_3551);
and U498 (N_498,In_1258,In_2593);
nand U499 (N_499,In_581,In_1551);
nor U500 (N_500,In_2615,In_788);
and U501 (N_501,In_4680,In_4756);
and U502 (N_502,In_1991,In_816);
xor U503 (N_503,In_2627,In_4073);
xnor U504 (N_504,In_3008,In_1041);
or U505 (N_505,In_1535,In_3607);
nor U506 (N_506,In_3137,In_1936);
and U507 (N_507,In_2548,In_3307);
and U508 (N_508,In_1146,In_2073);
xor U509 (N_509,In_2630,In_2361);
nor U510 (N_510,In_594,In_2426);
and U511 (N_511,In_2584,In_3782);
xor U512 (N_512,In_334,In_1875);
and U513 (N_513,In_3814,In_1673);
and U514 (N_514,In_2487,In_1978);
xor U515 (N_515,In_4335,In_377);
and U516 (N_516,In_1719,In_792);
nand U517 (N_517,In_3176,In_4875);
xnor U518 (N_518,In_2,In_3545);
or U519 (N_519,In_841,In_692);
and U520 (N_520,In_950,In_2747);
nor U521 (N_521,In_3014,In_4792);
nand U522 (N_522,In_2865,In_3480);
or U523 (N_523,In_374,In_4416);
xnor U524 (N_524,In_2368,In_4147);
xor U525 (N_525,In_4000,In_570);
xnor U526 (N_526,In_2236,In_2659);
xnor U527 (N_527,In_4914,In_4079);
nor U528 (N_528,In_3582,In_4374);
or U529 (N_529,In_1855,In_2753);
xnor U530 (N_530,In_2106,In_2313);
or U531 (N_531,In_4351,In_4749);
xor U532 (N_532,In_3771,In_106);
xor U533 (N_533,In_1237,In_4944);
xor U534 (N_534,In_16,In_4613);
xnor U535 (N_535,In_2757,In_153);
or U536 (N_536,In_1698,In_481);
and U537 (N_537,In_368,In_1561);
nor U538 (N_538,In_4372,In_2294);
xor U539 (N_539,In_487,In_1273);
nand U540 (N_540,In_4113,In_1367);
nand U541 (N_541,In_2823,In_1952);
nand U542 (N_542,In_2337,In_4412);
xnor U543 (N_543,In_3669,In_2137);
nand U544 (N_544,In_241,In_51);
or U545 (N_545,In_2725,In_1341);
nand U546 (N_546,In_641,In_3233);
xnor U547 (N_547,In_4537,In_2299);
nand U548 (N_548,In_4112,In_2101);
and U549 (N_549,In_1752,In_3026);
nor U550 (N_550,In_2618,In_2597);
and U551 (N_551,In_3098,In_246);
and U552 (N_552,In_409,In_976);
nand U553 (N_553,In_379,In_3088);
and U554 (N_554,In_4994,In_2249);
xnor U555 (N_555,In_4369,In_1677);
or U556 (N_556,In_1183,In_2681);
and U557 (N_557,In_4259,In_4486);
or U558 (N_558,In_3297,In_1835);
xnor U559 (N_559,In_2854,In_3179);
nand U560 (N_560,In_2507,In_3263);
or U561 (N_561,In_4048,In_4937);
or U562 (N_562,In_2353,In_1659);
xnor U563 (N_563,In_908,In_1475);
or U564 (N_564,In_3704,In_4510);
and U565 (N_565,In_605,In_4531);
xnor U566 (N_566,In_182,In_4828);
or U567 (N_567,In_2085,In_255);
or U568 (N_568,In_120,In_1170);
xnor U569 (N_569,In_2581,In_3538);
nand U570 (N_570,In_17,In_2992);
nand U571 (N_571,In_2133,In_114);
xnor U572 (N_572,In_2119,In_4557);
or U573 (N_573,In_2808,In_1605);
or U574 (N_574,In_2880,In_1084);
nor U575 (N_575,In_4501,In_2146);
or U576 (N_576,In_3166,In_3706);
nand U577 (N_577,In_3291,In_3409);
xnor U578 (N_578,In_2518,In_1650);
nor U579 (N_579,In_4380,In_189);
nor U580 (N_580,In_367,In_2892);
nand U581 (N_581,In_1407,In_2214);
and U582 (N_582,In_1857,In_3836);
nor U583 (N_583,In_3775,In_4817);
nor U584 (N_584,In_1430,In_2237);
or U585 (N_585,In_376,In_1289);
and U586 (N_586,In_1261,In_986);
xnor U587 (N_587,In_3698,In_1708);
nor U588 (N_588,In_4340,In_971);
xnor U589 (N_589,In_1086,In_4312);
nor U590 (N_590,In_10,In_2510);
nand U591 (N_591,In_1005,In_569);
nor U592 (N_592,In_4223,In_4007);
nor U593 (N_593,In_4121,In_2266);
nand U594 (N_594,In_1609,In_3185);
nor U595 (N_595,In_4563,In_733);
nor U596 (N_596,In_4926,In_676);
nor U597 (N_597,In_3058,In_401);
or U598 (N_598,In_4878,In_960);
nor U599 (N_599,In_2616,In_1397);
or U600 (N_600,In_2876,In_3312);
and U601 (N_601,In_2501,In_763);
xnor U602 (N_602,In_1860,In_4844);
nand U603 (N_603,In_2956,In_589);
or U604 (N_604,In_4838,In_1137);
nor U605 (N_605,In_572,In_1157);
and U606 (N_606,In_820,In_2031);
nor U607 (N_607,In_437,In_4812);
xor U608 (N_608,In_1524,In_724);
nor U609 (N_609,In_4720,In_4955);
and U610 (N_610,In_430,In_3436);
or U611 (N_611,In_1008,In_888);
nand U612 (N_612,In_76,In_4818);
or U613 (N_613,In_684,In_3380);
nand U614 (N_614,In_127,In_1276);
or U615 (N_615,In_3506,In_1627);
or U616 (N_616,In_2229,In_2614);
nand U617 (N_617,In_1144,In_3457);
nor U618 (N_618,In_1489,In_3353);
nor U619 (N_619,In_4564,In_1572);
nor U620 (N_620,In_3856,In_4986);
or U621 (N_621,In_3354,In_1147);
or U622 (N_622,In_2761,In_1861);
and U623 (N_623,In_38,In_2060);
and U624 (N_624,In_4134,In_1695);
nor U625 (N_625,In_3070,In_4067);
nand U626 (N_626,In_2473,In_3643);
or U627 (N_627,In_3874,In_3412);
or U628 (N_628,In_2453,In_4736);
nand U629 (N_629,In_1081,In_1235);
nor U630 (N_630,In_2363,In_3740);
xnor U631 (N_631,In_230,In_1926);
nand U632 (N_632,In_427,In_2578);
xor U633 (N_633,In_503,In_3906);
nand U634 (N_634,In_4631,In_2830);
xor U635 (N_635,In_4449,In_2869);
xor U636 (N_636,In_3280,In_149);
and U637 (N_637,In_1767,In_483);
or U638 (N_638,In_124,In_3172);
or U639 (N_639,In_2566,In_2429);
or U640 (N_640,In_4704,In_167);
xor U641 (N_641,In_2502,In_1747);
nand U642 (N_642,In_823,In_234);
xnor U643 (N_643,In_82,In_2638);
nor U644 (N_644,In_1807,In_435);
nor U645 (N_645,In_3552,In_550);
xnor U646 (N_646,In_4639,In_3352);
or U647 (N_647,In_3536,In_2609);
and U648 (N_648,In_1686,In_1642);
xor U649 (N_649,In_2967,In_1598);
and U650 (N_650,In_247,In_921);
nand U651 (N_651,In_3073,In_4246);
xnor U652 (N_652,In_3248,In_4107);
and U653 (N_653,In_3156,In_3739);
nand U654 (N_654,In_2541,In_4750);
nor U655 (N_655,In_817,In_4460);
nand U656 (N_656,In_2466,In_4163);
xor U657 (N_657,In_4580,In_2416);
or U658 (N_658,In_2921,In_1177);
nand U659 (N_659,In_4221,In_3985);
nand U660 (N_660,In_877,In_358);
nor U661 (N_661,In_2717,In_1159);
xnor U662 (N_662,In_4392,In_1998);
and U663 (N_663,In_3122,In_375);
nand U664 (N_664,In_2384,In_4254);
nor U665 (N_665,In_2858,In_3695);
and U666 (N_666,In_3089,In_4806);
xor U667 (N_667,In_2233,In_1589);
or U668 (N_668,In_1979,In_1483);
and U669 (N_669,In_3649,In_745);
nand U670 (N_670,In_4895,In_2986);
xor U671 (N_671,In_1584,In_2587);
nor U672 (N_672,In_1260,In_1257);
nand U673 (N_673,In_237,In_889);
nand U674 (N_674,In_1343,In_347);
nor U675 (N_675,In_2127,In_2920);
and U676 (N_676,In_1463,In_1520);
and U677 (N_677,In_2032,In_584);
nand U678 (N_678,In_1325,In_1741);
nor U679 (N_679,In_1628,In_2178);
xor U680 (N_680,In_671,In_1778);
nor U681 (N_681,In_2533,In_457);
nor U682 (N_682,In_2441,In_4671);
xor U683 (N_683,In_2081,In_2845);
or U684 (N_684,In_4341,In_903);
and U685 (N_685,In_4229,In_4967);
nand U686 (N_686,In_3523,In_2631);
xnor U687 (N_687,In_3790,In_270);
and U688 (N_688,In_4591,In_1155);
or U689 (N_689,In_3144,In_2881);
and U690 (N_690,In_933,In_2329);
and U691 (N_691,In_1648,In_1029);
nor U692 (N_692,In_2554,In_822);
nand U693 (N_693,In_1962,In_2588);
nand U694 (N_694,In_959,In_2765);
nand U695 (N_695,In_2620,In_1735);
or U696 (N_696,In_3381,In_2132);
xnor U697 (N_697,In_2055,In_4588);
or U698 (N_698,In_4118,In_195);
or U699 (N_699,In_4014,In_875);
and U700 (N_700,In_1751,In_36);
nor U701 (N_701,In_1451,In_3533);
nor U702 (N_702,In_1636,In_4689);
nand U703 (N_703,In_3454,In_1946);
nand U704 (N_704,In_1006,In_3576);
xor U705 (N_705,In_2097,In_65);
and U706 (N_706,In_2407,In_2782);
xor U707 (N_707,In_912,In_1418);
nor U708 (N_708,In_3999,In_662);
or U709 (N_709,In_784,In_4530);
xor U710 (N_710,In_3180,In_4762);
nand U711 (N_711,In_4643,In_3498);
or U712 (N_712,In_1439,In_4608);
nor U713 (N_713,In_455,In_3933);
or U714 (N_714,In_4890,In_3258);
nor U715 (N_715,In_3117,In_4892);
xnor U716 (N_716,In_4385,In_4462);
or U717 (N_717,In_2189,In_4975);
and U718 (N_718,In_4204,In_3475);
nand U719 (N_719,In_1417,In_2594);
and U720 (N_720,In_868,In_4471);
xor U721 (N_721,In_1211,In_2951);
and U722 (N_722,In_3237,In_953);
nand U723 (N_723,In_2612,In_3255);
nand U724 (N_724,In_1976,In_4321);
or U725 (N_725,In_1438,In_4296);
nor U726 (N_726,In_2629,In_2543);
and U727 (N_727,In_1910,In_942);
nand U728 (N_728,In_3639,In_2493);
or U729 (N_729,In_3651,In_2964);
or U730 (N_730,In_1990,In_1614);
and U731 (N_731,In_1838,In_962);
nand U732 (N_732,In_2538,In_2816);
xor U733 (N_733,In_1588,In_3844);
xor U734 (N_734,In_2335,In_1755);
or U735 (N_735,In_2821,In_2344);
nand U736 (N_736,In_1889,In_2191);
or U737 (N_737,In_2176,In_2932);
and U738 (N_738,In_3670,In_3373);
and U739 (N_739,In_4100,In_4609);
xnor U740 (N_740,In_3361,In_2475);
nand U741 (N_741,In_3797,In_4026);
or U742 (N_742,In_3920,In_4676);
xor U743 (N_743,In_3074,In_3148);
and U744 (N_744,In_4666,In_4461);
nor U745 (N_745,In_734,In_1599);
xor U746 (N_746,In_3217,In_1729);
xor U747 (N_747,In_4561,In_1034);
xnor U748 (N_748,In_3311,In_2326);
or U749 (N_749,In_225,In_1251);
or U750 (N_750,In_4516,In_1825);
nand U751 (N_751,In_4942,In_4657);
nand U752 (N_752,In_1384,In_1028);
xor U753 (N_753,In_3187,In_3369);
nand U754 (N_754,In_2701,In_4691);
or U755 (N_755,In_2435,In_1236);
nor U756 (N_756,In_343,In_3225);
nor U757 (N_757,In_4398,In_4545);
xnor U758 (N_758,In_398,In_4243);
and U759 (N_759,In_2159,In_4216);
and U760 (N_760,In_775,In_936);
or U761 (N_761,In_1383,In_3274);
or U762 (N_762,In_4777,In_4144);
nor U763 (N_763,In_847,In_2023);
or U764 (N_764,In_3375,In_3466);
nor U765 (N_765,In_2861,In_93);
xor U766 (N_766,In_3358,In_753);
xor U767 (N_767,In_2348,In_4910);
or U768 (N_768,In_3509,In_2252);
and U769 (N_769,In_4509,In_3232);
or U770 (N_770,In_4940,In_2472);
and U771 (N_771,In_864,In_64);
xor U772 (N_772,In_4880,In_203);
or U773 (N_773,In_505,In_4347);
and U774 (N_774,In_669,In_422);
nor U775 (N_775,In_1415,In_3825);
xnor U776 (N_776,In_4361,In_1591);
or U777 (N_777,In_4327,In_1680);
or U778 (N_778,In_4577,In_1196);
nor U779 (N_779,In_145,In_3377);
xor U780 (N_780,In_176,In_2644);
xor U781 (N_781,In_4434,In_130);
and U782 (N_782,In_2977,In_440);
or U783 (N_783,In_4070,In_4421);
or U784 (N_784,In_4368,In_1687);
nor U785 (N_785,In_4301,In_4323);
and U786 (N_786,In_3903,In_3724);
or U787 (N_787,In_2045,In_1443);
nor U788 (N_788,In_3881,In_2945);
nor U789 (N_789,In_851,In_340);
or U790 (N_790,In_2456,In_2423);
nand U791 (N_791,In_4206,In_2202);
nand U792 (N_792,In_4393,In_2632);
nor U793 (N_793,In_538,In_1169);
nor U794 (N_794,In_2109,In_319);
nand U795 (N_795,In_3081,In_4381);
nand U796 (N_796,In_832,In_4085);
nand U797 (N_797,In_2800,In_831);
xor U798 (N_798,In_4004,In_2973);
or U799 (N_799,In_529,In_2526);
and U800 (N_800,In_43,In_2674);
or U801 (N_801,In_4582,In_771);
and U802 (N_802,In_2307,In_2624);
nand U803 (N_803,In_1114,In_4814);
xnor U804 (N_804,In_1594,In_2551);
and U805 (N_805,In_394,In_531);
nand U806 (N_806,In_264,In_4020);
nor U807 (N_807,In_1240,In_2950);
nand U808 (N_808,In_3685,In_1401);
and U809 (N_809,In_97,In_3687);
or U810 (N_810,In_1180,In_2905);
or U811 (N_811,In_4106,In_2842);
nor U812 (N_812,In_1332,In_3319);
nor U813 (N_813,In_1500,In_4264);
or U814 (N_814,In_797,In_4400);
nand U815 (N_815,In_102,In_4864);
or U816 (N_816,In_4612,In_3678);
nor U817 (N_817,In_336,In_2070);
nor U818 (N_818,In_518,In_3201);
xnor U819 (N_819,In_3349,In_3883);
nand U820 (N_820,In_1997,In_1721);
nor U821 (N_821,In_1864,In_2295);
nor U822 (N_822,In_3046,In_2192);
xnor U823 (N_823,In_699,In_4857);
nand U824 (N_824,In_4445,In_4499);
or U825 (N_825,In_2001,In_337);
and U826 (N_826,In_3948,In_2103);
nor U827 (N_827,In_4757,In_2778);
or U828 (N_828,In_614,In_2712);
nand U829 (N_829,In_4784,In_107);
xor U830 (N_830,In_1020,In_1757);
xor U831 (N_831,In_3320,In_1110);
and U832 (N_832,In_386,In_2417);
nand U833 (N_833,In_1377,In_217);
or U834 (N_834,In_2488,In_3592);
xor U835 (N_835,In_3939,In_4917);
nor U836 (N_836,In_1505,In_1314);
xnor U837 (N_837,In_3347,In_819);
or U838 (N_838,In_2756,In_3292);
xor U839 (N_839,In_1286,In_2912);
nor U840 (N_840,In_2561,In_809);
xor U841 (N_841,In_3064,In_938);
or U842 (N_842,In_1239,In_3768);
nor U843 (N_843,In_1182,In_3393);
xor U844 (N_844,In_1986,In_1780);
xnor U845 (N_845,In_4463,In_1750);
nor U846 (N_846,In_339,In_2872);
nand U847 (N_847,In_2556,In_300);
xor U848 (N_848,In_2940,In_1366);
nand U849 (N_849,In_1399,In_2687);
and U850 (N_850,In_4711,In_1829);
and U851 (N_851,In_1293,In_470);
or U852 (N_852,In_4078,In_4726);
nor U853 (N_853,In_1466,In_3278);
nand U854 (N_854,In_4602,In_2499);
or U855 (N_855,In_1232,In_48);
or U856 (N_856,In_4999,In_3788);
or U857 (N_857,In_1915,In_3865);
nand U858 (N_858,In_2592,In_1789);
nand U859 (N_859,In_4746,In_601);
or U860 (N_860,In_4389,In_2959);
or U861 (N_861,In_126,In_365);
or U862 (N_862,In_2275,In_285);
nor U863 (N_863,In_1917,In_4865);
nand U864 (N_864,In_4088,In_2743);
xor U865 (N_865,In_3211,In_4138);
nor U866 (N_866,In_782,In_21);
xor U867 (N_867,In_1386,In_3013);
nand U868 (N_868,In_419,In_3054);
nand U869 (N_869,In_3520,In_2186);
xor U870 (N_870,In_4727,In_1176);
nor U871 (N_871,In_1333,In_403);
nor U872 (N_872,In_764,In_4198);
nor U873 (N_873,In_3252,In_1441);
and U874 (N_874,In_1459,In_4126);
nor U875 (N_875,In_1519,In_4252);
xor U876 (N_876,In_2013,In_4491);
nand U877 (N_877,In_3277,In_3542);
and U878 (N_878,In_2649,In_4109);
nor U879 (N_879,In_4266,In_3960);
xnor U880 (N_880,In_4480,In_2145);
or U881 (N_881,In_2623,In_1376);
or U882 (N_882,In_0,In_774);
nor U883 (N_883,In_2451,In_3386);
nand U884 (N_884,In_1315,In_4870);
nand U885 (N_885,In_1373,In_2947);
and U886 (N_886,In_3242,In_90);
and U887 (N_887,In_1381,In_2583);
nor U888 (N_888,In_3923,In_2810);
xnor U889 (N_889,In_4517,In_4422);
or U890 (N_890,In_146,In_3135);
xor U891 (N_891,In_3459,In_863);
xor U892 (N_892,In_1173,In_1852);
nor U893 (N_893,In_4105,In_289);
nor U894 (N_894,In_181,In_4200);
or U895 (N_895,In_651,In_2160);
nand U896 (N_896,In_2095,In_1433);
nand U897 (N_897,In_1192,In_4352);
xor U898 (N_898,In_3372,In_2071);
nor U899 (N_899,In_2848,In_4451);
nor U900 (N_900,In_4922,In_1632);
xor U901 (N_901,In_1713,In_1199);
nor U902 (N_902,In_4423,In_3256);
and U903 (N_903,In_4484,In_3859);
and U904 (N_904,In_144,In_2799);
nor U905 (N_905,In_2380,In_373);
or U906 (N_906,In_2775,In_388);
xnor U907 (N_907,In_4665,In_3025);
nand U908 (N_908,In_2748,In_3895);
and U909 (N_909,In_2149,In_3408);
and U910 (N_910,In_598,In_4559);
and U911 (N_911,In_3516,In_1775);
nor U912 (N_912,In_2185,In_4574);
and U913 (N_913,In_4581,In_1833);
and U914 (N_914,In_2866,In_3901);
or U915 (N_915,In_1464,In_3136);
xnor U916 (N_916,In_297,In_2610);
nand U917 (N_917,In_4348,In_2746);
xor U918 (N_918,In_2787,In_2056);
nor U919 (N_919,In_1347,In_1281);
or U920 (N_920,In_2619,In_4383);
or U921 (N_921,In_3676,In_2749);
and U922 (N_922,In_2835,In_4850);
nor U923 (N_923,In_588,In_3404);
xnor U924 (N_924,In_1901,In_1001);
nor U925 (N_925,In_2791,In_397);
nand U926 (N_926,In_3205,In_2759);
and U927 (N_927,In_4732,In_428);
or U928 (N_928,In_3223,In_2802);
nand U929 (N_929,In_2958,In_622);
or U930 (N_930,In_654,In_1823);
or U931 (N_931,In_2359,In_3218);
nand U932 (N_932,In_345,In_331);
xnor U933 (N_933,In_2422,In_694);
xor U934 (N_934,In_2302,In_3596);
and U935 (N_935,In_3100,In_3968);
nor U936 (N_936,In_3880,In_4042);
nand U937 (N_937,In_4003,In_4159);
nand U938 (N_938,In_3416,In_932);
or U939 (N_939,In_3147,In_3613);
nand U940 (N_940,In_454,In_1303);
nand U941 (N_941,In_1582,In_3527);
nor U942 (N_942,In_635,In_1539);
or U943 (N_943,In_385,In_1804);
nor U944 (N_944,In_1174,In_1205);
and U945 (N_945,In_3028,In_1390);
nor U946 (N_946,In_3652,In_2837);
xnor U947 (N_947,In_1067,In_2604);
nor U948 (N_948,In_853,In_1941);
and U949 (N_949,In_304,In_2894);
and U950 (N_950,In_3822,In_2304);
or U951 (N_951,In_2550,In_987);
or U952 (N_952,In_3085,In_4375);
xor U953 (N_953,In_715,In_410);
nor U954 (N_954,In_1327,In_3662);
nor U955 (N_955,In_315,In_2143);
and U956 (N_956,In_510,In_3103);
nand U957 (N_957,In_1882,In_4164);
or U958 (N_958,In_998,In_4544);
xor U959 (N_959,In_2534,In_2975);
nand U960 (N_960,In_2038,In_1787);
xnor U961 (N_961,In_105,In_2478);
nor U962 (N_962,In_4059,In_1208);
xor U963 (N_963,In_4050,In_4242);
xor U964 (N_964,In_2470,In_3555);
nor U965 (N_965,In_4045,In_2284);
nor U966 (N_966,In_4091,In_3987);
and U967 (N_967,In_4645,In_1949);
or U968 (N_968,In_2836,In_3870);
nor U969 (N_969,In_180,In_1815);
xor U970 (N_970,In_1014,In_806);
nor U971 (N_971,In_3476,In_3672);
or U972 (N_972,In_380,In_206);
nor U973 (N_973,In_3717,In_2987);
and U974 (N_974,In_4677,In_701);
xor U975 (N_975,In_4218,In_2455);
nor U976 (N_976,In_4409,In_2729);
nor U977 (N_977,In_3206,In_4915);
nand U978 (N_978,In_2122,In_3422);
or U979 (N_979,In_4173,In_1619);
nor U980 (N_980,In_4528,In_4148);
nor U981 (N_981,In_2528,In_555);
and U982 (N_982,In_1982,In_1575);
and U983 (N_983,In_4349,In_3414);
and U984 (N_984,In_2922,In_2278);
xnor U985 (N_985,In_3421,In_3017);
nor U986 (N_986,In_111,In_3744);
or U987 (N_987,In_2175,In_1370);
nand U988 (N_988,In_3402,In_871);
nor U989 (N_989,In_3023,In_4027);
nand U990 (N_990,In_624,In_534);
xor U991 (N_991,In_1802,In_1553);
nand U992 (N_992,In_4785,In_322);
or U993 (N_993,In_947,In_3068);
nor U994 (N_994,In_248,In_2292);
xor U995 (N_995,In_1563,In_2349);
nand U996 (N_996,In_3383,In_661);
or U997 (N_997,In_625,In_252);
nor U998 (N_998,In_4730,In_3007);
or U999 (N_999,In_3243,In_299);
and U1000 (N_1000,In_1133,In_1078);
nand U1001 (N_1001,In_4744,In_4931);
or U1002 (N_1002,In_2364,In_3299);
xnor U1003 (N_1003,N_761,In_3558);
xnor U1004 (N_1004,N_455,In_1821);
or U1005 (N_1005,In_3628,In_4178);
xor U1006 (N_1006,N_914,N_317);
nand U1007 (N_1007,In_1826,N_894);
and U1008 (N_1008,In_1168,In_3234);
xnor U1009 (N_1009,In_4411,In_2899);
nor U1010 (N_1010,In_2773,In_1543);
xor U1011 (N_1011,In_580,N_604);
and U1012 (N_1012,In_1414,In_4694);
xnor U1013 (N_1013,In_267,In_579);
nor U1014 (N_1014,N_89,In_638);
and U1015 (N_1015,In_4834,In_4887);
nand U1016 (N_1016,In_1973,In_1595);
and U1017 (N_1017,In_827,N_346);
nor U1018 (N_1018,In_667,In_2365);
or U1019 (N_1019,N_297,In_3719);
xnor U1020 (N_1020,In_4052,In_1808);
and U1021 (N_1021,In_2331,N_136);
and U1022 (N_1022,In_4222,In_707);
or U1023 (N_1023,In_350,In_4603);
xnor U1024 (N_1024,N_812,N_869);
xor U1025 (N_1025,In_3512,In_447);
nand U1026 (N_1026,N_359,In_3198);
nand U1027 (N_1027,In_3575,In_1017);
nor U1028 (N_1028,In_4758,In_780);
and U1029 (N_1029,In_316,N_755);
and U1030 (N_1030,In_172,In_3113);
nor U1031 (N_1031,N_788,In_1718);
nand U1032 (N_1032,N_548,In_4703);
or U1033 (N_1033,In_452,N_908);
and U1034 (N_1034,In_2432,N_306);
or U1035 (N_1035,N_101,In_3282);
nor U1036 (N_1036,In_1630,In_3186);
xor U1037 (N_1037,N_754,In_2481);
or U1038 (N_1038,In_4260,In_1453);
and U1039 (N_1039,In_46,In_1604);
nor U1040 (N_1040,N_827,N_453);
xor U1041 (N_1041,In_4863,In_742);
xor U1042 (N_1042,In_1658,N_35);
and U1043 (N_1043,In_890,In_4433);
nand U1044 (N_1044,In_4210,N_34);
xor U1045 (N_1045,In_1419,In_4883);
and U1046 (N_1046,N_750,In_119);
xor U1047 (N_1047,N_835,N_656);
nand U1048 (N_1048,N_610,In_3330);
xnor U1049 (N_1049,N_728,In_2420);
nand U1050 (N_1050,In_599,In_3992);
or U1051 (N_1051,N_266,In_1064);
xnor U1052 (N_1052,In_2131,In_3958);
and U1053 (N_1053,In_4929,In_3937);
nand U1054 (N_1054,In_2440,N_106);
nor U1055 (N_1055,N_232,In_3295);
nor U1056 (N_1056,In_2902,N_120);
nand U1057 (N_1057,In_1866,In_1421);
xor U1058 (N_1058,N_857,N_614);
or U1059 (N_1059,In_2167,In_3801);
and U1060 (N_1060,In_3579,In_3165);
or U1061 (N_1061,In_3455,In_3677);
and U1062 (N_1062,In_4981,In_566);
or U1063 (N_1063,In_2486,In_2230);
nand U1064 (N_1064,In_4290,In_2411);
and U1065 (N_1065,In_768,N_860);
and U1066 (N_1066,In_4961,In_3139);
nand U1067 (N_1067,In_1865,In_2918);
and U1068 (N_1068,In_3123,In_3097);
xnor U1069 (N_1069,In_2052,In_1607);
and U1070 (N_1070,N_249,N_37);
and U1071 (N_1071,In_2068,In_2650);
nand U1072 (N_1072,In_1913,In_3525);
xor U1073 (N_1073,In_1618,In_2904);
xor U1074 (N_1074,In_2371,In_4919);
nand U1075 (N_1075,In_630,In_597);
xnor U1076 (N_1076,In_3443,In_4830);
or U1077 (N_1077,In_424,In_3646);
or U1078 (N_1078,In_1810,N_83);
and U1079 (N_1079,In_974,In_4950);
or U1080 (N_1080,In_2670,In_2401);
and U1081 (N_1081,In_2900,N_39);
nand U1082 (N_1082,In_1126,N_131);
and U1083 (N_1083,In_291,In_3146);
or U1084 (N_1084,In_2148,In_4256);
nand U1085 (N_1085,In_1279,In_4733);
nor U1086 (N_1086,N_864,N_85);
and U1087 (N_1087,In_3333,In_1225);
xnor U1088 (N_1088,In_4002,N_344);
or U1089 (N_1089,N_684,In_2030);
xor U1090 (N_1090,In_517,In_1362);
and U1091 (N_1091,N_353,N_183);
xnor U1092 (N_1092,In_2040,N_231);
nor U1093 (N_1093,N_676,N_221);
nand U1094 (N_1094,In_4774,In_3212);
xnor U1095 (N_1095,In_4674,In_867);
and U1096 (N_1096,In_1634,In_1909);
nor U1097 (N_1097,N_688,In_262);
nor U1098 (N_1098,N_822,In_1492);
xnor U1099 (N_1099,In_3767,N_837);
and U1100 (N_1100,In_3753,In_1945);
and U1101 (N_1101,In_925,N_472);
or U1102 (N_1102,In_3701,In_2953);
nor U1103 (N_1103,N_867,In_3792);
nand U1104 (N_1104,N_14,In_1462);
and U1105 (N_1105,In_2930,In_4869);
or U1106 (N_1106,In_3163,In_686);
nand U1107 (N_1107,N_407,In_926);
nand U1108 (N_1108,In_2805,In_2645);
nand U1109 (N_1109,In_844,N_818);
or U1110 (N_1110,In_1087,In_4778);
nand U1111 (N_1111,In_1162,In_3449);
xnor U1112 (N_1112,In_4054,In_4598);
nand U1113 (N_1113,In_3452,In_825);
nand U1114 (N_1114,In_1354,In_66);
nand U1115 (N_1115,N_590,In_2037);
nor U1116 (N_1116,N_710,N_605);
nor U1117 (N_1117,In_3115,In_4824);
nor U1118 (N_1118,In_3411,N_782);
nor U1119 (N_1119,N_151,N_59);
or U1120 (N_1120,In_3431,In_4902);
xor U1121 (N_1121,In_4699,In_4015);
and U1122 (N_1122,In_4477,In_2154);
nor U1123 (N_1123,In_2882,In_1099);
nand U1124 (N_1124,In_3362,In_917);
and U1125 (N_1125,In_3427,N_391);
nor U1126 (N_1126,In_2323,In_1368);
nand U1127 (N_1127,N_110,In_2343);
or U1128 (N_1128,In_3642,In_1792);
nand U1129 (N_1129,In_3314,In_2098);
and U1130 (N_1130,In_730,In_4628);
nor U1131 (N_1131,In_218,In_615);
xor U1132 (N_1132,In_4633,N_795);
nand U1133 (N_1133,In_3839,In_201);
or U1134 (N_1134,In_1975,N_925);
nor U1135 (N_1135,In_1824,In_874);
or U1136 (N_1136,In_1771,In_425);
nand U1137 (N_1137,In_1250,In_2347);
and U1138 (N_1138,In_657,N_288);
or U1139 (N_1139,In_2024,In_2014);
nand U1140 (N_1140,N_916,In_1613);
nor U1141 (N_1141,In_1886,In_2996);
and U1142 (N_1142,In_3050,N_602);
xnor U1143 (N_1143,N_358,In_3647);
xnor U1144 (N_1144,In_3803,N_974);
nand U1145 (N_1145,In_2346,In_4058);
and U1146 (N_1146,In_141,N_663);
nand U1147 (N_1147,In_4205,N_435);
nor U1148 (N_1148,N_703,In_2428);
nand U1149 (N_1149,In_4862,N_920);
nor U1150 (N_1150,In_2999,In_1342);
and U1151 (N_1151,In_3365,N_304);
nor U1152 (N_1152,In_3710,In_3572);
or U1153 (N_1153,In_4490,N_281);
or U1154 (N_1154,In_2128,In_3134);
nand U1155 (N_1155,In_2065,N_592);
or U1156 (N_1156,In_3175,In_3770);
and U1157 (N_1157,In_15,In_3829);
and U1158 (N_1158,In_1666,N_479);
xor U1159 (N_1159,In_4378,In_2936);
nor U1160 (N_1160,N_712,In_421);
nor U1161 (N_1161,N_76,N_163);
and U1162 (N_1162,N_326,In_4277);
or U1163 (N_1163,N_92,N_118);
nor U1164 (N_1164,In_1398,N_253);
or U1165 (N_1165,N_112,In_4781);
nor U1166 (N_1166,In_3133,In_2461);
xnor U1167 (N_1167,N_467,N_899);
xor U1168 (N_1168,In_274,In_655);
nand U1169 (N_1169,N_865,In_4578);
nor U1170 (N_1170,In_3749,In_14);
and U1171 (N_1171,In_2935,In_2036);
nor U1172 (N_1172,In_4886,In_1266);
and U1173 (N_1173,In_4018,In_250);
or U1174 (N_1174,In_845,In_4364);
and U1175 (N_1175,In_4739,In_1523);
and U1176 (N_1176,In_3853,In_278);
or U1177 (N_1177,In_991,In_2373);
xnor U1178 (N_1178,In_4401,N_71);
nand U1179 (N_1179,N_17,N_124);
and U1180 (N_1180,In_642,In_3114);
or U1181 (N_1181,In_3511,In_4299);
nor U1182 (N_1182,In_3005,In_4945);
or U1183 (N_1183,N_157,N_481);
nor U1184 (N_1184,In_2287,In_4743);
or U1185 (N_1185,In_1047,In_261);
nand U1186 (N_1186,N_607,In_719);
or U1187 (N_1187,In_362,N_749);
or U1188 (N_1188,N_600,In_628);
nor U1189 (N_1189,In_992,In_2504);
or U1190 (N_1190,In_1080,In_2755);
xor U1191 (N_1191,In_3043,N_438);
xnor U1192 (N_1192,N_758,In_3360);
nor U1193 (N_1193,N_220,In_1674);
or U1194 (N_1194,In_3487,In_288);
xor U1195 (N_1195,In_4889,In_4555);
or U1196 (N_1196,In_3356,In_4738);
or U1197 (N_1197,N_651,In_4262);
or U1198 (N_1198,N_731,N_216);
and U1199 (N_1199,In_3539,In_1259);
or U1200 (N_1200,In_3195,In_4790);
nand U1201 (N_1201,In_306,In_4712);
or U1202 (N_1202,In_3598,N_978);
and U1203 (N_1203,In_3633,In_4371);
nor U1204 (N_1204,In_4535,In_2218);
xor U1205 (N_1205,In_3080,In_1623);
xnor U1206 (N_1206,N_973,In_4008);
or U1207 (N_1207,In_2362,In_4102);
nor U1208 (N_1208,In_519,In_2285);
and U1209 (N_1209,In_4320,In_1638);
nand U1210 (N_1210,In_2358,In_857);
xnor U1211 (N_1211,In_1951,In_2345);
nand U1212 (N_1212,In_3153,In_2889);
xnor U1213 (N_1213,In_732,N_967);
nand U1214 (N_1214,In_2508,N_342);
xnor U1215 (N_1215,In_1245,In_1685);
nor U1216 (N_1216,N_995,In_3780);
and U1217 (N_1217,In_922,In_736);
xor U1218 (N_1218,In_1479,In_4133);
nor U1219 (N_1219,In_1585,N_179);
nand U1220 (N_1220,In_1094,In_3947);
nand U1221 (N_1221,In_2445,In_2443);
xor U1222 (N_1222,In_446,In_551);
and U1223 (N_1223,In_955,In_477);
nor U1224 (N_1224,In_1733,In_2107);
xnor U1225 (N_1225,N_797,In_3149);
xnor U1226 (N_1226,In_502,In_4143);
nor U1227 (N_1227,In_770,In_2355);
nor U1228 (N_1228,In_1894,In_3056);
nand U1229 (N_1229,In_1790,In_3623);
xor U1230 (N_1230,N_635,In_2875);
or U1231 (N_1231,In_4729,In_3016);
nor U1232 (N_1232,N_982,N_31);
and U1233 (N_1233,In_3398,In_3914);
nor U1234 (N_1234,In_4356,In_2011);
or U1235 (N_1235,In_3627,In_2794);
or U1236 (N_1236,N_493,In_1890);
or U1237 (N_1237,In_1932,N_652);
nand U1238 (N_1238,In_4637,In_4403);
and U1239 (N_1239,In_1271,In_1646);
nand U1240 (N_1240,In_486,N_128);
xor U1241 (N_1241,In_2726,In_2675);
xor U1242 (N_1242,In_3935,In_4974);
nand U1243 (N_1243,N_764,In_2553);
nor U1244 (N_1244,In_4664,In_2141);
nand U1245 (N_1245,N_1,In_3925);
nor U1246 (N_1246,In_4215,In_2634);
or U1247 (N_1247,N_989,N_347);
nand U1248 (N_1248,N_903,In_2330);
xnor U1249 (N_1249,In_616,In_1899);
xnor U1250 (N_1250,N_971,In_1204);
or U1251 (N_1251,In_1683,N_148);
nand U1252 (N_1252,In_4120,N_813);
or U1253 (N_1253,In_3854,In_4379);
or U1254 (N_1254,In_140,In_2822);
xnor U1255 (N_1255,N_611,N_44);
xnor U1256 (N_1256,N_947,In_1338);
nand U1257 (N_1257,In_2733,In_1066);
or U1258 (N_1258,In_2784,In_4617);
nand U1259 (N_1259,N_91,In_4181);
and U1260 (N_1260,In_54,In_4991);
nor U1261 (N_1261,In_4124,In_954);
or U1262 (N_1262,In_1616,In_4185);
or U1263 (N_1263,In_4900,In_4154);
and U1264 (N_1264,N_489,In_3902);
nor U1265 (N_1265,N_318,In_4081);
nor U1266 (N_1266,In_1788,In_4095);
nor U1267 (N_1267,In_2639,N_631);
or U1268 (N_1268,In_1774,In_3732);
and U1269 (N_1269,In_4620,In_2691);
xor U1270 (N_1270,In_1119,In_2412);
nand U1271 (N_1271,In_1049,In_1763);
xor U1272 (N_1272,In_1597,In_1700);
xor U1273 (N_1273,N_274,In_1863);
nor U1274 (N_1274,In_3078,In_3599);
xnor U1275 (N_1275,In_1867,N_598);
nand U1276 (N_1276,N_494,In_3490);
and U1277 (N_1277,In_1344,N_936);
nand U1278 (N_1278,In_1213,N_441);
or U1279 (N_1279,In_3413,N_445);
or U1280 (N_1280,N_508,In_3641);
nor U1281 (N_1281,In_4410,In_3589);
nand U1282 (N_1282,In_1773,In_1502);
nor U1283 (N_1283,In_3052,In_1806);
nor U1284 (N_1284,In_4166,N_349);
xor U1285 (N_1285,In_4456,In_4169);
nand U1286 (N_1286,In_393,In_1264);
or U1287 (N_1287,In_4151,N_501);
nand U1288 (N_1288,N_82,In_3957);
or U1289 (N_1289,In_4273,N_307);
or U1290 (N_1290,In_4876,In_1966);
or U1291 (N_1291,N_802,In_2809);
or U1292 (N_1292,N_482,In_2780);
nand U1293 (N_1293,In_3996,N_627);
and U1294 (N_1294,In_4055,In_521);
nor U1295 (N_1295,In_3893,In_3382);
xnor U1296 (N_1296,In_3348,In_1324);
nor U1297 (N_1297,In_604,In_2839);
or U1298 (N_1298,In_99,N_310);
xor U1299 (N_1299,In_2890,In_2887);
or U1300 (N_1300,In_2317,N_986);
nand U1301 (N_1301,N_171,In_1444);
xor U1302 (N_1302,N_585,N_437);
nand U1303 (N_1303,In_1352,In_56);
and U1304 (N_1304,In_3863,In_2703);
and U1305 (N_1305,In_688,In_3502);
nor U1306 (N_1306,In_3079,In_308);
and U1307 (N_1307,In_286,In_1075);
nor U1308 (N_1308,In_143,N_889);
nand U1309 (N_1309,N_81,In_27);
xor U1310 (N_1310,In_103,In_861);
or U1311 (N_1311,In_2113,In_4074);
and U1312 (N_1312,In_2819,N_762);
and U1313 (N_1313,In_1644,In_235);
xnor U1314 (N_1314,In_4721,N_457);
nor U1315 (N_1315,N_397,N_242);
or U1316 (N_1316,In_4034,N_855);
or U1317 (N_1317,In_3783,N_256);
or U1318 (N_1318,In_4728,N_660);
nor U1319 (N_1319,In_796,In_767);
nor U1320 (N_1320,In_1925,In_1996);
nor U1321 (N_1321,In_3975,In_4288);
and U1322 (N_1322,In_3497,In_3858);
nand U1323 (N_1323,In_2262,In_3268);
and U1324 (N_1324,In_4325,In_3984);
or U1325 (N_1325,In_981,In_4985);
or U1326 (N_1326,N_569,In_108);
and U1327 (N_1327,In_4615,In_271);
nand U1328 (N_1328,In_1242,In_666);
xor U1329 (N_1329,In_2471,In_1004);
or U1330 (N_1330,In_2116,In_4570);
and U1331 (N_1331,N_531,In_3503);
nor U1332 (N_1332,In_3887,In_4780);
xnor U1333 (N_1333,In_4989,In_272);
nor U1334 (N_1334,N_186,In_3827);
and U1335 (N_1335,In_2886,In_1555);
or U1336 (N_1336,N_897,N_932);
or U1337 (N_1337,In_2818,In_35);
nand U1338 (N_1338,In_4796,In_3543);
or U1339 (N_1339,N_882,In_2562);
xnor U1340 (N_1340,In_1481,In_3787);
nor U1341 (N_1341,In_214,In_3471);
or U1342 (N_1342,In_4258,In_2301);
and U1343 (N_1343,In_2163,N_621);
nand U1344 (N_1344,In_3009,In_4599);
nand U1345 (N_1345,In_3450,In_1837);
and U1346 (N_1346,In_564,In_3334);
xnor U1347 (N_1347,In_3130,In_2789);
nor U1348 (N_1348,N_583,In_1233);
xnor U1349 (N_1349,N_449,N_204);
nand U1350 (N_1350,In_4983,N_144);
and U1351 (N_1351,In_3806,N_715);
xnor U1352 (N_1352,In_2648,In_2990);
xnor U1353 (N_1353,In_1339,In_1363);
and U1354 (N_1354,In_3387,N_972);
xor U1355 (N_1355,In_3981,In_1579);
nor U1356 (N_1356,N_773,N_167);
nand U1357 (N_1357,N_84,In_1970);
and U1358 (N_1358,In_4233,In_4959);
or U1359 (N_1359,N_460,N_706);
xor U1360 (N_1360,In_3355,N_454);
xor U1361 (N_1361,In_540,In_2008);
and U1362 (N_1362,N_362,In_4496);
xnor U1363 (N_1363,In_3847,N_536);
and U1364 (N_1364,In_3451,In_479);
or U1365 (N_1365,N_483,In_1216);
and U1366 (N_1366,In_4235,In_3837);
xor U1367 (N_1367,In_1153,N_841);
nand U1368 (N_1368,In_3742,N_846);
nand U1369 (N_1369,In_2657,N_96);
nor U1370 (N_1370,N_42,In_3557);
nand U1371 (N_1371,In_4066,N_667);
or U1372 (N_1372,In_4748,In_4437);
or U1373 (N_1373,In_1811,In_4232);
and U1374 (N_1374,In_1454,In_2424);
nor U1375 (N_1375,In_2989,In_4502);
nor U1376 (N_1376,N_690,N_57);
and U1377 (N_1377,In_3560,In_3821);
xnor U1378 (N_1378,N_64,In_4819);
nor U1379 (N_1379,In_3716,In_1947);
nand U1380 (N_1380,In_913,In_1786);
or U1381 (N_1381,In_1369,In_4685);
nand U1382 (N_1382,In_3245,In_2763);
or U1383 (N_1383,In_3585,In_2720);
xnor U1384 (N_1384,In_1313,In_1881);
xor U1385 (N_1385,In_418,N_28);
and U1386 (N_1386,N_783,In_3959);
or U1387 (N_1387,In_2909,In_4238);
xor U1388 (N_1388,In_4446,In_116);
nor U1389 (N_1389,In_2446,N_834);
and U1390 (N_1390,In_2088,In_3400);
or U1391 (N_1391,In_3945,N_284);
nor U1392 (N_1392,In_94,In_548);
or U1393 (N_1393,In_805,In_2633);
xnor U1394 (N_1394,In_4117,In_4584);
and U1395 (N_1395,N_988,In_1964);
and U1396 (N_1396,N_733,In_1003);
and U1397 (N_1397,N_294,In_3898);
and U1398 (N_1398,N_518,In_1887);
xnor U1399 (N_1399,In_1921,In_2982);
xor U1400 (N_1400,In_4707,In_4249);
or U1401 (N_1401,In_3666,In_2635);
nand U1402 (N_1402,N_471,N_836);
xor U1403 (N_1403,In_843,In_185);
nand U1404 (N_1404,In_493,In_931);
nor U1405 (N_1405,In_3886,In_4873);
or U1406 (N_1406,In_1843,In_305);
and U1407 (N_1407,In_2824,In_3833);
nor U1408 (N_1408,In_2273,In_4512);
nor U1409 (N_1409,N_142,In_904);
xnor U1410 (N_1410,In_215,N_674);
and U1411 (N_1411,N_431,In_445);
xor U1412 (N_1412,In_4334,In_4670);
or U1413 (N_1413,N_382,In_2671);
nor U1414 (N_1414,In_4572,In_2194);
or U1415 (N_1415,In_3940,N_228);
nand U1416 (N_1416,In_2768,In_1294);
and U1417 (N_1417,N_492,N_259);
nand U1418 (N_1418,In_2385,In_513);
and U1419 (N_1419,In_312,In_3253);
xnor U1420 (N_1420,In_748,In_2734);
and U1421 (N_1421,In_4529,In_1800);
nor U1422 (N_1422,N_201,In_207);
xor U1423 (N_1423,In_3692,In_3897);
xnor U1424 (N_1424,N_56,In_3273);
nor U1425 (N_1425,In_1203,In_1195);
nand U1426 (N_1426,In_1329,In_3456);
nand U1427 (N_1427,N_953,In_1131);
xor U1428 (N_1428,N_504,In_3885);
or U1429 (N_1429,In_3529,In_152);
and U1430 (N_1430,In_3066,In_1387);
or U1431 (N_1431,N_465,In_2796);
and U1432 (N_1432,In_948,In_2220);
nor U1433 (N_1433,In_583,In_2980);
and U1434 (N_1434,In_4855,In_2863);
and U1435 (N_1435,N_466,N_137);
nand U1436 (N_1436,In_2235,In_4475);
nor U1437 (N_1437,In_4183,In_3048);
nor U1438 (N_1438,In_1694,In_5);
xor U1439 (N_1439,In_2769,In_4647);
or U1440 (N_1440,In_2530,N_434);
nand U1441 (N_1441,In_3686,In_4224);
or U1442 (N_1442,In_3817,In_4626);
or U1443 (N_1443,In_3926,N_355);
and U1444 (N_1444,In_2340,In_3298);
nor U1445 (N_1445,In_2738,In_963);
xor U1446 (N_1446,In_2883,In_1457);
xnor U1447 (N_1447,N_245,In_3108);
xnor U1448 (N_1448,In_1392,In_3588);
nand U1449 (N_1449,In_2571,In_3702);
nor U1450 (N_1450,In_2457,In_1961);
or U1451 (N_1451,N_929,In_1304);
nand U1452 (N_1452,N_734,In_1596);
nor U1453 (N_1453,In_1645,N_45);
and U1454 (N_1454,In_311,In_1284);
nor U1455 (N_1455,In_1784,In_478);
and U1456 (N_1456,In_2519,N_994);
or U1457 (N_1457,N_608,In_55);
xnor U1458 (N_1458,In_4426,N_212);
and U1459 (N_1459,In_4938,In_1037);
nand U1460 (N_1460,In_371,In_3630);
nor U1461 (N_1461,N_283,In_668);
xnor U1462 (N_1462,N_478,N_909);
xor U1463 (N_1463,N_992,N_896);
xor U1464 (N_1464,In_405,In_1057);
nand U1465 (N_1465,In_1480,N_50);
or U1466 (N_1466,In_4860,In_3752);
and U1467 (N_1467,N_252,In_3581);
or U1468 (N_1468,In_2476,N_275);
xor U1469 (N_1469,In_349,In_3131);
or U1470 (N_1470,N_302,N_177);
nor U1471 (N_1471,In_3082,In_810);
nand U1472 (N_1472,In_3622,In_2503);
nor U1473 (N_1473,N_282,N_698);
or U1474 (N_1474,N_305,In_2383);
xnor U1475 (N_1475,In_2404,N_2);
nand U1476 (N_1476,In_354,In_4508);
or U1477 (N_1477,In_2942,N_744);
nor U1478 (N_1478,N_215,In_3689);
or U1479 (N_1479,In_3664,In_4500);
xnor U1480 (N_1480,In_1888,In_3505);
or U1481 (N_1481,In_1640,In_3580);
nor U1482 (N_1482,In_2170,In_2322);
nand U1483 (N_1483,In_1943,In_575);
nand U1484 (N_1484,In_1422,In_4809);
and U1485 (N_1485,In_4337,In_1340);
xnor U1486 (N_1486,N_890,N_559);
nor U1487 (N_1487,In_3120,In_557);
nor U1488 (N_1488,In_1120,In_3728);
nor U1489 (N_1489,In_3980,N_981);
nor U1490 (N_1490,In_1098,In_1907);
or U1491 (N_1491,In_4827,N_863);
and U1492 (N_1492,N_595,In_1512);
nor U1493 (N_1493,In_4267,N_459);
and U1494 (N_1494,In_2689,In_600);
nor U1495 (N_1495,In_2934,In_4548);
or U1496 (N_1496,In_3745,In_1870);
xor U1497 (N_1497,In_238,In_3251);
xor U1498 (N_1498,N_47,In_1762);
xnor U1499 (N_1499,In_4731,In_618);
xnor U1500 (N_1500,In_2850,In_221);
and U1501 (N_1501,In_1181,In_4619);
xnor U1502 (N_1502,In_3733,In_4505);
nor U1503 (N_1503,In_4845,In_4407);
xor U1504 (N_1504,In_1854,In_2529);
and U1505 (N_1505,In_2716,In_854);
or U1506 (N_1506,In_3834,N_425);
and U1507 (N_1507,N_521,In_7);
nor U1508 (N_1508,In_1060,N_119);
or U1509 (N_1509,In_1152,N_709);
nor U1510 (N_1510,In_672,In_1224);
and U1511 (N_1511,N_276,In_2736);
or U1512 (N_1512,N_99,In_4370);
xor U1513 (N_1513,In_4190,In_1136);
or U1514 (N_1514,N_60,In_204);
xnor U1515 (N_1515,In_3077,In_50);
or U1516 (N_1516,N_447,In_168);
and U1517 (N_1517,In_698,In_3504);
and U1518 (N_1518,In_3500,In_1402);
or U1519 (N_1519,N_700,N_944);
xor U1520 (N_1520,N_792,N_381);
or U1521 (N_1521,In_3907,N_826);
xnor U1522 (N_1522,In_2413,In_678);
nand U1523 (N_1523,In_4747,N_320);
and U1524 (N_1524,In_499,In_4333);
xnor U1525 (N_1525,In_909,N_643);
nor U1526 (N_1526,N_525,N_854);
nand U1527 (N_1527,In_4987,In_3648);
and U1528 (N_1528,In_2351,In_1472);
nand U1529 (N_1529,In_4125,In_4995);
nand U1530 (N_1530,N_286,In_3022);
xor U1531 (N_1531,In_3566,In_873);
nor U1532 (N_1532,In_4041,In_1908);
nor U1533 (N_1533,In_1486,In_3157);
and U1534 (N_1534,In_535,In_1069);
or U1535 (N_1535,N_557,In_3969);
xor U1536 (N_1536,In_1923,In_1059);
nor U1537 (N_1537,N_692,In_4303);
xor U1538 (N_1538,In_1331,In_3831);
nor U1539 (N_1539,N_311,In_3281);
nand U1540 (N_1540,In_3631,In_4696);
and U1541 (N_1541,In_4566,In_2983);
nor U1542 (N_1542,In_1118,N_922);
xor U1543 (N_1543,In_3321,N_32);
nand U1544 (N_1544,In_4001,In_3938);
nand U1545 (N_1545,In_2332,In_659);
nand U1546 (N_1546,In_4709,In_3403);
nand U1547 (N_1547,In_532,In_1356);
nor U1548 (N_1548,In_735,In_1601);
nor U1549 (N_1549,In_28,In_2324);
xnor U1550 (N_1550,In_762,In_2766);
or U1551 (N_1551,In_1536,N_390);
or U1552 (N_1552,In_2418,In_2077);
nand U1553 (N_1553,In_2467,In_23);
nor U1554 (N_1554,In_1409,In_3301);
or U1555 (N_1555,N_568,N_915);
nand U1556 (N_1556,N_161,In_3132);
or U1557 (N_1557,In_4655,In_675);
nand U1558 (N_1558,N_694,In_70);
xnor U1559 (N_1559,In_42,In_4786);
or U1560 (N_1560,In_3864,In_4269);
nand U1561 (N_1561,N_541,N_748);
nand U1562 (N_1562,In_3341,In_4839);
or U1563 (N_1563,In_958,In_3811);
nor U1564 (N_1564,In_2439,In_2086);
nand U1565 (N_1565,N_725,In_516);
or U1566 (N_1566,In_3244,In_3329);
or U1567 (N_1567,In_2280,In_1322);
nand U1568 (N_1568,In_1326,N_250);
or U1569 (N_1569,N_657,In_3316);
nor U1570 (N_1570,N_299,In_4906);
nor U1571 (N_1571,In_3595,In_3658);
nor U1572 (N_1572,In_4686,In_2102);
and U1573 (N_1573,In_3756,In_2080);
xnor U1574 (N_1574,In_3872,N_424);
nor U1575 (N_1575,In_4799,In_2190);
or U1576 (N_1576,N_19,In_3401);
nor U1577 (N_1577,N_243,In_2637);
nor U1578 (N_1578,In_3060,In_1988);
nand U1579 (N_1579,In_1077,In_3055);
xor U1580 (N_1580,In_3679,In_4387);
or U1581 (N_1581,In_2039,N_596);
xor U1582 (N_1582,In_691,In_4276);
xor U1583 (N_1583,In_2402,N_928);
or U1584 (N_1584,In_3604,In_4487);
and U1585 (N_1585,In_619,In_4586);
xor U1586 (N_1586,N_409,In_2642);
nor U1587 (N_1587,In_155,In_1856);
xnor U1588 (N_1588,In_536,In_273);
nand U1589 (N_1589,N_902,In_1518);
nand U1590 (N_1590,In_3761,In_1744);
nor U1591 (N_1591,In_898,In_3694);
xor U1592 (N_1592,In_2678,In_2438);
and U1593 (N_1593,In_743,In_1308);
xnor U1594 (N_1594,N_95,N_399);
nor U1595 (N_1595,In_2727,In_2437);
nand U1596 (N_1596,In_2688,In_3323);
xnor U1597 (N_1597,In_3823,In_2916);
xnor U1598 (N_1598,In_4152,In_2589);
xor U1599 (N_1599,In_85,In_848);
and U1600 (N_1600,In_4005,In_3667);
nand U1601 (N_1601,In_2517,In_1873);
xnor U1602 (N_1602,In_1749,In_175);
nor U1603 (N_1603,In_1554,N_440);
or U1604 (N_1604,In_700,N_885);
nand U1605 (N_1605,In_466,In_1431);
nand U1606 (N_1606,In_2545,In_1467);
xor U1607 (N_1607,N_159,N_969);
nand U1608 (N_1608,In_3324,N_999);
xnor U1609 (N_1609,In_4553,In_1550);
xnor U1610 (N_1610,N_218,In_2860);
nor U1611 (N_1611,In_2857,In_2035);
nand U1612 (N_1612,In_3983,In_456);
and U1613 (N_1613,In_4180,N_436);
xnor U1614 (N_1614,In_4286,N_670);
nor U1615 (N_1615,In_2647,In_1108);
or U1616 (N_1616,In_1010,N_785);
or U1617 (N_1617,In_4245,In_1185);
xnor U1618 (N_1618,In_2783,N_265);
and U1619 (N_1619,In_648,N_990);
nor U1620 (N_1620,In_1957,In_1018);
nand U1621 (N_1621,N_160,N_97);
nand U1622 (N_1622,In_61,In_4357);
xor U1623 (N_1623,N_668,In_2328);
and U1624 (N_1624,N_851,In_2342);
or U1625 (N_1625,In_3474,In_4946);
nor U1626 (N_1626,In_876,In_3779);
and U1627 (N_1627,In_1088,In_3035);
nand U1628 (N_1628,N_791,In_3731);
nand U1629 (N_1629,In_431,N_370);
and U1630 (N_1630,In_3001,N_907);
xnor U1631 (N_1631,In_4338,In_1042);
nor U1632 (N_1632,In_2797,N_589);
or U1633 (N_1633,N_904,In_3794);
or U1634 (N_1634,N_815,N_121);
and U1635 (N_1635,In_1522,In_1408);
nor U1636 (N_1636,In_4976,N_93);
nand U1637 (N_1637,In_754,In_627);
nand U1638 (N_1638,N_199,In_1148);
nor U1639 (N_1639,N_9,In_3750);
or U1640 (N_1640,In_4171,In_2096);
or U1641 (N_1641,In_2357,In_1795);
nand U1642 (N_1642,In_3696,In_3112);
xnor U1643 (N_1643,N_114,In_2399);
xnor U1644 (N_1644,In_4060,N_957);
and U1645 (N_1645,In_2506,N_552);
nand U1646 (N_1646,In_1125,In_3668);
nor U1647 (N_1647,N_832,In_1375);
xnor U1648 (N_1648,N_36,In_3259);
nor U1649 (N_1649,In_3214,In_404);
nor U1650 (N_1650,In_3367,N_72);
nand U1651 (N_1651,In_2715,In_3884);
xnor U1652 (N_1652,In_1590,In_711);
xor U1653 (N_1653,In_2139,In_4973);
xnor U1654 (N_1654,N_868,N_628);
and U1655 (N_1655,In_1031,N_686);
xor U1656 (N_1656,In_4408,N_43);
nor U1657 (N_1657,N_323,N_225);
nor U1658 (N_1658,In_935,In_2677);
or U1659 (N_1659,In_281,In_266);
or U1660 (N_1660,N_235,In_4718);
nor U1661 (N_1661,In_1705,In_2991);
nand U1662 (N_1662,N_650,In_3424);
nand U1663 (N_1663,In_2183,N_513);
nand U1664 (N_1664,In_4283,N_383);
nor U1665 (N_1665,In_4672,N_833);
nor U1666 (N_1666,N_681,In_4540);
and U1667 (N_1667,In_1797,In_2366);
and U1668 (N_1668,In_2104,In_4440);
and U1669 (N_1669,In_4435,In_3565);
or U1670 (N_1670,In_1633,In_3681);
xor U1671 (N_1671,In_996,In_2468);
or U1672 (N_1672,In_4339,In_3640);
nand U1673 (N_1673,In_295,In_866);
nor U1674 (N_1674,N_639,In_2043);
or U1675 (N_1675,N_227,In_3617);
nor U1676 (N_1676,N_222,In_2582);
nand U1677 (N_1677,In_2683,In_47);
or U1678 (N_1678,In_3210,In_2144);
and U1679 (N_1679,In_1403,In_2264);
nor U1680 (N_1680,In_2100,In_1143);
xor U1681 (N_1681,N_98,In_4971);
nor U1682 (N_1682,In_3541,In_2585);
xnor U1683 (N_1683,In_4167,N_843);
or U1684 (N_1684,N_529,N_713);
nor U1685 (N_1685,In_2607,In_4621);
xor U1686 (N_1686,N_470,In_3993);
xnor U1687 (N_1687,In_1434,In_165);
and U1688 (N_1688,In_2318,In_4656);
or U1689 (N_1689,In_3564,N_169);
xor U1690 (N_1690,In_1564,In_793);
nor U1691 (N_1691,In_3522,In_4454);
nor U1692 (N_1692,In_1704,In_1798);
and U1693 (N_1693,In_3286,N_330);
xor U1694 (N_1694,In_2997,N_763);
nor U1695 (N_1695,In_411,N_941);
xnor U1696 (N_1696,In_4251,In_460);
nand U1697 (N_1697,In_2525,In_577);
or U1698 (N_1698,In_4979,In_33);
xnor U1699 (N_1699,In_2051,In_1937);
nor U1700 (N_1700,In_3313,N_280);
and U1701 (N_1701,In_2256,In_4816);
and U1702 (N_1702,In_1079,In_2041);
or U1703 (N_1703,N_942,In_2263);
nor U1704 (N_1704,In_3909,N_133);
nor U1705 (N_1705,In_1664,In_3966);
or U1706 (N_1706,In_491,In_4797);
xnor U1707 (N_1707,In_1316,In_4069);
xor U1708 (N_1708,N_292,N_912);
or U1709 (N_1709,N_682,In_2213);
xnor U1710 (N_1710,In_4590,In_280);
nand U1711 (N_1711,In_138,In_1193);
or U1712 (N_1712,N_849,In_4284);
nor U1713 (N_1713,N_636,In_370);
xnor U1714 (N_1714,N_796,In_1030);
or U1715 (N_1715,In_2532,In_2245);
or U1716 (N_1716,N_830,In_4741);
xnor U1717 (N_1717,In_4533,In_1201);
or U1718 (N_1718,In_3524,In_2646);
and U1719 (N_1719,In_1684,In_4532);
and U1720 (N_1720,In_3774,In_353);
xor U1721 (N_1721,In_4103,In_88);
and U1722 (N_1722,In_3275,N_646);
or U1723 (N_1723,N_5,In_567);
and U1724 (N_1724,N_401,In_2197);
and U1725 (N_1725,N_328,In_4980);
xor U1726 (N_1726,In_1358,In_1484);
and U1727 (N_1727,In_3786,In_1954);
nor U1728 (N_1728,In_2270,N_3);
and U1729 (N_1729,In_3230,In_3272);
nand U1730 (N_1730,In_1282,In_2004);
xor U1731 (N_1731,In_1920,In_3328);
nor U1732 (N_1732,In_2704,N_473);
nor U1733 (N_1733,In_2224,In_697);
and U1734 (N_1734,In_716,In_355);
nor U1735 (N_1735,In_915,In_381);
nor U1736 (N_1736,In_3950,In_3260);
or U1737 (N_1737,N_324,In_1151);
nor U1738 (N_1738,In_1919,In_2907);
xor U1739 (N_1739,In_1371,In_2303);
or U1740 (N_1740,In_1394,In_1617);
xor U1741 (N_1741,In_4162,In_4866);
nor U1742 (N_1742,In_2414,In_2804);
or U1743 (N_1743,N_555,In_1218);
or U1744 (N_1744,In_1046,N_963);
xor U1745 (N_1745,In_951,In_4753);
and U1746 (N_1746,In_4525,N_152);
nand U1747 (N_1747,N_723,In_720);
and U1748 (N_1748,N_29,In_3546);
and U1749 (N_1749,N_366,N_803);
xnor U1750 (N_1750,In_2702,N_516);
and U1751 (N_1751,In_2268,N_285);
nor U1752 (N_1752,In_2243,In_2017);
nand U1753 (N_1753,In_3840,In_1212);
nand U1754 (N_1754,In_2613,In_1612);
or U1755 (N_1755,In_4417,In_3461);
and U1756 (N_1756,In_1903,In_1246);
xor U1757 (N_1757,In_4075,In_2879);
or U1758 (N_1758,In_3090,N_343);
nand U1759 (N_1759,In_3684,In_2020);
or U1760 (N_1760,In_1880,N_626);
nor U1761 (N_1761,In_2161,N_553);
and U1762 (N_1762,In_3145,In_1488);
and U1763 (N_1763,N_503,In_3093);
or U1764 (N_1764,N_214,In_2539);
and U1765 (N_1765,In_3530,In_1113);
xnor U1766 (N_1766,N_462,N_842);
nand U1767 (N_1767,In_3769,In_3279);
nor U1768 (N_1768,In_3391,N_189);
nand U1769 (N_1769,In_3846,In_333);
nor U1770 (N_1770,N_263,In_1933);
or U1771 (N_1771,In_4811,In_4128);
nor U1772 (N_1772,In_3754,N_759);
xnor U1773 (N_1773,In_2334,In_1799);
or U1774 (N_1774,In_3188,In_2590);
nand U1775 (N_1775,In_3644,N_499);
nor U1776 (N_1776,In_1672,In_3183);
and U1777 (N_1777,In_4068,N_586);
and U1778 (N_1778,In_1299,N_202);
xnor U1779 (N_1779,In_3015,N_955);
or U1780 (N_1780,In_91,In_2395);
nand U1781 (N_1781,In_1883,In_4282);
and U1782 (N_1782,In_4108,In_1074);
or U1783 (N_1783,N_884,In_1622);
or U1784 (N_1784,In_3418,In_2938);
xnor U1785 (N_1785,N_426,In_413);
nor U1786 (N_1786,In_3127,In_229);
nand U1787 (N_1787,In_1651,N_140);
or U1788 (N_1788,In_3059,In_807);
or U1789 (N_1789,In_3420,In_3723);
nand U1790 (N_1790,In_4365,In_4427);
nor U1791 (N_1791,In_1150,In_2390);
xor U1792 (N_1792,In_1781,In_4172);
or U1793 (N_1793,In_826,In_4993);
and U1794 (N_1794,In_4567,In_4459);
and U1795 (N_1795,N_450,In_4019);
nand U1796 (N_1796,In_2009,In_1012);
or U1797 (N_1797,In_3339,N_739);
nor U1798 (N_1798,N_798,In_3919);
or U1799 (N_1799,In_737,In_3465);
nor U1800 (N_1800,In_2434,In_4094);
xnor U1801 (N_1801,N_69,In_3250);
xnor U1802 (N_1802,In_2895,N_976);
and U1803 (N_1803,In_3309,N_487);
nand U1804 (N_1804,N_775,In_1312);
or U1805 (N_1805,In_2547,In_3930);
and U1806 (N_1806,N_574,In_2669);
or U1807 (N_1807,In_1139,In_2605);
nand U1808 (N_1808,In_1850,N_143);
nand U1809 (N_1809,In_3715,In_920);
nand U1810 (N_1810,N_429,In_4234);
and U1811 (N_1811,In_2151,In_4424);
nor U1812 (N_1812,N_334,In_2792);
and U1813 (N_1813,In_400,In_4737);
or U1814 (N_1814,In_222,In_1158);
nand U1815 (N_1815,In_2914,In_469);
or U1816 (N_1816,N_193,In_2169);
and U1817 (N_1817,In_4031,In_1189);
or U1818 (N_1818,In_4788,In_4040);
xnor U1819 (N_1819,In_1938,In_2090);
xnor U1820 (N_1820,In_977,In_1219);
and U1821 (N_1821,In_3229,N_594);
xor U1822 (N_1822,In_664,In_4202);
xor U1823 (N_1823,In_1184,In_1922);
or U1824 (N_1824,In_100,N_23);
nor U1825 (N_1825,N_393,In_3709);
nor U1826 (N_1826,In_3682,In_1891);
nand U1827 (N_1827,N_113,In_1045);
xor U1828 (N_1828,N_778,N_831);
nand U1829 (N_1829,In_4077,In_4279);
and U1830 (N_1830,In_361,In_3419);
nor U1831 (N_1831,In_3266,In_727);
xor U1832 (N_1832,N_261,In_1504);
xor U1833 (N_1833,N_774,In_2565);
or U1834 (N_1834,In_2931,N_194);
and U1835 (N_1835,In_453,N_273);
xor U1836 (N_1836,N_593,In_4367);
and U1837 (N_1837,N_55,N_634);
xor U1838 (N_1838,In_2386,N_428);
nand U1839 (N_1839,N_961,In_1128);
or U1840 (N_1840,In_3934,In_778);
xnor U1841 (N_1841,In_2834,In_2981);
xnor U1842 (N_1842,N_580,In_3737);
xnor U1843 (N_1843,In_1353,In_1608);
and U1844 (N_1844,In_3603,In_1024);
or U1845 (N_1845,In_3913,In_899);
and U1846 (N_1846,In_2923,In_3826);
xnor U1847 (N_1847,In_4658,In_3494);
nor U1848 (N_1848,In_3815,In_3061);
nor U1849 (N_1849,In_4575,In_174);
xor U1850 (N_1850,In_158,N_683);
nor U1851 (N_1851,In_761,In_463);
and U1852 (N_1852,N_549,In_4523);
and U1853 (N_1853,N_125,N_823);
xor U1854 (N_1854,In_4760,In_1135);
xor U1855 (N_1855,N_765,N_985);
and U1856 (N_1856,In_459,N_742);
xor U1857 (N_1857,In_4815,In_4562);
or U1858 (N_1858,In_4874,In_4132);
xor U1859 (N_1859,In_1268,N_198);
or U1860 (N_1860,In_916,In_1531);
nor U1861 (N_1861,N_737,In_4923);
nand U1862 (N_1862,N_87,In_644);
nor U1863 (N_1863,In_1009,In_1186);
nor U1864 (N_1864,N_746,In_3484);
or U1865 (N_1865,In_2596,In_4430);
nor U1866 (N_1866,N_181,N_267);
nand U1867 (N_1867,N_16,In_3799);
xor U1868 (N_1868,In_4893,N_781);
or U1869 (N_1869,In_1149,In_1578);
xnor U1870 (N_1870,In_4717,In_2611);
xnor U1871 (N_1871,In_1449,In_1016);
xor U1872 (N_1872,N_351,In_3594);
xor U1873 (N_1873,N_392,N_206);
nor U1874 (N_1874,In_4170,In_1230);
xnor U1875 (N_1875,In_4527,In_177);
and U1876 (N_1876,N_301,N_644);
and U1877 (N_1877,In_2764,In_2463);
xnor U1878 (N_1878,In_1981,In_4953);
or U1879 (N_1879,In_1360,In_4053);
nor U1880 (N_1880,N_801,In_136);
nand U1881 (N_1881,In_829,In_2450);
nor U1882 (N_1882,In_830,In_3300);
and U1883 (N_1883,In_1521,N_430);
nor U1884 (N_1884,In_1701,In_3296);
nor U1885 (N_1885,In_468,In_2381);
xor U1886 (N_1886,N_291,N_987);
and U1887 (N_1887,In_3447,In_2203);
xnor U1888 (N_1888,N_374,In_2089);
and U1889 (N_1889,In_4908,In_2403);
nand U1890 (N_1890,N_495,In_2253);
xor U1891 (N_1891,N_738,In_2998);
xor U1892 (N_1892,In_2354,N_962);
nand U1893 (N_1893,In_1892,In_2498);
or U1894 (N_1894,In_31,In_4667);
nor U1895 (N_1895,N_787,In_1549);
xnor U1896 (N_1896,In_3845,In_892);
and U1897 (N_1897,In_4962,In_2464);
or U1898 (N_1898,In_450,N_874);
nor U1899 (N_1899,In_1379,N_313);
or U1900 (N_1900,In_3170,In_4522);
or U1901 (N_1901,In_2667,In_4514);
nand U1902 (N_1902,N_80,N_70);
nand U1903 (N_1903,In_836,In_3593);
or U1904 (N_1904,In_2540,N_321);
or U1905 (N_1905,In_545,In_1039);
or U1906 (N_1906,In_582,In_3929);
and U1907 (N_1907,N_146,N_325);
or U1908 (N_1908,In_2568,In_4813);
xnor U1909 (N_1909,In_1625,In_1357);
and U1910 (N_1910,In_2762,In_2494);
and U1911 (N_1911,In_148,N_474);
or U1912 (N_1912,In_3759,N_895);
nand U1913 (N_1913,In_210,In_257);
xor U1914 (N_1914,N_845,In_4302);
xnor U1915 (N_1915,N_331,In_2115);
xor U1916 (N_1916,In_1765,In_4568);
or U1917 (N_1917,In_1641,N_939);
nand U1918 (N_1918,In_1091,In_1482);
nand U1919 (N_1919,In_524,In_910);
xnor U1920 (N_1920,N_887,In_1404);
nor U1921 (N_1921,In_2577,In_4795);
or U1922 (N_1922,In_3860,N_427);
nand U1923 (N_1923,In_4897,N_805);
nor U1924 (N_1924,In_882,N_640);
and U1925 (N_1925,In_4036,In_3289);
and U1926 (N_1926,In_1406,In_125);
and U1927 (N_1927,In_449,In_592);
or U1928 (N_1928,In_585,In_2138);
or U1929 (N_1929,In_1530,In_3977);
and U1930 (N_1930,In_3851,In_751);
or U1931 (N_1931,In_1779,In_2668);
nand U1932 (N_1932,In_2694,N_486);
or U1933 (N_1933,In_2251,In_1380);
or U1934 (N_1934,N_707,N_984);
or U1935 (N_1935,N_496,In_254);
nor U1936 (N_1936,In_4740,In_966);
nand U1937 (N_1937,In_1906,In_1221);
or U1938 (N_1938,In_3809,In_1022);
nor U1939 (N_1939,In_1309,In_1072);
nor U1940 (N_1940,In_2913,In_1248);
or U1941 (N_1941,In_3478,In_3238);
or U1942 (N_1942,In_4600,In_3031);
xnor U1943 (N_1943,In_4901,N_946);
xor U1944 (N_1944,In_4826,In_2208);
nor U1945 (N_1945,In_4344,In_63);
or U1946 (N_1946,In_4708,In_3965);
nand U1947 (N_1947,In_4519,In_72);
and U1948 (N_1948,N_200,In_2140);
xor U1949 (N_1949,N_500,In_2053);
nor U1950 (N_1950,In_3304,In_1844);
nand U1951 (N_1951,In_303,In_489);
nor U1952 (N_1952,In_1474,In_387);
or U1953 (N_1953,In_2409,N_878);
nor U1954 (N_1954,In_3556,In_2239);
xnor U1955 (N_1955,In_4131,In_329);
or U1956 (N_1956,N_394,N_675);
nor U1957 (N_1957,N_665,In_4023);
and U1958 (N_1958,In_4265,N_319);
nor U1959 (N_1959,In_1226,N_158);
xnor U1960 (N_1960,In_3673,N_524);
and U1961 (N_1961,N_398,In_4822);
nor U1962 (N_1962,N_380,N_664);
nand U1963 (N_1963,In_416,In_2376);
and U1964 (N_1964,In_940,In_492);
xnor U1965 (N_1965,In_4927,N_386);
xnor U1966 (N_1966,In_1270,In_546);
nand U1967 (N_1967,In_2452,In_3191);
nor U1968 (N_1968,N_463,In_2859);
nand U1969 (N_1969,In_895,N_735);
nand U1970 (N_1970,N_22,N_551);
xnor U1971 (N_1971,In_4029,In_2877);
xnor U1972 (N_1972,N_729,In_2469);
nor U1973 (N_1973,N_771,In_213);
or U1974 (N_1974,In_4662,N_192);
nand U1975 (N_1975,In_3625,N_111);
xnor U1976 (N_1976,In_1455,N_993);
or U1977 (N_1977,In_117,In_4287);
xor U1978 (N_1978,N_213,In_1841);
or U1979 (N_1979,In_3276,In_814);
nor U1980 (N_1980,In_25,In_4972);
and U1981 (N_1981,In_2851,In_1702);
or U1982 (N_1982,In_1526,In_4849);
or U1983 (N_1983,In_1592,N_316);
nand U1984 (N_1984,In_298,In_2480);
nor U1985 (N_1985,In_4916,N_601);
nand U1986 (N_1986,In_2491,In_649);
xnor U1987 (N_1987,In_4918,N_814);
nor U1988 (N_1988,In_4859,In_3932);
nand U1989 (N_1989,N_591,N_439);
and U1990 (N_1990,In_815,In_4013);
and U1991 (N_1991,In_4250,In_828);
nor U1992 (N_1992,In_363,In_1507);
or U1993 (N_1993,In_212,In_3936);
or U1994 (N_1994,In_4652,N_233);
xor U1995 (N_1995,In_4305,N_779);
nor U1996 (N_1996,In_500,In_4763);
nor U1997 (N_1997,N_701,In_607);
nor U1998 (N_1998,In_2572,N_360);
nand U1999 (N_1999,In_3171,N_724);
nand U2000 (N_2000,In_3982,In_2960);
nand U2001 (N_2001,In_4261,N_271);
or U2002 (N_2002,In_4941,In_2000);
nand U2003 (N_2003,N_277,In_2155);
and U2004 (N_2004,N_1267,In_2205);
xor U2005 (N_2005,In_1389,In_4573);
and U2006 (N_2006,N_1286,In_3892);
and U2007 (N_2007,In_412,In_2574);
and U2008 (N_2008,In_4319,In_2379);
nand U2009 (N_2009,In_3342,In_2527);
xor U2010 (N_2010,N_1292,N_880);
nand U2011 (N_2011,N_1554,N_244);
xnor U2012 (N_2012,N_879,In_1111);
and U2013 (N_2013,In_576,In_2067);
nor U2014 (N_2014,In_4715,In_3910);
and U2015 (N_2015,In_1993,N_1716);
nand U2016 (N_2016,N_178,N_1535);
nand U2017 (N_2017,In_1533,In_2901);
nor U2018 (N_2018,In_137,In_279);
nor U2019 (N_2019,In_4012,In_4823);
xnor U2020 (N_2020,N_1972,N_1622);
nor U2021 (N_2021,In_1812,In_4654);
or U2022 (N_2022,In_3989,N_673);
nor U2023 (N_2023,In_4935,N_132);
xnor U2024 (N_2024,N_442,In_3972);
or U2025 (N_2025,In_1513,In_4072);
nand U2026 (N_2026,N_1033,N_1195);
nand U2027 (N_2027,In_3470,In_60);
nor U2028 (N_2028,In_2573,N_168);
nand U2029 (N_2029,N_77,In_4888);
or U2030 (N_2030,In_2833,In_4856);
or U2031 (N_2031,In_1689,N_1547);
or U2032 (N_2032,In_4646,In_3442);
nor U2033 (N_2033,In_522,In_2027);
nand U2034 (N_2034,N_1281,N_998);
xnor U2035 (N_2035,In_1025,N_612);
or U2036 (N_2036,N_1369,N_1326);
nor U2037 (N_2037,N_1934,In_3203);
nor U2038 (N_2038,N_26,In_1283);
nor U2039 (N_2039,In_4428,In_4583);
or U2040 (N_2040,N_1865,In_2699);
and U2041 (N_2041,In_969,In_878);
nor U2042 (N_2042,N_1390,In_508);
or U2043 (N_2043,N_1666,In_4791);
nor U2044 (N_2044,N_711,In_879);
xnor U2045 (N_2045,N_340,N_1166);
nor U2046 (N_2046,N_776,In_1573);
and U2047 (N_2047,In_3501,N_129);
or U2048 (N_2048,N_1780,In_426);
and U2049 (N_2049,N_641,In_2911);
nor U2050 (N_2050,In_1346,N_1600);
nor U2051 (N_2051,N_1084,N_1140);
or U2052 (N_2052,N_1653,In_1746);
nand U2053 (N_2053,In_943,N_385);
or U2054 (N_2054,N_418,In_3586);
nor U2055 (N_2055,In_4722,N_251);
nand U2056 (N_2056,N_1417,In_2680);
nor U2057 (N_2057,N_1688,N_1465);
or U2058 (N_2058,N_75,N_1345);
or U2059 (N_2059,In_2852,N_1901);
and U2060 (N_2060,N_1146,In_4521);
or U2061 (N_2061,N_354,In_4635);
xnor U2062 (N_2062,In_2827,N_1476);
and U2063 (N_2063,In_2120,N_1661);
and U2064 (N_2064,N_1421,N_1889);
or U2065 (N_2065,N_361,N_1516);
xor U2066 (N_2066,N_377,In_2713);
nor U2067 (N_2067,N_1276,In_4457);
or U2068 (N_2068,In_1033,N_1840);
xnor U2069 (N_2069,N_1790,N_1233);
or U2070 (N_2070,N_1815,N_1308);
nor U2071 (N_2071,N_808,N_1518);
nand U2072 (N_2072,In_2719,In_4905);
or U2073 (N_2073,N_54,N_190);
nor U2074 (N_2074,N_671,N_1182);
xor U2075 (N_2075,In_439,N_1223);
xnor U2076 (N_2076,In_3246,In_473);
nor U2077 (N_2077,In_818,N_1114);
and U2078 (N_2078,N_65,In_1626);
nor U2079 (N_2079,In_112,N_1923);
nor U2080 (N_2080,N_1294,N_917);
nand U2081 (N_2081,N_1779,N_1933);
xnor U2082 (N_2082,In_4984,In_2290);
xor U2083 (N_2083,In_789,N_1939);
nand U2084 (N_2084,In_4831,In_1528);
xor U2085 (N_2085,In_4174,N_1279);
nand U2086 (N_2086,N_1966,N_900);
or U2087 (N_2087,In_556,In_3396);
xnor U2088 (N_2088,N_875,N_696);
nor U2089 (N_2089,In_1668,In_2737);
or U2090 (N_2090,N_514,N_1149);
nand U2091 (N_2091,N_810,N_368);
nand U2092 (N_2092,N_1491,N_1925);
nor U2093 (N_2093,In_292,N_848);
and U2094 (N_2094,N_1094,In_1766);
nand U2095 (N_2095,N_1654,In_3781);
nand U2096 (N_2096,In_1393,N_820);
and U2097 (N_2097,N_1976,N_238);
nor U2098 (N_2098,N_1379,In_4443);
and U2099 (N_2099,N_659,In_1134);
or U2100 (N_2100,N_138,N_272);
nor U2101 (N_2101,N_1360,N_7);
nor U2102 (N_2102,In_1000,In_1038);
and U2103 (N_2103,In_186,In_4649);
nor U2104 (N_2104,N_1576,In_1544);
nor U2105 (N_2105,N_1235,N_1499);
and U2106 (N_2106,N_870,N_816);
xnor U2107 (N_2107,In_1984,In_1021);
xor U2108 (N_2108,In_4140,N_1914);
nor U2109 (N_2109,N_1526,In_3399);
and U2110 (N_2110,In_1497,N_1536);
or U2111 (N_2111,In_3951,In_3485);
nand U2112 (N_2112,In_1190,In_4803);
and U2113 (N_2113,In_1450,In_674);
nand U2114 (N_2114,N_768,N_1480);
and U2115 (N_2115,N_421,N_770);
nor U2116 (N_2116,In_530,In_4061);
nor U2117 (N_2117,N_1703,In_498);
nor U2118 (N_2118,N_254,N_90);
and U2119 (N_2119,In_2874,In_2672);
and U2120 (N_2120,In_1832,N_717);
and U2121 (N_2121,In_1188,N_1568);
xor U2122 (N_2122,N_1471,N_333);
nand U2123 (N_2123,N_1960,In_1427);
and U2124 (N_2124,N_1411,In_4071);
or U2125 (N_2125,N_387,N_21);
nand U2126 (N_2126,In_4684,In_4122);
nand U2127 (N_2127,In_3370,N_339);
or U2128 (N_2128,In_2118,In_4943);
or U2129 (N_2129,In_1301,In_4175);
nor U2130 (N_2130,N_662,N_58);
or U2131 (N_2131,N_1642,In_2458);
nand U2132 (N_2132,In_2855,N_924);
or U2133 (N_2133,In_3891,N_1611);
nor U2134 (N_2134,In_4314,In_602);
and U2135 (N_2135,In_777,In_4853);
and U2136 (N_2136,N_208,N_1942);
xor U2137 (N_2137,In_3143,In_4415);
nand U2138 (N_2138,N_1122,In_191);
xor U2139 (N_2139,N_1738,N_1470);
nor U2140 (N_2140,In_1958,In_1348);
xor U2141 (N_2141,In_86,N_422);
or U2142 (N_2142,In_162,N_1340);
nand U2143 (N_2143,In_2333,N_1401);
xnor U2144 (N_2144,In_4956,N_1052);
xor U2145 (N_2145,In_3492,N_1207);
and U2146 (N_2146,In_3855,N_1435);
and U2147 (N_2147,In_2523,N_1228);
and U2148 (N_2148,N_624,In_84);
or U2149 (N_2149,In_3318,In_341);
nand U2150 (N_2150,In_2655,N_1630);
nor U2151 (N_2151,In_2628,In_512);
nor U2152 (N_2152,In_2924,In_4293);
and U2153 (N_2153,N_1724,In_1082);
xor U2154 (N_2154,N_1847,In_2906);
or U2155 (N_2155,In_330,In_2873);
and U2156 (N_2156,N_1561,N_1105);
xor U2157 (N_2157,In_4452,N_217);
and U2158 (N_2158,N_1265,In_2447);
or U2159 (N_2159,In_2535,In_660);
and U2160 (N_2160,In_1420,N_1605);
or U2161 (N_2161,In_713,N_1147);
and U2162 (N_2162,In_4723,In_3661);
nor U2163 (N_2163,In_4604,In_2142);
or U2164 (N_2164,In_3374,N_539);
nand U2165 (N_2165,In_2961,In_1902);
nor U2166 (N_2166,N_704,In_4391);
nor U2167 (N_2167,In_1753,In_897);
and U2168 (N_2168,N_1549,In_3918);
nor U2169 (N_2169,N_309,In_4057);
nand U2170 (N_2170,N_1846,In_1349);
xnor U2171 (N_2171,In_4359,N_116);
and U2172 (N_2172,N_1970,N_1701);
and U2173 (N_2173,N_1479,In_4782);
nand U2174 (N_2174,In_891,In_4761);
or U2175 (N_2175,N_1851,In_3072);
nor U2176 (N_2176,N_1525,N_1538);
xnor U2177 (N_2177,In_384,N_1174);
or U2178 (N_2178,In_2433,N_248);
and U2179 (N_2179,N_1603,In_3931);
nor U2180 (N_2180,In_4384,N_1203);
nor U2181 (N_2181,In_444,In_179);
or U2182 (N_2182,In_4714,N_687);
nand U2183 (N_2183,In_1851,In_2485);
xnor U2184 (N_2184,N_20,N_1287);
or U2185 (N_2185,N_402,N_258);
xnor U2186 (N_2186,N_1577,N_1719);
or U2187 (N_2187,N_777,In_1896);
and U2188 (N_2188,N_1310,In_2943);
and U2189 (N_2189,N_1139,N_1723);
xnor U2190 (N_2190,N_1836,N_858);
nand U2191 (N_2191,In_2598,N_727);
and U2192 (N_2192,In_3491,N_1819);
or U2193 (N_2193,N_1068,In_2730);
nor U2194 (N_2194,N_1800,In_1862);
nor U2195 (N_2195,In_232,N_1322);
and U2196 (N_2196,In_808,In_544);
or U2197 (N_2197,In_1916,In_4376);
and U2198 (N_2198,N_1542,In_1968);
nor U2199 (N_2199,In_1777,N_1284);
nand U2200 (N_2200,N_174,N_1928);
and U2201 (N_2201,In_4611,In_1432);
nand U2202 (N_2202,In_3990,In_1869);
or U2203 (N_2203,N_1615,N_1278);
xor U2204 (N_2204,In_542,In_1814);
or U2205 (N_2205,In_2536,N_977);
xor U2206 (N_2206,N_1989,N_1553);
nand U2207 (N_2207,In_4481,In_1738);
nor U2208 (N_2208,N_817,In_2489);
nor U2209 (N_2209,N_1692,N_1307);
xor U2210 (N_2210,N_1206,In_3423);
and U2211 (N_2211,N_1163,In_1491);
nor U2212 (N_2212,In_1063,In_2288);
nor U2213 (N_2213,N_1381,In_4798);
xor U2214 (N_2214,N_1250,In_4);
or U2215 (N_2215,In_110,N_1606);
nor U2216 (N_2216,N_1291,In_900);
or U2217 (N_2217,In_2135,N_1537);
or U2218 (N_2218,In_1649,N_1355);
xor U2219 (N_2219,N_1132,In_731);
nor U2220 (N_2220,N_1975,N_415);
or U2221 (N_2221,In_705,In_1036);
and U2222 (N_2222,N_1866,N_721);
nand U2223 (N_2223,N_732,In_1679);
nand U2224 (N_2224,N_1672,In_4313);
or U2225 (N_2225,N_1986,N_1468);
nand U2226 (N_2226,In_1739,In_3738);
or U2227 (N_2227,N_184,N_477);
nor U2228 (N_2228,In_1577,In_4678);
nand U2229 (N_2229,In_3904,In_2246);
or U2230 (N_2230,In_1905,In_1351);
or U2231 (N_2231,In_2781,In_4593);
nand U2232 (N_2232,N_1301,In_1247);
nand U2233 (N_2233,N_1757,N_1391);
nor U2234 (N_2234,In_4679,In_4624);
xor U2235 (N_2235,N_807,In_4660);
or U2236 (N_2236,N_1197,N_573);
or U2237 (N_2237,N_1930,In_1317);
xor U2238 (N_2238,N_1359,In_259);
or U2239 (N_2239,N_587,In_348);
or U2240 (N_2240,N_719,N_1073);
and U2241 (N_2241,N_1637,N_376);
nand U2242 (N_2242,In_749,In_4473);
and U2243 (N_2243,In_2786,In_4868);
xnor U2244 (N_2244,In_1761,In_1671);
xnor U2245 (N_2245,In_1785,In_1292);
xor U2246 (N_2246,N_1406,N_1985);
nor U2247 (N_2247,N_352,N_1596);
and U2248 (N_2248,In_4087,N_1208);
xor U2249 (N_2249,N_1969,In_1782);
and U2250 (N_2250,N_67,N_892);
and U2251 (N_2251,In_258,N_1014);
nand U2252 (N_2252,N_1720,In_840);
xnor U2253 (N_2253,In_4702,In_3876);
xor U2254 (N_2254,In_2398,In_703);
nand U2255 (N_2255,N_1978,N_1440);
nand U2256 (N_2256,N_1761,In_4345);
nand U2257 (N_2257,In_2179,In_2777);
xnor U2258 (N_2258,N_1604,In_2831);
or U2259 (N_2259,In_919,N_1474);
nand U2260 (N_2260,In_2093,N_1503);
xor U2261 (N_2261,In_1051,In_2188);
nor U2262 (N_2262,N_1919,N_1380);
and U2263 (N_2263,N_388,In_2061);
xor U2264 (N_2264,N_141,N_1570);
xor U2265 (N_2265,N_336,In_4543);
and U2266 (N_2266,N_669,In_2293);
nor U2267 (N_2267,In_3231,In_436);
xor U2268 (N_2268,In_2062,N_720);
or U2269 (N_2269,In_1026,In_849);
nand U2270 (N_2270,N_1082,N_806);
and U2271 (N_2271,N_956,N_1004);
nand U2272 (N_2272,In_2049,In_135);
and U2273 (N_2273,In_3665,N_1759);
xnor U2274 (N_2274,N_63,N_1735);
and U2275 (N_2275,N_1100,N_1609);
and U2276 (N_2276,N_1798,In_4821);
and U2277 (N_2277,N_1016,N_1261);
nand U2278 (N_2278,In_2971,In_2182);
xnor U2279 (N_2279,In_4745,In_1556);
nand U2280 (N_2280,In_1748,N_975);
nor U2281 (N_2281,N_1714,N_1694);
and U2282 (N_2282,N_581,In_2512);
nand U2283 (N_2283,N_935,In_3140);
or U2284 (N_2284,In_1101,In_3508);
nor U2285 (N_2285,In_4650,N_1224);
xor U2286 (N_2286,N_1253,In_287);
nor U2287 (N_2287,N_699,In_73);
or U2288 (N_2288,In_1364,N_1965);
nor U2289 (N_2289,In_4697,In_608);
nor U2290 (N_2290,In_2641,In_1178);
and U2291 (N_2291,N_1121,In_4431);
or U2292 (N_2292,N_1141,N_1160);
xor U2293 (N_2293,In_2767,In_609);
nor U2294 (N_2294,N_241,N_789);
and U2295 (N_2295,In_596,In_4513);
nand U2296 (N_2296,In_3363,N_1258);
xor U2297 (N_2297,In_4871,N_1677);
nor U2298 (N_2298,In_574,N_1523);
and U2299 (N_2299,N_866,N_1588);
or U2300 (N_2300,In_3857,N_1825);
nand U2301 (N_2301,In_1647,In_858);
nor U2302 (N_2302,In_2944,In_883);
nor U2303 (N_2303,N_1519,In_712);
xnor U2304 (N_2304,In_2864,In_4311);
xnor U2305 (N_2305,In_3219,N_1859);
and U2306 (N_2306,In_1558,In_1460);
and U2307 (N_2307,N_512,N_1240);
and U2308 (N_2308,In_3616,N_130);
xor U2309 (N_2309,N_1597,In_1496);
xor U2310 (N_2310,In_3657,N_1946);
nor U2311 (N_2311,In_4044,N_1656);
nor U2312 (N_2312,In_2754,In_96);
or U2313 (N_2313,N_107,In_4907);
and U2314 (N_2314,In_752,In_1423);
or U2315 (N_2315,N_1992,In_723);
nor U2316 (N_2316,N_337,In_2388);
xnor U2317 (N_2317,In_4382,In_978);
and U2318 (N_2318,N_1487,N_1091);
or U2319 (N_2319,N_853,N_1752);
nor U2320 (N_2320,In_3317,In_3660);
nor U2321 (N_2321,N_1217,N_154);
nand U2322 (N_2322,In_2903,N_1159);
nor U2323 (N_2323,In_163,N_1118);
and U2324 (N_2324,In_1690,In_2338);
xnor U2325 (N_2325,N_432,N_1900);
or U2326 (N_2326,N_1662,In_4913);
xor U2327 (N_2327,In_2124,N_1774);
or U2328 (N_2328,In_2801,N_1682);
or U2329 (N_2329,In_2979,In_3832);
and U2330 (N_2330,N_1438,In_4636);
xor U2331 (N_2331,In_1983,N_1710);
nor U2332 (N_2332,In_1109,In_150);
or U2333 (N_2333,In_3327,In_4156);
and U2334 (N_2334,N_1783,In_3306);
and U2335 (N_2335,In_3852,In_1345);
and U2336 (N_2336,In_1930,In_3118);
nand U2337 (N_2337,In_2111,In_2795);
nand U2338 (N_2338,In_646,N_1575);
xor U2339 (N_2339,In_1410,N_1056);
or U2340 (N_2340,N_1904,In_4928);
or U2341 (N_2341,N_25,In_690);
or U2342 (N_2342,N_1515,In_4661);
nand U2343 (N_2343,N_1070,N_1181);
xnor U2344 (N_2344,N_1612,In_1562);
or U2345 (N_2345,N_1830,N_819);
or U2346 (N_2346,In_611,N_743);
and U2347 (N_2347,N_918,In_3236);
xnor U2348 (N_2348,In_3194,In_746);
nor U2349 (N_2349,N_1886,In_3620);
nand U2350 (N_2350,N_1172,N_1095);
and U2351 (N_2351,In_2728,N_1559);
or U2352 (N_2352,In_4032,In_12);
nand U2353 (N_2353,N_1618,In_3288);
or U2354 (N_2354,N_542,In_4028);
and U2355 (N_2355,N_780,In_3151);
xor U2356 (N_2356,In_1007,In_3407);
nand U2357 (N_2357,In_4768,N_1120);
or U2358 (N_2358,In_4291,N_308);
and U2359 (N_2359,N_905,N_1257);
or U2360 (N_2360,N_1862,N_1348);
and U2361 (N_2361,N_1218,In_1994);
or U2362 (N_2362,N_1241,In_4082);
and U2363 (N_2363,N_1037,In_202);
nand U2364 (N_2364,In_957,In_1396);
xnor U2365 (N_2365,In_2250,In_2271);
nor U2366 (N_2366,In_2978,N_1044);
xnor U2367 (N_2367,N_420,In_233);
nand U2368 (N_2368,In_4047,In_2558);
or U2369 (N_2369,N_677,N_1760);
xnor U2370 (N_2370,N_1221,N_672);
nor U2371 (N_2371,N_1478,N_564);
and U2372 (N_2372,N_1884,In_1468);
nand U2373 (N_2373,In_3944,N_1638);
xnor U2374 (N_2374,In_3269,N_1729);
xnor U2375 (N_2375,In_2078,In_4285);
nand U2376 (N_2376,In_142,In_1853);
nor U2377 (N_2377,N_1329,In_52);
nor U2378 (N_2378,In_982,In_1717);
and U2379 (N_2379,N_1136,N_1717);
nor U2380 (N_2380,In_2225,N_1232);
or U2381 (N_2381,In_3900,In_632);
nor U2382 (N_2382,In_3796,N_1412);
and U2383 (N_2383,In_3075,In_1365);
nor U2384 (N_2384,N_1099,N_1351);
or U2385 (N_2385,In_2969,N_554);
nand U2386 (N_2386,In_3725,N_877);
or U2387 (N_2387,In_894,N_73);
xor U2388 (N_2388,N_538,In_2087);
nand U2389 (N_2389,N_416,In_4592);
or U2390 (N_2390,N_1874,N_246);
xnor U2391 (N_2391,In_1656,In_49);
nor U2392 (N_2392,In_4316,N_1955);
or U2393 (N_2393,N_505,In_2352);
nor U2394 (N_2394,In_884,N_1616);
nor U2395 (N_2395,In_2460,In_1297);
and U2396 (N_2396,N_527,N_784);
and U2397 (N_2397,N_1407,In_2770);
xor U2398 (N_2398,N_268,N_1086);
or U2399 (N_2399,In_3636,N_1442);
or U2400 (N_2400,In_563,N_224);
or U2401 (N_2401,N_940,N_1071);
xnor U2402 (N_2402,N_1051,In_3493);
or U2403 (N_2403,N_1180,In_4688);
or U2404 (N_2404,In_3003,N_303);
xnor U2405 (N_2405,N_1368,In_1089);
and U2406 (N_2406,N_1363,N_1896);
nand U2407 (N_2407,N_563,N_550);
xnor U2408 (N_2408,N_1187,In_3612);
xor U2409 (N_2409,In_881,N_1770);
nor U2410 (N_2410,N_1931,In_4904);
xor U2411 (N_2411,In_2259,In_3597);
or U2412 (N_2412,In_1661,In_1165);
and U2413 (N_2413,In_1465,N_1855);
or U2414 (N_2414,N_1842,N_1444);
nor U2415 (N_2415,In_3850,N_1185);
and U2416 (N_2416,In_2427,In_1660);
nor U2417 (N_2417,In_92,In_1166);
nand U2418 (N_2418,In_3294,N_1626);
or U2419 (N_2419,In_2779,N_745);
xor U2420 (N_2420,N_1303,In_722);
or U2421 (N_2421,N_1234,In_4397);
or U2422 (N_2422,In_3962,N_980);
and U2423 (N_2423,In_1027,In_3563);
or U2424 (N_2424,In_4996,N_1650);
and U2425 (N_2425,N_685,In_2261);
nor U2426 (N_2426,In_2177,In_3610);
xnor U2427 (N_2427,In_1093,In_983);
xnor U2428 (N_2428,N_247,N_1873);
xor U2429 (N_2429,N_926,In_2972);
and U2430 (N_2430,In_3039,N_1011);
or U2431 (N_2431,In_4101,N_1551);
and U2432 (N_2432,N_519,N_809);
nand U2433 (N_2433,In_251,In_2075);
nor U2434 (N_2434,N_1566,In_1707);
nor U2435 (N_2435,N_1385,In_999);
or U2436 (N_2436,In_2069,In_4236);
or U2437 (N_2437,In_3041,In_2949);
and U2438 (N_2438,In_3159,In_441);
and U2439 (N_2439,N_1010,In_245);
xnor U2440 (N_2440,N_1001,In_812);
nor U2441 (N_2441,In_3614,N_678);
nor U2442 (N_2442,In_1445,N_1562);
nand U2443 (N_2443,N_1041,N_1275);
or U2444 (N_2444,In_4735,N_88);
xnor U2445 (N_2445,In_4894,In_2662);
xnor U2446 (N_2446,N_1631,N_582);
nand U2447 (N_2447,N_1003,In_4618);
or U2448 (N_2448,In_1879,N_913);
nor U2449 (N_2449,N_1192,N_1212);
and U2450 (N_2450,N_1959,N_1722);
nor U2451 (N_2451,N_1450,N_1974);
xor U2452 (N_2452,In_952,N_1461);
nor U2453 (N_2453,N_1679,N_1582);
nand U2454 (N_2454,In_2079,In_3040);
and U2455 (N_2455,In_2341,N_1107);
nor U2456 (N_2456,In_2663,N_1602);
nand U2457 (N_2457,In_3109,In_1015);
nor U2458 (N_2458,In_3302,N_86);
nand U2459 (N_2459,N_446,In_3553);
or U2460 (N_2460,N_691,In_183);
nor U2461 (N_2461,In_2954,In_485);
xor U2462 (N_2462,N_927,In_2985);
and U2463 (N_2463,N_40,In_1323);
xor U2464 (N_2464,N_526,In_1874);
and U2465 (N_2465,In_4837,N_850);
and U2466 (N_2466,N_1778,N_1025);
and U2467 (N_2467,In_2522,N_560);
xor U2468 (N_2468,In_4769,In_2579);
or U2469 (N_2469,In_3703,In_3618);
xnor U2470 (N_2470,N_1860,N_1700);
or U2471 (N_2471,In_4227,In_2134);
or U2472 (N_2472,N_1718,N_1336);
xor U2473 (N_2473,In_2267,N_1804);
or U2474 (N_2474,In_129,N_575);
xnor U2475 (N_2475,N_1601,In_1999);
nor U2476 (N_2476,N_1020,N_400);
nor U2477 (N_2477,In_429,N_403);
nor U2478 (N_2478,N_1418,N_1687);
and U2479 (N_2479,N_1364,In_2425);
or U2480 (N_2480,In_3284,In_4241);
nor U2481 (N_2481,N_606,N_1318);
nor U2482 (N_2482,N_1592,In_1868);
or U2483 (N_2483,N_1254,In_4884);
nand U2484 (N_2484,N_1356,In_3712);
or U2485 (N_2485,In_3473,N_1295);
nand U2486 (N_2486,In_1337,In_4725);
or U2487 (N_2487,N_964,In_3956);
or U2488 (N_2488,N_1721,N_653);
nor U2489 (N_2489,In_1243,In_2105);
and U2490 (N_2490,N_979,N_12);
nor U2491 (N_2491,In_1955,In_4090);
or U2492 (N_2492,N_1106,In_3190);
nor U2493 (N_2493,N_1530,N_1222);
xor U2494 (N_2494,In_3208,In_4925);
nor U2495 (N_2495,In_4388,In_4692);
xnor U2496 (N_2496,In_464,N_1987);
xor U2497 (N_2497,N_468,N_570);
or U2498 (N_2498,In_3069,In_2321);
xor U2499 (N_2499,N_859,In_870);
nand U2500 (N_2500,N_1882,In_2820);
nand U2501 (N_2501,N_1373,In_3838);
xnor U2502 (N_2502,N_1127,N_166);
nor U2503 (N_2503,N_1230,N_1617);
nand U2504 (N_2504,In_1697,In_4700);
and U2505 (N_2505,In_3683,N_68);
nand U2506 (N_2506,In_4492,In_2878);
or U2507 (N_2507,N_736,In_2917);
nand U2508 (N_2508,N_1895,In_123);
nor U2509 (N_2509,In_3528,N_350);
nor U2510 (N_2510,In_2393,N_1386);
nand U2511 (N_2511,N_535,In_1231);
xor U2512 (N_2512,N_1484,N_996);
xnor U2513 (N_2513,In_3216,In_3591);
xor U2514 (N_2514,In_3002,N_484);
xnor U2515 (N_2515,In_928,In_645);
or U2516 (N_2516,In_2867,N_203);
or U2517 (N_2517,In_2957,N_1059);
xnor U2518 (N_2518,N_1186,In_3734);
xor U2519 (N_2519,N_1414,N_1319);
and U2520 (N_2520,In_3435,N_1008);
and U2521 (N_2521,In_3955,N_1488);
and U2522 (N_2522,In_1805,N_172);
xnor U2523 (N_2523,In_4724,In_738);
and U2524 (N_2524,N_1482,In_4641);
xor U2525 (N_2525,N_522,In_1568);
nand U2526 (N_2526,N_1891,N_1658);
nand U2527 (N_2527,N_1973,In_2751);
nor U2528 (N_2528,In_1452,N_1466);
and U2529 (N_2529,N_1756,In_3645);
or U2530 (N_2530,In_859,N_46);
or U2531 (N_2531,In_3861,N_1454);
and U2532 (N_2532,N_1881,In_4474);
nand U2533 (N_2533,N_1489,N_537);
xor U2534 (N_2534,In_4350,N_1814);
nor U2535 (N_2535,N_1625,N_1648);
xnor U2536 (N_2536,In_4458,In_344);
and U2537 (N_2537,N_1510,N_1633);
and U2538 (N_2538,N_1259,N_1501);
or U2539 (N_2539,N_1214,N_1990);
or U2540 (N_2540,In_4315,In_396);
and U2541 (N_2541,In_482,In_4982);
xor U2542 (N_2542,In_1234,In_4281);
nand U2543 (N_2543,N_799,N_104);
and U2544 (N_2544,N_811,N_1496);
nor U2545 (N_2545,N_960,N_1090);
and U2546 (N_2546,In_4418,In_3997);
nor U2547 (N_2547,N_1452,In_4872);
and U2548 (N_2548,N_1750,In_2888);
nand U2549 (N_2549,In_1734,N_1272);
nand U2550 (N_2550,In_4274,In_2774);
nand U2551 (N_2551,In_3922,In_2870);
and U2552 (N_2552,In_2695,N_176);
nand U2553 (N_2553,N_1342,N_1505);
xor U2554 (N_2554,N_633,N_1273);
and U2555 (N_2555,In_4330,In_4425);
and U2556 (N_2556,N_1198,N_1864);
or U2557 (N_2557,In_4552,In_1678);
xor U2558 (N_2558,N_1971,N_1337);
nor U2559 (N_2559,In_1429,In_1580);
xor U2560 (N_2560,N_49,In_1681);
or U2561 (N_2561,In_417,In_2110);
or U2562 (N_2562,N_1867,In_2108);
nor U2563 (N_2563,N_1045,N_1256);
or U2564 (N_2564,In_3820,In_1355);
or U2565 (N_2565,In_1244,In_4468);
nand U2566 (N_2566,N_898,In_1440);
nand U2567 (N_2567,In_1062,N_1619);
xnor U2568 (N_2568,In_4775,N_1054);
nand U2569 (N_2569,In_2369,In_2196);
nand U2570 (N_2570,N_1544,N_1164);
nand U2571 (N_2571,In_4668,In_3283);
or U2572 (N_2572,N_180,N_1080);
and U2573 (N_2573,N_66,In_3477);
nor U2574 (N_2574,N_1660,N_769);
and U2575 (N_2575,N_1227,N_1879);
nand U2576 (N_2576,N_226,N_411);
nor U2577 (N_2577,N_1811,In_2963);
and U2578 (N_2578,In_1606,In_591);
nor U2579 (N_2579,N_1175,N_53);
nor U2580 (N_2580,In_4390,N_1517);
nand U2581 (N_2581,In_3119,In_4194);
xnor U2582 (N_2582,In_4891,In_4504);
xnor U2583 (N_2583,In_3071,N_1290);
xnor U2584 (N_2584,In_4146,In_2599);
or U2585 (N_2585,N_1968,N_1154);
xor U2586 (N_2586,N_1772,N_1244);
and U2587 (N_2587,N_1393,In_2946);
xor U2588 (N_2588,N_1088,N_1205);
nand U2589 (N_2589,In_1667,In_3158);
xor U2590 (N_2590,N_1849,N_1196);
nand U2591 (N_2591,In_2698,In_4110);
or U2592 (N_2592,N_1956,In_4526);
or U2593 (N_2593,In_2760,In_1378);
xnor U2594 (N_2594,In_4270,In_2919);
xor U2595 (N_2595,N_6,N_654);
and U2596 (N_2596,In_3385,In_1567);
nor U2597 (N_2597,N_1331,N_544);
xor U2598 (N_2598,N_919,N_1424);
or U2599 (N_2599,N_838,N_1263);
nor U2600 (N_2600,In_1035,N_1170);
or U2601 (N_2601,In_3791,N_906);
or U2602 (N_2602,N_223,In_4184);
xor U2603 (N_2603,In_1950,In_4638);
and U2604 (N_2604,N_205,N_1485);
and U2605 (N_2605,In_2126,In_1485);
nand U2606 (N_2606,In_2015,In_679);
and U2607 (N_2607,In_3193,In_1723);
or U2608 (N_2608,In_803,In_606);
xor U2609 (N_2609,In_4099,In_1191);
and U2610 (N_2610,N_546,In_4534);
nand U2611 (N_2611,In_1527,N_357);
nand U2612 (N_2612,In_2130,N_1274);
nor U2613 (N_2613,In_1476,N_476);
or U2614 (N_2614,In_4644,N_1358);
nor U2615 (N_2615,In_3963,N_1998);
or U2616 (N_2616,In_3877,N_1305);
nor U2617 (N_2617,In_3691,In_2181);
nor U2618 (N_2618,N_1126,N_1076);
xnor U2619 (N_2619,N_404,N_1116);
nand U2620 (N_2620,In_2207,In_3569);
nor U2621 (N_2621,In_1400,N_1216);
xor U2622 (N_2622,In_656,N_490);
xor U2623 (N_2623,In_1138,N_4);
and U2624 (N_2624,In_706,N_117);
and U2625 (N_2625,N_1249,In_2372);
or U2626 (N_2626,N_413,In_2396);
and U2627 (N_2627,N_1243,In_1171);
or U2628 (N_2628,N_1028,N_1808);
nand U2629 (N_2629,In_3240,In_718);
nor U2630 (N_2630,In_1361,N_1853);
xnor U2631 (N_2631,N_1786,N_1740);
and U2632 (N_2632,In_3495,In_2209);
and U2633 (N_2633,N_945,N_48);
and U2634 (N_2634,N_1709,N_1529);
nor U2635 (N_2635,In_3882,In_4675);
and U2636 (N_2636,N_1572,N_1912);
nand U2637 (N_2637,N_1639,In_3721);
or U2638 (N_2638,N_1236,N_1908);
nor U2639 (N_2639,In_3053,In_961);
xnor U2640 (N_2640,N_507,In_4406);
nand U2641 (N_2641,In_26,In_3432);
nor U2642 (N_2642,In_3178,In_680);
or U2643 (N_2643,N_876,In_2812);
and U2644 (N_2644,In_856,N_523);
nor U2645 (N_2645,N_1793,N_1691);
xor U2646 (N_2646,In_1845,In_539);
nor U2647 (N_2647,In_3714,In_4439);
and U2648 (N_2648,In_475,N_62);
nor U2649 (N_2649,In_147,In_192);
and U2650 (N_2650,N_469,N_372);
xor U2651 (N_2651,N_1878,N_565);
nand U2652 (N_2652,In_1611,N_1297);
nand U2653 (N_2653,N_716,In_284);
and U2654 (N_2654,N_498,In_169);
or U2655 (N_2655,N_195,N_1560);
nor U2656 (N_2656,N_375,In_458);
and U2657 (N_2657,N_1892,In_1760);
nand U2658 (N_2658,N_921,In_2739);
and U2659 (N_2659,In_4695,N_1962);
nor U2660 (N_2660,N_1262,In_4324);
xor U2661 (N_2661,N_1455,N_1119);
nand U2662 (N_2662,N_695,N_1850);
and U2663 (N_2663,In_2305,In_1448);
and U2664 (N_2664,N_1967,N_1459);
or U2665 (N_2665,In_178,In_4141);
nor U2666 (N_2666,In_3619,In_81);
xnor U2667 (N_2667,In_1107,N_52);
nand U2668 (N_2668,In_369,In_3521);
nor U2669 (N_2669,N_1823,N_1089);
and U2670 (N_2670,In_53,N_1841);
or U2671 (N_2671,N_1947,In_4742);
nand U2672 (N_2672,N_74,In_4752);
xnor U2673 (N_2673,In_2283,N_433);
xnor U2674 (N_2674,In_725,N_1910);
or U2675 (N_2675,N_419,In_3315);
nand U2676 (N_2676,N_943,In_2282);
nand U2677 (N_2677,N_1269,N_1002);
or U2678 (N_2678,N_562,N_1888);
or U2679 (N_2679,N_804,N_348);
or U2680 (N_2680,N_1382,N_1796);
nor U2681 (N_2681,In_327,N_1728);
xnor U2682 (N_2682,In_855,N_27);
nor U2683 (N_2683,In_1849,N_1657);
nand U2684 (N_2684,In_4771,N_1574);
xnor U2685 (N_2685,In_4966,In_443);
nand U2686 (N_2686,N_1475,N_1453);
xnor U2687 (N_2687,In_1603,In_901);
or U2688 (N_2688,In_171,In_3063);
and U2689 (N_2689,N_1239,In_1663);
or U2690 (N_2690,N_1680,In_2965);
or U2691 (N_2691,In_4851,N_51);
and U2692 (N_2692,In_3816,In_4188);
xor U2693 (N_2693,In_650,N_1917);
nor U2694 (N_2694,In_4193,In_1044);
and U2695 (N_2695,In_2117,In_2898);
xnor U2696 (N_2696,N_1242,N_1248);
nor U2697 (N_2697,N_1781,N_1669);
nand U2698 (N_2698,N_1595,In_474);
nor U2699 (N_2699,N_451,N_1676);
or U2700 (N_2700,In_4836,N_1109);
xor U2701 (N_2701,In_2520,N_1670);
nand U2702 (N_2702,In_2829,N_1567);
and U2703 (N_2703,N_1508,In_4033);
nand U2704 (N_2704,N_1789,In_1828);
xnor U2705 (N_2705,In_4155,N_840);
nand U2706 (N_2706,In_3106,N_1101);
nor U2707 (N_2707,N_705,In_1654);
nor U2708 (N_2708,In_3570,N_597);
nand U2709 (N_2709,In_3941,In_1023);
or U2710 (N_2710,N_1271,In_1897);
and U2711 (N_2711,N_1826,In_1511);
or U2712 (N_2712,N_1110,In_1759);
and U2713 (N_2713,N_1247,N_1607);
or U2714 (N_2714,N_1394,In_3018);
or U2715 (N_2715,In_3430,In_811);
or U2716 (N_2716,N_1457,N_772);
and U2717 (N_2717,N_1695,In_4135);
nor U2718 (N_2718,N_1935,N_1134);
nor U2719 (N_2719,N_1032,N_584);
or U2720 (N_2720,In_156,In_3346);
or U2721 (N_2721,In_3027,N_1668);
nand U2722 (N_2722,In_2926,N_1795);
or U2723 (N_2723,N_1732,In_1210);
nand U2724 (N_2724,In_6,In_4355);
nor U2725 (N_2725,In_1643,In_1209);
nor U2726 (N_2726,N_1171,In_1716);
xnor U2727 (N_2727,N_1469,In_3463);
nor U2728 (N_2728,In_4192,N_1085);
nand U2729 (N_2729,N_365,In_3793);
xor U2730 (N_2730,In_3942,In_2724);
and U2731 (N_2731,N_1225,In_68);
nand U2732 (N_2732,N_1675,In_639);
and U2733 (N_2733,N_412,In_4429);
and U2734 (N_2734,In_3605,In_4968);
nand U2735 (N_2735,N_1995,N_1314);
and U2736 (N_2736,In_4093,In_2692);
or U2737 (N_2737,N_378,In_2531);
and U2738 (N_2738,In_3559,In_173);
nor U2739 (N_2739,In_184,In_3426);
or U2740 (N_2740,In_3177,N_1220);
nand U2741 (N_2741,In_1724,In_4861);
and U2742 (N_2742,In_4331,N_959);
or U2743 (N_2743,In_1263,N_888);
nor U2744 (N_2744,N_1871,N_1473);
xnor U2745 (N_2745,In_3161,In_2595);
or U2746 (N_2746,N_1880,N_260);
and U2747 (N_2747,N_620,N_1699);
xor U2748 (N_2748,N_1193,N_410);
nand U2749 (N_2749,N_332,N_1309);
nor U2750 (N_2750,In_4145,In_4177);
and U2751 (N_2751,N_356,N_1945);
nor U2752 (N_2752,N_534,In_1227);
and U2753 (N_2753,In_3818,N_1046);
nand U2754 (N_2754,N_196,N_609);
nand U2755 (N_2755,N_1027,In_1665);
nor U2756 (N_2756,N_1655,In_3107);
or U2757 (N_2757,N_269,N_13);
xor U2758 (N_2758,In_918,N_954);
nor U2759 (N_2759,In_677,In_3867);
nor U2760 (N_2760,N_1069,In_4681);
and U2761 (N_2761,N_255,N_1338);
or U2762 (N_2762,N_1246,N_881);
xnor U2763 (N_2763,N_1546,In_2772);
nor U2764 (N_2764,In_1200,N_156);
nor U2765 (N_2765,N_1805,N_1835);
and U2766 (N_2766,In_3835,N_1926);
xnor U2767 (N_2767,In_1977,N_1797);
and U2768 (N_2768,N_1477,In_3379);
xnor U2769 (N_2769,N_1036,N_1598);
nor U2770 (N_2770,In_525,In_434);
and U2771 (N_2771,In_1972,N_1321);
nand U2772 (N_2772,In_2129,N_1038);
nor U2773 (N_2773,N_1400,N_293);
nor U2774 (N_2774,N_714,In_1055);
or U2775 (N_2775,N_1252,N_335);
xor U2776 (N_2776,N_1812,N_149);
or U2777 (N_2777,N_1984,N_510);
xor U2778 (N_2778,N_886,N_1376);
nor U2779 (N_2779,N_1374,In_1424);
or U2780 (N_2780,N_1875,In_4594);
or U2781 (N_2781,In_1411,N_502);
or U2782 (N_2782,In_3830,N_444);
and U2783 (N_2783,N_1623,In_433);
nand U2784 (N_2784,In_4119,In_3086);
nor U2785 (N_2785,N_1906,In_1960);
nand U2786 (N_2786,In_2995,In_2064);
nor U2787 (N_2787,N_1361,N_1000);
or U2788 (N_2788,In_3758,In_4158);
xor U2789 (N_2789,N_1293,In_3537);
nor U2790 (N_2790,In_2255,N_396);
nand U2791 (N_2791,In_2709,In_3743);
nor U2792 (N_2792,N_1785,N_1674);
and U2793 (N_2793,N_287,N_1644);
nor U2794 (N_2794,N_1497,N_1981);
xor U2795 (N_2795,N_1636,In_930);
and U2796 (N_2796,In_2152,In_2993);
xor U2797 (N_2797,N_1548,In_1372);
nand U2798 (N_2798,N_1029,N_1277);
and U2799 (N_2799,In_4127,N_1005);
or U2800 (N_2800,N_1938,N_1748);
and U2801 (N_2801,N_219,In_2210);
or U2802 (N_2802,N_1238,In_3359);
nand U2803 (N_2803,In_4682,In_1942);
nor U2804 (N_2804,In_324,In_3766);
nand U2805 (N_2805,In_2735,N_790);
and U2806 (N_2806,In_989,In_2844);
and U2807 (N_2807,N_1833,In_2099);
xnor U2808 (N_2808,In_4021,N_1428);
nand U2809 (N_2809,N_1646,N_185);
or U2810 (N_2810,In_682,In_2974);
xor U2811 (N_2811,In_2310,In_3044);
xor U2812 (N_2812,N_1683,N_1034);
or U2813 (N_2813,N_61,N_1712);
nand U2814 (N_2814,In_4579,N_1168);
and U2815 (N_2815,In_1670,In_1179);
or U2816 (N_2816,N_1521,In_2193);
and U2817 (N_2817,N_264,In_3204);
or U2818 (N_2818,N_1635,In_3142);
or U2819 (N_2819,In_565,N_1705);
nor U2820 (N_2820,N_1219,N_1298);
or U2821 (N_2821,N_517,N_197);
xnor U2822 (N_2822,N_1017,N_757);
and U2823 (N_2823,In_2700,In_2896);
and U2824 (N_2824,N_1613,In_239);
and U2825 (N_2825,N_603,N_315);
or U2826 (N_2826,In_4329,In_356);
nand U2827 (N_2827,In_4149,In_1768);
nor U2828 (N_2828,N_619,N_862);
xor U2829 (N_2829,N_1741,In_4903);
and U2830 (N_2830,In_739,N_952);
or U2831 (N_2831,N_1404,N_844);
nor U2832 (N_2832,N_229,In_1980);
and U2833 (N_2833,N_236,In_4309);
xnor U2834 (N_2834,N_1325,N_458);
nor U2835 (N_2835,N_1200,N_1844);
nand U2836 (N_2836,In_2172,N_1854);
nand U2837 (N_2837,N_1743,In_2325);
xor U2838 (N_2838,N_1983,In_2497);
nand U2839 (N_2839,In_4546,N_718);
or U2840 (N_2840,N_38,N_520);
xor U2841 (N_2841,N_452,In_448);
xor U2842 (N_2842,N_1023,In_833);
nor U2843 (N_2843,In_2660,In_1732);
xnor U2844 (N_2844,N_617,In_1498);
and U2845 (N_2845,In_3303,In_2286);
nand U2846 (N_2846,In_4550,N_1148);
xnor U2847 (N_2847,In_3699,In_781);
xor U2848 (N_2848,N_1563,In_2033);
and U2849 (N_2849,N_1439,N_1067);
nor U2850 (N_2850,N_341,In_509);
and U2851 (N_2851,N_237,In_2026);
nand U2852 (N_2852,In_1691,N_1964);
xor U2853 (N_2853,In_1302,N_1921);
and U2854 (N_2854,In_1229,N_1767);
xor U2855 (N_2855,In_1730,In_154);
or U2856 (N_2856,In_1456,In_4217);
nand U2857 (N_2857,N_1997,N_1820);
or U2858 (N_2858,In_4920,N_1733);
or U2859 (N_2859,In_243,N_588);
nor U2860 (N_2860,In_1318,N_78);
or U2861 (N_2861,In_3584,In_3805);
nor U2862 (N_2862,N_615,In_3807);
xor U2863 (N_2863,In_2459,N_1532);
and U2864 (N_2864,In_4466,N_1583);
nor U2865 (N_2865,N_1788,N_314);
or U2866 (N_2866,N_1493,In_3573);
nand U2867 (N_2867,N_599,N_1145);
nor U2868 (N_2868,In_941,N_1370);
nand U2869 (N_2869,N_1378,N_1285);
or U2870 (N_2870,In_3974,In_79);
xnor U2871 (N_2871,In_3254,In_2586);
nor U2872 (N_2872,N_24,In_515);
or U2873 (N_2873,In_3351,In_3970);
or U2874 (N_2874,N_571,In_2166);
nand U2875 (N_2875,N_528,N_655);
xor U2876 (N_2876,N_1799,In_4373);
or U2877 (N_2877,In_4076,N_1357);
nor U2878 (N_2878,In_4161,N_1155);
or U2879 (N_2879,N_153,N_1150);
or U2880 (N_2880,In_4478,In_2544);
nand U2881 (N_2881,In_865,N_1097);
nor U2882 (N_2882,In_1586,N_1993);
nand U2883 (N_2883,In_4556,In_3795);
and U2884 (N_2884,N_475,In_3615);
or U2885 (N_2885,N_1514,N_1818);
xor U2886 (N_2886,N_1104,In_984);
nor U2887 (N_2887,N_155,In_3548);
or U2888 (N_2888,In_4453,N_1130);
or U2889 (N_2889,N_1031,In_2666);
nor U2890 (N_2890,In_2665,N_891);
and U2891 (N_2891,N_1204,N_578);
nand U2892 (N_2892,N_1664,In_4713);
nand U2893 (N_2893,In_3828,In_4800);
or U2894 (N_2894,In_949,N_1129);
nor U2895 (N_2895,In_3659,N_371);
xor U2896 (N_2896,In_3608,N_1058);
nand U2897 (N_2897,N_991,N_1199);
xnor U2898 (N_2898,N_0,In_4342);
nand U2899 (N_2899,In_9,N_1857);
or U2900 (N_2900,N_1902,In_721);
and U2901 (N_2901,N_1950,N_1977);
nand U2902 (N_2902,N_1915,In_432);
nand U2903 (N_2903,N_1429,N_18);
or U2904 (N_2904,In_3388,N_625);
and U2905 (N_2905,N_1632,N_1838);
and U2906 (N_2906,N_363,N_1827);
nor U2907 (N_2907,In_2838,N_910);
or U2908 (N_2908,N_1824,N_1671);
xnor U2909 (N_2909,N_871,N_1458);
nor U2910 (N_2910,N_1202,N_1922);
nor U2911 (N_2911,N_1334,In_3751);
and U2912 (N_2912,N_1446,N_1349);
nand U2913 (N_2913,N_209,In_2072);
and U2914 (N_2914,In_787,N_1317);
xnor U2915 (N_2915,N_1158,In_4783);
nand U2916 (N_2916,In_3486,In_2054);
nor U2917 (N_2917,In_2893,N_1941);
nor U2918 (N_2918,N_629,N_638);
and U2919 (N_2919,In_256,N_456);
nand U2920 (N_2920,In_4419,In_914);
nor U2921 (N_2921,In_800,N_1280);
and U2922 (N_2922,N_1640,In_1574);
xnor U2923 (N_2923,N_1524,N_1751);
or U2924 (N_2924,N_1111,In_4469);
nand U2925 (N_2925,In_1117,N_506);
and U2926 (N_2926,N_1913,In_1040);
nand U2927 (N_2927,In_760,N_30);
or U2928 (N_2928,N_1434,In_1965);
xnor U2929 (N_2929,In_1058,In_776);
nor U2930 (N_2930,N_1138,In_945);
nor U2931 (N_2931,In_3637,In_3720);
and U2932 (N_2932,In_4832,In_227);
nor U2933 (N_2933,N_1512,In_78);
and U2934 (N_2934,In_1944,N_1463);
nor U2935 (N_2935,N_1447,N_1079);
xnor U2936 (N_2936,In_2732,In_2112);
nand U2937 (N_2937,N_1769,In_1255);
nand U2938 (N_2938,In_3949,In_3510);
nor U2939 (N_2939,In_2741,N_295);
nand U2940 (N_2940,N_1384,N_852);
nand U2941 (N_2941,In_2217,N_1456);
or U2942 (N_2942,N_1948,In_1610);
and U2943 (N_2943,N_1062,In_869);
nor U2944 (N_2944,In_3890,In_4228);
nor U2945 (N_2945,N_1829,N_1684);
xor U2946 (N_2946,N_1545,In_3515);
and U2947 (N_2947,In_3227,In_3184);
nand U2948 (N_2948,In_631,In_629);
or U2949 (N_2949,In_3917,N_1344);
or U2950 (N_2950,In_4614,In_2742);
nand U2951 (N_2951,N_1087,In_4896);
xnor U2952 (N_2952,N_1845,In_4038);
nand U2953 (N_2953,N_1173,In_824);
nor U2954 (N_2954,N_1513,N_1313);
and U2955 (N_2955,N_1260,N_1775);
nor U2956 (N_2956,In_4065,In_3800);
nor U2957 (N_2957,In_4494,N_1663);
or U2958 (N_2958,N_1268,In_1736);
nor U2959 (N_2959,N_1809,N_1135);
xor U2960 (N_2960,N_1897,N_1383);
nand U2961 (N_2961,In_2382,N_173);
or U2962 (N_2962,N_1730,N_485);
nor U2963 (N_2963,N_1584,N_414);
nor U2964 (N_2964,In_2557,N_1299);
and U2965 (N_2965,N_1739,In_1711);
nor U2966 (N_2966,N_230,In_1985);
and U2967 (N_2967,In_3425,In_1935);
nand U2968 (N_2968,N_1861,N_1762);
or U2969 (N_2969,In_4854,N_1961);
nor U2970 (N_2970,In_495,N_1024);
and U2971 (N_2971,N_1422,N_1725);
nand U2972 (N_2972,In_1517,N_1282);
xnor U2973 (N_2973,N_234,N_345);
nand U2974 (N_2974,N_389,In_87);
xnor U2975 (N_2975,In_4960,N_1026);
xnor U2976 (N_2976,In_467,In_790);
nor U2977 (N_2977,In_1652,In_2843);
xor U2978 (N_2978,N_1426,In_1939);
nand U2979 (N_2979,In_2448,In_4852);
nand U2980 (N_2980,In_1699,N_1773);
xnor U2981 (N_2981,In_1217,In_2153);
nand U2982 (N_2982,In_3335,N_997);
nand U2983 (N_2983,In_159,N_1092);
or U2984 (N_2984,N_289,In_1934);
nand U2985 (N_2985,N_257,In_3862);
or U2986 (N_2986,In_2234,In_1898);
or U2987 (N_2987,N_1828,In_2462);
and U2988 (N_2988,N_1460,N_829);
or U2989 (N_2989,In_2195,N_1726);
xor U2990 (N_2990,In_2815,N_145);
xor U2991 (N_2991,N_1237,In_2308);
and U2992 (N_2992,In_372,N_1579);
and U2993 (N_2993,In_2300,In_2029);
nor U2994 (N_2994,In_2652,In_1566);
and U2995 (N_2995,In_4179,N_1988);
nand U2996 (N_2996,In_558,In_1974);
and U2997 (N_2997,N_1433,N_1890);
and U2998 (N_2998,In_1914,N_1893);
or U2999 (N_2999,N_515,In_3547);
xnor U3000 (N_3000,N_2899,N_2260);
or U3001 (N_3001,N_2906,N_135);
nor U3002 (N_3002,In_4489,In_2500);
xor U3003 (N_3003,N_2733,N_1652);
nor U3004 (N_3004,N_2585,In_1043);
or U3005 (N_3005,In_101,In_3927);
or U3006 (N_3006,N_1507,In_4153);
and U3007 (N_3007,N_2111,In_1859);
nand U3008 (N_3008,N_1430,N_2828);
nand U3009 (N_3009,N_1096,In_4444);
nor U3010 (N_3010,N_2890,N_2109);
nand U3011 (N_3011,N_576,N_367);
and U3012 (N_3012,N_1746,N_2724);
and U3013 (N_3013,N_1689,N_2292);
or U3014 (N_3014,In_3638,N_2017);
nor U3015 (N_3015,N_1372,In_4080);
nand U3016 (N_3016,In_382,N_1765);
and U3017 (N_3017,In_1737,In_4318);
nor U3018 (N_3018,In_3257,In_4263);
xor U3019 (N_3019,N_2567,N_2535);
or U3020 (N_3020,In_3019,N_2669);
and U3021 (N_3021,N_645,N_958);
nor U3022 (N_3022,N_2549,N_2168);
xor U3023 (N_3023,N_1316,In_4595);
or U3024 (N_3024,N_2423,N_464);
nand U3025 (N_3025,N_2678,N_1063);
xor U3026 (N_3026,In_2608,In_3998);
xnor U3027 (N_3027,In_1306,In_3600);
xnor U3028 (N_3028,N_1226,In_1547);
nor U3029 (N_3029,In_613,In_260);
nor U3030 (N_3030,N_567,N_2677);
or U3031 (N_3031,N_2758,N_2904);
nand U3032 (N_3032,In_1163,N_1371);
nor U3033 (N_3033,N_1509,N_2058);
nand U3034 (N_3034,In_1963,N_2238);
and U3035 (N_3035,N_1943,N_1634);
and U3036 (N_3036,In_2281,N_2694);
xnor U3037 (N_3037,N_752,N_2499);
nor U3038 (N_3038,N_2033,In_275);
xnor U3039 (N_3039,N_1113,N_2878);
xor U3040 (N_3040,N_1102,N_825);
and U3041 (N_3041,N_1448,N_2310);
nor U3042 (N_3042,In_3747,N_1587);
xnor U3043 (N_3043,In_415,N_2414);
nand U3044 (N_3044,N_2631,N_1123);
xnor U3045 (N_3045,N_1681,N_2096);
and U3046 (N_3046,N_2308,In_3033);
or U3047 (N_3047,N_2161,N_2152);
nor U3048 (N_3048,N_1144,N_1737);
nor U3049 (N_3049,In_4794,N_2075);
xor U3050 (N_3050,N_2916,N_1201);
nor U3051 (N_3051,N_2823,N_147);
xor U3052 (N_3052,N_637,N_730);
nand U3053 (N_3053,N_1231,N_2954);
xnor U3054 (N_3054,N_970,N_373);
nand U3055 (N_3055,N_1397,In_681);
or U3056 (N_3056,In_4825,In_1011);
xnor U3057 (N_3057,N_2520,N_2950);
xnor U3058 (N_3058,N_1049,N_1876);
and U3059 (N_3059,N_2117,N_2540);
nand U3060 (N_3060,N_1117,N_2287);
and U3061 (N_3061,N_480,N_2443);
xnor U3062 (N_3062,N_2449,In_4405);
or U3063 (N_3063,N_2780,N_2440);
or U3064 (N_3064,N_2723,N_2427);
xor U3065 (N_3065,N_1432,In_3653);
nand U3066 (N_3066,N_1431,N_2379);
and U3067 (N_3067,N_2953,In_3540);
and U3068 (N_3068,N_2072,N_1834);
or U3069 (N_3069,N_934,N_103);
or U3070 (N_3070,N_766,N_2660);
or U3071 (N_3071,N_278,N_2180);
nor U3072 (N_3072,N_2131,N_1296);
nand U3073 (N_3073,N_2162,In_3741);
or U3074 (N_3074,N_689,N_2857);
xnor U3075 (N_3075,N_2581,N_2612);
nand U3076 (N_3076,N_2958,N_2995);
xor U3077 (N_3077,N_1918,N_2842);
and U3078 (N_3078,In_3748,N_2836);
or U3079 (N_3079,N_2572,In_4116);
and U3080 (N_3080,N_2138,In_3602);
and U3081 (N_3081,N_2708,N_2876);
nand U3082 (N_3082,In_2711,N_2170);
and U3083 (N_3083,N_2227,N_2590);
nand U3084 (N_3084,N_1868,N_1169);
xnor U3085 (N_3085,N_1937,In_2223);
xnor U3086 (N_3086,In_1156,N_2433);
nand U3087 (N_3087,N_1362,In_4432);
nor U3088 (N_3088,N_2515,N_2425);
xnor U3089 (N_3089,N_2278,N_2177);
xnor U3090 (N_3090,N_2199,N_1586);
and U3091 (N_3091,In_2693,N_2882);
or U3092 (N_3092,N_2392,N_2453);
xnor U3093 (N_3093,N_2862,N_2101);
nor U3094 (N_3094,N_2243,N_2458);
or U3095 (N_3095,N_2785,N_2411);
nand U3096 (N_3096,N_2737,In_2710);
and U3097 (N_3097,N_965,N_2517);
or U3098 (N_3098,N_1936,N_122);
nor U3099 (N_3099,In_3010,N_1492);
or U3100 (N_3100,N_2750,In_653);
nand U3101 (N_3101,N_2040,N_1270);
xor U3102 (N_3102,N_2336,In_4064);
or U3103 (N_3103,In_1305,In_973);
nor U3104 (N_3104,N_2807,N_2468);
xnor U3105 (N_3105,In_4191,N_2455);
nor U3106 (N_3106,N_2060,N_2252);
or U3107 (N_3107,N_2139,In_1893);
nand U3108 (N_3108,N_2580,N_2805);
nor U3109 (N_3109,N_1332,N_165);
or U3110 (N_3110,N_2438,N_1131);
xnor U3111 (N_3111,N_1791,N_2447);
nand U3112 (N_3112,N_2487,N_2948);
xor U3113 (N_3113,N_2969,N_2276);
nand U3114 (N_3114,In_4885,N_630);
nor U3115 (N_3115,N_2229,N_2121);
and U3116 (N_3116,N_1288,N_2790);
and U3117 (N_3117,N_2932,N_622);
or U3118 (N_3118,N_2365,N_2930);
nand U3119 (N_3119,N_2241,N_2706);
or U3120 (N_3120,N_1304,In_821);
or U3121 (N_3121,N_2319,N_793);
xnor U3122 (N_3122,N_2989,In_161);
or U3123 (N_3123,N_2491,N_2735);
and U3124 (N_3124,N_2570,N_2952);
xnor U3125 (N_3125,N_1686,N_211);
nand U3126 (N_3126,N_2142,N_2843);
nor U3127 (N_3127,N_2542,N_1821);
xnor U3128 (N_3128,In_2265,N_1081);
nand U3129 (N_3129,In_839,N_1839);
nor U3130 (N_3130,N_2551,N_1013);
nor U3131 (N_3131,In_3587,N_2573);
nor U3132 (N_3132,N_2130,N_1481);
and U3133 (N_3133,N_2043,N_2657);
and U3134 (N_3134,In_139,N_2456);
xor U3135 (N_3135,In_3995,N_2061);
xor U3136 (N_3136,N_312,N_2010);
or U3137 (N_3137,N_2016,In_13);
nor U3138 (N_3138,N_2406,N_2098);
and U3139 (N_3139,N_2307,N_2064);
or U3140 (N_3140,N_1528,N_2746);
nor U3141 (N_3141,N_210,N_2982);
xnor U3142 (N_3142,N_2193,In_717);
nor U3143 (N_3143,N_2504,N_2335);
nor U3144 (N_3144,N_2321,N_2401);
nand U3145 (N_3145,N_2331,N_1697);
nor U3146 (N_3146,N_2511,N_1905);
or U3147 (N_3147,N_1564,N_2817);
or U3148 (N_3148,N_1015,In_132);
or U3149 (N_3149,N_2004,N_2065);
nor U3150 (N_3150,N_2727,N_1323);
nand U3151 (N_3151,In_1756,N_2159);
and U3152 (N_3152,N_2588,In_2076);
nor U3153 (N_3153,N_2176,N_2645);
xor U3154 (N_3154,N_2956,N_2315);
xor U3155 (N_3155,In_4104,In_1615);
and U3156 (N_3156,N_2407,N_2036);
or U3157 (N_3157,In_4196,In_4998);
nand U3158 (N_3158,In_3763,N_2866);
xor U3159 (N_3159,N_2768,N_930);
and U3160 (N_3160,In_634,N_2402);
nand U3161 (N_3161,N_2689,N_2639);
xnor U3162 (N_3162,N_1410,In_4114);
nand U3163 (N_3163,N_100,N_1074);
xnor U3164 (N_3164,N_2945,N_1124);
nand U3165 (N_3165,N_2211,N_2007);
and U3166 (N_3166,In_2788,In_1692);
nor U3167 (N_3167,N_1870,N_2002);
and U3168 (N_3168,N_1883,N_1832);
nor U3169 (N_3169,N_2085,N_2144);
nor U3170 (N_3170,In_2272,N_2000);
nor U3171 (N_3171,N_2502,N_2671);
nor U3172 (N_3172,N_2701,N_1178);
xor U3173 (N_3173,N_2726,N_2658);
and U3174 (N_3174,N_2963,N_2525);
nor U3175 (N_3175,N_2334,In_3776);
nor U3176 (N_3176,N_532,N_2532);
or U3177 (N_3177,N_2905,In_41);
xnor U3178 (N_3178,N_2314,In_620);
nand U3179 (N_3179,N_1328,N_2789);
or U3180 (N_3180,N_2546,N_2271);
xnor U3181 (N_3181,N_2195,N_658);
and U3182 (N_3182,In_18,In_553);
and U3183 (N_3183,In_1884,N_2595);
and U3184 (N_3184,N_2936,N_2845);
nand U3185 (N_3185,In_2825,N_2451);
xor U3186 (N_3186,N_2145,N_1413);
xnor U3187 (N_3187,N_191,N_2419);
and U3188 (N_3188,N_2739,In_552);
nand U3189 (N_3189,N_2964,N_2998);
or U3190 (N_3190,N_2666,N_679);
nand U3191 (N_3191,N_2943,N_2766);
nor U3192 (N_3192,N_2413,N_1731);
nand U3193 (N_3193,N_2970,N_2086);
or U3194 (N_3194,N_2757,N_2959);
xnor U3195 (N_3195,N_1527,N_937);
nand U3196 (N_3196,N_2891,N_2505);
and U3197 (N_3197,In_2291,N_2119);
and U3198 (N_3198,In_3366,N_1887);
nand U3199 (N_3199,N_2337,N_2333);
nand U3200 (N_3200,In_965,N_2089);
and U3201 (N_3201,N_2924,N_2068);
nand U3202 (N_3202,N_2863,N_2967);
and U3203 (N_3203,In_2868,In_1311);
and U3204 (N_3204,N_2630,N_2960);
xnor U3205 (N_3205,N_2434,N_545);
and U3206 (N_3206,N_1822,In_3675);
nand U3207 (N_3207,N_2695,N_861);
or U3208 (N_3208,N_2566,N_2417);
or U3209 (N_3209,N_1744,N_2593);
nor U3210 (N_3210,In_3978,N_2968);
or U3211 (N_3211,N_1556,N_2264);
nand U3212 (N_3212,In_2187,N_1581);
or U3213 (N_3213,In_1745,N_2731);
xnor U3214 (N_3214,N_2544,N_2233);
and U3215 (N_3215,N_1030,N_115);
and U3216 (N_3216,N_2594,N_2212);
xnor U3217 (N_3217,In_321,N_2338);
nor U3218 (N_3218,N_2776,In_3032);
xnor U3219 (N_3219,N_2272,N_2490);
and U3220 (N_3220,N_1552,N_1794);
nor U3221 (N_3221,N_1416,N_2647);
nand U3222 (N_3222,N_2404,N_1209);
or U3223 (N_3223,N_2095,In_253);
xnor U3224 (N_3224,N_2279,N_2342);
xnor U3225 (N_3225,N_2322,N_2420);
nor U3226 (N_3226,N_1852,In_1335);
and U3227 (N_3227,N_1932,N_1667);
nor U3228 (N_3228,N_108,N_2623);
nor U3229 (N_3229,N_175,N_2760);
nor U3230 (N_3230,N_2600,In_3464);
or U3231 (N_3231,N_2981,N_2340);
xor U3232 (N_3232,N_2054,N_613);
and U3233 (N_3233,In_1822,In_3371);
and U3234 (N_3234,N_751,N_2812);
or U3235 (N_3235,N_2178,N_1451);
and U3236 (N_3236,In_193,N_11);
and U3237 (N_3237,N_2576,In_1272);
and U3238 (N_3238,N_2752,N_2664);
nor U3239 (N_3239,In_3700,N_2734);
nor U3240 (N_3240,In_1090,In_747);
or U3241 (N_3241,In_3746,In_2449);
and U3242 (N_3242,N_2356,N_2318);
and U3243 (N_3243,N_2783,N_1885);
xor U3244 (N_3244,In_3397,N_2381);
nand U3245 (N_3245,In_3824,N_1443);
nor U3246 (N_3246,N_1047,N_2289);
nor U3247 (N_3247,N_1771,N_2556);
and U3248 (N_3248,N_1869,N_2399);
nand U3249 (N_3249,In_1541,In_3871);
and U3250 (N_3250,In_3707,N_2263);
and U3251 (N_3251,N_2545,N_2606);
nor U3252 (N_3252,N_2349,N_2284);
nand U3253 (N_3253,N_2351,N_1704);
or U3254 (N_3254,N_2185,N_2513);
nand U3255 (N_3255,N_1179,N_2224);
nand U3256 (N_3256,In_3517,N_1627);
nor U3257 (N_3257,N_2774,N_2104);
nand U3258 (N_3258,In_2082,N_2885);
or U3259 (N_3259,N_2112,In_3222);
xor U3260 (N_3260,N_2158,N_2787);
xor U3261 (N_3261,N_722,In_4275);
or U3262 (N_3262,N_2568,N_2353);
nor U3263 (N_3263,N_1927,N_2547);
nand U3264 (N_3264,N_1151,N_2872);
xnor U3265 (N_3265,In_2705,In_1388);
xnor U3266 (N_3266,N_1366,N_2853);
or U3267 (N_3267,N_1541,N_2083);
xnor U3268 (N_3268,N_2328,N_2716);
or U3269 (N_3269,N_2320,N_2925);
and U3270 (N_3270,N_1550,N_2803);
nor U3271 (N_3271,In_693,N_2756);
nand U3272 (N_3272,N_2796,N_1713);
nor U3273 (N_3273,N_2929,N_530);
nand U3274 (N_3274,N_2538,In_4115);
nor U3275 (N_3275,N_1367,N_1807);
nor U3276 (N_3276,N_2886,In_496);
or U3277 (N_3277,N_2821,N_2023);
xor U3278 (N_3278,In_944,N_1957);
or U3279 (N_3279,N_127,In_1918);
nand U3280 (N_3280,In_3729,N_2179);
nor U3281 (N_3281,N_2394,N_2865);
xor U3282 (N_3282,N_2509,N_2339);
and U3283 (N_3283,N_79,N_2076);
and U3284 (N_3284,In_1442,In_3384);
nor U3285 (N_3285,In_3429,In_1796);
and U3286 (N_3286,N_2592,N_2079);
or U3287 (N_3287,N_1980,N_2313);
and U3288 (N_3288,In_3084,In_2927);
and U3289 (N_3289,N_1289,N_1949);
nand U3290 (N_3290,In_3875,N_1698);
or U3291 (N_3291,N_2147,N_1659);
nand U3292 (N_3292,N_1580,N_2591);
and U3293 (N_3293,N_1324,N_509);
xor U3294 (N_3294,In_934,N_1050);
nand U3295 (N_3295,N_2745,N_2709);
nor U3296 (N_3296,N_1156,N_2019);
xor U3297 (N_3297,N_2445,N_2743);
xnor U3298 (N_3298,In_4640,In_1320);
nor U3299 (N_3299,In_1794,In_1122);
nor U3300 (N_3300,N_2978,In_4842);
and U3301 (N_3301,N_2316,N_1817);
nand U3302 (N_3302,N_2030,N_2071);
nor U3303 (N_3303,N_2767,N_1143);
or U3304 (N_3304,N_298,N_2245);
and U3305 (N_3305,In_714,N_2028);
or U3306 (N_3306,N_2405,In_3051);
and U3307 (N_3307,N_1387,N_2265);
and U3308 (N_3308,N_2648,N_767);
nand U3309 (N_3309,N_1540,N_2635);
or U3310 (N_3310,In_3499,N_1098);
xor U3311 (N_3311,N_1629,N_1843);
nand U3312 (N_3312,N_1060,In_2350);
or U3313 (N_3313,In_313,N_2685);
and U3314 (N_3314,N_2166,N_1768);
xnor U3315 (N_3315,N_2134,N_2661);
nor U3316 (N_3316,N_2908,N_2942);
nand U3317 (N_3317,In_3514,N_1504);
xor U3318 (N_3318,N_2298,In_979);
nor U3319 (N_3319,In_3460,N_1693);
xnor U3320 (N_3320,N_2081,In_801);
nor U3321 (N_3321,N_2188,In_4951);
xor U3322 (N_3322,In_1742,N_1075);
or U3323 (N_3323,N_2510,In_4807);
nand U3324 (N_3324,N_1066,N_2605);
or U3325 (N_3325,N_2991,N_2983);
nand U3326 (N_3326,N_2911,In_2483);
nand U3327 (N_3327,N_2627,N_2450);
nor U3328 (N_3328,In_2984,N_2385);
xor U3329 (N_3329,N_2364,N_2270);
xnor U3330 (N_3330,N_2962,N_1991);
nand U3331 (N_3331,N_2377,N_2643);
nor U3332 (N_3332,N_2347,In_3708);
nor U3333 (N_3333,In_2226,N_2940);
nor U3334 (N_3334,N_2601,In_3394);
nor U3335 (N_3335,N_2769,N_2692);
nor U3336 (N_3336,N_2831,N_2732);
nor U3337 (N_3337,N_2430,In_3577);
nand U3338 (N_3338,N_2389,N_15);
and U3339 (N_3339,N_2027,N_1464);
nor U3340 (N_3340,N_2558,N_2116);
or U3341 (N_3341,N_1621,In_1706);
xor U3342 (N_3342,N_2879,N_2395);
nand U3343 (N_3343,In_1061,In_2022);
and U3344 (N_3344,N_2775,N_102);
nor U3345 (N_3345,N_2840,N_2375);
or U3346 (N_3346,N_2782,N_2771);
or U3347 (N_3347,N_2688,N_1766);
nand U3348 (N_3348,N_1213,N_2755);
nand U3349 (N_3349,N_2784,N_2437);
nor U3350 (N_3350,In_4476,N_1764);
and U3351 (N_3351,N_2871,In_1948);
nor U3352 (N_3352,N_1315,N_800);
and U3353 (N_3353,N_2654,N_2242);
and U3354 (N_3354,In_3096,In_2248);
xor U3355 (N_3355,N_2469,In_3047);
xnor U3356 (N_3356,N_2175,N_2599);
and U3357 (N_3357,In_4990,N_2999);
nor U3358 (N_3358,N_543,N_405);
nand U3359 (N_3359,N_1565,In_1537);
or U3360 (N_3360,N_2408,N_747);
or U3361 (N_3361,In_804,In_2685);
or U3362 (N_3362,N_1782,N_1498);
and U3363 (N_3363,N_109,In_2653);
or U3364 (N_3364,N_2358,N_2299);
nand U3365 (N_3365,N_423,N_2257);
and U3366 (N_3366,N_2396,N_188);
nand U3367 (N_3367,In_134,N_2720);
or U3368 (N_3368,N_2670,N_2446);
nand U3369 (N_3369,In_4988,N_1255);
and U3370 (N_3370,N_2802,N_2359);
nor U3371 (N_3371,N_2182,N_1792);
nor U3372 (N_3372,N_2503,N_2398);
nand U3373 (N_3373,N_1916,In_2260);
nand U3374 (N_3374,N_1420,N_2136);
nor U3375 (N_3375,N_697,N_2873);
xor U3376 (N_3376,In_1583,N_2917);
nor U3377 (N_3377,N_824,N_2815);
and U3378 (N_3378,N_2014,N_1188);
or U3379 (N_3379,N_1006,N_2051);
nand U3380 (N_3380,N_2204,N_2108);
xnor U3381 (N_3381,N_2779,N_1152);
and U3382 (N_3382,In_2374,N_2258);
or U3383 (N_3383,N_2325,In_4952);
xor U3384 (N_3384,N_2997,N_2749);
nand U3385 (N_3385,N_2149,N_2721);
nand U3386 (N_3386,N_94,N_1531);
and U3387 (N_3387,N_1708,N_2093);
nand U3388 (N_3388,N_2039,N_786);
nand U3389 (N_3389,N_1350,N_1758);
nor U3390 (N_3390,N_1483,In_4438);
or U3391 (N_3391,N_2187,N_1951);
or U3392 (N_3392,In_45,N_2947);
xnor U3393 (N_3393,N_2526,N_2268);
nand U3394 (N_3394,N_1954,N_2624);
or U3395 (N_3395,N_2372,N_239);
and U3396 (N_3396,N_338,In_3239);
nor U3397 (N_3397,In_1096,In_3395);
nand U3398 (N_3398,N_2634,N_2105);
nand U3399 (N_3399,N_2579,In_4136);
nand U3400 (N_3400,N_1353,In_1769);
nor U3401 (N_3401,N_1500,N_2393);
nand U3402 (N_3402,N_1311,N_2067);
xnor U3403 (N_3403,N_2986,N_2818);
and U3404 (N_3404,N_2741,N_2120);
nand U3405 (N_3405,In_196,In_1253);
xor U3406 (N_3406,N_1053,N_1520);
and U3407 (N_3407,In_1682,In_1871);
nor U3408 (N_3408,N_207,N_2849);
and U3409 (N_3409,N_2690,N_2442);
or U3410 (N_3410,In_1172,In_4300);
nand U3411 (N_3411,N_2791,N_2323);
xor U3412 (N_3412,N_2388,N_2009);
xor U3413 (N_3413,In_3621,N_2889);
nor U3414 (N_3414,N_2839,In_4524);
and U3415 (N_3415,N_1065,N_2148);
or U3416 (N_3416,N_2632,In_328);
nor U3417 (N_3417,N_1012,N_1339);
nor U3418 (N_3418,N_2604,N_2683);
xnor U3419 (N_3419,N_2387,N_2584);
nand U3420 (N_3420,N_1522,N_2819);
and U3421 (N_3421,In_1992,N_666);
and U3422 (N_3422,N_2042,N_616);
or U3423 (N_3423,N_680,In_3128);
or U3424 (N_3424,N_1952,N_2100);
xor U3425 (N_3425,N_2516,N_2826);
and U3426 (N_3426,In_3322,In_4765);
xor U3427 (N_3427,N_2291,N_2957);
nand U3428 (N_3428,N_1591,In_1100);
nand U3429 (N_3429,N_1777,N_1251);
or U3430 (N_3430,N_2792,N_2485);
or U3431 (N_3431,N_577,In_3228);
nor U3432 (N_3432,In_3785,In_4160);
nand U3433 (N_3433,N_1555,In_1469);
and U3434 (N_3434,N_2073,N_2834);
nor U3435 (N_3435,N_1903,N_2697);
nand U3436 (N_3436,N_1571,N_2973);
nand U3437 (N_3437,In_4011,In_1731);
or U3438 (N_3438,In_2289,N_2901);
and U3439 (N_3439,N_2903,N_2341);
xor U3440 (N_3440,N_2435,N_648);
nand U3441 (N_3441,N_2975,N_1392);
xnor U3442 (N_3442,N_1673,In_2910);
xnor U3443 (N_3443,N_1831,N_1734);
or U3444 (N_3444,In_1070,N_2744);
nor U3445 (N_3445,N_1837,N_2018);
xnor U3446 (N_3446,N_2448,N_2534);
xor U3447 (N_3447,N_1685,N_968);
xor U3448 (N_3448,N_2705,N_2829);
nand U3449 (N_3449,N_1354,In_4306);
or U3450 (N_3450,N_951,N_901);
nor U3451 (N_3451,In_1858,N_2860);
nand U3452 (N_3452,In_302,N_693);
nand U3453 (N_3453,In_1602,N_2710);
nand U3454 (N_3454,In_623,In_1446);
or U3455 (N_3455,N_2665,N_2519);
or U3456 (N_3456,N_2496,In_3111);
nand U3457 (N_3457,N_2309,N_2919);
nand U3458 (N_3458,N_2077,N_2884);
or U3459 (N_3459,N_2011,In_1269);
xnor U3460 (N_3460,In_2640,N_1283);
and U3461 (N_3461,In_3121,N_2856);
xor U3462 (N_3462,N_2675,In_1330);
or U3463 (N_3463,In_1791,N_1191);
nor U3464 (N_3464,N_2066,N_1963);
nor U3465 (N_3465,N_162,In_2832);
xor U3466 (N_3466,N_2993,In_4808);
nor U3467 (N_3467,N_1229,N_2528);
xnor U3468 (N_3468,N_1920,In_2319);
nor U3469 (N_3469,N_270,N_1641);
or U3470 (N_3470,N_2137,N_1462);
nand U3471 (N_3471,N_2939,In_3911);
and U3472 (N_3472,N_708,N_1009);
xor U3473 (N_3473,N_2707,N_2762);
or U3474 (N_3474,N_760,N_2141);
nand U3475 (N_3475,N_1585,In_1655);
xnor U3476 (N_3476,In_2199,N_2126);
and U3477 (N_3477,N_1620,In_1290);
or U3478 (N_3478,In_4495,N_2459);
xor U3479 (N_3479,N_2808,In_3458);
nand U3480 (N_3480,In_3916,N_2236);
xnor U3481 (N_3481,In_1223,N_2736);
xor U3482 (N_3482,N_2603,In_4693);
nor U3483 (N_3483,N_2877,In_1639);
nand U3484 (N_3484,In_310,In_3440);
or U3485 (N_3485,In_4970,In_3095);
xnor U3486 (N_3486,In_3226,N_2928);
and U3487 (N_3487,N_1194,N_2326);
nand U3488 (N_3488,N_2092,In_391);
xor U3489 (N_3489,In_1295,N_2636);
and U3490 (N_3490,In_2826,N_1055);
nand U3491 (N_3491,N_2114,N_839);
xor U3492 (N_3492,N_1423,N_2467);
nand U3493 (N_3493,In_2387,In_2158);
nor U3494 (N_3494,In_1940,N_395);
xor U3495 (N_3495,N_2422,N_2247);
and U3496 (N_3496,In_993,N_2868);
and U3497 (N_3497,In_242,N_2206);
nand U3498 (N_3498,In_3390,In_3444);
or U3499 (N_3499,N_1539,In_236);
and U3500 (N_3500,N_1437,N_1210);
or U3501 (N_3501,N_2463,N_2329);
and U3502 (N_3502,N_2371,N_2223);
and U3503 (N_3503,N_2363,N_2129);
and U3504 (N_3504,N_1495,N_2921);
xor U3505 (N_3505,In_2994,N_2841);
nand U3506 (N_3506,N_2026,N_2470);
xor U3507 (N_3507,N_1643,N_2352);
nor U3508 (N_3508,In_3496,N_2205);
or U3509 (N_3509,N_2219,N_2565);
nand U3510 (N_3510,N_1727,N_2171);
xor U3511 (N_3511,N_2810,N_2063);
xnor U3512 (N_3512,N_2228,In_3544);
xnor U3513 (N_3513,N_1999,N_2234);
xnor U3514 (N_3514,N_2057,N_2679);
xnor U3515 (N_3515,N_2793,N_2931);
or U3516 (N_3516,In_3150,N_2160);
nand U3517 (N_3517,N_2163,In_4585);
nand U3518 (N_3518,N_1958,N_794);
or U3519 (N_3519,N_2777,In_4949);
and U3520 (N_3520,N_2941,In_3583);
or U3521 (N_3521,N_1395,N_2550);
or U3522 (N_3522,N_2354,N_2186);
xnor U3523 (N_3523,N_2539,N_2029);
nand U3524 (N_3524,In_3196,N_2497);
nand U3525 (N_3525,N_2987,N_1754);
or U3526 (N_3526,N_2412,N_2479);
and U3527 (N_3527,N_2713,N_2235);
or U3528 (N_3528,In_3160,N_2210);
nand U3529 (N_3529,N_2465,N_2722);
or U3530 (N_3530,N_2460,N_1128);
and U3531 (N_3531,N_2484,N_1806);
and U3532 (N_3532,N_2847,N_1506);
xnor U3533 (N_3533,N_2357,N_1165);
xnor U3534 (N_3534,In_2626,N_2914);
nand U3535 (N_3535,N_2306,N_2197);
xnor U3536 (N_3536,N_1755,N_2506);
xor U3537 (N_3537,N_2867,N_2869);
xnor U3538 (N_3538,N_2809,N_1803);
nand U3539 (N_3539,N_2718,N_1022);
and U3540 (N_3540,N_2274,N_2696);
nor U3541 (N_3541,N_2217,N_2432);
nor U3542 (N_3542,N_1810,N_1408);
and U3543 (N_3543,N_1157,N_2368);
or U3544 (N_3544,N_1696,N_2090);
xor U3545 (N_3545,N_2167,N_2103);
xnor U3546 (N_3546,N_2386,In_190);
nand U3547 (N_3547,N_2833,N_2800);
xnor U3548 (N_3548,N_702,N_1858);
and U3549 (N_3549,In_4396,N_911);
nor U3550 (N_3550,In_3711,N_1176);
nor U3551 (N_3551,N_2196,N_1183);
and U3552 (N_3552,N_1929,N_2001);
nor U3553 (N_3553,N_2518,N_1035);
nor U3554 (N_3554,N_2008,In_3152);
or U3555 (N_3555,N_33,N_2074);
and U3556 (N_3556,N_2439,In_2173);
xor U3557 (N_3557,In_3483,N_2949);
xor U3558 (N_3558,N_2597,In_612);
or U3559 (N_3559,N_1211,N_1093);
xor U3560 (N_3560,N_2403,In_1328);
or U3561 (N_3561,N_2898,N_2087);
or U3562 (N_3562,N_1486,N_2616);
or U3563 (N_3563,N_632,N_533);
and U3564 (N_3564,In_673,In_2034);
or U3565 (N_3565,N_2559,N_2742);
or U3566 (N_3566,In_985,N_2608);
or U3567 (N_3567,N_2367,N_2115);
nand U3568 (N_3568,N_2192,N_1533);
xnor U3569 (N_3569,N_2621,N_1077);
and U3570 (N_3570,In_3841,N_406);
nor U3571 (N_3571,In_224,N_2747);
nor U3572 (N_3572,N_2772,N_2135);
nand U3573 (N_3573,In_603,N_2586);
xnor U3574 (N_3574,N_1312,N_1335);
xnor U3575 (N_3575,N_2951,N_2348);
nand U3576 (N_3576,N_2838,N_948);
or U3577 (N_3577,N_2332,N_1494);
and U3578 (N_3578,N_1142,N_1994);
xor U3579 (N_3579,N_2044,In_2165);
nor U3580 (N_3580,N_2850,In_3261);
and U3581 (N_3581,N_2680,N_2536);
nand U3582 (N_3582,N_2641,N_2410);
xor U3583 (N_3583,N_2246,N_2786);
nand U3584 (N_3584,N_2582,In_364);
nand U3585 (N_3585,In_4017,In_3912);
nand U3586 (N_3586,In_1529,N_2283);
nand U3587 (N_3587,N_2288,In_1793);
or U3588 (N_3588,N_1594,N_2452);
and U3589 (N_3589,N_2140,In_4954);
nor U3590 (N_3590,N_2765,N_1245);
nor U3591 (N_3591,N_740,N_2216);
or U3592 (N_3592,N_2629,N_2844);
nand U3593 (N_3593,In_4213,N_1534);
nand U3594 (N_3594,In_896,N_2295);
nor U3595 (N_3595,N_2650,In_3705);
and U3596 (N_3596,In_911,N_1048);
or U3597 (N_3597,N_2429,N_2965);
and U3598 (N_3598,In_3262,In_4448);
xor U3599 (N_3599,N_2801,N_379);
xor U3600 (N_3600,N_1007,N_893);
nand U3601 (N_3601,N_1449,In_4097);
nand U3602 (N_3602,N_1306,In_4833);
and U3603 (N_3603,N_872,In_3310);
xnor U3604 (N_3604,N_1813,N_2421);
nor U3605 (N_3605,N_2620,N_1115);
nand U3606 (N_3606,N_2118,N_2330);
or U3607 (N_3607,In_643,In_282);
nor U3608 (N_3608,N_2198,N_547);
or U3609 (N_3609,N_2366,N_2032);
xnor U3610 (N_3610,In_294,N_1749);
nor U3611 (N_3611,N_2457,N_572);
or U3612 (N_3612,In_785,N_1403);
nor U3613 (N_3613,N_2855,N_1742);
nand U3614 (N_3614,In_4924,In_4498);
nor U3615 (N_3615,N_2207,N_2488);
nor U3616 (N_3616,In_4622,N_2495);
and U3617 (N_3617,N_2897,N_2021);
or U3618 (N_3618,N_2174,N_2031);
and U3619 (N_3619,N_2286,N_2715);
and U3620 (N_3620,N_1624,In_1895);
or U3621 (N_3621,In_3197,N_10);
nand U3622 (N_3622,In_2391,N_2293);
xor U3623 (N_3623,In_2084,In_4511);
xnor U3624 (N_3624,N_1103,N_2172);
nand U3625 (N_3625,N_2240,N_2049);
nand U3626 (N_3626,N_2611,N_1399);
nand U3627 (N_3627,N_1490,N_279);
and U3628 (N_3628,In_3629,In_880);
nand U3629 (N_3629,In_4322,In_3285);
nand U3630 (N_3630,N_2478,N_2183);
and U3631 (N_3631,N_2254,N_1940);
and U3632 (N_3632,N_2132,N_1162);
or U3633 (N_3633,N_1711,In_2601);
nor U3634 (N_3634,N_2222,N_2761);
and U3635 (N_3635,N_2225,N_2907);
or U3636 (N_3636,N_2827,N_461);
nand U3637 (N_3637,N_2237,N_2927);
nor U3638 (N_3638,N_497,N_1856);
or U3639 (N_3639,N_2926,N_2255);
nor U3640 (N_3640,In_3873,N_2994);
nand U3641 (N_3641,N_1215,N_2507);
or U3642 (N_3642,N_2253,N_2893);
xnor U3643 (N_3643,In_1770,N_2035);
nand U3644 (N_3644,N_726,N_2500);
nand U3645 (N_3645,N_2088,N_2269);
and U3646 (N_3646,N_2575,N_2454);
and U3647 (N_3647,N_1907,N_2646);
or U3648 (N_3648,N_1944,N_2091);
xnor U3649 (N_3649,N_2524,N_2913);
xnor U3650 (N_3650,N_540,N_2557);
nor U3651 (N_3651,N_2537,In_4442);
nand U3652 (N_3652,N_1072,In_2201);
nand U3653 (N_3653,N_2464,N_2343);
xnor U3654 (N_3654,N_856,In_2492);
nor U3655 (N_3655,N_1436,N_1589);
nor U3656 (N_3656,N_2625,In_2853);
nand U3657 (N_3657,N_2894,N_2239);
xor U3658 (N_3658,In_4467,N_2123);
xor U3659 (N_3659,In_4394,N_2202);
nand U3660 (N_3660,N_1707,N_2400);
and U3661 (N_3661,In_1056,In_1495);
nand U3662 (N_3662,N_2846,N_1396);
or U3663 (N_3663,N_2674,N_2788);
and U3664 (N_3664,In_3305,In_2421);
nor U3665 (N_3665,N_2609,N_2979);
and U3666 (N_3666,N_2012,In_2750);
xnor U3667 (N_3667,N_2038,N_2984);
and U3668 (N_3668,N_1333,In_3961);
nor U3669 (N_3669,In_1624,N_2005);
or U3670 (N_3670,N_2610,In_3899);
xor U3671 (N_3671,N_170,N_1573);
nand U3672 (N_3672,N_2191,N_1979);
nor U3673 (N_3673,N_2256,N_1343);
nor U3674 (N_3674,N_1801,In_937);
or U3675 (N_3675,N_2933,N_2208);
nand U3676 (N_3676,N_2751,N_618);
nor U3677 (N_3677,N_2146,N_649);
nand U3678 (N_3678,N_1599,N_1112);
and U3679 (N_3679,N_966,N_2267);
and U3680 (N_3680,In_4787,N_2700);
nor U3681 (N_3681,N_983,N_2615);
and U3682 (N_3682,N_2910,N_2436);
nand U3683 (N_3683,N_2431,N_2980);
nor U3684 (N_3684,N_2874,N_2346);
nor U3685 (N_3685,N_2428,N_2560);
or U3686 (N_3686,N_2226,N_2583);
nor U3687 (N_3687,In_351,N_2564);
and U3688 (N_3688,N_1784,N_2555);
nand U3689 (N_3689,N_2250,N_2618);
or U3690 (N_3690,In_3468,N_2041);
xnor U3691 (N_3691,In_389,In_740);
and U3692 (N_3692,N_417,In_2094);
and U3693 (N_3693,N_2056,N_2047);
or U3694 (N_3694,N_2870,In_3241);
or U3695 (N_3695,N_1511,In_3155);
nand U3696 (N_3696,N_1647,In_296);
xor U3697 (N_3697,N_2048,N_2482);
and U3698 (N_3698,In_1050,N_2376);
nand U3699 (N_3699,N_2173,N_2201);
or U3700 (N_3700,In_1776,In_4231);
nand U3701 (N_3701,N_2626,N_2738);
xor U3702 (N_3702,N_2441,N_2153);
xor U3703 (N_3703,N_2498,N_1747);
nand U3704 (N_3704,N_1593,N_873);
nand U3705 (N_3705,In_1693,In_157);
or U3706 (N_3706,N_2714,N_2107);
nor U3707 (N_3707,N_182,N_1039);
nand U3708 (N_3708,N_2691,N_2837);
and U3709 (N_3709,N_2996,N_2887);
xor U3710 (N_3710,In_507,N_2822);
nand U3711 (N_3711,N_1776,N_2543);
nor U3712 (N_3712,N_2303,N_2143);
and U3713 (N_3713,N_1445,N_2628);
xnor U3714 (N_3714,N_1608,N_2883);
xnor U3715 (N_3715,N_2561,N_2918);
xnor U3716 (N_3716,N_1377,N_2361);
or U3717 (N_3717,In_2658,N_2814);
nand U3718 (N_3718,In_3866,N_384);
and U3719 (N_3719,N_2426,N_2471);
nor U3720 (N_3720,N_1153,In_476);
or U3721 (N_3721,N_1863,N_2024);
or U3722 (N_3722,In_3441,N_2728);
nand U3723 (N_3723,N_2282,In_2465);
nand U3724 (N_3724,N_1402,In_573);
nand U3725 (N_3725,N_1346,In_2241);
and U3726 (N_3726,N_369,N_2391);
xnor U3727 (N_3727,N_2596,N_2462);
xor U3728 (N_3728,In_4226,N_2681);
nand U3729 (N_3729,In_3810,N_1341);
and U3730 (N_3730,N_126,In_4203);
or U3731 (N_3731,N_1706,N_938);
nand U3732 (N_3732,N_2554,N_950);
xor U3733 (N_3733,In_2948,N_2864);
nand U3734 (N_3734,N_1645,In_268);
and U3735 (N_3735,N_741,In_3434);
xnor U3736 (N_3736,N_2659,N_2244);
or U3737 (N_3737,N_2474,N_2296);
nor U3738 (N_3738,N_2266,N_642);
or U3739 (N_3739,N_1078,In_3655);
nand U3740 (N_3740,N_2770,N_2902);
xnor U3741 (N_3741,N_1167,N_1330);
nor U3742 (N_3742,N_2825,In_2790);
and U3743 (N_3743,N_949,N_821);
and U3744 (N_3744,N_2577,N_2571);
and U3745 (N_3745,In_4289,In_4936);
nor U3746 (N_3746,N_2151,In_2258);
xnor U3747 (N_3747,N_2311,N_2531);
and U3748 (N_3748,N_2698,N_2578);
xor U3749 (N_3749,N_1502,N_2686);
nor U3750 (N_3750,N_123,N_1816);
nor U3751 (N_3751,In_2430,N_1425);
nand U3752 (N_3752,N_2851,N_2230);
and U3753 (N_3753,N_2251,N_1021);
or U3754 (N_3754,N_2835,N_2476);
nand U3755 (N_3755,N_2297,N_2619);
nor U3756 (N_3756,N_2059,N_1375);
xor U3757 (N_3757,N_2194,N_1665);
nand U3758 (N_3758,In_2091,N_1405);
nand U3759 (N_3759,N_2662,N_2374);
or U3760 (N_3760,N_2684,N_2221);
nand U3761 (N_3761,In_3167,In_2988);
xnor U3762 (N_3762,N_2344,N_2300);
nor U3763 (N_3763,In_2377,N_1441);
or U3764 (N_3764,N_2966,N_1678);
nor U3765 (N_3765,N_443,In_1514);
xnor U3766 (N_3766,N_883,In_561);
nor U3767 (N_3767,N_1018,N_647);
nand U3768 (N_3768,In_4414,N_2880);
and U3769 (N_3769,In_383,N_2261);
nand U3770 (N_3770,N_2013,N_2290);
and U3771 (N_3771,N_2729,N_2409);
nand U3772 (N_3772,N_2080,In_115);
xor U3773 (N_3773,In_3928,N_1419);
nor U3774 (N_3774,In_4772,In_4569);
nand U3775 (N_3775,N_2362,In_4538);
nand U3776 (N_3776,In_4840,N_2656);
nor U3777 (N_3777,N_2006,N_2548);
and U3778 (N_3778,In_2316,N_2730);
nor U3779 (N_3779,N_2390,N_1898);
nand U3780 (N_3780,In_1635,N_2345);
xnor U3781 (N_3781,N_1899,N_2360);
and U3782 (N_3782,N_2530,N_2824);
or U3783 (N_3783,In_1900,N_2164);
xor U3784 (N_3784,N_1996,In_663);
or U3785 (N_3785,In_1570,N_364);
nand U3786 (N_3786,N_2909,N_2858);
and U3787 (N_3787,In_1032,N_164);
and U3788 (N_3788,N_566,In_2092);
and U3789 (N_3789,In_2296,N_2922);
nand U3790 (N_3790,In_562,N_2977);
nand U3791 (N_3791,In_1817,N_2165);
nand U3792 (N_3792,N_1877,N_2099);
nand U3793 (N_3793,N_1389,N_2859);
or U3794 (N_3794,N_2813,In_4083);
or U3795 (N_3795,N_322,N_2122);
xor U3796 (N_3796,In_4479,N_1909);
nor U3797 (N_3797,N_300,N_2231);
or U3798 (N_3798,N_2740,N_2301);
or U3799 (N_3799,N_2305,N_2037);
nand U3800 (N_3800,N_2370,In_2269);
or U3801 (N_3801,N_1264,N_2781);
nor U3802 (N_3802,N_2848,N_491);
nor U3803 (N_3803,N_1019,N_2533);
or U3804 (N_3804,N_2794,N_2324);
xnor U3805 (N_3805,In_3986,In_2915);
nand U3806 (N_3806,N_2613,N_2184);
xor U3807 (N_3807,In_1202,N_2811);
or U3808 (N_3808,N_558,N_2892);
nand U3809 (N_3809,N_1184,N_2383);
nor U3810 (N_3810,N_2480,In_1141);
or U3811 (N_3811,N_2203,In_2884);
and U3812 (N_3812,In_4129,N_561);
nand U3813 (N_3813,In_3878,In_4292);
and U3814 (N_3814,N_2055,N_2798);
or U3815 (N_3815,In_514,N_1569);
and U3816 (N_3816,In_2021,In_759);
nand U3817 (N_3817,In_1106,N_2189);
nand U3818 (N_3818,N_2200,N_2302);
and U3819 (N_3819,N_2473,N_2541);
or U3820 (N_3820,N_2444,In_1310);
or U3821 (N_3821,N_1578,In_1206);
nor U3822 (N_3822,N_2711,In_4360);
and U3823 (N_3823,N_2492,N_2213);
nand U3824 (N_3824,N_2992,In_1758);
xnor U3825 (N_3825,N_2699,In_3308);
xnor U3826 (N_3826,N_2702,N_2955);
xor U3827 (N_3827,N_2687,N_139);
or U3828 (N_3828,N_2804,N_2493);
and U3829 (N_3829,In_652,N_2587);
and U3830 (N_3830,In_795,N_2920);
nand U3831 (N_3831,N_2078,In_2606);
or U3832 (N_3832,N_2483,In_1819);
or U3833 (N_3833,In_4629,N_2418);
and U3834 (N_3834,N_2764,N_2832);
xnor U3835 (N_3835,N_2461,In_710);
or U3836 (N_3836,N_1628,N_2598);
nand U3837 (N_3837,N_2667,N_1347);
nor U3838 (N_3838,N_2416,N_1427);
nor U3839 (N_3839,N_1320,In_2807);
xor U3840 (N_3840,N_2633,N_1061);
or U3841 (N_3841,In_2242,In_2002);
and U3842 (N_3842,In_1703,In_3265);
or U3843 (N_3843,N_1040,In_670);
nand U3844 (N_3844,N_1125,N_2912);
nand U3845 (N_3845,N_2644,N_2852);
nor U3846 (N_3846,In_1,In_2419);
nor U3847 (N_3847,N_2128,N_2050);
and U3848 (N_3848,N_2475,N_1133);
nand U3849 (N_3849,N_1848,In_2025);
and U3850 (N_3850,N_2888,N_2988);
or U3851 (N_3851,In_1478,In_1461);
nor U3852 (N_3852,N_2285,N_2312);
xor U3853 (N_3853,N_2725,N_2380);
nand U3854 (N_3854,N_2327,N_2125);
xor U3855 (N_3855,In_2010,N_1189);
or U3856 (N_3856,N_2082,In_1552);
nand U3857 (N_3857,In_2125,N_2214);
nand U3858 (N_3858,N_2382,N_2514);
or U3859 (N_3859,N_2763,In_323);
nand U3860 (N_3860,N_2481,In_2952);
xor U3861 (N_3861,N_2900,N_2232);
or U3862 (N_3862,N_2673,N_2961);
nor U3863 (N_3863,N_2169,N_2717);
nor U3864 (N_3864,In_3168,In_1904);
or U3865 (N_3865,N_2778,N_756);
xnor U3866 (N_3866,N_623,N_2273);
or U3867 (N_3867,N_1649,N_2759);
or U3868 (N_3868,N_134,N_2355);
xnor U3869 (N_3869,N_828,N_1651);
or U3870 (N_3870,In_4212,N_329);
and U3871 (N_3871,N_933,N_2935);
xnor U3872 (N_3872,N_2003,In_783);
nor U3873 (N_3873,In_3343,N_1736);
and U3874 (N_3874,In_29,In_1953);
or U3875 (N_3875,N_2472,N_2522);
xnor U3876 (N_3876,N_1161,N_2106);
nand U3877 (N_3877,N_1108,N_1415);
or U3878 (N_3878,N_2946,In_4779);
and U3879 (N_3879,In_1969,N_2806);
nor U3880 (N_3880,N_2384,In_3611);
nor U3881 (N_3881,In_2114,N_2649);
nor U3882 (N_3882,N_1057,N_2154);
and U3883 (N_3883,In_2400,In_1187);
xnor U3884 (N_3884,N_2668,In_846);
or U3885 (N_3885,N_2378,N_1690);
nand U3886 (N_3886,N_2127,N_1300);
xnor U3887 (N_3887,N_847,N_408);
xor U3888 (N_3888,N_2676,N_2638);
and U3889 (N_3889,N_1590,N_1911);
nor U3890 (N_3890,N_448,N_1982);
nand U3891 (N_3891,N_2990,N_2773);
xnor U3892 (N_3892,N_2249,N_2944);
nor U3893 (N_3893,N_1558,N_1043);
xnor U3894 (N_3894,N_1715,N_2934);
and U3895 (N_3895,N_2501,N_1388);
xnor U3896 (N_3896,N_2052,In_1501);
nand U3897 (N_3897,N_2489,In_3437);
xnor U3898 (N_3898,N_2640,N_187);
xor U3899 (N_3899,N_2350,N_2563);
xnor U3900 (N_3900,In_2515,In_2664);
xnor U3901 (N_3901,In_1130,N_2820);
xor U3902 (N_3902,In_1783,N_2663);
and U3903 (N_3903,N_2124,N_2602);
nand U3904 (N_3904,N_1083,N_2248);
or U3905 (N_3905,N_1352,In_4483);
nand U3906 (N_3906,In_2542,N_2799);
nor U3907 (N_3907,N_1753,N_327);
nor U3908 (N_3908,N_1472,N_2712);
xor U3909 (N_3909,In_166,N_2070);
and U3910 (N_3910,N_2562,N_2614);
nand U3911 (N_3911,N_2693,N_1398);
or U3912 (N_3912,N_2304,N_2617);
nand U3913 (N_3913,N_2069,N_2397);
nand U3914 (N_3914,N_2642,N_2830);
or U3915 (N_3915,N_1763,N_2102);
nor U3916 (N_3916,N_2795,N_1302);
xor U3917 (N_3917,N_2215,N_2150);
or U3918 (N_3918,In_4789,N_2053);
nor U3919 (N_3919,N_1467,N_1787);
or U3920 (N_3920,N_105,In_997);
nor U3921 (N_3921,In_3138,In_2047);
xor U3922 (N_3922,N_8,N_2754);
nor U3923 (N_3923,In_1471,In_1754);
and U3924 (N_3924,In_3798,In_1715);
nand U3925 (N_3925,N_511,N_2097);
nor U3926 (N_3926,N_1064,In_2625);
nand U3927 (N_3927,In_1127,In_2442);
xnor U3928 (N_3928,N_2259,N_1872);
nor U3929 (N_3929,In_2603,N_2373);
xor U3930 (N_3930,N_2937,N_2529);
or U3931 (N_3931,N_1190,N_1557);
xor U3932 (N_3932,N_2477,N_2094);
nor U3933 (N_3933,N_2637,N_2972);
xnor U3934 (N_3934,In_2279,N_2466);
and U3935 (N_3935,N_2045,In_1956);
and U3936 (N_3936,N_2704,N_2022);
nor U3937 (N_3937,N_240,N_2589);
nor U3938 (N_3938,N_1953,N_2317);
nand U3939 (N_3939,N_2110,N_2523);
nor U3940 (N_3940,N_2607,N_2655);
and U3941 (N_3941,N_1894,N_2424);
nor U3942 (N_3942,N_1177,N_2923);
and U3943 (N_3943,N_2895,In_2976);
and U3944 (N_3944,N_753,In_3813);
nand U3945 (N_3945,N_2797,In_3042);
xnor U3946 (N_3946,N_290,N_2369);
nor U3947 (N_3947,In_4244,N_1409);
xor U3948 (N_3948,N_2672,N_262);
xor U3949 (N_3949,N_2622,N_1610);
nand U3950 (N_3950,N_2084,N_2703);
nor U3951 (N_3951,N_2133,N_2157);
nor U3952 (N_3952,N_2020,N_1614);
nand U3953 (N_3953,N_2854,N_2280);
or U3954 (N_3954,In_293,In_2941);
or U3955 (N_3955,N_923,N_2181);
nor U3956 (N_3956,N_2861,In_3578);
nor U3957 (N_3957,N_2682,N_2653);
and U3958 (N_3958,N_2652,In_4932);
or U3959 (N_3959,N_2553,N_1266);
or U3960 (N_3960,N_2062,In_1048);
nor U3961 (N_3961,N_2938,N_2985);
and U3962 (N_3962,N_579,N_2275);
nand U3963 (N_3963,In_633,In_4470);
nor U3964 (N_3964,In_709,N_2974);
or U3965 (N_3965,N_1543,N_2896);
or U3966 (N_3966,In_3249,In_4879);
and U3967 (N_3967,N_2113,N_931);
or U3968 (N_3968,In_1631,N_2574);
nand U3969 (N_3969,N_2281,N_2046);
or U3970 (N_3970,N_2294,N_2508);
and U3971 (N_3971,In_80,N_2277);
nand U3972 (N_3972,N_2753,N_1745);
nand U3973 (N_3973,N_1042,N_2262);
or U3974 (N_3974,N_2015,In_2327);
xnor U3975 (N_3975,N_661,N_2521);
nand U3976 (N_3976,In_4589,N_2552);
nand U3977 (N_3977,N_2156,In_4485);
nor U3978 (N_3978,N_2569,N_296);
nand U3979 (N_3979,In_160,N_41);
nor U3980 (N_3980,N_2025,N_2816);
nor U3981 (N_3981,In_226,In_4497);
nand U3982 (N_3982,In_3169,N_2527);
or U3983 (N_3983,N_2415,N_2651);
nor U3984 (N_3984,N_488,In_504);
nor U3985 (N_3985,N_2155,N_2881);
nand U3986 (N_3986,N_1924,N_2220);
nor U3987 (N_3987,N_1702,In_2389);
xnor U3988 (N_3988,In_366,In_3562);
and U3989 (N_3989,N_2976,N_2875);
nand U3990 (N_3990,N_2915,N_2486);
and U3991 (N_3991,N_2971,N_1327);
nor U3992 (N_3992,N_2218,N_150);
or U3993 (N_3993,In_3154,N_2209);
nor U3994 (N_3994,N_2034,N_556);
nor U3995 (N_3995,N_2494,N_2748);
and U3996 (N_3996,N_1802,In_1115);
xor U3997 (N_3997,In_3220,N_2190);
nand U3998 (N_3998,N_1137,N_2512);
and U3999 (N_3999,N_2719,N_1365);
nand U4000 (N_4000,N_3019,N_3933);
nand U4001 (N_4001,N_3832,N_3394);
nor U4002 (N_4002,N_3289,N_3906);
nand U4003 (N_4003,N_3664,N_3058);
and U4004 (N_4004,N_3255,N_3232);
and U4005 (N_4005,N_3699,N_3169);
and U4006 (N_4006,N_3754,N_3195);
nor U4007 (N_4007,N_3367,N_3780);
nor U4008 (N_4008,N_3273,N_3385);
nor U4009 (N_4009,N_3923,N_3763);
or U4010 (N_4010,N_3547,N_3485);
nand U4011 (N_4011,N_3454,N_3929);
and U4012 (N_4012,N_3839,N_3218);
and U4013 (N_4013,N_3194,N_3675);
xor U4014 (N_4014,N_3617,N_3348);
or U4015 (N_4015,N_3107,N_3503);
xor U4016 (N_4016,N_3198,N_3900);
nor U4017 (N_4017,N_3023,N_3850);
xor U4018 (N_4018,N_3057,N_3338);
nor U4019 (N_4019,N_3138,N_3036);
and U4020 (N_4020,N_3114,N_3949);
xnor U4021 (N_4021,N_3247,N_3251);
and U4022 (N_4022,N_3185,N_3126);
nor U4023 (N_4023,N_3256,N_3545);
nand U4024 (N_4024,N_3483,N_3531);
and U4025 (N_4025,N_3182,N_3868);
nor U4026 (N_4026,N_3679,N_3476);
and U4027 (N_4027,N_3712,N_3504);
and U4028 (N_4028,N_3027,N_3093);
or U4029 (N_4029,N_3134,N_3139);
nand U4030 (N_4030,N_3796,N_3276);
nor U4031 (N_4031,N_3004,N_3804);
nand U4032 (N_4032,N_3015,N_3172);
nand U4033 (N_4033,N_3197,N_3686);
or U4034 (N_4034,N_3970,N_3691);
nor U4035 (N_4035,N_3601,N_3698);
nand U4036 (N_4036,N_3452,N_3254);
and U4037 (N_4037,N_3755,N_3744);
nand U4038 (N_4038,N_3627,N_3075);
xor U4039 (N_4039,N_3189,N_3781);
and U4040 (N_4040,N_3302,N_3604);
nand U4041 (N_4041,N_3669,N_3438);
and U4042 (N_4042,N_3654,N_3646);
nor U4043 (N_4043,N_3620,N_3346);
nor U4044 (N_4044,N_3487,N_3040);
or U4045 (N_4045,N_3821,N_3161);
xor U4046 (N_4046,N_3061,N_3073);
or U4047 (N_4047,N_3739,N_3857);
or U4048 (N_4048,N_3365,N_3270);
and U4049 (N_4049,N_3773,N_3099);
nand U4050 (N_4050,N_3786,N_3459);
nor U4051 (N_4051,N_3767,N_3208);
and U4052 (N_4052,N_3676,N_3275);
nor U4053 (N_4053,N_3100,N_3074);
nor U4054 (N_4054,N_3635,N_3887);
and U4055 (N_4055,N_3037,N_3978);
and U4056 (N_4056,N_3340,N_3916);
xnor U4057 (N_4057,N_3315,N_3854);
or U4058 (N_4058,N_3445,N_3965);
or U4059 (N_4059,N_3966,N_3924);
and U4060 (N_4060,N_3648,N_3245);
nor U4061 (N_4061,N_3801,N_3407);
nor U4062 (N_4062,N_3615,N_3886);
nor U4063 (N_4063,N_3529,N_3294);
or U4064 (N_4064,N_3290,N_3008);
or U4065 (N_4065,N_3031,N_3539);
and U4066 (N_4066,N_3291,N_3947);
and U4067 (N_4067,N_3707,N_3910);
and U4068 (N_4068,N_3629,N_3964);
or U4069 (N_4069,N_3234,N_3889);
nor U4070 (N_4070,N_3769,N_3544);
or U4071 (N_4071,N_3848,N_3072);
or U4072 (N_4072,N_3077,N_3742);
nand U4073 (N_4073,N_3113,N_3395);
nand U4074 (N_4074,N_3064,N_3852);
and U4075 (N_4075,N_3472,N_3694);
or U4076 (N_4076,N_3990,N_3610);
xnor U4077 (N_4077,N_3591,N_3626);
and U4078 (N_4078,N_3761,N_3462);
xor U4079 (N_4079,N_3871,N_3378);
and U4080 (N_4080,N_3520,N_3860);
or U4081 (N_4081,N_3828,N_3749);
or U4082 (N_4082,N_3216,N_3103);
and U4083 (N_4083,N_3432,N_3693);
and U4084 (N_4084,N_3685,N_3044);
xnor U4085 (N_4085,N_3339,N_3342);
or U4086 (N_4086,N_3173,N_3587);
nor U4087 (N_4087,N_3643,N_3238);
nand U4088 (N_4088,N_3128,N_3489);
nand U4089 (N_4089,N_3830,N_3552);
or U4090 (N_4090,N_3250,N_3402);
or U4091 (N_4091,N_3533,N_3775);
nand U4092 (N_4092,N_3571,N_3778);
and U4093 (N_4093,N_3651,N_3311);
nor U4094 (N_4094,N_3437,N_3010);
and U4095 (N_4095,N_3084,N_3936);
or U4096 (N_4096,N_3033,N_3435);
or U4097 (N_4097,N_3145,N_3540);
nor U4098 (N_4098,N_3522,N_3988);
xnor U4099 (N_4099,N_3764,N_3463);
and U4100 (N_4100,N_3067,N_3710);
xnor U4101 (N_4101,N_3457,N_3969);
nor U4102 (N_4102,N_3049,N_3656);
nand U4103 (N_4103,N_3175,N_3295);
nand U4104 (N_4104,N_3841,N_3362);
and U4105 (N_4105,N_3876,N_3785);
xor U4106 (N_4106,N_3560,N_3500);
nand U4107 (N_4107,N_3371,N_3716);
or U4108 (N_4108,N_3375,N_3078);
or U4109 (N_4109,N_3230,N_3240);
xor U4110 (N_4110,N_3193,N_3129);
nor U4111 (N_4111,N_3757,N_3233);
or U4112 (N_4112,N_3538,N_3244);
nor U4113 (N_4113,N_3598,N_3762);
and U4114 (N_4114,N_3902,N_3605);
and U4115 (N_4115,N_3870,N_3895);
nand U4116 (N_4116,N_3260,N_3589);
xor U4117 (N_4117,N_3097,N_3680);
xnor U4118 (N_4118,N_3042,N_3011);
xor U4119 (N_4119,N_3105,N_3259);
nor U4120 (N_4120,N_3199,N_3810);
nor U4121 (N_4121,N_3746,N_3431);
xnor U4122 (N_4122,N_3364,N_3214);
xor U4123 (N_4123,N_3024,N_3131);
nand U4124 (N_4124,N_3579,N_3224);
nand U4125 (N_4125,N_3386,N_3471);
nand U4126 (N_4126,N_3133,N_3674);
and U4127 (N_4127,N_3312,N_3722);
or U4128 (N_4128,N_3771,N_3306);
xor U4129 (N_4129,N_3050,N_3249);
xnor U4130 (N_4130,N_3055,N_3650);
nor U4131 (N_4131,N_3086,N_3901);
xor U4132 (N_4132,N_3726,N_3162);
or U4133 (N_4133,N_3020,N_3115);
nor U4134 (N_4134,N_3409,N_3183);
xnor U4135 (N_4135,N_3192,N_3750);
nor U4136 (N_4136,N_3774,N_3649);
or U4137 (N_4137,N_3867,N_3071);
xor U4138 (N_4138,N_3989,N_3493);
and U4139 (N_4139,N_3140,N_3657);
nand U4140 (N_4140,N_3089,N_3516);
nand U4141 (N_4141,N_3932,N_3595);
or U4142 (N_4142,N_3800,N_3323);
nor U4143 (N_4143,N_3765,N_3748);
xor U4144 (N_4144,N_3287,N_3628);
nand U4145 (N_4145,N_3687,N_3013);
or U4146 (N_4146,N_3137,N_3150);
nand U4147 (N_4147,N_3802,N_3546);
nand U4148 (N_4148,N_3112,N_3207);
nor U4149 (N_4149,N_3388,N_3513);
nand U4150 (N_4150,N_3502,N_3599);
or U4151 (N_4151,N_3661,N_3678);
nor U4152 (N_4152,N_3704,N_3813);
xnor U4153 (N_4153,N_3844,N_3905);
xor U4154 (N_4154,N_3636,N_3743);
nor U4155 (N_4155,N_3341,N_3968);
xor U4156 (N_4156,N_3092,N_3630);
nand U4157 (N_4157,N_3701,N_3456);
and U4158 (N_4158,N_3724,N_3593);
and U4159 (N_4159,N_3066,N_3142);
or U4160 (N_4160,N_3110,N_3326);
or U4161 (N_4161,N_3580,N_3223);
or U4162 (N_4162,N_3586,N_3335);
xor U4163 (N_4163,N_3083,N_3009);
and U4164 (N_4164,N_3090,N_3959);
nor U4165 (N_4165,N_3891,N_3351);
and U4166 (N_4166,N_3337,N_3170);
xnor U4167 (N_4167,N_3148,N_3399);
nor U4168 (N_4168,N_3653,N_3448);
or U4169 (N_4169,N_3585,N_3235);
xnor U4170 (N_4170,N_3555,N_3515);
and U4171 (N_4171,N_3715,N_3242);
and U4172 (N_4172,N_3381,N_3479);
nand U4173 (N_4173,N_3795,N_3171);
or U4174 (N_4174,N_3683,N_3618);
nand U4175 (N_4175,N_3842,N_3915);
and U4176 (N_4176,N_3792,N_3590);
or U4177 (N_4177,N_3632,N_3144);
nand U4178 (N_4178,N_3440,N_3992);
xor U4179 (N_4179,N_3350,N_3288);
nor U4180 (N_4180,N_3467,N_3713);
nand U4181 (N_4181,N_3904,N_3612);
nand U4182 (N_4182,N_3411,N_3971);
or U4183 (N_4183,N_3534,N_3246);
nor U4184 (N_4184,N_3060,N_3510);
nand U4185 (N_4185,N_3805,N_3881);
and U4186 (N_4186,N_3327,N_3422);
nor U4187 (N_4187,N_3740,N_3400);
nand U4188 (N_4188,N_3280,N_3028);
and U4189 (N_4189,N_3321,N_3903);
nor U4190 (N_4190,N_3823,N_3644);
or U4191 (N_4191,N_3098,N_3731);
nor U4192 (N_4192,N_3186,N_3582);
or U4193 (N_4193,N_3486,N_3509);
nor U4194 (N_4194,N_3029,N_3007);
or U4195 (N_4195,N_3884,N_3997);
xnor U4196 (N_4196,N_3703,N_3942);
xnor U4197 (N_4197,N_3866,N_3861);
nand U4198 (N_4198,N_3859,N_3069);
nand U4199 (N_4199,N_3355,N_3553);
nand U4200 (N_4200,N_3568,N_3353);
nor U4201 (N_4201,N_3508,N_3753);
nand U4202 (N_4202,N_3621,N_3638);
or U4203 (N_4203,N_3718,N_3896);
nor U4204 (N_4204,N_3358,N_3951);
or U4205 (N_4205,N_3523,N_3322);
nor U4206 (N_4206,N_3705,N_3420);
nor U4207 (N_4207,N_3180,N_3833);
nand U4208 (N_4208,N_3414,N_3981);
xnor U4209 (N_4209,N_3877,N_3018);
and U4210 (N_4210,N_3885,N_3940);
nand U4211 (N_4211,N_3985,N_3106);
nor U4212 (N_4212,N_3541,N_3366);
xnor U4213 (N_4213,N_3984,N_3723);
nor U4214 (N_4214,N_3307,N_3392);
xnor U4215 (N_4215,N_3174,N_3677);
and U4216 (N_4216,N_3667,N_3583);
or U4217 (N_4217,N_3269,N_3888);
nor U4218 (N_4218,N_3943,N_3788);
and U4219 (N_4219,N_3334,N_3551);
and U4220 (N_4220,N_3633,N_3655);
nor U4221 (N_4221,N_3212,N_3542);
or U4222 (N_4222,N_3918,N_3954);
or U4223 (N_4223,N_3318,N_3853);
xor U4224 (N_4224,N_3770,N_3980);
nand U4225 (N_4225,N_3263,N_3660);
xnor U4226 (N_4226,N_3730,N_3054);
and U4227 (N_4227,N_3863,N_3458);
or U4228 (N_4228,N_3914,N_3447);
and U4229 (N_4229,N_3506,N_3473);
or U4230 (N_4230,N_3264,N_3639);
nand U4231 (N_4231,N_3324,N_3975);
nor U4232 (N_4232,N_3398,N_3917);
or U4233 (N_4233,N_3817,N_3536);
xor U4234 (N_4234,N_3257,N_3945);
xor U4235 (N_4235,N_3258,N_3221);
nor U4236 (N_4236,N_3228,N_3622);
xnor U4237 (N_4237,N_3397,N_3032);
or U4238 (N_4238,N_3899,N_3814);
and U4239 (N_4239,N_3229,N_3799);
or U4240 (N_4240,N_3897,N_3380);
and U4241 (N_4241,N_3436,N_3314);
nor U4242 (N_4242,N_3711,N_3825);
and U4243 (N_4243,N_3519,N_3594);
or U4244 (N_4244,N_3824,N_3014);
nor U4245 (N_4245,N_3478,N_3125);
or U4246 (N_4246,N_3776,N_3835);
xnor U4247 (N_4247,N_3132,N_3999);
xnor U4248 (N_4248,N_3892,N_3957);
xor U4249 (N_4249,N_3379,N_3157);
nor U4250 (N_4250,N_3231,N_3423);
or U4251 (N_4251,N_3127,N_3469);
or U4252 (N_4252,N_3045,N_3413);
nand U4253 (N_4253,N_3418,N_3446);
xor U4254 (N_4254,N_3526,N_3320);
nor U4255 (N_4255,N_3434,N_3453);
nand U4256 (N_4256,N_3282,N_3159);
and U4257 (N_4257,N_3424,N_3783);
and U4258 (N_4258,N_3682,N_3738);
nor U4259 (N_4259,N_3153,N_3393);
xnor U4260 (N_4260,N_3935,N_3672);
nor U4261 (N_4261,N_3470,N_3352);
and U4262 (N_4262,N_3872,N_3840);
xnor U4263 (N_4263,N_3564,N_3882);
nor U4264 (N_4264,N_3405,N_3236);
nand U4265 (N_4265,N_3963,N_3376);
or U4266 (N_4266,N_3268,N_3046);
nand U4267 (N_4267,N_3059,N_3165);
and U4268 (N_4268,N_3425,N_3645);
nor U4269 (N_4269,N_3220,N_3490);
or U4270 (N_4270,N_3298,N_3336);
or U4271 (N_4271,N_3475,N_3946);
and U4272 (N_4272,N_3427,N_3070);
xnor U4273 (N_4273,N_3634,N_3408);
nor U4274 (N_4274,N_3695,N_3973);
nor U4275 (N_4275,N_3363,N_3956);
nand U4276 (N_4276,N_3822,N_3444);
and U4277 (N_4277,N_3584,N_3967);
or U4278 (N_4278,N_3119,N_3313);
nand U4279 (N_4279,N_3869,N_3117);
nor U4280 (N_4280,N_3167,N_3567);
xor U4281 (N_4281,N_3569,N_3325);
xnor U4282 (N_4282,N_3816,N_3953);
nand U4283 (N_4283,N_3717,N_3625);
xnor U4284 (N_4284,N_3360,N_3330);
nand U4285 (N_4285,N_3297,N_3261);
and U4286 (N_4286,N_3152,N_3442);
and U4287 (N_4287,N_3637,N_3611);
nand U4288 (N_4288,N_3919,N_3370);
nand U4289 (N_4289,N_3986,N_3735);
and U4290 (N_4290,N_3300,N_3692);
xnor U4291 (N_4291,N_3184,N_3747);
nand U4292 (N_4292,N_3177,N_3797);
or U4293 (N_4293,N_3960,N_3433);
or U4294 (N_4294,N_3875,N_3017);
xor U4295 (N_4295,N_3168,N_3684);
xor U4296 (N_4296,N_3477,N_3554);
xnor U4297 (N_4297,N_3091,N_3349);
nand U4298 (N_4298,N_3791,N_3333);
nand U4299 (N_4299,N_3108,N_3053);
and U4300 (N_4300,N_3154,N_3271);
nand U4301 (N_4301,N_3211,N_3874);
nand U4302 (N_4302,N_3690,N_3124);
and U4303 (N_4303,N_3179,N_3237);
or U4304 (N_4304,N_3387,N_3521);
xnor U4305 (N_4305,N_3277,N_3826);
or U4306 (N_4306,N_3815,N_3272);
nor U4307 (N_4307,N_3441,N_3732);
nand U4308 (N_4308,N_3873,N_3666);
xnor U4309 (N_4309,N_3449,N_3697);
nand U4310 (N_4310,N_3266,N_3455);
nor U4311 (N_4311,N_3576,N_3203);
nor U4312 (N_4312,N_3081,N_3616);
xnor U4313 (N_4313,N_3623,N_3079);
and U4314 (N_4314,N_3354,N_3118);
or U4315 (N_4315,N_3931,N_3751);
and U4316 (N_4316,N_3494,N_3497);
or U4317 (N_4317,N_3429,N_3756);
nor U4318 (N_4318,N_3708,N_3213);
or U4319 (N_4319,N_3856,N_3619);
nand U4320 (N_4320,N_3880,N_3121);
xnor U4321 (N_4321,N_3451,N_3913);
or U4322 (N_4322,N_3831,N_3570);
and U4323 (N_4323,N_3518,N_3205);
nand U4324 (N_4324,N_3085,N_3329);
and U4325 (N_4325,N_3226,N_3227);
nand U4326 (N_4326,N_3845,N_3219);
and U4327 (N_4327,N_3721,N_3528);
nand U4328 (N_4328,N_3663,N_3111);
xor U4329 (N_4329,N_3846,N_3122);
xnor U4330 (N_4330,N_3994,N_3535);
or U4331 (N_4331,N_3331,N_3461);
or U4332 (N_4332,N_3838,N_3878);
xor U4333 (N_4333,N_3575,N_3995);
nor U4334 (N_4334,N_3790,N_3317);
or U4335 (N_4335,N_3720,N_3631);
and U4336 (N_4336,N_3415,N_3974);
nand U4337 (N_4337,N_3202,N_3286);
nor U4338 (N_4338,N_3927,N_3095);
nand U4339 (N_4339,N_3793,N_3076);
or U4340 (N_4340,N_3305,N_3345);
xor U4341 (N_4341,N_3204,N_3642);
or U4342 (N_4342,N_3566,N_3559);
xor U4343 (N_4343,N_3039,N_3498);
xor U4344 (N_4344,N_3301,N_3293);
nand U4345 (N_4345,N_3188,N_3096);
nand U4346 (N_4346,N_3777,N_3779);
nor U4347 (N_4347,N_3158,N_3401);
xnor U4348 (N_4348,N_3996,N_3026);
xor U4349 (N_4349,N_3241,N_3920);
xor U4350 (N_4350,N_3734,N_3789);
nor U4351 (N_4351,N_3668,N_3000);
or U4352 (N_4352,N_3784,N_3652);
or U4353 (N_4353,N_3592,N_3196);
xnor U4354 (N_4354,N_3279,N_3829);
or U4355 (N_4355,N_3016,N_3267);
or U4356 (N_4356,N_3404,N_3752);
or U4357 (N_4357,N_3819,N_3794);
nor U4358 (N_4358,N_3443,N_3530);
nor U4359 (N_4359,N_3962,N_3662);
nand U4360 (N_4360,N_3758,N_3480);
xnor U4361 (N_4361,N_3006,N_3416);
nor U4362 (N_4362,N_3149,N_3102);
nor U4363 (N_4363,N_3733,N_3807);
xor U4364 (N_4364,N_3038,N_3725);
and U4365 (N_4365,N_3041,N_3907);
nand U4366 (N_4366,N_3820,N_3958);
nand U4367 (N_4367,N_3412,N_3787);
nand U4368 (N_4368,N_3252,N_3310);
and U4369 (N_4369,N_3278,N_3556);
xnor U4370 (N_4370,N_3190,N_3603);
and U4371 (N_4371,N_3308,N_3572);
nor U4372 (N_4372,N_3088,N_3714);
and U4373 (N_4373,N_3265,N_3681);
xnor U4374 (N_4374,N_3135,N_3818);
nor U4375 (N_4375,N_3357,N_3396);
xor U4376 (N_4376,N_3658,N_3768);
nand U4377 (N_4377,N_3285,N_3602);
and U4378 (N_4378,N_3116,N_3562);
or U4379 (N_4379,N_3524,N_3403);
xnor U4380 (N_4380,N_3217,N_3166);
nand U4381 (N_4381,N_3670,N_3001);
nor U4382 (N_4382,N_3421,N_3883);
or U4383 (N_4383,N_3303,N_3745);
nor U4384 (N_4384,N_3406,N_3574);
and U4385 (N_4385,N_3858,N_3465);
or U4386 (N_4386,N_3491,N_3766);
nor U4387 (N_4387,N_3812,N_3222);
and U4388 (N_4388,N_3525,N_3501);
xnor U4389 (N_4389,N_3419,N_3048);
and U4390 (N_4390,N_3499,N_3191);
nor U4391 (N_4391,N_3944,N_3836);
and U4392 (N_4392,N_3296,N_3982);
nand U4393 (N_4393,N_3709,N_3543);
and U4394 (N_4394,N_3549,N_3082);
xnor U4395 (N_4395,N_3120,N_3359);
nor U4396 (N_4396,N_3532,N_3248);
xnor U4397 (N_4397,N_3736,N_3921);
nand U4398 (N_4398,N_3063,N_3760);
or U4399 (N_4399,N_3505,N_3808);
and U4400 (N_4400,N_3209,N_3909);
and U4401 (N_4401,N_3665,N_3737);
xnor U4402 (N_4402,N_3952,N_3147);
nor U4403 (N_4403,N_3484,N_3696);
and U4404 (N_4404,N_3806,N_3052);
and U4405 (N_4405,N_3151,N_3274);
nand U4406 (N_4406,N_3926,N_3130);
and U4407 (N_4407,N_3156,N_3062);
xnor U4408 (N_4408,N_3035,N_3215);
nor U4409 (N_4409,N_3851,N_3673);
or U4410 (N_4410,N_3080,N_3928);
nand U4411 (N_4411,N_3809,N_3608);
or U4412 (N_4412,N_3382,N_3343);
xnor U4413 (N_4413,N_3163,N_3056);
or U4414 (N_4414,N_3160,N_3460);
or U4415 (N_4415,N_3511,N_3281);
xnor U4416 (N_4416,N_3659,N_3597);
nor U4417 (N_4417,N_3136,N_3614);
nor U4418 (N_4418,N_3390,N_3930);
or U4419 (N_4419,N_3369,N_3759);
xnor U4420 (N_4420,N_3558,N_3284);
and U4421 (N_4421,N_3991,N_3563);
nand U4422 (N_4422,N_3328,N_3827);
xnor U4423 (N_4423,N_3176,N_3573);
and U4424 (N_4424,N_3640,N_3950);
or U4425 (N_4425,N_3937,N_3728);
nand U4426 (N_4426,N_3178,N_3292);
nor U4427 (N_4427,N_3210,N_3512);
or U4428 (N_4428,N_3243,N_3391);
xnor U4429 (N_4429,N_3578,N_3187);
xor U4430 (N_4430,N_3624,N_3022);
nor U4431 (N_4431,N_3374,N_3450);
xor U4432 (N_4432,N_3002,N_3347);
nor U4433 (N_4433,N_3565,N_3003);
nand U4434 (N_4434,N_3005,N_3934);
nor U4435 (N_4435,N_3025,N_3700);
nor U4436 (N_4436,N_3993,N_3983);
or U4437 (N_4437,N_3925,N_3051);
xor U4438 (N_4438,N_3976,N_3847);
and U4439 (N_4439,N_3972,N_3299);
and U4440 (N_4440,N_3862,N_3474);
and U4441 (N_4441,N_3922,N_3977);
nor U4442 (N_4442,N_3225,N_3109);
nor U4443 (N_4443,N_3262,N_3948);
nor U4444 (N_4444,N_3495,N_3332);
and U4445 (N_4445,N_3417,N_3941);
and U4446 (N_4446,N_3201,N_3987);
nand U4447 (N_4447,N_3426,N_3998);
nand U4448 (N_4448,N_3527,N_3143);
and U4449 (N_4449,N_3606,N_3898);
xor U4450 (N_4450,N_3043,N_3893);
nand U4451 (N_4451,N_3239,N_3389);
and U4452 (N_4452,N_3428,N_3410);
xor U4453 (N_4453,N_3068,N_3430);
nor U4454 (N_4454,N_3607,N_3496);
nor U4455 (N_4455,N_3319,N_3890);
and U4456 (N_4456,N_3641,N_3034);
xor U4457 (N_4457,N_3613,N_3101);
or U4458 (N_4458,N_3464,N_3577);
or U4459 (N_4459,N_3253,N_3912);
nor U4460 (N_4460,N_3384,N_3094);
xor U4461 (N_4461,N_3719,N_3849);
xnor U4462 (N_4462,N_3283,N_3837);
nand U4463 (N_4463,N_3200,N_3702);
xor U4464 (N_4464,N_3065,N_3309);
nand U4465 (N_4465,N_3537,N_3955);
or U4466 (N_4466,N_3843,N_3372);
and U4467 (N_4467,N_3141,N_3164);
and U4468 (N_4468,N_3514,N_3356);
and U4469 (N_4469,N_3087,N_3155);
nor U4470 (N_4470,N_3908,N_3689);
nor U4471 (N_4471,N_3688,N_3741);
nand U4472 (N_4472,N_3373,N_3482);
nand U4473 (N_4473,N_3517,N_3939);
or U4474 (N_4474,N_3961,N_3600);
nand U4475 (N_4475,N_3911,N_3492);
xnor U4476 (N_4476,N_3481,N_3466);
xor U4477 (N_4477,N_3803,N_3879);
xnor U4478 (N_4478,N_3368,N_3304);
or U4479 (N_4479,N_3811,N_3798);
nand U4480 (N_4480,N_3979,N_3727);
or U4481 (N_4481,N_3729,N_3938);
or U4482 (N_4482,N_3834,N_3146);
or U4483 (N_4483,N_3671,N_3012);
nand U4484 (N_4484,N_3596,N_3206);
or U4485 (N_4485,N_3047,N_3550);
nor U4486 (N_4486,N_3383,N_3104);
nand U4487 (N_4487,N_3609,N_3548);
and U4488 (N_4488,N_3557,N_3561);
or U4489 (N_4489,N_3588,N_3030);
nor U4490 (N_4490,N_3894,N_3647);
xnor U4491 (N_4491,N_3772,N_3377);
nand U4492 (N_4492,N_3468,N_3488);
nand U4493 (N_4493,N_3706,N_3344);
nor U4494 (N_4494,N_3021,N_3507);
nand U4495 (N_4495,N_3361,N_3865);
or U4496 (N_4496,N_3855,N_3581);
nand U4497 (N_4497,N_3316,N_3181);
nand U4498 (N_4498,N_3439,N_3864);
nand U4499 (N_4499,N_3782,N_3123);
nor U4500 (N_4500,N_3477,N_3351);
or U4501 (N_4501,N_3379,N_3918);
nor U4502 (N_4502,N_3833,N_3557);
xnor U4503 (N_4503,N_3662,N_3712);
nand U4504 (N_4504,N_3764,N_3099);
nor U4505 (N_4505,N_3441,N_3152);
nor U4506 (N_4506,N_3625,N_3012);
or U4507 (N_4507,N_3257,N_3703);
nand U4508 (N_4508,N_3784,N_3318);
and U4509 (N_4509,N_3757,N_3358);
nor U4510 (N_4510,N_3169,N_3368);
xnor U4511 (N_4511,N_3423,N_3969);
and U4512 (N_4512,N_3318,N_3025);
xnor U4513 (N_4513,N_3886,N_3895);
and U4514 (N_4514,N_3621,N_3985);
nor U4515 (N_4515,N_3963,N_3410);
and U4516 (N_4516,N_3639,N_3416);
nor U4517 (N_4517,N_3069,N_3836);
xor U4518 (N_4518,N_3390,N_3868);
nand U4519 (N_4519,N_3031,N_3156);
or U4520 (N_4520,N_3885,N_3135);
nand U4521 (N_4521,N_3690,N_3224);
and U4522 (N_4522,N_3850,N_3032);
or U4523 (N_4523,N_3345,N_3847);
or U4524 (N_4524,N_3709,N_3832);
nor U4525 (N_4525,N_3960,N_3784);
and U4526 (N_4526,N_3456,N_3599);
and U4527 (N_4527,N_3814,N_3396);
nor U4528 (N_4528,N_3706,N_3160);
nand U4529 (N_4529,N_3546,N_3957);
nand U4530 (N_4530,N_3208,N_3122);
xnor U4531 (N_4531,N_3637,N_3561);
nand U4532 (N_4532,N_3843,N_3946);
nor U4533 (N_4533,N_3974,N_3172);
nor U4534 (N_4534,N_3215,N_3815);
nor U4535 (N_4535,N_3211,N_3060);
nand U4536 (N_4536,N_3888,N_3107);
nand U4537 (N_4537,N_3356,N_3982);
and U4538 (N_4538,N_3550,N_3938);
xor U4539 (N_4539,N_3513,N_3870);
or U4540 (N_4540,N_3622,N_3306);
nand U4541 (N_4541,N_3640,N_3216);
xor U4542 (N_4542,N_3824,N_3310);
and U4543 (N_4543,N_3952,N_3668);
nand U4544 (N_4544,N_3502,N_3650);
nor U4545 (N_4545,N_3275,N_3699);
and U4546 (N_4546,N_3707,N_3279);
nand U4547 (N_4547,N_3386,N_3813);
and U4548 (N_4548,N_3281,N_3006);
xnor U4549 (N_4549,N_3008,N_3426);
nand U4550 (N_4550,N_3413,N_3210);
nor U4551 (N_4551,N_3284,N_3946);
xor U4552 (N_4552,N_3805,N_3666);
nand U4553 (N_4553,N_3206,N_3768);
nand U4554 (N_4554,N_3047,N_3820);
and U4555 (N_4555,N_3380,N_3792);
nand U4556 (N_4556,N_3944,N_3361);
xor U4557 (N_4557,N_3649,N_3762);
xor U4558 (N_4558,N_3969,N_3278);
nor U4559 (N_4559,N_3841,N_3077);
nand U4560 (N_4560,N_3343,N_3415);
or U4561 (N_4561,N_3805,N_3142);
xnor U4562 (N_4562,N_3298,N_3559);
nand U4563 (N_4563,N_3796,N_3200);
and U4564 (N_4564,N_3439,N_3004);
xnor U4565 (N_4565,N_3361,N_3276);
or U4566 (N_4566,N_3382,N_3803);
xor U4567 (N_4567,N_3803,N_3766);
nand U4568 (N_4568,N_3767,N_3689);
xor U4569 (N_4569,N_3647,N_3024);
nand U4570 (N_4570,N_3484,N_3083);
nor U4571 (N_4571,N_3054,N_3609);
or U4572 (N_4572,N_3367,N_3429);
and U4573 (N_4573,N_3277,N_3818);
xor U4574 (N_4574,N_3754,N_3445);
xor U4575 (N_4575,N_3646,N_3175);
and U4576 (N_4576,N_3115,N_3122);
xnor U4577 (N_4577,N_3703,N_3671);
xnor U4578 (N_4578,N_3651,N_3522);
xnor U4579 (N_4579,N_3669,N_3936);
nor U4580 (N_4580,N_3306,N_3254);
or U4581 (N_4581,N_3927,N_3794);
or U4582 (N_4582,N_3496,N_3366);
xor U4583 (N_4583,N_3844,N_3382);
nor U4584 (N_4584,N_3033,N_3236);
nor U4585 (N_4585,N_3787,N_3159);
or U4586 (N_4586,N_3537,N_3273);
nand U4587 (N_4587,N_3961,N_3876);
or U4588 (N_4588,N_3433,N_3697);
and U4589 (N_4589,N_3894,N_3241);
nor U4590 (N_4590,N_3552,N_3310);
nand U4591 (N_4591,N_3851,N_3155);
xnor U4592 (N_4592,N_3331,N_3951);
xnor U4593 (N_4593,N_3857,N_3401);
or U4594 (N_4594,N_3832,N_3643);
nor U4595 (N_4595,N_3492,N_3391);
and U4596 (N_4596,N_3035,N_3997);
xor U4597 (N_4597,N_3466,N_3095);
or U4598 (N_4598,N_3644,N_3546);
nor U4599 (N_4599,N_3430,N_3095);
xnor U4600 (N_4600,N_3894,N_3560);
and U4601 (N_4601,N_3339,N_3057);
and U4602 (N_4602,N_3687,N_3108);
or U4603 (N_4603,N_3474,N_3097);
or U4604 (N_4604,N_3506,N_3398);
xnor U4605 (N_4605,N_3326,N_3462);
nor U4606 (N_4606,N_3920,N_3992);
nand U4607 (N_4607,N_3758,N_3424);
or U4608 (N_4608,N_3059,N_3188);
or U4609 (N_4609,N_3642,N_3702);
nand U4610 (N_4610,N_3779,N_3352);
nand U4611 (N_4611,N_3711,N_3252);
nand U4612 (N_4612,N_3291,N_3807);
or U4613 (N_4613,N_3709,N_3814);
nor U4614 (N_4614,N_3408,N_3584);
nand U4615 (N_4615,N_3586,N_3333);
nor U4616 (N_4616,N_3850,N_3772);
and U4617 (N_4617,N_3213,N_3568);
and U4618 (N_4618,N_3970,N_3865);
nor U4619 (N_4619,N_3196,N_3497);
or U4620 (N_4620,N_3160,N_3059);
or U4621 (N_4621,N_3124,N_3473);
and U4622 (N_4622,N_3588,N_3570);
nor U4623 (N_4623,N_3127,N_3635);
nand U4624 (N_4624,N_3645,N_3809);
xnor U4625 (N_4625,N_3012,N_3835);
xor U4626 (N_4626,N_3507,N_3246);
nor U4627 (N_4627,N_3067,N_3019);
nor U4628 (N_4628,N_3638,N_3998);
nand U4629 (N_4629,N_3719,N_3134);
xor U4630 (N_4630,N_3469,N_3503);
and U4631 (N_4631,N_3556,N_3017);
xor U4632 (N_4632,N_3902,N_3624);
xor U4633 (N_4633,N_3620,N_3557);
xor U4634 (N_4634,N_3661,N_3373);
xnor U4635 (N_4635,N_3371,N_3749);
nor U4636 (N_4636,N_3756,N_3295);
and U4637 (N_4637,N_3779,N_3584);
nor U4638 (N_4638,N_3292,N_3754);
nand U4639 (N_4639,N_3165,N_3771);
and U4640 (N_4640,N_3852,N_3114);
nor U4641 (N_4641,N_3471,N_3636);
nand U4642 (N_4642,N_3446,N_3888);
nand U4643 (N_4643,N_3892,N_3890);
nand U4644 (N_4644,N_3207,N_3340);
nor U4645 (N_4645,N_3121,N_3678);
nor U4646 (N_4646,N_3073,N_3019);
and U4647 (N_4647,N_3090,N_3943);
nor U4648 (N_4648,N_3341,N_3454);
nor U4649 (N_4649,N_3965,N_3631);
or U4650 (N_4650,N_3372,N_3551);
nand U4651 (N_4651,N_3795,N_3263);
nor U4652 (N_4652,N_3155,N_3380);
or U4653 (N_4653,N_3340,N_3878);
nand U4654 (N_4654,N_3554,N_3862);
nor U4655 (N_4655,N_3344,N_3144);
or U4656 (N_4656,N_3508,N_3721);
nand U4657 (N_4657,N_3057,N_3039);
nand U4658 (N_4658,N_3951,N_3237);
nor U4659 (N_4659,N_3228,N_3420);
nand U4660 (N_4660,N_3448,N_3026);
nor U4661 (N_4661,N_3753,N_3082);
or U4662 (N_4662,N_3809,N_3041);
xor U4663 (N_4663,N_3248,N_3767);
nand U4664 (N_4664,N_3895,N_3398);
xnor U4665 (N_4665,N_3266,N_3279);
nand U4666 (N_4666,N_3922,N_3192);
nor U4667 (N_4667,N_3155,N_3833);
xor U4668 (N_4668,N_3871,N_3841);
and U4669 (N_4669,N_3422,N_3877);
xnor U4670 (N_4670,N_3838,N_3693);
or U4671 (N_4671,N_3993,N_3128);
nand U4672 (N_4672,N_3738,N_3775);
xor U4673 (N_4673,N_3831,N_3893);
nor U4674 (N_4674,N_3013,N_3658);
nand U4675 (N_4675,N_3215,N_3903);
xor U4676 (N_4676,N_3739,N_3909);
nand U4677 (N_4677,N_3142,N_3089);
xnor U4678 (N_4678,N_3360,N_3867);
or U4679 (N_4679,N_3204,N_3407);
nor U4680 (N_4680,N_3811,N_3543);
nand U4681 (N_4681,N_3817,N_3154);
or U4682 (N_4682,N_3808,N_3894);
and U4683 (N_4683,N_3421,N_3748);
or U4684 (N_4684,N_3459,N_3601);
or U4685 (N_4685,N_3023,N_3044);
xor U4686 (N_4686,N_3853,N_3659);
or U4687 (N_4687,N_3177,N_3442);
xor U4688 (N_4688,N_3979,N_3392);
nor U4689 (N_4689,N_3485,N_3037);
xnor U4690 (N_4690,N_3089,N_3009);
nor U4691 (N_4691,N_3771,N_3894);
nor U4692 (N_4692,N_3316,N_3566);
nand U4693 (N_4693,N_3513,N_3995);
and U4694 (N_4694,N_3151,N_3894);
nor U4695 (N_4695,N_3055,N_3618);
or U4696 (N_4696,N_3269,N_3285);
and U4697 (N_4697,N_3968,N_3576);
nor U4698 (N_4698,N_3679,N_3355);
and U4699 (N_4699,N_3964,N_3469);
xnor U4700 (N_4700,N_3931,N_3070);
xnor U4701 (N_4701,N_3974,N_3390);
or U4702 (N_4702,N_3548,N_3577);
xnor U4703 (N_4703,N_3993,N_3773);
and U4704 (N_4704,N_3179,N_3983);
xnor U4705 (N_4705,N_3250,N_3802);
nor U4706 (N_4706,N_3525,N_3034);
or U4707 (N_4707,N_3277,N_3627);
nor U4708 (N_4708,N_3453,N_3194);
and U4709 (N_4709,N_3137,N_3743);
nor U4710 (N_4710,N_3114,N_3685);
and U4711 (N_4711,N_3540,N_3286);
nor U4712 (N_4712,N_3267,N_3297);
and U4713 (N_4713,N_3514,N_3549);
xor U4714 (N_4714,N_3532,N_3261);
or U4715 (N_4715,N_3726,N_3320);
xor U4716 (N_4716,N_3018,N_3007);
nor U4717 (N_4717,N_3268,N_3482);
nor U4718 (N_4718,N_3751,N_3797);
nor U4719 (N_4719,N_3121,N_3504);
and U4720 (N_4720,N_3287,N_3234);
and U4721 (N_4721,N_3849,N_3071);
nor U4722 (N_4722,N_3452,N_3889);
nand U4723 (N_4723,N_3199,N_3444);
or U4724 (N_4724,N_3170,N_3239);
or U4725 (N_4725,N_3773,N_3127);
nand U4726 (N_4726,N_3495,N_3076);
and U4727 (N_4727,N_3772,N_3586);
nand U4728 (N_4728,N_3057,N_3104);
or U4729 (N_4729,N_3086,N_3681);
nor U4730 (N_4730,N_3242,N_3119);
nor U4731 (N_4731,N_3319,N_3194);
nand U4732 (N_4732,N_3847,N_3800);
xor U4733 (N_4733,N_3539,N_3033);
nor U4734 (N_4734,N_3660,N_3391);
xor U4735 (N_4735,N_3974,N_3778);
or U4736 (N_4736,N_3158,N_3354);
xor U4737 (N_4737,N_3326,N_3946);
nand U4738 (N_4738,N_3717,N_3384);
or U4739 (N_4739,N_3255,N_3040);
nor U4740 (N_4740,N_3618,N_3016);
nor U4741 (N_4741,N_3524,N_3628);
xnor U4742 (N_4742,N_3135,N_3693);
nor U4743 (N_4743,N_3258,N_3723);
nor U4744 (N_4744,N_3062,N_3944);
nand U4745 (N_4745,N_3140,N_3303);
and U4746 (N_4746,N_3671,N_3368);
nor U4747 (N_4747,N_3477,N_3605);
xnor U4748 (N_4748,N_3204,N_3471);
xor U4749 (N_4749,N_3543,N_3252);
xnor U4750 (N_4750,N_3352,N_3182);
xnor U4751 (N_4751,N_3625,N_3923);
or U4752 (N_4752,N_3360,N_3037);
nor U4753 (N_4753,N_3693,N_3483);
xnor U4754 (N_4754,N_3733,N_3741);
nor U4755 (N_4755,N_3156,N_3860);
xnor U4756 (N_4756,N_3383,N_3950);
xor U4757 (N_4757,N_3670,N_3272);
xor U4758 (N_4758,N_3119,N_3118);
xor U4759 (N_4759,N_3791,N_3672);
xor U4760 (N_4760,N_3306,N_3919);
and U4761 (N_4761,N_3435,N_3383);
and U4762 (N_4762,N_3702,N_3124);
or U4763 (N_4763,N_3386,N_3638);
and U4764 (N_4764,N_3320,N_3806);
xnor U4765 (N_4765,N_3647,N_3574);
nor U4766 (N_4766,N_3639,N_3220);
nor U4767 (N_4767,N_3417,N_3340);
and U4768 (N_4768,N_3146,N_3174);
nand U4769 (N_4769,N_3274,N_3610);
nand U4770 (N_4770,N_3290,N_3831);
or U4771 (N_4771,N_3688,N_3343);
or U4772 (N_4772,N_3014,N_3694);
nand U4773 (N_4773,N_3221,N_3841);
or U4774 (N_4774,N_3655,N_3585);
xnor U4775 (N_4775,N_3995,N_3027);
nand U4776 (N_4776,N_3004,N_3622);
nor U4777 (N_4777,N_3007,N_3304);
and U4778 (N_4778,N_3332,N_3861);
xnor U4779 (N_4779,N_3825,N_3485);
and U4780 (N_4780,N_3612,N_3203);
or U4781 (N_4781,N_3333,N_3950);
and U4782 (N_4782,N_3288,N_3559);
or U4783 (N_4783,N_3768,N_3935);
nand U4784 (N_4784,N_3690,N_3228);
or U4785 (N_4785,N_3493,N_3725);
nor U4786 (N_4786,N_3045,N_3374);
or U4787 (N_4787,N_3616,N_3463);
xor U4788 (N_4788,N_3340,N_3285);
or U4789 (N_4789,N_3800,N_3676);
nor U4790 (N_4790,N_3859,N_3910);
nor U4791 (N_4791,N_3091,N_3769);
nand U4792 (N_4792,N_3831,N_3959);
nor U4793 (N_4793,N_3015,N_3219);
and U4794 (N_4794,N_3341,N_3852);
nand U4795 (N_4795,N_3994,N_3337);
xor U4796 (N_4796,N_3568,N_3092);
nand U4797 (N_4797,N_3076,N_3986);
nand U4798 (N_4798,N_3616,N_3826);
nand U4799 (N_4799,N_3841,N_3691);
or U4800 (N_4800,N_3134,N_3729);
xnor U4801 (N_4801,N_3324,N_3197);
and U4802 (N_4802,N_3025,N_3978);
xnor U4803 (N_4803,N_3461,N_3508);
or U4804 (N_4804,N_3056,N_3789);
or U4805 (N_4805,N_3978,N_3936);
nor U4806 (N_4806,N_3796,N_3082);
or U4807 (N_4807,N_3474,N_3911);
xor U4808 (N_4808,N_3577,N_3503);
and U4809 (N_4809,N_3090,N_3792);
and U4810 (N_4810,N_3585,N_3804);
and U4811 (N_4811,N_3541,N_3909);
and U4812 (N_4812,N_3099,N_3417);
and U4813 (N_4813,N_3910,N_3227);
nand U4814 (N_4814,N_3814,N_3255);
and U4815 (N_4815,N_3466,N_3016);
and U4816 (N_4816,N_3000,N_3971);
and U4817 (N_4817,N_3230,N_3462);
xnor U4818 (N_4818,N_3383,N_3932);
and U4819 (N_4819,N_3199,N_3907);
and U4820 (N_4820,N_3509,N_3758);
nor U4821 (N_4821,N_3946,N_3335);
and U4822 (N_4822,N_3628,N_3069);
or U4823 (N_4823,N_3315,N_3152);
nand U4824 (N_4824,N_3732,N_3601);
and U4825 (N_4825,N_3722,N_3388);
nand U4826 (N_4826,N_3401,N_3310);
or U4827 (N_4827,N_3773,N_3204);
xnor U4828 (N_4828,N_3518,N_3123);
nand U4829 (N_4829,N_3190,N_3305);
or U4830 (N_4830,N_3266,N_3827);
nand U4831 (N_4831,N_3496,N_3991);
nor U4832 (N_4832,N_3720,N_3967);
nor U4833 (N_4833,N_3825,N_3823);
and U4834 (N_4834,N_3328,N_3600);
and U4835 (N_4835,N_3349,N_3586);
nand U4836 (N_4836,N_3746,N_3686);
nor U4837 (N_4837,N_3450,N_3382);
xor U4838 (N_4838,N_3269,N_3908);
and U4839 (N_4839,N_3450,N_3970);
and U4840 (N_4840,N_3105,N_3340);
nand U4841 (N_4841,N_3098,N_3483);
or U4842 (N_4842,N_3629,N_3301);
or U4843 (N_4843,N_3431,N_3365);
xnor U4844 (N_4844,N_3976,N_3500);
nor U4845 (N_4845,N_3158,N_3372);
nor U4846 (N_4846,N_3873,N_3572);
nor U4847 (N_4847,N_3355,N_3762);
nor U4848 (N_4848,N_3196,N_3527);
nand U4849 (N_4849,N_3859,N_3240);
nor U4850 (N_4850,N_3986,N_3702);
xnor U4851 (N_4851,N_3258,N_3709);
or U4852 (N_4852,N_3854,N_3313);
xor U4853 (N_4853,N_3048,N_3990);
nand U4854 (N_4854,N_3339,N_3945);
or U4855 (N_4855,N_3991,N_3705);
xor U4856 (N_4856,N_3861,N_3755);
or U4857 (N_4857,N_3084,N_3875);
nand U4858 (N_4858,N_3423,N_3857);
xnor U4859 (N_4859,N_3073,N_3467);
nor U4860 (N_4860,N_3349,N_3702);
nand U4861 (N_4861,N_3857,N_3008);
or U4862 (N_4862,N_3295,N_3434);
nand U4863 (N_4863,N_3259,N_3068);
nand U4864 (N_4864,N_3325,N_3938);
nor U4865 (N_4865,N_3635,N_3859);
xnor U4866 (N_4866,N_3186,N_3692);
or U4867 (N_4867,N_3431,N_3221);
nand U4868 (N_4868,N_3639,N_3025);
nor U4869 (N_4869,N_3508,N_3066);
nor U4870 (N_4870,N_3695,N_3546);
or U4871 (N_4871,N_3130,N_3760);
and U4872 (N_4872,N_3427,N_3215);
and U4873 (N_4873,N_3279,N_3109);
nand U4874 (N_4874,N_3561,N_3299);
nand U4875 (N_4875,N_3734,N_3765);
or U4876 (N_4876,N_3326,N_3763);
xor U4877 (N_4877,N_3304,N_3542);
and U4878 (N_4878,N_3420,N_3122);
xor U4879 (N_4879,N_3794,N_3966);
or U4880 (N_4880,N_3935,N_3366);
xnor U4881 (N_4881,N_3893,N_3781);
or U4882 (N_4882,N_3857,N_3927);
nand U4883 (N_4883,N_3939,N_3091);
or U4884 (N_4884,N_3439,N_3144);
or U4885 (N_4885,N_3706,N_3950);
nor U4886 (N_4886,N_3652,N_3518);
nor U4887 (N_4887,N_3417,N_3580);
xnor U4888 (N_4888,N_3068,N_3130);
nand U4889 (N_4889,N_3494,N_3517);
nor U4890 (N_4890,N_3859,N_3802);
and U4891 (N_4891,N_3999,N_3958);
xnor U4892 (N_4892,N_3267,N_3204);
nand U4893 (N_4893,N_3469,N_3275);
xnor U4894 (N_4894,N_3184,N_3053);
nand U4895 (N_4895,N_3944,N_3253);
nand U4896 (N_4896,N_3475,N_3683);
and U4897 (N_4897,N_3186,N_3262);
or U4898 (N_4898,N_3019,N_3587);
or U4899 (N_4899,N_3097,N_3543);
nand U4900 (N_4900,N_3446,N_3218);
and U4901 (N_4901,N_3259,N_3282);
xnor U4902 (N_4902,N_3349,N_3424);
or U4903 (N_4903,N_3063,N_3532);
or U4904 (N_4904,N_3800,N_3254);
and U4905 (N_4905,N_3283,N_3476);
or U4906 (N_4906,N_3146,N_3353);
nand U4907 (N_4907,N_3938,N_3228);
nor U4908 (N_4908,N_3751,N_3660);
or U4909 (N_4909,N_3636,N_3076);
xor U4910 (N_4910,N_3663,N_3723);
xnor U4911 (N_4911,N_3281,N_3453);
and U4912 (N_4912,N_3199,N_3804);
xor U4913 (N_4913,N_3822,N_3875);
nand U4914 (N_4914,N_3707,N_3130);
nand U4915 (N_4915,N_3584,N_3637);
xnor U4916 (N_4916,N_3947,N_3317);
nor U4917 (N_4917,N_3999,N_3913);
xnor U4918 (N_4918,N_3442,N_3997);
or U4919 (N_4919,N_3357,N_3923);
and U4920 (N_4920,N_3694,N_3635);
or U4921 (N_4921,N_3625,N_3588);
or U4922 (N_4922,N_3501,N_3865);
nand U4923 (N_4923,N_3787,N_3219);
nand U4924 (N_4924,N_3587,N_3748);
and U4925 (N_4925,N_3771,N_3102);
and U4926 (N_4926,N_3116,N_3683);
nand U4927 (N_4927,N_3485,N_3105);
xor U4928 (N_4928,N_3297,N_3770);
nand U4929 (N_4929,N_3974,N_3296);
or U4930 (N_4930,N_3769,N_3472);
or U4931 (N_4931,N_3632,N_3794);
or U4932 (N_4932,N_3055,N_3015);
or U4933 (N_4933,N_3132,N_3161);
or U4934 (N_4934,N_3539,N_3486);
nor U4935 (N_4935,N_3111,N_3042);
nor U4936 (N_4936,N_3324,N_3938);
xor U4937 (N_4937,N_3682,N_3039);
or U4938 (N_4938,N_3452,N_3068);
nand U4939 (N_4939,N_3042,N_3593);
nand U4940 (N_4940,N_3612,N_3762);
nor U4941 (N_4941,N_3522,N_3858);
or U4942 (N_4942,N_3624,N_3246);
nand U4943 (N_4943,N_3381,N_3572);
and U4944 (N_4944,N_3047,N_3816);
and U4945 (N_4945,N_3393,N_3935);
nand U4946 (N_4946,N_3916,N_3328);
xnor U4947 (N_4947,N_3037,N_3981);
nand U4948 (N_4948,N_3848,N_3641);
and U4949 (N_4949,N_3218,N_3866);
and U4950 (N_4950,N_3616,N_3419);
nor U4951 (N_4951,N_3879,N_3628);
nor U4952 (N_4952,N_3546,N_3195);
nor U4953 (N_4953,N_3048,N_3860);
nand U4954 (N_4954,N_3346,N_3696);
nor U4955 (N_4955,N_3023,N_3000);
xor U4956 (N_4956,N_3874,N_3611);
and U4957 (N_4957,N_3807,N_3631);
nand U4958 (N_4958,N_3621,N_3639);
or U4959 (N_4959,N_3077,N_3264);
nand U4960 (N_4960,N_3762,N_3559);
nor U4961 (N_4961,N_3651,N_3291);
xnor U4962 (N_4962,N_3031,N_3557);
or U4963 (N_4963,N_3863,N_3774);
xor U4964 (N_4964,N_3095,N_3980);
and U4965 (N_4965,N_3356,N_3551);
and U4966 (N_4966,N_3513,N_3193);
and U4967 (N_4967,N_3546,N_3708);
nor U4968 (N_4968,N_3794,N_3196);
and U4969 (N_4969,N_3247,N_3287);
nand U4970 (N_4970,N_3967,N_3860);
and U4971 (N_4971,N_3707,N_3486);
nand U4972 (N_4972,N_3791,N_3873);
or U4973 (N_4973,N_3341,N_3368);
or U4974 (N_4974,N_3056,N_3303);
or U4975 (N_4975,N_3377,N_3714);
or U4976 (N_4976,N_3358,N_3944);
nor U4977 (N_4977,N_3859,N_3419);
nand U4978 (N_4978,N_3095,N_3152);
or U4979 (N_4979,N_3949,N_3098);
xnor U4980 (N_4980,N_3930,N_3247);
and U4981 (N_4981,N_3815,N_3685);
xnor U4982 (N_4982,N_3464,N_3492);
nor U4983 (N_4983,N_3805,N_3698);
nand U4984 (N_4984,N_3560,N_3864);
or U4985 (N_4985,N_3312,N_3939);
or U4986 (N_4986,N_3882,N_3581);
or U4987 (N_4987,N_3692,N_3740);
nor U4988 (N_4988,N_3669,N_3760);
xor U4989 (N_4989,N_3779,N_3426);
and U4990 (N_4990,N_3281,N_3968);
and U4991 (N_4991,N_3657,N_3783);
xnor U4992 (N_4992,N_3808,N_3756);
nor U4993 (N_4993,N_3973,N_3398);
nand U4994 (N_4994,N_3151,N_3920);
and U4995 (N_4995,N_3423,N_3697);
and U4996 (N_4996,N_3348,N_3871);
nand U4997 (N_4997,N_3967,N_3853);
nand U4998 (N_4998,N_3033,N_3548);
or U4999 (N_4999,N_3312,N_3494);
and U5000 (N_5000,N_4390,N_4513);
nor U5001 (N_5001,N_4285,N_4635);
nand U5002 (N_5002,N_4738,N_4252);
xor U5003 (N_5003,N_4916,N_4152);
nand U5004 (N_5004,N_4510,N_4672);
xnor U5005 (N_5005,N_4524,N_4028);
and U5006 (N_5006,N_4288,N_4169);
and U5007 (N_5007,N_4348,N_4243);
xnor U5008 (N_5008,N_4291,N_4080);
nor U5009 (N_5009,N_4921,N_4257);
xnor U5010 (N_5010,N_4532,N_4332);
nand U5011 (N_5011,N_4274,N_4231);
xnor U5012 (N_5012,N_4782,N_4572);
or U5013 (N_5013,N_4036,N_4729);
or U5014 (N_5014,N_4439,N_4586);
xor U5015 (N_5015,N_4888,N_4181);
nand U5016 (N_5016,N_4937,N_4872);
and U5017 (N_5017,N_4177,N_4382);
nand U5018 (N_5018,N_4870,N_4170);
or U5019 (N_5019,N_4123,N_4262);
or U5020 (N_5020,N_4137,N_4237);
and U5021 (N_5021,N_4587,N_4551);
xnor U5022 (N_5022,N_4717,N_4681);
and U5023 (N_5023,N_4141,N_4780);
nor U5024 (N_5024,N_4037,N_4136);
xor U5025 (N_5025,N_4418,N_4887);
nand U5026 (N_5026,N_4186,N_4676);
and U5027 (N_5027,N_4135,N_4666);
nor U5028 (N_5028,N_4880,N_4634);
nor U5029 (N_5029,N_4308,N_4961);
xnor U5030 (N_5030,N_4515,N_4578);
or U5031 (N_5031,N_4046,N_4986);
nor U5032 (N_5032,N_4316,N_4310);
nand U5033 (N_5033,N_4817,N_4263);
and U5034 (N_5034,N_4727,N_4984);
or U5035 (N_5035,N_4172,N_4402);
nand U5036 (N_5036,N_4523,N_4313);
nor U5037 (N_5037,N_4525,N_4142);
nor U5038 (N_5038,N_4460,N_4454);
or U5039 (N_5039,N_4703,N_4520);
nand U5040 (N_5040,N_4816,N_4314);
or U5041 (N_5041,N_4254,N_4009);
or U5042 (N_5042,N_4238,N_4395);
xor U5043 (N_5043,N_4709,N_4248);
nor U5044 (N_5044,N_4176,N_4743);
or U5045 (N_5045,N_4424,N_4035);
and U5046 (N_5046,N_4095,N_4832);
and U5047 (N_5047,N_4958,N_4844);
nand U5048 (N_5048,N_4155,N_4718);
and U5049 (N_5049,N_4479,N_4754);
and U5050 (N_5050,N_4531,N_4350);
nand U5051 (N_5051,N_4226,N_4450);
nor U5052 (N_5052,N_4292,N_4922);
xnor U5053 (N_5053,N_4680,N_4850);
nand U5054 (N_5054,N_4442,N_4858);
or U5055 (N_5055,N_4225,N_4140);
nand U5056 (N_5056,N_4998,N_4069);
nor U5057 (N_5057,N_4939,N_4857);
nand U5058 (N_5058,N_4804,N_4309);
and U5059 (N_5059,N_4052,N_4983);
or U5060 (N_5060,N_4331,N_4210);
or U5061 (N_5061,N_4456,N_4938);
or U5062 (N_5062,N_4664,N_4497);
xor U5063 (N_5063,N_4247,N_4843);
xor U5064 (N_5064,N_4988,N_4603);
and U5065 (N_5065,N_4621,N_4649);
and U5066 (N_5066,N_4847,N_4143);
or U5067 (N_5067,N_4647,N_4588);
or U5068 (N_5068,N_4642,N_4926);
nor U5069 (N_5069,N_4550,N_4187);
or U5070 (N_5070,N_4777,N_4835);
and U5071 (N_5071,N_4697,N_4781);
or U5072 (N_5072,N_4656,N_4559);
nor U5073 (N_5073,N_4144,N_4400);
xnor U5074 (N_5074,N_4056,N_4971);
and U5075 (N_5075,N_4895,N_4467);
or U5076 (N_5076,N_4597,N_4084);
xnor U5077 (N_5077,N_4150,N_4808);
or U5078 (N_5078,N_4976,N_4256);
xor U5079 (N_5079,N_4665,N_4004);
nand U5080 (N_5080,N_4792,N_4434);
nor U5081 (N_5081,N_4326,N_4211);
nand U5082 (N_5082,N_4749,N_4432);
and U5083 (N_5083,N_4512,N_4890);
xor U5084 (N_5084,N_4742,N_4327);
nor U5085 (N_5085,N_4740,N_4829);
xor U5086 (N_5086,N_4825,N_4357);
and U5087 (N_5087,N_4239,N_4463);
nor U5088 (N_5088,N_4625,N_4616);
nor U5089 (N_5089,N_4813,N_4700);
nand U5090 (N_5090,N_4721,N_4407);
nor U5091 (N_5091,N_4093,N_4810);
nor U5092 (N_5092,N_4277,N_4077);
nor U5093 (N_5093,N_4115,N_4272);
nand U5094 (N_5094,N_4934,N_4695);
or U5095 (N_5095,N_4065,N_4959);
and U5096 (N_5096,N_4801,N_4392);
xor U5097 (N_5097,N_4509,N_4762);
nor U5098 (N_5098,N_4250,N_4406);
xnor U5099 (N_5099,N_4125,N_4923);
or U5100 (N_5100,N_4446,N_4683);
and U5101 (N_5101,N_4519,N_4105);
xor U5102 (N_5102,N_4799,N_4942);
nor U5103 (N_5103,N_4173,N_4894);
or U5104 (N_5104,N_4675,N_4386);
nand U5105 (N_5105,N_4655,N_4929);
nor U5106 (N_5106,N_4025,N_4469);
xnor U5107 (N_5107,N_4734,N_4241);
nor U5108 (N_5108,N_4830,N_4063);
and U5109 (N_5109,N_4162,N_4818);
or U5110 (N_5110,N_4696,N_4871);
or U5111 (N_5111,N_4295,N_4851);
nor U5112 (N_5112,N_4416,N_4071);
xor U5113 (N_5113,N_4911,N_4472);
xor U5114 (N_5114,N_4459,N_4444);
or U5115 (N_5115,N_4103,N_4537);
and U5116 (N_5116,N_4184,N_4637);
xnor U5117 (N_5117,N_4540,N_4965);
nand U5118 (N_5118,N_4278,N_4798);
and U5119 (N_5119,N_4158,N_4601);
or U5120 (N_5120,N_4583,N_4405);
nor U5121 (N_5121,N_4716,N_4950);
xnor U5122 (N_5122,N_4388,N_4945);
nand U5123 (N_5123,N_4110,N_4766);
xor U5124 (N_5124,N_4997,N_4612);
or U5125 (N_5125,N_4199,N_4318);
or U5126 (N_5126,N_4806,N_4599);
or U5127 (N_5127,N_4340,N_4306);
xnor U5128 (N_5128,N_4209,N_4555);
xnor U5129 (N_5129,N_4062,N_4886);
nor U5130 (N_5130,N_4974,N_4149);
xnor U5131 (N_5131,N_4884,N_4722);
xor U5132 (N_5132,N_4374,N_4329);
or U5133 (N_5133,N_4437,N_4617);
nor U5134 (N_5134,N_4061,N_4417);
nor U5135 (N_5135,N_4365,N_4967);
or U5136 (N_5136,N_4013,N_4016);
and U5137 (N_5137,N_4809,N_4842);
or U5138 (N_5138,N_4828,N_4498);
nor U5139 (N_5139,N_4440,N_4622);
xor U5140 (N_5140,N_4193,N_4678);
or U5141 (N_5141,N_4552,N_4714);
or U5142 (N_5142,N_4848,N_4478);
and U5143 (N_5143,N_4748,N_4430);
or U5144 (N_5144,N_4558,N_4756);
xor U5145 (N_5145,N_4644,N_4097);
nor U5146 (N_5146,N_4146,N_4132);
or U5147 (N_5147,N_4246,N_4452);
and U5148 (N_5148,N_4427,N_4885);
xor U5149 (N_5149,N_4117,N_4234);
xnor U5150 (N_5150,N_4863,N_4381);
nor U5151 (N_5151,N_4630,N_4204);
or U5152 (N_5152,N_4529,N_4701);
and U5153 (N_5153,N_4221,N_4378);
xor U5154 (N_5154,N_4739,N_4770);
nor U5155 (N_5155,N_4827,N_4541);
and U5156 (N_5156,N_4667,N_4445);
xnor U5157 (N_5157,N_4893,N_4133);
nor U5158 (N_5158,N_4567,N_4038);
or U5159 (N_5159,N_4506,N_4571);
and U5160 (N_5160,N_4026,N_4927);
or U5161 (N_5161,N_4546,N_4995);
or U5162 (N_5162,N_4342,N_4092);
nand U5163 (N_5163,N_4200,N_4154);
nor U5164 (N_5164,N_4129,N_4436);
xor U5165 (N_5165,N_4289,N_4359);
and U5166 (N_5166,N_4408,N_4414);
xnor U5167 (N_5167,N_4244,N_4494);
nand U5168 (N_5168,N_4966,N_4556);
and U5169 (N_5169,N_4480,N_4981);
nor U5170 (N_5170,N_4090,N_4968);
or U5171 (N_5171,N_4686,N_4705);
xnor U5172 (N_5172,N_4267,N_4131);
nand U5173 (N_5173,N_4972,N_4447);
or U5174 (N_5174,N_4502,N_4573);
xor U5175 (N_5175,N_4903,N_4702);
or U5176 (N_5176,N_4999,N_4086);
xor U5177 (N_5177,N_4048,N_4279);
and U5178 (N_5178,N_4661,N_4023);
xnor U5179 (N_5179,N_4726,N_4724);
xnor U5180 (N_5180,N_4778,N_4276);
xor U5181 (N_5181,N_4453,N_4604);
nand U5182 (N_5182,N_4865,N_4632);
and U5183 (N_5183,N_4773,N_4375);
nand U5184 (N_5184,N_4837,N_4083);
or U5185 (N_5185,N_4081,N_4130);
or U5186 (N_5186,N_4398,N_4946);
nand U5187 (N_5187,N_4167,N_4312);
and U5188 (N_5188,N_4031,N_4336);
or U5189 (N_5189,N_4220,N_4545);
xor U5190 (N_5190,N_4379,N_4539);
xnor U5191 (N_5191,N_4290,N_4600);
and U5192 (N_5192,N_4574,N_4047);
nand U5193 (N_5193,N_4643,N_4725);
nand U5194 (N_5194,N_4483,N_4528);
and U5195 (N_5195,N_4070,N_4297);
nand U5196 (N_5196,N_4042,N_4373);
nand U5197 (N_5197,N_4906,N_4055);
xor U5198 (N_5198,N_4753,N_4345);
and U5199 (N_5199,N_4917,N_4521);
and U5200 (N_5200,N_4698,N_4982);
or U5201 (N_5201,N_4299,N_4153);
and U5202 (N_5202,N_4836,N_4613);
nor U5203 (N_5203,N_4859,N_4720);
or U5204 (N_5204,N_4230,N_4100);
or U5205 (N_5205,N_4180,N_4928);
and U5206 (N_5206,N_4569,N_4404);
xnor U5207 (N_5207,N_4811,N_4735);
or U5208 (N_5208,N_4334,N_4205);
nor U5209 (N_5209,N_4122,N_4298);
nor U5210 (N_5210,N_4197,N_4800);
nand U5211 (N_5211,N_4328,N_4898);
and U5212 (N_5212,N_4860,N_4017);
or U5213 (N_5213,N_4323,N_4607);
xnor U5214 (N_5214,N_4987,N_4628);
xor U5215 (N_5215,N_4012,N_4458);
nand U5216 (N_5216,N_4905,N_4296);
nor U5217 (N_5217,N_4228,N_4420);
nor U5218 (N_5218,N_4448,N_4320);
xnor U5219 (N_5219,N_4783,N_4779);
nand U5220 (N_5220,N_4639,N_4692);
xor U5221 (N_5221,N_4371,N_4774);
nor U5222 (N_5222,N_4339,N_4087);
or U5223 (N_5223,N_4719,N_4271);
xor U5224 (N_5224,N_4235,N_4875);
nor U5225 (N_5225,N_4183,N_4864);
and U5226 (N_5226,N_4422,N_4768);
xnor U5227 (N_5227,N_4208,N_4824);
or U5228 (N_5228,N_4251,N_4912);
and U5229 (N_5229,N_4213,N_4560);
xor U5230 (N_5230,N_4648,N_4301);
nor U5231 (N_5231,N_4820,N_4699);
xnor U5232 (N_5232,N_4608,N_4951);
or U5233 (N_5233,N_4954,N_4415);
nor U5234 (N_5234,N_4947,N_4641);
and U5235 (N_5235,N_4687,N_4901);
xor U5236 (N_5236,N_4088,N_4078);
or U5237 (N_5237,N_4490,N_4147);
or U5238 (N_5238,N_4980,N_4428);
and U5239 (N_5239,N_4401,N_4669);
and U5240 (N_5240,N_4102,N_4387);
and U5241 (N_5241,N_4451,N_4011);
and U5242 (N_5242,N_4112,N_4054);
nand U5243 (N_5243,N_4684,N_4812);
xor U5244 (N_5244,N_4557,N_4711);
xor U5245 (N_5245,N_4931,N_4629);
and U5246 (N_5246,N_4367,N_4505);
nand U5247 (N_5247,N_4554,N_4157);
and U5248 (N_5248,N_4736,N_4041);
or U5249 (N_5249,N_4355,N_4646);
or U5250 (N_5250,N_4178,N_4443);
and U5251 (N_5251,N_4626,N_4281);
nand U5252 (N_5252,N_4996,N_4412);
nor U5253 (N_5253,N_4366,N_4021);
or U5254 (N_5254,N_4364,N_4099);
or U5255 (N_5255,N_4384,N_4882);
nand U5256 (N_5256,N_4032,N_4685);
xnor U5257 (N_5257,N_4689,N_4435);
and U5258 (N_5258,N_4145,N_4485);
nand U5259 (N_5259,N_4192,N_4815);
nor U5260 (N_5260,N_4068,N_4764);
nand U5261 (N_5261,N_4772,N_4470);
xnor U5262 (N_5262,N_4826,N_4671);
or U5263 (N_5263,N_4438,N_4191);
nand U5264 (N_5264,N_4960,N_4148);
xnor U5265 (N_5265,N_4091,N_4807);
nand U5266 (N_5266,N_4000,N_4179);
nand U5267 (N_5267,N_4232,N_4050);
or U5268 (N_5268,N_4462,N_4846);
xor U5269 (N_5269,N_4253,N_4360);
nor U5270 (N_5270,N_4730,N_4581);
nor U5271 (N_5271,N_4659,N_4979);
or U5272 (N_5272,N_4611,N_4330);
or U5273 (N_5273,N_4259,N_4198);
or U5274 (N_5274,N_4631,N_4341);
xnor U5275 (N_5275,N_4358,N_4707);
nand U5276 (N_5276,N_4838,N_4185);
and U5277 (N_5277,N_4431,N_4589);
and U5278 (N_5278,N_4503,N_4385);
or U5279 (N_5279,N_4879,N_4138);
and U5280 (N_5280,N_4650,N_4925);
or U5281 (N_5281,N_4005,N_4892);
nand U5282 (N_5282,N_4269,N_4166);
nor U5283 (N_5283,N_4245,N_4883);
or U5284 (N_5284,N_4171,N_4803);
nor U5285 (N_5285,N_4723,N_4118);
nor U5286 (N_5286,N_4433,N_4317);
nand U5287 (N_5287,N_4514,N_4516);
nor U5288 (N_5288,N_4473,N_4109);
nand U5289 (N_5289,N_4902,N_4457);
nand U5290 (N_5290,N_4704,N_4163);
or U5291 (N_5291,N_4214,N_4731);
nand U5292 (N_5292,N_4620,N_4508);
or U5293 (N_5293,N_4845,N_4920);
and U5294 (N_5294,N_4866,N_4106);
or U5295 (N_5295,N_4805,N_4264);
nor U5296 (N_5296,N_4370,N_4595);
and U5297 (N_5297,N_4159,N_4580);
or U5298 (N_5298,N_4027,N_4732);
nand U5299 (N_5299,N_4034,N_4862);
and U5300 (N_5300,N_4590,N_4488);
or U5301 (N_5301,N_4258,N_4001);
and U5302 (N_5302,N_4763,N_4944);
nor U5303 (N_5303,N_4303,N_4691);
nand U5304 (N_5304,N_4394,N_4900);
nor U5305 (N_5305,N_4755,N_4127);
and U5306 (N_5306,N_4814,N_4391);
and U5307 (N_5307,N_4399,N_4182);
nor U5308 (N_5308,N_4913,N_4104);
xor U5309 (N_5309,N_4195,N_4728);
nor U5310 (N_5310,N_4881,N_4854);
xnor U5311 (N_5311,N_4833,N_4582);
or U5312 (N_5312,N_4305,N_4051);
xor U5313 (N_5313,N_4821,N_4940);
or U5314 (N_5314,N_4116,N_4376);
xor U5315 (N_5315,N_4168,N_4111);
and U5316 (N_5316,N_4108,N_4565);
nand U5317 (N_5317,N_4789,N_4802);
nor U5318 (N_5318,N_4273,N_4658);
nand U5319 (N_5319,N_4561,N_4674);
nor U5320 (N_5320,N_4598,N_4349);
xor U5321 (N_5321,N_4975,N_4495);
nand U5322 (N_5322,N_4831,N_4533);
nand U5323 (N_5323,N_4955,N_4236);
nor U5324 (N_5324,N_4839,N_4134);
xnor U5325 (N_5325,N_4948,N_4287);
nand U5326 (N_5326,N_4008,N_4484);
or U5327 (N_5327,N_4060,N_4527);
xor U5328 (N_5328,N_4769,N_4352);
or U5329 (N_5329,N_4156,N_4007);
nand U5330 (N_5330,N_4215,N_4190);
nand U5331 (N_5331,N_4160,N_4429);
and U5332 (N_5332,N_4354,N_4591);
xnor U5333 (N_5333,N_4657,N_4496);
xor U5334 (N_5334,N_4227,N_4403);
nand U5335 (N_5335,N_4393,N_4899);
nand U5336 (N_5336,N_4909,N_4468);
nor U5337 (N_5337,N_4896,N_4841);
or U5338 (N_5338,N_4619,N_4098);
and U5339 (N_5339,N_4553,N_4268);
and U5340 (N_5340,N_4029,N_4936);
and U5341 (N_5341,N_4377,N_4030);
nor U5342 (N_5342,N_4823,N_4543);
and U5343 (N_5343,N_4610,N_4602);
nand U5344 (N_5344,N_4229,N_4423);
nor U5345 (N_5345,N_4522,N_4217);
or U5346 (N_5346,N_4544,N_4507);
xor U5347 (N_5347,N_4304,N_4605);
nand U5348 (N_5348,N_4526,N_4534);
nor U5349 (N_5349,N_4941,N_4175);
nor U5350 (N_5350,N_4203,N_4663);
xor U5351 (N_5351,N_4795,N_4464);
xnor U5352 (N_5352,N_4002,N_4856);
and U5353 (N_5353,N_4662,N_4489);
xor U5354 (N_5354,N_4511,N_4877);
nor U5355 (N_5355,N_4849,N_4867);
nand U5356 (N_5356,N_4346,N_4492);
and U5357 (N_5357,N_4094,N_4202);
or U5358 (N_5358,N_4380,N_4549);
and U5359 (N_5359,N_4530,N_4067);
or U5360 (N_5360,N_4410,N_4322);
nand U5361 (N_5361,N_4594,N_4189);
or U5362 (N_5362,N_4564,N_4633);
or U5363 (N_5363,N_4609,N_4425);
and U5364 (N_5364,N_4072,N_4990);
or U5365 (N_5365,N_4282,N_4618);
xor U5366 (N_5366,N_4043,N_4744);
xnor U5367 (N_5367,N_4383,N_4741);
nand U5368 (N_5368,N_4481,N_4563);
nand U5369 (N_5369,N_4889,N_4019);
and U5370 (N_5370,N_4347,N_4351);
nand U5371 (N_5371,N_4126,N_4333);
or U5372 (N_5372,N_4465,N_4338);
and U5373 (N_5373,N_4712,N_4904);
and U5374 (N_5374,N_4219,N_4690);
or U5375 (N_5375,N_4499,N_4688);
nand U5376 (N_5376,N_4861,N_4834);
and U5377 (N_5377,N_4421,N_4977);
and U5378 (N_5378,N_4280,N_4010);
nand U5379 (N_5379,N_4640,N_4461);
or U5380 (N_5380,N_4787,N_4049);
nor U5381 (N_5381,N_4670,N_4441);
nand U5382 (N_5382,N_4284,N_4784);
xor U5383 (N_5383,N_4518,N_4164);
nor U5384 (N_5384,N_4985,N_4708);
and U5385 (N_5385,N_4989,N_4015);
or U5386 (N_5386,N_4788,N_4869);
nand U5387 (N_5387,N_4372,N_4767);
and U5388 (N_5388,N_4542,N_4082);
xor U5389 (N_5389,N_4242,N_4096);
nand U5390 (N_5390,N_4915,N_4694);
nor U5391 (N_5391,N_4076,N_4786);
and U5392 (N_5392,N_4223,N_4353);
xnor U5393 (N_5393,N_4745,N_4449);
or U5394 (N_5394,N_4576,N_4040);
nand U5395 (N_5395,N_4174,N_4113);
or U5396 (N_5396,N_4878,N_4249);
xor U5397 (N_5397,N_4797,N_4891);
nand U5398 (N_5398,N_4566,N_4324);
nor U5399 (N_5399,N_4224,N_4750);
and U5400 (N_5400,N_4361,N_4579);
and U5401 (N_5401,N_4261,N_4057);
nor U5402 (N_5402,N_4079,N_4335);
nand U5403 (N_5403,N_4319,N_4119);
or U5404 (N_5404,N_4500,N_4693);
or U5405 (N_5405,N_4165,N_4957);
nor U5406 (N_5406,N_4682,N_4970);
or U5407 (N_5407,N_4538,N_4994);
xnor U5408 (N_5408,N_4233,N_4952);
xnor U5409 (N_5409,N_4652,N_4746);
nor U5410 (N_5410,N_4255,N_4907);
or U5411 (N_5411,N_4222,N_4747);
xor U5412 (N_5412,N_4300,N_4074);
xor U5413 (N_5413,N_4275,N_4466);
and U5414 (N_5414,N_4368,N_4822);
and U5415 (N_5415,N_4194,N_4897);
nand U5416 (N_5416,N_4614,N_4908);
nand U5417 (N_5417,N_4627,N_4409);
nor U5418 (N_5418,N_4064,N_4853);
xnor U5419 (N_5419,N_4973,N_4120);
or U5420 (N_5420,N_4426,N_4733);
nand U5421 (N_5421,N_4419,N_4978);
or U5422 (N_5422,N_4910,N_4638);
and U5423 (N_5423,N_4568,N_4053);
nand U5424 (N_5424,N_4024,N_4389);
xnor U5425 (N_5425,N_4039,N_4932);
nand U5426 (N_5426,N_4949,N_4033);
nor U5427 (N_5427,N_4018,N_4776);
or U5428 (N_5428,N_4311,N_4653);
or U5429 (N_5429,N_4673,N_4482);
xor U5430 (N_5430,N_4791,N_4593);
nand U5431 (N_5431,N_4216,N_4536);
or U5432 (N_5432,N_4758,N_4114);
nor U5433 (N_5433,N_4991,N_4765);
nand U5434 (N_5434,N_4501,N_4369);
nand U5435 (N_5435,N_4584,N_4188);
nand U5436 (N_5436,N_4151,N_4760);
or U5437 (N_5437,N_4260,N_4124);
and U5438 (N_5438,N_4623,N_4876);
and U5439 (N_5439,N_4286,N_4715);
xor U5440 (N_5440,N_4562,N_4212);
xor U5441 (N_5441,N_4710,N_4636);
nor U5442 (N_5442,N_4058,N_4493);
nand U5443 (N_5443,N_4993,N_4963);
and U5444 (N_5444,N_4266,N_4796);
nor U5445 (N_5445,N_4855,N_4679);
nand U5446 (N_5446,N_4592,N_4362);
and U5447 (N_5447,N_4014,N_4486);
and U5448 (N_5448,N_4073,N_4321);
xor U5449 (N_5449,N_4547,N_4411);
or U5450 (N_5450,N_4840,N_4660);
nand U5451 (N_5451,N_4668,N_4852);
and U5452 (N_5452,N_4022,N_4962);
or U5453 (N_5453,N_4356,N_4476);
xor U5454 (N_5454,N_4161,N_4517);
nand U5455 (N_5455,N_4914,N_4477);
xnor U5456 (N_5456,N_4307,N_4874);
and U5457 (N_5457,N_4752,N_4956);
and U5458 (N_5458,N_4651,N_4785);
nor U5459 (N_5459,N_4771,N_4196);
nor U5460 (N_5460,N_4059,N_4455);
xnor U5461 (N_5461,N_4487,N_4101);
xor U5462 (N_5462,N_4294,N_4868);
nor U5463 (N_5463,N_4570,N_4003);
and U5464 (N_5464,N_4873,N_4793);
nor U5465 (N_5465,N_4413,N_4270);
nand U5466 (N_5466,N_4240,N_4089);
nand U5467 (N_5467,N_4964,N_4471);
xnor U5468 (N_5468,N_4535,N_4128);
and U5469 (N_5469,N_4759,N_4992);
nand U5470 (N_5470,N_4677,N_4751);
or U5471 (N_5471,N_4085,N_4302);
nor U5472 (N_5472,N_4344,N_4713);
xor U5473 (N_5473,N_4325,N_4397);
nand U5474 (N_5474,N_4761,N_4206);
nor U5475 (N_5475,N_4596,N_4575);
xnor U5476 (N_5476,N_4918,N_4606);
or U5477 (N_5477,N_4066,N_4107);
and U5478 (N_5478,N_4315,N_4645);
nand U5479 (N_5479,N_4474,N_4218);
or U5480 (N_5480,N_4943,N_4737);
nor U5481 (N_5481,N_4283,N_4775);
xnor U5482 (N_5482,N_4006,N_4139);
nand U5483 (N_5483,N_4045,N_4396);
and U5484 (N_5484,N_4337,N_4293);
nor U5485 (N_5485,N_4819,N_4121);
or U5486 (N_5486,N_4504,N_4201);
or U5487 (N_5487,N_4265,N_4794);
nand U5488 (N_5488,N_4930,N_4044);
xnor U5489 (N_5489,N_4585,N_4953);
or U5490 (N_5490,N_4933,N_4935);
xnor U5491 (N_5491,N_4757,N_4790);
and U5492 (N_5492,N_4075,N_4207);
nand U5493 (N_5493,N_4343,N_4969);
nand U5494 (N_5494,N_4363,N_4706);
and U5495 (N_5495,N_4020,N_4548);
or U5496 (N_5496,N_4919,N_4577);
and U5497 (N_5497,N_4491,N_4624);
or U5498 (N_5498,N_4924,N_4475);
or U5499 (N_5499,N_4615,N_4654);
xnor U5500 (N_5500,N_4026,N_4360);
or U5501 (N_5501,N_4178,N_4865);
nand U5502 (N_5502,N_4027,N_4207);
or U5503 (N_5503,N_4409,N_4658);
and U5504 (N_5504,N_4823,N_4925);
xor U5505 (N_5505,N_4420,N_4936);
nand U5506 (N_5506,N_4407,N_4394);
or U5507 (N_5507,N_4723,N_4726);
xor U5508 (N_5508,N_4780,N_4254);
and U5509 (N_5509,N_4700,N_4889);
xor U5510 (N_5510,N_4543,N_4714);
nor U5511 (N_5511,N_4289,N_4807);
nand U5512 (N_5512,N_4235,N_4005);
nor U5513 (N_5513,N_4027,N_4956);
xor U5514 (N_5514,N_4659,N_4868);
nor U5515 (N_5515,N_4111,N_4205);
xnor U5516 (N_5516,N_4101,N_4916);
nor U5517 (N_5517,N_4649,N_4305);
and U5518 (N_5518,N_4303,N_4663);
nor U5519 (N_5519,N_4139,N_4792);
nor U5520 (N_5520,N_4920,N_4930);
xor U5521 (N_5521,N_4596,N_4222);
and U5522 (N_5522,N_4810,N_4529);
nor U5523 (N_5523,N_4486,N_4616);
and U5524 (N_5524,N_4098,N_4109);
and U5525 (N_5525,N_4685,N_4528);
nand U5526 (N_5526,N_4314,N_4119);
and U5527 (N_5527,N_4999,N_4117);
nor U5528 (N_5528,N_4047,N_4521);
or U5529 (N_5529,N_4905,N_4128);
and U5530 (N_5530,N_4289,N_4411);
or U5531 (N_5531,N_4380,N_4234);
or U5532 (N_5532,N_4835,N_4327);
and U5533 (N_5533,N_4828,N_4347);
xor U5534 (N_5534,N_4466,N_4096);
xor U5535 (N_5535,N_4265,N_4670);
xor U5536 (N_5536,N_4389,N_4182);
nor U5537 (N_5537,N_4304,N_4784);
and U5538 (N_5538,N_4872,N_4180);
nand U5539 (N_5539,N_4124,N_4214);
nand U5540 (N_5540,N_4344,N_4188);
or U5541 (N_5541,N_4296,N_4258);
nand U5542 (N_5542,N_4963,N_4687);
nor U5543 (N_5543,N_4504,N_4037);
xor U5544 (N_5544,N_4650,N_4360);
nor U5545 (N_5545,N_4019,N_4113);
or U5546 (N_5546,N_4926,N_4520);
xor U5547 (N_5547,N_4392,N_4810);
xnor U5548 (N_5548,N_4190,N_4235);
nor U5549 (N_5549,N_4255,N_4177);
or U5550 (N_5550,N_4330,N_4981);
or U5551 (N_5551,N_4125,N_4116);
nor U5552 (N_5552,N_4123,N_4603);
or U5553 (N_5553,N_4268,N_4137);
xnor U5554 (N_5554,N_4510,N_4993);
nand U5555 (N_5555,N_4970,N_4159);
xnor U5556 (N_5556,N_4594,N_4134);
nand U5557 (N_5557,N_4556,N_4421);
or U5558 (N_5558,N_4864,N_4766);
nand U5559 (N_5559,N_4820,N_4292);
xnor U5560 (N_5560,N_4391,N_4573);
xor U5561 (N_5561,N_4538,N_4509);
nand U5562 (N_5562,N_4594,N_4517);
and U5563 (N_5563,N_4880,N_4358);
or U5564 (N_5564,N_4519,N_4903);
nand U5565 (N_5565,N_4926,N_4301);
nand U5566 (N_5566,N_4378,N_4048);
nor U5567 (N_5567,N_4469,N_4720);
xor U5568 (N_5568,N_4488,N_4194);
nand U5569 (N_5569,N_4560,N_4816);
xor U5570 (N_5570,N_4768,N_4377);
nor U5571 (N_5571,N_4235,N_4824);
nor U5572 (N_5572,N_4173,N_4731);
or U5573 (N_5573,N_4898,N_4737);
or U5574 (N_5574,N_4100,N_4481);
nor U5575 (N_5575,N_4251,N_4906);
xor U5576 (N_5576,N_4522,N_4107);
nand U5577 (N_5577,N_4195,N_4820);
xor U5578 (N_5578,N_4910,N_4903);
nor U5579 (N_5579,N_4970,N_4271);
and U5580 (N_5580,N_4134,N_4468);
and U5581 (N_5581,N_4799,N_4700);
xor U5582 (N_5582,N_4393,N_4397);
xor U5583 (N_5583,N_4582,N_4487);
xnor U5584 (N_5584,N_4590,N_4140);
and U5585 (N_5585,N_4099,N_4809);
or U5586 (N_5586,N_4389,N_4797);
or U5587 (N_5587,N_4547,N_4638);
and U5588 (N_5588,N_4992,N_4113);
and U5589 (N_5589,N_4271,N_4161);
and U5590 (N_5590,N_4362,N_4013);
nor U5591 (N_5591,N_4481,N_4113);
or U5592 (N_5592,N_4836,N_4029);
or U5593 (N_5593,N_4604,N_4276);
and U5594 (N_5594,N_4228,N_4778);
and U5595 (N_5595,N_4428,N_4432);
and U5596 (N_5596,N_4013,N_4384);
xor U5597 (N_5597,N_4840,N_4464);
nor U5598 (N_5598,N_4215,N_4761);
and U5599 (N_5599,N_4594,N_4192);
and U5600 (N_5600,N_4557,N_4171);
nor U5601 (N_5601,N_4956,N_4670);
nand U5602 (N_5602,N_4429,N_4383);
xnor U5603 (N_5603,N_4407,N_4302);
nand U5604 (N_5604,N_4466,N_4835);
nand U5605 (N_5605,N_4926,N_4281);
nor U5606 (N_5606,N_4233,N_4338);
or U5607 (N_5607,N_4830,N_4413);
xor U5608 (N_5608,N_4980,N_4139);
and U5609 (N_5609,N_4528,N_4373);
or U5610 (N_5610,N_4271,N_4117);
nand U5611 (N_5611,N_4887,N_4896);
nor U5612 (N_5612,N_4146,N_4307);
xnor U5613 (N_5613,N_4351,N_4653);
or U5614 (N_5614,N_4534,N_4289);
nor U5615 (N_5615,N_4527,N_4228);
and U5616 (N_5616,N_4962,N_4970);
and U5617 (N_5617,N_4400,N_4338);
xnor U5618 (N_5618,N_4085,N_4665);
or U5619 (N_5619,N_4896,N_4569);
or U5620 (N_5620,N_4834,N_4441);
nor U5621 (N_5621,N_4027,N_4253);
nor U5622 (N_5622,N_4063,N_4442);
xor U5623 (N_5623,N_4795,N_4347);
and U5624 (N_5624,N_4361,N_4243);
nand U5625 (N_5625,N_4767,N_4528);
nand U5626 (N_5626,N_4804,N_4159);
xnor U5627 (N_5627,N_4520,N_4646);
xnor U5628 (N_5628,N_4945,N_4903);
nand U5629 (N_5629,N_4468,N_4348);
nor U5630 (N_5630,N_4056,N_4320);
and U5631 (N_5631,N_4407,N_4718);
and U5632 (N_5632,N_4340,N_4044);
nand U5633 (N_5633,N_4944,N_4461);
xor U5634 (N_5634,N_4291,N_4713);
nand U5635 (N_5635,N_4004,N_4763);
nand U5636 (N_5636,N_4902,N_4023);
and U5637 (N_5637,N_4740,N_4746);
xor U5638 (N_5638,N_4427,N_4556);
nand U5639 (N_5639,N_4601,N_4386);
nand U5640 (N_5640,N_4658,N_4382);
or U5641 (N_5641,N_4173,N_4762);
and U5642 (N_5642,N_4109,N_4760);
and U5643 (N_5643,N_4682,N_4735);
nor U5644 (N_5644,N_4681,N_4635);
and U5645 (N_5645,N_4750,N_4841);
xnor U5646 (N_5646,N_4559,N_4155);
nor U5647 (N_5647,N_4861,N_4518);
nand U5648 (N_5648,N_4122,N_4265);
and U5649 (N_5649,N_4735,N_4196);
nor U5650 (N_5650,N_4228,N_4247);
and U5651 (N_5651,N_4591,N_4162);
and U5652 (N_5652,N_4773,N_4359);
nor U5653 (N_5653,N_4852,N_4897);
nand U5654 (N_5654,N_4723,N_4203);
nand U5655 (N_5655,N_4701,N_4164);
and U5656 (N_5656,N_4427,N_4779);
or U5657 (N_5657,N_4738,N_4499);
nor U5658 (N_5658,N_4873,N_4668);
xnor U5659 (N_5659,N_4207,N_4825);
or U5660 (N_5660,N_4957,N_4629);
nand U5661 (N_5661,N_4476,N_4532);
and U5662 (N_5662,N_4950,N_4546);
nor U5663 (N_5663,N_4156,N_4562);
or U5664 (N_5664,N_4842,N_4909);
xnor U5665 (N_5665,N_4808,N_4912);
or U5666 (N_5666,N_4383,N_4761);
xor U5667 (N_5667,N_4266,N_4359);
xnor U5668 (N_5668,N_4162,N_4059);
nand U5669 (N_5669,N_4082,N_4935);
or U5670 (N_5670,N_4688,N_4412);
and U5671 (N_5671,N_4690,N_4909);
nand U5672 (N_5672,N_4151,N_4187);
nor U5673 (N_5673,N_4422,N_4888);
and U5674 (N_5674,N_4202,N_4018);
and U5675 (N_5675,N_4185,N_4520);
nand U5676 (N_5676,N_4365,N_4476);
and U5677 (N_5677,N_4243,N_4744);
nor U5678 (N_5678,N_4159,N_4623);
and U5679 (N_5679,N_4151,N_4504);
nand U5680 (N_5680,N_4826,N_4279);
nor U5681 (N_5681,N_4722,N_4771);
nand U5682 (N_5682,N_4471,N_4869);
nor U5683 (N_5683,N_4259,N_4315);
or U5684 (N_5684,N_4385,N_4761);
and U5685 (N_5685,N_4228,N_4122);
nor U5686 (N_5686,N_4374,N_4293);
xnor U5687 (N_5687,N_4073,N_4496);
or U5688 (N_5688,N_4631,N_4110);
nand U5689 (N_5689,N_4251,N_4274);
nor U5690 (N_5690,N_4038,N_4137);
and U5691 (N_5691,N_4448,N_4933);
nand U5692 (N_5692,N_4596,N_4643);
nor U5693 (N_5693,N_4319,N_4375);
or U5694 (N_5694,N_4515,N_4810);
and U5695 (N_5695,N_4173,N_4767);
or U5696 (N_5696,N_4732,N_4354);
nor U5697 (N_5697,N_4506,N_4347);
nand U5698 (N_5698,N_4856,N_4015);
or U5699 (N_5699,N_4970,N_4939);
nor U5700 (N_5700,N_4840,N_4778);
nor U5701 (N_5701,N_4673,N_4662);
nand U5702 (N_5702,N_4667,N_4228);
nor U5703 (N_5703,N_4858,N_4880);
xor U5704 (N_5704,N_4028,N_4541);
or U5705 (N_5705,N_4890,N_4808);
or U5706 (N_5706,N_4152,N_4909);
and U5707 (N_5707,N_4666,N_4322);
or U5708 (N_5708,N_4353,N_4303);
nor U5709 (N_5709,N_4017,N_4614);
nor U5710 (N_5710,N_4198,N_4986);
nor U5711 (N_5711,N_4823,N_4111);
and U5712 (N_5712,N_4110,N_4976);
nor U5713 (N_5713,N_4890,N_4397);
nand U5714 (N_5714,N_4592,N_4387);
nand U5715 (N_5715,N_4078,N_4045);
nand U5716 (N_5716,N_4103,N_4196);
or U5717 (N_5717,N_4147,N_4649);
and U5718 (N_5718,N_4391,N_4304);
xnor U5719 (N_5719,N_4600,N_4762);
and U5720 (N_5720,N_4884,N_4577);
or U5721 (N_5721,N_4858,N_4235);
or U5722 (N_5722,N_4048,N_4203);
nand U5723 (N_5723,N_4270,N_4163);
xor U5724 (N_5724,N_4576,N_4248);
nand U5725 (N_5725,N_4807,N_4556);
nand U5726 (N_5726,N_4616,N_4823);
nor U5727 (N_5727,N_4032,N_4910);
xnor U5728 (N_5728,N_4374,N_4392);
or U5729 (N_5729,N_4884,N_4487);
or U5730 (N_5730,N_4569,N_4797);
nand U5731 (N_5731,N_4242,N_4738);
nand U5732 (N_5732,N_4639,N_4931);
xnor U5733 (N_5733,N_4313,N_4414);
nor U5734 (N_5734,N_4872,N_4897);
nor U5735 (N_5735,N_4152,N_4389);
nand U5736 (N_5736,N_4151,N_4112);
nand U5737 (N_5737,N_4331,N_4151);
nand U5738 (N_5738,N_4512,N_4034);
nor U5739 (N_5739,N_4123,N_4524);
and U5740 (N_5740,N_4703,N_4405);
nor U5741 (N_5741,N_4491,N_4452);
or U5742 (N_5742,N_4356,N_4696);
or U5743 (N_5743,N_4297,N_4700);
xor U5744 (N_5744,N_4250,N_4480);
or U5745 (N_5745,N_4779,N_4036);
nor U5746 (N_5746,N_4048,N_4131);
nor U5747 (N_5747,N_4662,N_4771);
nor U5748 (N_5748,N_4338,N_4278);
or U5749 (N_5749,N_4663,N_4391);
and U5750 (N_5750,N_4685,N_4912);
nand U5751 (N_5751,N_4570,N_4106);
and U5752 (N_5752,N_4825,N_4773);
nand U5753 (N_5753,N_4158,N_4458);
nand U5754 (N_5754,N_4675,N_4586);
or U5755 (N_5755,N_4245,N_4386);
nand U5756 (N_5756,N_4394,N_4380);
and U5757 (N_5757,N_4475,N_4361);
and U5758 (N_5758,N_4055,N_4429);
or U5759 (N_5759,N_4957,N_4510);
or U5760 (N_5760,N_4618,N_4747);
nor U5761 (N_5761,N_4584,N_4897);
or U5762 (N_5762,N_4019,N_4432);
nand U5763 (N_5763,N_4798,N_4302);
nor U5764 (N_5764,N_4341,N_4604);
or U5765 (N_5765,N_4837,N_4265);
nor U5766 (N_5766,N_4668,N_4562);
nor U5767 (N_5767,N_4786,N_4278);
nor U5768 (N_5768,N_4810,N_4390);
or U5769 (N_5769,N_4731,N_4549);
nor U5770 (N_5770,N_4198,N_4894);
xor U5771 (N_5771,N_4284,N_4884);
and U5772 (N_5772,N_4485,N_4633);
nand U5773 (N_5773,N_4925,N_4101);
and U5774 (N_5774,N_4156,N_4529);
and U5775 (N_5775,N_4505,N_4948);
xnor U5776 (N_5776,N_4440,N_4967);
nor U5777 (N_5777,N_4937,N_4491);
nor U5778 (N_5778,N_4826,N_4883);
or U5779 (N_5779,N_4606,N_4646);
or U5780 (N_5780,N_4078,N_4076);
or U5781 (N_5781,N_4240,N_4623);
nand U5782 (N_5782,N_4320,N_4306);
and U5783 (N_5783,N_4834,N_4556);
nand U5784 (N_5784,N_4808,N_4174);
nand U5785 (N_5785,N_4214,N_4199);
xor U5786 (N_5786,N_4625,N_4632);
or U5787 (N_5787,N_4937,N_4124);
nor U5788 (N_5788,N_4423,N_4947);
nand U5789 (N_5789,N_4050,N_4324);
and U5790 (N_5790,N_4037,N_4434);
xor U5791 (N_5791,N_4323,N_4162);
nand U5792 (N_5792,N_4530,N_4184);
or U5793 (N_5793,N_4312,N_4316);
nand U5794 (N_5794,N_4035,N_4718);
nor U5795 (N_5795,N_4773,N_4334);
nor U5796 (N_5796,N_4982,N_4194);
and U5797 (N_5797,N_4657,N_4398);
nor U5798 (N_5798,N_4890,N_4078);
nand U5799 (N_5799,N_4287,N_4780);
xnor U5800 (N_5800,N_4732,N_4580);
nand U5801 (N_5801,N_4097,N_4048);
nand U5802 (N_5802,N_4129,N_4948);
nand U5803 (N_5803,N_4167,N_4030);
or U5804 (N_5804,N_4567,N_4688);
nand U5805 (N_5805,N_4658,N_4564);
nand U5806 (N_5806,N_4072,N_4466);
nor U5807 (N_5807,N_4956,N_4372);
and U5808 (N_5808,N_4536,N_4151);
xnor U5809 (N_5809,N_4681,N_4662);
xor U5810 (N_5810,N_4540,N_4766);
and U5811 (N_5811,N_4078,N_4510);
or U5812 (N_5812,N_4650,N_4812);
xnor U5813 (N_5813,N_4871,N_4172);
nand U5814 (N_5814,N_4445,N_4081);
nor U5815 (N_5815,N_4575,N_4632);
xnor U5816 (N_5816,N_4317,N_4329);
xnor U5817 (N_5817,N_4557,N_4624);
or U5818 (N_5818,N_4023,N_4639);
or U5819 (N_5819,N_4811,N_4808);
and U5820 (N_5820,N_4574,N_4740);
nor U5821 (N_5821,N_4946,N_4391);
or U5822 (N_5822,N_4214,N_4376);
and U5823 (N_5823,N_4676,N_4695);
or U5824 (N_5824,N_4366,N_4024);
nor U5825 (N_5825,N_4755,N_4912);
nor U5826 (N_5826,N_4709,N_4184);
nor U5827 (N_5827,N_4021,N_4828);
nand U5828 (N_5828,N_4396,N_4380);
and U5829 (N_5829,N_4543,N_4839);
and U5830 (N_5830,N_4816,N_4227);
xor U5831 (N_5831,N_4969,N_4490);
or U5832 (N_5832,N_4458,N_4968);
xnor U5833 (N_5833,N_4270,N_4457);
and U5834 (N_5834,N_4002,N_4919);
or U5835 (N_5835,N_4218,N_4698);
xnor U5836 (N_5836,N_4023,N_4125);
or U5837 (N_5837,N_4735,N_4326);
nand U5838 (N_5838,N_4425,N_4191);
nand U5839 (N_5839,N_4433,N_4031);
nand U5840 (N_5840,N_4504,N_4775);
or U5841 (N_5841,N_4846,N_4531);
or U5842 (N_5842,N_4019,N_4006);
nand U5843 (N_5843,N_4131,N_4849);
nor U5844 (N_5844,N_4210,N_4347);
or U5845 (N_5845,N_4678,N_4745);
or U5846 (N_5846,N_4563,N_4273);
nor U5847 (N_5847,N_4980,N_4166);
nand U5848 (N_5848,N_4181,N_4987);
and U5849 (N_5849,N_4233,N_4029);
xor U5850 (N_5850,N_4435,N_4775);
nor U5851 (N_5851,N_4735,N_4538);
nor U5852 (N_5852,N_4665,N_4624);
xnor U5853 (N_5853,N_4553,N_4862);
and U5854 (N_5854,N_4936,N_4208);
or U5855 (N_5855,N_4156,N_4390);
nor U5856 (N_5856,N_4476,N_4955);
xor U5857 (N_5857,N_4189,N_4909);
nor U5858 (N_5858,N_4402,N_4275);
or U5859 (N_5859,N_4834,N_4930);
or U5860 (N_5860,N_4420,N_4078);
and U5861 (N_5861,N_4204,N_4782);
nand U5862 (N_5862,N_4121,N_4266);
xnor U5863 (N_5863,N_4836,N_4273);
nand U5864 (N_5864,N_4969,N_4537);
or U5865 (N_5865,N_4130,N_4212);
or U5866 (N_5866,N_4534,N_4811);
nand U5867 (N_5867,N_4878,N_4062);
nor U5868 (N_5868,N_4042,N_4553);
nand U5869 (N_5869,N_4004,N_4165);
nand U5870 (N_5870,N_4919,N_4607);
nor U5871 (N_5871,N_4065,N_4458);
xnor U5872 (N_5872,N_4726,N_4304);
nor U5873 (N_5873,N_4056,N_4167);
and U5874 (N_5874,N_4395,N_4804);
nor U5875 (N_5875,N_4908,N_4188);
nor U5876 (N_5876,N_4686,N_4357);
xor U5877 (N_5877,N_4442,N_4089);
xor U5878 (N_5878,N_4885,N_4954);
xnor U5879 (N_5879,N_4326,N_4819);
or U5880 (N_5880,N_4806,N_4868);
nor U5881 (N_5881,N_4376,N_4063);
nor U5882 (N_5882,N_4265,N_4650);
or U5883 (N_5883,N_4494,N_4993);
xor U5884 (N_5884,N_4181,N_4077);
xnor U5885 (N_5885,N_4367,N_4061);
nand U5886 (N_5886,N_4807,N_4841);
nor U5887 (N_5887,N_4167,N_4391);
nor U5888 (N_5888,N_4912,N_4594);
nor U5889 (N_5889,N_4219,N_4070);
xor U5890 (N_5890,N_4947,N_4150);
and U5891 (N_5891,N_4246,N_4921);
and U5892 (N_5892,N_4554,N_4169);
or U5893 (N_5893,N_4408,N_4011);
nor U5894 (N_5894,N_4000,N_4565);
or U5895 (N_5895,N_4684,N_4371);
and U5896 (N_5896,N_4639,N_4851);
or U5897 (N_5897,N_4633,N_4146);
and U5898 (N_5898,N_4971,N_4440);
nor U5899 (N_5899,N_4536,N_4688);
or U5900 (N_5900,N_4299,N_4673);
nor U5901 (N_5901,N_4931,N_4231);
nand U5902 (N_5902,N_4120,N_4018);
and U5903 (N_5903,N_4483,N_4715);
and U5904 (N_5904,N_4972,N_4863);
and U5905 (N_5905,N_4964,N_4539);
xnor U5906 (N_5906,N_4102,N_4891);
or U5907 (N_5907,N_4681,N_4205);
xor U5908 (N_5908,N_4210,N_4647);
and U5909 (N_5909,N_4954,N_4173);
and U5910 (N_5910,N_4733,N_4986);
and U5911 (N_5911,N_4070,N_4501);
nand U5912 (N_5912,N_4054,N_4144);
xnor U5913 (N_5913,N_4873,N_4535);
or U5914 (N_5914,N_4744,N_4858);
nor U5915 (N_5915,N_4151,N_4623);
xor U5916 (N_5916,N_4907,N_4363);
nor U5917 (N_5917,N_4404,N_4312);
xor U5918 (N_5918,N_4085,N_4532);
nand U5919 (N_5919,N_4490,N_4714);
xnor U5920 (N_5920,N_4469,N_4506);
nand U5921 (N_5921,N_4898,N_4582);
nor U5922 (N_5922,N_4105,N_4102);
nor U5923 (N_5923,N_4170,N_4055);
nand U5924 (N_5924,N_4443,N_4199);
or U5925 (N_5925,N_4895,N_4208);
xnor U5926 (N_5926,N_4973,N_4430);
or U5927 (N_5927,N_4920,N_4617);
nand U5928 (N_5928,N_4854,N_4669);
or U5929 (N_5929,N_4212,N_4302);
nor U5930 (N_5930,N_4415,N_4891);
nor U5931 (N_5931,N_4154,N_4936);
or U5932 (N_5932,N_4173,N_4181);
nor U5933 (N_5933,N_4511,N_4619);
nor U5934 (N_5934,N_4478,N_4766);
or U5935 (N_5935,N_4841,N_4394);
nand U5936 (N_5936,N_4556,N_4523);
nor U5937 (N_5937,N_4878,N_4747);
nand U5938 (N_5938,N_4948,N_4150);
and U5939 (N_5939,N_4420,N_4639);
and U5940 (N_5940,N_4168,N_4579);
and U5941 (N_5941,N_4660,N_4111);
and U5942 (N_5942,N_4035,N_4445);
nand U5943 (N_5943,N_4408,N_4417);
xnor U5944 (N_5944,N_4487,N_4898);
and U5945 (N_5945,N_4168,N_4167);
or U5946 (N_5946,N_4195,N_4539);
xnor U5947 (N_5947,N_4060,N_4569);
xnor U5948 (N_5948,N_4268,N_4188);
or U5949 (N_5949,N_4506,N_4682);
and U5950 (N_5950,N_4251,N_4493);
nor U5951 (N_5951,N_4245,N_4328);
or U5952 (N_5952,N_4336,N_4131);
and U5953 (N_5953,N_4062,N_4858);
and U5954 (N_5954,N_4682,N_4288);
or U5955 (N_5955,N_4866,N_4776);
or U5956 (N_5956,N_4054,N_4058);
or U5957 (N_5957,N_4307,N_4519);
xor U5958 (N_5958,N_4291,N_4457);
xor U5959 (N_5959,N_4407,N_4002);
or U5960 (N_5960,N_4263,N_4607);
nand U5961 (N_5961,N_4331,N_4600);
or U5962 (N_5962,N_4349,N_4127);
xor U5963 (N_5963,N_4170,N_4686);
nand U5964 (N_5964,N_4287,N_4435);
nor U5965 (N_5965,N_4431,N_4856);
nor U5966 (N_5966,N_4806,N_4640);
nor U5967 (N_5967,N_4472,N_4794);
nor U5968 (N_5968,N_4249,N_4326);
nand U5969 (N_5969,N_4361,N_4838);
nand U5970 (N_5970,N_4198,N_4597);
and U5971 (N_5971,N_4446,N_4498);
or U5972 (N_5972,N_4339,N_4904);
nand U5973 (N_5973,N_4826,N_4200);
nor U5974 (N_5974,N_4361,N_4060);
or U5975 (N_5975,N_4739,N_4837);
xor U5976 (N_5976,N_4089,N_4520);
nor U5977 (N_5977,N_4701,N_4896);
or U5978 (N_5978,N_4233,N_4644);
nand U5979 (N_5979,N_4063,N_4638);
xnor U5980 (N_5980,N_4673,N_4588);
or U5981 (N_5981,N_4838,N_4009);
nand U5982 (N_5982,N_4711,N_4760);
or U5983 (N_5983,N_4307,N_4974);
nor U5984 (N_5984,N_4574,N_4910);
nand U5985 (N_5985,N_4674,N_4817);
nor U5986 (N_5986,N_4534,N_4069);
nand U5987 (N_5987,N_4716,N_4050);
xor U5988 (N_5988,N_4916,N_4103);
nor U5989 (N_5989,N_4376,N_4940);
nor U5990 (N_5990,N_4260,N_4629);
xnor U5991 (N_5991,N_4316,N_4955);
nand U5992 (N_5992,N_4455,N_4580);
nor U5993 (N_5993,N_4807,N_4443);
or U5994 (N_5994,N_4439,N_4702);
xnor U5995 (N_5995,N_4134,N_4303);
and U5996 (N_5996,N_4881,N_4571);
nand U5997 (N_5997,N_4493,N_4955);
or U5998 (N_5998,N_4793,N_4081);
nand U5999 (N_5999,N_4108,N_4164);
nor U6000 (N_6000,N_5752,N_5136);
nor U6001 (N_6001,N_5268,N_5109);
nor U6002 (N_6002,N_5923,N_5809);
nand U6003 (N_6003,N_5726,N_5714);
xor U6004 (N_6004,N_5771,N_5783);
xor U6005 (N_6005,N_5501,N_5585);
and U6006 (N_6006,N_5756,N_5139);
xor U6007 (N_6007,N_5987,N_5527);
nand U6008 (N_6008,N_5369,N_5272);
and U6009 (N_6009,N_5006,N_5488);
or U6010 (N_6010,N_5031,N_5759);
or U6011 (N_6011,N_5789,N_5490);
or U6012 (N_6012,N_5038,N_5449);
nor U6013 (N_6013,N_5371,N_5480);
and U6014 (N_6014,N_5803,N_5266);
or U6015 (N_6015,N_5703,N_5248);
nor U6016 (N_6016,N_5012,N_5039);
nor U6017 (N_6017,N_5652,N_5740);
nand U6018 (N_6018,N_5440,N_5320);
nand U6019 (N_6019,N_5225,N_5680);
nand U6020 (N_6020,N_5066,N_5681);
nand U6021 (N_6021,N_5676,N_5938);
nand U6022 (N_6022,N_5285,N_5532);
nor U6023 (N_6023,N_5370,N_5707);
nor U6024 (N_6024,N_5884,N_5297);
xor U6025 (N_6025,N_5090,N_5725);
nand U6026 (N_6026,N_5723,N_5454);
or U6027 (N_6027,N_5858,N_5169);
nand U6028 (N_6028,N_5633,N_5436);
xor U6029 (N_6029,N_5889,N_5439);
or U6030 (N_6030,N_5104,N_5607);
xnor U6031 (N_6031,N_5750,N_5015);
or U6032 (N_6032,N_5940,N_5893);
xor U6033 (N_6033,N_5985,N_5002);
or U6034 (N_6034,N_5388,N_5409);
or U6035 (N_6035,N_5042,N_5170);
xnor U6036 (N_6036,N_5308,N_5534);
or U6037 (N_6037,N_5686,N_5850);
or U6038 (N_6038,N_5129,N_5928);
nand U6039 (N_6039,N_5566,N_5905);
and U6040 (N_6040,N_5577,N_5797);
or U6041 (N_6041,N_5291,N_5852);
and U6042 (N_6042,N_5559,N_5970);
nor U6043 (N_6043,N_5616,N_5205);
nand U6044 (N_6044,N_5380,N_5262);
nor U6045 (N_6045,N_5653,N_5084);
and U6046 (N_6046,N_5802,N_5043);
nand U6047 (N_6047,N_5727,N_5739);
xor U6048 (N_6048,N_5922,N_5080);
xor U6049 (N_6049,N_5337,N_5619);
xor U6050 (N_6050,N_5103,N_5896);
and U6051 (N_6051,N_5310,N_5267);
nor U6052 (N_6052,N_5142,N_5845);
or U6053 (N_6053,N_5419,N_5798);
nand U6054 (N_6054,N_5097,N_5368);
and U6055 (N_6055,N_5351,N_5235);
xnor U6056 (N_6056,N_5751,N_5432);
nand U6057 (N_6057,N_5975,N_5834);
or U6058 (N_6058,N_5383,N_5018);
nor U6059 (N_6059,N_5426,N_5515);
nand U6060 (N_6060,N_5886,N_5996);
and U6061 (N_6061,N_5269,N_5067);
nor U6062 (N_6062,N_5167,N_5332);
nor U6063 (N_6063,N_5499,N_5019);
nor U6064 (N_6064,N_5322,N_5247);
and U6065 (N_6065,N_5945,N_5780);
or U6066 (N_6066,N_5132,N_5154);
nor U6067 (N_6067,N_5529,N_5004);
xnor U6068 (N_6068,N_5563,N_5784);
xor U6069 (N_6069,N_5448,N_5656);
xor U6070 (N_6070,N_5230,N_5222);
or U6071 (N_6071,N_5513,N_5500);
xnor U6072 (N_6072,N_5251,N_5962);
or U6073 (N_6073,N_5863,N_5821);
xor U6074 (N_6074,N_5149,N_5530);
or U6075 (N_6075,N_5462,N_5484);
xor U6076 (N_6076,N_5979,N_5531);
nor U6077 (N_6077,N_5143,N_5433);
and U6078 (N_6078,N_5977,N_5904);
nand U6079 (N_6079,N_5754,N_5564);
xor U6080 (N_6080,N_5976,N_5869);
or U6081 (N_6081,N_5441,N_5762);
nand U6082 (N_6082,N_5549,N_5278);
nand U6083 (N_6083,N_5284,N_5711);
xor U6084 (N_6084,N_5952,N_5187);
nor U6085 (N_6085,N_5698,N_5325);
and U6086 (N_6086,N_5258,N_5941);
and U6087 (N_6087,N_5650,N_5181);
or U6088 (N_6088,N_5437,N_5227);
xor U6089 (N_6089,N_5662,N_5110);
nor U6090 (N_6090,N_5746,N_5315);
xnor U6091 (N_6091,N_5827,N_5483);
nor U6092 (N_6092,N_5024,N_5197);
nand U6093 (N_6093,N_5156,N_5603);
and U6094 (N_6094,N_5548,N_5728);
xnor U6095 (N_6095,N_5620,N_5636);
xor U6096 (N_6096,N_5206,N_5316);
and U6097 (N_6097,N_5423,N_5157);
and U6098 (N_6098,N_5737,N_5891);
nand U6099 (N_6099,N_5849,N_5554);
nor U6100 (N_6100,N_5243,N_5874);
nand U6101 (N_6101,N_5425,N_5776);
nand U6102 (N_6102,N_5763,N_5062);
nand U6103 (N_6103,N_5856,N_5647);
nand U6104 (N_6104,N_5398,N_5733);
xor U6105 (N_6105,N_5931,N_5822);
and U6106 (N_6106,N_5175,N_5796);
and U6107 (N_6107,N_5379,N_5870);
and U6108 (N_6108,N_5343,N_5161);
xnor U6109 (N_6109,N_5048,N_5086);
xor U6110 (N_6110,N_5010,N_5866);
nor U6111 (N_6111,N_5583,N_5516);
and U6112 (N_6112,N_5994,N_5663);
and U6113 (N_6113,N_5775,N_5117);
xnor U6114 (N_6114,N_5805,N_5178);
and U6115 (N_6115,N_5311,N_5667);
xor U6116 (N_6116,N_5831,N_5787);
xor U6117 (N_6117,N_5344,N_5966);
nand U6118 (N_6118,N_5690,N_5326);
xor U6119 (N_6119,N_5608,N_5151);
nand U6120 (N_6120,N_5214,N_5670);
or U6121 (N_6121,N_5778,N_5936);
nand U6122 (N_6122,N_5918,N_5921);
nor U6123 (N_6123,N_5446,N_5742);
nand U6124 (N_6124,N_5618,N_5535);
nor U6125 (N_6125,N_5735,N_5150);
or U6126 (N_6126,N_5321,N_5826);
or U6127 (N_6127,N_5333,N_5438);
and U6128 (N_6128,N_5832,N_5494);
or U6129 (N_6129,N_5871,N_5260);
nand U6130 (N_6130,N_5777,N_5068);
or U6131 (N_6131,N_5592,N_5328);
or U6132 (N_6132,N_5173,N_5298);
xnor U6133 (N_6133,N_5242,N_5948);
or U6134 (N_6134,N_5729,N_5466);
nand U6135 (N_6135,N_5875,N_5696);
nor U6136 (N_6136,N_5479,N_5894);
nand U6137 (N_6137,N_5610,N_5883);
nor U6138 (N_6138,N_5401,N_5281);
xor U6139 (N_6139,N_5482,N_5359);
or U6140 (N_6140,N_5906,N_5949);
nor U6141 (N_6141,N_5393,N_5946);
xnor U6142 (N_6142,N_5558,N_5145);
nand U6143 (N_6143,N_5634,N_5828);
nor U6144 (N_6144,N_5163,N_5572);
or U6145 (N_6145,N_5353,N_5836);
xnor U6146 (N_6146,N_5933,N_5541);
nor U6147 (N_6147,N_5410,N_5288);
or U6148 (N_6148,N_5624,N_5890);
nor U6149 (N_6149,N_5003,N_5571);
nand U6150 (N_6150,N_5715,N_5271);
nand U6151 (N_6151,N_5747,N_5105);
nand U6152 (N_6152,N_5580,N_5102);
or U6153 (N_6153,N_5615,N_5493);
nor U6154 (N_6154,N_5509,N_5280);
xnor U6155 (N_6155,N_5233,N_5396);
or U6156 (N_6156,N_5293,N_5005);
nand U6157 (N_6157,N_5518,N_5342);
xor U6158 (N_6158,N_5391,N_5605);
nand U6159 (N_6159,N_5362,N_5492);
or U6160 (N_6160,N_5338,N_5144);
xor U6161 (N_6161,N_5877,N_5191);
nor U6162 (N_6162,N_5304,N_5035);
nor U6163 (N_6163,N_5357,N_5567);
or U6164 (N_6164,N_5460,N_5404);
nor U6165 (N_6165,N_5000,N_5033);
nand U6166 (N_6166,N_5372,N_5443);
or U6167 (N_6167,N_5963,N_5622);
xnor U6168 (N_6168,N_5220,N_5470);
nand U6169 (N_6169,N_5349,N_5734);
nand U6170 (N_6170,N_5758,N_5261);
nor U6171 (N_6171,N_5160,N_5244);
xor U6172 (N_6172,N_5793,N_5504);
or U6173 (N_6173,N_5761,N_5327);
xor U6174 (N_6174,N_5617,N_5137);
or U6175 (N_6175,N_5825,N_5407);
nor U6176 (N_6176,N_5376,N_5378);
and U6177 (N_6177,N_5782,N_5553);
or U6178 (N_6178,N_5234,N_5275);
or U6179 (N_6179,N_5700,N_5017);
and U6180 (N_6180,N_5444,N_5898);
nor U6181 (N_6181,N_5960,N_5324);
nor U6182 (N_6182,N_5971,N_5190);
xnor U6183 (N_6183,N_5279,N_5168);
and U6184 (N_6184,N_5375,N_5427);
and U6185 (N_6185,N_5697,N_5318);
nor U6186 (N_6186,N_5679,N_5844);
nand U6187 (N_6187,N_5645,N_5286);
nor U6188 (N_6188,N_5568,N_5202);
nor U6189 (N_6189,N_5228,N_5910);
nor U6190 (N_6190,N_5596,N_5467);
xnor U6191 (N_6191,N_5064,N_5442);
and U6192 (N_6192,N_5589,N_5087);
and U6193 (N_6193,N_5245,N_5118);
and U6194 (N_6194,N_5702,N_5902);
nor U6195 (N_6195,N_5341,N_5126);
xor U6196 (N_6196,N_5853,N_5599);
or U6197 (N_6197,N_5111,N_5346);
nand U6198 (N_6198,N_5195,N_5766);
nor U6199 (N_6199,N_5112,N_5508);
nor U6200 (N_6200,N_5699,N_5788);
xnor U6201 (N_6201,N_5146,N_5299);
or U6202 (N_6202,N_5988,N_5287);
nor U6203 (N_6203,N_5289,N_5100);
nand U6204 (N_6204,N_5037,N_5053);
xor U6205 (N_6205,N_5842,N_5709);
and U6206 (N_6206,N_5528,N_5431);
or U6207 (N_6207,N_5034,N_5198);
xnor U6208 (N_6208,N_5974,N_5843);
and U6209 (N_6209,N_5485,N_5913);
or U6210 (N_6210,N_5473,N_5632);
nor U6211 (N_6211,N_5331,N_5623);
nand U6212 (N_6212,N_5795,N_5303);
and U6213 (N_6213,N_5395,N_5521);
xor U6214 (N_6214,N_5744,N_5141);
and U6215 (N_6215,N_5965,N_5808);
nor U6216 (N_6216,N_5107,N_5045);
nor U6217 (N_6217,N_5159,N_5629);
or U6218 (N_6218,N_5989,N_5174);
and U6219 (N_6219,N_5040,N_5718);
nor U6220 (N_6220,N_5550,N_5429);
and U6221 (N_6221,N_5791,N_5123);
xnor U6222 (N_6222,N_5131,N_5212);
nor U6223 (N_6223,N_5800,N_5957);
or U6224 (N_6224,N_5408,N_5022);
xnor U6225 (N_6225,N_5319,N_5188);
and U6226 (N_6226,N_5811,N_5323);
xnor U6227 (N_6227,N_5124,N_5211);
nor U6228 (N_6228,N_5475,N_5172);
nor U6229 (N_6229,N_5049,N_5955);
xnor U6230 (N_6230,N_5867,N_5745);
xnor U6231 (N_6231,N_5030,N_5959);
nand U6232 (N_6232,N_5611,N_5706);
nor U6233 (N_6233,N_5929,N_5785);
xor U6234 (N_6234,N_5179,N_5011);
nor U6235 (N_6235,N_5070,N_5678);
nor U6236 (N_6236,N_5660,N_5336);
and U6237 (N_6237,N_5073,N_5602);
nand U6238 (N_6238,N_5095,N_5916);
and U6239 (N_6239,N_5468,N_5519);
nor U6240 (N_6240,N_5542,N_5586);
xnor U6241 (N_6241,N_5947,N_5226);
nand U6242 (N_6242,N_5912,N_5593);
nand U6243 (N_6243,N_5236,N_5063);
xnor U6244 (N_6244,N_5814,N_5083);
nand U6245 (N_6245,N_5522,N_5738);
nand U6246 (N_6246,N_5972,N_5694);
nor U6247 (N_6247,N_5847,N_5184);
or U6248 (N_6248,N_5390,N_5356);
and U6249 (N_6249,N_5930,N_5330);
xor U6250 (N_6250,N_5786,N_5773);
nand U6251 (N_6251,N_5223,N_5790);
xor U6252 (N_6252,N_5807,N_5524);
and U6253 (N_6253,N_5021,N_5654);
nand U6254 (N_6254,N_5186,N_5920);
nand U6255 (N_6255,N_5249,N_5743);
nand U6256 (N_6256,N_5465,N_5254);
xor U6257 (N_6257,N_5628,N_5876);
or U6258 (N_6258,N_5007,N_5273);
nor U6259 (N_6259,N_5968,N_5630);
xnor U6260 (N_6260,N_5329,N_5525);
nand U6261 (N_6261,N_5116,N_5882);
or U6262 (N_6262,N_5093,N_5969);
or U6263 (N_6263,N_5666,N_5301);
nor U6264 (N_6264,N_5153,N_5639);
nand U6265 (N_6265,N_5020,N_5682);
nor U6266 (N_6266,N_5907,N_5428);
nor U6267 (N_6267,N_5052,N_5373);
and U6268 (N_6268,N_5259,N_5282);
nor U6269 (N_6269,N_5794,N_5792);
nand U6270 (N_6270,N_5387,N_5246);
and U6271 (N_6271,N_5270,N_5025);
or U6272 (N_6272,N_5489,N_5865);
nand U6273 (N_6273,N_5481,N_5935);
nor U6274 (N_6274,N_5685,N_5908);
or U6275 (N_6275,N_5594,N_5609);
xnor U6276 (N_6276,N_5354,N_5815);
and U6277 (N_6277,N_5673,N_5998);
nand U6278 (N_6278,N_5452,N_5027);
nor U6279 (N_6279,N_5665,N_5964);
nor U6280 (N_6280,N_5241,N_5731);
nand U6281 (N_6281,N_5981,N_5218);
and U6282 (N_6282,N_5309,N_5445);
xor U6283 (N_6283,N_5637,N_5641);
xnor U6284 (N_6284,N_5956,N_5047);
nand U6285 (N_6285,N_5833,N_5999);
nor U6286 (N_6286,N_5755,N_5512);
and U6287 (N_6287,N_5416,N_5290);
nand U6288 (N_6288,N_5879,N_5418);
xnor U6289 (N_6289,N_5505,N_5415);
and U6290 (N_6290,N_5810,N_5597);
nor U6291 (N_6291,N_5413,N_5355);
nand U6292 (N_6292,N_5732,N_5455);
or U6293 (N_6293,N_5127,N_5135);
nor U6294 (N_6294,N_5712,N_5887);
nor U6295 (N_6295,N_5061,N_5403);
nor U6296 (N_6296,N_5098,N_5717);
xnor U6297 (N_6297,N_5201,N_5082);
nand U6298 (N_6298,N_5768,N_5899);
nand U6299 (N_6299,N_5240,N_5672);
or U6300 (N_6300,N_5925,N_5453);
nand U6301 (N_6301,N_5598,N_5683);
and U6302 (N_6302,N_5540,N_5350);
and U6303 (N_6303,N_5892,N_5231);
and U6304 (N_6304,N_5417,N_5026);
or U6305 (N_6305,N_5292,N_5400);
nor U6306 (N_6306,N_5182,N_5753);
and U6307 (N_6307,N_5399,N_5526);
nor U6308 (N_6308,N_5757,N_5995);
and U6309 (N_6309,N_5074,N_5180);
and U6310 (N_6310,N_5250,N_5069);
xnor U6311 (N_6311,N_5644,N_5997);
nand U6312 (N_6312,N_5177,N_5199);
or U6313 (N_6313,N_5217,N_5502);
nand U6314 (N_6314,N_5691,N_5461);
xnor U6315 (N_6315,N_5614,N_5774);
nor U6316 (N_6316,N_5885,N_5591);
and U6317 (N_6317,N_5770,N_5089);
or U6318 (N_6318,N_5265,N_5424);
nand U6319 (N_6319,N_5878,N_5340);
and U6320 (N_6320,N_5171,N_5381);
xor U6321 (N_6321,N_5943,N_5576);
xnor U6322 (N_6322,N_5911,N_5895);
and U6323 (N_6323,N_5352,N_5560);
nand U6324 (N_6324,N_5434,N_5239);
nor U6325 (N_6325,N_5059,N_5613);
and U6326 (N_6326,N_5451,N_5919);
xor U6327 (N_6327,N_5651,N_5295);
or U6328 (N_6328,N_5219,N_5119);
nand U6329 (N_6329,N_5978,N_5075);
and U6330 (N_6330,N_5961,N_5347);
nor U6331 (N_6331,N_5713,N_5307);
xor U6332 (N_6332,N_5386,N_5057);
nand U6333 (N_6333,N_5009,N_5973);
nand U6334 (N_6334,N_5574,N_5868);
nand U6335 (N_6335,N_5716,N_5194);
xor U6336 (N_6336,N_5649,N_5993);
xor U6337 (N_6337,N_5846,N_5088);
xor U6338 (N_6338,N_5224,N_5054);
or U6339 (N_6339,N_5538,N_5058);
xnor U6340 (N_6340,N_5575,N_5498);
and U6341 (N_6341,N_5779,N_5873);
and U6342 (N_6342,N_5569,N_5950);
or U6343 (N_6343,N_5101,N_5909);
nor U6344 (N_6344,N_5096,N_5203);
nand U6345 (N_6345,N_5207,N_5402);
or U6346 (N_6346,N_5365,N_5487);
and U6347 (N_6347,N_5345,N_5570);
xnor U6348 (N_6348,N_5183,N_5937);
and U6349 (N_6349,N_5176,N_5990);
nand U6350 (N_6350,N_5506,N_5300);
nor U6351 (N_6351,N_5412,N_5196);
nand U6352 (N_6352,N_5621,N_5823);
xnor U6353 (N_6353,N_5561,N_5927);
and U6354 (N_6354,N_5028,N_5704);
nor U6355 (N_6355,N_5824,N_5626);
nand U6356 (N_6356,N_5276,N_5544);
nor U6357 (N_6357,N_5189,N_5769);
xor U6358 (N_6358,N_5001,N_5121);
nand U6359 (N_6359,N_5719,N_5692);
or U6360 (N_6360,N_5851,N_5363);
nand U6361 (N_6361,N_5926,N_5819);
and U6362 (N_6362,N_5274,N_5263);
xor U6363 (N_6363,N_5335,N_5838);
nand U6364 (N_6364,N_5491,N_5748);
xor U6365 (N_6365,N_5812,N_5152);
nor U6366 (N_6366,N_5646,N_5032);
nand U6367 (N_6367,N_5511,N_5749);
nor U6368 (N_6368,N_5317,N_5606);
nand U6369 (N_6369,N_5830,N_5953);
and U6370 (N_6370,N_5642,N_5185);
nand U6371 (N_6371,N_5625,N_5060);
and U6372 (N_6372,N_5817,N_5801);
xnor U6373 (N_6373,N_5669,N_5765);
nand U6374 (N_6374,N_5557,N_5469);
nand U6375 (N_6375,N_5724,N_5684);
nand U6376 (N_6376,N_5474,N_5587);
xor U6377 (N_6377,N_5208,N_5533);
xor U6378 (N_6378,N_5255,N_5507);
and U6379 (N_6379,N_5983,N_5166);
or U6380 (N_6380,N_5115,N_5215);
nor U6381 (N_6381,N_5108,N_5939);
nand U6382 (N_6382,N_5164,N_5361);
nand U6383 (N_6383,N_5671,N_5781);
and U6384 (N_6384,N_5552,N_5901);
xor U6385 (N_6385,N_5991,N_5495);
xor U6386 (N_6386,N_5539,N_5471);
and U6387 (N_6387,N_5982,N_5076);
xnor U6388 (N_6388,N_5209,N_5503);
xnor U6389 (N_6389,N_5612,N_5720);
or U6390 (N_6390,N_5253,N_5463);
xor U6391 (N_6391,N_5496,N_5394);
nor U6392 (N_6392,N_5458,N_5600);
or U6393 (N_6393,N_5165,N_5545);
or U6394 (N_6394,N_5556,N_5221);
nand U6395 (N_6395,N_5459,N_5595);
or U6396 (N_6396,N_5133,N_5008);
nand U6397 (N_6397,N_5079,N_5421);
nand U6398 (N_6398,N_5536,N_5829);
nand U6399 (N_6399,N_5581,N_5857);
nand U6400 (N_6400,N_5954,N_5120);
and U6401 (N_6401,N_5200,N_5520);
nand U6402 (N_6402,N_5476,N_5050);
nand U6403 (N_6403,N_5277,N_5130);
or U6404 (N_6404,N_5640,N_5114);
xor U6405 (N_6405,N_5693,N_5162);
nor U6406 (N_6406,N_5687,N_5364);
and U6407 (N_6407,N_5138,N_5296);
and U6408 (N_6408,N_5314,N_5113);
nor U6409 (N_6409,N_5367,N_5377);
or U6410 (N_6410,N_5430,N_5457);
nor U6411 (N_6411,N_5204,N_5701);
nand U6412 (N_6412,N_5565,N_5730);
or U6413 (N_6413,N_5590,N_5635);
xor U6414 (N_6414,N_5839,N_5841);
nand U6415 (N_6415,N_5767,N_5992);
and U6416 (N_6416,N_5213,N_5689);
and U6417 (N_6417,N_5880,N_5664);
xor U6418 (N_6418,N_5543,N_5252);
and U6419 (N_6419,N_5631,N_5721);
xnor U6420 (N_6420,N_5478,N_5806);
nor U6421 (N_6421,N_5951,N_5804);
nor U6422 (N_6422,N_5081,N_5555);
and U6423 (N_6423,N_5405,N_5125);
nand U6424 (N_6424,N_5422,N_5710);
or U6425 (N_6425,N_5435,N_5897);
nand U6426 (N_6426,N_5818,N_5257);
or U6427 (N_6427,N_5385,N_5638);
nand U6428 (N_6428,N_5914,N_5588);
or U6429 (N_6429,N_5967,N_5094);
and U6430 (N_6430,N_5382,N_5643);
xnor U6431 (N_6431,N_5464,N_5934);
xor U6432 (N_6432,N_5456,N_5772);
nand U6433 (N_6433,N_5741,N_5551);
and U6434 (N_6434,N_5389,N_5514);
or U6435 (N_6435,N_5216,N_5888);
nor U6436 (N_6436,N_5392,N_5799);
xnor U6437 (N_6437,N_5044,N_5374);
nor U6438 (N_6438,N_5859,N_5736);
and U6439 (N_6439,N_5722,N_5562);
and U6440 (N_6440,N_5764,N_5036);
xor U6441 (N_6441,N_5579,N_5046);
or U6442 (N_6442,N_5312,N_5155);
and U6443 (N_6443,N_5237,N_5283);
nor U6444 (N_6444,N_5041,N_5232);
nand U6445 (N_6445,N_5128,N_5302);
nor U6446 (N_6446,N_5547,N_5148);
nor U6447 (N_6447,N_5029,N_5980);
nand U6448 (N_6448,N_5659,N_5305);
or U6449 (N_6449,N_5537,N_5106);
nand U6450 (N_6450,N_5816,N_5192);
and U6451 (N_6451,N_5134,N_5861);
xnor U6452 (N_6452,N_5140,N_5472);
nor U6453 (N_6453,N_5091,N_5486);
nor U6454 (N_6454,N_5414,N_5864);
and U6455 (N_6455,N_5013,N_5099);
nor U6456 (N_6456,N_5210,N_5658);
and U6457 (N_6457,N_5334,N_5674);
nor U6458 (N_6458,N_5820,N_5601);
nand U6459 (N_6459,N_5051,N_5411);
or U6460 (N_6460,N_5397,N_5056);
xnor U6461 (N_6461,N_5450,N_5627);
xor U6462 (N_6462,N_5984,N_5313);
xor U6463 (N_6463,N_5604,N_5675);
and U6464 (N_6464,N_5688,N_5147);
and U6465 (N_6465,N_5077,N_5497);
nand U6466 (N_6466,N_5055,N_5855);
xnor U6467 (N_6467,N_5306,N_5092);
and U6468 (N_6468,N_5915,N_5578);
xnor U6469 (N_6469,N_5986,N_5708);
xor U6470 (N_6470,N_5813,N_5229);
or U6471 (N_6471,N_5193,N_5510);
and U6472 (N_6472,N_5677,N_5860);
nand U6473 (N_6473,N_5264,N_5573);
xnor U6474 (N_6474,N_5942,N_5085);
nor U6475 (N_6475,N_5072,N_5023);
nor U6476 (N_6476,N_5705,N_5661);
or U6477 (N_6477,N_5238,N_5014);
and U6478 (N_6478,N_5760,N_5881);
or U6479 (N_6479,N_5523,N_5584);
xor U6480 (N_6480,N_5840,N_5655);
or U6481 (N_6481,N_5872,N_5294);
nand U6482 (N_6482,N_5420,N_5358);
or U6483 (N_6483,N_5348,N_5944);
nor U6484 (N_6484,N_5657,N_5835);
and U6485 (N_6485,N_5668,N_5071);
nand U6486 (N_6486,N_5903,N_5065);
xnor U6487 (N_6487,N_5360,N_5862);
or U6488 (N_6488,N_5848,N_5517);
xor U6489 (N_6489,N_5447,N_5477);
or U6490 (N_6490,N_5854,N_5924);
nor U6491 (N_6491,N_5648,N_5016);
xor U6492 (N_6492,N_5837,N_5900);
xor U6493 (N_6493,N_5932,N_5958);
or U6494 (N_6494,N_5582,N_5078);
and U6495 (N_6495,N_5384,N_5406);
xor U6496 (N_6496,N_5256,N_5158);
nor U6497 (N_6497,N_5546,N_5366);
xor U6498 (N_6498,N_5122,N_5695);
xor U6499 (N_6499,N_5339,N_5917);
nand U6500 (N_6500,N_5205,N_5374);
nor U6501 (N_6501,N_5830,N_5053);
nand U6502 (N_6502,N_5763,N_5991);
or U6503 (N_6503,N_5766,N_5417);
nor U6504 (N_6504,N_5808,N_5212);
nor U6505 (N_6505,N_5318,N_5484);
or U6506 (N_6506,N_5521,N_5072);
or U6507 (N_6507,N_5641,N_5211);
or U6508 (N_6508,N_5998,N_5613);
and U6509 (N_6509,N_5924,N_5071);
xor U6510 (N_6510,N_5336,N_5328);
nor U6511 (N_6511,N_5803,N_5407);
or U6512 (N_6512,N_5103,N_5546);
nor U6513 (N_6513,N_5445,N_5580);
xor U6514 (N_6514,N_5631,N_5193);
xor U6515 (N_6515,N_5608,N_5000);
and U6516 (N_6516,N_5515,N_5577);
nor U6517 (N_6517,N_5356,N_5975);
nand U6518 (N_6518,N_5156,N_5041);
and U6519 (N_6519,N_5616,N_5489);
nor U6520 (N_6520,N_5931,N_5852);
nand U6521 (N_6521,N_5077,N_5661);
or U6522 (N_6522,N_5628,N_5663);
nand U6523 (N_6523,N_5353,N_5310);
nand U6524 (N_6524,N_5723,N_5852);
xnor U6525 (N_6525,N_5188,N_5562);
and U6526 (N_6526,N_5621,N_5203);
nor U6527 (N_6527,N_5943,N_5363);
or U6528 (N_6528,N_5757,N_5693);
nand U6529 (N_6529,N_5325,N_5877);
and U6530 (N_6530,N_5787,N_5465);
nand U6531 (N_6531,N_5687,N_5209);
nand U6532 (N_6532,N_5121,N_5612);
nor U6533 (N_6533,N_5506,N_5129);
or U6534 (N_6534,N_5071,N_5934);
or U6535 (N_6535,N_5957,N_5783);
xnor U6536 (N_6536,N_5274,N_5835);
nor U6537 (N_6537,N_5288,N_5201);
or U6538 (N_6538,N_5229,N_5278);
nor U6539 (N_6539,N_5110,N_5523);
and U6540 (N_6540,N_5716,N_5407);
xnor U6541 (N_6541,N_5085,N_5806);
and U6542 (N_6542,N_5105,N_5704);
nor U6543 (N_6543,N_5648,N_5735);
or U6544 (N_6544,N_5620,N_5305);
and U6545 (N_6545,N_5118,N_5040);
nand U6546 (N_6546,N_5563,N_5011);
nor U6547 (N_6547,N_5383,N_5750);
or U6548 (N_6548,N_5886,N_5554);
or U6549 (N_6549,N_5014,N_5108);
xor U6550 (N_6550,N_5944,N_5569);
nand U6551 (N_6551,N_5226,N_5705);
and U6552 (N_6552,N_5298,N_5382);
nor U6553 (N_6553,N_5064,N_5353);
nor U6554 (N_6554,N_5131,N_5016);
nor U6555 (N_6555,N_5313,N_5816);
nor U6556 (N_6556,N_5754,N_5166);
or U6557 (N_6557,N_5800,N_5817);
and U6558 (N_6558,N_5167,N_5590);
or U6559 (N_6559,N_5708,N_5226);
or U6560 (N_6560,N_5964,N_5308);
nor U6561 (N_6561,N_5518,N_5227);
xor U6562 (N_6562,N_5855,N_5465);
or U6563 (N_6563,N_5466,N_5923);
nor U6564 (N_6564,N_5660,N_5665);
xor U6565 (N_6565,N_5228,N_5386);
or U6566 (N_6566,N_5866,N_5667);
nor U6567 (N_6567,N_5278,N_5699);
nor U6568 (N_6568,N_5146,N_5282);
xor U6569 (N_6569,N_5789,N_5922);
or U6570 (N_6570,N_5962,N_5368);
nand U6571 (N_6571,N_5356,N_5308);
or U6572 (N_6572,N_5152,N_5034);
xnor U6573 (N_6573,N_5467,N_5339);
nand U6574 (N_6574,N_5029,N_5933);
nand U6575 (N_6575,N_5299,N_5976);
xnor U6576 (N_6576,N_5213,N_5628);
and U6577 (N_6577,N_5072,N_5071);
nand U6578 (N_6578,N_5216,N_5785);
and U6579 (N_6579,N_5416,N_5984);
and U6580 (N_6580,N_5013,N_5737);
xnor U6581 (N_6581,N_5855,N_5462);
and U6582 (N_6582,N_5684,N_5763);
xor U6583 (N_6583,N_5936,N_5570);
xor U6584 (N_6584,N_5884,N_5281);
xnor U6585 (N_6585,N_5786,N_5249);
nor U6586 (N_6586,N_5846,N_5622);
nand U6587 (N_6587,N_5232,N_5356);
nor U6588 (N_6588,N_5869,N_5310);
nor U6589 (N_6589,N_5994,N_5869);
or U6590 (N_6590,N_5515,N_5429);
nand U6591 (N_6591,N_5501,N_5238);
nor U6592 (N_6592,N_5828,N_5324);
xor U6593 (N_6593,N_5182,N_5250);
nor U6594 (N_6594,N_5765,N_5857);
nor U6595 (N_6595,N_5575,N_5714);
and U6596 (N_6596,N_5463,N_5064);
nor U6597 (N_6597,N_5548,N_5070);
and U6598 (N_6598,N_5438,N_5686);
xor U6599 (N_6599,N_5098,N_5930);
xnor U6600 (N_6600,N_5748,N_5927);
xor U6601 (N_6601,N_5167,N_5048);
nand U6602 (N_6602,N_5321,N_5315);
nand U6603 (N_6603,N_5179,N_5158);
xnor U6604 (N_6604,N_5974,N_5872);
nand U6605 (N_6605,N_5344,N_5368);
or U6606 (N_6606,N_5790,N_5402);
or U6607 (N_6607,N_5482,N_5819);
and U6608 (N_6608,N_5631,N_5143);
or U6609 (N_6609,N_5860,N_5709);
nand U6610 (N_6610,N_5839,N_5308);
nand U6611 (N_6611,N_5070,N_5830);
or U6612 (N_6612,N_5820,N_5152);
xnor U6613 (N_6613,N_5215,N_5779);
or U6614 (N_6614,N_5783,N_5330);
xnor U6615 (N_6615,N_5966,N_5824);
or U6616 (N_6616,N_5059,N_5015);
and U6617 (N_6617,N_5508,N_5743);
and U6618 (N_6618,N_5131,N_5867);
or U6619 (N_6619,N_5833,N_5521);
xor U6620 (N_6620,N_5948,N_5598);
nor U6621 (N_6621,N_5548,N_5793);
nand U6622 (N_6622,N_5810,N_5774);
xnor U6623 (N_6623,N_5505,N_5349);
nand U6624 (N_6624,N_5442,N_5246);
nor U6625 (N_6625,N_5105,N_5092);
and U6626 (N_6626,N_5376,N_5943);
xnor U6627 (N_6627,N_5118,N_5517);
nor U6628 (N_6628,N_5122,N_5051);
nor U6629 (N_6629,N_5264,N_5114);
nand U6630 (N_6630,N_5755,N_5764);
xnor U6631 (N_6631,N_5092,N_5321);
or U6632 (N_6632,N_5413,N_5468);
and U6633 (N_6633,N_5559,N_5332);
nor U6634 (N_6634,N_5980,N_5046);
nand U6635 (N_6635,N_5077,N_5756);
xnor U6636 (N_6636,N_5275,N_5162);
nand U6637 (N_6637,N_5567,N_5644);
xnor U6638 (N_6638,N_5905,N_5375);
xor U6639 (N_6639,N_5991,N_5166);
nand U6640 (N_6640,N_5867,N_5778);
and U6641 (N_6641,N_5609,N_5246);
and U6642 (N_6642,N_5761,N_5002);
nor U6643 (N_6643,N_5033,N_5093);
xor U6644 (N_6644,N_5189,N_5313);
xor U6645 (N_6645,N_5846,N_5328);
and U6646 (N_6646,N_5696,N_5782);
or U6647 (N_6647,N_5212,N_5496);
nor U6648 (N_6648,N_5560,N_5612);
nor U6649 (N_6649,N_5109,N_5137);
nor U6650 (N_6650,N_5654,N_5097);
and U6651 (N_6651,N_5322,N_5436);
or U6652 (N_6652,N_5172,N_5463);
or U6653 (N_6653,N_5401,N_5277);
or U6654 (N_6654,N_5165,N_5473);
nand U6655 (N_6655,N_5266,N_5461);
xnor U6656 (N_6656,N_5100,N_5692);
or U6657 (N_6657,N_5711,N_5992);
or U6658 (N_6658,N_5399,N_5406);
nand U6659 (N_6659,N_5052,N_5692);
nor U6660 (N_6660,N_5132,N_5863);
or U6661 (N_6661,N_5642,N_5861);
nand U6662 (N_6662,N_5415,N_5387);
and U6663 (N_6663,N_5121,N_5105);
xnor U6664 (N_6664,N_5169,N_5989);
xor U6665 (N_6665,N_5218,N_5306);
or U6666 (N_6666,N_5843,N_5795);
or U6667 (N_6667,N_5776,N_5866);
xnor U6668 (N_6668,N_5623,N_5923);
nand U6669 (N_6669,N_5847,N_5389);
nor U6670 (N_6670,N_5406,N_5993);
nand U6671 (N_6671,N_5321,N_5977);
nand U6672 (N_6672,N_5059,N_5295);
nand U6673 (N_6673,N_5728,N_5361);
or U6674 (N_6674,N_5126,N_5661);
and U6675 (N_6675,N_5214,N_5385);
and U6676 (N_6676,N_5348,N_5594);
or U6677 (N_6677,N_5470,N_5995);
nand U6678 (N_6678,N_5538,N_5578);
or U6679 (N_6679,N_5802,N_5078);
nand U6680 (N_6680,N_5066,N_5575);
and U6681 (N_6681,N_5687,N_5943);
xnor U6682 (N_6682,N_5053,N_5538);
nand U6683 (N_6683,N_5135,N_5182);
xor U6684 (N_6684,N_5764,N_5653);
and U6685 (N_6685,N_5317,N_5394);
xor U6686 (N_6686,N_5726,N_5502);
xnor U6687 (N_6687,N_5059,N_5035);
nand U6688 (N_6688,N_5904,N_5457);
xor U6689 (N_6689,N_5376,N_5325);
or U6690 (N_6690,N_5360,N_5264);
or U6691 (N_6691,N_5533,N_5114);
nor U6692 (N_6692,N_5876,N_5904);
nand U6693 (N_6693,N_5449,N_5876);
or U6694 (N_6694,N_5449,N_5022);
or U6695 (N_6695,N_5011,N_5746);
nand U6696 (N_6696,N_5475,N_5125);
xor U6697 (N_6697,N_5256,N_5822);
nand U6698 (N_6698,N_5485,N_5688);
and U6699 (N_6699,N_5929,N_5153);
and U6700 (N_6700,N_5655,N_5399);
nor U6701 (N_6701,N_5253,N_5313);
or U6702 (N_6702,N_5454,N_5560);
nor U6703 (N_6703,N_5673,N_5197);
or U6704 (N_6704,N_5389,N_5380);
nand U6705 (N_6705,N_5272,N_5979);
nand U6706 (N_6706,N_5060,N_5773);
xnor U6707 (N_6707,N_5250,N_5521);
xnor U6708 (N_6708,N_5843,N_5311);
nand U6709 (N_6709,N_5525,N_5745);
and U6710 (N_6710,N_5829,N_5704);
nand U6711 (N_6711,N_5029,N_5057);
nor U6712 (N_6712,N_5837,N_5256);
nand U6713 (N_6713,N_5275,N_5524);
nor U6714 (N_6714,N_5704,N_5544);
nand U6715 (N_6715,N_5419,N_5425);
or U6716 (N_6716,N_5931,N_5486);
xnor U6717 (N_6717,N_5629,N_5882);
nor U6718 (N_6718,N_5170,N_5356);
or U6719 (N_6719,N_5373,N_5779);
and U6720 (N_6720,N_5911,N_5918);
or U6721 (N_6721,N_5845,N_5823);
or U6722 (N_6722,N_5720,N_5311);
nor U6723 (N_6723,N_5262,N_5686);
or U6724 (N_6724,N_5191,N_5939);
nor U6725 (N_6725,N_5185,N_5944);
or U6726 (N_6726,N_5793,N_5308);
or U6727 (N_6727,N_5271,N_5229);
and U6728 (N_6728,N_5351,N_5782);
xor U6729 (N_6729,N_5803,N_5155);
or U6730 (N_6730,N_5719,N_5400);
or U6731 (N_6731,N_5652,N_5553);
nor U6732 (N_6732,N_5515,N_5456);
nor U6733 (N_6733,N_5904,N_5833);
and U6734 (N_6734,N_5639,N_5289);
nor U6735 (N_6735,N_5497,N_5679);
nand U6736 (N_6736,N_5432,N_5447);
xnor U6737 (N_6737,N_5361,N_5787);
and U6738 (N_6738,N_5972,N_5122);
or U6739 (N_6739,N_5039,N_5748);
and U6740 (N_6740,N_5523,N_5329);
or U6741 (N_6741,N_5199,N_5551);
xnor U6742 (N_6742,N_5996,N_5446);
nand U6743 (N_6743,N_5534,N_5228);
nor U6744 (N_6744,N_5351,N_5636);
nand U6745 (N_6745,N_5764,N_5972);
or U6746 (N_6746,N_5690,N_5766);
and U6747 (N_6747,N_5655,N_5753);
xnor U6748 (N_6748,N_5775,N_5778);
nand U6749 (N_6749,N_5216,N_5384);
or U6750 (N_6750,N_5644,N_5650);
nand U6751 (N_6751,N_5737,N_5933);
xor U6752 (N_6752,N_5873,N_5190);
nand U6753 (N_6753,N_5852,N_5471);
and U6754 (N_6754,N_5354,N_5800);
and U6755 (N_6755,N_5746,N_5217);
or U6756 (N_6756,N_5159,N_5444);
nor U6757 (N_6757,N_5926,N_5551);
nand U6758 (N_6758,N_5421,N_5465);
xor U6759 (N_6759,N_5912,N_5180);
and U6760 (N_6760,N_5299,N_5581);
and U6761 (N_6761,N_5787,N_5109);
nand U6762 (N_6762,N_5528,N_5023);
and U6763 (N_6763,N_5191,N_5865);
or U6764 (N_6764,N_5021,N_5391);
and U6765 (N_6765,N_5430,N_5668);
or U6766 (N_6766,N_5335,N_5445);
nor U6767 (N_6767,N_5444,N_5105);
or U6768 (N_6768,N_5550,N_5770);
xnor U6769 (N_6769,N_5061,N_5440);
xor U6770 (N_6770,N_5464,N_5329);
nand U6771 (N_6771,N_5019,N_5216);
xor U6772 (N_6772,N_5374,N_5738);
and U6773 (N_6773,N_5881,N_5151);
or U6774 (N_6774,N_5440,N_5408);
xor U6775 (N_6775,N_5347,N_5738);
nand U6776 (N_6776,N_5558,N_5902);
and U6777 (N_6777,N_5729,N_5894);
xor U6778 (N_6778,N_5794,N_5940);
nor U6779 (N_6779,N_5740,N_5801);
or U6780 (N_6780,N_5467,N_5889);
nor U6781 (N_6781,N_5453,N_5448);
xnor U6782 (N_6782,N_5871,N_5024);
nand U6783 (N_6783,N_5493,N_5861);
or U6784 (N_6784,N_5465,N_5837);
xor U6785 (N_6785,N_5297,N_5301);
nor U6786 (N_6786,N_5297,N_5333);
or U6787 (N_6787,N_5432,N_5013);
xor U6788 (N_6788,N_5083,N_5802);
or U6789 (N_6789,N_5120,N_5893);
or U6790 (N_6790,N_5103,N_5983);
or U6791 (N_6791,N_5853,N_5978);
xor U6792 (N_6792,N_5132,N_5960);
nor U6793 (N_6793,N_5783,N_5017);
nor U6794 (N_6794,N_5813,N_5940);
xor U6795 (N_6795,N_5545,N_5220);
xnor U6796 (N_6796,N_5733,N_5008);
and U6797 (N_6797,N_5644,N_5258);
xor U6798 (N_6798,N_5664,N_5569);
nor U6799 (N_6799,N_5516,N_5095);
and U6800 (N_6800,N_5468,N_5586);
nor U6801 (N_6801,N_5559,N_5749);
nor U6802 (N_6802,N_5193,N_5733);
xor U6803 (N_6803,N_5138,N_5724);
xor U6804 (N_6804,N_5583,N_5782);
nor U6805 (N_6805,N_5860,N_5820);
nand U6806 (N_6806,N_5893,N_5895);
nor U6807 (N_6807,N_5856,N_5915);
and U6808 (N_6808,N_5077,N_5076);
xnor U6809 (N_6809,N_5335,N_5757);
or U6810 (N_6810,N_5821,N_5989);
and U6811 (N_6811,N_5328,N_5064);
nand U6812 (N_6812,N_5622,N_5442);
nand U6813 (N_6813,N_5994,N_5957);
and U6814 (N_6814,N_5273,N_5111);
nor U6815 (N_6815,N_5198,N_5779);
or U6816 (N_6816,N_5848,N_5683);
xor U6817 (N_6817,N_5448,N_5383);
or U6818 (N_6818,N_5716,N_5630);
nand U6819 (N_6819,N_5712,N_5869);
nand U6820 (N_6820,N_5661,N_5476);
and U6821 (N_6821,N_5978,N_5536);
xnor U6822 (N_6822,N_5309,N_5389);
nand U6823 (N_6823,N_5943,N_5756);
xnor U6824 (N_6824,N_5559,N_5647);
nand U6825 (N_6825,N_5357,N_5998);
and U6826 (N_6826,N_5296,N_5416);
nand U6827 (N_6827,N_5853,N_5235);
or U6828 (N_6828,N_5366,N_5708);
or U6829 (N_6829,N_5604,N_5348);
xor U6830 (N_6830,N_5261,N_5397);
nand U6831 (N_6831,N_5963,N_5509);
and U6832 (N_6832,N_5127,N_5811);
and U6833 (N_6833,N_5569,N_5043);
xnor U6834 (N_6834,N_5642,N_5310);
or U6835 (N_6835,N_5483,N_5707);
and U6836 (N_6836,N_5740,N_5852);
or U6837 (N_6837,N_5664,N_5861);
or U6838 (N_6838,N_5460,N_5534);
xor U6839 (N_6839,N_5999,N_5096);
xnor U6840 (N_6840,N_5418,N_5249);
xnor U6841 (N_6841,N_5413,N_5471);
xnor U6842 (N_6842,N_5729,N_5573);
xnor U6843 (N_6843,N_5866,N_5564);
nor U6844 (N_6844,N_5924,N_5325);
xor U6845 (N_6845,N_5769,N_5043);
xnor U6846 (N_6846,N_5887,N_5978);
and U6847 (N_6847,N_5787,N_5833);
nor U6848 (N_6848,N_5183,N_5701);
or U6849 (N_6849,N_5960,N_5144);
or U6850 (N_6850,N_5771,N_5696);
or U6851 (N_6851,N_5045,N_5503);
nor U6852 (N_6852,N_5462,N_5067);
and U6853 (N_6853,N_5254,N_5083);
and U6854 (N_6854,N_5236,N_5367);
nor U6855 (N_6855,N_5488,N_5776);
and U6856 (N_6856,N_5668,N_5943);
xnor U6857 (N_6857,N_5099,N_5211);
and U6858 (N_6858,N_5714,N_5626);
nand U6859 (N_6859,N_5731,N_5569);
xor U6860 (N_6860,N_5951,N_5510);
or U6861 (N_6861,N_5927,N_5108);
or U6862 (N_6862,N_5905,N_5771);
and U6863 (N_6863,N_5377,N_5230);
or U6864 (N_6864,N_5123,N_5606);
xnor U6865 (N_6865,N_5402,N_5316);
xnor U6866 (N_6866,N_5807,N_5489);
xor U6867 (N_6867,N_5418,N_5784);
nor U6868 (N_6868,N_5304,N_5397);
and U6869 (N_6869,N_5345,N_5290);
or U6870 (N_6870,N_5477,N_5412);
and U6871 (N_6871,N_5052,N_5572);
xor U6872 (N_6872,N_5963,N_5031);
and U6873 (N_6873,N_5275,N_5051);
nand U6874 (N_6874,N_5467,N_5150);
and U6875 (N_6875,N_5988,N_5972);
xor U6876 (N_6876,N_5076,N_5959);
nand U6877 (N_6877,N_5003,N_5530);
xor U6878 (N_6878,N_5608,N_5832);
or U6879 (N_6879,N_5904,N_5503);
xor U6880 (N_6880,N_5859,N_5111);
nand U6881 (N_6881,N_5824,N_5669);
xnor U6882 (N_6882,N_5540,N_5413);
xnor U6883 (N_6883,N_5485,N_5723);
or U6884 (N_6884,N_5306,N_5087);
or U6885 (N_6885,N_5197,N_5848);
or U6886 (N_6886,N_5038,N_5555);
xor U6887 (N_6887,N_5572,N_5240);
nand U6888 (N_6888,N_5644,N_5956);
nor U6889 (N_6889,N_5540,N_5453);
xor U6890 (N_6890,N_5876,N_5514);
nand U6891 (N_6891,N_5538,N_5891);
nand U6892 (N_6892,N_5116,N_5885);
xnor U6893 (N_6893,N_5925,N_5754);
and U6894 (N_6894,N_5845,N_5591);
and U6895 (N_6895,N_5124,N_5181);
nor U6896 (N_6896,N_5273,N_5209);
nor U6897 (N_6897,N_5477,N_5512);
nand U6898 (N_6898,N_5151,N_5459);
and U6899 (N_6899,N_5032,N_5082);
nand U6900 (N_6900,N_5806,N_5658);
or U6901 (N_6901,N_5752,N_5767);
or U6902 (N_6902,N_5078,N_5155);
and U6903 (N_6903,N_5078,N_5475);
xor U6904 (N_6904,N_5649,N_5463);
nor U6905 (N_6905,N_5123,N_5683);
nand U6906 (N_6906,N_5977,N_5522);
xnor U6907 (N_6907,N_5685,N_5020);
xor U6908 (N_6908,N_5842,N_5583);
xor U6909 (N_6909,N_5461,N_5563);
and U6910 (N_6910,N_5554,N_5921);
xnor U6911 (N_6911,N_5975,N_5016);
xor U6912 (N_6912,N_5093,N_5626);
nor U6913 (N_6913,N_5667,N_5328);
xnor U6914 (N_6914,N_5702,N_5917);
or U6915 (N_6915,N_5345,N_5979);
and U6916 (N_6916,N_5510,N_5289);
nor U6917 (N_6917,N_5029,N_5792);
nor U6918 (N_6918,N_5417,N_5262);
or U6919 (N_6919,N_5830,N_5089);
nor U6920 (N_6920,N_5708,N_5349);
xor U6921 (N_6921,N_5998,N_5185);
xor U6922 (N_6922,N_5667,N_5308);
xor U6923 (N_6923,N_5995,N_5693);
xnor U6924 (N_6924,N_5515,N_5931);
nand U6925 (N_6925,N_5683,N_5190);
nand U6926 (N_6926,N_5728,N_5302);
nand U6927 (N_6927,N_5078,N_5237);
xor U6928 (N_6928,N_5993,N_5356);
xnor U6929 (N_6929,N_5013,N_5497);
nand U6930 (N_6930,N_5258,N_5159);
nor U6931 (N_6931,N_5202,N_5487);
or U6932 (N_6932,N_5811,N_5579);
nor U6933 (N_6933,N_5393,N_5460);
xnor U6934 (N_6934,N_5166,N_5653);
nand U6935 (N_6935,N_5392,N_5267);
and U6936 (N_6936,N_5018,N_5590);
nor U6937 (N_6937,N_5731,N_5623);
or U6938 (N_6938,N_5951,N_5288);
nand U6939 (N_6939,N_5300,N_5755);
nor U6940 (N_6940,N_5176,N_5264);
nor U6941 (N_6941,N_5240,N_5345);
nand U6942 (N_6942,N_5976,N_5682);
or U6943 (N_6943,N_5762,N_5829);
or U6944 (N_6944,N_5348,N_5704);
and U6945 (N_6945,N_5198,N_5302);
xnor U6946 (N_6946,N_5784,N_5865);
nor U6947 (N_6947,N_5410,N_5294);
nor U6948 (N_6948,N_5071,N_5364);
nand U6949 (N_6949,N_5164,N_5536);
xor U6950 (N_6950,N_5092,N_5774);
or U6951 (N_6951,N_5220,N_5565);
nand U6952 (N_6952,N_5153,N_5017);
or U6953 (N_6953,N_5887,N_5061);
and U6954 (N_6954,N_5415,N_5640);
and U6955 (N_6955,N_5783,N_5015);
xor U6956 (N_6956,N_5993,N_5594);
nand U6957 (N_6957,N_5479,N_5790);
nor U6958 (N_6958,N_5672,N_5616);
or U6959 (N_6959,N_5515,N_5421);
and U6960 (N_6960,N_5521,N_5150);
nor U6961 (N_6961,N_5843,N_5484);
and U6962 (N_6962,N_5980,N_5059);
nand U6963 (N_6963,N_5475,N_5103);
nand U6964 (N_6964,N_5011,N_5243);
nand U6965 (N_6965,N_5667,N_5179);
nand U6966 (N_6966,N_5871,N_5041);
or U6967 (N_6967,N_5630,N_5749);
nor U6968 (N_6968,N_5613,N_5747);
nor U6969 (N_6969,N_5689,N_5086);
nand U6970 (N_6970,N_5413,N_5559);
or U6971 (N_6971,N_5154,N_5357);
nor U6972 (N_6972,N_5801,N_5268);
and U6973 (N_6973,N_5936,N_5799);
nor U6974 (N_6974,N_5659,N_5984);
nor U6975 (N_6975,N_5221,N_5773);
nor U6976 (N_6976,N_5247,N_5771);
nor U6977 (N_6977,N_5500,N_5020);
nand U6978 (N_6978,N_5882,N_5535);
or U6979 (N_6979,N_5013,N_5946);
xor U6980 (N_6980,N_5523,N_5210);
nor U6981 (N_6981,N_5796,N_5500);
nor U6982 (N_6982,N_5488,N_5446);
or U6983 (N_6983,N_5199,N_5769);
xor U6984 (N_6984,N_5487,N_5120);
or U6985 (N_6985,N_5149,N_5559);
or U6986 (N_6986,N_5577,N_5086);
or U6987 (N_6987,N_5548,N_5590);
and U6988 (N_6988,N_5852,N_5177);
and U6989 (N_6989,N_5695,N_5219);
and U6990 (N_6990,N_5570,N_5610);
nor U6991 (N_6991,N_5607,N_5462);
xor U6992 (N_6992,N_5959,N_5336);
or U6993 (N_6993,N_5968,N_5919);
nand U6994 (N_6994,N_5803,N_5633);
nand U6995 (N_6995,N_5437,N_5065);
xor U6996 (N_6996,N_5624,N_5949);
nand U6997 (N_6997,N_5090,N_5970);
and U6998 (N_6998,N_5984,N_5241);
or U6999 (N_6999,N_5144,N_5931);
or U7000 (N_7000,N_6117,N_6667);
nand U7001 (N_7001,N_6610,N_6477);
and U7002 (N_7002,N_6339,N_6185);
or U7003 (N_7003,N_6332,N_6001);
nor U7004 (N_7004,N_6343,N_6545);
nor U7005 (N_7005,N_6944,N_6769);
nand U7006 (N_7006,N_6213,N_6181);
xor U7007 (N_7007,N_6814,N_6523);
xnor U7008 (N_7008,N_6945,N_6015);
or U7009 (N_7009,N_6754,N_6377);
and U7010 (N_7010,N_6927,N_6497);
nand U7011 (N_7011,N_6660,N_6065);
nand U7012 (N_7012,N_6883,N_6128);
nand U7013 (N_7013,N_6305,N_6723);
and U7014 (N_7014,N_6369,N_6420);
nor U7015 (N_7015,N_6300,N_6784);
and U7016 (N_7016,N_6929,N_6159);
or U7017 (N_7017,N_6187,N_6672);
nand U7018 (N_7018,N_6245,N_6834);
nand U7019 (N_7019,N_6280,N_6857);
and U7020 (N_7020,N_6625,N_6830);
nor U7021 (N_7021,N_6718,N_6948);
nand U7022 (N_7022,N_6078,N_6094);
nand U7023 (N_7023,N_6768,N_6992);
or U7024 (N_7024,N_6861,N_6234);
nand U7025 (N_7025,N_6100,N_6049);
nand U7026 (N_7026,N_6736,N_6169);
nand U7027 (N_7027,N_6445,N_6961);
or U7028 (N_7028,N_6017,N_6429);
xnor U7029 (N_7029,N_6743,N_6330);
or U7030 (N_7030,N_6876,N_6634);
nand U7031 (N_7031,N_6451,N_6557);
or U7032 (N_7032,N_6592,N_6644);
and U7033 (N_7033,N_6681,N_6030);
xnor U7034 (N_7034,N_6647,N_6337);
or U7035 (N_7035,N_6528,N_6400);
nor U7036 (N_7036,N_6033,N_6608);
nor U7037 (N_7037,N_6721,N_6527);
and U7038 (N_7038,N_6309,N_6967);
nand U7039 (N_7039,N_6771,N_6886);
nor U7040 (N_7040,N_6498,N_6387);
and U7041 (N_7041,N_6188,N_6285);
and U7042 (N_7042,N_6818,N_6071);
xnor U7043 (N_7043,N_6690,N_6887);
xnor U7044 (N_7044,N_6151,N_6266);
and U7045 (N_7045,N_6877,N_6101);
or U7046 (N_7046,N_6711,N_6686);
nor U7047 (N_7047,N_6202,N_6352);
xnor U7048 (N_7048,N_6542,N_6095);
and U7049 (N_7049,N_6798,N_6006);
xnor U7050 (N_7050,N_6239,N_6888);
nor U7051 (N_7051,N_6493,N_6930);
nand U7052 (N_7052,N_6620,N_6119);
nor U7053 (N_7053,N_6727,N_6765);
or U7054 (N_7054,N_6042,N_6990);
and U7055 (N_7055,N_6507,N_6054);
nand U7056 (N_7056,N_6916,N_6260);
nor U7057 (N_7057,N_6465,N_6406);
xnor U7058 (N_7058,N_6565,N_6298);
nor U7059 (N_7059,N_6136,N_6749);
xor U7060 (N_7060,N_6212,N_6748);
and U7061 (N_7061,N_6601,N_6165);
and U7062 (N_7062,N_6589,N_6342);
and U7063 (N_7063,N_6132,N_6518);
xnor U7064 (N_7064,N_6413,N_6824);
or U7065 (N_7065,N_6085,N_6368);
xnor U7066 (N_7066,N_6700,N_6841);
or U7067 (N_7067,N_6879,N_6444);
xor U7068 (N_7068,N_6316,N_6147);
and U7069 (N_7069,N_6904,N_6863);
and U7070 (N_7070,N_6198,N_6770);
nor U7071 (N_7071,N_6963,N_6899);
nand U7072 (N_7072,N_6050,N_6773);
or U7073 (N_7073,N_6433,N_6763);
and U7074 (N_7074,N_6885,N_6868);
and U7075 (N_7075,N_6027,N_6709);
or U7076 (N_7076,N_6520,N_6115);
and U7077 (N_7077,N_6227,N_6687);
and U7078 (N_7078,N_6402,N_6106);
or U7079 (N_7079,N_6999,N_6807);
xnor U7080 (N_7080,N_6262,N_6203);
xnor U7081 (N_7081,N_6673,N_6813);
or U7082 (N_7082,N_6446,N_6210);
or U7083 (N_7083,N_6215,N_6612);
xor U7084 (N_7084,N_6591,N_6574);
and U7085 (N_7085,N_6781,N_6725);
or U7086 (N_7086,N_6416,N_6192);
nor U7087 (N_7087,N_6167,N_6907);
xor U7088 (N_7088,N_6541,N_6606);
or U7089 (N_7089,N_6615,N_6423);
nor U7090 (N_7090,N_6326,N_6750);
nand U7091 (N_7091,N_6645,N_6256);
or U7092 (N_7092,N_6597,N_6636);
nor U7093 (N_7093,N_6800,N_6914);
xnor U7094 (N_7094,N_6452,N_6123);
nand U7095 (N_7095,N_6252,N_6583);
xnor U7096 (N_7096,N_6981,N_6832);
or U7097 (N_7097,N_6380,N_6469);
or U7098 (N_7098,N_6087,N_6678);
or U7099 (N_7099,N_6120,N_6910);
and U7100 (N_7100,N_6270,N_6261);
nand U7101 (N_7101,N_6255,N_6531);
or U7102 (N_7102,N_6079,N_6959);
xnor U7103 (N_7103,N_6741,N_6635);
nor U7104 (N_7104,N_6640,N_6535);
nor U7105 (N_7105,N_6848,N_6873);
xnor U7106 (N_7106,N_6683,N_6793);
xor U7107 (N_7107,N_6061,N_6180);
or U7108 (N_7108,N_6013,N_6826);
nand U7109 (N_7109,N_6066,N_6787);
xor U7110 (N_7110,N_6953,N_6627);
and U7111 (N_7111,N_6447,N_6599);
nand U7112 (N_7112,N_6011,N_6418);
nor U7113 (N_7113,N_6383,N_6467);
xnor U7114 (N_7114,N_6072,N_6797);
and U7115 (N_7115,N_6211,N_6568);
nor U7116 (N_7116,N_6143,N_6614);
nor U7117 (N_7117,N_6836,N_6121);
xnor U7118 (N_7118,N_6384,N_6464);
nor U7119 (N_7119,N_6980,N_6827);
or U7120 (N_7120,N_6733,N_6555);
and U7121 (N_7121,N_6391,N_6297);
nor U7122 (N_7122,N_6294,N_6140);
nand U7123 (N_7123,N_6398,N_6379);
or U7124 (N_7124,N_6319,N_6291);
xnor U7125 (N_7125,N_6840,N_6746);
xnor U7126 (N_7126,N_6516,N_6225);
xnor U7127 (N_7127,N_6704,N_6460);
or U7128 (N_7128,N_6127,N_6373);
nor U7129 (N_7129,N_6880,N_6590);
and U7130 (N_7130,N_6903,N_6160);
xor U7131 (N_7131,N_6974,N_6064);
nor U7132 (N_7132,N_6110,N_6549);
nand U7133 (N_7133,N_6412,N_6524);
nand U7134 (N_7134,N_6329,N_6149);
nor U7135 (N_7135,N_6485,N_6053);
or U7136 (N_7136,N_6805,N_6772);
nand U7137 (N_7137,N_6462,N_6175);
and U7138 (N_7138,N_6442,N_6569);
nor U7139 (N_7139,N_6321,N_6775);
and U7140 (N_7140,N_6970,N_6706);
nor U7141 (N_7141,N_6367,N_6108);
nor U7142 (N_7142,N_6891,N_6751);
or U7143 (N_7143,N_6005,N_6401);
nand U7144 (N_7144,N_6244,N_6925);
and U7145 (N_7145,N_6098,N_6301);
nor U7146 (N_7146,N_6675,N_6920);
and U7147 (N_7147,N_6074,N_6652);
xnor U7148 (N_7148,N_6338,N_6278);
nand U7149 (N_7149,N_6694,N_6734);
or U7150 (N_7150,N_6443,N_6633);
xnor U7151 (N_7151,N_6676,N_6405);
nand U7152 (N_7152,N_6866,N_6157);
and U7153 (N_7153,N_6272,N_6014);
xnor U7154 (N_7154,N_6954,N_6637);
nand U7155 (N_7155,N_6372,N_6985);
nor U7156 (N_7156,N_6209,N_6511);
or U7157 (N_7157,N_6825,N_6533);
and U7158 (N_7158,N_6839,N_6314);
or U7159 (N_7159,N_6624,N_6317);
nor U7160 (N_7160,N_6302,N_6327);
nand U7161 (N_7161,N_6560,N_6141);
and U7162 (N_7162,N_6801,N_6055);
or U7163 (N_7163,N_6928,N_6996);
or U7164 (N_7164,N_6295,N_6796);
nand U7165 (N_7165,N_6747,N_6695);
nor U7166 (N_7166,N_6231,N_6938);
or U7167 (N_7167,N_6414,N_6148);
and U7168 (N_7168,N_6193,N_6434);
or U7169 (N_7169,N_6435,N_6578);
nand U7170 (N_7170,N_6243,N_6788);
xor U7171 (N_7171,N_6281,N_6501);
nor U7172 (N_7172,N_6154,N_6968);
and U7173 (N_7173,N_6259,N_6835);
nor U7174 (N_7174,N_6171,N_6605);
xor U7175 (N_7175,N_6097,N_6570);
and U7176 (N_7176,N_6922,N_6410);
xnor U7177 (N_7177,N_6290,N_6942);
nand U7178 (N_7178,N_6395,N_6470);
nand U7179 (N_7179,N_6018,N_6086);
nand U7180 (N_7180,N_6911,N_6490);
or U7181 (N_7181,N_6240,N_6287);
and U7182 (N_7182,N_6719,N_6688);
xnor U7183 (N_7183,N_6525,N_6728);
nor U7184 (N_7184,N_6463,N_6973);
or U7185 (N_7185,N_6292,N_6726);
xnor U7186 (N_7186,N_6993,N_6691);
nor U7187 (N_7187,N_6284,N_6932);
or U7188 (N_7188,N_6921,N_6514);
or U7189 (N_7189,N_6776,N_6440);
nand U7190 (N_7190,N_6360,N_6096);
nand U7191 (N_7191,N_6919,N_6851);
xnor U7192 (N_7192,N_6038,N_6817);
nand U7193 (N_7193,N_6865,N_6466);
nand U7194 (N_7194,N_6665,N_6481);
xnor U7195 (N_7195,N_6092,N_6575);
and U7196 (N_7196,N_6035,N_6492);
or U7197 (N_7197,N_6168,N_6254);
xor U7198 (N_7198,N_6714,N_6965);
nor U7199 (N_7199,N_6803,N_6204);
or U7200 (N_7200,N_6226,N_6902);
xor U7201 (N_7201,N_6689,N_6764);
nand U7202 (N_7202,N_6331,N_6924);
and U7203 (N_7203,N_6178,N_6145);
xnor U7204 (N_7204,N_6219,N_6347);
nand U7205 (N_7205,N_6346,N_6562);
and U7206 (N_7206,N_6758,N_6333);
xnor U7207 (N_7207,N_6238,N_6829);
nand U7208 (N_7208,N_6941,N_6271);
nor U7209 (N_7209,N_6311,N_6220);
and U7210 (N_7210,N_6617,N_6604);
nor U7211 (N_7211,N_6454,N_6125);
nor U7212 (N_7212,N_6618,N_6532);
nor U7213 (N_7213,N_6517,N_6376);
nor U7214 (N_7214,N_6002,N_6642);
or U7215 (N_7215,N_6815,N_6025);
or U7216 (N_7216,N_6559,N_6708);
or U7217 (N_7217,N_6623,N_6896);
nor U7218 (N_7218,N_6988,N_6872);
nand U7219 (N_7219,N_6643,N_6007);
nor U7220 (N_7220,N_6289,N_6579);
xor U7221 (N_7221,N_6735,N_6046);
nand U7222 (N_7222,N_6890,N_6389);
and U7223 (N_7223,N_6200,N_6712);
or U7224 (N_7224,N_6739,N_6176);
or U7225 (N_7225,N_6744,N_6685);
or U7226 (N_7226,N_6947,N_6804);
nor U7227 (N_7227,N_6207,N_6931);
xnor U7228 (N_7228,N_6611,N_6340);
and U7229 (N_7229,N_6546,N_6503);
nor U7230 (N_7230,N_6051,N_6453);
or U7231 (N_7231,N_6653,N_6091);
or U7232 (N_7232,N_6581,N_6162);
nand U7233 (N_7233,N_6842,N_6431);
or U7234 (N_7234,N_6553,N_6052);
and U7235 (N_7235,N_6142,N_6926);
xnor U7236 (N_7236,N_6461,N_6702);
nand U7237 (N_7237,N_6631,N_6161);
nand U7238 (N_7238,N_6519,N_6320);
nand U7239 (N_7239,N_6940,N_6247);
xor U7240 (N_7240,N_6021,N_6875);
nand U7241 (N_7241,N_6296,N_6855);
xnor U7242 (N_7242,N_6669,N_6044);
or U7243 (N_7243,N_6224,N_6566);
and U7244 (N_7244,N_6774,N_6135);
nand U7245 (N_7245,N_6201,N_6551);
nor U7246 (N_7246,N_6828,N_6915);
nor U7247 (N_7247,N_6056,N_6126);
nand U7248 (N_7248,N_6595,N_6757);
or U7249 (N_7249,N_6138,N_6441);
and U7250 (N_7250,N_6205,N_6859);
or U7251 (N_7251,N_6365,N_6472);
nand U7252 (N_7252,N_6697,N_6471);
xnor U7253 (N_7253,N_6102,N_6680);
and U7254 (N_7254,N_6268,N_6286);
and U7255 (N_7255,N_6600,N_6698);
and U7256 (N_7256,N_6458,N_6629);
or U7257 (N_7257,N_6639,N_6577);
and U7258 (N_7258,N_6273,N_6455);
nor U7259 (N_7259,N_6449,N_6468);
xnor U7260 (N_7260,N_6567,N_6515);
or U7261 (N_7261,N_6955,N_6731);
nand U7262 (N_7262,N_6960,N_6076);
nand U7263 (N_7263,N_6073,N_6923);
nand U7264 (N_7264,N_6847,N_6808);
nor U7265 (N_7265,N_6693,N_6109);
or U7266 (N_7266,N_6217,N_6022);
xor U7267 (N_7267,N_6664,N_6303);
nand U7268 (N_7268,N_6118,N_6889);
and U7269 (N_7269,N_6190,N_6821);
nand U7270 (N_7270,N_6388,N_6392);
and U7271 (N_7271,N_6032,N_6208);
xor U7272 (N_7272,N_6436,N_6191);
nand U7273 (N_7273,N_6075,N_6062);
and U7274 (N_7274,N_6279,N_6170);
nand U7275 (N_7275,N_6802,N_6315);
nand U7276 (N_7276,N_6473,N_6177);
nor U7277 (N_7277,N_6584,N_6666);
xnor U7278 (N_7278,N_6133,N_6060);
xnor U7279 (N_7279,N_6031,N_6674);
nand U7280 (N_7280,N_6103,N_6554);
nor U7281 (N_7281,N_6753,N_6586);
nand U7282 (N_7282,N_6283,N_6358);
nor U7283 (N_7283,N_6632,N_6760);
and U7284 (N_7284,N_6040,N_6496);
or U7285 (N_7285,N_6166,N_6396);
and U7286 (N_7286,N_6799,N_6513);
xnor U7287 (N_7287,N_6385,N_6856);
nor U7288 (N_7288,N_6587,N_6696);
nor U7289 (N_7289,N_6901,N_6082);
nor U7290 (N_7290,N_6487,N_6048);
nand U7291 (N_7291,N_6214,N_6415);
and U7292 (N_7292,N_6703,N_6083);
nor U7293 (N_7293,N_6732,N_6036);
xnor U7294 (N_7294,N_6233,N_6322);
and U7295 (N_7295,N_6229,N_6364);
or U7296 (N_7296,N_6081,N_6806);
and U7297 (N_7297,N_6510,N_6752);
and U7298 (N_7298,N_6494,N_6670);
or U7299 (N_7299,N_6218,N_6276);
or U7300 (N_7300,N_6112,N_6241);
and U7301 (N_7301,N_6619,N_6235);
and U7302 (N_7302,N_6277,N_6113);
nor U7303 (N_7303,N_6543,N_6646);
or U7304 (N_7304,N_6616,N_6716);
xor U7305 (N_7305,N_6648,N_6016);
nand U7306 (N_7306,N_6088,N_6020);
or U7307 (N_7307,N_6194,N_6762);
or U7308 (N_7308,N_6246,N_6009);
xor U7309 (N_7309,N_6898,N_6474);
and U7310 (N_7310,N_6846,N_6344);
nor U7311 (N_7311,N_6304,N_6484);
nor U7312 (N_7312,N_6263,N_6966);
nor U7313 (N_7313,N_6371,N_6386);
xnor U7314 (N_7314,N_6596,N_6172);
nor U7315 (N_7315,N_6399,N_6068);
or U7316 (N_7316,N_6023,N_6351);
and U7317 (N_7317,N_6867,N_6356);
nand U7318 (N_7318,N_6375,N_6004);
or U7319 (N_7319,N_6849,N_6782);
xnor U7320 (N_7320,N_6977,N_6390);
and U7321 (N_7321,N_6656,N_6958);
and U7322 (N_7322,N_6534,N_6488);
nor U7323 (N_7323,N_6738,N_6174);
and U7324 (N_7324,N_6745,N_6427);
and U7325 (N_7325,N_6905,N_6323);
nor U7326 (N_7326,N_6370,N_6978);
nand U7327 (N_7327,N_6328,N_6936);
and U7328 (N_7328,N_6838,N_6158);
nor U7329 (N_7329,N_6104,N_6306);
xnor U7330 (N_7330,N_6107,N_6251);
nand U7331 (N_7331,N_6090,N_6508);
nor U7332 (N_7332,N_6037,N_6593);
or U7333 (N_7333,N_6459,N_6854);
nor U7334 (N_7334,N_6724,N_6003);
nor U7335 (N_7335,N_6114,N_6893);
nor U7336 (N_7336,N_6144,N_6348);
and U7337 (N_7337,N_6506,N_6236);
nor U7338 (N_7338,N_6341,N_6428);
or U7339 (N_7339,N_6495,N_6408);
or U7340 (N_7340,N_6070,N_6195);
xor U7341 (N_7341,N_6785,N_6288);
xnor U7342 (N_7342,N_6638,N_6318);
nor U7343 (N_7343,N_6491,N_6779);
xor U7344 (N_7344,N_6173,N_6199);
nand U7345 (N_7345,N_6819,N_6561);
xor U7346 (N_7346,N_6994,N_6935);
nor U7347 (N_7347,N_6912,N_6852);
and U7348 (N_7348,N_6892,N_6478);
and U7349 (N_7349,N_6823,N_6984);
or U7350 (N_7350,N_6979,N_6057);
nand U7351 (N_7351,N_6809,N_6661);
xnor U7352 (N_7352,N_6426,N_6182);
nor U7353 (N_7353,N_6995,N_6603);
nor U7354 (N_7354,N_6184,N_6918);
xnor U7355 (N_7355,N_6982,N_6430);
and U7356 (N_7356,N_6780,N_6164);
and U7357 (N_7357,N_6312,N_6345);
nor U7358 (N_7358,N_6336,N_6437);
nand U7359 (N_7359,N_6621,N_6105);
nand U7360 (N_7360,N_6684,N_6419);
xor U7361 (N_7361,N_6221,N_6335);
nor U7362 (N_7362,N_6794,N_6655);
or U7363 (N_7363,N_6662,N_6130);
xor U7364 (N_7364,N_6366,N_6382);
nand U7365 (N_7365,N_6269,N_6862);
and U7366 (N_7366,N_6964,N_6833);
and U7367 (N_7367,N_6650,N_6869);
nor U7368 (N_7368,N_6715,N_6539);
nor U7369 (N_7369,N_6179,N_6206);
and U7370 (N_7370,N_6069,N_6124);
or U7371 (N_7371,N_6908,N_6536);
and U7372 (N_7372,N_6786,N_6699);
and U7373 (N_7373,N_6357,N_6626);
nor U7374 (N_7374,N_6576,N_6730);
and U7375 (N_7375,N_6755,N_6394);
and U7376 (N_7376,N_6475,N_6223);
xnor U7377 (N_7377,N_6939,N_6080);
and U7378 (N_7378,N_6537,N_6111);
and U7379 (N_7379,N_6264,N_6909);
nand U7380 (N_7380,N_6480,N_6767);
or U7381 (N_7381,N_6933,N_6010);
nor U7382 (N_7382,N_6265,N_6232);
and U7383 (N_7383,N_6237,N_6099);
and U7384 (N_7384,N_6630,N_6654);
xor U7385 (N_7385,N_6063,N_6155);
nor U7386 (N_7386,N_6267,N_6024);
xnor U7387 (N_7387,N_6409,N_6969);
or U7388 (N_7388,N_6355,N_6564);
and U7389 (N_7389,N_6489,N_6189);
nand U7390 (N_7390,N_6622,N_6822);
nand U7391 (N_7391,N_6354,N_6540);
and U7392 (N_7392,N_6359,N_6729);
and U7393 (N_7393,N_6526,N_6811);
and U7394 (N_7394,N_6722,N_6677);
xnor U7395 (N_7395,N_6843,N_6607);
nor U7396 (N_7396,N_6810,N_6361);
nor U7397 (N_7397,N_6432,N_6242);
xnor U7398 (N_7398,N_6448,N_6282);
nand U7399 (N_7399,N_6831,N_6183);
or U7400 (N_7400,N_6084,N_6222);
or U7401 (N_7401,N_6663,N_6350);
or U7402 (N_7402,N_6353,N_6783);
or U7403 (N_7403,N_6791,N_6882);
xnor U7404 (N_7404,N_6906,N_6740);
nand U7405 (N_7405,N_6059,N_6609);
xnor U7406 (N_7406,N_6766,N_6668);
xor U7407 (N_7407,N_6613,N_6482);
xnor U7408 (N_7408,N_6778,N_6486);
or U7409 (N_7409,N_6934,N_6000);
xnor U7410 (N_7410,N_6334,N_6972);
or U7411 (N_7411,N_6742,N_6324);
and U7412 (N_7412,N_6790,N_6381);
or U7413 (N_7413,N_6393,N_6837);
or U7414 (N_7414,N_6820,N_6864);
and U7415 (N_7415,N_6950,N_6710);
or U7416 (N_7416,N_6047,N_6571);
or U7417 (N_7417,N_6129,N_6156);
nor U7418 (N_7418,N_6844,N_6761);
and U7419 (N_7419,N_6956,N_6012);
nor U7420 (N_7420,N_6884,N_6558);
nor U7421 (N_7421,N_6483,N_6310);
and U7422 (N_7422,N_6067,N_6937);
nand U7423 (N_7423,N_6530,N_6991);
nand U7424 (N_7424,N_6045,N_6216);
nand U7425 (N_7425,N_6499,N_6682);
or U7426 (N_7426,N_6858,N_6572);
nand U7427 (N_7427,N_6248,N_6362);
and U7428 (N_7428,N_6756,N_6089);
nor U7429 (N_7429,N_6792,N_6547);
nor U7430 (N_7430,N_6957,N_6504);
or U7431 (N_7431,N_6186,N_6580);
xnor U7432 (N_7432,N_6152,N_6522);
nand U7433 (N_7433,N_6308,N_6895);
nand U7434 (N_7434,N_6421,N_6422);
nor U7435 (N_7435,N_6573,N_6594);
nand U7436 (N_7436,N_6476,N_6363);
nand U7437 (N_7437,N_6093,N_6325);
xnor U7438 (N_7438,N_6692,N_6249);
and U7439 (N_7439,N_6008,N_6917);
nor U7440 (N_7440,N_6812,N_6258);
or U7441 (N_7441,N_6707,N_6986);
nor U7442 (N_7442,N_6424,N_6439);
nor U7443 (N_7443,N_6479,N_6552);
xor U7444 (N_7444,N_6795,N_6043);
and U7445 (N_7445,N_6041,N_6456);
xor U7446 (N_7446,N_6989,N_6871);
nor U7447 (N_7447,N_6962,N_6860);
or U7448 (N_7448,N_6897,N_6556);
nand U7449 (N_7449,N_6197,N_6987);
xor U7450 (N_7450,N_6307,N_6538);
xor U7451 (N_7451,N_6874,N_6137);
and U7452 (N_7452,N_6228,N_6500);
nand U7453 (N_7453,N_6313,N_6878);
and U7454 (N_7454,N_6713,N_6529);
or U7455 (N_7455,N_6975,N_6998);
nor U7456 (N_7456,N_6582,N_6275);
or U7457 (N_7457,N_6628,N_6705);
nand U7458 (N_7458,N_6026,N_6509);
and U7459 (N_7459,N_6900,N_6983);
xnor U7460 (N_7460,N_6777,N_6657);
xnor U7461 (N_7461,N_6374,N_6034);
nand U7462 (N_7462,N_6971,N_6403);
or U7463 (N_7463,N_6585,N_6163);
nand U7464 (N_7464,N_6505,N_6122);
or U7465 (N_7465,N_6378,N_6146);
nand U7466 (N_7466,N_6274,N_6134);
and U7467 (N_7467,N_6028,N_6425);
xnor U7468 (N_7468,N_6139,N_6450);
and U7469 (N_7469,N_6548,N_6720);
or U7470 (N_7470,N_6943,N_6976);
or U7471 (N_7471,N_6651,N_6913);
xnor U7472 (N_7472,N_6077,N_6997);
nor U7473 (N_7473,N_6230,N_6397);
and U7474 (N_7474,N_6457,N_6293);
nor U7475 (N_7475,N_6521,N_6701);
nor U7476 (N_7476,N_6257,N_6641);
and U7477 (N_7477,N_6588,N_6658);
xor U7478 (N_7478,N_6131,N_6299);
and U7479 (N_7479,N_6512,N_6649);
xor U7480 (N_7480,N_6881,N_6550);
nand U7481 (N_7481,N_6659,N_6853);
xnor U7482 (N_7482,N_6150,N_6438);
and U7483 (N_7483,N_6816,N_6952);
nor U7484 (N_7484,N_6153,N_6951);
xnor U7485 (N_7485,N_6946,N_6671);
xnor U7486 (N_7486,N_6404,N_6759);
nor U7487 (N_7487,N_6019,N_6407);
nand U7488 (N_7488,N_6417,N_6845);
xor U7489 (N_7489,N_6850,N_6544);
and U7490 (N_7490,N_6679,N_6116);
xor U7491 (N_7491,N_6717,N_6039);
or U7492 (N_7492,N_6502,N_6563);
nand U7493 (N_7493,N_6196,N_6894);
nor U7494 (N_7494,N_6029,N_6250);
nand U7495 (N_7495,N_6870,N_6349);
xor U7496 (N_7496,N_6949,N_6058);
or U7497 (N_7497,N_6789,N_6411);
and U7498 (N_7498,N_6598,N_6602);
and U7499 (N_7499,N_6253,N_6737);
or U7500 (N_7500,N_6640,N_6954);
nand U7501 (N_7501,N_6201,N_6659);
nor U7502 (N_7502,N_6398,N_6824);
xor U7503 (N_7503,N_6580,N_6309);
xor U7504 (N_7504,N_6811,N_6477);
nand U7505 (N_7505,N_6181,N_6732);
nand U7506 (N_7506,N_6291,N_6121);
nand U7507 (N_7507,N_6120,N_6443);
nand U7508 (N_7508,N_6662,N_6436);
nor U7509 (N_7509,N_6169,N_6160);
xnor U7510 (N_7510,N_6828,N_6523);
xor U7511 (N_7511,N_6853,N_6794);
nor U7512 (N_7512,N_6324,N_6744);
nor U7513 (N_7513,N_6677,N_6220);
nor U7514 (N_7514,N_6477,N_6422);
or U7515 (N_7515,N_6267,N_6545);
nand U7516 (N_7516,N_6212,N_6529);
nor U7517 (N_7517,N_6333,N_6980);
nand U7518 (N_7518,N_6446,N_6500);
nor U7519 (N_7519,N_6129,N_6050);
xor U7520 (N_7520,N_6170,N_6589);
xnor U7521 (N_7521,N_6002,N_6839);
nand U7522 (N_7522,N_6674,N_6819);
and U7523 (N_7523,N_6560,N_6947);
nor U7524 (N_7524,N_6254,N_6296);
nand U7525 (N_7525,N_6685,N_6729);
nor U7526 (N_7526,N_6205,N_6538);
xnor U7527 (N_7527,N_6803,N_6878);
and U7528 (N_7528,N_6910,N_6707);
nand U7529 (N_7529,N_6284,N_6356);
and U7530 (N_7530,N_6207,N_6162);
or U7531 (N_7531,N_6694,N_6808);
and U7532 (N_7532,N_6230,N_6897);
and U7533 (N_7533,N_6593,N_6178);
xnor U7534 (N_7534,N_6505,N_6586);
nor U7535 (N_7535,N_6752,N_6558);
nand U7536 (N_7536,N_6122,N_6328);
or U7537 (N_7537,N_6958,N_6186);
nand U7538 (N_7538,N_6666,N_6754);
nand U7539 (N_7539,N_6996,N_6731);
xor U7540 (N_7540,N_6867,N_6653);
nand U7541 (N_7541,N_6060,N_6131);
nand U7542 (N_7542,N_6093,N_6632);
and U7543 (N_7543,N_6529,N_6981);
xnor U7544 (N_7544,N_6529,N_6016);
nor U7545 (N_7545,N_6872,N_6597);
xor U7546 (N_7546,N_6466,N_6560);
nand U7547 (N_7547,N_6767,N_6604);
and U7548 (N_7548,N_6224,N_6078);
nand U7549 (N_7549,N_6265,N_6807);
xnor U7550 (N_7550,N_6114,N_6686);
and U7551 (N_7551,N_6615,N_6058);
or U7552 (N_7552,N_6526,N_6802);
nor U7553 (N_7553,N_6772,N_6713);
nor U7554 (N_7554,N_6992,N_6921);
nor U7555 (N_7555,N_6283,N_6118);
or U7556 (N_7556,N_6736,N_6157);
nor U7557 (N_7557,N_6044,N_6509);
nand U7558 (N_7558,N_6451,N_6746);
nand U7559 (N_7559,N_6686,N_6396);
nor U7560 (N_7560,N_6843,N_6787);
or U7561 (N_7561,N_6057,N_6507);
or U7562 (N_7562,N_6267,N_6110);
or U7563 (N_7563,N_6804,N_6676);
and U7564 (N_7564,N_6428,N_6108);
xor U7565 (N_7565,N_6229,N_6367);
nor U7566 (N_7566,N_6082,N_6598);
xor U7567 (N_7567,N_6439,N_6522);
xor U7568 (N_7568,N_6542,N_6921);
nand U7569 (N_7569,N_6937,N_6014);
or U7570 (N_7570,N_6744,N_6376);
nand U7571 (N_7571,N_6001,N_6193);
nand U7572 (N_7572,N_6161,N_6305);
nand U7573 (N_7573,N_6488,N_6999);
xnor U7574 (N_7574,N_6336,N_6167);
nor U7575 (N_7575,N_6630,N_6721);
or U7576 (N_7576,N_6201,N_6457);
nor U7577 (N_7577,N_6781,N_6609);
nor U7578 (N_7578,N_6772,N_6283);
and U7579 (N_7579,N_6650,N_6752);
nor U7580 (N_7580,N_6440,N_6638);
or U7581 (N_7581,N_6352,N_6099);
and U7582 (N_7582,N_6745,N_6407);
nor U7583 (N_7583,N_6312,N_6087);
or U7584 (N_7584,N_6632,N_6265);
nor U7585 (N_7585,N_6400,N_6643);
nor U7586 (N_7586,N_6038,N_6992);
and U7587 (N_7587,N_6568,N_6877);
or U7588 (N_7588,N_6352,N_6072);
and U7589 (N_7589,N_6915,N_6373);
and U7590 (N_7590,N_6519,N_6597);
nand U7591 (N_7591,N_6868,N_6736);
or U7592 (N_7592,N_6588,N_6064);
nand U7593 (N_7593,N_6919,N_6178);
xor U7594 (N_7594,N_6357,N_6771);
nor U7595 (N_7595,N_6893,N_6842);
nor U7596 (N_7596,N_6556,N_6193);
xnor U7597 (N_7597,N_6679,N_6563);
and U7598 (N_7598,N_6069,N_6784);
nor U7599 (N_7599,N_6915,N_6935);
and U7600 (N_7600,N_6270,N_6392);
xnor U7601 (N_7601,N_6296,N_6760);
or U7602 (N_7602,N_6609,N_6439);
nor U7603 (N_7603,N_6945,N_6452);
nand U7604 (N_7604,N_6947,N_6239);
xnor U7605 (N_7605,N_6758,N_6997);
and U7606 (N_7606,N_6702,N_6066);
and U7607 (N_7607,N_6099,N_6406);
nor U7608 (N_7608,N_6462,N_6212);
nor U7609 (N_7609,N_6076,N_6311);
and U7610 (N_7610,N_6251,N_6275);
nand U7611 (N_7611,N_6941,N_6824);
or U7612 (N_7612,N_6633,N_6447);
and U7613 (N_7613,N_6305,N_6683);
xnor U7614 (N_7614,N_6907,N_6716);
nor U7615 (N_7615,N_6174,N_6239);
nand U7616 (N_7616,N_6942,N_6268);
nor U7617 (N_7617,N_6300,N_6602);
nand U7618 (N_7618,N_6733,N_6323);
nor U7619 (N_7619,N_6842,N_6302);
nor U7620 (N_7620,N_6726,N_6970);
xnor U7621 (N_7621,N_6919,N_6346);
nor U7622 (N_7622,N_6535,N_6994);
and U7623 (N_7623,N_6522,N_6036);
xnor U7624 (N_7624,N_6237,N_6421);
or U7625 (N_7625,N_6751,N_6953);
nor U7626 (N_7626,N_6931,N_6835);
and U7627 (N_7627,N_6447,N_6557);
and U7628 (N_7628,N_6905,N_6153);
xor U7629 (N_7629,N_6349,N_6358);
nor U7630 (N_7630,N_6380,N_6764);
nand U7631 (N_7631,N_6216,N_6669);
nor U7632 (N_7632,N_6496,N_6528);
xor U7633 (N_7633,N_6235,N_6681);
nand U7634 (N_7634,N_6738,N_6958);
nor U7635 (N_7635,N_6480,N_6056);
nand U7636 (N_7636,N_6141,N_6518);
xor U7637 (N_7637,N_6861,N_6847);
and U7638 (N_7638,N_6448,N_6775);
xnor U7639 (N_7639,N_6689,N_6224);
nand U7640 (N_7640,N_6167,N_6161);
and U7641 (N_7641,N_6460,N_6737);
xnor U7642 (N_7642,N_6788,N_6335);
or U7643 (N_7643,N_6342,N_6389);
nand U7644 (N_7644,N_6258,N_6328);
xor U7645 (N_7645,N_6523,N_6162);
nor U7646 (N_7646,N_6922,N_6596);
nand U7647 (N_7647,N_6794,N_6793);
or U7648 (N_7648,N_6374,N_6444);
or U7649 (N_7649,N_6525,N_6683);
xnor U7650 (N_7650,N_6058,N_6497);
xor U7651 (N_7651,N_6004,N_6297);
nor U7652 (N_7652,N_6099,N_6120);
or U7653 (N_7653,N_6456,N_6491);
nand U7654 (N_7654,N_6475,N_6769);
xnor U7655 (N_7655,N_6179,N_6228);
or U7656 (N_7656,N_6400,N_6545);
and U7657 (N_7657,N_6046,N_6021);
xor U7658 (N_7658,N_6584,N_6345);
nand U7659 (N_7659,N_6027,N_6434);
and U7660 (N_7660,N_6837,N_6842);
and U7661 (N_7661,N_6840,N_6317);
nand U7662 (N_7662,N_6749,N_6046);
nor U7663 (N_7663,N_6828,N_6755);
and U7664 (N_7664,N_6366,N_6812);
or U7665 (N_7665,N_6696,N_6967);
or U7666 (N_7666,N_6771,N_6197);
or U7667 (N_7667,N_6238,N_6467);
and U7668 (N_7668,N_6268,N_6622);
xnor U7669 (N_7669,N_6048,N_6488);
nor U7670 (N_7670,N_6334,N_6871);
nor U7671 (N_7671,N_6796,N_6407);
and U7672 (N_7672,N_6099,N_6423);
nand U7673 (N_7673,N_6200,N_6361);
or U7674 (N_7674,N_6360,N_6715);
nor U7675 (N_7675,N_6681,N_6690);
and U7676 (N_7676,N_6433,N_6654);
xnor U7677 (N_7677,N_6049,N_6230);
nand U7678 (N_7678,N_6015,N_6489);
nand U7679 (N_7679,N_6229,N_6216);
and U7680 (N_7680,N_6009,N_6232);
nor U7681 (N_7681,N_6579,N_6210);
nor U7682 (N_7682,N_6437,N_6529);
and U7683 (N_7683,N_6685,N_6931);
xnor U7684 (N_7684,N_6712,N_6890);
or U7685 (N_7685,N_6407,N_6841);
nor U7686 (N_7686,N_6170,N_6130);
or U7687 (N_7687,N_6117,N_6780);
nand U7688 (N_7688,N_6557,N_6067);
xor U7689 (N_7689,N_6470,N_6582);
or U7690 (N_7690,N_6806,N_6787);
nand U7691 (N_7691,N_6324,N_6062);
nand U7692 (N_7692,N_6861,N_6100);
or U7693 (N_7693,N_6698,N_6012);
xnor U7694 (N_7694,N_6065,N_6123);
xnor U7695 (N_7695,N_6318,N_6148);
xor U7696 (N_7696,N_6189,N_6735);
or U7697 (N_7697,N_6916,N_6855);
xor U7698 (N_7698,N_6346,N_6751);
nand U7699 (N_7699,N_6960,N_6783);
nor U7700 (N_7700,N_6553,N_6076);
xnor U7701 (N_7701,N_6353,N_6199);
and U7702 (N_7702,N_6791,N_6278);
and U7703 (N_7703,N_6773,N_6346);
and U7704 (N_7704,N_6342,N_6999);
nor U7705 (N_7705,N_6285,N_6961);
and U7706 (N_7706,N_6398,N_6617);
or U7707 (N_7707,N_6298,N_6646);
and U7708 (N_7708,N_6406,N_6230);
xnor U7709 (N_7709,N_6487,N_6566);
xor U7710 (N_7710,N_6099,N_6542);
nand U7711 (N_7711,N_6653,N_6931);
and U7712 (N_7712,N_6010,N_6342);
nor U7713 (N_7713,N_6564,N_6845);
xnor U7714 (N_7714,N_6326,N_6576);
nand U7715 (N_7715,N_6164,N_6117);
nand U7716 (N_7716,N_6706,N_6165);
and U7717 (N_7717,N_6960,N_6114);
nor U7718 (N_7718,N_6447,N_6602);
xnor U7719 (N_7719,N_6706,N_6977);
and U7720 (N_7720,N_6356,N_6383);
xor U7721 (N_7721,N_6945,N_6644);
xor U7722 (N_7722,N_6717,N_6321);
and U7723 (N_7723,N_6662,N_6415);
or U7724 (N_7724,N_6501,N_6263);
xnor U7725 (N_7725,N_6729,N_6574);
nand U7726 (N_7726,N_6630,N_6280);
or U7727 (N_7727,N_6264,N_6269);
nand U7728 (N_7728,N_6529,N_6587);
and U7729 (N_7729,N_6050,N_6170);
and U7730 (N_7730,N_6547,N_6921);
nor U7731 (N_7731,N_6870,N_6018);
nor U7732 (N_7732,N_6368,N_6831);
or U7733 (N_7733,N_6839,N_6118);
xnor U7734 (N_7734,N_6549,N_6761);
or U7735 (N_7735,N_6353,N_6771);
or U7736 (N_7736,N_6499,N_6299);
and U7737 (N_7737,N_6325,N_6103);
xor U7738 (N_7738,N_6025,N_6985);
nand U7739 (N_7739,N_6713,N_6092);
xnor U7740 (N_7740,N_6149,N_6200);
nor U7741 (N_7741,N_6948,N_6063);
or U7742 (N_7742,N_6014,N_6935);
nor U7743 (N_7743,N_6088,N_6575);
nand U7744 (N_7744,N_6049,N_6420);
or U7745 (N_7745,N_6209,N_6143);
xor U7746 (N_7746,N_6738,N_6140);
nor U7747 (N_7747,N_6404,N_6901);
and U7748 (N_7748,N_6740,N_6677);
nor U7749 (N_7749,N_6647,N_6017);
and U7750 (N_7750,N_6781,N_6300);
nand U7751 (N_7751,N_6987,N_6525);
nor U7752 (N_7752,N_6179,N_6277);
nor U7753 (N_7753,N_6456,N_6000);
and U7754 (N_7754,N_6133,N_6347);
nor U7755 (N_7755,N_6831,N_6058);
xnor U7756 (N_7756,N_6896,N_6206);
nor U7757 (N_7757,N_6525,N_6978);
xnor U7758 (N_7758,N_6272,N_6451);
nand U7759 (N_7759,N_6042,N_6182);
nor U7760 (N_7760,N_6927,N_6836);
nand U7761 (N_7761,N_6427,N_6295);
and U7762 (N_7762,N_6218,N_6946);
nand U7763 (N_7763,N_6963,N_6475);
nand U7764 (N_7764,N_6168,N_6615);
or U7765 (N_7765,N_6610,N_6718);
or U7766 (N_7766,N_6326,N_6211);
nand U7767 (N_7767,N_6189,N_6159);
nor U7768 (N_7768,N_6784,N_6880);
nor U7769 (N_7769,N_6895,N_6803);
xor U7770 (N_7770,N_6256,N_6724);
xnor U7771 (N_7771,N_6931,N_6807);
or U7772 (N_7772,N_6521,N_6320);
nor U7773 (N_7773,N_6655,N_6056);
nand U7774 (N_7774,N_6205,N_6264);
nor U7775 (N_7775,N_6348,N_6819);
or U7776 (N_7776,N_6035,N_6417);
nand U7777 (N_7777,N_6105,N_6036);
xnor U7778 (N_7778,N_6524,N_6150);
nand U7779 (N_7779,N_6611,N_6796);
or U7780 (N_7780,N_6247,N_6191);
nor U7781 (N_7781,N_6167,N_6013);
nor U7782 (N_7782,N_6230,N_6626);
nor U7783 (N_7783,N_6919,N_6883);
nand U7784 (N_7784,N_6586,N_6129);
nand U7785 (N_7785,N_6528,N_6357);
xor U7786 (N_7786,N_6791,N_6046);
xor U7787 (N_7787,N_6322,N_6469);
nor U7788 (N_7788,N_6575,N_6470);
nand U7789 (N_7789,N_6228,N_6590);
and U7790 (N_7790,N_6509,N_6016);
nand U7791 (N_7791,N_6908,N_6795);
and U7792 (N_7792,N_6696,N_6603);
nor U7793 (N_7793,N_6217,N_6753);
or U7794 (N_7794,N_6922,N_6640);
or U7795 (N_7795,N_6190,N_6374);
nor U7796 (N_7796,N_6238,N_6012);
nor U7797 (N_7797,N_6699,N_6851);
nor U7798 (N_7798,N_6583,N_6811);
and U7799 (N_7799,N_6258,N_6185);
nand U7800 (N_7800,N_6686,N_6647);
nand U7801 (N_7801,N_6514,N_6080);
or U7802 (N_7802,N_6993,N_6288);
or U7803 (N_7803,N_6366,N_6633);
or U7804 (N_7804,N_6630,N_6285);
nor U7805 (N_7805,N_6866,N_6679);
xor U7806 (N_7806,N_6184,N_6791);
xor U7807 (N_7807,N_6760,N_6213);
xnor U7808 (N_7808,N_6613,N_6037);
nand U7809 (N_7809,N_6065,N_6619);
or U7810 (N_7810,N_6317,N_6949);
nand U7811 (N_7811,N_6846,N_6644);
or U7812 (N_7812,N_6003,N_6586);
nand U7813 (N_7813,N_6152,N_6036);
nand U7814 (N_7814,N_6932,N_6962);
or U7815 (N_7815,N_6057,N_6493);
xor U7816 (N_7816,N_6299,N_6850);
or U7817 (N_7817,N_6457,N_6014);
nor U7818 (N_7818,N_6451,N_6656);
and U7819 (N_7819,N_6379,N_6789);
xnor U7820 (N_7820,N_6499,N_6177);
nor U7821 (N_7821,N_6946,N_6040);
nor U7822 (N_7822,N_6630,N_6535);
xnor U7823 (N_7823,N_6172,N_6449);
nor U7824 (N_7824,N_6992,N_6941);
or U7825 (N_7825,N_6625,N_6638);
nor U7826 (N_7826,N_6914,N_6152);
nor U7827 (N_7827,N_6330,N_6097);
or U7828 (N_7828,N_6393,N_6927);
and U7829 (N_7829,N_6023,N_6976);
nor U7830 (N_7830,N_6905,N_6603);
nand U7831 (N_7831,N_6405,N_6661);
nor U7832 (N_7832,N_6152,N_6716);
and U7833 (N_7833,N_6950,N_6164);
nor U7834 (N_7834,N_6190,N_6088);
nor U7835 (N_7835,N_6643,N_6231);
or U7836 (N_7836,N_6799,N_6879);
xnor U7837 (N_7837,N_6701,N_6318);
nand U7838 (N_7838,N_6499,N_6139);
xor U7839 (N_7839,N_6466,N_6357);
and U7840 (N_7840,N_6787,N_6943);
xor U7841 (N_7841,N_6751,N_6301);
xnor U7842 (N_7842,N_6351,N_6593);
xnor U7843 (N_7843,N_6433,N_6347);
xnor U7844 (N_7844,N_6136,N_6374);
nor U7845 (N_7845,N_6221,N_6735);
nand U7846 (N_7846,N_6562,N_6841);
xor U7847 (N_7847,N_6895,N_6075);
or U7848 (N_7848,N_6514,N_6983);
nand U7849 (N_7849,N_6965,N_6486);
nor U7850 (N_7850,N_6385,N_6630);
nand U7851 (N_7851,N_6402,N_6584);
and U7852 (N_7852,N_6647,N_6527);
nand U7853 (N_7853,N_6235,N_6455);
nor U7854 (N_7854,N_6104,N_6541);
or U7855 (N_7855,N_6253,N_6759);
xor U7856 (N_7856,N_6433,N_6382);
xnor U7857 (N_7857,N_6908,N_6738);
or U7858 (N_7858,N_6161,N_6002);
or U7859 (N_7859,N_6542,N_6426);
xnor U7860 (N_7860,N_6784,N_6230);
nor U7861 (N_7861,N_6285,N_6735);
and U7862 (N_7862,N_6579,N_6768);
and U7863 (N_7863,N_6924,N_6893);
xnor U7864 (N_7864,N_6748,N_6505);
nor U7865 (N_7865,N_6538,N_6270);
xnor U7866 (N_7866,N_6249,N_6884);
and U7867 (N_7867,N_6377,N_6315);
nor U7868 (N_7868,N_6775,N_6552);
xor U7869 (N_7869,N_6356,N_6233);
nor U7870 (N_7870,N_6647,N_6092);
nor U7871 (N_7871,N_6542,N_6927);
nor U7872 (N_7872,N_6973,N_6718);
and U7873 (N_7873,N_6508,N_6877);
nor U7874 (N_7874,N_6801,N_6984);
or U7875 (N_7875,N_6113,N_6688);
or U7876 (N_7876,N_6155,N_6995);
nor U7877 (N_7877,N_6486,N_6205);
or U7878 (N_7878,N_6546,N_6972);
nor U7879 (N_7879,N_6620,N_6628);
xnor U7880 (N_7880,N_6656,N_6618);
nand U7881 (N_7881,N_6197,N_6884);
or U7882 (N_7882,N_6700,N_6616);
nor U7883 (N_7883,N_6514,N_6838);
or U7884 (N_7884,N_6451,N_6916);
and U7885 (N_7885,N_6561,N_6180);
or U7886 (N_7886,N_6181,N_6621);
or U7887 (N_7887,N_6592,N_6096);
and U7888 (N_7888,N_6681,N_6221);
xor U7889 (N_7889,N_6966,N_6913);
nor U7890 (N_7890,N_6167,N_6311);
and U7891 (N_7891,N_6421,N_6269);
xor U7892 (N_7892,N_6900,N_6865);
nor U7893 (N_7893,N_6723,N_6798);
nor U7894 (N_7894,N_6000,N_6774);
and U7895 (N_7895,N_6815,N_6281);
nand U7896 (N_7896,N_6836,N_6040);
nor U7897 (N_7897,N_6126,N_6066);
or U7898 (N_7898,N_6302,N_6234);
xnor U7899 (N_7899,N_6441,N_6452);
xor U7900 (N_7900,N_6136,N_6154);
nand U7901 (N_7901,N_6829,N_6270);
xnor U7902 (N_7902,N_6338,N_6484);
or U7903 (N_7903,N_6217,N_6682);
nand U7904 (N_7904,N_6020,N_6805);
xor U7905 (N_7905,N_6567,N_6578);
nor U7906 (N_7906,N_6077,N_6252);
and U7907 (N_7907,N_6042,N_6717);
nor U7908 (N_7908,N_6209,N_6879);
nor U7909 (N_7909,N_6353,N_6117);
nand U7910 (N_7910,N_6650,N_6483);
xor U7911 (N_7911,N_6600,N_6515);
xor U7912 (N_7912,N_6161,N_6698);
nor U7913 (N_7913,N_6639,N_6879);
or U7914 (N_7914,N_6683,N_6955);
and U7915 (N_7915,N_6817,N_6435);
nand U7916 (N_7916,N_6672,N_6616);
nor U7917 (N_7917,N_6800,N_6178);
or U7918 (N_7918,N_6202,N_6424);
xor U7919 (N_7919,N_6199,N_6800);
or U7920 (N_7920,N_6144,N_6595);
or U7921 (N_7921,N_6391,N_6668);
or U7922 (N_7922,N_6448,N_6410);
nand U7923 (N_7923,N_6818,N_6753);
or U7924 (N_7924,N_6770,N_6308);
or U7925 (N_7925,N_6286,N_6529);
and U7926 (N_7926,N_6287,N_6391);
nor U7927 (N_7927,N_6432,N_6877);
or U7928 (N_7928,N_6081,N_6708);
nand U7929 (N_7929,N_6623,N_6133);
or U7930 (N_7930,N_6761,N_6578);
and U7931 (N_7931,N_6470,N_6765);
and U7932 (N_7932,N_6059,N_6179);
xnor U7933 (N_7933,N_6842,N_6722);
nand U7934 (N_7934,N_6550,N_6480);
nand U7935 (N_7935,N_6545,N_6404);
and U7936 (N_7936,N_6204,N_6911);
xor U7937 (N_7937,N_6718,N_6324);
nand U7938 (N_7938,N_6953,N_6411);
nand U7939 (N_7939,N_6909,N_6049);
xor U7940 (N_7940,N_6085,N_6544);
nand U7941 (N_7941,N_6445,N_6147);
nor U7942 (N_7942,N_6039,N_6613);
and U7943 (N_7943,N_6144,N_6992);
nor U7944 (N_7944,N_6345,N_6637);
xor U7945 (N_7945,N_6553,N_6265);
nand U7946 (N_7946,N_6287,N_6026);
and U7947 (N_7947,N_6217,N_6930);
xor U7948 (N_7948,N_6648,N_6109);
nand U7949 (N_7949,N_6802,N_6047);
nand U7950 (N_7950,N_6855,N_6483);
nand U7951 (N_7951,N_6990,N_6473);
or U7952 (N_7952,N_6771,N_6756);
xor U7953 (N_7953,N_6560,N_6502);
nor U7954 (N_7954,N_6203,N_6232);
or U7955 (N_7955,N_6722,N_6631);
and U7956 (N_7956,N_6309,N_6743);
xnor U7957 (N_7957,N_6647,N_6600);
nor U7958 (N_7958,N_6115,N_6711);
nor U7959 (N_7959,N_6220,N_6838);
nor U7960 (N_7960,N_6027,N_6609);
and U7961 (N_7961,N_6148,N_6590);
and U7962 (N_7962,N_6285,N_6754);
xor U7963 (N_7963,N_6722,N_6838);
nand U7964 (N_7964,N_6773,N_6968);
nand U7965 (N_7965,N_6335,N_6412);
or U7966 (N_7966,N_6461,N_6206);
xnor U7967 (N_7967,N_6344,N_6124);
xnor U7968 (N_7968,N_6154,N_6937);
nand U7969 (N_7969,N_6557,N_6820);
and U7970 (N_7970,N_6026,N_6535);
and U7971 (N_7971,N_6723,N_6909);
nor U7972 (N_7972,N_6564,N_6006);
and U7973 (N_7973,N_6040,N_6092);
and U7974 (N_7974,N_6437,N_6030);
xor U7975 (N_7975,N_6885,N_6188);
or U7976 (N_7976,N_6746,N_6596);
nand U7977 (N_7977,N_6917,N_6399);
nand U7978 (N_7978,N_6715,N_6861);
or U7979 (N_7979,N_6984,N_6915);
nor U7980 (N_7980,N_6658,N_6951);
or U7981 (N_7981,N_6214,N_6341);
nand U7982 (N_7982,N_6990,N_6804);
nor U7983 (N_7983,N_6448,N_6434);
xnor U7984 (N_7984,N_6313,N_6509);
or U7985 (N_7985,N_6798,N_6129);
nor U7986 (N_7986,N_6151,N_6232);
and U7987 (N_7987,N_6904,N_6344);
nand U7988 (N_7988,N_6243,N_6323);
and U7989 (N_7989,N_6192,N_6884);
nand U7990 (N_7990,N_6531,N_6157);
xnor U7991 (N_7991,N_6890,N_6657);
or U7992 (N_7992,N_6679,N_6029);
nand U7993 (N_7993,N_6139,N_6846);
xor U7994 (N_7994,N_6372,N_6486);
xor U7995 (N_7995,N_6036,N_6903);
nor U7996 (N_7996,N_6388,N_6905);
xor U7997 (N_7997,N_6855,N_6333);
xnor U7998 (N_7998,N_6985,N_6250);
xor U7999 (N_7999,N_6464,N_6683);
nand U8000 (N_8000,N_7737,N_7910);
or U8001 (N_8001,N_7818,N_7641);
or U8002 (N_8002,N_7928,N_7843);
nand U8003 (N_8003,N_7494,N_7350);
nor U8004 (N_8004,N_7044,N_7352);
and U8005 (N_8005,N_7619,N_7095);
nor U8006 (N_8006,N_7330,N_7835);
xnor U8007 (N_8007,N_7200,N_7883);
xnor U8008 (N_8008,N_7812,N_7823);
nor U8009 (N_8009,N_7216,N_7436);
or U8010 (N_8010,N_7639,N_7250);
xor U8011 (N_8011,N_7107,N_7672);
nand U8012 (N_8012,N_7713,N_7614);
nand U8013 (N_8013,N_7645,N_7132);
or U8014 (N_8014,N_7934,N_7886);
or U8015 (N_8015,N_7307,N_7926);
or U8016 (N_8016,N_7485,N_7417);
xnor U8017 (N_8017,N_7675,N_7163);
xnor U8018 (N_8018,N_7852,N_7535);
or U8019 (N_8019,N_7468,N_7961);
or U8020 (N_8020,N_7727,N_7210);
nor U8021 (N_8021,N_7997,N_7377);
and U8022 (N_8022,N_7915,N_7402);
xor U8023 (N_8023,N_7676,N_7253);
or U8024 (N_8024,N_7504,N_7702);
and U8025 (N_8025,N_7491,N_7159);
nand U8026 (N_8026,N_7257,N_7018);
xnor U8027 (N_8027,N_7596,N_7691);
xor U8028 (N_8028,N_7890,N_7325);
and U8029 (N_8029,N_7813,N_7597);
nor U8030 (N_8030,N_7828,N_7310);
xnor U8031 (N_8031,N_7769,N_7804);
nor U8032 (N_8032,N_7223,N_7233);
xor U8033 (N_8033,N_7892,N_7052);
and U8034 (N_8034,N_7924,N_7483);
xor U8035 (N_8035,N_7930,N_7488);
nand U8036 (N_8036,N_7746,N_7955);
nand U8037 (N_8037,N_7141,N_7005);
xor U8038 (N_8038,N_7879,N_7001);
or U8039 (N_8039,N_7004,N_7124);
nor U8040 (N_8040,N_7336,N_7887);
xor U8041 (N_8041,N_7166,N_7304);
xor U8042 (N_8042,N_7321,N_7602);
nand U8043 (N_8043,N_7161,N_7680);
nor U8044 (N_8044,N_7635,N_7416);
and U8045 (N_8045,N_7145,N_7134);
nor U8046 (N_8046,N_7882,N_7598);
nand U8047 (N_8047,N_7471,N_7326);
nand U8048 (N_8048,N_7220,N_7408);
nor U8049 (N_8049,N_7858,N_7857);
and U8050 (N_8050,N_7573,N_7207);
nand U8051 (N_8051,N_7411,N_7987);
or U8052 (N_8052,N_7293,N_7604);
and U8053 (N_8053,N_7829,N_7793);
nor U8054 (N_8054,N_7153,N_7372);
and U8055 (N_8055,N_7757,N_7654);
xor U8056 (N_8056,N_7825,N_7206);
nor U8057 (N_8057,N_7795,N_7611);
or U8058 (N_8058,N_7152,N_7148);
or U8059 (N_8059,N_7418,N_7292);
or U8060 (N_8060,N_7324,N_7996);
nor U8061 (N_8061,N_7923,N_7677);
xor U8062 (N_8062,N_7547,N_7553);
nand U8063 (N_8063,N_7301,N_7357);
nand U8064 (N_8064,N_7105,N_7659);
xor U8065 (N_8065,N_7985,N_7642);
nand U8066 (N_8066,N_7164,N_7264);
xnor U8067 (N_8067,N_7461,N_7601);
xnor U8068 (N_8068,N_7475,N_7388);
nand U8069 (N_8069,N_7067,N_7271);
and U8070 (N_8070,N_7782,N_7419);
nor U8071 (N_8071,N_7374,N_7640);
and U8072 (N_8072,N_7169,N_7306);
xor U8073 (N_8073,N_7329,N_7409);
xnor U8074 (N_8074,N_7748,N_7281);
xor U8075 (N_8075,N_7668,N_7221);
nand U8076 (N_8076,N_7120,N_7068);
and U8077 (N_8077,N_7239,N_7744);
and U8078 (N_8078,N_7734,N_7397);
xor U8079 (N_8079,N_7021,N_7690);
or U8080 (N_8080,N_7447,N_7730);
nand U8081 (N_8081,N_7122,N_7929);
xor U8082 (N_8082,N_7552,N_7123);
and U8083 (N_8083,N_7229,N_7781);
and U8084 (N_8084,N_7384,N_7541);
xor U8085 (N_8085,N_7248,N_7354);
nand U8086 (N_8086,N_7674,N_7809);
nand U8087 (N_8087,N_7722,N_7567);
nand U8088 (N_8088,N_7038,N_7231);
nor U8089 (N_8089,N_7341,N_7007);
and U8090 (N_8090,N_7988,N_7479);
or U8091 (N_8091,N_7342,N_7087);
xnor U8092 (N_8092,N_7884,N_7945);
nor U8093 (N_8093,N_7976,N_7845);
and U8094 (N_8094,N_7562,N_7867);
nand U8095 (N_8095,N_7158,N_7539);
and U8096 (N_8096,N_7951,N_7992);
xor U8097 (N_8097,N_7740,N_7735);
nor U8098 (N_8098,N_7392,N_7056);
xnor U8099 (N_8099,N_7282,N_7453);
and U8100 (N_8100,N_7527,N_7054);
and U8101 (N_8101,N_7034,N_7061);
nor U8102 (N_8102,N_7836,N_7308);
nand U8103 (N_8103,N_7362,N_7279);
nor U8104 (N_8104,N_7623,N_7580);
nand U8105 (N_8105,N_7941,N_7305);
xor U8106 (N_8106,N_7393,N_7978);
xor U8107 (N_8107,N_7710,N_7665);
and U8108 (N_8108,N_7142,N_7805);
nor U8109 (N_8109,N_7450,N_7331);
and U8110 (N_8110,N_7741,N_7186);
and U8111 (N_8111,N_7811,N_7643);
nor U8112 (N_8112,N_7509,N_7344);
or U8113 (N_8113,N_7517,N_7464);
and U8114 (N_8114,N_7266,N_7631);
nor U8115 (N_8115,N_7480,N_7252);
or U8116 (N_8116,N_7833,N_7270);
xnor U8117 (N_8117,N_7143,N_7222);
or U8118 (N_8118,N_7947,N_7489);
nor U8119 (N_8119,N_7522,N_7177);
and U8120 (N_8120,N_7856,N_7872);
nand U8121 (N_8121,N_7794,N_7669);
nor U8122 (N_8122,N_7888,N_7002);
nand U8123 (N_8123,N_7940,N_7942);
or U8124 (N_8124,N_7209,N_7360);
and U8125 (N_8125,N_7891,N_7082);
and U8126 (N_8126,N_7777,N_7014);
nand U8127 (N_8127,N_7628,N_7719);
and U8128 (N_8128,N_7606,N_7398);
nand U8129 (N_8129,N_7172,N_7484);
and U8130 (N_8130,N_7729,N_7455);
nor U8131 (N_8131,N_7295,N_7017);
or U8132 (N_8132,N_7822,N_7171);
and U8133 (N_8133,N_7118,N_7931);
nor U8134 (N_8134,N_7170,N_7065);
nor U8135 (N_8135,N_7759,N_7133);
nor U8136 (N_8136,N_7974,N_7587);
or U8137 (N_8137,N_7277,N_7303);
nand U8138 (N_8138,N_7898,N_7115);
xnor U8139 (N_8139,N_7981,N_7919);
nor U8140 (N_8140,N_7268,N_7078);
xor U8141 (N_8141,N_7138,N_7626);
xnor U8142 (N_8142,N_7911,N_7851);
nor U8143 (N_8143,N_7473,N_7050);
xor U8144 (N_8144,N_7554,N_7199);
nand U8145 (N_8145,N_7335,N_7294);
nand U8146 (N_8146,N_7678,N_7590);
nor U8147 (N_8147,N_7998,N_7874);
or U8148 (N_8148,N_7426,N_7055);
or U8149 (N_8149,N_7712,N_7663);
nand U8150 (N_8150,N_7525,N_7178);
nand U8151 (N_8151,N_7218,N_7693);
nor U8152 (N_8152,N_7391,N_7516);
or U8153 (N_8153,N_7476,N_7600);
nand U8154 (N_8154,N_7045,N_7470);
or U8155 (N_8155,N_7296,N_7816);
xor U8156 (N_8156,N_7185,N_7954);
xor U8157 (N_8157,N_7049,N_7842);
nand U8158 (N_8158,N_7815,N_7979);
xor U8159 (N_8159,N_7080,N_7400);
and U8160 (N_8160,N_7280,N_7456);
nand U8161 (N_8161,N_7093,N_7214);
nor U8162 (N_8162,N_7756,N_7071);
nand U8163 (N_8163,N_7237,N_7254);
nor U8164 (N_8164,N_7963,N_7658);
nand U8165 (N_8165,N_7916,N_7188);
xnor U8166 (N_8166,N_7708,N_7059);
nor U8167 (N_8167,N_7909,N_7104);
nand U8168 (N_8168,N_7984,N_7739);
or U8169 (N_8169,N_7644,N_7927);
nand U8170 (N_8170,N_7878,N_7512);
nand U8171 (N_8171,N_7555,N_7550);
xor U8172 (N_8172,N_7116,N_7260);
xnor U8173 (N_8173,N_7273,N_7181);
nor U8174 (N_8174,N_7810,N_7943);
or U8175 (N_8175,N_7462,N_7316);
nand U8176 (N_8176,N_7538,N_7047);
xnor U8177 (N_8177,N_7551,N_7238);
xnor U8178 (N_8178,N_7463,N_7956);
xnor U8179 (N_8179,N_7083,N_7610);
and U8180 (N_8180,N_7434,N_7820);
or U8181 (N_8181,N_7106,N_7340);
nand U8182 (N_8182,N_7807,N_7932);
or U8183 (N_8183,N_7784,N_7297);
and U8184 (N_8184,N_7351,N_7768);
xor U8185 (N_8185,N_7556,N_7053);
nand U8186 (N_8186,N_7236,N_7022);
nand U8187 (N_8187,N_7969,N_7037);
xnor U8188 (N_8188,N_7908,N_7399);
nand U8189 (N_8189,N_7276,N_7629);
nand U8190 (N_8190,N_7278,N_7515);
nor U8191 (N_8191,N_7286,N_7339);
nand U8192 (N_8192,N_7348,N_7994);
or U8193 (N_8193,N_7798,N_7745);
nor U8194 (N_8194,N_7896,N_7819);
nand U8195 (N_8195,N_7960,N_7315);
or U8196 (N_8196,N_7179,N_7195);
and U8197 (N_8197,N_7474,N_7460);
nand U8198 (N_8198,N_7009,N_7786);
xor U8199 (N_8199,N_7318,N_7492);
or U8200 (N_8200,N_7760,N_7285);
nor U8201 (N_8201,N_7424,N_7086);
nor U8202 (N_8202,N_7761,N_7300);
xor U8203 (N_8203,N_7160,N_7689);
or U8204 (N_8204,N_7466,N_7935);
or U8205 (N_8205,N_7799,N_7103);
or U8206 (N_8206,N_7752,N_7211);
and U8207 (N_8207,N_7792,N_7897);
xnor U8208 (N_8208,N_7019,N_7048);
nand U8209 (N_8209,N_7032,N_7187);
xnor U8210 (N_8210,N_7043,N_7309);
xor U8211 (N_8211,N_7472,N_7648);
nor U8212 (N_8212,N_7989,N_7905);
xor U8213 (N_8213,N_7383,N_7767);
nor U8214 (N_8214,N_7420,N_7803);
xor U8215 (N_8215,N_7202,N_7684);
nor U8216 (N_8216,N_7208,N_7006);
xnor U8217 (N_8217,N_7111,N_7345);
or U8218 (N_8218,N_7182,N_7151);
nor U8219 (N_8219,N_7778,N_7228);
nand U8220 (N_8220,N_7859,N_7312);
xor U8221 (N_8221,N_7736,N_7251);
xor U8222 (N_8222,N_7594,N_7687);
and U8223 (N_8223,N_7502,N_7565);
or U8224 (N_8224,N_7196,N_7521);
nor U8225 (N_8225,N_7881,N_7999);
and U8226 (N_8226,N_7622,N_7421);
or U8227 (N_8227,N_7333,N_7081);
nor U8228 (N_8228,N_7946,N_7201);
xnor U8229 (N_8229,N_7670,N_7013);
and U8230 (N_8230,N_7557,N_7526);
nor U8231 (N_8231,N_7094,N_7718);
or U8232 (N_8232,N_7993,N_7405);
and U8233 (N_8233,N_7838,N_7854);
nor U8234 (N_8234,N_7742,N_7849);
or U8235 (N_8235,N_7267,N_7030);
nor U8236 (N_8236,N_7853,N_7477);
nand U8237 (N_8237,N_7386,N_7832);
nand U8238 (N_8238,N_7288,N_7518);
and U8239 (N_8239,N_7790,N_7395);
and U8240 (N_8240,N_7366,N_7682);
nor U8241 (N_8241,N_7764,N_7334);
nor U8242 (N_8242,N_7057,N_7564);
xor U8243 (N_8243,N_7291,N_7673);
nor U8244 (N_8244,N_7226,N_7242);
nor U8245 (N_8245,N_7438,N_7039);
and U8246 (N_8246,N_7481,N_7800);
or U8247 (N_8247,N_7871,N_7532);
nor U8248 (N_8248,N_7099,N_7848);
nor U8249 (N_8249,N_7446,N_7802);
or U8250 (N_8250,N_7519,N_7412);
nand U8251 (N_8251,N_7637,N_7983);
xnor U8252 (N_8252,N_7575,N_7724);
xnor U8253 (N_8253,N_7040,N_7119);
and U8254 (N_8254,N_7721,N_7363);
nor U8255 (N_8255,N_7826,N_7130);
or U8256 (N_8256,N_7902,N_7632);
xnor U8257 (N_8257,N_7443,N_7454);
or U8258 (N_8258,N_7112,N_7382);
and U8259 (N_8259,N_7387,N_7096);
xor U8260 (N_8260,N_7146,N_7574);
or U8261 (N_8261,N_7824,N_7868);
and U8262 (N_8262,N_7486,N_7789);
or U8263 (N_8263,N_7865,N_7660);
and U8264 (N_8264,N_7197,N_7776);
and U8265 (N_8265,N_7364,N_7864);
xnor U8266 (N_8266,N_7085,N_7577);
nand U8267 (N_8267,N_7369,N_7566);
xor U8268 (N_8268,N_7709,N_7404);
or U8269 (N_8269,N_7679,N_7968);
nand U8270 (N_8270,N_7970,N_7375);
nor U8271 (N_8271,N_7174,N_7413);
and U8272 (N_8272,N_7389,N_7863);
nor U8273 (N_8273,N_7010,N_7558);
and U8274 (N_8274,N_7311,N_7064);
nand U8275 (N_8275,N_7072,N_7332);
xnor U8276 (N_8276,N_7102,N_7568);
and U8277 (N_8277,N_7584,N_7284);
and U8278 (N_8278,N_7618,N_7136);
nor U8279 (N_8279,N_7579,N_7088);
nor U8280 (N_8280,N_7731,N_7150);
and U8281 (N_8281,N_7203,N_7542);
nand U8282 (N_8282,N_7060,N_7771);
nand U8283 (N_8283,N_7075,N_7227);
nand U8284 (N_8284,N_7011,N_7507);
nand U8285 (N_8285,N_7320,N_7873);
nor U8286 (N_8286,N_7036,N_7847);
nor U8287 (N_8287,N_7026,N_7696);
and U8288 (N_8288,N_7452,N_7796);
nand U8289 (N_8289,N_7529,N_7378);
xor U8290 (N_8290,N_7023,N_7487);
nand U8291 (N_8291,N_7243,N_7633);
xor U8292 (N_8292,N_7763,N_7936);
xor U8293 (N_8293,N_7885,N_7814);
nor U8294 (N_8294,N_7298,N_7385);
or U8295 (N_8295,N_7900,N_7355);
and U8296 (N_8296,N_7358,N_7493);
nand U8297 (N_8297,N_7613,N_7063);
and U8298 (N_8298,N_7431,N_7949);
xnor U8299 (N_8299,N_7025,N_7995);
nand U8300 (N_8300,N_7770,N_7499);
or U8301 (N_8301,N_7346,N_7373);
and U8302 (N_8302,N_7563,N_7451);
and U8303 (N_8303,N_7356,N_7918);
or U8304 (N_8304,N_7168,N_7437);
xnor U8305 (N_8305,N_7272,N_7365);
nand U8306 (N_8306,N_7962,N_7540);
xor U8307 (N_8307,N_7184,N_7167);
and U8308 (N_8308,N_7445,N_7194);
or U8309 (N_8309,N_7508,N_7189);
xor U8310 (N_8310,N_7390,N_7097);
nand U8311 (N_8311,N_7583,N_7559);
and U8312 (N_8312,N_7965,N_7531);
nor U8313 (N_8313,N_7840,N_7754);
and U8314 (N_8314,N_7113,N_7703);
xnor U8315 (N_8315,N_7681,N_7046);
and U8316 (N_8316,N_7062,N_7302);
and U8317 (N_8317,N_7975,N_7662);
nor U8318 (N_8318,N_7255,N_7371);
nand U8319 (N_8319,N_7287,N_7175);
xnor U8320 (N_8320,N_7091,N_7035);
nand U8321 (N_8321,N_7860,N_7593);
nor U8322 (N_8322,N_7544,N_7647);
xor U8323 (N_8323,N_7704,N_7353);
and U8324 (N_8324,N_7073,N_7198);
and U8325 (N_8325,N_7520,N_7127);
or U8326 (N_8326,N_7008,N_7449);
xor U8327 (N_8327,N_7459,N_7808);
xor U8328 (N_8328,N_7139,N_7821);
xor U8329 (N_8329,N_7801,N_7000);
xor U8330 (N_8330,N_7290,N_7367);
xor U8331 (N_8331,N_7543,N_7289);
xor U8332 (N_8332,N_7560,N_7627);
nor U8333 (N_8333,N_7785,N_7343);
xor U8334 (N_8334,N_7876,N_7850);
and U8335 (N_8335,N_7889,N_7429);
and U8336 (N_8336,N_7548,N_7991);
nand U8337 (N_8337,N_7726,N_7621);
xnor U8338 (N_8338,N_7505,N_7572);
or U8339 (N_8339,N_7234,N_7396);
and U8340 (N_8340,N_7215,N_7204);
or U8341 (N_8341,N_7368,N_7578);
nor U8342 (N_8342,N_7755,N_7448);
or U8343 (N_8343,N_7317,N_7683);
nand U8344 (N_8344,N_7249,N_7031);
nand U8345 (N_8345,N_7089,N_7074);
xnor U8346 (N_8346,N_7925,N_7866);
or U8347 (N_8347,N_7381,N_7765);
and U8348 (N_8348,N_7422,N_7137);
xnor U8349 (N_8349,N_7880,N_7894);
nor U8350 (N_8350,N_7114,N_7612);
xnor U8351 (N_8351,N_7269,N_7967);
and U8352 (N_8352,N_7615,N_7523);
or U8353 (N_8353,N_7183,N_7775);
xnor U8354 (N_8354,N_7066,N_7588);
and U8355 (N_8355,N_7435,N_7723);
nand U8356 (N_8356,N_7265,N_7176);
or U8357 (N_8357,N_7585,N_7700);
or U8358 (N_8358,N_7904,N_7439);
and U8359 (N_8359,N_7140,N_7753);
and U8360 (N_8360,N_7938,N_7939);
nand U8361 (N_8361,N_7686,N_7241);
nand U8362 (N_8362,N_7192,N_7444);
nor U8363 (N_8363,N_7698,N_7870);
xor U8364 (N_8364,N_7920,N_7869);
or U8365 (N_8365,N_7569,N_7666);
or U8366 (N_8366,N_7831,N_7797);
nand U8367 (N_8367,N_7787,N_7503);
and U8368 (N_8368,N_7156,N_7749);
nand U8369 (N_8369,N_7609,N_7501);
and U8370 (N_8370,N_7070,N_7977);
xor U8371 (N_8371,N_7617,N_7616);
xor U8372 (N_8372,N_7497,N_7256);
or U8373 (N_8373,N_7469,N_7425);
nor U8374 (N_8374,N_7359,N_7135);
nor U8375 (N_8375,N_7570,N_7524);
nor U8376 (N_8376,N_7990,N_7240);
nor U8377 (N_8377,N_7651,N_7478);
nor U8378 (N_8378,N_7245,N_7957);
nand U8379 (N_8379,N_7457,N_7766);
xnor U8380 (N_8380,N_7982,N_7440);
or U8381 (N_8381,N_7958,N_7003);
nand U8382 (N_8382,N_7084,N_7762);
nand U8383 (N_8383,N_7155,N_7774);
xnor U8384 (N_8384,N_7685,N_7545);
or U8385 (N_8385,N_7692,N_7079);
xnor U8386 (N_8386,N_7027,N_7129);
and U8387 (N_8387,N_7128,N_7537);
or U8388 (N_8388,N_7758,N_7661);
xnor U8389 (N_8389,N_7607,N_7534);
or U8390 (N_8390,N_7733,N_7834);
xnor U8391 (N_8391,N_7728,N_7069);
nor U8392 (N_8392,N_7791,N_7020);
or U8393 (N_8393,N_7263,N_7899);
nor U8394 (N_8394,N_7376,N_7817);
or U8395 (N_8395,N_7205,N_7903);
or U8396 (N_8396,N_7608,N_7714);
xor U8397 (N_8397,N_7656,N_7495);
nor U8398 (N_8398,N_7953,N_7980);
nand U8399 (N_8399,N_7513,N_7780);
and U8400 (N_8400,N_7028,N_7401);
nor U8401 (N_8401,N_7012,N_7051);
xnor U8402 (N_8402,N_7015,N_7147);
nor U8403 (N_8403,N_7349,N_7699);
xnor U8404 (N_8404,N_7090,N_7971);
and U8405 (N_8405,N_7844,N_7788);
and U8406 (N_8406,N_7948,N_7620);
nand U8407 (N_8407,N_7506,N_7646);
nor U8408 (N_8408,N_7695,N_7423);
or U8409 (N_8409,N_7952,N_7694);
nand U8410 (N_8410,N_7624,N_7299);
nand U8411 (N_8411,N_7536,N_7514);
nor U8412 (N_8412,N_7747,N_7193);
and U8413 (N_8413,N_7922,N_7595);
nor U8414 (N_8414,N_7110,N_7907);
nand U8415 (N_8415,N_7592,N_7258);
and U8416 (N_8416,N_7750,N_7986);
and U8417 (N_8417,N_7126,N_7893);
xor U8418 (N_8418,N_7259,N_7649);
or U8419 (N_8419,N_7244,N_7846);
and U8420 (N_8420,N_7246,N_7275);
nor U8421 (N_8421,N_7274,N_7964);
nand U8422 (N_8422,N_7561,N_7743);
nor U8423 (N_8423,N_7033,N_7906);
and U8424 (N_8424,N_7715,N_7191);
nor U8425 (N_8425,N_7839,N_7261);
xnor U8426 (N_8426,N_7530,N_7433);
and U8427 (N_8427,N_7546,N_7427);
and U8428 (N_8428,N_7338,N_7830);
nand U8429 (N_8429,N_7157,N_7973);
nor U8430 (N_8430,N_7041,N_7212);
or U8431 (N_8431,N_7664,N_7586);
xor U8432 (N_8432,N_7467,N_7313);
nand U8433 (N_8433,N_7162,N_7630);
nand U8434 (N_8434,N_7652,N_7458);
nand U8435 (N_8435,N_7582,N_7430);
or U8436 (N_8436,N_7862,N_7328);
nand U8437 (N_8437,N_7914,N_7283);
xor U8438 (N_8438,N_7589,N_7190);
or U8439 (N_8439,N_7549,N_7861);
and U8440 (N_8440,N_7125,N_7603);
or U8441 (N_8441,N_7653,N_7533);
nor U8442 (N_8442,N_7732,N_7751);
nor U8443 (N_8443,N_7496,N_7707);
and U8444 (N_8444,N_7855,N_7465);
nand U8445 (N_8445,N_7414,N_7441);
and U8446 (N_8446,N_7576,N_7720);
nor U8447 (N_8447,N_7841,N_7432);
and U8448 (N_8448,N_7901,N_7235);
or U8449 (N_8449,N_7108,N_7117);
or U8450 (N_8450,N_7837,N_7109);
and U8451 (N_8451,N_7697,N_7688);
or U8452 (N_8452,N_7029,N_7092);
nand U8453 (N_8453,N_7428,N_7511);
xor U8454 (N_8454,N_7042,N_7605);
nand U8455 (N_8455,N_7394,N_7717);
nand U8456 (N_8456,N_7482,N_7917);
nor U8457 (N_8457,N_7772,N_7370);
or U8458 (N_8458,N_7706,N_7406);
nand U8459 (N_8459,N_7403,N_7410);
nor U8460 (N_8460,N_7650,N_7154);
xor U8461 (N_8461,N_7327,N_7076);
xnor U8462 (N_8462,N_7219,N_7667);
or U8463 (N_8463,N_7528,N_7407);
or U8464 (N_8464,N_7959,N_7230);
xor U8465 (N_8465,N_7173,N_7016);
nand U8466 (N_8466,N_7725,N_7131);
nand U8467 (N_8467,N_7716,N_7950);
nor U8468 (N_8468,N_7972,N_7912);
xnor U8469 (N_8469,N_7500,N_7705);
nand U8470 (N_8470,N_7165,N_7636);
nor U8471 (N_8471,N_7933,N_7895);
nor U8472 (N_8472,N_7149,N_7323);
nand U8473 (N_8473,N_7655,N_7379);
nor U8474 (N_8474,N_7711,N_7581);
nor U8475 (N_8475,N_7827,N_7101);
and U8476 (N_8476,N_7058,N_7180);
or U8477 (N_8477,N_7217,N_7337);
nor U8478 (N_8478,N_7121,N_7098);
nand U8479 (N_8479,N_7634,N_7510);
nor U8480 (N_8480,N_7657,N_7944);
nand U8481 (N_8481,N_7314,N_7599);
xor U8482 (N_8482,N_7773,N_7806);
nand U8483 (N_8483,N_7262,N_7738);
xnor U8484 (N_8484,N_7877,N_7213);
or U8485 (N_8485,N_7625,N_7225);
xor U8486 (N_8486,N_7875,N_7361);
or U8487 (N_8487,N_7100,N_7024);
xnor U8488 (N_8488,N_7701,N_7966);
or U8489 (N_8489,N_7442,N_7571);
and U8490 (N_8490,N_7921,N_7415);
nor U8491 (N_8491,N_7232,N_7779);
nor U8492 (N_8492,N_7671,N_7913);
nor U8493 (N_8493,N_7144,N_7937);
nand U8494 (N_8494,N_7247,N_7347);
nand U8495 (N_8495,N_7224,N_7638);
xnor U8496 (N_8496,N_7077,N_7591);
nor U8497 (N_8497,N_7498,N_7490);
or U8498 (N_8498,N_7380,N_7783);
nor U8499 (N_8499,N_7322,N_7319);
or U8500 (N_8500,N_7089,N_7091);
nand U8501 (N_8501,N_7818,N_7670);
nand U8502 (N_8502,N_7474,N_7364);
and U8503 (N_8503,N_7645,N_7574);
nor U8504 (N_8504,N_7865,N_7156);
nand U8505 (N_8505,N_7398,N_7045);
or U8506 (N_8506,N_7408,N_7607);
nor U8507 (N_8507,N_7674,N_7048);
nor U8508 (N_8508,N_7516,N_7079);
and U8509 (N_8509,N_7251,N_7258);
xor U8510 (N_8510,N_7092,N_7279);
nor U8511 (N_8511,N_7771,N_7271);
and U8512 (N_8512,N_7024,N_7081);
and U8513 (N_8513,N_7863,N_7514);
or U8514 (N_8514,N_7253,N_7783);
nor U8515 (N_8515,N_7085,N_7731);
or U8516 (N_8516,N_7020,N_7312);
xor U8517 (N_8517,N_7431,N_7650);
nor U8518 (N_8518,N_7512,N_7769);
xor U8519 (N_8519,N_7450,N_7088);
xor U8520 (N_8520,N_7911,N_7526);
and U8521 (N_8521,N_7682,N_7391);
and U8522 (N_8522,N_7982,N_7513);
nor U8523 (N_8523,N_7881,N_7173);
xor U8524 (N_8524,N_7689,N_7472);
nand U8525 (N_8525,N_7168,N_7116);
or U8526 (N_8526,N_7234,N_7819);
nor U8527 (N_8527,N_7627,N_7481);
and U8528 (N_8528,N_7189,N_7646);
or U8529 (N_8529,N_7241,N_7109);
and U8530 (N_8530,N_7444,N_7495);
nand U8531 (N_8531,N_7123,N_7150);
and U8532 (N_8532,N_7105,N_7703);
xor U8533 (N_8533,N_7738,N_7053);
and U8534 (N_8534,N_7988,N_7525);
and U8535 (N_8535,N_7444,N_7546);
nor U8536 (N_8536,N_7036,N_7480);
or U8537 (N_8537,N_7544,N_7847);
and U8538 (N_8538,N_7394,N_7580);
or U8539 (N_8539,N_7428,N_7332);
nor U8540 (N_8540,N_7008,N_7689);
nor U8541 (N_8541,N_7391,N_7712);
or U8542 (N_8542,N_7983,N_7726);
xor U8543 (N_8543,N_7150,N_7918);
xnor U8544 (N_8544,N_7176,N_7361);
nand U8545 (N_8545,N_7039,N_7926);
or U8546 (N_8546,N_7129,N_7174);
or U8547 (N_8547,N_7991,N_7347);
and U8548 (N_8548,N_7353,N_7713);
nand U8549 (N_8549,N_7498,N_7771);
nor U8550 (N_8550,N_7455,N_7073);
and U8551 (N_8551,N_7420,N_7542);
xor U8552 (N_8552,N_7959,N_7397);
or U8553 (N_8553,N_7708,N_7516);
or U8554 (N_8554,N_7392,N_7075);
and U8555 (N_8555,N_7019,N_7332);
or U8556 (N_8556,N_7869,N_7876);
or U8557 (N_8557,N_7065,N_7098);
nand U8558 (N_8558,N_7413,N_7131);
and U8559 (N_8559,N_7978,N_7310);
xnor U8560 (N_8560,N_7242,N_7461);
xor U8561 (N_8561,N_7702,N_7410);
nand U8562 (N_8562,N_7750,N_7619);
and U8563 (N_8563,N_7750,N_7153);
nand U8564 (N_8564,N_7318,N_7806);
xnor U8565 (N_8565,N_7562,N_7899);
and U8566 (N_8566,N_7176,N_7871);
and U8567 (N_8567,N_7745,N_7185);
nor U8568 (N_8568,N_7675,N_7604);
xor U8569 (N_8569,N_7221,N_7247);
and U8570 (N_8570,N_7489,N_7522);
or U8571 (N_8571,N_7990,N_7601);
or U8572 (N_8572,N_7647,N_7743);
and U8573 (N_8573,N_7014,N_7916);
nand U8574 (N_8574,N_7122,N_7615);
nand U8575 (N_8575,N_7150,N_7739);
or U8576 (N_8576,N_7503,N_7437);
nand U8577 (N_8577,N_7873,N_7100);
xor U8578 (N_8578,N_7081,N_7186);
and U8579 (N_8579,N_7317,N_7592);
xor U8580 (N_8580,N_7267,N_7096);
or U8581 (N_8581,N_7976,N_7551);
nor U8582 (N_8582,N_7670,N_7466);
xnor U8583 (N_8583,N_7440,N_7822);
and U8584 (N_8584,N_7073,N_7120);
and U8585 (N_8585,N_7969,N_7753);
nor U8586 (N_8586,N_7165,N_7409);
or U8587 (N_8587,N_7830,N_7745);
or U8588 (N_8588,N_7924,N_7786);
nor U8589 (N_8589,N_7602,N_7907);
xor U8590 (N_8590,N_7076,N_7177);
nand U8591 (N_8591,N_7050,N_7807);
or U8592 (N_8592,N_7632,N_7139);
or U8593 (N_8593,N_7497,N_7275);
and U8594 (N_8594,N_7805,N_7626);
and U8595 (N_8595,N_7963,N_7640);
nor U8596 (N_8596,N_7125,N_7670);
nand U8597 (N_8597,N_7302,N_7488);
or U8598 (N_8598,N_7671,N_7956);
nor U8599 (N_8599,N_7828,N_7671);
and U8600 (N_8600,N_7044,N_7305);
and U8601 (N_8601,N_7978,N_7939);
nor U8602 (N_8602,N_7038,N_7886);
nand U8603 (N_8603,N_7776,N_7942);
nor U8604 (N_8604,N_7844,N_7199);
nor U8605 (N_8605,N_7074,N_7435);
or U8606 (N_8606,N_7534,N_7064);
and U8607 (N_8607,N_7250,N_7875);
nor U8608 (N_8608,N_7235,N_7955);
or U8609 (N_8609,N_7154,N_7306);
nor U8610 (N_8610,N_7294,N_7826);
and U8611 (N_8611,N_7295,N_7508);
or U8612 (N_8612,N_7026,N_7166);
and U8613 (N_8613,N_7095,N_7528);
xnor U8614 (N_8614,N_7521,N_7855);
xor U8615 (N_8615,N_7626,N_7190);
xor U8616 (N_8616,N_7217,N_7806);
nor U8617 (N_8617,N_7743,N_7785);
and U8618 (N_8618,N_7727,N_7369);
nor U8619 (N_8619,N_7602,N_7557);
and U8620 (N_8620,N_7655,N_7342);
nand U8621 (N_8621,N_7166,N_7459);
and U8622 (N_8622,N_7912,N_7068);
or U8623 (N_8623,N_7019,N_7733);
nand U8624 (N_8624,N_7677,N_7681);
nor U8625 (N_8625,N_7326,N_7624);
and U8626 (N_8626,N_7698,N_7263);
and U8627 (N_8627,N_7589,N_7439);
nor U8628 (N_8628,N_7798,N_7590);
and U8629 (N_8629,N_7898,N_7369);
xnor U8630 (N_8630,N_7177,N_7803);
xnor U8631 (N_8631,N_7582,N_7081);
nor U8632 (N_8632,N_7418,N_7048);
and U8633 (N_8633,N_7559,N_7870);
or U8634 (N_8634,N_7879,N_7206);
nand U8635 (N_8635,N_7840,N_7706);
nand U8636 (N_8636,N_7495,N_7047);
nor U8637 (N_8637,N_7518,N_7991);
or U8638 (N_8638,N_7117,N_7710);
and U8639 (N_8639,N_7376,N_7768);
and U8640 (N_8640,N_7223,N_7745);
xor U8641 (N_8641,N_7089,N_7364);
or U8642 (N_8642,N_7464,N_7776);
nor U8643 (N_8643,N_7472,N_7273);
nand U8644 (N_8644,N_7797,N_7438);
nor U8645 (N_8645,N_7263,N_7851);
or U8646 (N_8646,N_7719,N_7901);
xnor U8647 (N_8647,N_7904,N_7566);
nor U8648 (N_8648,N_7240,N_7334);
nor U8649 (N_8649,N_7034,N_7950);
nor U8650 (N_8650,N_7251,N_7554);
or U8651 (N_8651,N_7098,N_7735);
and U8652 (N_8652,N_7055,N_7060);
and U8653 (N_8653,N_7421,N_7859);
nor U8654 (N_8654,N_7952,N_7401);
or U8655 (N_8655,N_7890,N_7621);
or U8656 (N_8656,N_7608,N_7304);
nand U8657 (N_8657,N_7713,N_7626);
or U8658 (N_8658,N_7317,N_7022);
nor U8659 (N_8659,N_7686,N_7334);
xnor U8660 (N_8660,N_7876,N_7925);
nor U8661 (N_8661,N_7369,N_7045);
xnor U8662 (N_8662,N_7916,N_7082);
xor U8663 (N_8663,N_7684,N_7156);
nand U8664 (N_8664,N_7640,N_7240);
or U8665 (N_8665,N_7271,N_7780);
nor U8666 (N_8666,N_7056,N_7984);
and U8667 (N_8667,N_7005,N_7050);
xnor U8668 (N_8668,N_7292,N_7125);
and U8669 (N_8669,N_7904,N_7724);
or U8670 (N_8670,N_7448,N_7909);
xnor U8671 (N_8671,N_7570,N_7480);
and U8672 (N_8672,N_7776,N_7641);
nor U8673 (N_8673,N_7754,N_7318);
nor U8674 (N_8674,N_7057,N_7668);
xor U8675 (N_8675,N_7003,N_7992);
nor U8676 (N_8676,N_7060,N_7324);
and U8677 (N_8677,N_7641,N_7570);
nor U8678 (N_8678,N_7469,N_7898);
or U8679 (N_8679,N_7700,N_7215);
nand U8680 (N_8680,N_7816,N_7889);
nand U8681 (N_8681,N_7629,N_7546);
or U8682 (N_8682,N_7228,N_7971);
or U8683 (N_8683,N_7647,N_7073);
or U8684 (N_8684,N_7855,N_7007);
and U8685 (N_8685,N_7516,N_7001);
xor U8686 (N_8686,N_7793,N_7200);
or U8687 (N_8687,N_7257,N_7412);
or U8688 (N_8688,N_7187,N_7026);
nor U8689 (N_8689,N_7385,N_7628);
or U8690 (N_8690,N_7352,N_7057);
nand U8691 (N_8691,N_7386,N_7128);
and U8692 (N_8692,N_7706,N_7522);
or U8693 (N_8693,N_7394,N_7150);
or U8694 (N_8694,N_7228,N_7699);
or U8695 (N_8695,N_7548,N_7472);
xor U8696 (N_8696,N_7317,N_7427);
nor U8697 (N_8697,N_7340,N_7825);
or U8698 (N_8698,N_7847,N_7066);
xor U8699 (N_8699,N_7334,N_7324);
and U8700 (N_8700,N_7998,N_7287);
and U8701 (N_8701,N_7070,N_7237);
and U8702 (N_8702,N_7148,N_7733);
xor U8703 (N_8703,N_7901,N_7392);
and U8704 (N_8704,N_7311,N_7231);
and U8705 (N_8705,N_7611,N_7926);
nand U8706 (N_8706,N_7651,N_7181);
nand U8707 (N_8707,N_7634,N_7541);
xor U8708 (N_8708,N_7154,N_7596);
nand U8709 (N_8709,N_7454,N_7548);
nor U8710 (N_8710,N_7839,N_7451);
or U8711 (N_8711,N_7234,N_7049);
and U8712 (N_8712,N_7970,N_7663);
xnor U8713 (N_8713,N_7768,N_7733);
and U8714 (N_8714,N_7266,N_7392);
and U8715 (N_8715,N_7416,N_7032);
and U8716 (N_8716,N_7925,N_7150);
nor U8717 (N_8717,N_7781,N_7878);
and U8718 (N_8718,N_7148,N_7063);
or U8719 (N_8719,N_7564,N_7343);
nand U8720 (N_8720,N_7684,N_7567);
and U8721 (N_8721,N_7052,N_7974);
or U8722 (N_8722,N_7869,N_7298);
and U8723 (N_8723,N_7221,N_7712);
nand U8724 (N_8724,N_7569,N_7641);
or U8725 (N_8725,N_7242,N_7220);
nand U8726 (N_8726,N_7014,N_7860);
nand U8727 (N_8727,N_7716,N_7643);
or U8728 (N_8728,N_7287,N_7316);
or U8729 (N_8729,N_7992,N_7987);
and U8730 (N_8730,N_7893,N_7596);
nor U8731 (N_8731,N_7375,N_7425);
and U8732 (N_8732,N_7555,N_7056);
and U8733 (N_8733,N_7520,N_7638);
and U8734 (N_8734,N_7412,N_7461);
and U8735 (N_8735,N_7350,N_7127);
nor U8736 (N_8736,N_7399,N_7866);
xor U8737 (N_8737,N_7280,N_7516);
nor U8738 (N_8738,N_7647,N_7781);
nand U8739 (N_8739,N_7923,N_7472);
and U8740 (N_8740,N_7166,N_7804);
nand U8741 (N_8741,N_7037,N_7989);
nor U8742 (N_8742,N_7423,N_7658);
nor U8743 (N_8743,N_7332,N_7835);
nand U8744 (N_8744,N_7307,N_7832);
nor U8745 (N_8745,N_7661,N_7669);
nor U8746 (N_8746,N_7730,N_7927);
and U8747 (N_8747,N_7913,N_7176);
xnor U8748 (N_8748,N_7821,N_7207);
or U8749 (N_8749,N_7984,N_7846);
and U8750 (N_8750,N_7381,N_7622);
nand U8751 (N_8751,N_7261,N_7907);
nor U8752 (N_8752,N_7954,N_7744);
nor U8753 (N_8753,N_7580,N_7876);
and U8754 (N_8754,N_7221,N_7013);
or U8755 (N_8755,N_7343,N_7689);
and U8756 (N_8756,N_7059,N_7893);
or U8757 (N_8757,N_7713,N_7631);
xnor U8758 (N_8758,N_7593,N_7384);
nor U8759 (N_8759,N_7441,N_7287);
xnor U8760 (N_8760,N_7521,N_7566);
and U8761 (N_8761,N_7003,N_7525);
xor U8762 (N_8762,N_7496,N_7439);
or U8763 (N_8763,N_7660,N_7756);
or U8764 (N_8764,N_7881,N_7648);
and U8765 (N_8765,N_7715,N_7452);
xor U8766 (N_8766,N_7620,N_7225);
nand U8767 (N_8767,N_7484,N_7614);
nor U8768 (N_8768,N_7839,N_7160);
and U8769 (N_8769,N_7020,N_7010);
xnor U8770 (N_8770,N_7137,N_7538);
nand U8771 (N_8771,N_7636,N_7697);
nand U8772 (N_8772,N_7109,N_7341);
nand U8773 (N_8773,N_7636,N_7744);
xnor U8774 (N_8774,N_7766,N_7197);
and U8775 (N_8775,N_7743,N_7585);
and U8776 (N_8776,N_7766,N_7686);
nand U8777 (N_8777,N_7391,N_7759);
nand U8778 (N_8778,N_7063,N_7024);
or U8779 (N_8779,N_7410,N_7152);
or U8780 (N_8780,N_7531,N_7795);
xnor U8781 (N_8781,N_7869,N_7266);
and U8782 (N_8782,N_7492,N_7459);
and U8783 (N_8783,N_7124,N_7086);
or U8784 (N_8784,N_7184,N_7460);
and U8785 (N_8785,N_7432,N_7667);
nand U8786 (N_8786,N_7248,N_7322);
nand U8787 (N_8787,N_7253,N_7332);
and U8788 (N_8788,N_7374,N_7330);
and U8789 (N_8789,N_7856,N_7515);
nand U8790 (N_8790,N_7750,N_7841);
xor U8791 (N_8791,N_7555,N_7055);
and U8792 (N_8792,N_7476,N_7493);
xnor U8793 (N_8793,N_7699,N_7842);
xor U8794 (N_8794,N_7974,N_7209);
nor U8795 (N_8795,N_7038,N_7100);
nor U8796 (N_8796,N_7659,N_7837);
or U8797 (N_8797,N_7561,N_7984);
nor U8798 (N_8798,N_7203,N_7211);
nand U8799 (N_8799,N_7681,N_7746);
nand U8800 (N_8800,N_7862,N_7437);
xor U8801 (N_8801,N_7622,N_7695);
xnor U8802 (N_8802,N_7567,N_7292);
xor U8803 (N_8803,N_7635,N_7537);
or U8804 (N_8804,N_7645,N_7353);
nor U8805 (N_8805,N_7846,N_7712);
xor U8806 (N_8806,N_7357,N_7468);
nor U8807 (N_8807,N_7411,N_7307);
or U8808 (N_8808,N_7894,N_7243);
nand U8809 (N_8809,N_7407,N_7579);
and U8810 (N_8810,N_7536,N_7315);
and U8811 (N_8811,N_7551,N_7827);
nand U8812 (N_8812,N_7514,N_7531);
xor U8813 (N_8813,N_7748,N_7143);
xor U8814 (N_8814,N_7964,N_7186);
and U8815 (N_8815,N_7505,N_7675);
nor U8816 (N_8816,N_7486,N_7327);
nor U8817 (N_8817,N_7009,N_7807);
and U8818 (N_8818,N_7507,N_7307);
xnor U8819 (N_8819,N_7587,N_7761);
or U8820 (N_8820,N_7106,N_7180);
or U8821 (N_8821,N_7604,N_7014);
or U8822 (N_8822,N_7635,N_7371);
or U8823 (N_8823,N_7817,N_7577);
xnor U8824 (N_8824,N_7029,N_7440);
xnor U8825 (N_8825,N_7979,N_7920);
or U8826 (N_8826,N_7819,N_7461);
nand U8827 (N_8827,N_7538,N_7423);
and U8828 (N_8828,N_7256,N_7164);
nor U8829 (N_8829,N_7505,N_7160);
or U8830 (N_8830,N_7759,N_7988);
nand U8831 (N_8831,N_7237,N_7355);
nor U8832 (N_8832,N_7567,N_7979);
nand U8833 (N_8833,N_7862,N_7935);
nand U8834 (N_8834,N_7151,N_7244);
and U8835 (N_8835,N_7079,N_7152);
and U8836 (N_8836,N_7787,N_7988);
and U8837 (N_8837,N_7681,N_7794);
xor U8838 (N_8838,N_7910,N_7350);
xor U8839 (N_8839,N_7237,N_7762);
and U8840 (N_8840,N_7408,N_7619);
nand U8841 (N_8841,N_7249,N_7765);
nor U8842 (N_8842,N_7350,N_7044);
xor U8843 (N_8843,N_7562,N_7613);
xnor U8844 (N_8844,N_7566,N_7027);
nand U8845 (N_8845,N_7794,N_7005);
xnor U8846 (N_8846,N_7655,N_7144);
or U8847 (N_8847,N_7986,N_7886);
xor U8848 (N_8848,N_7732,N_7593);
nor U8849 (N_8849,N_7150,N_7071);
nand U8850 (N_8850,N_7110,N_7562);
xnor U8851 (N_8851,N_7665,N_7777);
or U8852 (N_8852,N_7829,N_7347);
nand U8853 (N_8853,N_7031,N_7121);
nor U8854 (N_8854,N_7486,N_7644);
nor U8855 (N_8855,N_7942,N_7442);
nor U8856 (N_8856,N_7961,N_7964);
nand U8857 (N_8857,N_7560,N_7083);
or U8858 (N_8858,N_7669,N_7940);
nor U8859 (N_8859,N_7501,N_7393);
xor U8860 (N_8860,N_7676,N_7217);
or U8861 (N_8861,N_7487,N_7357);
and U8862 (N_8862,N_7965,N_7141);
or U8863 (N_8863,N_7918,N_7543);
and U8864 (N_8864,N_7897,N_7129);
xor U8865 (N_8865,N_7739,N_7716);
and U8866 (N_8866,N_7718,N_7299);
xor U8867 (N_8867,N_7105,N_7125);
xnor U8868 (N_8868,N_7389,N_7283);
and U8869 (N_8869,N_7055,N_7499);
nor U8870 (N_8870,N_7163,N_7381);
or U8871 (N_8871,N_7056,N_7320);
nand U8872 (N_8872,N_7175,N_7293);
nor U8873 (N_8873,N_7740,N_7469);
nor U8874 (N_8874,N_7787,N_7834);
xor U8875 (N_8875,N_7786,N_7246);
xnor U8876 (N_8876,N_7158,N_7452);
and U8877 (N_8877,N_7850,N_7481);
nor U8878 (N_8878,N_7185,N_7344);
xor U8879 (N_8879,N_7512,N_7171);
and U8880 (N_8880,N_7858,N_7582);
or U8881 (N_8881,N_7716,N_7177);
xnor U8882 (N_8882,N_7040,N_7339);
nand U8883 (N_8883,N_7891,N_7534);
xor U8884 (N_8884,N_7835,N_7839);
or U8885 (N_8885,N_7120,N_7779);
nor U8886 (N_8886,N_7076,N_7515);
nand U8887 (N_8887,N_7639,N_7104);
xor U8888 (N_8888,N_7538,N_7777);
and U8889 (N_8889,N_7513,N_7077);
and U8890 (N_8890,N_7001,N_7899);
nor U8891 (N_8891,N_7326,N_7658);
nor U8892 (N_8892,N_7565,N_7705);
nand U8893 (N_8893,N_7803,N_7610);
xnor U8894 (N_8894,N_7430,N_7886);
or U8895 (N_8895,N_7367,N_7597);
nor U8896 (N_8896,N_7968,N_7421);
or U8897 (N_8897,N_7786,N_7334);
nor U8898 (N_8898,N_7968,N_7193);
and U8899 (N_8899,N_7067,N_7694);
xor U8900 (N_8900,N_7868,N_7220);
xor U8901 (N_8901,N_7376,N_7182);
nor U8902 (N_8902,N_7024,N_7253);
or U8903 (N_8903,N_7073,N_7741);
nand U8904 (N_8904,N_7239,N_7590);
nand U8905 (N_8905,N_7637,N_7829);
nand U8906 (N_8906,N_7800,N_7769);
or U8907 (N_8907,N_7607,N_7083);
and U8908 (N_8908,N_7295,N_7149);
xor U8909 (N_8909,N_7890,N_7048);
nand U8910 (N_8910,N_7551,N_7889);
nand U8911 (N_8911,N_7234,N_7359);
and U8912 (N_8912,N_7326,N_7299);
nor U8913 (N_8913,N_7253,N_7651);
nor U8914 (N_8914,N_7232,N_7639);
nand U8915 (N_8915,N_7921,N_7239);
nand U8916 (N_8916,N_7920,N_7095);
nor U8917 (N_8917,N_7438,N_7674);
xor U8918 (N_8918,N_7273,N_7645);
nand U8919 (N_8919,N_7728,N_7044);
nor U8920 (N_8920,N_7160,N_7829);
nor U8921 (N_8921,N_7367,N_7227);
xor U8922 (N_8922,N_7374,N_7395);
or U8923 (N_8923,N_7452,N_7559);
or U8924 (N_8924,N_7013,N_7420);
or U8925 (N_8925,N_7959,N_7336);
nor U8926 (N_8926,N_7258,N_7187);
xnor U8927 (N_8927,N_7802,N_7689);
nor U8928 (N_8928,N_7041,N_7019);
and U8929 (N_8929,N_7527,N_7141);
or U8930 (N_8930,N_7578,N_7993);
nor U8931 (N_8931,N_7653,N_7247);
xor U8932 (N_8932,N_7647,N_7870);
nand U8933 (N_8933,N_7167,N_7259);
nand U8934 (N_8934,N_7924,N_7379);
xor U8935 (N_8935,N_7590,N_7107);
nor U8936 (N_8936,N_7182,N_7488);
or U8937 (N_8937,N_7161,N_7183);
xor U8938 (N_8938,N_7930,N_7703);
xnor U8939 (N_8939,N_7098,N_7971);
or U8940 (N_8940,N_7134,N_7625);
nor U8941 (N_8941,N_7662,N_7410);
nand U8942 (N_8942,N_7302,N_7748);
nor U8943 (N_8943,N_7227,N_7536);
and U8944 (N_8944,N_7714,N_7198);
or U8945 (N_8945,N_7855,N_7936);
nand U8946 (N_8946,N_7043,N_7127);
xor U8947 (N_8947,N_7931,N_7675);
nand U8948 (N_8948,N_7287,N_7582);
xnor U8949 (N_8949,N_7552,N_7440);
or U8950 (N_8950,N_7689,N_7427);
and U8951 (N_8951,N_7083,N_7090);
or U8952 (N_8952,N_7222,N_7220);
xor U8953 (N_8953,N_7738,N_7568);
and U8954 (N_8954,N_7338,N_7367);
xnor U8955 (N_8955,N_7496,N_7837);
nor U8956 (N_8956,N_7393,N_7076);
and U8957 (N_8957,N_7614,N_7822);
nand U8958 (N_8958,N_7229,N_7114);
xor U8959 (N_8959,N_7944,N_7089);
nand U8960 (N_8960,N_7615,N_7835);
or U8961 (N_8961,N_7501,N_7223);
nand U8962 (N_8962,N_7055,N_7174);
and U8963 (N_8963,N_7948,N_7538);
or U8964 (N_8964,N_7499,N_7178);
or U8965 (N_8965,N_7956,N_7564);
xor U8966 (N_8966,N_7169,N_7501);
or U8967 (N_8967,N_7820,N_7665);
nand U8968 (N_8968,N_7033,N_7601);
or U8969 (N_8969,N_7678,N_7041);
or U8970 (N_8970,N_7656,N_7095);
or U8971 (N_8971,N_7916,N_7886);
or U8972 (N_8972,N_7440,N_7515);
or U8973 (N_8973,N_7409,N_7302);
or U8974 (N_8974,N_7045,N_7251);
xnor U8975 (N_8975,N_7878,N_7834);
nor U8976 (N_8976,N_7159,N_7077);
and U8977 (N_8977,N_7104,N_7407);
and U8978 (N_8978,N_7481,N_7941);
and U8979 (N_8979,N_7222,N_7138);
nor U8980 (N_8980,N_7489,N_7501);
xnor U8981 (N_8981,N_7449,N_7520);
or U8982 (N_8982,N_7082,N_7176);
and U8983 (N_8983,N_7384,N_7637);
and U8984 (N_8984,N_7607,N_7754);
nand U8985 (N_8985,N_7289,N_7910);
nor U8986 (N_8986,N_7553,N_7076);
xor U8987 (N_8987,N_7248,N_7504);
nand U8988 (N_8988,N_7454,N_7721);
xnor U8989 (N_8989,N_7017,N_7196);
nand U8990 (N_8990,N_7652,N_7805);
and U8991 (N_8991,N_7321,N_7888);
nor U8992 (N_8992,N_7517,N_7667);
xor U8993 (N_8993,N_7533,N_7076);
xnor U8994 (N_8994,N_7718,N_7891);
nor U8995 (N_8995,N_7434,N_7239);
xnor U8996 (N_8996,N_7533,N_7330);
nor U8997 (N_8997,N_7590,N_7901);
and U8998 (N_8998,N_7746,N_7303);
nor U8999 (N_8999,N_7006,N_7881);
nor U9000 (N_9000,N_8456,N_8032);
nor U9001 (N_9001,N_8700,N_8674);
and U9002 (N_9002,N_8633,N_8308);
xor U9003 (N_9003,N_8647,N_8194);
nand U9004 (N_9004,N_8412,N_8475);
nand U9005 (N_9005,N_8084,N_8454);
nand U9006 (N_9006,N_8075,N_8330);
nand U9007 (N_9007,N_8711,N_8112);
xor U9008 (N_9008,N_8147,N_8615);
and U9009 (N_9009,N_8855,N_8940);
nand U9010 (N_9010,N_8728,N_8152);
xnor U9011 (N_9011,N_8684,N_8737);
nor U9012 (N_9012,N_8401,N_8122);
xor U9013 (N_9013,N_8842,N_8587);
and U9014 (N_9014,N_8971,N_8759);
or U9015 (N_9015,N_8227,N_8080);
xor U9016 (N_9016,N_8963,N_8572);
nor U9017 (N_9017,N_8616,N_8988);
xor U9018 (N_9018,N_8070,N_8025);
nand U9019 (N_9019,N_8607,N_8492);
and U9020 (N_9020,N_8861,N_8409);
and U9021 (N_9021,N_8528,N_8134);
nor U9022 (N_9022,N_8160,N_8329);
nand U9023 (N_9023,N_8441,N_8175);
nor U9024 (N_9024,N_8305,N_8664);
and U9025 (N_9025,N_8127,N_8012);
or U9026 (N_9026,N_8369,N_8884);
xor U9027 (N_9027,N_8229,N_8179);
or U9028 (N_9028,N_8508,N_8877);
nand U9029 (N_9029,N_8818,N_8773);
nand U9030 (N_9030,N_8746,N_8280);
and U9031 (N_9031,N_8310,N_8217);
or U9032 (N_9032,N_8094,N_8361);
nand U9033 (N_9033,N_8610,N_8091);
xnor U9034 (N_9034,N_8594,N_8778);
and U9035 (N_9035,N_8619,N_8126);
and U9036 (N_9036,N_8891,N_8827);
or U9037 (N_9037,N_8709,N_8923);
xor U9038 (N_9038,N_8113,N_8105);
or U9039 (N_9039,N_8398,N_8964);
xnor U9040 (N_9040,N_8789,N_8244);
and U9041 (N_9041,N_8564,N_8052);
xor U9042 (N_9042,N_8506,N_8394);
and U9043 (N_9043,N_8035,N_8557);
and U9044 (N_9044,N_8829,N_8912);
and U9045 (N_9045,N_8274,N_8540);
and U9046 (N_9046,N_8416,N_8031);
nand U9047 (N_9047,N_8747,N_8464);
xnor U9048 (N_9048,N_8267,N_8142);
and U9049 (N_9049,N_8872,N_8887);
and U9050 (N_9050,N_8439,N_8016);
xnor U9051 (N_9051,N_8799,N_8103);
or U9052 (N_9052,N_8751,N_8804);
nand U9053 (N_9053,N_8212,N_8284);
and U9054 (N_9054,N_8694,N_8762);
nand U9055 (N_9055,N_8967,N_8365);
nor U9056 (N_9056,N_8748,N_8315);
nand U9057 (N_9057,N_8422,N_8362);
xor U9058 (N_9058,N_8187,N_8965);
and U9059 (N_9059,N_8661,N_8133);
xnor U9060 (N_9060,N_8955,N_8867);
and U9061 (N_9061,N_8874,N_8438);
nor U9062 (N_9062,N_8022,N_8523);
nor U9063 (N_9063,N_8620,N_8485);
nand U9064 (N_9064,N_8073,N_8155);
and U9065 (N_9065,N_8929,N_8268);
nor U9066 (N_9066,N_8351,N_8192);
nand U9067 (N_9067,N_8801,N_8513);
nor U9068 (N_9068,N_8333,N_8800);
nand U9069 (N_9069,N_8776,N_8784);
xnor U9070 (N_9070,N_8288,N_8332);
nand U9071 (N_9071,N_8995,N_8770);
nand U9072 (N_9072,N_8430,N_8658);
nor U9073 (N_9073,N_8823,N_8785);
nand U9074 (N_9074,N_8273,N_8937);
nor U9075 (N_9075,N_8612,N_8418);
and U9076 (N_9076,N_8889,N_8825);
and U9077 (N_9077,N_8260,N_8791);
or U9078 (N_9078,N_8370,N_8426);
xnor U9079 (N_9079,N_8579,N_8393);
nor U9080 (N_9080,N_8580,N_8111);
xor U9081 (N_9081,N_8742,N_8519);
and U9082 (N_9082,N_8537,N_8072);
or U9083 (N_9083,N_8752,N_8974);
nor U9084 (N_9084,N_8359,N_8435);
or U9085 (N_9085,N_8253,N_8191);
nor U9086 (N_9086,N_8527,N_8905);
and U9087 (N_9087,N_8314,N_8851);
xor U9088 (N_9088,N_8136,N_8036);
nor U9089 (N_9089,N_8856,N_8657);
or U9090 (N_9090,N_8681,N_8379);
nor U9091 (N_9091,N_8337,N_8037);
nand U9092 (N_9092,N_8881,N_8535);
nor U9093 (N_9093,N_8555,N_8685);
and U9094 (N_9094,N_8900,N_8691);
nor U9095 (N_9095,N_8138,N_8821);
nor U9096 (N_9096,N_8522,N_8899);
or U9097 (N_9097,N_8950,N_8407);
nand U9098 (N_9098,N_8767,N_8734);
nand U9099 (N_9099,N_8001,N_8882);
or U9100 (N_9100,N_8859,N_8902);
nand U9101 (N_9101,N_8830,N_8278);
and U9102 (N_9102,N_8713,N_8511);
nor U9103 (N_9103,N_8088,N_8654);
xnor U9104 (N_9104,N_8547,N_8993);
and U9105 (N_9105,N_8312,N_8196);
nand U9106 (N_9106,N_8245,N_8125);
nor U9107 (N_9107,N_8053,N_8501);
xor U9108 (N_9108,N_8864,N_8741);
or U9109 (N_9109,N_8857,N_8195);
nand U9110 (N_9110,N_8771,N_8590);
and U9111 (N_9111,N_8660,N_8099);
or U9112 (N_9112,N_8903,N_8478);
or U9113 (N_9113,N_8530,N_8832);
or U9114 (N_9114,N_8353,N_8836);
nor U9115 (N_9115,N_8679,N_8917);
and U9116 (N_9116,N_8833,N_8328);
xnor U9117 (N_9117,N_8690,N_8976);
and U9118 (N_9118,N_8671,N_8895);
xnor U9119 (N_9119,N_8300,N_8597);
and U9120 (N_9120,N_8999,N_8434);
nor U9121 (N_9121,N_8500,N_8045);
nand U9122 (N_9122,N_8461,N_8603);
nor U9123 (N_9123,N_8687,N_8556);
nor U9124 (N_9124,N_8712,N_8287);
xnor U9125 (N_9125,N_8391,N_8890);
nand U9126 (N_9126,N_8472,N_8197);
nor U9127 (N_9127,N_8371,N_8958);
or U9128 (N_9128,N_8468,N_8169);
nor U9129 (N_9129,N_8521,N_8460);
or U9130 (N_9130,N_8384,N_8349);
xor U9131 (N_9131,N_8683,N_8060);
xor U9132 (N_9132,N_8813,N_8865);
nor U9133 (N_9133,N_8516,N_8699);
nand U9134 (N_9134,N_8517,N_8390);
or U9135 (N_9135,N_8188,N_8056);
nand U9136 (N_9136,N_8172,N_8893);
nand U9137 (N_9137,N_8583,N_8512);
xnor U9138 (N_9138,N_8628,N_8130);
or U9139 (N_9139,N_8471,N_8225);
nand U9140 (N_9140,N_8841,N_8098);
nand U9141 (N_9141,N_8562,N_8726);
xnor U9142 (N_9142,N_8210,N_8296);
xnor U9143 (N_9143,N_8824,N_8624);
nand U9144 (N_9144,N_8845,N_8843);
xor U9145 (N_9145,N_8062,N_8885);
nand U9146 (N_9146,N_8490,N_8121);
nand U9147 (N_9147,N_8896,N_8402);
xor U9148 (N_9148,N_8381,N_8289);
xor U9149 (N_9149,N_8419,N_8208);
and U9150 (N_9150,N_8935,N_8008);
and U9151 (N_9151,N_8246,N_8835);
and U9152 (N_9152,N_8352,N_8497);
nand U9153 (N_9153,N_8163,N_8588);
xnor U9154 (N_9154,N_8334,N_8151);
nand U9155 (N_9155,N_8545,N_8368);
nand U9156 (N_9156,N_8215,N_8346);
nand U9157 (N_9157,N_8421,N_8814);
or U9158 (N_9158,N_8886,N_8470);
and U9159 (N_9159,N_8584,N_8614);
xor U9160 (N_9160,N_8875,N_8449);
or U9161 (N_9161,N_8910,N_8499);
nor U9162 (N_9162,N_8986,N_8730);
nor U9163 (N_9163,N_8367,N_8846);
and U9164 (N_9164,N_8772,N_8577);
or U9165 (N_9165,N_8915,N_8880);
nor U9166 (N_9166,N_8768,N_8107);
and U9167 (N_9167,N_8922,N_8931);
xor U9168 (N_9168,N_8644,N_8014);
nand U9169 (N_9169,N_8567,N_8838);
nor U9170 (N_9170,N_8676,N_8445);
nand U9171 (N_9171,N_8815,N_8481);
nand U9172 (N_9172,N_8114,N_8677);
or U9173 (N_9173,N_8313,N_8951);
and U9174 (N_9174,N_8451,N_8901);
nand U9175 (N_9175,N_8085,N_8593);
nand U9176 (N_9176,N_8326,N_8631);
nor U9177 (N_9177,N_8236,N_8059);
nand U9178 (N_9178,N_8729,N_8532);
xor U9179 (N_9179,N_8578,N_8442);
and U9180 (N_9180,N_8303,N_8488);
nand U9181 (N_9181,N_8656,N_8159);
nor U9182 (N_9182,N_8718,N_8242);
nand U9183 (N_9183,N_8183,N_8042);
nor U9184 (N_9184,N_8000,N_8655);
nand U9185 (N_9185,N_8299,N_8224);
and U9186 (N_9186,N_8808,N_8727);
or U9187 (N_9187,N_8281,N_8604);
nor U9188 (N_9188,N_8831,N_8788);
and U9189 (N_9189,N_8186,N_8177);
and U9190 (N_9190,N_8695,N_8854);
or U9191 (N_9191,N_8176,N_8339);
xor U9192 (N_9192,N_8714,N_8263);
nor U9193 (N_9193,N_8097,N_8476);
and U9194 (N_9194,N_8463,N_8820);
nand U9195 (N_9195,N_8092,N_8642);
nor U9196 (N_9196,N_8926,N_8675);
nand U9197 (N_9197,N_8802,N_8710);
nor U9198 (N_9198,N_8238,N_8182);
or U9199 (N_9199,N_8109,N_8009);
nor U9200 (N_9200,N_8262,N_8888);
nand U9201 (N_9201,N_8150,N_8425);
and U9202 (N_9202,N_8558,N_8010);
or U9203 (N_9203,N_8474,N_8913);
or U9204 (N_9204,N_8252,N_8455);
nor U9205 (N_9205,N_8693,N_8906);
nor U9206 (N_9206,N_8331,N_8118);
xnor U9207 (N_9207,N_8248,N_8431);
nand U9208 (N_9208,N_8291,N_8387);
nand U9209 (N_9209,N_8108,N_8483);
and U9210 (N_9210,N_8294,N_8921);
nand U9211 (N_9211,N_8206,N_8071);
and U9212 (N_9212,N_8209,N_8443);
and U9213 (N_9213,N_8780,N_8892);
nand U9214 (N_9214,N_8319,N_8672);
nand U9215 (N_9215,N_8703,N_8322);
or U9216 (N_9216,N_8436,N_8722);
and U9217 (N_9217,N_8645,N_8302);
xor U9218 (N_9218,N_8247,N_8848);
and U9219 (N_9219,N_8626,N_8634);
nand U9220 (N_9220,N_8731,N_8744);
and U9221 (N_9221,N_8171,N_8058);
xnor U9222 (N_9222,N_8286,N_8592);
nor U9223 (N_9223,N_8417,N_8222);
nor U9224 (N_9224,N_8423,N_8806);
or U9225 (N_9225,N_8199,N_8599);
nand U9226 (N_9226,N_8862,N_8297);
or U9227 (N_9227,N_8311,N_8357);
and U9228 (N_9228,N_8953,N_8480);
and U9229 (N_9229,N_8484,N_8458);
xnor U9230 (N_9230,N_8374,N_8397);
and U9231 (N_9231,N_8618,N_8621);
nor U9232 (N_9232,N_8601,N_8665);
nor U9233 (N_9233,N_8004,N_8948);
nand U9234 (N_9234,N_8574,N_8595);
nor U9235 (N_9235,N_8341,N_8894);
nor U9236 (N_9236,N_8448,N_8934);
and U9237 (N_9237,N_8283,N_8447);
and U9238 (N_9238,N_8927,N_8998);
nand U9239 (N_9239,N_8749,N_8076);
nand U9240 (N_9240,N_8720,N_8064);
nand U9241 (N_9241,N_8026,N_8724);
nand U9242 (N_9242,N_8941,N_8975);
nand U9243 (N_9243,N_8266,N_8055);
and U9244 (N_9244,N_8561,N_8154);
xor U9245 (N_9245,N_8822,N_8198);
and U9246 (N_9246,N_8414,N_8798);
nor U9247 (N_9247,N_8306,N_8548);
nor U9248 (N_9248,N_8068,N_8648);
and U9249 (N_9249,N_8170,N_8494);
and U9250 (N_9250,N_8873,N_8120);
nand U9251 (N_9251,N_8493,N_8486);
and U9252 (N_9252,N_8598,N_8507);
nand U9253 (N_9253,N_8812,N_8290);
nor U9254 (N_9254,N_8013,N_8538);
nand U9255 (N_9255,N_8652,N_8201);
nor U9256 (N_9256,N_8017,N_8137);
nor U9257 (N_9257,N_8256,N_8174);
or U9258 (N_9258,N_8704,N_8809);
xor U9259 (N_9259,N_8868,N_8504);
or U9260 (N_9260,N_8817,N_8144);
and U9261 (N_9261,N_8735,N_8943);
or U9262 (N_9262,N_8968,N_8207);
and U9263 (N_9263,N_8143,N_8420);
nand U9264 (N_9264,N_8944,N_8553);
xnor U9265 (N_9265,N_8750,N_8003);
xnor U9266 (N_9266,N_8057,N_8372);
and U9267 (N_9267,N_8404,N_8219);
xnor U9268 (N_9268,N_8979,N_8632);
or U9269 (N_9269,N_8366,N_8259);
nand U9270 (N_9270,N_8119,N_8793);
xor U9271 (N_9271,N_8688,N_8358);
nor U9272 (N_9272,N_8128,N_8395);
xor U9273 (N_9273,N_8354,N_8295);
nand U9274 (N_9274,N_8503,N_8041);
nand U9275 (N_9275,N_8226,N_8293);
nand U9276 (N_9276,N_8095,N_8011);
and U9277 (N_9277,N_8518,N_8282);
nand U9278 (N_9278,N_8043,N_8309);
nor U9279 (N_9279,N_8651,N_8969);
xor U9280 (N_9280,N_8608,N_8705);
and U9281 (N_9281,N_8849,N_8081);
or U9282 (N_9282,N_8093,N_8870);
or U9283 (N_9283,N_8063,N_8396);
and U9284 (N_9284,N_8863,N_8498);
xor U9285 (N_9285,N_8932,N_8650);
or U9286 (N_9286,N_8181,N_8204);
nor U9287 (N_9287,N_8909,N_8637);
xor U9288 (N_9288,N_8272,N_8686);
xnor U9289 (N_9289,N_8106,N_8415);
or U9290 (N_9290,N_8465,N_8104);
nand U9291 (N_9291,N_8939,N_8110);
and U9292 (N_9292,N_8536,N_8065);
nand U9293 (N_9293,N_8231,N_8027);
nand U9294 (N_9294,N_8596,N_8725);
and U9295 (N_9295,N_8549,N_8129);
nor U9296 (N_9296,N_8585,N_8796);
nor U9297 (N_9297,N_8764,N_8689);
and U9298 (N_9298,N_8066,N_8533);
or U9299 (N_9299,N_8961,N_8586);
and U9300 (N_9300,N_8324,N_8141);
nor U9301 (N_9301,N_8230,N_8509);
nand U9302 (N_9302,N_8040,N_8925);
nand U9303 (N_9303,N_8020,N_8344);
or U9304 (N_9304,N_8707,N_8980);
and U9305 (N_9305,N_8444,N_8525);
or U9306 (N_9306,N_8054,N_8023);
or U9307 (N_9307,N_8738,N_8433);
xnor U9308 (N_9308,N_8156,N_8323);
xnor U9309 (N_9309,N_8839,N_8167);
or U9310 (N_9310,N_8347,N_8149);
nand U9311 (N_9311,N_8706,N_8432);
xor U9312 (N_9312,N_8745,N_8466);
and U9313 (N_9313,N_8692,N_8970);
xor U9314 (N_9314,N_8589,N_8716);
and U9315 (N_9315,N_8570,N_8258);
or U9316 (N_9316,N_8928,N_8542);
nor U9317 (N_9317,N_8479,N_8406);
and U9318 (N_9318,N_8050,N_8203);
xor U9319 (N_9319,N_8904,N_8942);
xnor U9320 (N_9320,N_8617,N_8911);
nor U9321 (N_9321,N_8996,N_8606);
or U9322 (N_9322,N_8505,N_8193);
nand U9323 (N_9323,N_8794,N_8541);
nor U9324 (N_9324,N_8457,N_8218);
and U9325 (N_9325,N_8898,N_8879);
or U9326 (N_9326,N_8719,N_8239);
xnor U9327 (N_9327,N_8277,N_8405);
nor U9328 (N_9328,N_8807,N_8257);
or U9329 (N_9329,N_8697,N_8667);
nor U9330 (N_9330,N_8756,N_8200);
xor U9331 (N_9331,N_8984,N_8006);
nor U9332 (N_9332,N_8145,N_8049);
nand U9333 (N_9333,N_8382,N_8205);
and U9334 (N_9334,N_8496,N_8760);
and U9335 (N_9335,N_8321,N_8166);
nand U9336 (N_9336,N_8779,N_8816);
xor U9337 (N_9337,N_8966,N_8721);
nand U9338 (N_9338,N_8304,N_8837);
nand U9339 (N_9339,N_8467,N_8795);
or U9340 (N_9340,N_8757,N_8930);
xnor U9341 (N_9341,N_8786,N_8947);
xnor U9342 (N_9342,N_8271,N_8213);
nor U9343 (N_9343,N_8221,N_8086);
nand U9344 (N_9344,N_8639,N_8437);
nand U9345 (N_9345,N_8340,N_8514);
or U9346 (N_9346,N_8625,N_8452);
nand U9347 (N_9347,N_8853,N_8858);
nor U9348 (N_9348,N_8413,N_8429);
and U9349 (N_9349,N_8317,N_8918);
nand U9350 (N_9350,N_8543,N_8325);
or U9351 (N_9351,N_8990,N_8916);
or U9352 (N_9352,N_8034,N_8701);
and U9353 (N_9353,N_8410,N_8834);
xor U9354 (N_9354,N_8101,N_8754);
and U9355 (N_9355,N_8960,N_8180);
xor U9356 (N_9356,N_8670,N_8473);
and U9357 (N_9357,N_8285,N_8569);
nand U9358 (N_9358,N_8100,N_8811);
xnor U9359 (N_9359,N_8005,N_8241);
xnor U9360 (N_9360,N_8350,N_8377);
nand U9361 (N_9361,N_8919,N_8202);
xnor U9362 (N_9362,N_8047,N_8972);
xnor U9363 (N_9363,N_8847,N_8019);
or U9364 (N_9364,N_8232,N_8733);
nor U9365 (N_9365,N_8659,N_8028);
nor U9366 (N_9366,N_8261,N_8860);
nand U9367 (N_9367,N_8061,N_8680);
and U9368 (N_9368,N_8949,N_8678);
and U9369 (N_9369,N_8487,N_8938);
xor U9370 (N_9370,N_8534,N_8852);
or U9371 (N_9371,N_8563,N_8327);
nand U9372 (N_9372,N_8082,N_8878);
or U9373 (N_9373,N_8605,N_8029);
or U9374 (N_9374,N_8985,N_8573);
or U9375 (N_9375,N_8168,N_8866);
or U9376 (N_9376,N_8636,N_8345);
nor U9377 (N_9377,N_8761,N_8453);
or U9378 (N_9378,N_8551,N_8717);
and U9379 (N_9379,N_8077,N_8264);
nor U9380 (N_9380,N_8575,N_8758);
xor U9381 (N_9381,N_8783,N_8805);
nor U9382 (N_9382,N_8131,N_8609);
and U9383 (N_9383,N_8276,N_8380);
nand U9384 (N_9384,N_8571,N_8529);
nor U9385 (N_9385,N_8462,N_8320);
nor U9386 (N_9386,N_8769,N_8933);
or U9387 (N_9387,N_8385,N_8907);
and U9388 (N_9388,N_8959,N_8044);
or U9389 (N_9389,N_8775,N_8184);
and U9390 (N_9390,N_8840,N_8069);
nand U9391 (N_9391,N_8002,N_8450);
xnor U9392 (N_9392,N_8030,N_8223);
nand U9393 (N_9393,N_8336,N_8038);
xor U9394 (N_9394,N_8946,N_8662);
and U9395 (N_9395,N_8048,N_8810);
and U9396 (N_9396,N_8153,N_8559);
or U9397 (N_9397,N_8243,N_8446);
or U9398 (N_9398,N_8781,N_8292);
xor U9399 (N_9399,N_8790,N_8146);
nand U9400 (N_9400,N_8024,N_8954);
nor U9401 (N_9401,N_8869,N_8356);
or U9402 (N_9402,N_8702,N_8338);
nor U9403 (N_9403,N_8997,N_8161);
nor U9404 (N_9404,N_8576,N_8673);
nor U9405 (N_9405,N_8386,N_8682);
nor U9406 (N_9406,N_8235,N_8623);
nand U9407 (N_9407,N_8973,N_8550);
or U9408 (N_9408,N_8469,N_8335);
nor U9409 (N_9409,N_8477,N_8774);
nand U9410 (N_9410,N_8039,N_8007);
nor U9411 (N_9411,N_8920,N_8270);
nor U9412 (N_9412,N_8178,N_8117);
nand U9413 (N_9413,N_8135,N_8740);
xor U9414 (N_9414,N_8755,N_8428);
or U9415 (N_9415,N_8568,N_8627);
nor U9416 (N_9416,N_8234,N_8945);
and U9417 (N_9417,N_8364,N_8360);
and U9418 (N_9418,N_8565,N_8373);
nor U9419 (N_9419,N_8250,N_8526);
nand U9420 (N_9420,N_8090,N_8240);
and U9421 (N_9421,N_8819,N_8826);
nor U9422 (N_9422,N_8515,N_8307);
xnor U9423 (N_9423,N_8763,N_8992);
or U9424 (N_9424,N_8994,N_8696);
xor U9425 (N_9425,N_8643,N_8348);
xnor U9426 (N_9426,N_8539,N_8638);
xnor U9427 (N_9427,N_8981,N_8237);
nand U9428 (N_9428,N_8777,N_8228);
and U9429 (N_9429,N_8427,N_8924);
or U9430 (N_9430,N_8298,N_8622);
and U9431 (N_9431,N_8411,N_8115);
nor U9432 (N_9432,N_8736,N_8962);
and U9433 (N_9433,N_8897,N_8275);
nor U9434 (N_9434,N_8316,N_8591);
xnor U9435 (N_9435,N_8318,N_8502);
nor U9436 (N_9436,N_8765,N_8083);
and U9437 (N_9437,N_8560,N_8124);
nor U9438 (N_9438,N_8033,N_8046);
nor U9439 (N_9439,N_8668,N_8666);
nand U9440 (N_9440,N_8342,N_8797);
nand U9441 (N_9441,N_8546,N_8343);
and U9442 (N_9442,N_8520,N_8723);
or U9443 (N_9443,N_8871,N_8613);
xor U9444 (N_9444,N_8189,N_8440);
nor U9445 (N_9445,N_8977,N_8355);
nor U9446 (N_9446,N_8403,N_8646);
or U9447 (N_9447,N_8495,N_8978);
nor U9448 (N_9448,N_8635,N_8482);
or U9449 (N_9449,N_8400,N_8363);
nand U9450 (N_9450,N_8408,N_8732);
and U9451 (N_9451,N_8582,N_8708);
xor U9452 (N_9452,N_8123,N_8641);
and U9453 (N_9453,N_8376,N_8255);
xnor U9454 (N_9454,N_8162,N_8956);
nand U9455 (N_9455,N_8139,N_8883);
nand U9456 (N_9456,N_8378,N_8743);
nor U9457 (N_9457,N_8792,N_8216);
and U9458 (N_9458,N_8489,N_8249);
xnor U9459 (N_9459,N_8787,N_8383);
nand U9460 (N_9460,N_8018,N_8078);
nand U9461 (N_9461,N_8089,N_8987);
or U9462 (N_9462,N_8640,N_8254);
nor U9463 (N_9463,N_8491,N_8051);
nand U9464 (N_9464,N_8301,N_8388);
xnor U9465 (N_9465,N_8164,N_8581);
nand U9466 (N_9466,N_8269,N_8265);
nor U9467 (N_9467,N_8936,N_8140);
nor U9468 (N_9468,N_8698,N_8600);
xor U9469 (N_9469,N_8663,N_8079);
or U9470 (N_9470,N_8279,N_8611);
nor U9471 (N_9471,N_8116,N_8982);
nor U9472 (N_9472,N_8629,N_8991);
nand U9473 (N_9473,N_8067,N_8251);
xor U9474 (N_9474,N_8828,N_8165);
nor U9475 (N_9475,N_8908,N_8389);
and U9476 (N_9476,N_8566,N_8715);
nand U9477 (N_9477,N_8649,N_8148);
and U9478 (N_9478,N_8375,N_8957);
or U9479 (N_9479,N_8850,N_8602);
or U9480 (N_9480,N_8653,N_8544);
and U9481 (N_9481,N_8989,N_8510);
and U9482 (N_9482,N_8102,N_8074);
nor U9483 (N_9483,N_8739,N_8190);
and U9484 (N_9484,N_8021,N_8630);
and U9485 (N_9485,N_8844,N_8173);
xnor U9486 (N_9486,N_8531,N_8211);
and U9487 (N_9487,N_8157,N_8983);
nor U9488 (N_9488,N_8782,N_8015);
nand U9489 (N_9489,N_8669,N_8096);
and U9490 (N_9490,N_8914,N_8132);
and U9491 (N_9491,N_8554,N_8185);
or U9492 (N_9492,N_8459,N_8552);
or U9493 (N_9493,N_8214,N_8524);
and U9494 (N_9494,N_8392,N_8158);
or U9495 (N_9495,N_8876,N_8087);
xor U9496 (N_9496,N_8803,N_8220);
nand U9497 (N_9497,N_8233,N_8753);
or U9498 (N_9498,N_8952,N_8766);
and U9499 (N_9499,N_8399,N_8424);
or U9500 (N_9500,N_8916,N_8489);
or U9501 (N_9501,N_8120,N_8715);
or U9502 (N_9502,N_8754,N_8492);
nand U9503 (N_9503,N_8331,N_8192);
nor U9504 (N_9504,N_8104,N_8608);
or U9505 (N_9505,N_8510,N_8015);
nand U9506 (N_9506,N_8056,N_8149);
and U9507 (N_9507,N_8438,N_8467);
and U9508 (N_9508,N_8634,N_8942);
nor U9509 (N_9509,N_8872,N_8477);
nand U9510 (N_9510,N_8080,N_8190);
and U9511 (N_9511,N_8639,N_8291);
xnor U9512 (N_9512,N_8177,N_8495);
and U9513 (N_9513,N_8785,N_8025);
xor U9514 (N_9514,N_8820,N_8159);
nor U9515 (N_9515,N_8598,N_8319);
and U9516 (N_9516,N_8078,N_8387);
xor U9517 (N_9517,N_8018,N_8229);
nand U9518 (N_9518,N_8618,N_8405);
and U9519 (N_9519,N_8291,N_8733);
and U9520 (N_9520,N_8078,N_8919);
nor U9521 (N_9521,N_8018,N_8082);
xnor U9522 (N_9522,N_8031,N_8098);
and U9523 (N_9523,N_8453,N_8139);
nand U9524 (N_9524,N_8839,N_8903);
xor U9525 (N_9525,N_8426,N_8636);
nor U9526 (N_9526,N_8166,N_8975);
nand U9527 (N_9527,N_8074,N_8889);
nand U9528 (N_9528,N_8838,N_8938);
xnor U9529 (N_9529,N_8501,N_8027);
nand U9530 (N_9530,N_8507,N_8320);
xnor U9531 (N_9531,N_8735,N_8039);
or U9532 (N_9532,N_8997,N_8070);
or U9533 (N_9533,N_8591,N_8195);
xnor U9534 (N_9534,N_8785,N_8328);
nand U9535 (N_9535,N_8104,N_8096);
nand U9536 (N_9536,N_8654,N_8949);
xnor U9537 (N_9537,N_8510,N_8169);
or U9538 (N_9538,N_8484,N_8369);
nand U9539 (N_9539,N_8173,N_8883);
or U9540 (N_9540,N_8522,N_8072);
and U9541 (N_9541,N_8597,N_8548);
nor U9542 (N_9542,N_8789,N_8522);
xnor U9543 (N_9543,N_8650,N_8138);
xor U9544 (N_9544,N_8238,N_8848);
nand U9545 (N_9545,N_8433,N_8666);
nand U9546 (N_9546,N_8953,N_8506);
nand U9547 (N_9547,N_8932,N_8489);
and U9548 (N_9548,N_8117,N_8758);
xnor U9549 (N_9549,N_8789,N_8914);
nor U9550 (N_9550,N_8025,N_8419);
nand U9551 (N_9551,N_8794,N_8248);
nand U9552 (N_9552,N_8610,N_8107);
or U9553 (N_9553,N_8912,N_8178);
nor U9554 (N_9554,N_8570,N_8743);
nor U9555 (N_9555,N_8950,N_8108);
xor U9556 (N_9556,N_8202,N_8418);
or U9557 (N_9557,N_8357,N_8111);
xor U9558 (N_9558,N_8786,N_8617);
nor U9559 (N_9559,N_8397,N_8033);
nand U9560 (N_9560,N_8336,N_8517);
nand U9561 (N_9561,N_8708,N_8406);
xnor U9562 (N_9562,N_8064,N_8146);
nand U9563 (N_9563,N_8750,N_8230);
and U9564 (N_9564,N_8956,N_8652);
nand U9565 (N_9565,N_8371,N_8014);
or U9566 (N_9566,N_8261,N_8886);
and U9567 (N_9567,N_8389,N_8489);
nand U9568 (N_9568,N_8793,N_8327);
nand U9569 (N_9569,N_8362,N_8043);
nor U9570 (N_9570,N_8064,N_8202);
nand U9571 (N_9571,N_8393,N_8275);
nor U9572 (N_9572,N_8825,N_8368);
xnor U9573 (N_9573,N_8826,N_8541);
nor U9574 (N_9574,N_8888,N_8785);
or U9575 (N_9575,N_8552,N_8336);
xor U9576 (N_9576,N_8384,N_8377);
nor U9577 (N_9577,N_8502,N_8215);
and U9578 (N_9578,N_8176,N_8525);
nand U9579 (N_9579,N_8714,N_8991);
or U9580 (N_9580,N_8300,N_8197);
xor U9581 (N_9581,N_8834,N_8909);
or U9582 (N_9582,N_8356,N_8063);
or U9583 (N_9583,N_8134,N_8609);
nand U9584 (N_9584,N_8074,N_8780);
nand U9585 (N_9585,N_8070,N_8856);
nand U9586 (N_9586,N_8347,N_8181);
nand U9587 (N_9587,N_8609,N_8349);
nand U9588 (N_9588,N_8690,N_8637);
or U9589 (N_9589,N_8028,N_8258);
or U9590 (N_9590,N_8885,N_8337);
or U9591 (N_9591,N_8900,N_8122);
and U9592 (N_9592,N_8568,N_8449);
nand U9593 (N_9593,N_8839,N_8987);
and U9594 (N_9594,N_8691,N_8877);
nand U9595 (N_9595,N_8422,N_8010);
nor U9596 (N_9596,N_8872,N_8244);
and U9597 (N_9597,N_8893,N_8094);
or U9598 (N_9598,N_8805,N_8203);
nand U9599 (N_9599,N_8363,N_8230);
xnor U9600 (N_9600,N_8810,N_8256);
and U9601 (N_9601,N_8753,N_8371);
nor U9602 (N_9602,N_8355,N_8775);
and U9603 (N_9603,N_8075,N_8055);
or U9604 (N_9604,N_8481,N_8804);
or U9605 (N_9605,N_8777,N_8794);
xnor U9606 (N_9606,N_8267,N_8907);
or U9607 (N_9607,N_8646,N_8896);
nor U9608 (N_9608,N_8505,N_8019);
xnor U9609 (N_9609,N_8086,N_8546);
nor U9610 (N_9610,N_8912,N_8537);
nor U9611 (N_9611,N_8621,N_8256);
xnor U9612 (N_9612,N_8951,N_8085);
xnor U9613 (N_9613,N_8116,N_8403);
nand U9614 (N_9614,N_8571,N_8276);
or U9615 (N_9615,N_8590,N_8083);
or U9616 (N_9616,N_8776,N_8361);
and U9617 (N_9617,N_8714,N_8473);
nand U9618 (N_9618,N_8750,N_8712);
nor U9619 (N_9619,N_8321,N_8021);
xnor U9620 (N_9620,N_8307,N_8690);
xnor U9621 (N_9621,N_8520,N_8925);
nor U9622 (N_9622,N_8065,N_8074);
xor U9623 (N_9623,N_8165,N_8563);
or U9624 (N_9624,N_8769,N_8601);
or U9625 (N_9625,N_8893,N_8260);
nor U9626 (N_9626,N_8736,N_8517);
and U9627 (N_9627,N_8918,N_8384);
or U9628 (N_9628,N_8466,N_8141);
or U9629 (N_9629,N_8639,N_8400);
xnor U9630 (N_9630,N_8520,N_8913);
xor U9631 (N_9631,N_8290,N_8361);
nand U9632 (N_9632,N_8904,N_8217);
nand U9633 (N_9633,N_8850,N_8170);
nand U9634 (N_9634,N_8532,N_8355);
nand U9635 (N_9635,N_8593,N_8525);
nor U9636 (N_9636,N_8564,N_8708);
and U9637 (N_9637,N_8964,N_8082);
and U9638 (N_9638,N_8804,N_8020);
and U9639 (N_9639,N_8051,N_8149);
or U9640 (N_9640,N_8797,N_8488);
and U9641 (N_9641,N_8549,N_8915);
nor U9642 (N_9642,N_8753,N_8166);
xor U9643 (N_9643,N_8136,N_8349);
and U9644 (N_9644,N_8696,N_8136);
xnor U9645 (N_9645,N_8696,N_8065);
or U9646 (N_9646,N_8785,N_8897);
xor U9647 (N_9647,N_8638,N_8043);
nor U9648 (N_9648,N_8091,N_8799);
or U9649 (N_9649,N_8263,N_8709);
and U9650 (N_9650,N_8373,N_8269);
nand U9651 (N_9651,N_8048,N_8285);
and U9652 (N_9652,N_8550,N_8715);
and U9653 (N_9653,N_8529,N_8570);
nand U9654 (N_9654,N_8473,N_8069);
or U9655 (N_9655,N_8975,N_8853);
nor U9656 (N_9656,N_8924,N_8611);
nand U9657 (N_9657,N_8447,N_8989);
nor U9658 (N_9658,N_8743,N_8992);
nand U9659 (N_9659,N_8671,N_8003);
xor U9660 (N_9660,N_8905,N_8449);
nor U9661 (N_9661,N_8332,N_8978);
or U9662 (N_9662,N_8048,N_8220);
and U9663 (N_9663,N_8255,N_8308);
nand U9664 (N_9664,N_8552,N_8549);
nand U9665 (N_9665,N_8373,N_8350);
or U9666 (N_9666,N_8809,N_8463);
or U9667 (N_9667,N_8291,N_8833);
or U9668 (N_9668,N_8159,N_8008);
nor U9669 (N_9669,N_8564,N_8906);
xnor U9670 (N_9670,N_8828,N_8385);
or U9671 (N_9671,N_8833,N_8877);
xnor U9672 (N_9672,N_8418,N_8638);
nor U9673 (N_9673,N_8451,N_8136);
xnor U9674 (N_9674,N_8586,N_8337);
nor U9675 (N_9675,N_8714,N_8183);
nand U9676 (N_9676,N_8113,N_8922);
nor U9677 (N_9677,N_8982,N_8751);
and U9678 (N_9678,N_8297,N_8231);
nor U9679 (N_9679,N_8909,N_8540);
or U9680 (N_9680,N_8501,N_8239);
xnor U9681 (N_9681,N_8095,N_8270);
nand U9682 (N_9682,N_8958,N_8809);
nand U9683 (N_9683,N_8158,N_8376);
and U9684 (N_9684,N_8889,N_8268);
and U9685 (N_9685,N_8526,N_8410);
nand U9686 (N_9686,N_8472,N_8010);
nor U9687 (N_9687,N_8316,N_8215);
nor U9688 (N_9688,N_8316,N_8251);
or U9689 (N_9689,N_8319,N_8997);
nor U9690 (N_9690,N_8039,N_8440);
nor U9691 (N_9691,N_8419,N_8070);
nand U9692 (N_9692,N_8758,N_8152);
nor U9693 (N_9693,N_8719,N_8376);
or U9694 (N_9694,N_8271,N_8182);
and U9695 (N_9695,N_8729,N_8220);
or U9696 (N_9696,N_8632,N_8783);
nor U9697 (N_9697,N_8376,N_8922);
nor U9698 (N_9698,N_8438,N_8361);
nand U9699 (N_9699,N_8443,N_8051);
nor U9700 (N_9700,N_8276,N_8117);
nand U9701 (N_9701,N_8644,N_8175);
and U9702 (N_9702,N_8901,N_8500);
xnor U9703 (N_9703,N_8472,N_8361);
or U9704 (N_9704,N_8558,N_8251);
nor U9705 (N_9705,N_8467,N_8465);
nand U9706 (N_9706,N_8614,N_8988);
nor U9707 (N_9707,N_8950,N_8448);
nor U9708 (N_9708,N_8324,N_8638);
nor U9709 (N_9709,N_8376,N_8934);
nand U9710 (N_9710,N_8034,N_8917);
xnor U9711 (N_9711,N_8916,N_8392);
nor U9712 (N_9712,N_8660,N_8056);
nor U9713 (N_9713,N_8626,N_8803);
and U9714 (N_9714,N_8650,N_8508);
nor U9715 (N_9715,N_8925,N_8608);
nand U9716 (N_9716,N_8719,N_8048);
or U9717 (N_9717,N_8646,N_8312);
xnor U9718 (N_9718,N_8283,N_8083);
xnor U9719 (N_9719,N_8173,N_8797);
nand U9720 (N_9720,N_8172,N_8273);
and U9721 (N_9721,N_8026,N_8071);
xnor U9722 (N_9722,N_8951,N_8905);
and U9723 (N_9723,N_8925,N_8543);
xnor U9724 (N_9724,N_8245,N_8865);
nor U9725 (N_9725,N_8034,N_8427);
or U9726 (N_9726,N_8409,N_8794);
nand U9727 (N_9727,N_8459,N_8222);
nand U9728 (N_9728,N_8437,N_8760);
and U9729 (N_9729,N_8978,N_8223);
xor U9730 (N_9730,N_8101,N_8670);
nor U9731 (N_9731,N_8136,N_8208);
and U9732 (N_9732,N_8642,N_8990);
or U9733 (N_9733,N_8061,N_8408);
or U9734 (N_9734,N_8542,N_8927);
xnor U9735 (N_9735,N_8875,N_8381);
and U9736 (N_9736,N_8288,N_8465);
nand U9737 (N_9737,N_8109,N_8370);
and U9738 (N_9738,N_8380,N_8698);
nor U9739 (N_9739,N_8193,N_8270);
nor U9740 (N_9740,N_8821,N_8587);
or U9741 (N_9741,N_8937,N_8174);
nor U9742 (N_9742,N_8027,N_8969);
and U9743 (N_9743,N_8541,N_8314);
xor U9744 (N_9744,N_8774,N_8048);
xor U9745 (N_9745,N_8530,N_8217);
nor U9746 (N_9746,N_8713,N_8499);
or U9747 (N_9747,N_8505,N_8955);
nor U9748 (N_9748,N_8402,N_8214);
nand U9749 (N_9749,N_8754,N_8451);
xor U9750 (N_9750,N_8342,N_8542);
nor U9751 (N_9751,N_8604,N_8632);
xor U9752 (N_9752,N_8062,N_8429);
xnor U9753 (N_9753,N_8119,N_8758);
xor U9754 (N_9754,N_8249,N_8070);
xnor U9755 (N_9755,N_8699,N_8684);
nand U9756 (N_9756,N_8408,N_8675);
or U9757 (N_9757,N_8151,N_8878);
or U9758 (N_9758,N_8617,N_8270);
xnor U9759 (N_9759,N_8499,N_8152);
nor U9760 (N_9760,N_8911,N_8797);
xnor U9761 (N_9761,N_8743,N_8196);
xnor U9762 (N_9762,N_8400,N_8675);
nor U9763 (N_9763,N_8674,N_8773);
xor U9764 (N_9764,N_8068,N_8724);
nand U9765 (N_9765,N_8835,N_8895);
xnor U9766 (N_9766,N_8925,N_8071);
or U9767 (N_9767,N_8905,N_8115);
nand U9768 (N_9768,N_8362,N_8263);
or U9769 (N_9769,N_8259,N_8288);
or U9770 (N_9770,N_8079,N_8912);
xor U9771 (N_9771,N_8510,N_8632);
and U9772 (N_9772,N_8637,N_8755);
xor U9773 (N_9773,N_8277,N_8368);
or U9774 (N_9774,N_8668,N_8047);
and U9775 (N_9775,N_8675,N_8734);
or U9776 (N_9776,N_8302,N_8185);
xnor U9777 (N_9777,N_8635,N_8924);
nand U9778 (N_9778,N_8070,N_8347);
nand U9779 (N_9779,N_8660,N_8277);
xnor U9780 (N_9780,N_8346,N_8923);
xnor U9781 (N_9781,N_8919,N_8607);
nand U9782 (N_9782,N_8803,N_8260);
xnor U9783 (N_9783,N_8877,N_8874);
or U9784 (N_9784,N_8575,N_8119);
xnor U9785 (N_9785,N_8676,N_8309);
nand U9786 (N_9786,N_8329,N_8269);
and U9787 (N_9787,N_8377,N_8951);
xor U9788 (N_9788,N_8262,N_8284);
and U9789 (N_9789,N_8084,N_8485);
and U9790 (N_9790,N_8503,N_8032);
xor U9791 (N_9791,N_8568,N_8728);
and U9792 (N_9792,N_8471,N_8318);
nor U9793 (N_9793,N_8465,N_8122);
and U9794 (N_9794,N_8396,N_8602);
and U9795 (N_9795,N_8583,N_8693);
xnor U9796 (N_9796,N_8474,N_8152);
nand U9797 (N_9797,N_8158,N_8835);
nand U9798 (N_9798,N_8331,N_8945);
nor U9799 (N_9799,N_8910,N_8546);
xor U9800 (N_9800,N_8642,N_8194);
or U9801 (N_9801,N_8758,N_8148);
or U9802 (N_9802,N_8794,N_8561);
xnor U9803 (N_9803,N_8521,N_8266);
nor U9804 (N_9804,N_8542,N_8753);
or U9805 (N_9805,N_8320,N_8599);
or U9806 (N_9806,N_8414,N_8728);
nand U9807 (N_9807,N_8155,N_8266);
nor U9808 (N_9808,N_8599,N_8169);
xor U9809 (N_9809,N_8866,N_8213);
nand U9810 (N_9810,N_8336,N_8846);
xnor U9811 (N_9811,N_8213,N_8111);
nand U9812 (N_9812,N_8035,N_8628);
and U9813 (N_9813,N_8342,N_8743);
and U9814 (N_9814,N_8540,N_8956);
nor U9815 (N_9815,N_8491,N_8553);
and U9816 (N_9816,N_8291,N_8738);
nor U9817 (N_9817,N_8599,N_8290);
and U9818 (N_9818,N_8758,N_8981);
nor U9819 (N_9819,N_8774,N_8922);
and U9820 (N_9820,N_8903,N_8312);
xor U9821 (N_9821,N_8010,N_8764);
or U9822 (N_9822,N_8429,N_8367);
and U9823 (N_9823,N_8090,N_8833);
and U9824 (N_9824,N_8996,N_8765);
or U9825 (N_9825,N_8101,N_8429);
xor U9826 (N_9826,N_8818,N_8316);
and U9827 (N_9827,N_8852,N_8542);
nand U9828 (N_9828,N_8866,N_8028);
nor U9829 (N_9829,N_8217,N_8596);
or U9830 (N_9830,N_8138,N_8223);
nor U9831 (N_9831,N_8345,N_8946);
xor U9832 (N_9832,N_8224,N_8656);
nor U9833 (N_9833,N_8651,N_8602);
and U9834 (N_9834,N_8414,N_8026);
nor U9835 (N_9835,N_8244,N_8318);
or U9836 (N_9836,N_8122,N_8788);
or U9837 (N_9837,N_8491,N_8276);
nand U9838 (N_9838,N_8992,N_8213);
xor U9839 (N_9839,N_8848,N_8103);
and U9840 (N_9840,N_8266,N_8679);
nor U9841 (N_9841,N_8294,N_8416);
nand U9842 (N_9842,N_8834,N_8564);
or U9843 (N_9843,N_8913,N_8223);
xor U9844 (N_9844,N_8419,N_8363);
nand U9845 (N_9845,N_8419,N_8882);
nand U9846 (N_9846,N_8203,N_8916);
nor U9847 (N_9847,N_8296,N_8455);
or U9848 (N_9848,N_8576,N_8570);
nand U9849 (N_9849,N_8418,N_8190);
and U9850 (N_9850,N_8240,N_8810);
nor U9851 (N_9851,N_8844,N_8005);
nand U9852 (N_9852,N_8098,N_8194);
nor U9853 (N_9853,N_8670,N_8295);
and U9854 (N_9854,N_8201,N_8677);
or U9855 (N_9855,N_8790,N_8890);
nand U9856 (N_9856,N_8855,N_8811);
and U9857 (N_9857,N_8816,N_8839);
nor U9858 (N_9858,N_8076,N_8078);
and U9859 (N_9859,N_8613,N_8827);
or U9860 (N_9860,N_8695,N_8296);
or U9861 (N_9861,N_8489,N_8327);
or U9862 (N_9862,N_8005,N_8060);
xnor U9863 (N_9863,N_8394,N_8383);
nand U9864 (N_9864,N_8516,N_8742);
nand U9865 (N_9865,N_8418,N_8986);
nand U9866 (N_9866,N_8233,N_8291);
or U9867 (N_9867,N_8307,N_8578);
nor U9868 (N_9868,N_8933,N_8002);
xor U9869 (N_9869,N_8232,N_8608);
nand U9870 (N_9870,N_8237,N_8650);
nand U9871 (N_9871,N_8609,N_8085);
and U9872 (N_9872,N_8113,N_8772);
and U9873 (N_9873,N_8840,N_8435);
nand U9874 (N_9874,N_8424,N_8669);
xnor U9875 (N_9875,N_8954,N_8747);
nand U9876 (N_9876,N_8461,N_8133);
nor U9877 (N_9877,N_8129,N_8339);
nand U9878 (N_9878,N_8671,N_8453);
and U9879 (N_9879,N_8141,N_8547);
and U9880 (N_9880,N_8180,N_8362);
nor U9881 (N_9881,N_8144,N_8103);
or U9882 (N_9882,N_8038,N_8663);
or U9883 (N_9883,N_8134,N_8728);
nor U9884 (N_9884,N_8055,N_8549);
xor U9885 (N_9885,N_8202,N_8181);
and U9886 (N_9886,N_8061,N_8225);
nor U9887 (N_9887,N_8325,N_8186);
and U9888 (N_9888,N_8430,N_8056);
and U9889 (N_9889,N_8181,N_8017);
or U9890 (N_9890,N_8190,N_8723);
or U9891 (N_9891,N_8169,N_8834);
and U9892 (N_9892,N_8818,N_8874);
or U9893 (N_9893,N_8150,N_8802);
and U9894 (N_9894,N_8986,N_8212);
nand U9895 (N_9895,N_8590,N_8789);
or U9896 (N_9896,N_8384,N_8705);
nor U9897 (N_9897,N_8239,N_8740);
nor U9898 (N_9898,N_8545,N_8181);
and U9899 (N_9899,N_8609,N_8769);
nand U9900 (N_9900,N_8479,N_8063);
nand U9901 (N_9901,N_8363,N_8725);
nor U9902 (N_9902,N_8431,N_8849);
xnor U9903 (N_9903,N_8797,N_8594);
nand U9904 (N_9904,N_8803,N_8419);
xnor U9905 (N_9905,N_8385,N_8272);
nand U9906 (N_9906,N_8104,N_8348);
or U9907 (N_9907,N_8692,N_8162);
nand U9908 (N_9908,N_8872,N_8496);
xnor U9909 (N_9909,N_8494,N_8799);
or U9910 (N_9910,N_8292,N_8389);
or U9911 (N_9911,N_8378,N_8695);
xnor U9912 (N_9912,N_8693,N_8514);
and U9913 (N_9913,N_8053,N_8485);
and U9914 (N_9914,N_8858,N_8938);
and U9915 (N_9915,N_8628,N_8048);
nand U9916 (N_9916,N_8324,N_8019);
nor U9917 (N_9917,N_8526,N_8754);
xnor U9918 (N_9918,N_8327,N_8124);
or U9919 (N_9919,N_8735,N_8179);
or U9920 (N_9920,N_8889,N_8472);
and U9921 (N_9921,N_8838,N_8271);
or U9922 (N_9922,N_8143,N_8842);
xor U9923 (N_9923,N_8990,N_8730);
or U9924 (N_9924,N_8437,N_8494);
nand U9925 (N_9925,N_8408,N_8936);
xnor U9926 (N_9926,N_8090,N_8160);
nand U9927 (N_9927,N_8136,N_8290);
xor U9928 (N_9928,N_8456,N_8669);
or U9929 (N_9929,N_8470,N_8187);
xnor U9930 (N_9930,N_8022,N_8020);
nor U9931 (N_9931,N_8475,N_8254);
or U9932 (N_9932,N_8455,N_8386);
xnor U9933 (N_9933,N_8330,N_8911);
or U9934 (N_9934,N_8717,N_8294);
and U9935 (N_9935,N_8306,N_8738);
or U9936 (N_9936,N_8654,N_8644);
nand U9937 (N_9937,N_8739,N_8415);
xnor U9938 (N_9938,N_8907,N_8185);
and U9939 (N_9939,N_8438,N_8035);
and U9940 (N_9940,N_8734,N_8661);
nor U9941 (N_9941,N_8145,N_8844);
nor U9942 (N_9942,N_8908,N_8489);
and U9943 (N_9943,N_8067,N_8197);
or U9944 (N_9944,N_8250,N_8560);
and U9945 (N_9945,N_8261,N_8656);
xor U9946 (N_9946,N_8944,N_8734);
nor U9947 (N_9947,N_8647,N_8517);
and U9948 (N_9948,N_8788,N_8346);
nand U9949 (N_9949,N_8395,N_8117);
or U9950 (N_9950,N_8910,N_8308);
nand U9951 (N_9951,N_8716,N_8761);
and U9952 (N_9952,N_8603,N_8241);
nor U9953 (N_9953,N_8858,N_8142);
nor U9954 (N_9954,N_8284,N_8541);
nand U9955 (N_9955,N_8657,N_8495);
and U9956 (N_9956,N_8796,N_8480);
nor U9957 (N_9957,N_8272,N_8101);
xnor U9958 (N_9958,N_8938,N_8169);
or U9959 (N_9959,N_8949,N_8008);
nor U9960 (N_9960,N_8807,N_8328);
or U9961 (N_9961,N_8542,N_8162);
nor U9962 (N_9962,N_8778,N_8964);
or U9963 (N_9963,N_8704,N_8183);
nor U9964 (N_9964,N_8738,N_8381);
xor U9965 (N_9965,N_8240,N_8383);
nor U9966 (N_9966,N_8276,N_8131);
xnor U9967 (N_9967,N_8773,N_8344);
nand U9968 (N_9968,N_8422,N_8198);
xnor U9969 (N_9969,N_8582,N_8691);
and U9970 (N_9970,N_8548,N_8799);
nor U9971 (N_9971,N_8533,N_8316);
or U9972 (N_9972,N_8924,N_8492);
or U9973 (N_9973,N_8329,N_8484);
or U9974 (N_9974,N_8843,N_8117);
nand U9975 (N_9975,N_8017,N_8239);
nor U9976 (N_9976,N_8989,N_8169);
and U9977 (N_9977,N_8342,N_8788);
xnor U9978 (N_9978,N_8737,N_8568);
or U9979 (N_9979,N_8079,N_8045);
nor U9980 (N_9980,N_8900,N_8679);
nor U9981 (N_9981,N_8282,N_8051);
nor U9982 (N_9982,N_8197,N_8950);
or U9983 (N_9983,N_8870,N_8830);
or U9984 (N_9984,N_8357,N_8611);
or U9985 (N_9985,N_8519,N_8092);
xnor U9986 (N_9986,N_8075,N_8292);
or U9987 (N_9987,N_8755,N_8167);
xor U9988 (N_9988,N_8979,N_8164);
xnor U9989 (N_9989,N_8514,N_8451);
nand U9990 (N_9990,N_8115,N_8223);
or U9991 (N_9991,N_8714,N_8851);
nand U9992 (N_9992,N_8274,N_8557);
or U9993 (N_9993,N_8256,N_8836);
nand U9994 (N_9994,N_8957,N_8527);
and U9995 (N_9995,N_8379,N_8453);
and U9996 (N_9996,N_8740,N_8946);
nand U9997 (N_9997,N_8843,N_8651);
xnor U9998 (N_9998,N_8342,N_8995);
or U9999 (N_9999,N_8807,N_8414);
nor U10000 (N_10000,N_9420,N_9207);
xnor U10001 (N_10001,N_9561,N_9558);
nor U10002 (N_10002,N_9651,N_9368);
nor U10003 (N_10003,N_9168,N_9028);
nor U10004 (N_10004,N_9304,N_9442);
xor U10005 (N_10005,N_9091,N_9810);
and U10006 (N_10006,N_9332,N_9241);
nor U10007 (N_10007,N_9968,N_9783);
or U10008 (N_10008,N_9125,N_9223);
or U10009 (N_10009,N_9599,N_9699);
xnor U10010 (N_10010,N_9343,N_9197);
nand U10011 (N_10011,N_9250,N_9871);
or U10012 (N_10012,N_9855,N_9767);
and U10013 (N_10013,N_9696,N_9627);
nand U10014 (N_10014,N_9307,N_9615);
and U10015 (N_10015,N_9794,N_9977);
xnor U10016 (N_10016,N_9647,N_9576);
and U10017 (N_10017,N_9392,N_9879);
nor U10018 (N_10018,N_9349,N_9580);
xor U10019 (N_10019,N_9698,N_9920);
and U10020 (N_10020,N_9625,N_9875);
nor U10021 (N_10021,N_9406,N_9903);
nand U10022 (N_10022,N_9916,N_9876);
nand U10023 (N_10023,N_9531,N_9019);
nor U10024 (N_10024,N_9428,N_9693);
and U10025 (N_10025,N_9983,N_9537);
or U10026 (N_10026,N_9416,N_9085);
nor U10027 (N_10027,N_9723,N_9052);
nor U10028 (N_10028,N_9475,N_9710);
xnor U10029 (N_10029,N_9581,N_9287);
nand U10030 (N_10030,N_9954,N_9433);
or U10031 (N_10031,N_9787,N_9351);
and U10032 (N_10032,N_9186,N_9672);
and U10033 (N_10033,N_9275,N_9452);
or U10034 (N_10034,N_9214,N_9541);
and U10035 (N_10035,N_9515,N_9538);
and U10036 (N_10036,N_9098,N_9032);
nor U10037 (N_10037,N_9917,N_9593);
and U10038 (N_10038,N_9555,N_9260);
or U10039 (N_10039,N_9112,N_9825);
xor U10040 (N_10040,N_9634,N_9553);
or U10041 (N_10041,N_9901,N_9722);
and U10042 (N_10042,N_9739,N_9451);
xnor U10043 (N_10043,N_9549,N_9444);
nand U10044 (N_10044,N_9623,N_9161);
nor U10045 (N_10045,N_9743,N_9725);
xnor U10046 (N_10046,N_9193,N_9919);
or U10047 (N_10047,N_9545,N_9302);
nor U10048 (N_10048,N_9109,N_9745);
nand U10049 (N_10049,N_9323,N_9219);
xnor U10050 (N_10050,N_9014,N_9422);
xor U10051 (N_10051,N_9807,N_9746);
nand U10052 (N_10052,N_9866,N_9128);
nand U10053 (N_10053,N_9678,N_9359);
and U10054 (N_10054,N_9708,N_9820);
nor U10055 (N_10055,N_9024,N_9753);
nand U10056 (N_10056,N_9614,N_9873);
or U10057 (N_10057,N_9863,N_9700);
xnor U10058 (N_10058,N_9078,N_9652);
and U10059 (N_10059,N_9730,N_9832);
or U10060 (N_10060,N_9211,N_9813);
nor U10061 (N_10061,N_9377,N_9099);
or U10062 (N_10062,N_9675,N_9571);
or U10063 (N_10063,N_9791,N_9987);
or U10064 (N_10064,N_9591,N_9837);
and U10065 (N_10065,N_9643,N_9227);
and U10066 (N_10066,N_9347,N_9947);
or U10067 (N_10067,N_9117,N_9777);
and U10068 (N_10068,N_9311,N_9759);
and U10069 (N_10069,N_9847,N_9044);
and U10070 (N_10070,N_9528,N_9003);
nand U10071 (N_10071,N_9264,N_9862);
and U10072 (N_10072,N_9205,N_9185);
nand U10073 (N_10073,N_9828,N_9566);
nor U10074 (N_10074,N_9628,N_9718);
or U10075 (N_10075,N_9882,N_9105);
xor U10076 (N_10076,N_9291,N_9149);
xor U10077 (N_10077,N_9841,N_9738);
and U10078 (N_10078,N_9731,N_9846);
and U10079 (N_10079,N_9153,N_9575);
nand U10080 (N_10080,N_9023,N_9897);
nand U10081 (N_10081,N_9017,N_9221);
or U10082 (N_10082,N_9027,N_9001);
or U10083 (N_10083,N_9237,N_9450);
nor U10084 (N_10084,N_9512,N_9673);
xnor U10085 (N_10085,N_9865,N_9174);
or U10086 (N_10086,N_9621,N_9907);
nand U10087 (N_10087,N_9612,N_9732);
xor U10088 (N_10088,N_9329,N_9069);
or U10089 (N_10089,N_9034,N_9141);
and U10090 (N_10090,N_9856,N_9279);
and U10091 (N_10091,N_9140,N_9683);
and U10092 (N_10092,N_9939,N_9839);
and U10093 (N_10093,N_9529,N_9735);
xor U10094 (N_10094,N_9077,N_9640);
nor U10095 (N_10095,N_9579,N_9456);
nor U10096 (N_10096,N_9253,N_9251);
xor U10097 (N_10097,N_9570,N_9196);
nand U10098 (N_10098,N_9844,N_9244);
nand U10099 (N_10099,N_9543,N_9247);
nand U10100 (N_10100,N_9355,N_9995);
nor U10101 (N_10101,N_9022,N_9381);
nor U10102 (N_10102,N_9484,N_9997);
and U10103 (N_10103,N_9518,N_9124);
xor U10104 (N_10104,N_9478,N_9948);
nand U10105 (N_10105,N_9402,N_9333);
nor U10106 (N_10106,N_9962,N_9031);
nor U10107 (N_10107,N_9497,N_9938);
xor U10108 (N_10108,N_9177,N_9754);
nor U10109 (N_10109,N_9375,N_9799);
xnor U10110 (N_10110,N_9306,N_9602);
and U10111 (N_10111,N_9975,N_9976);
nor U10112 (N_10112,N_9138,N_9455);
and U10113 (N_10113,N_9814,N_9891);
nor U10114 (N_10114,N_9165,N_9559);
nor U10115 (N_10115,N_9180,N_9946);
xor U10116 (N_10116,N_9271,N_9812);
nor U10117 (N_10117,N_9396,N_9296);
nor U10118 (N_10118,N_9895,N_9702);
or U10119 (N_10119,N_9072,N_9586);
xnor U10120 (N_10120,N_9064,N_9273);
nor U10121 (N_10121,N_9148,N_9413);
and U10122 (N_10122,N_9073,N_9344);
xor U10123 (N_10123,N_9051,N_9904);
nand U10124 (N_10124,N_9945,N_9363);
and U10125 (N_10125,N_9386,N_9990);
nand U10126 (N_10126,N_9403,N_9494);
or U10127 (N_10127,N_9564,N_9927);
or U10128 (N_10128,N_9853,N_9009);
nand U10129 (N_10129,N_9719,N_9885);
nand U10130 (N_10130,N_9358,N_9802);
or U10131 (N_10131,N_9806,N_9395);
or U10132 (N_10132,N_9005,N_9058);
or U10133 (N_10133,N_9682,N_9274);
or U10134 (N_10134,N_9100,N_9957);
xnor U10135 (N_10135,N_9485,N_9330);
or U10136 (N_10136,N_9937,N_9991);
nand U10137 (N_10137,N_9025,N_9313);
or U10138 (N_10138,N_9061,N_9277);
xor U10139 (N_10139,N_9691,N_9546);
nor U10140 (N_10140,N_9134,N_9487);
or U10141 (N_10141,N_9522,N_9823);
and U10142 (N_10142,N_9793,N_9298);
and U10143 (N_10143,N_9638,N_9257);
xor U10144 (N_10144,N_9055,N_9163);
nand U10145 (N_10145,N_9026,N_9658);
nor U10146 (N_10146,N_9335,N_9889);
and U10147 (N_10147,N_9744,N_9039);
nor U10148 (N_10148,N_9690,N_9108);
nand U10149 (N_10149,N_9239,N_9974);
nand U10150 (N_10150,N_9784,N_9408);
nor U10151 (N_10151,N_9521,N_9076);
or U10152 (N_10152,N_9637,N_9910);
or U10153 (N_10153,N_9079,N_9902);
or U10154 (N_10154,N_9131,N_9648);
nor U10155 (N_10155,N_9129,N_9256);
nor U10156 (N_10156,N_9183,N_9817);
nor U10157 (N_10157,N_9081,N_9175);
nand U10158 (N_10158,N_9789,N_9655);
xor U10159 (N_10159,N_9797,N_9431);
xnor U10160 (N_10160,N_9988,N_9821);
nand U10161 (N_10161,N_9574,N_9914);
nand U10162 (N_10162,N_9785,N_9301);
xor U10163 (N_10163,N_9082,N_9912);
nor U10164 (N_10164,N_9636,N_9006);
nand U10165 (N_10165,N_9000,N_9146);
nand U10166 (N_10166,N_9049,N_9981);
and U10167 (N_10167,N_9373,N_9181);
xnor U10168 (N_10168,N_9860,N_9258);
nor U10169 (N_10169,N_9858,N_9387);
nor U10170 (N_10170,N_9116,N_9401);
nand U10171 (N_10171,N_9701,N_9065);
xor U10172 (N_10172,N_9519,N_9342);
and U10173 (N_10173,N_9805,N_9630);
nand U10174 (N_10174,N_9782,N_9070);
or U10175 (N_10175,N_9374,N_9463);
or U10176 (N_10176,N_9776,N_9419);
and U10177 (N_10177,N_9840,N_9246);
or U10178 (N_10178,N_9268,N_9763);
nor U10179 (N_10179,N_9182,N_9607);
and U10180 (N_10180,N_9911,N_9960);
xor U10181 (N_10181,N_9203,N_9404);
or U10182 (N_10182,N_9299,N_9908);
xnor U10183 (N_10183,N_9610,N_9712);
and U10184 (N_10184,N_9479,N_9978);
xnor U10185 (N_10185,N_9905,N_9235);
and U10186 (N_10186,N_9476,N_9276);
nand U10187 (N_10187,N_9290,N_9899);
nor U10188 (N_10188,N_9770,N_9795);
nand U10189 (N_10189,N_9715,N_9752);
and U10190 (N_10190,N_9362,N_9151);
nand U10191 (N_10191,N_9520,N_9315);
and U10192 (N_10192,N_9393,N_9861);
or U10193 (N_10193,N_9953,N_9798);
nor U10194 (N_10194,N_9540,N_9650);
or U10195 (N_10195,N_9616,N_9724);
and U10196 (N_10196,N_9043,N_9389);
nor U10197 (N_10197,N_9721,N_9378);
or U10198 (N_10198,N_9573,N_9316);
xnor U10199 (N_10199,N_9286,N_9191);
nand U10200 (N_10200,N_9132,N_9868);
nor U10201 (N_10201,N_9002,N_9517);
or U10202 (N_10202,N_9900,N_9471);
or U10203 (N_10203,N_9755,N_9461);
nand U10204 (N_10204,N_9762,N_9300);
and U10205 (N_10205,N_9880,N_9980);
or U10206 (N_10206,N_9166,N_9626);
nor U10207 (N_10207,N_9733,N_9004);
nor U10208 (N_10208,N_9350,N_9348);
xnor U10209 (N_10209,N_9040,N_9266);
and U10210 (N_10210,N_9356,N_9331);
nor U10211 (N_10211,N_9411,N_9303);
nor U10212 (N_10212,N_9936,N_9326);
nand U10213 (N_10213,N_9327,N_9262);
nor U10214 (N_10214,N_9989,N_9867);
and U10215 (N_10215,N_9322,N_9281);
and U10216 (N_10216,N_9737,N_9984);
nor U10217 (N_10217,N_9944,N_9265);
xor U10218 (N_10218,N_9489,N_9506);
or U10219 (N_10219,N_9152,N_9102);
xor U10220 (N_10220,N_9282,N_9680);
and U10221 (N_10221,N_9622,N_9749);
nor U10222 (N_10222,N_9457,N_9421);
nor U10223 (N_10223,N_9063,N_9534);
or U10224 (N_10224,N_9544,N_9585);
or U10225 (N_10225,N_9441,N_9269);
or U10226 (N_10226,N_9011,N_9928);
and U10227 (N_10227,N_9417,N_9226);
or U10228 (N_10228,N_9748,N_9964);
or U10229 (N_10229,N_9337,N_9971);
xor U10230 (N_10230,N_9649,N_9179);
or U10231 (N_10231,N_9458,N_9909);
nor U10232 (N_10232,N_9943,N_9554);
and U10233 (N_10233,N_9669,N_9781);
or U10234 (N_10234,N_9982,N_9493);
nand U10235 (N_10235,N_9569,N_9385);
or U10236 (N_10236,N_9836,N_9604);
and U10237 (N_10237,N_9926,N_9156);
and U10238 (N_10238,N_9229,N_9523);
nand U10239 (N_10239,N_9341,N_9923);
and U10240 (N_10240,N_9292,N_9764);
xor U10241 (N_10241,N_9309,N_9438);
xnor U10242 (N_10242,N_9881,N_9371);
nand U10243 (N_10243,N_9220,N_9532);
xor U10244 (N_10244,N_9288,N_9328);
xor U10245 (N_10245,N_9113,N_9560);
nor U10246 (N_10246,N_9896,N_9961);
and U10247 (N_10247,N_9418,N_9407);
xnor U10248 (N_10248,N_9225,N_9788);
and U10249 (N_10249,N_9635,N_9459);
nand U10250 (N_10250,N_9446,N_9503);
nor U10251 (N_10251,N_9619,N_9432);
and U10252 (N_10252,N_9270,N_9760);
xnor U10253 (N_10253,N_9436,N_9357);
xnor U10254 (N_10254,N_9206,N_9147);
and U10255 (N_10255,N_9854,N_9819);
nand U10256 (N_10256,N_9704,N_9103);
or U10257 (N_10257,N_9941,N_9222);
and U10258 (N_10258,N_9956,N_9369);
xnor U10259 (N_10259,N_9556,N_9178);
and U10260 (N_10260,N_9285,N_9720);
xor U10261 (N_10261,N_9567,N_9707);
xnor U10262 (N_10262,N_9066,N_9613);
or U10263 (N_10263,N_9790,N_9188);
nand U10264 (N_10264,N_9824,N_9490);
or U10265 (N_10265,N_9668,N_9167);
and U10266 (N_10266,N_9804,N_9979);
xor U10267 (N_10267,N_9123,N_9200);
and U10268 (N_10268,N_9843,N_9059);
nor U10269 (N_10269,N_9851,N_9925);
or U10270 (N_10270,N_9139,N_9194);
nand U10271 (N_10271,N_9596,N_9884);
xnor U10272 (N_10272,N_9931,N_9533);
or U10273 (N_10273,N_9671,N_9325);
xor U10274 (N_10274,N_9234,N_9486);
nor U10275 (N_10275,N_9453,N_9133);
nor U10276 (N_10276,N_9513,N_9029);
or U10277 (N_10277,N_9199,N_9670);
nor U10278 (N_10278,N_9992,N_9435);
nor U10279 (N_10279,N_9967,N_9826);
or U10280 (N_10280,N_9190,N_9773);
or U10281 (N_10281,N_9445,N_9477);
or U10282 (N_10282,N_9158,N_9539);
or U10283 (N_10283,N_9398,N_9423);
xnor U10284 (N_10284,N_9852,N_9189);
or U10285 (N_10285,N_9526,N_9632);
or U10286 (N_10286,N_9831,N_9611);
nand U10287 (N_10287,N_9624,N_9894);
xnor U10288 (N_10288,N_9424,N_9934);
xor U10289 (N_10289,N_9999,N_9481);
xor U10290 (N_10290,N_9815,N_9293);
and U10291 (N_10291,N_9890,N_9716);
or U10292 (N_10292,N_9259,N_9464);
nor U10293 (N_10293,N_9067,N_9500);
and U10294 (N_10294,N_9973,N_9448);
and U10295 (N_10295,N_9012,N_9473);
and U10296 (N_10296,N_9676,N_9434);
or U10297 (N_10297,N_9769,N_9405);
nor U10298 (N_10298,N_9187,N_9686);
xor U10299 (N_10299,N_9321,N_9958);
nor U10300 (N_10300,N_9157,N_9877);
and U10301 (N_10301,N_9491,N_9430);
or U10302 (N_10302,N_9425,N_9859);
xor U10303 (N_10303,N_9530,N_9587);
xor U10304 (N_10304,N_9050,N_9703);
xnor U10305 (N_10305,N_9060,N_9045);
nand U10306 (N_10306,N_9583,N_9106);
nor U10307 (N_10307,N_9524,N_9644);
xor U10308 (N_10308,N_9527,N_9935);
xnor U10309 (N_10309,N_9850,N_9808);
or U10310 (N_10310,N_9361,N_9071);
or U10311 (N_10311,N_9339,N_9366);
and U10312 (N_10312,N_9572,N_9792);
xnor U10313 (N_10313,N_9874,N_9849);
nor U10314 (N_10314,N_9209,N_9758);
and U10315 (N_10315,N_9390,N_9563);
or U10316 (N_10316,N_9388,N_9845);
nor U10317 (N_10317,N_9037,N_9728);
xnor U10318 (N_10318,N_9740,N_9483);
nand U10319 (N_10319,N_9940,N_9629);
nor U10320 (N_10320,N_9033,N_9775);
and U10321 (N_10321,N_9741,N_9231);
nand U10322 (N_10322,N_9516,N_9665);
nand U10323 (N_10323,N_9996,N_9352);
xnor U10324 (N_10324,N_9383,N_9713);
xnor U10325 (N_10325,N_9057,N_9122);
xor U10326 (N_10326,N_9312,N_9013);
xnor U10327 (N_10327,N_9089,N_9232);
nor U10328 (N_10328,N_9084,N_9319);
nand U10329 (N_10329,N_9667,N_9557);
nand U10330 (N_10330,N_9454,N_9310);
or U10331 (N_10331,N_9757,N_9460);
and U10332 (N_10332,N_9482,N_9094);
xor U10333 (N_10333,N_9075,N_9245);
nand U10334 (N_10334,N_9240,N_9261);
nor U10335 (N_10335,N_9663,N_9092);
or U10336 (N_10336,N_9093,N_9878);
nor U10337 (N_10337,N_9657,N_9169);
or U10338 (N_10338,N_9437,N_9466);
xor U10339 (N_10339,N_9150,N_9692);
xor U10340 (N_10340,N_9653,N_9771);
or U10341 (N_10341,N_9048,N_9121);
xnor U10342 (N_10342,N_9742,N_9525);
nand U10343 (N_10343,N_9848,N_9159);
xor U10344 (N_10344,N_9414,N_9394);
xnor U10345 (N_10345,N_9397,N_9086);
nor U10346 (N_10346,N_9143,N_9536);
and U10347 (N_10347,N_9210,N_9498);
xnor U10348 (N_10348,N_9320,N_9198);
and U10349 (N_10349,N_9830,N_9470);
nand U10350 (N_10350,N_9354,N_9765);
and U10351 (N_10351,N_9747,N_9694);
nor U10352 (N_10352,N_9508,N_9324);
nor U10353 (N_10353,N_9213,N_9184);
xnor U10354 (N_10354,N_9924,N_9509);
or U10355 (N_10355,N_9501,N_9510);
and U10356 (N_10356,N_9601,N_9308);
and U10357 (N_10357,N_9111,N_9443);
or U10358 (N_10358,N_9857,N_9228);
nand U10359 (N_10359,N_9780,N_9970);
xnor U10360 (N_10360,N_9986,N_9933);
and U10361 (N_10361,N_9047,N_9689);
or U10362 (N_10362,N_9969,N_9248);
or U10363 (N_10363,N_9215,N_9230);
xnor U10364 (N_10364,N_9447,N_9115);
nor U10365 (N_10365,N_9144,N_9212);
nor U10366 (N_10366,N_9609,N_9294);
xnor U10367 (N_10367,N_9993,N_9679);
xor U10368 (N_10368,N_9042,N_9550);
and U10369 (N_10369,N_9488,N_9734);
and U10370 (N_10370,N_9317,N_9062);
nand U10371 (N_10371,N_9097,N_9127);
or U10372 (N_10372,N_9864,N_9372);
or U10373 (N_10373,N_9041,N_9204);
xor U10374 (N_10374,N_9729,N_9822);
nor U10375 (N_10375,N_9499,N_9913);
or U10376 (N_10376,N_9681,N_9562);
or U10377 (N_10377,N_9620,N_9617);
xnor U10378 (N_10378,N_9380,N_9577);
and U10379 (N_10379,N_9496,N_9502);
nor U10380 (N_10380,N_9966,N_9829);
and U10381 (N_10381,N_9176,N_9136);
and U10382 (N_10382,N_9120,N_9535);
nand U10383 (N_10383,N_9376,N_9888);
or U10384 (N_10384,N_9467,N_9818);
and U10385 (N_10385,N_9353,N_9126);
xnor U10386 (N_10386,N_9095,N_9963);
xor U10387 (N_10387,N_9007,N_9932);
xor U10388 (N_10388,N_9654,N_9687);
and U10389 (N_10389,N_9118,N_9726);
nor U10390 (N_10390,N_9589,N_9192);
nor U10391 (N_10391,N_9018,N_9440);
or U10392 (N_10392,N_9751,N_9803);
xor U10393 (N_10393,N_9918,N_9314);
or U10394 (N_10394,N_9582,N_9409);
and U10395 (N_10395,N_9706,N_9170);
nand U10396 (N_10396,N_9838,N_9162);
nand U10397 (N_10397,N_9674,N_9284);
nor U10398 (N_10398,N_9505,N_9834);
and U10399 (N_10399,N_9297,N_9021);
and U10400 (N_10400,N_9243,N_9038);
and U10401 (N_10401,N_9603,N_9796);
and U10402 (N_10402,N_9208,N_9685);
nor U10403 (N_10403,N_9597,N_9272);
nor U10404 (N_10404,N_9468,N_9083);
nand U10405 (N_10405,N_9779,N_9252);
nand U10406 (N_10406,N_9036,N_9705);
or U10407 (N_10407,N_9160,N_9410);
nor U10408 (N_10408,N_9915,N_9449);
nand U10409 (N_10409,N_9255,N_9426);
nor U10410 (N_10410,N_9633,N_9233);
or U10411 (N_10411,N_9107,N_9594);
or U10412 (N_10412,N_9114,N_9631);
nand U10413 (N_10413,N_9346,N_9068);
xnor U10414 (N_10414,N_9427,N_9088);
xor U10415 (N_10415,N_9280,N_9588);
nand U10416 (N_10416,N_9659,N_9382);
nand U10417 (N_10417,N_9886,N_9090);
and U10418 (N_10418,N_9552,N_9736);
and U10419 (N_10419,N_9216,N_9469);
and U10420 (N_10420,N_9872,N_9642);
or U10421 (N_10421,N_9883,N_9278);
xor U10422 (N_10422,N_9930,N_9504);
nand U10423 (N_10423,N_9008,N_9786);
nor U10424 (N_10424,N_9869,N_9020);
and U10425 (N_10425,N_9336,N_9074);
nand U10426 (N_10426,N_9360,N_9495);
or U10427 (N_10427,N_9547,N_9365);
or U10428 (N_10428,N_9254,N_9507);
or U10429 (N_10429,N_9283,N_9661);
and U10430 (N_10430,N_9606,N_9994);
or U10431 (N_10431,N_9054,N_9816);
xnor U10432 (N_10432,N_9542,N_9898);
and U10433 (N_10433,N_9870,N_9155);
nor U10434 (N_10434,N_9046,N_9318);
or U10435 (N_10435,N_9384,N_9774);
xor U10436 (N_10436,N_9766,N_9289);
nand U10437 (N_10437,N_9010,N_9511);
or U10438 (N_10438,N_9202,N_9985);
nand U10439 (N_10439,N_9750,N_9201);
nor U10440 (N_10440,N_9101,N_9236);
and U10441 (N_10441,N_9639,N_9334);
or U10442 (N_10442,N_9242,N_9224);
nand U10443 (N_10443,N_9592,N_9605);
and U10444 (N_10444,N_9172,N_9772);
and U10445 (N_10445,N_9267,N_9811);
xor U10446 (N_10446,N_9835,N_9080);
xor U10447 (N_10447,N_9688,N_9548);
or U10448 (N_10448,N_9399,N_9087);
xor U10449 (N_10449,N_9660,N_9295);
xor U10450 (N_10450,N_9217,N_9514);
nand U10451 (N_10451,N_9218,N_9249);
nand U10452 (N_10452,N_9238,N_9130);
and U10453 (N_10453,N_9950,N_9697);
and U10454 (N_10454,N_9263,N_9415);
nand U10455 (N_10455,N_9015,N_9833);
or U10456 (N_10456,N_9664,N_9965);
nor U10457 (N_10457,N_9137,N_9590);
nor U10458 (N_10458,N_9104,N_9391);
or U10459 (N_10459,N_9778,N_9922);
nor U10460 (N_10460,N_9480,N_9662);
or U10461 (N_10461,N_9565,N_9584);
and U10462 (N_10462,N_9154,N_9600);
or U10463 (N_10463,N_9800,N_9016);
nand U10464 (N_10464,N_9711,N_9887);
nand U10465 (N_10465,N_9641,N_9465);
nand U10466 (N_10466,N_9809,N_9646);
nand U10467 (N_10467,N_9578,N_9598);
nand U10468 (N_10468,N_9717,N_9714);
and U10469 (N_10469,N_9952,N_9842);
and U10470 (N_10470,N_9608,N_9998);
xnor U10471 (N_10471,N_9893,N_9955);
nor U10472 (N_10472,N_9827,N_9709);
and U10473 (N_10473,N_9656,N_9801);
or U10474 (N_10474,N_9056,N_9756);
nand U10475 (N_10475,N_9951,N_9462);
nand U10476 (N_10476,N_9338,N_9035);
xor U10477 (N_10477,N_9684,N_9949);
or U10478 (N_10478,N_9340,N_9645);
or U10479 (N_10479,N_9727,N_9695);
and U10480 (N_10480,N_9959,N_9110);
nand U10481 (N_10481,N_9568,N_9768);
or U10482 (N_10482,N_9972,N_9474);
or U10483 (N_10483,N_9119,N_9921);
or U10484 (N_10484,N_9135,N_9364);
nand U10485 (N_10485,N_9439,N_9761);
nand U10486 (N_10486,N_9429,N_9142);
xnor U10487 (N_10487,N_9164,N_9096);
nand U10488 (N_10488,N_9677,N_9345);
xnor U10489 (N_10489,N_9492,N_9595);
or U10490 (N_10490,N_9906,N_9892);
and U10491 (N_10491,N_9472,N_9618);
and U10492 (N_10492,N_9171,N_9145);
nor U10493 (N_10493,N_9367,N_9173);
or U10494 (N_10494,N_9666,N_9551);
or U10495 (N_10495,N_9929,N_9030);
and U10496 (N_10496,N_9370,N_9379);
or U10497 (N_10497,N_9412,N_9195);
nor U10498 (N_10498,N_9305,N_9053);
nor U10499 (N_10499,N_9942,N_9400);
or U10500 (N_10500,N_9188,N_9958);
and U10501 (N_10501,N_9534,N_9005);
xnor U10502 (N_10502,N_9512,N_9078);
and U10503 (N_10503,N_9462,N_9322);
nor U10504 (N_10504,N_9620,N_9634);
xnor U10505 (N_10505,N_9493,N_9589);
and U10506 (N_10506,N_9142,N_9158);
or U10507 (N_10507,N_9195,N_9997);
and U10508 (N_10508,N_9589,N_9126);
xor U10509 (N_10509,N_9525,N_9864);
nor U10510 (N_10510,N_9597,N_9518);
nor U10511 (N_10511,N_9955,N_9168);
and U10512 (N_10512,N_9633,N_9297);
nand U10513 (N_10513,N_9914,N_9316);
nor U10514 (N_10514,N_9741,N_9496);
nor U10515 (N_10515,N_9692,N_9677);
or U10516 (N_10516,N_9620,N_9213);
or U10517 (N_10517,N_9697,N_9966);
or U10518 (N_10518,N_9898,N_9395);
or U10519 (N_10519,N_9215,N_9243);
nand U10520 (N_10520,N_9263,N_9805);
nor U10521 (N_10521,N_9316,N_9797);
xor U10522 (N_10522,N_9830,N_9682);
and U10523 (N_10523,N_9563,N_9603);
or U10524 (N_10524,N_9923,N_9336);
nand U10525 (N_10525,N_9238,N_9500);
nor U10526 (N_10526,N_9131,N_9751);
nand U10527 (N_10527,N_9943,N_9420);
xor U10528 (N_10528,N_9534,N_9402);
nor U10529 (N_10529,N_9056,N_9704);
nor U10530 (N_10530,N_9623,N_9860);
or U10531 (N_10531,N_9377,N_9517);
xor U10532 (N_10532,N_9595,N_9550);
nand U10533 (N_10533,N_9554,N_9041);
xor U10534 (N_10534,N_9256,N_9388);
or U10535 (N_10535,N_9806,N_9618);
nand U10536 (N_10536,N_9376,N_9719);
and U10537 (N_10537,N_9314,N_9517);
and U10538 (N_10538,N_9575,N_9805);
nand U10539 (N_10539,N_9191,N_9973);
nand U10540 (N_10540,N_9860,N_9692);
xnor U10541 (N_10541,N_9966,N_9830);
nand U10542 (N_10542,N_9434,N_9457);
nor U10543 (N_10543,N_9792,N_9912);
nor U10544 (N_10544,N_9948,N_9044);
nand U10545 (N_10545,N_9128,N_9581);
nand U10546 (N_10546,N_9063,N_9724);
xor U10547 (N_10547,N_9698,N_9400);
nand U10548 (N_10548,N_9477,N_9357);
xnor U10549 (N_10549,N_9037,N_9386);
or U10550 (N_10550,N_9194,N_9693);
nor U10551 (N_10551,N_9068,N_9403);
nor U10552 (N_10552,N_9753,N_9149);
nand U10553 (N_10553,N_9319,N_9192);
or U10554 (N_10554,N_9547,N_9320);
nor U10555 (N_10555,N_9369,N_9016);
xnor U10556 (N_10556,N_9604,N_9552);
nor U10557 (N_10557,N_9320,N_9977);
nand U10558 (N_10558,N_9970,N_9618);
and U10559 (N_10559,N_9998,N_9417);
nor U10560 (N_10560,N_9616,N_9271);
and U10561 (N_10561,N_9105,N_9659);
nand U10562 (N_10562,N_9000,N_9450);
nand U10563 (N_10563,N_9123,N_9887);
nor U10564 (N_10564,N_9019,N_9201);
and U10565 (N_10565,N_9056,N_9821);
nand U10566 (N_10566,N_9828,N_9958);
nand U10567 (N_10567,N_9428,N_9045);
or U10568 (N_10568,N_9903,N_9173);
nor U10569 (N_10569,N_9131,N_9982);
xor U10570 (N_10570,N_9701,N_9689);
nor U10571 (N_10571,N_9294,N_9457);
and U10572 (N_10572,N_9621,N_9660);
or U10573 (N_10573,N_9844,N_9346);
nand U10574 (N_10574,N_9201,N_9240);
and U10575 (N_10575,N_9995,N_9530);
nor U10576 (N_10576,N_9455,N_9480);
or U10577 (N_10577,N_9227,N_9499);
xnor U10578 (N_10578,N_9523,N_9025);
nor U10579 (N_10579,N_9466,N_9225);
nand U10580 (N_10580,N_9799,N_9020);
nor U10581 (N_10581,N_9670,N_9837);
nand U10582 (N_10582,N_9055,N_9365);
nor U10583 (N_10583,N_9139,N_9402);
or U10584 (N_10584,N_9526,N_9452);
xor U10585 (N_10585,N_9437,N_9974);
xor U10586 (N_10586,N_9645,N_9924);
or U10587 (N_10587,N_9445,N_9683);
and U10588 (N_10588,N_9404,N_9811);
and U10589 (N_10589,N_9991,N_9743);
nand U10590 (N_10590,N_9293,N_9207);
or U10591 (N_10591,N_9663,N_9065);
xnor U10592 (N_10592,N_9884,N_9686);
xnor U10593 (N_10593,N_9765,N_9348);
or U10594 (N_10594,N_9550,N_9543);
xor U10595 (N_10595,N_9726,N_9778);
nand U10596 (N_10596,N_9266,N_9270);
nand U10597 (N_10597,N_9832,N_9451);
nand U10598 (N_10598,N_9431,N_9716);
and U10599 (N_10599,N_9294,N_9889);
and U10600 (N_10600,N_9352,N_9076);
nand U10601 (N_10601,N_9149,N_9323);
nand U10602 (N_10602,N_9156,N_9031);
and U10603 (N_10603,N_9388,N_9957);
nand U10604 (N_10604,N_9268,N_9563);
or U10605 (N_10605,N_9927,N_9394);
xnor U10606 (N_10606,N_9591,N_9180);
xor U10607 (N_10607,N_9005,N_9506);
or U10608 (N_10608,N_9669,N_9797);
nand U10609 (N_10609,N_9890,N_9415);
xor U10610 (N_10610,N_9463,N_9575);
nor U10611 (N_10611,N_9601,N_9925);
and U10612 (N_10612,N_9410,N_9449);
xnor U10613 (N_10613,N_9813,N_9987);
xnor U10614 (N_10614,N_9588,N_9872);
and U10615 (N_10615,N_9375,N_9066);
xor U10616 (N_10616,N_9524,N_9676);
and U10617 (N_10617,N_9455,N_9500);
and U10618 (N_10618,N_9377,N_9539);
or U10619 (N_10619,N_9900,N_9082);
and U10620 (N_10620,N_9686,N_9349);
nor U10621 (N_10621,N_9334,N_9494);
or U10622 (N_10622,N_9425,N_9688);
xor U10623 (N_10623,N_9208,N_9686);
and U10624 (N_10624,N_9272,N_9385);
and U10625 (N_10625,N_9853,N_9544);
xor U10626 (N_10626,N_9086,N_9454);
and U10627 (N_10627,N_9939,N_9778);
or U10628 (N_10628,N_9546,N_9456);
and U10629 (N_10629,N_9591,N_9714);
nor U10630 (N_10630,N_9533,N_9575);
xnor U10631 (N_10631,N_9334,N_9275);
xnor U10632 (N_10632,N_9011,N_9063);
nor U10633 (N_10633,N_9360,N_9694);
or U10634 (N_10634,N_9202,N_9939);
xnor U10635 (N_10635,N_9132,N_9404);
or U10636 (N_10636,N_9390,N_9070);
and U10637 (N_10637,N_9289,N_9682);
nor U10638 (N_10638,N_9673,N_9449);
nor U10639 (N_10639,N_9453,N_9920);
xnor U10640 (N_10640,N_9796,N_9821);
xor U10641 (N_10641,N_9749,N_9782);
nand U10642 (N_10642,N_9494,N_9327);
xor U10643 (N_10643,N_9846,N_9551);
nor U10644 (N_10644,N_9960,N_9379);
and U10645 (N_10645,N_9169,N_9943);
nand U10646 (N_10646,N_9538,N_9739);
xnor U10647 (N_10647,N_9446,N_9760);
nand U10648 (N_10648,N_9092,N_9144);
or U10649 (N_10649,N_9231,N_9657);
xnor U10650 (N_10650,N_9609,N_9523);
or U10651 (N_10651,N_9222,N_9285);
nand U10652 (N_10652,N_9342,N_9914);
xnor U10653 (N_10653,N_9709,N_9019);
or U10654 (N_10654,N_9676,N_9224);
or U10655 (N_10655,N_9462,N_9117);
nor U10656 (N_10656,N_9695,N_9928);
nand U10657 (N_10657,N_9996,N_9391);
nand U10658 (N_10658,N_9081,N_9226);
nor U10659 (N_10659,N_9947,N_9231);
nand U10660 (N_10660,N_9296,N_9552);
or U10661 (N_10661,N_9198,N_9359);
nand U10662 (N_10662,N_9918,N_9989);
and U10663 (N_10663,N_9452,N_9668);
or U10664 (N_10664,N_9574,N_9178);
nor U10665 (N_10665,N_9892,N_9210);
nand U10666 (N_10666,N_9272,N_9781);
nand U10667 (N_10667,N_9764,N_9754);
or U10668 (N_10668,N_9482,N_9921);
nand U10669 (N_10669,N_9666,N_9008);
nor U10670 (N_10670,N_9473,N_9292);
nor U10671 (N_10671,N_9675,N_9209);
and U10672 (N_10672,N_9205,N_9761);
xor U10673 (N_10673,N_9528,N_9048);
xnor U10674 (N_10674,N_9789,N_9408);
xor U10675 (N_10675,N_9574,N_9552);
and U10676 (N_10676,N_9031,N_9808);
nor U10677 (N_10677,N_9707,N_9317);
nor U10678 (N_10678,N_9265,N_9632);
nand U10679 (N_10679,N_9427,N_9094);
nor U10680 (N_10680,N_9813,N_9775);
xor U10681 (N_10681,N_9970,N_9982);
or U10682 (N_10682,N_9815,N_9531);
xnor U10683 (N_10683,N_9902,N_9142);
or U10684 (N_10684,N_9035,N_9592);
nor U10685 (N_10685,N_9177,N_9601);
nor U10686 (N_10686,N_9690,N_9954);
nor U10687 (N_10687,N_9269,N_9816);
nor U10688 (N_10688,N_9338,N_9604);
xor U10689 (N_10689,N_9875,N_9532);
and U10690 (N_10690,N_9924,N_9882);
and U10691 (N_10691,N_9021,N_9416);
nor U10692 (N_10692,N_9847,N_9845);
or U10693 (N_10693,N_9361,N_9666);
and U10694 (N_10694,N_9057,N_9652);
nor U10695 (N_10695,N_9034,N_9024);
and U10696 (N_10696,N_9098,N_9368);
or U10697 (N_10697,N_9680,N_9018);
and U10698 (N_10698,N_9060,N_9069);
or U10699 (N_10699,N_9062,N_9788);
and U10700 (N_10700,N_9932,N_9199);
or U10701 (N_10701,N_9174,N_9496);
xnor U10702 (N_10702,N_9201,N_9649);
nor U10703 (N_10703,N_9278,N_9809);
xnor U10704 (N_10704,N_9508,N_9248);
and U10705 (N_10705,N_9652,N_9732);
and U10706 (N_10706,N_9444,N_9742);
xnor U10707 (N_10707,N_9483,N_9183);
and U10708 (N_10708,N_9162,N_9566);
xor U10709 (N_10709,N_9569,N_9823);
or U10710 (N_10710,N_9363,N_9922);
nor U10711 (N_10711,N_9043,N_9346);
xor U10712 (N_10712,N_9477,N_9338);
nand U10713 (N_10713,N_9352,N_9903);
nor U10714 (N_10714,N_9298,N_9552);
or U10715 (N_10715,N_9358,N_9025);
and U10716 (N_10716,N_9336,N_9033);
nand U10717 (N_10717,N_9988,N_9959);
xnor U10718 (N_10718,N_9672,N_9602);
xor U10719 (N_10719,N_9493,N_9597);
nor U10720 (N_10720,N_9644,N_9566);
or U10721 (N_10721,N_9222,N_9042);
nand U10722 (N_10722,N_9160,N_9257);
or U10723 (N_10723,N_9565,N_9381);
or U10724 (N_10724,N_9439,N_9606);
nand U10725 (N_10725,N_9973,N_9334);
and U10726 (N_10726,N_9903,N_9524);
nor U10727 (N_10727,N_9880,N_9270);
or U10728 (N_10728,N_9889,N_9298);
or U10729 (N_10729,N_9233,N_9427);
nand U10730 (N_10730,N_9217,N_9962);
or U10731 (N_10731,N_9727,N_9059);
and U10732 (N_10732,N_9277,N_9568);
xor U10733 (N_10733,N_9521,N_9182);
nand U10734 (N_10734,N_9317,N_9976);
nand U10735 (N_10735,N_9067,N_9111);
xnor U10736 (N_10736,N_9540,N_9853);
or U10737 (N_10737,N_9979,N_9201);
nor U10738 (N_10738,N_9123,N_9810);
and U10739 (N_10739,N_9505,N_9987);
xor U10740 (N_10740,N_9167,N_9383);
and U10741 (N_10741,N_9482,N_9674);
nor U10742 (N_10742,N_9445,N_9450);
nand U10743 (N_10743,N_9770,N_9354);
or U10744 (N_10744,N_9738,N_9432);
and U10745 (N_10745,N_9522,N_9892);
xor U10746 (N_10746,N_9914,N_9528);
xnor U10747 (N_10747,N_9181,N_9624);
nand U10748 (N_10748,N_9853,N_9471);
xnor U10749 (N_10749,N_9632,N_9975);
nor U10750 (N_10750,N_9892,N_9499);
nor U10751 (N_10751,N_9343,N_9935);
and U10752 (N_10752,N_9218,N_9777);
or U10753 (N_10753,N_9383,N_9774);
or U10754 (N_10754,N_9686,N_9975);
nand U10755 (N_10755,N_9474,N_9319);
nand U10756 (N_10756,N_9657,N_9604);
xor U10757 (N_10757,N_9719,N_9797);
nand U10758 (N_10758,N_9794,N_9052);
nand U10759 (N_10759,N_9595,N_9452);
nor U10760 (N_10760,N_9360,N_9697);
xnor U10761 (N_10761,N_9448,N_9134);
nand U10762 (N_10762,N_9470,N_9342);
or U10763 (N_10763,N_9565,N_9133);
nor U10764 (N_10764,N_9503,N_9591);
nand U10765 (N_10765,N_9395,N_9883);
or U10766 (N_10766,N_9248,N_9466);
nand U10767 (N_10767,N_9467,N_9652);
nand U10768 (N_10768,N_9052,N_9611);
xnor U10769 (N_10769,N_9223,N_9345);
nor U10770 (N_10770,N_9660,N_9186);
nor U10771 (N_10771,N_9487,N_9957);
or U10772 (N_10772,N_9045,N_9149);
xor U10773 (N_10773,N_9797,N_9461);
or U10774 (N_10774,N_9635,N_9963);
nor U10775 (N_10775,N_9449,N_9075);
or U10776 (N_10776,N_9177,N_9167);
xor U10777 (N_10777,N_9151,N_9353);
nand U10778 (N_10778,N_9676,N_9694);
nand U10779 (N_10779,N_9417,N_9145);
xor U10780 (N_10780,N_9125,N_9603);
xnor U10781 (N_10781,N_9669,N_9025);
and U10782 (N_10782,N_9993,N_9490);
nor U10783 (N_10783,N_9262,N_9103);
xnor U10784 (N_10784,N_9293,N_9757);
and U10785 (N_10785,N_9344,N_9581);
and U10786 (N_10786,N_9897,N_9501);
and U10787 (N_10787,N_9820,N_9451);
nand U10788 (N_10788,N_9784,N_9358);
nand U10789 (N_10789,N_9597,N_9675);
and U10790 (N_10790,N_9056,N_9162);
and U10791 (N_10791,N_9510,N_9033);
nor U10792 (N_10792,N_9060,N_9837);
xor U10793 (N_10793,N_9154,N_9462);
xor U10794 (N_10794,N_9779,N_9960);
nor U10795 (N_10795,N_9196,N_9424);
or U10796 (N_10796,N_9811,N_9882);
and U10797 (N_10797,N_9788,N_9790);
and U10798 (N_10798,N_9717,N_9319);
nand U10799 (N_10799,N_9334,N_9715);
xor U10800 (N_10800,N_9815,N_9647);
xor U10801 (N_10801,N_9868,N_9612);
or U10802 (N_10802,N_9118,N_9253);
nor U10803 (N_10803,N_9021,N_9590);
and U10804 (N_10804,N_9774,N_9419);
nand U10805 (N_10805,N_9030,N_9414);
xor U10806 (N_10806,N_9008,N_9374);
or U10807 (N_10807,N_9645,N_9879);
or U10808 (N_10808,N_9924,N_9944);
xnor U10809 (N_10809,N_9477,N_9722);
nand U10810 (N_10810,N_9812,N_9869);
nand U10811 (N_10811,N_9300,N_9328);
nand U10812 (N_10812,N_9992,N_9390);
or U10813 (N_10813,N_9883,N_9675);
xnor U10814 (N_10814,N_9269,N_9628);
nor U10815 (N_10815,N_9054,N_9303);
nand U10816 (N_10816,N_9188,N_9139);
nor U10817 (N_10817,N_9120,N_9176);
and U10818 (N_10818,N_9016,N_9398);
nor U10819 (N_10819,N_9387,N_9248);
nand U10820 (N_10820,N_9921,N_9589);
nand U10821 (N_10821,N_9123,N_9576);
nand U10822 (N_10822,N_9361,N_9704);
and U10823 (N_10823,N_9033,N_9709);
and U10824 (N_10824,N_9003,N_9352);
xnor U10825 (N_10825,N_9068,N_9955);
and U10826 (N_10826,N_9692,N_9588);
or U10827 (N_10827,N_9649,N_9512);
nor U10828 (N_10828,N_9385,N_9701);
and U10829 (N_10829,N_9971,N_9063);
and U10830 (N_10830,N_9498,N_9591);
nand U10831 (N_10831,N_9576,N_9594);
nor U10832 (N_10832,N_9753,N_9189);
nor U10833 (N_10833,N_9551,N_9977);
nor U10834 (N_10834,N_9116,N_9258);
and U10835 (N_10835,N_9292,N_9834);
or U10836 (N_10836,N_9164,N_9392);
xor U10837 (N_10837,N_9584,N_9931);
or U10838 (N_10838,N_9124,N_9376);
xnor U10839 (N_10839,N_9084,N_9135);
nor U10840 (N_10840,N_9079,N_9631);
nor U10841 (N_10841,N_9391,N_9926);
xnor U10842 (N_10842,N_9230,N_9126);
and U10843 (N_10843,N_9331,N_9982);
xnor U10844 (N_10844,N_9117,N_9072);
and U10845 (N_10845,N_9410,N_9279);
xor U10846 (N_10846,N_9882,N_9322);
and U10847 (N_10847,N_9191,N_9563);
xor U10848 (N_10848,N_9834,N_9673);
and U10849 (N_10849,N_9183,N_9945);
nor U10850 (N_10850,N_9215,N_9036);
or U10851 (N_10851,N_9727,N_9871);
xnor U10852 (N_10852,N_9555,N_9992);
nor U10853 (N_10853,N_9803,N_9175);
nand U10854 (N_10854,N_9785,N_9363);
nor U10855 (N_10855,N_9887,N_9521);
or U10856 (N_10856,N_9975,N_9966);
xnor U10857 (N_10857,N_9612,N_9138);
nor U10858 (N_10858,N_9263,N_9008);
or U10859 (N_10859,N_9500,N_9051);
nand U10860 (N_10860,N_9159,N_9886);
xnor U10861 (N_10861,N_9069,N_9009);
and U10862 (N_10862,N_9560,N_9157);
xnor U10863 (N_10863,N_9161,N_9282);
and U10864 (N_10864,N_9272,N_9106);
nor U10865 (N_10865,N_9274,N_9303);
xor U10866 (N_10866,N_9802,N_9130);
nand U10867 (N_10867,N_9176,N_9313);
or U10868 (N_10868,N_9644,N_9103);
nand U10869 (N_10869,N_9020,N_9155);
xor U10870 (N_10870,N_9636,N_9236);
or U10871 (N_10871,N_9559,N_9011);
or U10872 (N_10872,N_9928,N_9390);
nand U10873 (N_10873,N_9978,N_9653);
or U10874 (N_10874,N_9151,N_9550);
or U10875 (N_10875,N_9315,N_9087);
and U10876 (N_10876,N_9498,N_9519);
xor U10877 (N_10877,N_9875,N_9491);
nor U10878 (N_10878,N_9900,N_9196);
nand U10879 (N_10879,N_9145,N_9630);
and U10880 (N_10880,N_9219,N_9380);
xor U10881 (N_10881,N_9548,N_9492);
nor U10882 (N_10882,N_9242,N_9080);
xor U10883 (N_10883,N_9805,N_9563);
nand U10884 (N_10884,N_9390,N_9167);
and U10885 (N_10885,N_9757,N_9039);
nor U10886 (N_10886,N_9419,N_9560);
xnor U10887 (N_10887,N_9351,N_9309);
nand U10888 (N_10888,N_9228,N_9478);
nand U10889 (N_10889,N_9440,N_9947);
xnor U10890 (N_10890,N_9282,N_9983);
nand U10891 (N_10891,N_9525,N_9895);
nand U10892 (N_10892,N_9955,N_9060);
nand U10893 (N_10893,N_9753,N_9029);
and U10894 (N_10894,N_9689,N_9563);
or U10895 (N_10895,N_9355,N_9536);
and U10896 (N_10896,N_9279,N_9390);
or U10897 (N_10897,N_9276,N_9692);
xor U10898 (N_10898,N_9437,N_9764);
or U10899 (N_10899,N_9753,N_9823);
xnor U10900 (N_10900,N_9476,N_9987);
or U10901 (N_10901,N_9891,N_9713);
nand U10902 (N_10902,N_9622,N_9575);
and U10903 (N_10903,N_9213,N_9850);
or U10904 (N_10904,N_9378,N_9643);
nand U10905 (N_10905,N_9954,N_9979);
and U10906 (N_10906,N_9374,N_9688);
or U10907 (N_10907,N_9070,N_9308);
or U10908 (N_10908,N_9689,N_9346);
or U10909 (N_10909,N_9940,N_9878);
nand U10910 (N_10910,N_9528,N_9329);
xor U10911 (N_10911,N_9428,N_9175);
nand U10912 (N_10912,N_9838,N_9038);
nand U10913 (N_10913,N_9315,N_9016);
xor U10914 (N_10914,N_9451,N_9567);
nand U10915 (N_10915,N_9775,N_9276);
or U10916 (N_10916,N_9398,N_9322);
nand U10917 (N_10917,N_9922,N_9985);
or U10918 (N_10918,N_9358,N_9965);
nor U10919 (N_10919,N_9997,N_9938);
nand U10920 (N_10920,N_9309,N_9025);
nand U10921 (N_10921,N_9853,N_9581);
nand U10922 (N_10922,N_9568,N_9257);
or U10923 (N_10923,N_9216,N_9100);
and U10924 (N_10924,N_9355,N_9096);
xor U10925 (N_10925,N_9718,N_9331);
nor U10926 (N_10926,N_9384,N_9258);
and U10927 (N_10927,N_9858,N_9973);
nand U10928 (N_10928,N_9681,N_9425);
or U10929 (N_10929,N_9616,N_9161);
nand U10930 (N_10930,N_9855,N_9345);
nor U10931 (N_10931,N_9909,N_9989);
nor U10932 (N_10932,N_9336,N_9904);
xor U10933 (N_10933,N_9187,N_9562);
or U10934 (N_10934,N_9895,N_9715);
nor U10935 (N_10935,N_9008,N_9169);
nand U10936 (N_10936,N_9880,N_9467);
and U10937 (N_10937,N_9368,N_9944);
nor U10938 (N_10938,N_9378,N_9418);
and U10939 (N_10939,N_9098,N_9363);
nand U10940 (N_10940,N_9352,N_9481);
or U10941 (N_10941,N_9442,N_9897);
or U10942 (N_10942,N_9330,N_9523);
xor U10943 (N_10943,N_9117,N_9857);
nand U10944 (N_10944,N_9237,N_9451);
or U10945 (N_10945,N_9820,N_9288);
or U10946 (N_10946,N_9989,N_9232);
xnor U10947 (N_10947,N_9610,N_9810);
xor U10948 (N_10948,N_9201,N_9554);
and U10949 (N_10949,N_9427,N_9447);
nand U10950 (N_10950,N_9096,N_9491);
and U10951 (N_10951,N_9170,N_9633);
xor U10952 (N_10952,N_9930,N_9416);
nand U10953 (N_10953,N_9602,N_9455);
and U10954 (N_10954,N_9314,N_9651);
xor U10955 (N_10955,N_9962,N_9514);
nand U10956 (N_10956,N_9519,N_9893);
xnor U10957 (N_10957,N_9161,N_9588);
and U10958 (N_10958,N_9556,N_9125);
nor U10959 (N_10959,N_9503,N_9811);
xor U10960 (N_10960,N_9024,N_9475);
nor U10961 (N_10961,N_9578,N_9142);
or U10962 (N_10962,N_9498,N_9388);
nor U10963 (N_10963,N_9954,N_9085);
or U10964 (N_10964,N_9160,N_9229);
or U10965 (N_10965,N_9126,N_9509);
nand U10966 (N_10966,N_9540,N_9775);
or U10967 (N_10967,N_9160,N_9458);
or U10968 (N_10968,N_9269,N_9352);
nor U10969 (N_10969,N_9258,N_9263);
and U10970 (N_10970,N_9382,N_9405);
or U10971 (N_10971,N_9381,N_9129);
nand U10972 (N_10972,N_9560,N_9589);
or U10973 (N_10973,N_9396,N_9922);
nand U10974 (N_10974,N_9285,N_9374);
nand U10975 (N_10975,N_9049,N_9218);
and U10976 (N_10976,N_9458,N_9952);
nor U10977 (N_10977,N_9096,N_9077);
nand U10978 (N_10978,N_9052,N_9838);
and U10979 (N_10979,N_9518,N_9956);
nor U10980 (N_10980,N_9061,N_9372);
and U10981 (N_10981,N_9647,N_9626);
and U10982 (N_10982,N_9644,N_9669);
nand U10983 (N_10983,N_9383,N_9033);
nor U10984 (N_10984,N_9302,N_9228);
xor U10985 (N_10985,N_9302,N_9271);
xor U10986 (N_10986,N_9107,N_9595);
and U10987 (N_10987,N_9143,N_9723);
nor U10988 (N_10988,N_9777,N_9201);
xor U10989 (N_10989,N_9374,N_9010);
or U10990 (N_10990,N_9665,N_9511);
or U10991 (N_10991,N_9078,N_9619);
or U10992 (N_10992,N_9289,N_9922);
nand U10993 (N_10993,N_9782,N_9178);
nor U10994 (N_10994,N_9657,N_9835);
xor U10995 (N_10995,N_9092,N_9808);
and U10996 (N_10996,N_9508,N_9789);
and U10997 (N_10997,N_9338,N_9077);
or U10998 (N_10998,N_9299,N_9463);
nor U10999 (N_10999,N_9346,N_9193);
nor U11000 (N_11000,N_10075,N_10052);
xnor U11001 (N_11001,N_10005,N_10679);
xnor U11002 (N_11002,N_10788,N_10066);
xnor U11003 (N_11003,N_10069,N_10212);
nand U11004 (N_11004,N_10874,N_10503);
xnor U11005 (N_11005,N_10269,N_10281);
xor U11006 (N_11006,N_10932,N_10665);
nand U11007 (N_11007,N_10782,N_10222);
nand U11008 (N_11008,N_10636,N_10850);
nand U11009 (N_11009,N_10260,N_10012);
xnor U11010 (N_11010,N_10629,N_10225);
or U11011 (N_11011,N_10266,N_10504);
or U11012 (N_11012,N_10578,N_10904);
xor U11013 (N_11013,N_10599,N_10735);
xnor U11014 (N_11014,N_10179,N_10477);
xor U11015 (N_11015,N_10660,N_10466);
or U11016 (N_11016,N_10505,N_10417);
or U11017 (N_11017,N_10536,N_10923);
or U11018 (N_11018,N_10635,N_10241);
or U11019 (N_11019,N_10166,N_10007);
xor U11020 (N_11020,N_10998,N_10018);
and U11021 (N_11021,N_10667,N_10813);
nand U11022 (N_11022,N_10529,N_10887);
nand U11023 (N_11023,N_10458,N_10375);
nand U11024 (N_11024,N_10471,N_10893);
or U11025 (N_11025,N_10791,N_10221);
xnor U11026 (N_11026,N_10767,N_10470);
xor U11027 (N_11027,N_10848,N_10950);
or U11028 (N_11028,N_10934,N_10806);
or U11029 (N_11029,N_10803,N_10755);
or U11030 (N_11030,N_10410,N_10734);
or U11031 (N_11031,N_10634,N_10334);
and U11032 (N_11032,N_10015,N_10844);
xor U11033 (N_11033,N_10406,N_10078);
nand U11034 (N_11034,N_10652,N_10176);
and U11035 (N_11035,N_10839,N_10303);
and U11036 (N_11036,N_10983,N_10374);
nand U11037 (N_11037,N_10698,N_10645);
or U11038 (N_11038,N_10008,N_10832);
nand U11039 (N_11039,N_10656,N_10242);
xnor U11040 (N_11040,N_10521,N_10684);
xor U11041 (N_11041,N_10963,N_10984);
xnor U11042 (N_11042,N_10270,N_10366);
xor U11043 (N_11043,N_10863,N_10830);
nor U11044 (N_11044,N_10921,N_10423);
or U11045 (N_11045,N_10319,N_10740);
xor U11046 (N_11046,N_10165,N_10610);
xor U11047 (N_11047,N_10535,N_10388);
xnor U11048 (N_11048,N_10870,N_10168);
or U11049 (N_11049,N_10231,N_10025);
and U11050 (N_11050,N_10373,N_10886);
nand U11051 (N_11051,N_10455,N_10418);
nand U11052 (N_11052,N_10939,N_10871);
and U11053 (N_11053,N_10064,N_10948);
xnor U11054 (N_11054,N_10172,N_10632);
or U11055 (N_11055,N_10031,N_10764);
nand U11056 (N_11056,N_10738,N_10262);
and U11057 (N_11057,N_10872,N_10710);
xnor U11058 (N_11058,N_10343,N_10603);
xor U11059 (N_11059,N_10726,N_10279);
nor U11060 (N_11060,N_10670,N_10256);
nand U11061 (N_11061,N_10962,N_10092);
nor U11062 (N_11062,N_10058,N_10902);
nor U11063 (N_11063,N_10822,N_10054);
xor U11064 (N_11064,N_10158,N_10719);
xnor U11065 (N_11065,N_10145,N_10416);
or U11066 (N_11066,N_10879,N_10237);
and U11067 (N_11067,N_10690,N_10481);
nor U11068 (N_11068,N_10633,N_10233);
xor U11069 (N_11069,N_10271,N_10508);
nand U11070 (N_11070,N_10510,N_10011);
xor U11071 (N_11071,N_10713,N_10286);
nand U11072 (N_11072,N_10506,N_10261);
and U11073 (N_11073,N_10197,N_10894);
xnor U11074 (N_11074,N_10252,N_10802);
and U11075 (N_11075,N_10640,N_10370);
nand U11076 (N_11076,N_10982,N_10105);
nor U11077 (N_11077,N_10084,N_10760);
nand U11078 (N_11078,N_10428,N_10680);
and U11079 (N_11079,N_10593,N_10773);
nor U11080 (N_11080,N_10947,N_10193);
xor U11081 (N_11081,N_10924,N_10573);
nor U11082 (N_11082,N_10461,N_10407);
and U11083 (N_11083,N_10930,N_10309);
nor U11084 (N_11084,N_10562,N_10707);
nand U11085 (N_11085,N_10293,N_10780);
nand U11086 (N_11086,N_10208,N_10553);
nand U11087 (N_11087,N_10459,N_10519);
or U11088 (N_11088,N_10327,N_10202);
or U11089 (N_11089,N_10322,N_10487);
or U11090 (N_11090,N_10475,N_10490);
nand U11091 (N_11091,N_10751,N_10859);
and U11092 (N_11092,N_10037,N_10446);
and U11093 (N_11093,N_10558,N_10958);
or U11094 (N_11094,N_10686,N_10841);
xor U11095 (N_11095,N_10729,N_10439);
or U11096 (N_11096,N_10612,N_10127);
and U11097 (N_11097,N_10986,N_10400);
and U11098 (N_11098,N_10047,N_10706);
or U11099 (N_11099,N_10150,N_10170);
and U11100 (N_11100,N_10689,N_10067);
xnor U11101 (N_11101,N_10071,N_10700);
and U11102 (N_11102,N_10912,N_10372);
nor U11103 (N_11103,N_10673,N_10033);
xnor U11104 (N_11104,N_10595,N_10659);
nor U11105 (N_11105,N_10026,N_10332);
nor U11106 (N_11106,N_10027,N_10435);
or U11107 (N_11107,N_10929,N_10385);
xor U11108 (N_11108,N_10325,N_10393);
nor U11109 (N_11109,N_10587,N_10377);
nor U11110 (N_11110,N_10720,N_10215);
or U11111 (N_11111,N_10885,N_10901);
or U11112 (N_11112,N_10248,N_10449);
nand U11113 (N_11113,N_10541,N_10837);
nor U11114 (N_11114,N_10216,N_10081);
and U11115 (N_11115,N_10364,N_10961);
xor U11116 (N_11116,N_10232,N_10443);
nand U11117 (N_11117,N_10224,N_10928);
or U11118 (N_11118,N_10509,N_10711);
xnor U11119 (N_11119,N_10151,N_10049);
nor U11120 (N_11120,N_10174,N_10565);
or U11121 (N_11121,N_10144,N_10997);
nor U11122 (N_11122,N_10717,N_10588);
nor U11123 (N_11123,N_10688,N_10655);
or U11124 (N_11124,N_10055,N_10491);
and U11125 (N_11125,N_10826,N_10810);
or U11126 (N_11126,N_10793,N_10537);
or U11127 (N_11127,N_10605,N_10299);
nor U11128 (N_11128,N_10157,N_10315);
and U11129 (N_11129,N_10563,N_10978);
or U11130 (N_11130,N_10001,N_10692);
or U11131 (N_11131,N_10265,N_10163);
or U11132 (N_11132,N_10219,N_10792);
nand U11133 (N_11133,N_10228,N_10161);
xnor U11134 (N_11134,N_10906,N_10080);
or U11135 (N_11135,N_10354,N_10359);
and U11136 (N_11136,N_10355,N_10728);
and U11137 (N_11137,N_10852,N_10577);
or U11138 (N_11138,N_10630,N_10429);
and U11139 (N_11139,N_10290,N_10936);
nand U11140 (N_11140,N_10646,N_10824);
nor U11141 (N_11141,N_10651,N_10213);
nand U11142 (N_11142,N_10444,N_10474);
nand U11143 (N_11143,N_10827,N_10494);
xnor U11144 (N_11144,N_10095,N_10387);
or U11145 (N_11145,N_10568,N_10989);
nand U11146 (N_11146,N_10153,N_10101);
nor U11147 (N_11147,N_10549,N_10668);
nor U11148 (N_11148,N_10324,N_10203);
nand U11149 (N_11149,N_10142,N_10909);
or U11150 (N_11150,N_10292,N_10583);
xor U11151 (N_11151,N_10102,N_10194);
nor U11152 (N_11152,N_10952,N_10951);
or U11153 (N_11153,N_10479,N_10701);
and U11154 (N_11154,N_10123,N_10496);
nor U11155 (N_11155,N_10762,N_10169);
xnor U11156 (N_11156,N_10083,N_10524);
nor U11157 (N_11157,N_10516,N_10278);
and U11158 (N_11158,N_10484,N_10148);
nor U11159 (N_11159,N_10189,N_10235);
or U11160 (N_11160,N_10079,N_10747);
xnor U11161 (N_11161,N_10511,N_10274);
nand U11162 (N_11162,N_10009,N_10816);
xnor U11163 (N_11163,N_10333,N_10472);
or U11164 (N_11164,N_10677,N_10838);
or U11165 (N_11165,N_10335,N_10920);
and U11166 (N_11166,N_10399,N_10575);
or U11167 (N_11167,N_10528,N_10768);
nor U11168 (N_11168,N_10899,N_10182);
nor U11169 (N_11169,N_10386,N_10908);
and U11170 (N_11170,N_10103,N_10187);
or U11171 (N_11171,N_10088,N_10674);
nor U11172 (N_11172,N_10514,N_10363);
nand U11173 (N_11173,N_10561,N_10229);
nand U11174 (N_11174,N_10462,N_10425);
xor U11175 (N_11175,N_10448,N_10905);
and U11176 (N_11176,N_10382,N_10115);
nand U11177 (N_11177,N_10135,N_10916);
or U11178 (N_11178,N_10704,N_10815);
nand U11179 (N_11179,N_10727,N_10104);
or U11180 (N_11180,N_10041,N_10703);
nand U11181 (N_11181,N_10849,N_10451);
or U11182 (N_11182,N_10938,N_10730);
and U11183 (N_11183,N_10970,N_10831);
nand U11184 (N_11184,N_10570,N_10507);
and U11185 (N_11185,N_10132,N_10356);
nand U11186 (N_11186,N_10898,N_10137);
and U11187 (N_11187,N_10096,N_10757);
nand U11188 (N_11188,N_10206,N_10620);
or U11189 (N_11189,N_10533,N_10149);
nand U11190 (N_11190,N_10238,N_10403);
xor U11191 (N_11191,N_10427,N_10090);
or U11192 (N_11192,N_10006,N_10124);
nor U11193 (N_11193,N_10609,N_10942);
nand U11194 (N_11194,N_10990,N_10236);
xor U11195 (N_11195,N_10050,N_10596);
nor U11196 (N_11196,N_10136,N_10489);
and U11197 (N_11197,N_10846,N_10348);
and U11198 (N_11198,N_10051,N_10621);
nor U11199 (N_11199,N_10664,N_10336);
nor U11200 (N_11200,N_10540,N_10211);
nor U11201 (N_11201,N_10809,N_10777);
and U11202 (N_11202,N_10941,N_10944);
nand U11203 (N_11203,N_10914,N_10736);
and U11204 (N_11204,N_10087,N_10833);
xor U11205 (N_11205,N_10666,N_10116);
nand U11206 (N_11206,N_10010,N_10878);
nand U11207 (N_11207,N_10074,N_10807);
xor U11208 (N_11208,N_10152,N_10129);
nor U11209 (N_11209,N_10209,N_10714);
xnor U11210 (N_11210,N_10973,N_10880);
and U11211 (N_11211,N_10766,N_10121);
and U11212 (N_11212,N_10744,N_10441);
and U11213 (N_11213,N_10367,N_10369);
or U11214 (N_11214,N_10126,N_10955);
nor U11215 (N_11215,N_10404,N_10437);
or U11216 (N_11216,N_10550,N_10527);
and U11217 (N_11217,N_10845,N_10625);
and U11218 (N_11218,N_10752,N_10316);
nor U11219 (N_11219,N_10042,N_10089);
xor U11220 (N_11220,N_10731,N_10113);
or U11221 (N_11221,N_10285,N_10086);
or U11222 (N_11222,N_10927,N_10284);
nand U11223 (N_11223,N_10606,N_10053);
nand U11224 (N_11224,N_10781,N_10882);
or U11225 (N_11225,N_10300,N_10681);
nand U11226 (N_11226,N_10709,N_10812);
nor U11227 (N_11227,N_10226,N_10493);
xnor U11228 (N_11228,N_10177,N_10987);
nor U11229 (N_11229,N_10118,N_10301);
nand U11230 (N_11230,N_10994,N_10028);
nor U11231 (N_11231,N_10227,N_10992);
xor U11232 (N_11232,N_10492,N_10522);
nand U11233 (N_11233,N_10384,N_10305);
nand U11234 (N_11234,N_10184,N_10530);
and U11235 (N_11235,N_10964,N_10753);
or U11236 (N_11236,N_10122,N_10217);
and U11237 (N_11237,N_10501,N_10949);
nand U11238 (N_11238,N_10467,N_10682);
and U11239 (N_11239,N_10624,N_10817);
or U11240 (N_11240,N_10016,N_10555);
xnor U11241 (N_11241,N_10304,N_10342);
nor U11242 (N_11242,N_10314,N_10943);
nor U11243 (N_11243,N_10068,N_10945);
and U11244 (N_11244,N_10552,N_10060);
xnor U11245 (N_11245,N_10035,N_10450);
xnor U11246 (N_11246,N_10130,N_10974);
xnor U11247 (N_11247,N_10985,N_10750);
or U11248 (N_11248,N_10043,N_10523);
nor U11249 (N_11249,N_10705,N_10685);
xor U11250 (N_11250,N_10862,N_10725);
nor U11251 (N_11251,N_10557,N_10447);
xor U11252 (N_11252,N_10210,N_10323);
xor U11253 (N_11253,N_10259,N_10585);
and U11254 (N_11254,N_10469,N_10650);
nand U11255 (N_11255,N_10953,N_10412);
or U11256 (N_11256,N_10046,N_10631);
xnor U11257 (N_11257,N_10861,N_10133);
xnor U11258 (N_11258,N_10485,N_10560);
nand U11259 (N_11259,N_10057,N_10676);
xor U11260 (N_11260,N_10254,N_10162);
and U11261 (N_11261,N_10828,N_10933);
nor U11262 (N_11262,N_10107,N_10351);
and U11263 (N_11263,N_10935,N_10897);
and U11264 (N_11264,N_10072,N_10967);
nand U11265 (N_11265,N_10240,N_10787);
nor U11266 (N_11266,N_10622,N_10062);
nand U11267 (N_11267,N_10192,N_10772);
nor U11268 (N_11268,N_10272,N_10979);
xor U11269 (N_11269,N_10498,N_10742);
and U11270 (N_11270,N_10581,N_10662);
xnor U11271 (N_11271,N_10821,N_10854);
nand U11272 (N_11272,N_10675,N_10312);
nand U11273 (N_11273,N_10545,N_10413);
nor U11274 (N_11274,N_10584,N_10737);
xor U11275 (N_11275,N_10977,N_10805);
xnor U11276 (N_11276,N_10340,N_10649);
nand U11277 (N_11277,N_10289,N_10098);
or U11278 (N_11278,N_10420,N_10716);
nor U11279 (N_11279,N_10065,N_10036);
or U11280 (N_11280,N_10980,N_10070);
nor U11281 (N_11281,N_10154,N_10601);
nand U11282 (N_11282,N_10432,N_10889);
nor U11283 (N_11283,N_10811,N_10185);
nor U11284 (N_11284,N_10480,N_10464);
xor U11285 (N_11285,N_10627,N_10171);
and U11286 (N_11286,N_10564,N_10347);
nor U11287 (N_11287,N_10532,N_10223);
nand U11288 (N_11288,N_10460,N_10250);
nand U11289 (N_11289,N_10294,N_10454);
nor U11290 (N_11290,N_10296,N_10547);
nand U11291 (N_11291,N_10275,N_10257);
and U11292 (N_11292,N_10199,N_10453);
or U11293 (N_11293,N_10867,N_10117);
and U11294 (N_11294,N_10181,N_10981);
nor U11295 (N_11295,N_10770,N_10842);
nand U11296 (N_11296,N_10186,N_10253);
or U11297 (N_11297,N_10038,N_10851);
nor U11298 (N_11298,N_10648,N_10543);
nand U11299 (N_11299,N_10834,N_10797);
nand U11300 (N_11300,N_10436,N_10799);
or U11301 (N_11301,N_10167,N_10566);
nor U11302 (N_11302,N_10247,N_10869);
nor U11303 (N_11303,N_10311,N_10741);
nand U11304 (N_11304,N_10972,N_10919);
nor U11305 (N_11305,N_10531,N_10749);
xor U11306 (N_11306,N_10892,N_10559);
or U11307 (N_11307,N_10891,N_10754);
xor U11308 (N_11308,N_10338,N_10112);
nor U11309 (N_11309,N_10804,N_10903);
and U11310 (N_11310,N_10263,N_10695);
or U11311 (N_11311,N_10258,N_10672);
and U11312 (N_11312,N_10108,N_10383);
nor U11313 (N_11313,N_10654,N_10877);
nor U11314 (N_11314,N_10623,N_10534);
and U11315 (N_11315,N_10794,N_10442);
nand U11316 (N_11316,N_10282,N_10991);
xor U11317 (N_11317,N_10765,N_10718);
and U11318 (N_11318,N_10093,N_10954);
and U11319 (N_11319,N_10800,N_10307);
nor U11320 (N_11320,N_10776,N_10313);
or U11321 (N_11321,N_10440,N_10337);
nand U11322 (N_11322,N_10497,N_10708);
nand U11323 (N_11323,N_10361,N_10733);
or U11324 (N_11324,N_10180,N_10795);
nor U11325 (N_11325,N_10789,N_10607);
nor U11326 (N_11326,N_10959,N_10995);
and U11327 (N_11327,N_10106,N_10330);
nor U11328 (N_11328,N_10756,N_10156);
and U11329 (N_11329,N_10518,N_10389);
nor U11330 (N_11330,N_10683,N_10138);
xor U11331 (N_11331,N_10976,N_10234);
nor U11332 (N_11332,N_10020,N_10395);
or U11333 (N_11333,N_10539,N_10191);
xor U11334 (N_11334,N_10456,N_10380);
nand U11335 (N_11335,N_10888,N_10918);
nand U11336 (N_11336,N_10993,N_10975);
nor U11337 (N_11337,N_10567,N_10111);
and U11338 (N_11338,N_10019,N_10840);
and U11339 (N_11339,N_10590,N_10002);
or U11340 (N_11340,N_10843,N_10243);
or U11341 (N_11341,N_10743,N_10207);
nand U11342 (N_11342,N_10045,N_10426);
nor U11343 (N_11343,N_10349,N_10239);
or U11344 (N_11344,N_10452,N_10589);
and U11345 (N_11345,N_10597,N_10819);
nor U11346 (N_11346,N_10966,N_10771);
nand U11347 (N_11347,N_10661,N_10960);
and U11348 (N_11348,N_10619,N_10702);
nor U11349 (N_11349,N_10611,N_10814);
xor U11350 (N_11350,N_10044,N_10723);
xor U11351 (N_11351,N_10353,N_10774);
xor U11352 (N_11352,N_10626,N_10745);
nor U11353 (N_11353,N_10200,N_10542);
or U11354 (N_11354,N_10937,N_10628);
xor U11355 (N_11355,N_10957,N_10178);
or U11356 (N_11356,N_10000,N_10173);
nor U11357 (N_11357,N_10120,N_10415);
xnor U11358 (N_11358,N_10582,N_10586);
nand U11359 (N_11359,N_10280,N_10687);
nand U11360 (N_11360,N_10783,N_10820);
nand U11361 (N_11361,N_10097,N_10344);
and U11362 (N_11362,N_10457,N_10183);
xor U11363 (N_11363,N_10571,N_10671);
xor U11364 (N_11364,N_10004,N_10779);
and U11365 (N_11365,N_10617,N_10288);
nor U11366 (N_11366,N_10056,N_10155);
nor U11367 (N_11367,N_10317,N_10268);
xor U11368 (N_11368,N_10297,N_10357);
and U11369 (N_11369,N_10500,N_10273);
and U11370 (N_11370,N_10775,N_10143);
nand U11371 (N_11371,N_10604,N_10085);
or U11372 (N_11372,N_10579,N_10956);
nor U11373 (N_11373,N_10131,N_10034);
xor U11374 (N_11374,N_10580,N_10411);
nor U11375 (N_11375,N_10022,N_10146);
nand U11376 (N_11376,N_10855,N_10048);
nor U11377 (N_11377,N_10678,N_10551);
nor U11378 (N_11378,N_10875,N_10401);
and U11379 (N_11379,N_10402,N_10638);
nand U11380 (N_11380,N_10341,N_10915);
xnor U11381 (N_11381,N_10653,N_10544);
and U11382 (N_11382,N_10040,N_10134);
and U11383 (N_11383,N_10431,N_10201);
nand U11384 (N_11384,N_10438,N_10911);
or U11385 (N_11385,N_10077,N_10109);
xor U11386 (N_11386,N_10548,N_10287);
and U11387 (N_11387,N_10013,N_10023);
nand U11388 (N_11388,N_10881,N_10414);
nand U11389 (N_11389,N_10345,N_10785);
or U11390 (N_11390,N_10128,N_10784);
and U11391 (N_11391,N_10091,N_10613);
or U11392 (N_11392,N_10251,N_10430);
and U11393 (N_11393,N_10396,N_10864);
xnor U11394 (N_11394,N_10073,N_10796);
xor U11395 (N_11395,N_10318,N_10245);
or U11396 (N_11396,N_10499,N_10835);
and U11397 (N_11397,N_10482,N_10378);
nand U11398 (N_11398,N_10669,N_10546);
or U11399 (N_11399,N_10473,N_10032);
and U11400 (N_11400,N_10836,N_10913);
or U11401 (N_11401,N_10119,N_10647);
nand U11402 (N_11402,N_10295,N_10159);
nand U11403 (N_11403,N_10657,N_10569);
nor U11404 (N_11404,N_10890,N_10868);
xor U11405 (N_11405,N_10424,N_10847);
or U11406 (N_11406,N_10576,N_10866);
nor U11407 (N_11407,N_10030,N_10512);
xor U11408 (N_11408,N_10398,N_10615);
or U11409 (N_11409,N_10059,N_10362);
or U11410 (N_11410,N_10465,N_10003);
or U11411 (N_11411,N_10476,N_10488);
nand U11412 (N_11412,N_10188,N_10264);
and U11413 (N_11413,N_10759,N_10405);
xor U11414 (N_11414,N_10365,N_10922);
and U11415 (N_11415,N_10926,N_10198);
xnor U11416 (N_11416,N_10358,N_10526);
nor U11417 (N_11417,N_10592,N_10147);
nor U11418 (N_11418,N_10790,N_10220);
or U11419 (N_11419,N_10376,N_10715);
nand U11420 (N_11420,N_10538,N_10408);
nor U11421 (N_11421,N_10644,N_10965);
nand U11422 (N_11422,N_10371,N_10988);
or U11423 (N_11423,N_10691,N_10230);
nor U11424 (N_11424,N_10391,N_10291);
nor U11425 (N_11425,N_10808,N_10298);
xor U11426 (N_11426,N_10495,N_10463);
or U11427 (N_11427,N_10468,N_10190);
and U11428 (N_11428,N_10277,N_10856);
xor U11429 (N_11429,N_10699,N_10876);
and U11430 (N_11430,N_10602,N_10255);
or U11431 (N_11431,N_10572,N_10419);
and U11432 (N_11432,N_10829,N_10663);
xnor U11433 (N_11433,N_10642,N_10125);
xnor U11434 (N_11434,N_10598,N_10249);
or U11435 (N_11435,N_10818,N_10082);
nand U11436 (N_11436,N_10825,N_10141);
and U11437 (N_11437,N_10798,N_10515);
or U11438 (N_11438,N_10017,N_10917);
and U11439 (N_11439,N_10326,N_10712);
nor U11440 (N_11440,N_10339,N_10860);
or U11441 (N_11441,N_10556,N_10641);
and U11442 (N_11442,N_10946,N_10276);
nor U11443 (N_11443,N_10308,N_10352);
and U11444 (N_11444,N_10999,N_10608);
nand U11445 (N_11445,N_10024,N_10346);
and U11446 (N_11446,N_10968,N_10328);
xnor U11447 (N_11447,N_10196,N_10204);
or U11448 (N_11448,N_10761,N_10483);
and U11449 (N_11449,N_10940,N_10513);
or U11450 (N_11450,N_10160,N_10021);
nand U11451 (N_11451,N_10591,N_10724);
nor U11452 (N_11452,N_10397,N_10360);
nor U11453 (N_11453,N_10076,N_10693);
nand U11454 (N_11454,N_10883,N_10320);
nand U11455 (N_11455,N_10267,N_10637);
nand U11456 (N_11456,N_10858,N_10329);
xnor U11457 (N_11457,N_10525,N_10422);
and U11458 (N_11458,N_10421,N_10907);
nand U11459 (N_11459,N_10574,N_10218);
nor U11460 (N_11460,N_10639,N_10094);
xor U11461 (N_11461,N_10971,N_10321);
and U11462 (N_11462,N_10786,N_10896);
nor U11463 (N_11463,N_10643,N_10925);
xor U11464 (N_11464,N_10394,N_10502);
and U11465 (N_11465,N_10114,N_10658);
or U11466 (N_11466,N_10381,N_10873);
or U11467 (N_11467,N_10368,N_10618);
xnor U11468 (N_11468,N_10616,N_10769);
xor U11469 (N_11469,N_10110,N_10517);
nand U11470 (N_11470,N_10306,N_10246);
or U11471 (N_11471,N_10748,N_10694);
or U11472 (N_11472,N_10721,N_10746);
nor U11473 (N_11473,N_10520,N_10486);
nor U11474 (N_11474,N_10433,N_10350);
nand U11475 (N_11475,N_10139,N_10283);
or U11476 (N_11476,N_10823,N_10801);
or U11477 (N_11477,N_10910,N_10445);
nand U11478 (N_11478,N_10600,N_10039);
or U11479 (N_11479,N_10732,N_10205);
xnor U11480 (N_11480,N_10696,N_10214);
and U11481 (N_11481,N_10063,N_10778);
nor U11482 (N_11482,N_10164,N_10739);
xnor U11483 (N_11483,N_10554,N_10931);
and U11484 (N_11484,N_10853,N_10900);
xor U11485 (N_11485,N_10969,N_10884);
xnor U11486 (N_11486,N_10244,N_10175);
or U11487 (N_11487,N_10722,N_10697);
nand U11488 (N_11488,N_10310,N_10014);
nand U11489 (N_11489,N_10331,N_10594);
xnor U11490 (N_11490,N_10478,N_10857);
nand U11491 (N_11491,N_10392,N_10758);
nand U11492 (N_11492,N_10099,N_10029);
and U11493 (N_11493,N_10996,N_10434);
xor U11494 (N_11494,N_10140,N_10763);
nand U11495 (N_11495,N_10379,N_10614);
or U11496 (N_11496,N_10061,N_10390);
nor U11497 (N_11497,N_10409,N_10865);
or U11498 (N_11498,N_10895,N_10100);
nand U11499 (N_11499,N_10302,N_10195);
and U11500 (N_11500,N_10931,N_10165);
xnor U11501 (N_11501,N_10684,N_10513);
xor U11502 (N_11502,N_10347,N_10852);
and U11503 (N_11503,N_10626,N_10020);
nor U11504 (N_11504,N_10389,N_10732);
nor U11505 (N_11505,N_10536,N_10332);
xor U11506 (N_11506,N_10736,N_10867);
or U11507 (N_11507,N_10934,N_10562);
nor U11508 (N_11508,N_10719,N_10879);
nand U11509 (N_11509,N_10625,N_10060);
xor U11510 (N_11510,N_10258,N_10838);
and U11511 (N_11511,N_10731,N_10728);
or U11512 (N_11512,N_10629,N_10011);
nand U11513 (N_11513,N_10597,N_10006);
nand U11514 (N_11514,N_10893,N_10847);
or U11515 (N_11515,N_10338,N_10787);
nand U11516 (N_11516,N_10479,N_10858);
xor U11517 (N_11517,N_10406,N_10057);
nand U11518 (N_11518,N_10193,N_10430);
nor U11519 (N_11519,N_10301,N_10349);
or U11520 (N_11520,N_10105,N_10382);
nand U11521 (N_11521,N_10638,N_10481);
nand U11522 (N_11522,N_10647,N_10159);
xor U11523 (N_11523,N_10156,N_10042);
nor U11524 (N_11524,N_10643,N_10920);
xor U11525 (N_11525,N_10510,N_10320);
nor U11526 (N_11526,N_10391,N_10913);
or U11527 (N_11527,N_10812,N_10150);
xnor U11528 (N_11528,N_10582,N_10439);
or U11529 (N_11529,N_10791,N_10949);
or U11530 (N_11530,N_10533,N_10067);
nor U11531 (N_11531,N_10712,N_10570);
xor U11532 (N_11532,N_10296,N_10154);
and U11533 (N_11533,N_10544,N_10055);
or U11534 (N_11534,N_10708,N_10054);
and U11535 (N_11535,N_10418,N_10672);
nor U11536 (N_11536,N_10574,N_10532);
or U11537 (N_11537,N_10884,N_10816);
nor U11538 (N_11538,N_10997,N_10099);
nand U11539 (N_11539,N_10962,N_10890);
and U11540 (N_11540,N_10984,N_10705);
nor U11541 (N_11541,N_10878,N_10264);
xor U11542 (N_11542,N_10882,N_10618);
xnor U11543 (N_11543,N_10954,N_10621);
or U11544 (N_11544,N_10903,N_10885);
nand U11545 (N_11545,N_10209,N_10973);
or U11546 (N_11546,N_10700,N_10087);
and U11547 (N_11547,N_10767,N_10353);
xnor U11548 (N_11548,N_10270,N_10012);
nor U11549 (N_11549,N_10923,N_10653);
or U11550 (N_11550,N_10964,N_10553);
and U11551 (N_11551,N_10229,N_10462);
or U11552 (N_11552,N_10960,N_10615);
or U11553 (N_11553,N_10545,N_10721);
and U11554 (N_11554,N_10986,N_10301);
xor U11555 (N_11555,N_10884,N_10510);
or U11556 (N_11556,N_10571,N_10257);
nor U11557 (N_11557,N_10346,N_10700);
nor U11558 (N_11558,N_10748,N_10030);
or U11559 (N_11559,N_10047,N_10906);
or U11560 (N_11560,N_10769,N_10943);
and U11561 (N_11561,N_10766,N_10889);
or U11562 (N_11562,N_10060,N_10197);
nand U11563 (N_11563,N_10953,N_10929);
xnor U11564 (N_11564,N_10849,N_10045);
and U11565 (N_11565,N_10697,N_10526);
xnor U11566 (N_11566,N_10651,N_10828);
nand U11567 (N_11567,N_10811,N_10222);
nand U11568 (N_11568,N_10094,N_10857);
and U11569 (N_11569,N_10721,N_10438);
or U11570 (N_11570,N_10669,N_10629);
nand U11571 (N_11571,N_10832,N_10705);
or U11572 (N_11572,N_10868,N_10844);
nor U11573 (N_11573,N_10751,N_10672);
nand U11574 (N_11574,N_10911,N_10804);
nor U11575 (N_11575,N_10074,N_10632);
xor U11576 (N_11576,N_10296,N_10026);
nand U11577 (N_11577,N_10672,N_10769);
xor U11578 (N_11578,N_10550,N_10646);
nor U11579 (N_11579,N_10961,N_10075);
nand U11580 (N_11580,N_10054,N_10811);
xor U11581 (N_11581,N_10191,N_10659);
nand U11582 (N_11582,N_10555,N_10812);
nor U11583 (N_11583,N_10710,N_10037);
xnor U11584 (N_11584,N_10242,N_10064);
xnor U11585 (N_11585,N_10826,N_10157);
or U11586 (N_11586,N_10106,N_10913);
nand U11587 (N_11587,N_10232,N_10600);
nor U11588 (N_11588,N_10131,N_10560);
nor U11589 (N_11589,N_10569,N_10565);
and U11590 (N_11590,N_10099,N_10273);
and U11591 (N_11591,N_10393,N_10948);
and U11592 (N_11592,N_10889,N_10869);
or U11593 (N_11593,N_10199,N_10331);
nand U11594 (N_11594,N_10242,N_10989);
nand U11595 (N_11595,N_10930,N_10506);
or U11596 (N_11596,N_10109,N_10551);
nand U11597 (N_11597,N_10370,N_10782);
nor U11598 (N_11598,N_10764,N_10435);
and U11599 (N_11599,N_10055,N_10589);
or U11600 (N_11600,N_10706,N_10882);
xor U11601 (N_11601,N_10273,N_10666);
nand U11602 (N_11602,N_10842,N_10689);
xor U11603 (N_11603,N_10520,N_10916);
and U11604 (N_11604,N_10580,N_10058);
nor U11605 (N_11605,N_10163,N_10068);
xnor U11606 (N_11606,N_10678,N_10400);
xor U11607 (N_11607,N_10891,N_10391);
nor U11608 (N_11608,N_10997,N_10454);
or U11609 (N_11609,N_10131,N_10806);
and U11610 (N_11610,N_10725,N_10048);
nand U11611 (N_11611,N_10330,N_10213);
and U11612 (N_11612,N_10632,N_10756);
nand U11613 (N_11613,N_10994,N_10619);
xor U11614 (N_11614,N_10003,N_10152);
xor U11615 (N_11615,N_10375,N_10024);
and U11616 (N_11616,N_10488,N_10361);
and U11617 (N_11617,N_10846,N_10814);
or U11618 (N_11618,N_10450,N_10961);
or U11619 (N_11619,N_10013,N_10202);
and U11620 (N_11620,N_10952,N_10547);
nor U11621 (N_11621,N_10269,N_10682);
xnor U11622 (N_11622,N_10809,N_10080);
or U11623 (N_11623,N_10571,N_10184);
or U11624 (N_11624,N_10552,N_10231);
nor U11625 (N_11625,N_10922,N_10383);
nor U11626 (N_11626,N_10800,N_10139);
or U11627 (N_11627,N_10452,N_10357);
nor U11628 (N_11628,N_10699,N_10948);
xnor U11629 (N_11629,N_10854,N_10520);
nor U11630 (N_11630,N_10210,N_10793);
and U11631 (N_11631,N_10516,N_10270);
nand U11632 (N_11632,N_10937,N_10513);
xnor U11633 (N_11633,N_10046,N_10311);
or U11634 (N_11634,N_10477,N_10499);
xnor U11635 (N_11635,N_10750,N_10815);
xnor U11636 (N_11636,N_10428,N_10562);
and U11637 (N_11637,N_10981,N_10800);
and U11638 (N_11638,N_10392,N_10062);
nand U11639 (N_11639,N_10889,N_10760);
nand U11640 (N_11640,N_10497,N_10570);
nor U11641 (N_11641,N_10072,N_10222);
or U11642 (N_11642,N_10896,N_10088);
or U11643 (N_11643,N_10610,N_10996);
and U11644 (N_11644,N_10653,N_10862);
xnor U11645 (N_11645,N_10530,N_10585);
nand U11646 (N_11646,N_10872,N_10671);
nand U11647 (N_11647,N_10086,N_10515);
nand U11648 (N_11648,N_10447,N_10609);
nor U11649 (N_11649,N_10562,N_10059);
or U11650 (N_11650,N_10863,N_10588);
or U11651 (N_11651,N_10322,N_10125);
nand U11652 (N_11652,N_10458,N_10543);
nor U11653 (N_11653,N_10776,N_10100);
xnor U11654 (N_11654,N_10364,N_10526);
or U11655 (N_11655,N_10233,N_10168);
nor U11656 (N_11656,N_10221,N_10043);
nor U11657 (N_11657,N_10317,N_10361);
xor U11658 (N_11658,N_10973,N_10419);
nor U11659 (N_11659,N_10818,N_10440);
and U11660 (N_11660,N_10776,N_10701);
nand U11661 (N_11661,N_10483,N_10648);
xnor U11662 (N_11662,N_10703,N_10875);
and U11663 (N_11663,N_10920,N_10599);
or U11664 (N_11664,N_10019,N_10359);
and U11665 (N_11665,N_10031,N_10116);
or U11666 (N_11666,N_10672,N_10577);
nor U11667 (N_11667,N_10966,N_10670);
nor U11668 (N_11668,N_10726,N_10540);
nand U11669 (N_11669,N_10405,N_10287);
xnor U11670 (N_11670,N_10747,N_10070);
nor U11671 (N_11671,N_10749,N_10351);
nor U11672 (N_11672,N_10314,N_10834);
nand U11673 (N_11673,N_10173,N_10865);
or U11674 (N_11674,N_10854,N_10458);
and U11675 (N_11675,N_10776,N_10331);
or U11676 (N_11676,N_10870,N_10761);
nor U11677 (N_11677,N_10415,N_10532);
and U11678 (N_11678,N_10794,N_10991);
nor U11679 (N_11679,N_10458,N_10672);
nand U11680 (N_11680,N_10301,N_10098);
xnor U11681 (N_11681,N_10123,N_10964);
nor U11682 (N_11682,N_10814,N_10848);
nand U11683 (N_11683,N_10196,N_10687);
and U11684 (N_11684,N_10890,N_10572);
nor U11685 (N_11685,N_10761,N_10078);
or U11686 (N_11686,N_10506,N_10113);
xnor U11687 (N_11687,N_10267,N_10503);
nand U11688 (N_11688,N_10758,N_10731);
and U11689 (N_11689,N_10716,N_10927);
and U11690 (N_11690,N_10583,N_10841);
or U11691 (N_11691,N_10001,N_10046);
xor U11692 (N_11692,N_10675,N_10514);
nand U11693 (N_11693,N_10611,N_10044);
xor U11694 (N_11694,N_10171,N_10106);
xor U11695 (N_11695,N_10038,N_10619);
and U11696 (N_11696,N_10708,N_10854);
nand U11697 (N_11697,N_10126,N_10120);
or U11698 (N_11698,N_10612,N_10873);
and U11699 (N_11699,N_10433,N_10170);
or U11700 (N_11700,N_10601,N_10261);
nand U11701 (N_11701,N_10157,N_10057);
nor U11702 (N_11702,N_10069,N_10225);
or U11703 (N_11703,N_10385,N_10689);
nand U11704 (N_11704,N_10225,N_10915);
xnor U11705 (N_11705,N_10757,N_10281);
and U11706 (N_11706,N_10268,N_10325);
and U11707 (N_11707,N_10287,N_10738);
nor U11708 (N_11708,N_10988,N_10028);
xor U11709 (N_11709,N_10061,N_10430);
xnor U11710 (N_11710,N_10953,N_10923);
or U11711 (N_11711,N_10508,N_10332);
or U11712 (N_11712,N_10713,N_10512);
xor U11713 (N_11713,N_10694,N_10393);
nor U11714 (N_11714,N_10037,N_10327);
and U11715 (N_11715,N_10668,N_10796);
nor U11716 (N_11716,N_10085,N_10454);
nor U11717 (N_11717,N_10033,N_10354);
nor U11718 (N_11718,N_10322,N_10310);
xnor U11719 (N_11719,N_10328,N_10528);
and U11720 (N_11720,N_10948,N_10161);
or U11721 (N_11721,N_10294,N_10327);
or U11722 (N_11722,N_10626,N_10629);
nand U11723 (N_11723,N_10106,N_10018);
and U11724 (N_11724,N_10400,N_10560);
nand U11725 (N_11725,N_10763,N_10153);
nand U11726 (N_11726,N_10647,N_10675);
and U11727 (N_11727,N_10372,N_10321);
and U11728 (N_11728,N_10994,N_10711);
nor U11729 (N_11729,N_10706,N_10950);
or U11730 (N_11730,N_10090,N_10526);
nor U11731 (N_11731,N_10927,N_10045);
xnor U11732 (N_11732,N_10143,N_10235);
xnor U11733 (N_11733,N_10925,N_10949);
nand U11734 (N_11734,N_10102,N_10453);
or U11735 (N_11735,N_10227,N_10522);
nand U11736 (N_11736,N_10182,N_10891);
xnor U11737 (N_11737,N_10876,N_10150);
and U11738 (N_11738,N_10853,N_10864);
or U11739 (N_11739,N_10760,N_10341);
or U11740 (N_11740,N_10981,N_10815);
nor U11741 (N_11741,N_10443,N_10658);
nor U11742 (N_11742,N_10292,N_10513);
and U11743 (N_11743,N_10944,N_10585);
nand U11744 (N_11744,N_10780,N_10394);
and U11745 (N_11745,N_10038,N_10722);
or U11746 (N_11746,N_10152,N_10891);
nand U11747 (N_11747,N_10492,N_10639);
nand U11748 (N_11748,N_10264,N_10046);
and U11749 (N_11749,N_10243,N_10349);
or U11750 (N_11750,N_10421,N_10563);
nand U11751 (N_11751,N_10468,N_10861);
nor U11752 (N_11752,N_10584,N_10832);
nor U11753 (N_11753,N_10687,N_10514);
and U11754 (N_11754,N_10767,N_10526);
and U11755 (N_11755,N_10196,N_10081);
nor U11756 (N_11756,N_10629,N_10812);
or U11757 (N_11757,N_10576,N_10888);
or U11758 (N_11758,N_10501,N_10150);
and U11759 (N_11759,N_10832,N_10419);
xor U11760 (N_11760,N_10512,N_10435);
or U11761 (N_11761,N_10422,N_10228);
or U11762 (N_11762,N_10740,N_10280);
or U11763 (N_11763,N_10042,N_10670);
nor U11764 (N_11764,N_10482,N_10466);
or U11765 (N_11765,N_10913,N_10108);
and U11766 (N_11766,N_10829,N_10865);
or U11767 (N_11767,N_10656,N_10049);
nand U11768 (N_11768,N_10807,N_10767);
xnor U11769 (N_11769,N_10900,N_10248);
or U11770 (N_11770,N_10659,N_10886);
xor U11771 (N_11771,N_10864,N_10376);
nor U11772 (N_11772,N_10834,N_10821);
and U11773 (N_11773,N_10349,N_10021);
and U11774 (N_11774,N_10974,N_10360);
or U11775 (N_11775,N_10547,N_10482);
nand U11776 (N_11776,N_10216,N_10280);
nor U11777 (N_11777,N_10790,N_10150);
nand U11778 (N_11778,N_10001,N_10712);
nand U11779 (N_11779,N_10337,N_10710);
xnor U11780 (N_11780,N_10887,N_10467);
and U11781 (N_11781,N_10641,N_10394);
nor U11782 (N_11782,N_10543,N_10349);
xnor U11783 (N_11783,N_10498,N_10238);
xor U11784 (N_11784,N_10739,N_10258);
or U11785 (N_11785,N_10092,N_10693);
nor U11786 (N_11786,N_10803,N_10435);
nor U11787 (N_11787,N_10625,N_10507);
nand U11788 (N_11788,N_10671,N_10080);
nor U11789 (N_11789,N_10937,N_10742);
or U11790 (N_11790,N_10474,N_10892);
nand U11791 (N_11791,N_10665,N_10821);
nor U11792 (N_11792,N_10433,N_10871);
nor U11793 (N_11793,N_10917,N_10288);
or U11794 (N_11794,N_10454,N_10876);
nor U11795 (N_11795,N_10233,N_10420);
nand U11796 (N_11796,N_10697,N_10241);
nor U11797 (N_11797,N_10158,N_10394);
nor U11798 (N_11798,N_10168,N_10663);
and U11799 (N_11799,N_10428,N_10211);
and U11800 (N_11800,N_10911,N_10711);
or U11801 (N_11801,N_10514,N_10005);
nand U11802 (N_11802,N_10097,N_10989);
and U11803 (N_11803,N_10923,N_10779);
xnor U11804 (N_11804,N_10301,N_10568);
nor U11805 (N_11805,N_10818,N_10746);
nor U11806 (N_11806,N_10862,N_10683);
or U11807 (N_11807,N_10150,N_10302);
or U11808 (N_11808,N_10488,N_10567);
nor U11809 (N_11809,N_10965,N_10144);
nand U11810 (N_11810,N_10696,N_10170);
and U11811 (N_11811,N_10853,N_10403);
and U11812 (N_11812,N_10335,N_10473);
nor U11813 (N_11813,N_10425,N_10266);
and U11814 (N_11814,N_10760,N_10363);
nand U11815 (N_11815,N_10468,N_10788);
or U11816 (N_11816,N_10911,N_10103);
or U11817 (N_11817,N_10494,N_10090);
nand U11818 (N_11818,N_10413,N_10429);
nand U11819 (N_11819,N_10587,N_10817);
and U11820 (N_11820,N_10207,N_10775);
nand U11821 (N_11821,N_10052,N_10386);
nand U11822 (N_11822,N_10936,N_10226);
and U11823 (N_11823,N_10115,N_10241);
xnor U11824 (N_11824,N_10017,N_10785);
and U11825 (N_11825,N_10633,N_10060);
and U11826 (N_11826,N_10847,N_10269);
nor U11827 (N_11827,N_10038,N_10860);
and U11828 (N_11828,N_10186,N_10336);
nand U11829 (N_11829,N_10909,N_10148);
xnor U11830 (N_11830,N_10676,N_10135);
or U11831 (N_11831,N_10183,N_10692);
or U11832 (N_11832,N_10763,N_10308);
nand U11833 (N_11833,N_10045,N_10799);
and U11834 (N_11834,N_10124,N_10451);
and U11835 (N_11835,N_10481,N_10426);
nor U11836 (N_11836,N_10532,N_10466);
xnor U11837 (N_11837,N_10943,N_10721);
xnor U11838 (N_11838,N_10632,N_10700);
and U11839 (N_11839,N_10630,N_10354);
or U11840 (N_11840,N_10210,N_10825);
and U11841 (N_11841,N_10159,N_10172);
nor U11842 (N_11842,N_10823,N_10425);
and U11843 (N_11843,N_10748,N_10894);
xor U11844 (N_11844,N_10535,N_10262);
nor U11845 (N_11845,N_10946,N_10162);
nor U11846 (N_11846,N_10208,N_10115);
and U11847 (N_11847,N_10167,N_10432);
xnor U11848 (N_11848,N_10957,N_10035);
nand U11849 (N_11849,N_10738,N_10001);
nor U11850 (N_11850,N_10474,N_10861);
nand U11851 (N_11851,N_10955,N_10441);
nor U11852 (N_11852,N_10331,N_10916);
nand U11853 (N_11853,N_10250,N_10171);
xor U11854 (N_11854,N_10230,N_10843);
or U11855 (N_11855,N_10088,N_10401);
nand U11856 (N_11856,N_10975,N_10618);
or U11857 (N_11857,N_10942,N_10046);
nand U11858 (N_11858,N_10129,N_10431);
xnor U11859 (N_11859,N_10092,N_10070);
nand U11860 (N_11860,N_10959,N_10073);
or U11861 (N_11861,N_10433,N_10809);
nor U11862 (N_11862,N_10927,N_10149);
nor U11863 (N_11863,N_10890,N_10387);
and U11864 (N_11864,N_10608,N_10321);
nand U11865 (N_11865,N_10852,N_10468);
and U11866 (N_11866,N_10327,N_10383);
xor U11867 (N_11867,N_10289,N_10374);
nand U11868 (N_11868,N_10002,N_10216);
and U11869 (N_11869,N_10691,N_10817);
or U11870 (N_11870,N_10693,N_10990);
and U11871 (N_11871,N_10730,N_10130);
and U11872 (N_11872,N_10322,N_10446);
nand U11873 (N_11873,N_10641,N_10651);
and U11874 (N_11874,N_10370,N_10006);
nand U11875 (N_11875,N_10784,N_10909);
or U11876 (N_11876,N_10661,N_10922);
nor U11877 (N_11877,N_10125,N_10060);
or U11878 (N_11878,N_10198,N_10704);
and U11879 (N_11879,N_10602,N_10985);
nand U11880 (N_11880,N_10418,N_10416);
and U11881 (N_11881,N_10215,N_10995);
or U11882 (N_11882,N_10020,N_10189);
xor U11883 (N_11883,N_10223,N_10503);
nand U11884 (N_11884,N_10728,N_10553);
nor U11885 (N_11885,N_10544,N_10542);
and U11886 (N_11886,N_10201,N_10203);
xor U11887 (N_11887,N_10571,N_10421);
and U11888 (N_11888,N_10320,N_10661);
xor U11889 (N_11889,N_10460,N_10506);
nand U11890 (N_11890,N_10232,N_10170);
and U11891 (N_11891,N_10510,N_10092);
xnor U11892 (N_11892,N_10922,N_10311);
or U11893 (N_11893,N_10668,N_10604);
or U11894 (N_11894,N_10961,N_10588);
xor U11895 (N_11895,N_10306,N_10378);
nor U11896 (N_11896,N_10301,N_10786);
nor U11897 (N_11897,N_10741,N_10301);
nand U11898 (N_11898,N_10072,N_10421);
and U11899 (N_11899,N_10555,N_10445);
nor U11900 (N_11900,N_10145,N_10771);
xor U11901 (N_11901,N_10793,N_10327);
and U11902 (N_11902,N_10398,N_10714);
nand U11903 (N_11903,N_10057,N_10564);
and U11904 (N_11904,N_10141,N_10382);
and U11905 (N_11905,N_10441,N_10300);
and U11906 (N_11906,N_10037,N_10623);
xnor U11907 (N_11907,N_10965,N_10121);
and U11908 (N_11908,N_10839,N_10666);
nor U11909 (N_11909,N_10284,N_10130);
xor U11910 (N_11910,N_10463,N_10401);
nand U11911 (N_11911,N_10710,N_10846);
xnor U11912 (N_11912,N_10375,N_10521);
nor U11913 (N_11913,N_10914,N_10209);
xnor U11914 (N_11914,N_10371,N_10118);
nand U11915 (N_11915,N_10279,N_10227);
nand U11916 (N_11916,N_10323,N_10948);
and U11917 (N_11917,N_10301,N_10882);
or U11918 (N_11918,N_10716,N_10614);
nand U11919 (N_11919,N_10982,N_10573);
or U11920 (N_11920,N_10557,N_10738);
and U11921 (N_11921,N_10932,N_10958);
or U11922 (N_11922,N_10581,N_10366);
nand U11923 (N_11923,N_10765,N_10705);
and U11924 (N_11924,N_10781,N_10836);
or U11925 (N_11925,N_10004,N_10756);
or U11926 (N_11926,N_10259,N_10603);
or U11927 (N_11927,N_10369,N_10683);
nand U11928 (N_11928,N_10880,N_10062);
xnor U11929 (N_11929,N_10089,N_10108);
and U11930 (N_11930,N_10316,N_10142);
nand U11931 (N_11931,N_10559,N_10269);
nor U11932 (N_11932,N_10102,N_10756);
or U11933 (N_11933,N_10369,N_10456);
or U11934 (N_11934,N_10757,N_10128);
nor U11935 (N_11935,N_10220,N_10178);
xnor U11936 (N_11936,N_10975,N_10525);
or U11937 (N_11937,N_10909,N_10618);
and U11938 (N_11938,N_10316,N_10322);
and U11939 (N_11939,N_10414,N_10285);
or U11940 (N_11940,N_10639,N_10704);
and U11941 (N_11941,N_10851,N_10598);
and U11942 (N_11942,N_10063,N_10473);
or U11943 (N_11943,N_10639,N_10892);
nor U11944 (N_11944,N_10681,N_10703);
or U11945 (N_11945,N_10992,N_10280);
and U11946 (N_11946,N_10034,N_10120);
and U11947 (N_11947,N_10187,N_10031);
xnor U11948 (N_11948,N_10616,N_10058);
xnor U11949 (N_11949,N_10821,N_10423);
xor U11950 (N_11950,N_10474,N_10002);
nand U11951 (N_11951,N_10435,N_10417);
and U11952 (N_11952,N_10213,N_10542);
nor U11953 (N_11953,N_10591,N_10024);
and U11954 (N_11954,N_10184,N_10597);
nor U11955 (N_11955,N_10425,N_10698);
nor U11956 (N_11956,N_10510,N_10542);
nand U11957 (N_11957,N_10906,N_10706);
and U11958 (N_11958,N_10290,N_10953);
xor U11959 (N_11959,N_10083,N_10443);
or U11960 (N_11960,N_10363,N_10364);
nor U11961 (N_11961,N_10277,N_10222);
or U11962 (N_11962,N_10758,N_10374);
and U11963 (N_11963,N_10569,N_10160);
xnor U11964 (N_11964,N_10652,N_10382);
or U11965 (N_11965,N_10999,N_10976);
xor U11966 (N_11966,N_10579,N_10406);
and U11967 (N_11967,N_10701,N_10629);
xnor U11968 (N_11968,N_10455,N_10057);
nor U11969 (N_11969,N_10614,N_10037);
nand U11970 (N_11970,N_10062,N_10972);
nand U11971 (N_11971,N_10752,N_10609);
or U11972 (N_11972,N_10826,N_10469);
nand U11973 (N_11973,N_10646,N_10341);
nand U11974 (N_11974,N_10698,N_10095);
or U11975 (N_11975,N_10426,N_10950);
or U11976 (N_11976,N_10919,N_10403);
and U11977 (N_11977,N_10257,N_10782);
and U11978 (N_11978,N_10876,N_10048);
nor U11979 (N_11979,N_10841,N_10833);
xor U11980 (N_11980,N_10642,N_10725);
nor U11981 (N_11981,N_10067,N_10483);
or U11982 (N_11982,N_10199,N_10178);
nand U11983 (N_11983,N_10020,N_10530);
or U11984 (N_11984,N_10541,N_10079);
and U11985 (N_11985,N_10712,N_10963);
and U11986 (N_11986,N_10956,N_10991);
or U11987 (N_11987,N_10905,N_10907);
nor U11988 (N_11988,N_10582,N_10014);
nand U11989 (N_11989,N_10749,N_10793);
or U11990 (N_11990,N_10655,N_10689);
and U11991 (N_11991,N_10885,N_10524);
or U11992 (N_11992,N_10714,N_10829);
and U11993 (N_11993,N_10959,N_10489);
and U11994 (N_11994,N_10888,N_10977);
xnor U11995 (N_11995,N_10710,N_10432);
nor U11996 (N_11996,N_10097,N_10750);
and U11997 (N_11997,N_10577,N_10332);
nand U11998 (N_11998,N_10672,N_10291);
and U11999 (N_11999,N_10474,N_10882);
xnor U12000 (N_12000,N_11038,N_11520);
nand U12001 (N_12001,N_11161,N_11508);
nor U12002 (N_12002,N_11361,N_11286);
or U12003 (N_12003,N_11192,N_11719);
nor U12004 (N_12004,N_11316,N_11403);
or U12005 (N_12005,N_11321,N_11611);
or U12006 (N_12006,N_11069,N_11681);
and U12007 (N_12007,N_11685,N_11747);
and U12008 (N_12008,N_11770,N_11895);
and U12009 (N_12009,N_11813,N_11310);
nor U12010 (N_12010,N_11757,N_11975);
nand U12011 (N_12011,N_11124,N_11208);
and U12012 (N_12012,N_11226,N_11665);
or U12013 (N_12013,N_11198,N_11515);
xnor U12014 (N_12014,N_11004,N_11015);
xor U12015 (N_12015,N_11847,N_11604);
or U12016 (N_12016,N_11011,N_11993);
nand U12017 (N_12017,N_11119,N_11866);
and U12018 (N_12018,N_11439,N_11413);
nand U12019 (N_12019,N_11697,N_11320);
nor U12020 (N_12020,N_11898,N_11746);
or U12021 (N_12021,N_11818,N_11451);
xnor U12022 (N_12022,N_11894,N_11752);
and U12023 (N_12023,N_11315,N_11715);
and U12024 (N_12024,N_11741,N_11743);
or U12025 (N_12025,N_11978,N_11142);
and U12026 (N_12026,N_11998,N_11060);
nor U12027 (N_12027,N_11381,N_11420);
xor U12028 (N_12028,N_11750,N_11678);
and U12029 (N_12029,N_11332,N_11127);
or U12030 (N_12030,N_11964,N_11560);
nand U12031 (N_12031,N_11425,N_11905);
and U12032 (N_12032,N_11382,N_11174);
nor U12033 (N_12033,N_11555,N_11917);
nor U12034 (N_12034,N_11667,N_11612);
nor U12035 (N_12035,N_11630,N_11085);
and U12036 (N_12036,N_11787,N_11772);
nor U12037 (N_12037,N_11704,N_11564);
or U12038 (N_12038,N_11372,N_11729);
xnor U12039 (N_12039,N_11029,N_11991);
xnor U12040 (N_12040,N_11789,N_11846);
or U12041 (N_12041,N_11351,N_11014);
nand U12042 (N_12042,N_11405,N_11983);
or U12043 (N_12043,N_11243,N_11220);
nor U12044 (N_12044,N_11553,N_11362);
or U12045 (N_12045,N_11797,N_11404);
or U12046 (N_12046,N_11341,N_11094);
nand U12047 (N_12047,N_11526,N_11945);
nand U12048 (N_12048,N_11650,N_11102);
nand U12049 (N_12049,N_11597,N_11954);
and U12050 (N_12050,N_11644,N_11334);
or U12051 (N_12051,N_11767,N_11911);
nand U12052 (N_12052,N_11521,N_11875);
or U12053 (N_12053,N_11242,N_11231);
or U12054 (N_12054,N_11516,N_11354);
xor U12055 (N_12055,N_11497,N_11267);
xnor U12056 (N_12056,N_11578,N_11478);
xnor U12057 (N_12057,N_11620,N_11036);
or U12058 (N_12058,N_11798,N_11180);
and U12059 (N_12059,N_11135,N_11854);
nor U12060 (N_12060,N_11962,N_11549);
nor U12061 (N_12061,N_11328,N_11087);
nor U12062 (N_12062,N_11322,N_11380);
nand U12063 (N_12063,N_11754,N_11724);
nand U12064 (N_12064,N_11392,N_11622);
and U12065 (N_12065,N_11988,N_11475);
nand U12066 (N_12066,N_11112,N_11456);
nor U12067 (N_12067,N_11594,N_11663);
xnor U12068 (N_12068,N_11244,N_11901);
nor U12069 (N_12069,N_11929,N_11337);
xor U12070 (N_12070,N_11708,N_11369);
or U12071 (N_12071,N_11502,N_11995);
xor U12072 (N_12072,N_11629,N_11646);
nor U12073 (N_12073,N_11093,N_11671);
nor U12074 (N_12074,N_11336,N_11982);
or U12075 (N_12075,N_11677,N_11571);
xor U12076 (N_12076,N_11169,N_11976);
xor U12077 (N_12077,N_11997,N_11842);
nand U12078 (N_12078,N_11951,N_11047);
nand U12079 (N_12079,N_11943,N_11915);
xor U12080 (N_12080,N_11907,N_11299);
or U12081 (N_12081,N_11494,N_11805);
nor U12082 (N_12082,N_11430,N_11376);
nor U12083 (N_12083,N_11079,N_11283);
or U12084 (N_12084,N_11407,N_11638);
nand U12085 (N_12085,N_11931,N_11680);
xor U12086 (N_12086,N_11327,N_11305);
nor U12087 (N_12087,N_11543,N_11324);
nand U12088 (N_12088,N_11281,N_11709);
and U12089 (N_12089,N_11730,N_11696);
or U12090 (N_12090,N_11936,N_11554);
or U12091 (N_12091,N_11821,N_11768);
nand U12092 (N_12092,N_11209,N_11500);
and U12093 (N_12093,N_11904,N_11733);
nor U12094 (N_12094,N_11482,N_11261);
nor U12095 (N_12095,N_11265,N_11559);
nor U12096 (N_12096,N_11517,N_11486);
nand U12097 (N_12097,N_11593,N_11417);
or U12098 (N_12098,N_11230,N_11609);
and U12099 (N_12099,N_11375,N_11177);
and U12100 (N_12100,N_11817,N_11984);
nor U12101 (N_12101,N_11247,N_11736);
nand U12102 (N_12102,N_11223,N_11173);
or U12103 (N_12103,N_11147,N_11022);
nor U12104 (N_12104,N_11833,N_11355);
nand U12105 (N_12105,N_11883,N_11097);
or U12106 (N_12106,N_11170,N_11419);
and U12107 (N_12107,N_11062,N_11289);
or U12108 (N_12108,N_11167,N_11181);
nor U12109 (N_12109,N_11437,N_11987);
nor U12110 (N_12110,N_11676,N_11568);
nand U12111 (N_12111,N_11657,N_11352);
nor U12112 (N_12112,N_11675,N_11734);
nor U12113 (N_12113,N_11184,N_11445);
and U12114 (N_12114,N_11346,N_11207);
nor U12115 (N_12115,N_11851,N_11980);
and U12116 (N_12116,N_11706,N_11623);
nand U12117 (N_12117,N_11021,N_11303);
or U12118 (N_12118,N_11211,N_11460);
or U12119 (N_12119,N_11870,N_11891);
nor U12120 (N_12120,N_11151,N_11467);
nand U12121 (N_12121,N_11879,N_11115);
or U12122 (N_12122,N_11602,N_11892);
nand U12123 (N_12123,N_11458,N_11105);
and U12124 (N_12124,N_11826,N_11273);
nor U12125 (N_12125,N_11459,N_11044);
nand U12126 (N_12126,N_11534,N_11791);
and U12127 (N_12127,N_11807,N_11994);
and U12128 (N_12128,N_11596,N_11471);
or U12129 (N_12129,N_11288,N_11738);
xor U12130 (N_12130,N_11318,N_11873);
xor U12131 (N_12131,N_11258,N_11009);
or U12132 (N_12132,N_11503,N_11587);
xor U12133 (N_12133,N_11284,N_11837);
or U12134 (N_12134,N_11639,N_11057);
xor U12135 (N_12135,N_11902,N_11777);
nand U12136 (N_12136,N_11579,N_11956);
nand U12137 (N_12137,N_11013,N_11916);
xnor U12138 (N_12138,N_11974,N_11280);
or U12139 (N_12139,N_11156,N_11477);
xnor U12140 (N_12140,N_11003,N_11969);
or U12141 (N_12141,N_11695,N_11563);
xor U12142 (N_12142,N_11507,N_11979);
nor U12143 (N_12143,N_11130,N_11148);
nor U12144 (N_12144,N_11914,N_11290);
and U12145 (N_12145,N_11399,N_11766);
and U12146 (N_12146,N_11006,N_11199);
xor U12147 (N_12147,N_11925,N_11648);
xnor U12148 (N_12148,N_11292,N_11692);
nor U12149 (N_12149,N_11647,N_11653);
or U12150 (N_12150,N_11074,N_11531);
nand U12151 (N_12151,N_11282,N_11927);
or U12152 (N_12152,N_11092,N_11589);
xor U12153 (N_12153,N_11252,N_11890);
nand U12154 (N_12154,N_11213,N_11628);
or U12155 (N_12155,N_11479,N_11463);
or U12156 (N_12156,N_11095,N_11919);
nor U12157 (N_12157,N_11137,N_11547);
or U12158 (N_12158,N_11809,N_11504);
xor U12159 (N_12159,N_11260,N_11251);
nand U12160 (N_12160,N_11640,N_11388);
nand U12161 (N_12161,N_11353,N_11365);
xor U12162 (N_12162,N_11838,N_11725);
and U12163 (N_12163,N_11576,N_11253);
nor U12164 (N_12164,N_11977,N_11990);
and U12165 (N_12165,N_11468,N_11270);
or U12166 (N_12166,N_11435,N_11558);
and U12167 (N_12167,N_11073,N_11162);
and U12168 (N_12168,N_11737,N_11548);
or U12169 (N_12169,N_11820,N_11026);
xnor U12170 (N_12170,N_11091,N_11501);
xor U12171 (N_12171,N_11386,N_11368);
nor U12172 (N_12172,N_11783,N_11586);
xor U12173 (N_12173,N_11072,N_11157);
nand U12174 (N_12174,N_11635,N_11924);
nor U12175 (N_12175,N_11212,N_11016);
or U12176 (N_12176,N_11721,N_11236);
nand U12177 (N_12177,N_11309,N_11858);
nor U12178 (N_12178,N_11195,N_11947);
nor U12179 (N_12179,N_11032,N_11776);
nand U12180 (N_12180,N_11132,N_11512);
nand U12181 (N_12181,N_11686,N_11900);
nor U12182 (N_12182,N_11317,N_11514);
xor U12183 (N_12183,N_11771,N_11371);
xnor U12184 (N_12184,N_11155,N_11331);
nor U12185 (N_12185,N_11567,N_11800);
or U12186 (N_12186,N_11410,N_11271);
xor U12187 (N_12187,N_11849,N_11224);
nand U12188 (N_12188,N_11160,N_11228);
or U12189 (N_12189,N_11020,N_11918);
nand U12190 (N_12190,N_11786,N_11227);
xor U12191 (N_12191,N_11631,N_11498);
nor U12192 (N_12192,N_11489,N_11138);
nand U12193 (N_12193,N_11436,N_11163);
nand U12194 (N_12194,N_11496,N_11774);
nor U12195 (N_12195,N_11525,N_11189);
or U12196 (N_12196,N_11523,N_11679);
and U12197 (N_12197,N_11366,N_11557);
xor U12198 (N_12198,N_11356,N_11625);
and U12199 (N_12199,N_11136,N_11054);
or U12200 (N_12200,N_11100,N_11176);
or U12201 (N_12201,N_11035,N_11856);
nand U12202 (N_12202,N_11325,N_11803);
nor U12203 (N_12203,N_11530,N_11225);
or U12204 (N_12204,N_11277,N_11484);
xnor U12205 (N_12205,N_11519,N_11864);
xor U12206 (N_12206,N_11763,N_11887);
or U12207 (N_12207,N_11125,N_11159);
or U12208 (N_12208,N_11705,N_11999);
nand U12209 (N_12209,N_11397,N_11179);
and U12210 (N_12210,N_11215,N_11524);
nor U12211 (N_12211,N_11045,N_11882);
and U12212 (N_12212,N_11688,N_11010);
or U12213 (N_12213,N_11835,N_11963);
xor U12214 (N_12214,N_11699,N_11206);
xor U12215 (N_12215,N_11400,N_11043);
xor U12216 (N_12216,N_11845,N_11164);
xnor U12217 (N_12217,N_11432,N_11232);
nor U12218 (N_12218,N_11664,N_11098);
and U12219 (N_12219,N_11808,N_11731);
or U12220 (N_12220,N_11753,N_11541);
or U12221 (N_12221,N_11745,N_11465);
nor U12222 (N_12222,N_11831,N_11030);
and U12223 (N_12223,N_11391,N_11390);
xnor U12224 (N_12224,N_11150,N_11840);
or U12225 (N_12225,N_11201,N_11298);
and U12226 (N_12226,N_11690,N_11421);
or U12227 (N_12227,N_11001,N_11930);
nor U12228 (N_12228,N_11339,N_11063);
nor U12229 (N_12229,N_11480,N_11867);
nor U12230 (N_12230,N_11606,N_11565);
and U12231 (N_12231,N_11165,N_11735);
xor U12232 (N_12232,N_11145,N_11689);
nor U12233 (N_12233,N_11701,N_11275);
xor U12234 (N_12234,N_11510,N_11575);
or U12235 (N_12235,N_11308,N_11881);
nand U12236 (N_12236,N_11605,N_11241);
nor U12237 (N_12237,N_11957,N_11264);
or U12238 (N_12238,N_11522,N_11384);
nand U12239 (N_12239,N_11312,N_11133);
or U12240 (N_12240,N_11333,N_11438);
xor U12241 (N_12241,N_11815,N_11556);
and U12242 (N_12242,N_11483,N_11473);
xor U12243 (N_12243,N_11075,N_11246);
nand U12244 (N_12244,N_11285,N_11728);
nor U12245 (N_12245,N_11238,N_11722);
nand U12246 (N_12246,N_11046,N_11450);
nor U12247 (N_12247,N_11960,N_11139);
and U12248 (N_12248,N_11389,N_11023);
nand U12249 (N_12249,N_11633,N_11114);
and U12250 (N_12250,N_11717,N_11442);
xor U12251 (N_12251,N_11117,N_11345);
nor U12252 (N_12252,N_11792,N_11017);
and U12253 (N_12253,N_11278,N_11053);
or U12254 (N_12254,N_11823,N_11446);
and U12255 (N_12255,N_11595,N_11779);
nor U12256 (N_12256,N_11204,N_11096);
and U12257 (N_12257,N_11058,N_11052);
xnor U12258 (N_12258,N_11235,N_11518);
nor U12259 (N_12259,N_11217,N_11064);
and U12260 (N_12260,N_11935,N_11412);
or U12261 (N_12261,N_11641,N_11319);
nand U12262 (N_12262,N_11584,N_11617);
xnor U12263 (N_12263,N_11490,N_11784);
or U12264 (N_12264,N_11153,N_11423);
nor U12265 (N_12265,N_11222,N_11799);
nor U12266 (N_12266,N_11440,N_11387);
and U12267 (N_12267,N_11788,N_11666);
xnor U12268 (N_12268,N_11810,N_11670);
or U12269 (N_12269,N_11330,N_11953);
or U12270 (N_12270,N_11700,N_11297);
or U12271 (N_12271,N_11028,N_11909);
or U12272 (N_12272,N_11920,N_11506);
nand U12273 (N_12273,N_11812,N_11528);
nor U12274 (N_12274,N_11535,N_11269);
or U12275 (N_12275,N_11966,N_11027);
and U12276 (N_12276,N_11128,N_11830);
or U12277 (N_12277,N_11476,N_11785);
nand U12278 (N_12278,N_11279,N_11066);
or U12279 (N_12279,N_11110,N_11056);
and U12280 (N_12280,N_11860,N_11744);
and U12281 (N_12281,N_11068,N_11373);
xor U12282 (N_12282,N_11893,N_11886);
xnor U12283 (N_12283,N_11726,N_11684);
nor U12284 (N_12284,N_11740,N_11577);
nand U12285 (N_12285,N_11711,N_11775);
or U12286 (N_12286,N_11411,N_11034);
or U12287 (N_12287,N_11104,N_11229);
nand U12288 (N_12288,N_11108,N_11844);
xnor U12289 (N_12289,N_11985,N_11580);
or U12290 (N_12290,N_11972,N_11424);
nand U12291 (N_12291,N_11196,N_11616);
xnor U12292 (N_12292,N_11374,N_11455);
and U12293 (N_12293,N_11592,N_11089);
and U12294 (N_12294,N_11470,N_11143);
or U12295 (N_12295,N_11566,N_11154);
nor U12296 (N_12296,N_11827,N_11078);
nor U12297 (N_12297,N_11989,N_11487);
nor U12298 (N_12298,N_11673,N_11829);
xor U12299 (N_12299,N_11296,N_11140);
xnor U12300 (N_12300,N_11658,N_11219);
nor U12301 (N_12301,N_11019,N_11338);
and U12302 (N_12302,N_11903,N_11872);
and U12303 (N_12303,N_11913,N_11344);
nand U12304 (N_12304,N_11632,N_11481);
nand U12305 (N_12305,N_11878,N_11544);
nor U12306 (N_12306,N_11287,N_11614);
nor U12307 (N_12307,N_11464,N_11537);
xnor U12308 (N_12308,N_11533,N_11065);
or U12309 (N_12309,N_11950,N_11107);
or U12310 (N_12310,N_11581,N_11570);
or U12311 (N_12311,N_11839,N_11342);
and U12312 (N_12312,N_11645,N_11652);
xnor U12313 (N_12313,N_11123,N_11937);
nand U12314 (N_12314,N_11216,N_11959);
nand U12315 (N_12315,N_11532,N_11536);
xnor U12316 (N_12316,N_11472,N_11551);
nor U12317 (N_12317,N_11949,N_11041);
nand U12318 (N_12318,N_11939,N_11912);
nor U12319 (N_12319,N_11152,N_11245);
xnor U12320 (N_12320,N_11769,N_11801);
nand U12321 (N_12321,N_11585,N_11274);
and U12322 (N_12322,N_11178,N_11134);
nand U12323 (N_12323,N_11185,N_11707);
nand U12324 (N_12324,N_11843,N_11340);
nand U12325 (N_12325,N_11718,N_11773);
xor U12326 (N_12326,N_11923,N_11910);
nand U12327 (N_12327,N_11254,N_11329);
xor U12328 (N_12328,N_11590,N_11461);
or U12329 (N_12329,N_11335,N_11509);
nand U12330 (N_12330,N_11656,N_11061);
nand U12331 (N_12331,N_11965,N_11434);
or U12332 (N_12332,N_11859,N_11781);
xnor U12333 (N_12333,N_11562,N_11116);
xor U12334 (N_12334,N_11627,N_11702);
or U12335 (N_12335,N_11710,N_11493);
nor U12336 (N_12336,N_11025,N_11214);
nand U12337 (N_12337,N_11203,N_11669);
and U12338 (N_12338,N_11414,N_11349);
nor U12339 (N_12339,N_11377,N_11841);
xor U12340 (N_12340,N_11166,N_11070);
or U12341 (N_12341,N_11000,N_11857);
xnor U12342 (N_12342,N_11651,N_11008);
xnor U12343 (N_12343,N_11126,N_11921);
nand U12344 (N_12344,N_11444,N_11357);
or U12345 (N_12345,N_11158,N_11952);
or U12346 (N_12346,N_11938,N_11396);
xnor U12347 (N_12347,N_11491,N_11661);
xnor U12348 (N_12348,N_11416,N_11233);
and U12349 (N_12349,N_11002,N_11762);
or U12350 (N_12350,N_11326,N_11683);
nor U12351 (N_12351,N_11121,N_11941);
and U12352 (N_12352,N_11462,N_11113);
nand U12353 (N_12353,N_11863,N_11379);
or U12354 (N_12354,N_11819,N_11869);
or U12355 (N_12355,N_11083,N_11759);
nor U12356 (N_12356,N_11539,N_11732);
nand U12357 (N_12357,N_11449,N_11861);
nor U12358 (N_12358,N_11573,N_11933);
xnor U12359 (N_12359,N_11469,N_11865);
or U12360 (N_12360,N_11037,N_11853);
and U12361 (N_12361,N_11761,N_11120);
nand U12362 (N_12362,N_11615,N_11816);
nand U12363 (N_12363,N_11794,N_11802);
or U12364 (N_12364,N_11218,N_11603);
or U12365 (N_12365,N_11790,N_11109);
or U12366 (N_12366,N_11545,N_11687);
xnor U12367 (N_12367,N_11234,N_11583);
or U12368 (N_12368,N_11239,N_11415);
nand U12369 (N_12369,N_11529,N_11655);
nor U12370 (N_12370,N_11885,N_11649);
xnor U12371 (N_12371,N_11401,N_11183);
and U12372 (N_12372,N_11601,N_11452);
or U12373 (N_12373,N_11848,N_11996);
nor U12374 (N_12374,N_11877,N_11634);
xnor U12375 (N_12375,N_11946,N_11048);
and U12376 (N_12376,N_11221,N_11888);
and U12377 (N_12377,N_11934,N_11050);
nand U12378 (N_12378,N_11765,N_11505);
nand U12379 (N_12379,N_11492,N_11538);
and U12380 (N_12380,N_11262,N_11406);
and U12381 (N_12381,N_11090,N_11301);
xor U12382 (N_12382,N_11742,N_11051);
and U12383 (N_12383,N_11621,N_11550);
nor U12384 (N_12384,N_11402,N_11370);
and U12385 (N_12385,N_11144,N_11383);
xnor U12386 (N_12386,N_11850,N_11122);
xor U12387 (N_12387,N_11986,N_11168);
nand U12388 (N_12388,N_11118,N_11276);
or U12389 (N_12389,N_11076,N_11080);
nor U12390 (N_12390,N_11572,N_11307);
and U12391 (N_12391,N_11205,N_11398);
xor U12392 (N_12392,N_11237,N_11928);
nor U12393 (N_12393,N_11499,N_11714);
xor U12394 (N_12394,N_11202,N_11457);
or U12395 (N_12395,N_11932,N_11598);
xor U12396 (N_12396,N_11485,N_11591);
nand U12397 (N_12397,N_11059,N_11200);
and U12398 (N_12398,N_11188,N_11782);
xnor U12399 (N_12399,N_11268,N_11992);
or U12400 (N_12400,N_11466,N_11613);
and U12401 (N_12401,N_11855,N_11693);
nand U12402 (N_12402,N_11306,N_11257);
xor U12403 (N_12403,N_11955,N_11662);
nand U12404 (N_12404,N_11973,N_11018);
nand U12405 (N_12405,N_11896,N_11131);
nor U12406 (N_12406,N_11088,N_11948);
xnor U12407 (N_12407,N_11637,N_11190);
xnor U12408 (N_12408,N_11323,N_11347);
and U12409 (N_12409,N_11447,N_11716);
nor U12410 (N_12410,N_11182,N_11042);
or U12411 (N_12411,N_11049,N_11084);
or U12412 (N_12412,N_11778,N_11582);
xor U12413 (N_12413,N_11795,N_11433);
nand U12414 (N_12414,N_11723,N_11314);
xnor U12415 (N_12415,N_11897,N_11958);
nor U12416 (N_12416,N_11540,N_11454);
xor U12417 (N_12417,N_11643,N_11824);
or U12418 (N_12418,N_11378,N_11364);
and U12419 (N_12419,N_11682,N_11348);
nor U12420 (N_12420,N_11626,N_11739);
xnor U12421 (N_12421,N_11618,N_11197);
nor U12422 (N_12422,N_11495,N_11129);
and U12423 (N_12423,N_11968,N_11852);
or U12424 (N_12424,N_11111,N_11619);
or U12425 (N_12425,N_11822,N_11141);
xnor U12426 (N_12426,N_11146,N_11249);
and U12427 (N_12427,N_11713,N_11263);
nor U12428 (N_12428,N_11961,N_11385);
and U12429 (N_12429,N_11636,N_11748);
nand U12430 (N_12430,N_11302,N_11828);
nor U12431 (N_12431,N_11876,N_11024);
xor U12432 (N_12432,N_11005,N_11428);
nor U12433 (N_12433,N_11106,N_11569);
xnor U12434 (N_12434,N_11031,N_11552);
nand U12435 (N_12435,N_11868,N_11443);
or U12436 (N_12436,N_11659,N_11294);
or U12437 (N_12437,N_11055,N_11874);
xnor U12438 (N_12438,N_11393,N_11033);
xor U12439 (N_12439,N_11250,N_11720);
and U12440 (N_12440,N_11077,N_11311);
nand U12441 (N_12441,N_11040,N_11814);
nor U12442 (N_12442,N_11453,N_11187);
and U12443 (N_12443,N_11880,N_11513);
and U12444 (N_12444,N_11363,N_11359);
nand U12445 (N_12445,N_11942,N_11608);
nand U12446 (N_12446,N_11511,N_11304);
and U12447 (N_12447,N_11674,N_11408);
or U12448 (N_12448,N_11967,N_11793);
nor U12449 (N_12449,N_11703,N_11099);
or U12450 (N_12450,N_11193,N_11691);
xor U12451 (N_12451,N_11429,N_11940);
nor U12452 (N_12452,N_11908,N_11186);
xor U12453 (N_12453,N_11588,N_11836);
xor U12454 (N_12454,N_11422,N_11474);
or U12455 (N_12455,N_11749,N_11394);
xnor U12456 (N_12456,N_11542,N_11210);
and U12457 (N_12457,N_11358,N_11295);
nor U12458 (N_12458,N_11796,N_11431);
or U12459 (N_12459,N_11610,N_11624);
xnor U12460 (N_12460,N_11780,N_11071);
or U12461 (N_12461,N_11367,N_11668);
and U12462 (N_12462,N_11395,N_11712);
xor U12463 (N_12463,N_11527,N_11427);
nand U12464 (N_12464,N_11081,N_11654);
or U12465 (N_12465,N_11804,N_11149);
and U12466 (N_12466,N_11760,N_11266);
and U12467 (N_12467,N_11832,N_11448);
nor U12468 (N_12468,N_11012,N_11922);
and U12469 (N_12469,N_11811,N_11350);
nor U12470 (N_12470,N_11694,N_11103);
nand U12471 (N_12471,N_11862,N_11889);
xor U12472 (N_12472,N_11067,N_11259);
xnor U12473 (N_12473,N_11291,N_11561);
nor U12474 (N_12474,N_11758,N_11599);
xor U12475 (N_12475,N_11884,N_11764);
or U12476 (N_12476,N_11418,N_11926);
nand U12477 (N_12477,N_11086,N_11194);
nand U12478 (N_12478,N_11672,N_11899);
or U12479 (N_12479,N_11727,N_11806);
nand U12480 (N_12480,N_11607,N_11409);
nor U12481 (N_12481,N_11971,N_11171);
nand U12482 (N_12482,N_11546,N_11756);
nor U12483 (N_12483,N_11240,N_11970);
and U12484 (N_12484,N_11248,N_11360);
xor U12485 (N_12485,N_11944,N_11698);
nor U12486 (N_12486,N_11313,N_11441);
nand U12487 (N_12487,N_11574,N_11834);
xnor U12488 (N_12488,N_11825,N_11255);
and U12489 (N_12489,N_11039,N_11191);
and U12490 (N_12490,N_11007,N_11082);
nor U12491 (N_12491,N_11642,N_11300);
xor U12492 (N_12492,N_11600,N_11755);
xor U12493 (N_12493,N_11293,N_11272);
and U12494 (N_12494,N_11172,N_11488);
or U12495 (N_12495,N_11426,N_11660);
nor U12496 (N_12496,N_11175,N_11906);
or U12497 (N_12497,N_11751,N_11101);
xor U12498 (N_12498,N_11256,N_11871);
nand U12499 (N_12499,N_11981,N_11343);
and U12500 (N_12500,N_11169,N_11368);
or U12501 (N_12501,N_11803,N_11789);
xor U12502 (N_12502,N_11833,N_11810);
nand U12503 (N_12503,N_11008,N_11014);
nand U12504 (N_12504,N_11545,N_11923);
nand U12505 (N_12505,N_11499,N_11526);
or U12506 (N_12506,N_11276,N_11935);
xor U12507 (N_12507,N_11296,N_11270);
and U12508 (N_12508,N_11671,N_11774);
nand U12509 (N_12509,N_11456,N_11559);
nand U12510 (N_12510,N_11053,N_11590);
xnor U12511 (N_12511,N_11805,N_11214);
nor U12512 (N_12512,N_11581,N_11165);
nand U12513 (N_12513,N_11262,N_11241);
nand U12514 (N_12514,N_11194,N_11139);
nand U12515 (N_12515,N_11141,N_11242);
xor U12516 (N_12516,N_11554,N_11439);
xnor U12517 (N_12517,N_11142,N_11048);
and U12518 (N_12518,N_11141,N_11385);
nand U12519 (N_12519,N_11662,N_11046);
and U12520 (N_12520,N_11650,N_11416);
nor U12521 (N_12521,N_11201,N_11079);
and U12522 (N_12522,N_11339,N_11197);
xor U12523 (N_12523,N_11019,N_11332);
xor U12524 (N_12524,N_11950,N_11898);
nor U12525 (N_12525,N_11015,N_11468);
xor U12526 (N_12526,N_11758,N_11896);
nor U12527 (N_12527,N_11635,N_11654);
and U12528 (N_12528,N_11384,N_11164);
xor U12529 (N_12529,N_11436,N_11845);
and U12530 (N_12530,N_11611,N_11923);
and U12531 (N_12531,N_11487,N_11095);
and U12532 (N_12532,N_11455,N_11092);
xor U12533 (N_12533,N_11771,N_11695);
nand U12534 (N_12534,N_11475,N_11413);
nand U12535 (N_12535,N_11061,N_11910);
nand U12536 (N_12536,N_11796,N_11292);
or U12537 (N_12537,N_11113,N_11836);
nor U12538 (N_12538,N_11119,N_11883);
or U12539 (N_12539,N_11581,N_11008);
nand U12540 (N_12540,N_11754,N_11350);
nor U12541 (N_12541,N_11985,N_11408);
and U12542 (N_12542,N_11064,N_11404);
nand U12543 (N_12543,N_11091,N_11862);
xor U12544 (N_12544,N_11224,N_11018);
xor U12545 (N_12545,N_11350,N_11671);
and U12546 (N_12546,N_11180,N_11944);
xor U12547 (N_12547,N_11654,N_11082);
or U12548 (N_12548,N_11838,N_11068);
xor U12549 (N_12549,N_11521,N_11283);
nor U12550 (N_12550,N_11883,N_11995);
or U12551 (N_12551,N_11039,N_11873);
xnor U12552 (N_12552,N_11613,N_11531);
nand U12553 (N_12553,N_11811,N_11612);
nor U12554 (N_12554,N_11896,N_11941);
nand U12555 (N_12555,N_11975,N_11166);
xor U12556 (N_12556,N_11858,N_11755);
nand U12557 (N_12557,N_11905,N_11379);
or U12558 (N_12558,N_11408,N_11730);
and U12559 (N_12559,N_11442,N_11451);
nand U12560 (N_12560,N_11296,N_11336);
nor U12561 (N_12561,N_11641,N_11111);
nor U12562 (N_12562,N_11085,N_11784);
xnor U12563 (N_12563,N_11352,N_11089);
or U12564 (N_12564,N_11492,N_11630);
and U12565 (N_12565,N_11880,N_11935);
xnor U12566 (N_12566,N_11721,N_11904);
and U12567 (N_12567,N_11461,N_11451);
or U12568 (N_12568,N_11698,N_11797);
nor U12569 (N_12569,N_11116,N_11006);
or U12570 (N_12570,N_11629,N_11336);
xnor U12571 (N_12571,N_11556,N_11114);
nor U12572 (N_12572,N_11169,N_11691);
nand U12573 (N_12573,N_11408,N_11379);
or U12574 (N_12574,N_11960,N_11538);
or U12575 (N_12575,N_11982,N_11965);
and U12576 (N_12576,N_11026,N_11489);
nor U12577 (N_12577,N_11757,N_11354);
and U12578 (N_12578,N_11776,N_11702);
nor U12579 (N_12579,N_11158,N_11736);
xnor U12580 (N_12580,N_11545,N_11119);
nand U12581 (N_12581,N_11031,N_11043);
xnor U12582 (N_12582,N_11725,N_11879);
nor U12583 (N_12583,N_11944,N_11524);
and U12584 (N_12584,N_11021,N_11603);
xor U12585 (N_12585,N_11660,N_11832);
and U12586 (N_12586,N_11077,N_11987);
nor U12587 (N_12587,N_11402,N_11211);
or U12588 (N_12588,N_11522,N_11717);
and U12589 (N_12589,N_11419,N_11651);
nand U12590 (N_12590,N_11407,N_11216);
nand U12591 (N_12591,N_11631,N_11059);
or U12592 (N_12592,N_11561,N_11461);
nand U12593 (N_12593,N_11369,N_11944);
xor U12594 (N_12594,N_11050,N_11295);
and U12595 (N_12595,N_11270,N_11548);
or U12596 (N_12596,N_11265,N_11242);
xnor U12597 (N_12597,N_11016,N_11096);
and U12598 (N_12598,N_11484,N_11121);
nand U12599 (N_12599,N_11307,N_11668);
nor U12600 (N_12600,N_11898,N_11859);
nand U12601 (N_12601,N_11850,N_11115);
nand U12602 (N_12602,N_11222,N_11247);
and U12603 (N_12603,N_11375,N_11426);
nor U12604 (N_12604,N_11538,N_11364);
xnor U12605 (N_12605,N_11949,N_11706);
or U12606 (N_12606,N_11103,N_11895);
and U12607 (N_12607,N_11598,N_11069);
nand U12608 (N_12608,N_11545,N_11507);
nor U12609 (N_12609,N_11291,N_11367);
nor U12610 (N_12610,N_11738,N_11951);
or U12611 (N_12611,N_11772,N_11746);
nand U12612 (N_12612,N_11538,N_11087);
and U12613 (N_12613,N_11285,N_11846);
and U12614 (N_12614,N_11216,N_11772);
or U12615 (N_12615,N_11985,N_11358);
nor U12616 (N_12616,N_11819,N_11613);
nand U12617 (N_12617,N_11052,N_11545);
xor U12618 (N_12618,N_11376,N_11561);
nand U12619 (N_12619,N_11373,N_11060);
xor U12620 (N_12620,N_11823,N_11417);
and U12621 (N_12621,N_11780,N_11287);
xnor U12622 (N_12622,N_11811,N_11607);
nor U12623 (N_12623,N_11296,N_11381);
or U12624 (N_12624,N_11131,N_11748);
and U12625 (N_12625,N_11336,N_11293);
and U12626 (N_12626,N_11653,N_11646);
nand U12627 (N_12627,N_11474,N_11384);
and U12628 (N_12628,N_11718,N_11291);
or U12629 (N_12629,N_11748,N_11379);
nand U12630 (N_12630,N_11508,N_11249);
nor U12631 (N_12631,N_11577,N_11136);
nand U12632 (N_12632,N_11551,N_11386);
nor U12633 (N_12633,N_11487,N_11656);
nor U12634 (N_12634,N_11703,N_11162);
and U12635 (N_12635,N_11046,N_11706);
or U12636 (N_12636,N_11184,N_11792);
xor U12637 (N_12637,N_11256,N_11096);
or U12638 (N_12638,N_11961,N_11045);
nor U12639 (N_12639,N_11765,N_11773);
nor U12640 (N_12640,N_11511,N_11582);
nand U12641 (N_12641,N_11100,N_11252);
nand U12642 (N_12642,N_11849,N_11903);
nor U12643 (N_12643,N_11053,N_11721);
xnor U12644 (N_12644,N_11012,N_11010);
and U12645 (N_12645,N_11323,N_11598);
or U12646 (N_12646,N_11728,N_11679);
and U12647 (N_12647,N_11466,N_11895);
and U12648 (N_12648,N_11255,N_11173);
nor U12649 (N_12649,N_11297,N_11868);
nand U12650 (N_12650,N_11710,N_11812);
nor U12651 (N_12651,N_11798,N_11842);
nand U12652 (N_12652,N_11976,N_11285);
nor U12653 (N_12653,N_11951,N_11018);
nand U12654 (N_12654,N_11604,N_11453);
nor U12655 (N_12655,N_11797,N_11901);
xnor U12656 (N_12656,N_11288,N_11609);
xor U12657 (N_12657,N_11911,N_11477);
or U12658 (N_12658,N_11620,N_11705);
nor U12659 (N_12659,N_11245,N_11071);
nor U12660 (N_12660,N_11479,N_11610);
nand U12661 (N_12661,N_11802,N_11095);
and U12662 (N_12662,N_11389,N_11517);
nor U12663 (N_12663,N_11816,N_11068);
nand U12664 (N_12664,N_11013,N_11831);
xor U12665 (N_12665,N_11680,N_11270);
xor U12666 (N_12666,N_11392,N_11932);
nor U12667 (N_12667,N_11668,N_11901);
and U12668 (N_12668,N_11032,N_11316);
and U12669 (N_12669,N_11115,N_11709);
xnor U12670 (N_12670,N_11453,N_11873);
xnor U12671 (N_12671,N_11895,N_11053);
and U12672 (N_12672,N_11864,N_11873);
or U12673 (N_12673,N_11718,N_11698);
or U12674 (N_12674,N_11955,N_11222);
or U12675 (N_12675,N_11616,N_11050);
nor U12676 (N_12676,N_11865,N_11056);
xnor U12677 (N_12677,N_11345,N_11686);
nand U12678 (N_12678,N_11900,N_11427);
nand U12679 (N_12679,N_11566,N_11852);
xor U12680 (N_12680,N_11926,N_11992);
nor U12681 (N_12681,N_11851,N_11253);
nand U12682 (N_12682,N_11675,N_11614);
nor U12683 (N_12683,N_11071,N_11911);
or U12684 (N_12684,N_11293,N_11138);
or U12685 (N_12685,N_11192,N_11893);
nand U12686 (N_12686,N_11419,N_11049);
nor U12687 (N_12687,N_11942,N_11459);
or U12688 (N_12688,N_11297,N_11663);
and U12689 (N_12689,N_11638,N_11064);
xor U12690 (N_12690,N_11546,N_11281);
or U12691 (N_12691,N_11546,N_11086);
nand U12692 (N_12692,N_11099,N_11850);
nand U12693 (N_12693,N_11947,N_11307);
nand U12694 (N_12694,N_11607,N_11420);
and U12695 (N_12695,N_11574,N_11774);
and U12696 (N_12696,N_11569,N_11286);
or U12697 (N_12697,N_11541,N_11564);
or U12698 (N_12698,N_11987,N_11579);
or U12699 (N_12699,N_11840,N_11404);
or U12700 (N_12700,N_11502,N_11443);
or U12701 (N_12701,N_11781,N_11416);
nand U12702 (N_12702,N_11614,N_11381);
or U12703 (N_12703,N_11368,N_11708);
and U12704 (N_12704,N_11793,N_11692);
or U12705 (N_12705,N_11761,N_11939);
xnor U12706 (N_12706,N_11814,N_11809);
xnor U12707 (N_12707,N_11749,N_11642);
and U12708 (N_12708,N_11752,N_11427);
or U12709 (N_12709,N_11582,N_11205);
nor U12710 (N_12710,N_11669,N_11174);
nand U12711 (N_12711,N_11469,N_11931);
or U12712 (N_12712,N_11850,N_11987);
or U12713 (N_12713,N_11592,N_11305);
xnor U12714 (N_12714,N_11573,N_11028);
nor U12715 (N_12715,N_11549,N_11006);
and U12716 (N_12716,N_11442,N_11137);
xor U12717 (N_12717,N_11036,N_11723);
or U12718 (N_12718,N_11870,N_11338);
nor U12719 (N_12719,N_11453,N_11769);
or U12720 (N_12720,N_11400,N_11060);
and U12721 (N_12721,N_11750,N_11349);
nor U12722 (N_12722,N_11213,N_11444);
or U12723 (N_12723,N_11936,N_11053);
or U12724 (N_12724,N_11571,N_11794);
nor U12725 (N_12725,N_11150,N_11950);
nand U12726 (N_12726,N_11449,N_11095);
xor U12727 (N_12727,N_11990,N_11010);
xor U12728 (N_12728,N_11683,N_11002);
nand U12729 (N_12729,N_11808,N_11550);
or U12730 (N_12730,N_11759,N_11777);
and U12731 (N_12731,N_11701,N_11388);
and U12732 (N_12732,N_11188,N_11529);
or U12733 (N_12733,N_11997,N_11204);
or U12734 (N_12734,N_11467,N_11358);
nor U12735 (N_12735,N_11367,N_11907);
nand U12736 (N_12736,N_11026,N_11097);
or U12737 (N_12737,N_11177,N_11889);
or U12738 (N_12738,N_11730,N_11697);
and U12739 (N_12739,N_11918,N_11341);
nor U12740 (N_12740,N_11086,N_11262);
or U12741 (N_12741,N_11007,N_11891);
and U12742 (N_12742,N_11373,N_11513);
nor U12743 (N_12743,N_11160,N_11171);
nand U12744 (N_12744,N_11210,N_11091);
nor U12745 (N_12745,N_11039,N_11464);
nor U12746 (N_12746,N_11359,N_11628);
xnor U12747 (N_12747,N_11103,N_11138);
nand U12748 (N_12748,N_11895,N_11286);
nand U12749 (N_12749,N_11678,N_11795);
nand U12750 (N_12750,N_11187,N_11749);
nor U12751 (N_12751,N_11609,N_11613);
nor U12752 (N_12752,N_11959,N_11155);
and U12753 (N_12753,N_11931,N_11446);
xor U12754 (N_12754,N_11801,N_11662);
nor U12755 (N_12755,N_11867,N_11508);
xor U12756 (N_12756,N_11337,N_11949);
nor U12757 (N_12757,N_11352,N_11362);
and U12758 (N_12758,N_11316,N_11876);
or U12759 (N_12759,N_11774,N_11452);
nor U12760 (N_12760,N_11267,N_11682);
or U12761 (N_12761,N_11848,N_11144);
or U12762 (N_12762,N_11726,N_11023);
nor U12763 (N_12763,N_11372,N_11866);
nor U12764 (N_12764,N_11222,N_11759);
xor U12765 (N_12765,N_11988,N_11163);
nor U12766 (N_12766,N_11442,N_11350);
xnor U12767 (N_12767,N_11751,N_11480);
nand U12768 (N_12768,N_11026,N_11248);
nor U12769 (N_12769,N_11950,N_11574);
and U12770 (N_12770,N_11209,N_11641);
and U12771 (N_12771,N_11584,N_11192);
xnor U12772 (N_12772,N_11159,N_11899);
xnor U12773 (N_12773,N_11246,N_11288);
xor U12774 (N_12774,N_11484,N_11236);
xor U12775 (N_12775,N_11097,N_11182);
xnor U12776 (N_12776,N_11007,N_11470);
or U12777 (N_12777,N_11901,N_11236);
nand U12778 (N_12778,N_11978,N_11781);
and U12779 (N_12779,N_11053,N_11126);
and U12780 (N_12780,N_11459,N_11677);
nor U12781 (N_12781,N_11586,N_11547);
or U12782 (N_12782,N_11817,N_11536);
xnor U12783 (N_12783,N_11066,N_11226);
or U12784 (N_12784,N_11633,N_11249);
xnor U12785 (N_12785,N_11242,N_11338);
nand U12786 (N_12786,N_11394,N_11088);
nand U12787 (N_12787,N_11516,N_11164);
nand U12788 (N_12788,N_11347,N_11722);
and U12789 (N_12789,N_11492,N_11709);
or U12790 (N_12790,N_11193,N_11950);
and U12791 (N_12791,N_11132,N_11238);
xnor U12792 (N_12792,N_11676,N_11953);
and U12793 (N_12793,N_11223,N_11432);
xnor U12794 (N_12794,N_11200,N_11322);
xnor U12795 (N_12795,N_11516,N_11815);
nor U12796 (N_12796,N_11733,N_11589);
nor U12797 (N_12797,N_11549,N_11392);
xnor U12798 (N_12798,N_11959,N_11031);
nand U12799 (N_12799,N_11623,N_11163);
nor U12800 (N_12800,N_11198,N_11932);
xnor U12801 (N_12801,N_11389,N_11852);
and U12802 (N_12802,N_11912,N_11528);
or U12803 (N_12803,N_11802,N_11924);
nor U12804 (N_12804,N_11273,N_11750);
and U12805 (N_12805,N_11795,N_11518);
nand U12806 (N_12806,N_11625,N_11554);
xnor U12807 (N_12807,N_11096,N_11967);
nor U12808 (N_12808,N_11345,N_11222);
xor U12809 (N_12809,N_11963,N_11141);
and U12810 (N_12810,N_11453,N_11175);
and U12811 (N_12811,N_11420,N_11877);
nand U12812 (N_12812,N_11059,N_11530);
xnor U12813 (N_12813,N_11565,N_11545);
xnor U12814 (N_12814,N_11238,N_11392);
nor U12815 (N_12815,N_11961,N_11969);
xnor U12816 (N_12816,N_11084,N_11086);
or U12817 (N_12817,N_11179,N_11762);
and U12818 (N_12818,N_11540,N_11131);
nand U12819 (N_12819,N_11352,N_11539);
or U12820 (N_12820,N_11865,N_11914);
or U12821 (N_12821,N_11501,N_11315);
or U12822 (N_12822,N_11600,N_11457);
and U12823 (N_12823,N_11023,N_11187);
xor U12824 (N_12824,N_11328,N_11820);
nor U12825 (N_12825,N_11595,N_11459);
xor U12826 (N_12826,N_11598,N_11743);
nand U12827 (N_12827,N_11653,N_11284);
xnor U12828 (N_12828,N_11306,N_11564);
nor U12829 (N_12829,N_11331,N_11679);
xnor U12830 (N_12830,N_11222,N_11327);
nor U12831 (N_12831,N_11870,N_11486);
or U12832 (N_12832,N_11031,N_11741);
nand U12833 (N_12833,N_11480,N_11085);
xor U12834 (N_12834,N_11777,N_11687);
and U12835 (N_12835,N_11238,N_11572);
and U12836 (N_12836,N_11481,N_11103);
nor U12837 (N_12837,N_11221,N_11230);
or U12838 (N_12838,N_11438,N_11564);
nand U12839 (N_12839,N_11945,N_11268);
nor U12840 (N_12840,N_11657,N_11747);
nor U12841 (N_12841,N_11202,N_11859);
or U12842 (N_12842,N_11677,N_11079);
xnor U12843 (N_12843,N_11162,N_11301);
xor U12844 (N_12844,N_11485,N_11920);
nor U12845 (N_12845,N_11217,N_11104);
nand U12846 (N_12846,N_11689,N_11577);
nor U12847 (N_12847,N_11489,N_11003);
xnor U12848 (N_12848,N_11234,N_11633);
xor U12849 (N_12849,N_11871,N_11776);
nor U12850 (N_12850,N_11146,N_11295);
nand U12851 (N_12851,N_11776,N_11237);
xor U12852 (N_12852,N_11489,N_11059);
and U12853 (N_12853,N_11166,N_11434);
and U12854 (N_12854,N_11063,N_11922);
nor U12855 (N_12855,N_11799,N_11746);
nand U12856 (N_12856,N_11582,N_11241);
nand U12857 (N_12857,N_11985,N_11221);
nor U12858 (N_12858,N_11578,N_11189);
or U12859 (N_12859,N_11276,N_11009);
and U12860 (N_12860,N_11903,N_11007);
and U12861 (N_12861,N_11989,N_11021);
nand U12862 (N_12862,N_11224,N_11114);
nand U12863 (N_12863,N_11373,N_11958);
nand U12864 (N_12864,N_11448,N_11070);
and U12865 (N_12865,N_11317,N_11412);
nor U12866 (N_12866,N_11644,N_11605);
nor U12867 (N_12867,N_11190,N_11945);
and U12868 (N_12868,N_11799,N_11383);
or U12869 (N_12869,N_11034,N_11442);
xnor U12870 (N_12870,N_11063,N_11990);
nor U12871 (N_12871,N_11467,N_11434);
nor U12872 (N_12872,N_11644,N_11359);
and U12873 (N_12873,N_11348,N_11956);
and U12874 (N_12874,N_11841,N_11038);
or U12875 (N_12875,N_11158,N_11949);
xor U12876 (N_12876,N_11076,N_11387);
nand U12877 (N_12877,N_11194,N_11308);
xnor U12878 (N_12878,N_11588,N_11488);
nor U12879 (N_12879,N_11745,N_11097);
nor U12880 (N_12880,N_11769,N_11912);
xnor U12881 (N_12881,N_11636,N_11771);
or U12882 (N_12882,N_11904,N_11523);
nand U12883 (N_12883,N_11721,N_11785);
nand U12884 (N_12884,N_11123,N_11636);
nor U12885 (N_12885,N_11094,N_11774);
nor U12886 (N_12886,N_11637,N_11305);
or U12887 (N_12887,N_11446,N_11040);
nand U12888 (N_12888,N_11267,N_11464);
nand U12889 (N_12889,N_11316,N_11642);
or U12890 (N_12890,N_11250,N_11724);
and U12891 (N_12891,N_11459,N_11428);
xor U12892 (N_12892,N_11939,N_11426);
and U12893 (N_12893,N_11515,N_11350);
xor U12894 (N_12894,N_11187,N_11355);
xor U12895 (N_12895,N_11462,N_11701);
and U12896 (N_12896,N_11685,N_11455);
nor U12897 (N_12897,N_11548,N_11509);
nand U12898 (N_12898,N_11344,N_11712);
and U12899 (N_12899,N_11180,N_11498);
xor U12900 (N_12900,N_11557,N_11715);
nor U12901 (N_12901,N_11678,N_11144);
and U12902 (N_12902,N_11754,N_11699);
or U12903 (N_12903,N_11988,N_11651);
or U12904 (N_12904,N_11366,N_11006);
and U12905 (N_12905,N_11033,N_11067);
nand U12906 (N_12906,N_11803,N_11233);
xor U12907 (N_12907,N_11601,N_11746);
xor U12908 (N_12908,N_11686,N_11888);
and U12909 (N_12909,N_11374,N_11851);
nor U12910 (N_12910,N_11921,N_11867);
or U12911 (N_12911,N_11790,N_11509);
and U12912 (N_12912,N_11524,N_11146);
nor U12913 (N_12913,N_11912,N_11192);
nand U12914 (N_12914,N_11639,N_11726);
or U12915 (N_12915,N_11239,N_11854);
and U12916 (N_12916,N_11617,N_11321);
nand U12917 (N_12917,N_11900,N_11269);
or U12918 (N_12918,N_11639,N_11698);
nand U12919 (N_12919,N_11724,N_11538);
nor U12920 (N_12920,N_11125,N_11410);
nand U12921 (N_12921,N_11915,N_11884);
or U12922 (N_12922,N_11801,N_11744);
nor U12923 (N_12923,N_11019,N_11831);
nand U12924 (N_12924,N_11755,N_11725);
or U12925 (N_12925,N_11046,N_11770);
nor U12926 (N_12926,N_11003,N_11052);
and U12927 (N_12927,N_11037,N_11080);
nor U12928 (N_12928,N_11686,N_11633);
and U12929 (N_12929,N_11889,N_11816);
or U12930 (N_12930,N_11851,N_11773);
nand U12931 (N_12931,N_11099,N_11679);
xnor U12932 (N_12932,N_11622,N_11422);
and U12933 (N_12933,N_11918,N_11877);
xor U12934 (N_12934,N_11252,N_11329);
or U12935 (N_12935,N_11073,N_11881);
and U12936 (N_12936,N_11689,N_11061);
xor U12937 (N_12937,N_11725,N_11418);
nand U12938 (N_12938,N_11633,N_11651);
or U12939 (N_12939,N_11827,N_11444);
or U12940 (N_12940,N_11292,N_11686);
nor U12941 (N_12941,N_11663,N_11132);
and U12942 (N_12942,N_11729,N_11975);
nand U12943 (N_12943,N_11684,N_11868);
xnor U12944 (N_12944,N_11635,N_11666);
xor U12945 (N_12945,N_11325,N_11226);
nand U12946 (N_12946,N_11195,N_11869);
and U12947 (N_12947,N_11332,N_11553);
xnor U12948 (N_12948,N_11394,N_11945);
nand U12949 (N_12949,N_11620,N_11391);
xnor U12950 (N_12950,N_11983,N_11230);
or U12951 (N_12951,N_11827,N_11872);
nand U12952 (N_12952,N_11646,N_11846);
nor U12953 (N_12953,N_11791,N_11013);
nor U12954 (N_12954,N_11109,N_11954);
nor U12955 (N_12955,N_11836,N_11370);
and U12956 (N_12956,N_11509,N_11469);
and U12957 (N_12957,N_11409,N_11648);
nor U12958 (N_12958,N_11010,N_11913);
and U12959 (N_12959,N_11705,N_11324);
nand U12960 (N_12960,N_11446,N_11791);
or U12961 (N_12961,N_11781,N_11646);
and U12962 (N_12962,N_11732,N_11152);
nand U12963 (N_12963,N_11347,N_11093);
or U12964 (N_12964,N_11461,N_11538);
and U12965 (N_12965,N_11032,N_11761);
or U12966 (N_12966,N_11666,N_11366);
and U12967 (N_12967,N_11648,N_11331);
nor U12968 (N_12968,N_11612,N_11445);
nor U12969 (N_12969,N_11188,N_11984);
and U12970 (N_12970,N_11139,N_11996);
or U12971 (N_12971,N_11707,N_11097);
nor U12972 (N_12972,N_11730,N_11002);
nand U12973 (N_12973,N_11411,N_11094);
and U12974 (N_12974,N_11970,N_11346);
and U12975 (N_12975,N_11602,N_11601);
nor U12976 (N_12976,N_11358,N_11827);
or U12977 (N_12977,N_11129,N_11163);
or U12978 (N_12978,N_11251,N_11360);
nor U12979 (N_12979,N_11643,N_11658);
xnor U12980 (N_12980,N_11228,N_11164);
or U12981 (N_12981,N_11590,N_11671);
or U12982 (N_12982,N_11205,N_11635);
nor U12983 (N_12983,N_11872,N_11633);
nor U12984 (N_12984,N_11146,N_11648);
nand U12985 (N_12985,N_11226,N_11827);
and U12986 (N_12986,N_11506,N_11638);
and U12987 (N_12987,N_11367,N_11011);
xor U12988 (N_12988,N_11937,N_11241);
nand U12989 (N_12989,N_11952,N_11990);
and U12990 (N_12990,N_11604,N_11039);
nor U12991 (N_12991,N_11037,N_11102);
and U12992 (N_12992,N_11375,N_11108);
or U12993 (N_12993,N_11700,N_11216);
nor U12994 (N_12994,N_11368,N_11055);
nor U12995 (N_12995,N_11686,N_11229);
nand U12996 (N_12996,N_11339,N_11190);
nand U12997 (N_12997,N_11299,N_11035);
and U12998 (N_12998,N_11535,N_11605);
xor U12999 (N_12999,N_11513,N_11680);
nor U13000 (N_13000,N_12262,N_12703);
nand U13001 (N_13001,N_12815,N_12868);
and U13002 (N_13002,N_12316,N_12491);
xnor U13003 (N_13003,N_12554,N_12538);
and U13004 (N_13004,N_12921,N_12680);
nand U13005 (N_13005,N_12704,N_12798);
nor U13006 (N_13006,N_12292,N_12970);
nor U13007 (N_13007,N_12080,N_12525);
and U13008 (N_13008,N_12698,N_12419);
and U13009 (N_13009,N_12682,N_12863);
nor U13010 (N_13010,N_12786,N_12655);
or U13011 (N_13011,N_12206,N_12599);
nor U13012 (N_13012,N_12991,N_12629);
and U13013 (N_13013,N_12070,N_12841);
nand U13014 (N_13014,N_12013,N_12595);
xnor U13015 (N_13015,N_12651,N_12090);
xnor U13016 (N_13016,N_12221,N_12039);
xor U13017 (N_13017,N_12318,N_12127);
or U13018 (N_13018,N_12691,N_12010);
nand U13019 (N_13019,N_12839,N_12073);
nand U13020 (N_13020,N_12467,N_12185);
nand U13021 (N_13021,N_12081,N_12353);
or U13022 (N_13022,N_12883,N_12575);
xnor U13023 (N_13023,N_12140,N_12861);
nor U13024 (N_13024,N_12796,N_12279);
or U13025 (N_13025,N_12097,N_12520);
and U13026 (N_13026,N_12373,N_12535);
and U13027 (N_13027,N_12465,N_12674);
nand U13028 (N_13028,N_12986,N_12645);
xnor U13029 (N_13029,N_12952,N_12802);
and U13030 (N_13030,N_12499,N_12440);
nor U13031 (N_13031,N_12893,N_12098);
nand U13032 (N_13032,N_12570,N_12222);
or U13033 (N_13033,N_12055,N_12483);
and U13034 (N_13034,N_12679,N_12082);
or U13035 (N_13035,N_12992,N_12613);
xnor U13036 (N_13036,N_12668,N_12175);
and U13037 (N_13037,N_12038,N_12665);
or U13038 (N_13038,N_12287,N_12845);
and U13039 (N_13039,N_12050,N_12409);
or U13040 (N_13040,N_12226,N_12233);
and U13041 (N_13041,N_12166,N_12650);
nand U13042 (N_13042,N_12450,N_12813);
and U13043 (N_13043,N_12941,N_12909);
and U13044 (N_13044,N_12454,N_12609);
and U13045 (N_13045,N_12623,N_12755);
and U13046 (N_13046,N_12531,N_12980);
nand U13047 (N_13047,N_12943,N_12549);
nor U13048 (N_13048,N_12296,N_12835);
nor U13049 (N_13049,N_12514,N_12299);
or U13050 (N_13050,N_12134,N_12333);
nand U13051 (N_13051,N_12870,N_12572);
xor U13052 (N_13052,N_12319,N_12960);
nor U13053 (N_13053,N_12824,N_12357);
and U13054 (N_13054,N_12740,N_12334);
nand U13055 (N_13055,N_12984,N_12717);
or U13056 (N_13056,N_12005,N_12168);
nand U13057 (N_13057,N_12577,N_12945);
xor U13058 (N_13058,N_12396,N_12302);
and U13059 (N_13059,N_12508,N_12335);
nor U13060 (N_13060,N_12643,N_12751);
xor U13061 (N_13061,N_12593,N_12632);
nor U13062 (N_13062,N_12042,N_12120);
and U13063 (N_13063,N_12722,N_12971);
nor U13064 (N_13064,N_12585,N_12817);
and U13065 (N_13065,N_12821,N_12877);
nor U13066 (N_13066,N_12311,N_12076);
nand U13067 (N_13067,N_12582,N_12580);
nor U13068 (N_13068,N_12460,N_12425);
nor U13069 (N_13069,N_12488,N_12383);
and U13070 (N_13070,N_12181,N_12170);
nor U13071 (N_13071,N_12763,N_12126);
nor U13072 (N_13072,N_12154,N_12325);
or U13073 (N_13073,N_12563,N_12115);
nor U13074 (N_13074,N_12114,N_12551);
and U13075 (N_13075,N_12244,N_12118);
nand U13076 (N_13076,N_12972,N_12574);
nor U13077 (N_13077,N_12735,N_12283);
and U13078 (N_13078,N_12162,N_12420);
and U13079 (N_13079,N_12374,N_12102);
and U13080 (N_13080,N_12035,N_12280);
nor U13081 (N_13081,N_12928,N_12686);
or U13082 (N_13082,N_12022,N_12478);
nand U13083 (N_13083,N_12128,N_12300);
nand U13084 (N_13084,N_12509,N_12477);
or U13085 (N_13085,N_12112,N_12875);
nand U13086 (N_13086,N_12539,N_12922);
nand U13087 (N_13087,N_12489,N_12034);
xor U13088 (N_13088,N_12148,N_12809);
or U13089 (N_13089,N_12129,N_12231);
and U13090 (N_13090,N_12448,N_12392);
xnor U13091 (N_13091,N_12537,N_12003);
xor U13092 (N_13092,N_12130,N_12739);
or U13093 (N_13093,N_12495,N_12581);
or U13094 (N_13094,N_12517,N_12339);
and U13095 (N_13095,N_12219,N_12622);
and U13096 (N_13096,N_12726,N_12471);
xnor U13097 (N_13097,N_12548,N_12664);
or U13098 (N_13098,N_12503,N_12286);
and U13099 (N_13099,N_12345,N_12519);
nor U13100 (N_13100,N_12201,N_12305);
xor U13101 (N_13101,N_12193,N_12721);
nor U13102 (N_13102,N_12442,N_12436);
xnor U13103 (N_13103,N_12230,N_12844);
nor U13104 (N_13104,N_12406,N_12389);
nand U13105 (N_13105,N_12935,N_12167);
nand U13106 (N_13106,N_12249,N_12387);
nor U13107 (N_13107,N_12513,N_12094);
nand U13108 (N_13108,N_12207,N_12312);
or U13109 (N_13109,N_12269,N_12638);
and U13110 (N_13110,N_12072,N_12901);
or U13111 (N_13111,N_12526,N_12764);
xor U13112 (N_13112,N_12304,N_12153);
xor U13113 (N_13113,N_12368,N_12033);
or U13114 (N_13114,N_12736,N_12036);
or U13115 (N_13115,N_12028,N_12957);
xnor U13116 (N_13116,N_12847,N_12902);
or U13117 (N_13117,N_12485,N_12025);
nor U13118 (N_13118,N_12745,N_12395);
nor U13119 (N_13119,N_12246,N_12214);
and U13120 (N_13120,N_12248,N_12079);
nand U13121 (N_13121,N_12662,N_12948);
nor U13122 (N_13122,N_12779,N_12053);
or U13123 (N_13123,N_12136,N_12458);
xnor U13124 (N_13124,N_12349,N_12242);
or U13125 (N_13125,N_12727,N_12288);
or U13126 (N_13126,N_12566,N_12694);
xor U13127 (N_13127,N_12274,N_12794);
and U13128 (N_13128,N_12133,N_12761);
nor U13129 (N_13129,N_12051,N_12189);
xnor U13130 (N_13130,N_12838,N_12329);
or U13131 (N_13131,N_12423,N_12731);
xor U13132 (N_13132,N_12336,N_12507);
and U13133 (N_13133,N_12927,N_12437);
xnor U13134 (N_13134,N_12697,N_12894);
or U13135 (N_13135,N_12381,N_12007);
nor U13136 (N_13136,N_12372,N_12530);
xnor U13137 (N_13137,N_12769,N_12669);
nand U13138 (N_13138,N_12770,N_12444);
and U13139 (N_13139,N_12546,N_12752);
nand U13140 (N_13140,N_12108,N_12846);
or U13141 (N_13141,N_12684,N_12424);
nand U13142 (N_13142,N_12364,N_12994);
and U13143 (N_13143,N_12936,N_12734);
or U13144 (N_13144,N_12216,N_12270);
nor U13145 (N_13145,N_12621,N_12848);
and U13146 (N_13146,N_12502,N_12597);
and U13147 (N_13147,N_12188,N_12382);
nand U13148 (N_13148,N_12750,N_12925);
xnor U13149 (N_13149,N_12330,N_12250);
xor U13150 (N_13150,N_12856,N_12583);
and U13151 (N_13151,N_12399,N_12031);
or U13152 (N_13152,N_12807,N_12947);
and U13153 (N_13153,N_12747,N_12552);
nor U13154 (N_13154,N_12592,N_12482);
nand U13155 (N_13155,N_12152,N_12604);
and U13156 (N_13156,N_12203,N_12121);
nand U13157 (N_13157,N_12606,N_12047);
nand U13158 (N_13158,N_12759,N_12787);
or U13159 (N_13159,N_12982,N_12619);
or U13160 (N_13160,N_12317,N_12874);
nor U13161 (N_13161,N_12290,N_12378);
and U13162 (N_13162,N_12869,N_12481);
and U13163 (N_13163,N_12681,N_12147);
or U13164 (N_13164,N_12107,N_12493);
or U13165 (N_13165,N_12562,N_12394);
xnor U13166 (N_13166,N_12565,N_12295);
or U13167 (N_13167,N_12032,N_12511);
nand U13168 (N_13168,N_12522,N_12777);
xnor U13169 (N_13169,N_12365,N_12431);
or U13170 (N_13170,N_12393,N_12291);
nand U13171 (N_13171,N_12975,N_12321);
nor U13172 (N_13172,N_12161,N_12989);
nor U13173 (N_13173,N_12658,N_12271);
xnor U13174 (N_13174,N_12560,N_12920);
or U13175 (N_13175,N_12995,N_12781);
nand U13176 (N_13176,N_12433,N_12117);
nand U13177 (N_13177,N_12294,N_12545);
nor U13178 (N_13178,N_12576,N_12380);
nor U13179 (N_13179,N_12654,N_12146);
xor U13180 (N_13180,N_12404,N_12195);
xnor U13181 (N_13181,N_12640,N_12008);
nand U13182 (N_13182,N_12924,N_12462);
nor U13183 (N_13183,N_12015,N_12176);
and U13184 (N_13184,N_12852,N_12265);
and U13185 (N_13185,N_12347,N_12182);
and U13186 (N_13186,N_12940,N_12806);
nand U13187 (N_13187,N_12111,N_12385);
or U13188 (N_13188,N_12801,N_12155);
nand U13189 (N_13189,N_12765,N_12964);
xor U13190 (N_13190,N_12137,N_12463);
or U13191 (N_13191,N_12174,N_12962);
xnor U13192 (N_13192,N_12904,N_12422);
and U13193 (N_13193,N_12238,N_12190);
or U13194 (N_13194,N_12307,N_12067);
nand U13195 (N_13195,N_12093,N_12427);
nor U13196 (N_13196,N_12931,N_12479);
nand U13197 (N_13197,N_12515,N_12224);
nor U13198 (N_13198,N_12790,N_12359);
xor U13199 (N_13199,N_12435,N_12879);
and U13200 (N_13200,N_12284,N_12521);
xnor U13201 (N_13201,N_12949,N_12625);
or U13202 (N_13202,N_12278,N_12832);
or U13203 (N_13203,N_12607,N_12834);
and U13204 (N_13204,N_12403,N_12961);
nand U13205 (N_13205,N_12315,N_12459);
and U13206 (N_13206,N_12884,N_12990);
nor U13207 (N_13207,N_12159,N_12470);
nand U13208 (N_13208,N_12797,N_12601);
nand U13209 (N_13209,N_12528,N_12512);
nor U13210 (N_13210,N_12612,N_12062);
nand U13211 (N_13211,N_12211,N_12075);
nand U13212 (N_13212,N_12516,N_12376);
nand U13213 (N_13213,N_12194,N_12830);
xnor U13214 (N_13214,N_12938,N_12309);
nand U13215 (N_13215,N_12784,N_12687);
or U13216 (N_13216,N_12390,N_12840);
nand U13217 (N_13217,N_12569,N_12343);
and U13218 (N_13218,N_12873,N_12466);
xnor U13219 (N_13219,N_12445,N_12584);
or U13220 (N_13220,N_12354,N_12639);
xnor U13221 (N_13221,N_12441,N_12125);
nand U13222 (N_13222,N_12710,N_12012);
nand U13223 (N_13223,N_12139,N_12124);
and U13224 (N_13224,N_12110,N_12266);
xor U13225 (N_13225,N_12558,N_12586);
and U13226 (N_13226,N_12149,N_12542);
xnor U13227 (N_13227,N_12054,N_12232);
xor U13228 (N_13228,N_12864,N_12808);
nand U13229 (N_13229,N_12375,N_12965);
and U13230 (N_13230,N_12910,N_12065);
xor U13231 (N_13231,N_12472,N_12780);
xor U13232 (N_13232,N_12892,N_12059);
and U13233 (N_13233,N_12138,N_12527);
and U13234 (N_13234,N_12898,N_12878);
nor U13235 (N_13235,N_12760,N_12297);
nand U13236 (N_13236,N_12496,N_12078);
xnor U13237 (N_13237,N_12741,N_12918);
xnor U13238 (N_13238,N_12827,N_12712);
and U13239 (N_13239,N_12122,N_12273);
xor U13240 (N_13240,N_12532,N_12713);
xnor U13241 (N_13241,N_12135,N_12657);
nand U13242 (N_13242,N_12708,N_12473);
or U13243 (N_13243,N_12851,N_12618);
nor U13244 (N_13244,N_12733,N_12023);
and U13245 (N_13245,N_12652,N_12958);
xnor U13246 (N_13246,N_12430,N_12020);
or U13247 (N_13247,N_12087,N_12896);
nor U13248 (N_13248,N_12324,N_12701);
or U13249 (N_13249,N_12700,N_12872);
nand U13250 (N_13250,N_12706,N_12282);
or U13251 (N_13251,N_12589,N_12092);
or U13252 (N_13252,N_12408,N_12105);
or U13253 (N_13253,N_12037,N_12578);
xor U13254 (N_13254,N_12644,N_12268);
nand U13255 (N_13255,N_12646,N_12800);
and U13256 (N_13256,N_12886,N_12084);
xnor U13257 (N_13257,N_12142,N_12002);
and U13258 (N_13258,N_12338,N_12457);
xor U13259 (N_13259,N_12171,N_12150);
nand U13260 (N_13260,N_12379,N_12064);
nor U13261 (N_13261,N_12659,N_12942);
or U13262 (N_13262,N_12843,N_12702);
nand U13263 (N_13263,N_12398,N_12447);
nor U13264 (N_13264,N_12748,N_12647);
xnor U13265 (N_13265,N_12151,N_12919);
or U13266 (N_13266,N_12636,N_12591);
xor U13267 (N_13267,N_12377,N_12497);
or U13268 (N_13268,N_12160,N_12068);
nand U13269 (N_13269,N_12308,N_12344);
xor U13270 (N_13270,N_12649,N_12428);
and U13271 (N_13271,N_12814,N_12077);
or U13272 (N_13272,N_12220,N_12453);
nor U13273 (N_13273,N_12215,N_12363);
and U13274 (N_13274,N_12783,N_12811);
nand U13275 (N_13275,N_12416,N_12985);
xnor U13276 (N_13276,N_12825,N_12568);
and U13277 (N_13277,N_12716,N_12446);
and U13278 (N_13278,N_12685,N_12907);
and U13279 (N_13279,N_12556,N_12871);
nand U13280 (N_13280,N_12810,N_12561);
nand U13281 (N_13281,N_12983,N_12218);
nand U13282 (N_13282,N_12069,N_12116);
or U13283 (N_13283,N_12772,N_12199);
xor U13284 (N_13284,N_12474,N_12086);
or U13285 (N_13285,N_12778,N_12768);
nand U13286 (N_13286,N_12045,N_12754);
nand U13287 (N_13287,N_12724,N_12326);
or U13288 (N_13288,N_12775,N_12746);
nor U13289 (N_13289,N_12163,N_12946);
nor U13290 (N_13290,N_12004,N_12923);
and U13291 (N_13291,N_12822,N_12251);
and U13292 (N_13292,N_12854,N_12074);
and U13293 (N_13293,N_12819,N_12384);
nor U13294 (N_13294,N_12944,N_12988);
and U13295 (N_13295,N_12720,N_12977);
xor U13296 (N_13296,N_12916,N_12277);
xor U13297 (N_13297,N_12314,N_12366);
and U13298 (N_13298,N_12667,N_12881);
nand U13299 (N_13299,N_12719,N_12429);
nor U13300 (N_13300,N_12917,N_12298);
xor U13301 (N_13301,N_12504,N_12782);
or U13302 (N_13302,N_12937,N_12805);
nor U13303 (N_13303,N_12564,N_12633);
nor U13304 (N_13304,N_12434,N_12723);
nand U13305 (N_13305,N_12738,N_12743);
nand U13306 (N_13306,N_12494,N_12099);
xnor U13307 (N_13307,N_12006,N_12867);
xnor U13308 (N_13308,N_12891,N_12888);
or U13309 (N_13309,N_12293,N_12276);
nand U13310 (N_13310,N_12415,N_12753);
xnor U13311 (N_13311,N_12860,N_12468);
nand U13312 (N_13312,N_12241,N_12411);
and U13313 (N_13313,N_12289,N_12967);
or U13314 (N_13314,N_12024,N_12518);
and U13315 (N_13315,N_12355,N_12027);
and U13316 (N_13316,N_12410,N_12475);
nand U13317 (N_13317,N_12367,N_12693);
xnor U13318 (N_13318,N_12930,N_12200);
and U13319 (N_13319,N_12011,N_12208);
nor U13320 (N_13320,N_12849,N_12063);
and U13321 (N_13321,N_12158,N_12223);
nand U13322 (N_13322,N_12058,N_12362);
or U13323 (N_13323,N_12959,N_12788);
or U13324 (N_13324,N_12795,N_12642);
and U13325 (N_13325,N_12456,N_12187);
nand U13326 (N_13326,N_12313,N_12978);
or U13327 (N_13327,N_12974,N_12956);
and U13328 (N_13328,N_12275,N_12085);
xnor U13329 (N_13329,N_12091,N_12254);
xnor U13330 (N_13330,N_12263,N_12332);
nand U13331 (N_13331,N_12145,N_12536);
nor U13332 (N_13332,N_12837,N_12903);
and U13333 (N_13333,N_12976,N_12631);
xor U13334 (N_13334,N_12661,N_12842);
nor U13335 (N_13335,N_12486,N_12178);
or U13336 (N_13336,N_12157,N_12183);
or U13337 (N_13337,N_12829,N_12057);
xnor U13338 (N_13338,N_12413,N_12331);
nand U13339 (N_13339,N_12998,N_12596);
and U13340 (N_13340,N_12767,N_12337);
nand U13341 (N_13341,N_12954,N_12202);
nor U13342 (N_13342,N_12043,N_12533);
xnor U13343 (N_13343,N_12156,N_12401);
nor U13344 (N_13344,N_12113,N_12323);
and U13345 (N_13345,N_12826,N_12934);
nor U13346 (N_13346,N_12432,N_12831);
nor U13347 (N_13347,N_12310,N_12557);
xnor U13348 (N_13348,N_12358,N_12529);
nand U13349 (N_13349,N_12227,N_12555);
xor U13350 (N_13350,N_12993,N_12553);
xnor U13351 (N_13351,N_12885,N_12953);
and U13352 (N_13352,N_12132,N_12418);
xor U13353 (N_13353,N_12550,N_12255);
and U13354 (N_13354,N_12887,N_12253);
nor U13355 (N_13355,N_12610,N_12240);
nor U13356 (N_13356,N_12352,N_12257);
and U13357 (N_13357,N_12912,N_12019);
and U13358 (N_13358,N_12348,N_12616);
and U13359 (N_13359,N_12041,N_12600);
and U13360 (N_13360,N_12350,N_12191);
and U13361 (N_13361,N_12342,N_12212);
nand U13362 (N_13362,N_12198,N_12973);
and U13363 (N_13363,N_12803,N_12501);
nor U13364 (N_13364,N_12547,N_12452);
and U13365 (N_13365,N_12793,N_12758);
nand U13366 (N_13366,N_12611,N_12523);
and U13367 (N_13367,N_12997,N_12234);
and U13368 (N_13368,N_12812,N_12179);
xor U13369 (N_13369,N_12172,N_12505);
xnor U13370 (N_13370,N_12672,N_12624);
and U13371 (N_13371,N_12370,N_12356);
nand U13372 (N_13372,N_12966,N_12400);
and U13373 (N_13373,N_12267,N_12071);
nand U13374 (N_13374,N_12260,N_12524);
xor U13375 (N_13375,N_12637,N_12026);
nor U13376 (N_13376,N_12728,N_12361);
and U13377 (N_13377,N_12707,N_12256);
and U13378 (N_13378,N_12897,N_12774);
nand U13379 (N_13379,N_12438,N_12673);
xor U13380 (N_13380,N_12030,N_12715);
nand U13381 (N_13381,N_12173,N_12950);
nand U13382 (N_13382,N_12169,N_12048);
nor U13383 (N_13383,N_12913,N_12000);
or U13384 (N_13384,N_12890,N_12052);
or U13385 (N_13385,N_12029,N_12484);
nor U13386 (N_13386,N_12303,N_12951);
nand U13387 (N_13387,N_12857,N_12259);
and U13388 (N_13388,N_12705,N_12165);
xnor U13389 (N_13389,N_12939,N_12590);
nand U13390 (N_13390,N_12828,N_12369);
or U13391 (N_13391,N_12534,N_12689);
nor U13392 (N_13392,N_12285,N_12602);
xor U13393 (N_13393,N_12627,N_12725);
nor U13394 (N_13394,N_12776,N_12742);
xor U13395 (N_13395,N_12653,N_12184);
xnor U13396 (N_13396,N_12926,N_12328);
xor U13397 (N_13397,N_12677,N_12101);
nand U13398 (N_13398,N_12177,N_12678);
nand U13399 (N_13399,N_12660,N_12785);
or U13400 (N_13400,N_12046,N_12690);
or U13401 (N_13401,N_12327,N_12608);
nand U13402 (N_13402,N_12594,N_12180);
nor U13403 (N_13403,N_12141,N_12351);
or U13404 (N_13404,N_12209,N_12749);
nand U13405 (N_13405,N_12213,N_12617);
or U13406 (N_13406,N_12882,N_12088);
xor U13407 (N_13407,N_12963,N_12889);
xor U13408 (N_13408,N_12696,N_12480);
xor U13409 (N_13409,N_12588,N_12692);
or U13410 (N_13410,N_12634,N_12143);
xnor U13411 (N_13411,N_12421,N_12487);
nand U13412 (N_13412,N_12932,N_12855);
and U13413 (N_13413,N_12630,N_12833);
nand U13414 (N_13414,N_12322,N_12414);
or U13415 (N_13415,N_12235,N_12217);
and U13416 (N_13416,N_12862,N_12492);
and U13417 (N_13417,N_12320,N_12164);
or U13418 (N_13418,N_12605,N_12104);
nand U13419 (N_13419,N_12009,N_12301);
xnor U13420 (N_13420,N_12229,N_12709);
nand U13421 (N_13421,N_12103,N_12899);
or U13422 (N_13422,N_12853,N_12264);
and U13423 (N_13423,N_12587,N_12464);
nor U13424 (N_13424,N_12017,N_12670);
nand U13425 (N_13425,N_12981,N_12573);
nor U13426 (N_13426,N_12858,N_12391);
nand U13427 (N_13427,N_12018,N_12598);
and U13428 (N_13428,N_12791,N_12131);
and U13429 (N_13429,N_12915,N_12210);
or U13430 (N_13430,N_12955,N_12490);
and U13431 (N_13431,N_12979,N_12061);
and U13432 (N_13432,N_12820,N_12186);
or U13433 (N_13433,N_12196,N_12818);
and U13434 (N_13434,N_12744,N_12968);
xor U13435 (N_13435,N_12407,N_12641);
and U13436 (N_13436,N_12237,N_12245);
or U13437 (N_13437,N_12044,N_12771);
xor U13438 (N_13438,N_12439,N_12614);
or U13439 (N_13439,N_12272,N_12247);
nor U13440 (N_13440,N_12461,N_12239);
nor U13441 (N_13441,N_12757,N_12900);
or U13442 (N_13442,N_12192,N_12197);
and U13443 (N_13443,N_12066,N_12397);
and U13444 (N_13444,N_12730,N_12014);
and U13445 (N_13445,N_12695,N_12106);
nor U13446 (N_13446,N_12766,N_12671);
and U13447 (N_13447,N_12865,N_12756);
or U13448 (N_13448,N_12498,N_12729);
nor U13449 (N_13449,N_12620,N_12850);
or U13450 (N_13450,N_12049,N_12500);
nor U13451 (N_13451,N_12906,N_12675);
and U13452 (N_13452,N_12449,N_12123);
xnor U13453 (N_13453,N_12252,N_12683);
or U13454 (N_13454,N_12083,N_12100);
nor U13455 (N_13455,N_12880,N_12243);
xor U13456 (N_13456,N_12417,N_12628);
and U13457 (N_13457,N_12096,N_12914);
or U13458 (N_13458,N_12228,N_12799);
xor U13459 (N_13459,N_12543,N_12340);
nor U13460 (N_13460,N_12789,N_12999);
nand U13461 (N_13461,N_12908,N_12089);
and U13462 (N_13462,N_12426,N_12021);
xor U13463 (N_13463,N_12455,N_12016);
and U13464 (N_13464,N_12060,N_12933);
nand U13465 (N_13465,N_12371,N_12402);
nor U13466 (N_13466,N_12895,N_12929);
and U13467 (N_13467,N_12714,N_12540);
nand U13468 (N_13468,N_12443,N_12119);
xnor U13469 (N_13469,N_12205,N_12969);
nor U13470 (N_13470,N_12911,N_12699);
and U13471 (N_13471,N_12510,N_12476);
xnor U13472 (N_13472,N_12905,N_12656);
nor U13473 (N_13473,N_12204,N_12506);
nor U13474 (N_13474,N_12663,N_12109);
nand U13475 (N_13475,N_12341,N_12346);
nand U13476 (N_13476,N_12732,N_12258);
and U13477 (N_13477,N_12866,N_12571);
xor U13478 (N_13478,N_12996,N_12635);
and U13479 (N_13479,N_12144,N_12876);
nor U13480 (N_13480,N_12823,N_12762);
xor U13481 (N_13481,N_12095,N_12676);
and U13482 (N_13482,N_12541,N_12603);
and U13483 (N_13483,N_12412,N_12737);
xnor U13484 (N_13484,N_12388,N_12626);
and U13485 (N_13485,N_12666,N_12804);
nor U13486 (N_13486,N_12451,N_12648);
nand U13487 (N_13487,N_12386,N_12236);
or U13488 (N_13488,N_12306,N_12859);
xor U13489 (N_13489,N_12773,N_12711);
and U13490 (N_13490,N_12360,N_12001);
and U13491 (N_13491,N_12615,N_12836);
nand U13492 (N_13492,N_12405,N_12040);
xnor U13493 (N_13493,N_12544,N_12056);
and U13494 (N_13494,N_12816,N_12792);
xnor U13495 (N_13495,N_12579,N_12688);
or U13496 (N_13496,N_12469,N_12718);
nor U13497 (N_13497,N_12987,N_12559);
nand U13498 (N_13498,N_12281,N_12225);
nor U13499 (N_13499,N_12567,N_12261);
xnor U13500 (N_13500,N_12237,N_12000);
and U13501 (N_13501,N_12596,N_12443);
or U13502 (N_13502,N_12333,N_12150);
or U13503 (N_13503,N_12439,N_12121);
xor U13504 (N_13504,N_12633,N_12998);
nand U13505 (N_13505,N_12074,N_12893);
xor U13506 (N_13506,N_12549,N_12065);
and U13507 (N_13507,N_12913,N_12764);
or U13508 (N_13508,N_12685,N_12880);
and U13509 (N_13509,N_12184,N_12079);
nand U13510 (N_13510,N_12379,N_12643);
or U13511 (N_13511,N_12977,N_12633);
nor U13512 (N_13512,N_12708,N_12135);
nor U13513 (N_13513,N_12502,N_12453);
or U13514 (N_13514,N_12761,N_12711);
xnor U13515 (N_13515,N_12800,N_12215);
xor U13516 (N_13516,N_12863,N_12679);
nand U13517 (N_13517,N_12167,N_12770);
and U13518 (N_13518,N_12702,N_12570);
nand U13519 (N_13519,N_12346,N_12935);
xnor U13520 (N_13520,N_12383,N_12517);
xnor U13521 (N_13521,N_12048,N_12781);
or U13522 (N_13522,N_12834,N_12267);
and U13523 (N_13523,N_12177,N_12225);
or U13524 (N_13524,N_12068,N_12261);
and U13525 (N_13525,N_12613,N_12328);
or U13526 (N_13526,N_12332,N_12589);
nand U13527 (N_13527,N_12393,N_12824);
xnor U13528 (N_13528,N_12299,N_12177);
and U13529 (N_13529,N_12699,N_12084);
and U13530 (N_13530,N_12962,N_12396);
xnor U13531 (N_13531,N_12954,N_12500);
xor U13532 (N_13532,N_12250,N_12626);
and U13533 (N_13533,N_12719,N_12541);
nor U13534 (N_13534,N_12323,N_12936);
or U13535 (N_13535,N_12508,N_12476);
nor U13536 (N_13536,N_12862,N_12387);
xnor U13537 (N_13537,N_12992,N_12944);
xnor U13538 (N_13538,N_12195,N_12545);
nand U13539 (N_13539,N_12009,N_12237);
nand U13540 (N_13540,N_12059,N_12598);
and U13541 (N_13541,N_12362,N_12766);
or U13542 (N_13542,N_12613,N_12757);
or U13543 (N_13543,N_12407,N_12736);
and U13544 (N_13544,N_12958,N_12743);
or U13545 (N_13545,N_12652,N_12355);
or U13546 (N_13546,N_12782,N_12356);
nor U13547 (N_13547,N_12640,N_12419);
nor U13548 (N_13548,N_12070,N_12136);
nand U13549 (N_13549,N_12320,N_12736);
nand U13550 (N_13550,N_12755,N_12264);
nand U13551 (N_13551,N_12289,N_12739);
or U13552 (N_13552,N_12285,N_12939);
nand U13553 (N_13553,N_12259,N_12699);
nand U13554 (N_13554,N_12054,N_12943);
nand U13555 (N_13555,N_12797,N_12232);
or U13556 (N_13556,N_12137,N_12895);
nor U13557 (N_13557,N_12553,N_12546);
nor U13558 (N_13558,N_12007,N_12899);
and U13559 (N_13559,N_12898,N_12965);
or U13560 (N_13560,N_12993,N_12758);
nor U13561 (N_13561,N_12541,N_12839);
and U13562 (N_13562,N_12156,N_12445);
and U13563 (N_13563,N_12765,N_12137);
and U13564 (N_13564,N_12966,N_12024);
nor U13565 (N_13565,N_12404,N_12569);
nand U13566 (N_13566,N_12526,N_12250);
or U13567 (N_13567,N_12797,N_12201);
xnor U13568 (N_13568,N_12559,N_12604);
nand U13569 (N_13569,N_12756,N_12698);
nor U13570 (N_13570,N_12318,N_12136);
and U13571 (N_13571,N_12369,N_12919);
or U13572 (N_13572,N_12901,N_12349);
nor U13573 (N_13573,N_12204,N_12973);
and U13574 (N_13574,N_12948,N_12873);
nor U13575 (N_13575,N_12949,N_12229);
nor U13576 (N_13576,N_12456,N_12913);
xnor U13577 (N_13577,N_12195,N_12970);
nand U13578 (N_13578,N_12108,N_12061);
or U13579 (N_13579,N_12719,N_12986);
and U13580 (N_13580,N_12042,N_12184);
or U13581 (N_13581,N_12648,N_12829);
nor U13582 (N_13582,N_12211,N_12243);
nor U13583 (N_13583,N_12857,N_12119);
and U13584 (N_13584,N_12211,N_12792);
or U13585 (N_13585,N_12691,N_12568);
xnor U13586 (N_13586,N_12819,N_12608);
or U13587 (N_13587,N_12162,N_12051);
and U13588 (N_13588,N_12433,N_12413);
nand U13589 (N_13589,N_12511,N_12316);
nand U13590 (N_13590,N_12688,N_12960);
or U13591 (N_13591,N_12035,N_12100);
xnor U13592 (N_13592,N_12530,N_12797);
xor U13593 (N_13593,N_12142,N_12216);
or U13594 (N_13594,N_12758,N_12604);
nor U13595 (N_13595,N_12469,N_12926);
nor U13596 (N_13596,N_12155,N_12891);
nand U13597 (N_13597,N_12766,N_12220);
and U13598 (N_13598,N_12091,N_12798);
xor U13599 (N_13599,N_12983,N_12512);
and U13600 (N_13600,N_12542,N_12511);
xor U13601 (N_13601,N_12557,N_12550);
and U13602 (N_13602,N_12891,N_12172);
nand U13603 (N_13603,N_12052,N_12798);
xnor U13604 (N_13604,N_12697,N_12115);
nor U13605 (N_13605,N_12077,N_12473);
or U13606 (N_13606,N_12048,N_12415);
nor U13607 (N_13607,N_12254,N_12017);
or U13608 (N_13608,N_12879,N_12399);
or U13609 (N_13609,N_12699,N_12743);
or U13610 (N_13610,N_12800,N_12542);
or U13611 (N_13611,N_12695,N_12438);
and U13612 (N_13612,N_12905,N_12802);
and U13613 (N_13613,N_12663,N_12525);
nand U13614 (N_13614,N_12787,N_12851);
and U13615 (N_13615,N_12568,N_12308);
nand U13616 (N_13616,N_12182,N_12919);
and U13617 (N_13617,N_12907,N_12644);
nor U13618 (N_13618,N_12635,N_12379);
xor U13619 (N_13619,N_12449,N_12145);
and U13620 (N_13620,N_12925,N_12181);
nor U13621 (N_13621,N_12803,N_12820);
and U13622 (N_13622,N_12103,N_12973);
nor U13623 (N_13623,N_12459,N_12440);
or U13624 (N_13624,N_12182,N_12747);
and U13625 (N_13625,N_12737,N_12692);
or U13626 (N_13626,N_12149,N_12101);
xor U13627 (N_13627,N_12322,N_12875);
xnor U13628 (N_13628,N_12836,N_12722);
xor U13629 (N_13629,N_12184,N_12390);
nand U13630 (N_13630,N_12837,N_12518);
and U13631 (N_13631,N_12962,N_12454);
and U13632 (N_13632,N_12643,N_12418);
and U13633 (N_13633,N_12303,N_12095);
xnor U13634 (N_13634,N_12216,N_12146);
nor U13635 (N_13635,N_12348,N_12937);
nor U13636 (N_13636,N_12620,N_12601);
and U13637 (N_13637,N_12653,N_12892);
and U13638 (N_13638,N_12595,N_12489);
nand U13639 (N_13639,N_12676,N_12534);
nand U13640 (N_13640,N_12209,N_12178);
nand U13641 (N_13641,N_12029,N_12409);
and U13642 (N_13642,N_12003,N_12093);
nand U13643 (N_13643,N_12098,N_12794);
xor U13644 (N_13644,N_12654,N_12663);
xor U13645 (N_13645,N_12265,N_12124);
xnor U13646 (N_13646,N_12618,N_12534);
and U13647 (N_13647,N_12512,N_12423);
nor U13648 (N_13648,N_12155,N_12135);
xor U13649 (N_13649,N_12768,N_12351);
nor U13650 (N_13650,N_12268,N_12027);
nand U13651 (N_13651,N_12199,N_12943);
or U13652 (N_13652,N_12265,N_12579);
xor U13653 (N_13653,N_12768,N_12032);
xnor U13654 (N_13654,N_12070,N_12268);
nor U13655 (N_13655,N_12740,N_12379);
nor U13656 (N_13656,N_12555,N_12152);
nor U13657 (N_13657,N_12348,N_12659);
nor U13658 (N_13658,N_12063,N_12582);
nor U13659 (N_13659,N_12621,N_12870);
and U13660 (N_13660,N_12644,N_12899);
nand U13661 (N_13661,N_12186,N_12427);
or U13662 (N_13662,N_12568,N_12157);
nor U13663 (N_13663,N_12465,N_12841);
xnor U13664 (N_13664,N_12172,N_12239);
and U13665 (N_13665,N_12145,N_12194);
nor U13666 (N_13666,N_12381,N_12679);
and U13667 (N_13667,N_12981,N_12461);
xor U13668 (N_13668,N_12163,N_12405);
or U13669 (N_13669,N_12361,N_12293);
and U13670 (N_13670,N_12310,N_12832);
nor U13671 (N_13671,N_12009,N_12156);
nor U13672 (N_13672,N_12553,N_12348);
nor U13673 (N_13673,N_12529,N_12162);
or U13674 (N_13674,N_12019,N_12498);
nor U13675 (N_13675,N_12709,N_12199);
or U13676 (N_13676,N_12569,N_12697);
and U13677 (N_13677,N_12830,N_12234);
or U13678 (N_13678,N_12093,N_12871);
or U13679 (N_13679,N_12414,N_12314);
nor U13680 (N_13680,N_12204,N_12097);
or U13681 (N_13681,N_12763,N_12176);
xor U13682 (N_13682,N_12990,N_12474);
xnor U13683 (N_13683,N_12550,N_12442);
or U13684 (N_13684,N_12901,N_12861);
xor U13685 (N_13685,N_12513,N_12821);
nor U13686 (N_13686,N_12762,N_12414);
nand U13687 (N_13687,N_12097,N_12931);
nand U13688 (N_13688,N_12099,N_12672);
and U13689 (N_13689,N_12175,N_12643);
and U13690 (N_13690,N_12182,N_12258);
xnor U13691 (N_13691,N_12906,N_12419);
nor U13692 (N_13692,N_12899,N_12780);
nand U13693 (N_13693,N_12916,N_12850);
or U13694 (N_13694,N_12872,N_12328);
xnor U13695 (N_13695,N_12987,N_12354);
or U13696 (N_13696,N_12934,N_12288);
and U13697 (N_13697,N_12135,N_12157);
nor U13698 (N_13698,N_12365,N_12267);
nor U13699 (N_13699,N_12966,N_12074);
nand U13700 (N_13700,N_12480,N_12100);
nor U13701 (N_13701,N_12583,N_12852);
nand U13702 (N_13702,N_12622,N_12833);
nor U13703 (N_13703,N_12073,N_12863);
nand U13704 (N_13704,N_12623,N_12351);
nand U13705 (N_13705,N_12143,N_12833);
nor U13706 (N_13706,N_12844,N_12637);
or U13707 (N_13707,N_12184,N_12915);
or U13708 (N_13708,N_12910,N_12515);
or U13709 (N_13709,N_12289,N_12974);
nor U13710 (N_13710,N_12885,N_12164);
xnor U13711 (N_13711,N_12228,N_12052);
or U13712 (N_13712,N_12194,N_12491);
nor U13713 (N_13713,N_12349,N_12032);
xnor U13714 (N_13714,N_12403,N_12314);
xor U13715 (N_13715,N_12775,N_12247);
nor U13716 (N_13716,N_12557,N_12952);
nor U13717 (N_13717,N_12007,N_12280);
nand U13718 (N_13718,N_12955,N_12064);
or U13719 (N_13719,N_12020,N_12242);
or U13720 (N_13720,N_12056,N_12147);
xnor U13721 (N_13721,N_12776,N_12065);
or U13722 (N_13722,N_12035,N_12869);
nor U13723 (N_13723,N_12917,N_12784);
or U13724 (N_13724,N_12618,N_12978);
xnor U13725 (N_13725,N_12245,N_12644);
nand U13726 (N_13726,N_12592,N_12167);
or U13727 (N_13727,N_12984,N_12925);
xnor U13728 (N_13728,N_12835,N_12162);
nor U13729 (N_13729,N_12177,N_12063);
xor U13730 (N_13730,N_12085,N_12778);
xnor U13731 (N_13731,N_12969,N_12735);
nor U13732 (N_13732,N_12850,N_12613);
nor U13733 (N_13733,N_12154,N_12919);
nand U13734 (N_13734,N_12013,N_12992);
xnor U13735 (N_13735,N_12533,N_12243);
xnor U13736 (N_13736,N_12810,N_12587);
xnor U13737 (N_13737,N_12330,N_12785);
or U13738 (N_13738,N_12400,N_12281);
or U13739 (N_13739,N_12018,N_12169);
xnor U13740 (N_13740,N_12562,N_12292);
or U13741 (N_13741,N_12194,N_12541);
or U13742 (N_13742,N_12790,N_12205);
nand U13743 (N_13743,N_12768,N_12753);
nor U13744 (N_13744,N_12183,N_12372);
or U13745 (N_13745,N_12583,N_12029);
or U13746 (N_13746,N_12702,N_12958);
or U13747 (N_13747,N_12915,N_12739);
nand U13748 (N_13748,N_12532,N_12153);
and U13749 (N_13749,N_12741,N_12883);
or U13750 (N_13750,N_12223,N_12800);
or U13751 (N_13751,N_12419,N_12990);
and U13752 (N_13752,N_12223,N_12472);
xor U13753 (N_13753,N_12194,N_12297);
and U13754 (N_13754,N_12540,N_12357);
xor U13755 (N_13755,N_12495,N_12976);
xnor U13756 (N_13756,N_12430,N_12285);
and U13757 (N_13757,N_12410,N_12923);
nand U13758 (N_13758,N_12212,N_12555);
or U13759 (N_13759,N_12841,N_12510);
xor U13760 (N_13760,N_12122,N_12662);
nand U13761 (N_13761,N_12628,N_12440);
and U13762 (N_13762,N_12607,N_12642);
and U13763 (N_13763,N_12468,N_12312);
and U13764 (N_13764,N_12317,N_12291);
or U13765 (N_13765,N_12044,N_12656);
or U13766 (N_13766,N_12388,N_12462);
xnor U13767 (N_13767,N_12670,N_12165);
xnor U13768 (N_13768,N_12131,N_12875);
and U13769 (N_13769,N_12506,N_12818);
nor U13770 (N_13770,N_12037,N_12429);
nand U13771 (N_13771,N_12608,N_12582);
nor U13772 (N_13772,N_12439,N_12431);
nand U13773 (N_13773,N_12677,N_12116);
xor U13774 (N_13774,N_12313,N_12067);
or U13775 (N_13775,N_12115,N_12551);
or U13776 (N_13776,N_12972,N_12628);
xor U13777 (N_13777,N_12288,N_12575);
and U13778 (N_13778,N_12869,N_12522);
or U13779 (N_13779,N_12148,N_12479);
nand U13780 (N_13780,N_12871,N_12195);
or U13781 (N_13781,N_12877,N_12047);
nor U13782 (N_13782,N_12491,N_12721);
nor U13783 (N_13783,N_12242,N_12578);
nand U13784 (N_13784,N_12465,N_12009);
nor U13785 (N_13785,N_12437,N_12113);
or U13786 (N_13786,N_12858,N_12497);
nor U13787 (N_13787,N_12638,N_12077);
xnor U13788 (N_13788,N_12131,N_12953);
nand U13789 (N_13789,N_12012,N_12371);
nor U13790 (N_13790,N_12953,N_12959);
and U13791 (N_13791,N_12749,N_12277);
and U13792 (N_13792,N_12466,N_12158);
nand U13793 (N_13793,N_12493,N_12934);
and U13794 (N_13794,N_12193,N_12741);
xnor U13795 (N_13795,N_12933,N_12402);
xnor U13796 (N_13796,N_12325,N_12599);
or U13797 (N_13797,N_12096,N_12186);
nor U13798 (N_13798,N_12392,N_12954);
or U13799 (N_13799,N_12081,N_12819);
and U13800 (N_13800,N_12678,N_12045);
nor U13801 (N_13801,N_12601,N_12534);
or U13802 (N_13802,N_12322,N_12753);
xor U13803 (N_13803,N_12282,N_12768);
xnor U13804 (N_13804,N_12898,N_12283);
xor U13805 (N_13805,N_12998,N_12791);
and U13806 (N_13806,N_12627,N_12239);
nand U13807 (N_13807,N_12842,N_12274);
xor U13808 (N_13808,N_12194,N_12391);
xnor U13809 (N_13809,N_12012,N_12320);
nor U13810 (N_13810,N_12378,N_12333);
and U13811 (N_13811,N_12098,N_12237);
or U13812 (N_13812,N_12414,N_12604);
nand U13813 (N_13813,N_12657,N_12622);
or U13814 (N_13814,N_12612,N_12389);
or U13815 (N_13815,N_12058,N_12226);
or U13816 (N_13816,N_12197,N_12834);
and U13817 (N_13817,N_12870,N_12490);
and U13818 (N_13818,N_12612,N_12282);
nor U13819 (N_13819,N_12735,N_12573);
nand U13820 (N_13820,N_12027,N_12512);
xor U13821 (N_13821,N_12550,N_12756);
and U13822 (N_13822,N_12621,N_12550);
and U13823 (N_13823,N_12912,N_12207);
or U13824 (N_13824,N_12800,N_12966);
and U13825 (N_13825,N_12613,N_12493);
nand U13826 (N_13826,N_12665,N_12182);
xor U13827 (N_13827,N_12755,N_12192);
and U13828 (N_13828,N_12773,N_12491);
nand U13829 (N_13829,N_12312,N_12943);
or U13830 (N_13830,N_12065,N_12467);
nor U13831 (N_13831,N_12574,N_12318);
nand U13832 (N_13832,N_12392,N_12345);
nor U13833 (N_13833,N_12281,N_12290);
nand U13834 (N_13834,N_12039,N_12279);
or U13835 (N_13835,N_12773,N_12684);
and U13836 (N_13836,N_12583,N_12737);
nor U13837 (N_13837,N_12969,N_12197);
nand U13838 (N_13838,N_12519,N_12818);
or U13839 (N_13839,N_12397,N_12118);
or U13840 (N_13840,N_12442,N_12670);
or U13841 (N_13841,N_12946,N_12397);
and U13842 (N_13842,N_12538,N_12606);
and U13843 (N_13843,N_12691,N_12643);
nand U13844 (N_13844,N_12907,N_12106);
or U13845 (N_13845,N_12419,N_12836);
and U13846 (N_13846,N_12773,N_12751);
nand U13847 (N_13847,N_12894,N_12254);
nor U13848 (N_13848,N_12855,N_12959);
xor U13849 (N_13849,N_12591,N_12660);
xnor U13850 (N_13850,N_12235,N_12992);
and U13851 (N_13851,N_12949,N_12174);
nor U13852 (N_13852,N_12967,N_12037);
xnor U13853 (N_13853,N_12210,N_12743);
or U13854 (N_13854,N_12663,N_12086);
nand U13855 (N_13855,N_12009,N_12282);
or U13856 (N_13856,N_12913,N_12250);
and U13857 (N_13857,N_12269,N_12316);
and U13858 (N_13858,N_12360,N_12342);
xnor U13859 (N_13859,N_12348,N_12135);
nand U13860 (N_13860,N_12238,N_12590);
xor U13861 (N_13861,N_12216,N_12491);
and U13862 (N_13862,N_12935,N_12734);
nor U13863 (N_13863,N_12285,N_12210);
or U13864 (N_13864,N_12018,N_12676);
or U13865 (N_13865,N_12958,N_12763);
xnor U13866 (N_13866,N_12098,N_12666);
or U13867 (N_13867,N_12776,N_12448);
and U13868 (N_13868,N_12478,N_12541);
or U13869 (N_13869,N_12111,N_12746);
nor U13870 (N_13870,N_12628,N_12172);
or U13871 (N_13871,N_12612,N_12531);
and U13872 (N_13872,N_12737,N_12740);
nand U13873 (N_13873,N_12009,N_12379);
nor U13874 (N_13874,N_12857,N_12883);
or U13875 (N_13875,N_12151,N_12190);
xor U13876 (N_13876,N_12488,N_12909);
nor U13877 (N_13877,N_12846,N_12662);
nand U13878 (N_13878,N_12041,N_12441);
and U13879 (N_13879,N_12760,N_12930);
xnor U13880 (N_13880,N_12576,N_12682);
and U13881 (N_13881,N_12347,N_12786);
nand U13882 (N_13882,N_12138,N_12603);
xor U13883 (N_13883,N_12760,N_12681);
or U13884 (N_13884,N_12604,N_12627);
and U13885 (N_13885,N_12297,N_12233);
nor U13886 (N_13886,N_12941,N_12035);
nor U13887 (N_13887,N_12478,N_12586);
or U13888 (N_13888,N_12244,N_12170);
and U13889 (N_13889,N_12612,N_12962);
xor U13890 (N_13890,N_12218,N_12781);
and U13891 (N_13891,N_12324,N_12887);
nor U13892 (N_13892,N_12396,N_12887);
and U13893 (N_13893,N_12563,N_12256);
and U13894 (N_13894,N_12019,N_12807);
nor U13895 (N_13895,N_12132,N_12703);
nand U13896 (N_13896,N_12697,N_12355);
nor U13897 (N_13897,N_12658,N_12985);
xnor U13898 (N_13898,N_12789,N_12240);
xor U13899 (N_13899,N_12783,N_12760);
xnor U13900 (N_13900,N_12789,N_12084);
xor U13901 (N_13901,N_12934,N_12454);
nor U13902 (N_13902,N_12573,N_12889);
nor U13903 (N_13903,N_12458,N_12917);
nand U13904 (N_13904,N_12738,N_12814);
and U13905 (N_13905,N_12263,N_12053);
nand U13906 (N_13906,N_12293,N_12584);
nand U13907 (N_13907,N_12663,N_12069);
and U13908 (N_13908,N_12313,N_12495);
nor U13909 (N_13909,N_12719,N_12163);
or U13910 (N_13910,N_12340,N_12330);
or U13911 (N_13911,N_12365,N_12027);
nand U13912 (N_13912,N_12387,N_12382);
nand U13913 (N_13913,N_12712,N_12210);
xor U13914 (N_13914,N_12367,N_12725);
xor U13915 (N_13915,N_12103,N_12179);
nand U13916 (N_13916,N_12485,N_12309);
xor U13917 (N_13917,N_12308,N_12202);
nand U13918 (N_13918,N_12832,N_12725);
or U13919 (N_13919,N_12028,N_12201);
nor U13920 (N_13920,N_12356,N_12498);
xnor U13921 (N_13921,N_12233,N_12580);
nor U13922 (N_13922,N_12457,N_12194);
xor U13923 (N_13923,N_12486,N_12975);
nor U13924 (N_13924,N_12246,N_12151);
or U13925 (N_13925,N_12974,N_12881);
nand U13926 (N_13926,N_12115,N_12735);
nor U13927 (N_13927,N_12150,N_12859);
and U13928 (N_13928,N_12757,N_12839);
and U13929 (N_13929,N_12825,N_12991);
nor U13930 (N_13930,N_12212,N_12526);
xnor U13931 (N_13931,N_12496,N_12157);
and U13932 (N_13932,N_12648,N_12004);
nand U13933 (N_13933,N_12866,N_12761);
or U13934 (N_13934,N_12030,N_12559);
nor U13935 (N_13935,N_12376,N_12467);
nor U13936 (N_13936,N_12941,N_12624);
xor U13937 (N_13937,N_12712,N_12774);
or U13938 (N_13938,N_12014,N_12801);
and U13939 (N_13939,N_12460,N_12154);
xor U13940 (N_13940,N_12841,N_12360);
xnor U13941 (N_13941,N_12356,N_12770);
and U13942 (N_13942,N_12296,N_12334);
or U13943 (N_13943,N_12795,N_12839);
and U13944 (N_13944,N_12562,N_12552);
nand U13945 (N_13945,N_12065,N_12787);
and U13946 (N_13946,N_12867,N_12437);
and U13947 (N_13947,N_12177,N_12071);
xor U13948 (N_13948,N_12741,N_12087);
and U13949 (N_13949,N_12450,N_12276);
and U13950 (N_13950,N_12430,N_12878);
nand U13951 (N_13951,N_12249,N_12256);
nor U13952 (N_13952,N_12532,N_12900);
nor U13953 (N_13953,N_12704,N_12102);
nor U13954 (N_13954,N_12821,N_12708);
xor U13955 (N_13955,N_12046,N_12564);
nor U13956 (N_13956,N_12837,N_12080);
or U13957 (N_13957,N_12838,N_12723);
nor U13958 (N_13958,N_12984,N_12674);
or U13959 (N_13959,N_12459,N_12002);
xor U13960 (N_13960,N_12971,N_12595);
xor U13961 (N_13961,N_12035,N_12184);
and U13962 (N_13962,N_12472,N_12395);
nand U13963 (N_13963,N_12503,N_12365);
nand U13964 (N_13964,N_12716,N_12132);
xnor U13965 (N_13965,N_12008,N_12577);
xnor U13966 (N_13966,N_12195,N_12295);
or U13967 (N_13967,N_12477,N_12865);
nand U13968 (N_13968,N_12624,N_12548);
nor U13969 (N_13969,N_12385,N_12937);
xnor U13970 (N_13970,N_12236,N_12631);
xnor U13971 (N_13971,N_12568,N_12818);
and U13972 (N_13972,N_12898,N_12873);
or U13973 (N_13973,N_12491,N_12245);
nor U13974 (N_13974,N_12629,N_12048);
xor U13975 (N_13975,N_12664,N_12075);
nor U13976 (N_13976,N_12407,N_12305);
and U13977 (N_13977,N_12203,N_12486);
nand U13978 (N_13978,N_12761,N_12854);
nor U13979 (N_13979,N_12807,N_12733);
nor U13980 (N_13980,N_12460,N_12080);
xnor U13981 (N_13981,N_12546,N_12396);
xor U13982 (N_13982,N_12686,N_12003);
or U13983 (N_13983,N_12543,N_12553);
nand U13984 (N_13984,N_12683,N_12744);
and U13985 (N_13985,N_12681,N_12534);
nand U13986 (N_13986,N_12473,N_12540);
xor U13987 (N_13987,N_12391,N_12912);
xor U13988 (N_13988,N_12458,N_12496);
nand U13989 (N_13989,N_12612,N_12537);
and U13990 (N_13990,N_12609,N_12626);
and U13991 (N_13991,N_12052,N_12272);
nand U13992 (N_13992,N_12979,N_12385);
xnor U13993 (N_13993,N_12660,N_12407);
xnor U13994 (N_13994,N_12552,N_12490);
xnor U13995 (N_13995,N_12756,N_12010);
xnor U13996 (N_13996,N_12477,N_12316);
nor U13997 (N_13997,N_12443,N_12029);
xor U13998 (N_13998,N_12337,N_12550);
or U13999 (N_13999,N_12167,N_12096);
or U14000 (N_14000,N_13910,N_13527);
xnor U14001 (N_14001,N_13508,N_13178);
or U14002 (N_14002,N_13501,N_13451);
nand U14003 (N_14003,N_13430,N_13194);
and U14004 (N_14004,N_13116,N_13391);
xor U14005 (N_14005,N_13084,N_13512);
xor U14006 (N_14006,N_13760,N_13039);
xnor U14007 (N_14007,N_13573,N_13268);
nand U14008 (N_14008,N_13970,N_13074);
nand U14009 (N_14009,N_13955,N_13563);
xnor U14010 (N_14010,N_13727,N_13920);
xor U14011 (N_14011,N_13153,N_13419);
xnor U14012 (N_14012,N_13219,N_13759);
nand U14013 (N_14013,N_13120,N_13250);
nand U14014 (N_14014,N_13701,N_13063);
and U14015 (N_14015,N_13246,N_13318);
nand U14016 (N_14016,N_13119,N_13911);
nand U14017 (N_14017,N_13572,N_13005);
nor U14018 (N_14018,N_13413,N_13693);
xor U14019 (N_14019,N_13638,N_13981);
or U14020 (N_14020,N_13748,N_13598);
xor U14021 (N_14021,N_13353,N_13372);
nand U14022 (N_14022,N_13043,N_13105);
and U14023 (N_14023,N_13912,N_13800);
and U14024 (N_14024,N_13624,N_13183);
nor U14025 (N_14025,N_13238,N_13146);
xnor U14026 (N_14026,N_13409,N_13228);
nand U14027 (N_14027,N_13042,N_13832);
xnor U14028 (N_14028,N_13266,N_13869);
nor U14029 (N_14029,N_13552,N_13035);
nand U14030 (N_14030,N_13079,N_13725);
nor U14031 (N_14031,N_13616,N_13252);
nand U14032 (N_14032,N_13464,N_13886);
or U14033 (N_14033,N_13987,N_13967);
nand U14034 (N_14034,N_13744,N_13431);
nand U14035 (N_14035,N_13921,N_13668);
nand U14036 (N_14036,N_13386,N_13775);
nand U14037 (N_14037,N_13139,N_13015);
nand U14038 (N_14038,N_13352,N_13368);
nor U14039 (N_14039,N_13485,N_13135);
and U14040 (N_14040,N_13847,N_13164);
or U14041 (N_14041,N_13296,N_13033);
nor U14042 (N_14042,N_13816,N_13576);
nor U14043 (N_14043,N_13992,N_13198);
and U14044 (N_14044,N_13018,N_13048);
or U14045 (N_14045,N_13160,N_13503);
and U14046 (N_14046,N_13067,N_13533);
and U14047 (N_14047,N_13637,N_13754);
xnor U14048 (N_14048,N_13136,N_13762);
nand U14049 (N_14049,N_13627,N_13123);
xnor U14050 (N_14050,N_13118,N_13375);
nor U14051 (N_14051,N_13176,N_13940);
nor U14052 (N_14052,N_13764,N_13271);
xor U14053 (N_14053,N_13507,N_13931);
and U14054 (N_14054,N_13144,N_13787);
nor U14055 (N_14055,N_13009,N_13289);
or U14056 (N_14056,N_13639,N_13003);
and U14057 (N_14057,N_13640,N_13203);
nand U14058 (N_14058,N_13614,N_13393);
or U14059 (N_14059,N_13729,N_13661);
or U14060 (N_14060,N_13620,N_13613);
and U14061 (N_14061,N_13215,N_13845);
and U14062 (N_14062,N_13114,N_13104);
or U14063 (N_14063,N_13685,N_13364);
xnor U14064 (N_14064,N_13423,N_13954);
nor U14065 (N_14065,N_13878,N_13898);
or U14066 (N_14066,N_13418,N_13773);
or U14067 (N_14067,N_13389,N_13392);
xor U14068 (N_14068,N_13076,N_13989);
nand U14069 (N_14069,N_13736,N_13702);
nor U14070 (N_14070,N_13703,N_13936);
or U14071 (N_14071,N_13166,N_13276);
nor U14072 (N_14072,N_13578,N_13601);
xnor U14073 (N_14073,N_13195,N_13712);
nor U14074 (N_14074,N_13677,N_13997);
and U14075 (N_14075,N_13542,N_13926);
xnor U14076 (N_14076,N_13836,N_13486);
and U14077 (N_14077,N_13458,N_13723);
xnor U14078 (N_14078,N_13843,N_13522);
or U14079 (N_14079,N_13355,N_13444);
xor U14080 (N_14080,N_13167,N_13185);
and U14081 (N_14081,N_13567,N_13377);
and U14082 (N_14082,N_13795,N_13647);
xor U14083 (N_14083,N_13779,N_13579);
nand U14084 (N_14084,N_13628,N_13047);
or U14085 (N_14085,N_13087,N_13498);
xnor U14086 (N_14086,N_13959,N_13256);
nor U14087 (N_14087,N_13900,N_13496);
nand U14088 (N_14088,N_13312,N_13150);
nor U14089 (N_14089,N_13516,N_13095);
xnor U14090 (N_14090,N_13864,N_13839);
nor U14091 (N_14091,N_13283,N_13259);
nand U14092 (N_14092,N_13958,N_13983);
xnor U14093 (N_14093,N_13093,N_13460);
or U14094 (N_14094,N_13667,N_13680);
nor U14095 (N_14095,N_13991,N_13143);
nand U14096 (N_14096,N_13265,N_13478);
xor U14097 (N_14097,N_13088,N_13811);
or U14098 (N_14098,N_13604,N_13100);
nor U14099 (N_14099,N_13326,N_13124);
and U14100 (N_14100,N_13761,N_13913);
nand U14101 (N_14101,N_13121,N_13255);
xor U14102 (N_14102,N_13092,N_13536);
or U14103 (N_14103,N_13110,N_13867);
nand U14104 (N_14104,N_13013,N_13710);
nor U14105 (N_14105,N_13949,N_13891);
and U14106 (N_14106,N_13626,N_13681);
nand U14107 (N_14107,N_13101,N_13887);
nand U14108 (N_14108,N_13052,N_13127);
or U14109 (N_14109,N_13551,N_13417);
or U14110 (N_14110,N_13996,N_13490);
and U14111 (N_14111,N_13059,N_13062);
nor U14112 (N_14112,N_13367,N_13530);
xnor U14113 (N_14113,N_13137,N_13995);
xnor U14114 (N_14114,N_13466,N_13607);
nand U14115 (N_14115,N_13874,N_13592);
or U14116 (N_14116,N_13260,N_13141);
nor U14117 (N_14117,N_13528,N_13525);
nor U14118 (N_14118,N_13644,N_13243);
nor U14119 (N_14119,N_13611,N_13347);
or U14120 (N_14120,N_13140,N_13286);
and U14121 (N_14121,N_13863,N_13837);
or U14122 (N_14122,N_13481,N_13814);
nand U14123 (N_14123,N_13133,N_13986);
nor U14124 (N_14124,N_13502,N_13189);
xor U14125 (N_14125,N_13310,N_13763);
or U14126 (N_14126,N_13969,N_13558);
nand U14127 (N_14127,N_13044,N_13051);
or U14128 (N_14128,N_13196,N_13232);
nor U14129 (N_14129,N_13830,N_13817);
or U14130 (N_14130,N_13077,N_13623);
nor U14131 (N_14131,N_13977,N_13138);
and U14132 (N_14132,N_13309,N_13669);
nor U14133 (N_14133,N_13828,N_13365);
xor U14134 (N_14134,N_13511,N_13709);
nand U14135 (N_14135,N_13161,N_13155);
and U14136 (N_14136,N_13295,N_13565);
and U14137 (N_14137,N_13350,N_13621);
or U14138 (N_14138,N_13274,N_13381);
or U14139 (N_14139,N_13450,N_13899);
xor U14140 (N_14140,N_13071,N_13069);
nor U14141 (N_14141,N_13017,N_13468);
or U14142 (N_14142,N_13738,N_13348);
nor U14143 (N_14143,N_13467,N_13461);
nor U14144 (N_14144,N_13299,N_13169);
or U14145 (N_14145,N_13794,N_13534);
xor U14146 (N_14146,N_13943,N_13732);
xnor U14147 (N_14147,N_13242,N_13745);
or U14148 (N_14148,N_13798,N_13019);
nor U14149 (N_14149,N_13718,N_13157);
nand U14150 (N_14150,N_13251,N_13390);
or U14151 (N_14151,N_13765,N_13889);
nand U14152 (N_14152,N_13494,N_13739);
nor U14153 (N_14153,N_13756,N_13480);
nand U14154 (N_14154,N_13923,N_13788);
nor U14155 (N_14155,N_13865,N_13394);
and U14156 (N_14156,N_13369,N_13148);
or U14157 (N_14157,N_13323,N_13441);
and U14158 (N_14158,N_13434,N_13181);
nor U14159 (N_14159,N_13649,N_13154);
nand U14160 (N_14160,N_13520,N_13491);
xnor U14161 (N_14161,N_13320,N_13014);
nand U14162 (N_14162,N_13514,N_13708);
or U14163 (N_14163,N_13191,N_13281);
nand U14164 (N_14164,N_13403,N_13646);
nand U14165 (N_14165,N_13683,N_13332);
or U14166 (N_14166,N_13257,N_13747);
nand U14167 (N_14167,N_13550,N_13346);
nor U14168 (N_14168,N_13999,N_13218);
or U14169 (N_14169,N_13933,N_13134);
nand U14170 (N_14170,N_13605,N_13792);
nand U14171 (N_14171,N_13325,N_13882);
nand U14172 (N_14172,N_13472,N_13408);
xor U14173 (N_14173,N_13860,N_13094);
nor U14174 (N_14174,N_13329,N_13262);
nor U14175 (N_14175,N_13666,N_13894);
nor U14176 (N_14176,N_13509,N_13938);
xor U14177 (N_14177,N_13045,N_13258);
xnor U14178 (N_14178,N_13953,N_13674);
and U14179 (N_14179,N_13713,N_13755);
nor U14180 (N_14180,N_13208,N_13657);
nor U14181 (N_14181,N_13635,N_13929);
or U14182 (N_14182,N_13826,N_13179);
nor U14183 (N_14183,N_13149,N_13361);
and U14184 (N_14184,N_13803,N_13791);
xor U14185 (N_14185,N_13342,N_13223);
nor U14186 (N_14186,N_13777,N_13385);
nand U14187 (N_14187,N_13532,N_13396);
nand U14188 (N_14188,N_13807,N_13584);
nand U14189 (N_14189,N_13948,N_13696);
xnor U14190 (N_14190,N_13632,N_13589);
and U14191 (N_14191,N_13880,N_13964);
xor U14192 (N_14192,N_13724,N_13619);
or U14193 (N_14193,N_13307,N_13993);
nor U14194 (N_14194,N_13022,N_13446);
nor U14195 (N_14195,N_13881,N_13500);
nand U14196 (N_14196,N_13021,N_13927);
nor U14197 (N_14197,N_13041,N_13694);
nor U14198 (N_14198,N_13590,N_13147);
nand U14199 (N_14199,N_13050,N_13965);
and U14200 (N_14200,N_13870,N_13379);
nand U14201 (N_14201,N_13304,N_13278);
or U14202 (N_14202,N_13539,N_13400);
nor U14203 (N_14203,N_13631,N_13495);
and U14204 (N_14204,N_13730,N_13952);
nor U14205 (N_14205,N_13156,N_13142);
xor U14206 (N_14206,N_13175,N_13410);
nand U14207 (N_14207,N_13239,N_13673);
and U14208 (N_14208,N_13227,N_13893);
nor U14209 (N_14209,N_13414,N_13914);
xnor U14210 (N_14210,N_13825,N_13126);
nor U14211 (N_14211,N_13554,N_13388);
xnor U14212 (N_14212,N_13335,N_13838);
or U14213 (N_14213,N_13324,N_13688);
xor U14214 (N_14214,N_13222,N_13433);
xnor U14215 (N_14215,N_13924,N_13122);
and U14216 (N_14216,N_13820,N_13850);
or U14217 (N_14217,N_13518,N_13772);
nor U14218 (N_14218,N_13474,N_13753);
or U14219 (N_14219,N_13109,N_13813);
xor U14220 (N_14220,N_13333,N_13054);
xnor U14221 (N_14221,N_13848,N_13658);
and U14222 (N_14222,N_13767,N_13602);
and U14223 (N_14223,N_13363,N_13700);
nand U14224 (N_14224,N_13231,N_13892);
xor U14225 (N_14225,N_13793,N_13538);
nor U14226 (N_14226,N_13244,N_13210);
nor U14227 (N_14227,N_13734,N_13782);
nand U14228 (N_14228,N_13334,N_13315);
xor U14229 (N_14229,N_13901,N_13275);
nand U14230 (N_14230,N_13654,N_13254);
xnor U14231 (N_14231,N_13004,N_13586);
or U14232 (N_14232,N_13883,N_13078);
nor U14233 (N_14233,N_13086,N_13676);
nor U14234 (N_14234,N_13188,N_13888);
and U14235 (N_14235,N_13984,N_13636);
and U14236 (N_14236,N_13769,N_13523);
or U14237 (N_14237,N_13543,N_13566);
xnor U14238 (N_14238,N_13766,N_13002);
xor U14239 (N_14239,N_13440,N_13719);
nand U14240 (N_14240,N_13085,N_13497);
nor U14241 (N_14241,N_13297,N_13159);
nor U14242 (N_14242,N_13402,N_13200);
nand U14243 (N_14243,N_13944,N_13302);
and U14244 (N_14244,N_13192,N_13588);
nor U14245 (N_14245,N_13505,N_13822);
nor U14246 (N_14246,N_13107,N_13854);
xor U14247 (N_14247,N_13337,N_13934);
or U14248 (N_14248,N_13399,N_13199);
xor U14249 (N_14249,N_13055,N_13540);
nand U14250 (N_14250,N_13061,N_13305);
or U14251 (N_14251,N_13974,N_13233);
xor U14252 (N_14252,N_13277,N_13449);
nand U14253 (N_14253,N_13561,N_13416);
or U14254 (N_14254,N_13629,N_13317);
and U14255 (N_14255,N_13207,N_13331);
or U14256 (N_14256,N_13343,N_13455);
nand U14257 (N_14257,N_13922,N_13341);
nor U14258 (N_14258,N_13224,N_13438);
xnor U14259 (N_14259,N_13270,N_13098);
and U14260 (N_14260,N_13130,N_13282);
nand U14261 (N_14261,N_13932,N_13306);
and U14262 (N_14262,N_13383,N_13090);
xnor U14263 (N_14263,N_13594,N_13966);
and U14264 (N_14264,N_13939,N_13956);
and U14265 (N_14265,N_13930,N_13855);
nor U14266 (N_14266,N_13960,N_13612);
xnor U14267 (N_14267,N_13735,N_13526);
or U14268 (N_14268,N_13452,N_13571);
nor U14269 (N_14269,N_13454,N_13065);
xor U14270 (N_14270,N_13663,N_13432);
xor U14271 (N_14271,N_13327,N_13988);
nor U14272 (N_14272,N_13961,N_13597);
or U14273 (N_14273,N_13174,N_13687);
and U14274 (N_14274,N_13699,N_13670);
nor U14275 (N_14275,N_13979,N_13583);
xnor U14276 (N_14276,N_13235,N_13345);
or U14277 (N_14277,N_13475,N_13802);
xor U14278 (N_14278,N_13796,N_13294);
and U14279 (N_14279,N_13717,N_13273);
and U14280 (N_14280,N_13715,N_13338);
nand U14281 (N_14281,N_13875,N_13284);
or U14282 (N_14282,N_13113,N_13513);
xnor U14283 (N_14283,N_13751,N_13264);
xnor U14284 (N_14284,N_13316,N_13405);
xnor U14285 (N_14285,N_13942,N_13716);
nand U14286 (N_14286,N_13840,N_13902);
and U14287 (N_14287,N_13737,N_13556);
and U14288 (N_14288,N_13547,N_13099);
and U14289 (N_14289,N_13908,N_13706);
xor U14290 (N_14290,N_13746,N_13951);
or U14291 (N_14291,N_13027,N_13907);
nor U14292 (N_14292,N_13267,N_13428);
nor U14293 (N_14293,N_13682,N_13241);
and U14294 (N_14294,N_13036,N_13553);
xor U14295 (N_14295,N_13941,N_13422);
or U14296 (N_14296,N_13871,N_13544);
and U14297 (N_14297,N_13280,N_13557);
nand U14298 (N_14298,N_13487,N_13378);
nor U14299 (N_14299,N_13660,N_13492);
and U14300 (N_14300,N_13453,N_13785);
and U14301 (N_14301,N_13443,N_13128);
or U14302 (N_14302,N_13030,N_13978);
and U14303 (N_14303,N_13226,N_13023);
xnor U14304 (N_14304,N_13844,N_13517);
nand U14305 (N_14305,N_13132,N_13585);
or U14306 (N_14306,N_13288,N_13925);
nand U14307 (N_14307,N_13852,N_13291);
xnor U14308 (N_14308,N_13555,N_13293);
nor U14309 (N_14309,N_13482,N_13469);
nor U14310 (N_14310,N_13398,N_13415);
and U14311 (N_14311,N_13784,N_13873);
xor U14312 (N_14312,N_13645,N_13476);
nor U14313 (N_14313,N_13531,N_13285);
and U14314 (N_14314,N_13722,N_13070);
nor U14315 (N_14315,N_13499,N_13998);
or U14316 (N_14316,N_13362,N_13108);
and U14317 (N_14317,N_13945,N_13648);
and U14318 (N_14318,N_13906,N_13008);
nor U14319 (N_14319,N_13780,N_13537);
or U14320 (N_14320,N_13720,N_13568);
nor U14321 (N_14321,N_13439,N_13075);
nor U14322 (N_14322,N_13985,N_13245);
nor U14323 (N_14323,N_13359,N_13221);
nand U14324 (N_14324,N_13225,N_13456);
nor U14325 (N_14325,N_13115,N_13479);
and U14326 (N_14326,N_13812,N_13424);
xnor U14327 (N_14327,N_13397,N_13382);
xor U14328 (N_14328,N_13229,N_13664);
nand U14329 (N_14329,N_13918,N_13704);
xnor U14330 (N_14330,N_13833,N_13690);
xnor U14331 (N_14331,N_13506,N_13301);
and U14332 (N_14332,N_13373,N_13808);
nand U14333 (N_14333,N_13020,N_13356);
or U14334 (N_14334,N_13170,N_13809);
and U14335 (N_14335,N_13609,N_13308);
nor U14336 (N_14336,N_13937,N_13615);
nand U14337 (N_14337,N_13319,N_13994);
or U14338 (N_14338,N_13376,N_13504);
xor U14339 (N_14339,N_13484,N_13919);
or U14340 (N_14340,N_13692,N_13560);
and U14341 (N_14341,N_13064,N_13240);
or U14342 (N_14342,N_13786,N_13928);
nand U14343 (N_14343,N_13213,N_13351);
nand U14344 (N_14344,N_13728,N_13824);
xor U14345 (N_14345,N_13016,N_13314);
xor U14346 (N_14346,N_13072,N_13651);
or U14347 (N_14347,N_13292,N_13968);
nor U14348 (N_14348,N_13608,N_13354);
nand U14349 (N_14349,N_13053,N_13510);
xnor U14350 (N_14350,N_13884,N_13435);
and U14351 (N_14351,N_13581,N_13757);
and U14352 (N_14352,N_13407,N_13829);
xnor U14353 (N_14353,N_13957,N_13618);
or U14354 (N_14354,N_13106,N_13726);
nand U14355 (N_14355,N_13743,N_13470);
xnor U14356 (N_14356,N_13797,N_13007);
and U14357 (N_14357,N_13406,N_13591);
nand U14358 (N_14358,N_13695,N_13742);
nand U14359 (N_14359,N_13653,N_13524);
or U14360 (N_14360,N_13990,N_13436);
and U14361 (N_14361,N_13321,N_13298);
xor U14362 (N_14362,N_13789,N_13896);
or U14363 (N_14363,N_13112,N_13425);
xnor U14364 (N_14364,N_13749,N_13272);
or U14365 (N_14365,N_13129,N_13603);
or U14366 (N_14366,N_13483,N_13574);
nand U14367 (N_14367,N_13905,N_13916);
and U14368 (N_14368,N_13214,N_13721);
or U14369 (N_14369,N_13360,N_13165);
xor U14370 (N_14370,N_13197,N_13890);
and U14371 (N_14371,N_13493,N_13903);
nand U14372 (N_14372,N_13209,N_13339);
or U14373 (N_14373,N_13125,N_13862);
nand U14374 (N_14374,N_13287,N_13650);
nor U14375 (N_14375,N_13655,N_13783);
nor U14376 (N_14376,N_13263,N_13853);
nor U14377 (N_14377,N_13387,N_13401);
and U14378 (N_14378,N_13366,N_13740);
xor U14379 (N_14379,N_13117,N_13404);
nor U14380 (N_14380,N_13752,N_13322);
nand U14381 (N_14381,N_13473,N_13025);
or U14382 (N_14382,N_13290,N_13672);
nand U14383 (N_14383,N_13678,N_13935);
nand U14384 (N_14384,N_13575,N_13230);
and U14385 (N_14385,N_13212,N_13714);
xnor U14386 (N_14386,N_13617,N_13488);
or U14387 (N_14387,N_13577,N_13193);
and U14388 (N_14388,N_13380,N_13823);
xor U14389 (N_14389,N_13340,N_13841);
nand U14390 (N_14390,N_13336,N_13068);
or U14391 (N_14391,N_13012,N_13859);
and U14392 (N_14392,N_13972,N_13201);
nor U14393 (N_14393,N_13031,N_13976);
xor U14394 (N_14394,N_13963,N_13037);
xor U14395 (N_14395,N_13058,N_13546);
nor U14396 (N_14396,N_13758,N_13630);
nor U14397 (N_14397,N_13834,N_13060);
xnor U14398 (N_14398,N_13187,N_13384);
xor U14399 (N_14399,N_13519,N_13876);
or U14400 (N_14400,N_13562,N_13778);
nor U14401 (N_14401,N_13622,N_13858);
xnor U14402 (N_14402,N_13006,N_13868);
nor U14403 (N_14403,N_13580,N_13950);
or U14404 (N_14404,N_13371,N_13489);
nand U14405 (N_14405,N_13034,N_13818);
nand U14406 (N_14406,N_13349,N_13973);
nand U14407 (N_14407,N_13249,N_13705);
or U14408 (N_14408,N_13915,N_13559);
and U14409 (N_14409,N_13711,N_13083);
xor U14410 (N_14410,N_13570,N_13781);
xor U14411 (N_14411,N_13776,N_13427);
and U14412 (N_14412,N_13172,N_13815);
xnor U14413 (N_14413,N_13861,N_13857);
nand U14414 (N_14414,N_13421,N_13202);
nor U14415 (N_14415,N_13011,N_13463);
nor U14416 (N_14416,N_13600,N_13529);
nor U14417 (N_14417,N_13145,N_13459);
xnor U14418 (N_14418,N_13593,N_13872);
nor U14419 (N_14419,N_13096,N_13545);
or U14420 (N_14420,N_13541,N_13131);
xnor U14421 (N_14421,N_13163,N_13049);
xnor U14422 (N_14422,N_13689,N_13186);
nor U14423 (N_14423,N_13885,N_13686);
and U14424 (N_14424,N_13253,N_13810);
nor U14425 (N_14425,N_13980,N_13827);
and U14426 (N_14426,N_13158,N_13733);
or U14427 (N_14427,N_13103,N_13102);
nand U14428 (N_14428,N_13633,N_13247);
or U14429 (N_14429,N_13057,N_13206);
and U14430 (N_14430,N_13205,N_13426);
nor U14431 (N_14431,N_13835,N_13741);
nand U14432 (N_14432,N_13162,N_13248);
nand U14433 (N_14433,N_13866,N_13947);
nand U14434 (N_14434,N_13080,N_13081);
nand U14435 (N_14435,N_13750,N_13173);
xnor U14436 (N_14436,N_13768,N_13831);
and U14437 (N_14437,N_13671,N_13731);
nor U14438 (N_14438,N_13975,N_13056);
nor U14439 (N_14439,N_13851,N_13445);
nor U14440 (N_14440,N_13066,N_13684);
and U14441 (N_14441,N_13790,N_13842);
xnor U14442 (N_14442,N_13024,N_13895);
xor U14443 (N_14443,N_13535,N_13625);
nand U14444 (N_14444,N_13182,N_13001);
xnor U14445 (N_14445,N_13799,N_13643);
or U14446 (N_14446,N_13448,N_13641);
or U14447 (N_14447,N_13089,N_13211);
xor U14448 (N_14448,N_13564,N_13521);
nor U14449 (N_14449,N_13656,N_13634);
or U14450 (N_14450,N_13804,N_13515);
xor U14451 (N_14451,N_13046,N_13819);
and U14452 (N_14452,N_13204,N_13269);
and U14453 (N_14453,N_13236,N_13040);
xnor U14454 (N_14454,N_13707,N_13599);
nor U14455 (N_14455,N_13462,N_13856);
nand U14456 (N_14456,N_13477,N_13190);
or U14457 (N_14457,N_13471,N_13442);
nand U14458 (N_14458,N_13982,N_13904);
xnor U14459 (N_14459,N_13805,N_13849);
nor U14460 (N_14460,N_13082,N_13659);
nor U14461 (N_14461,N_13595,N_13642);
or U14462 (N_14462,N_13457,N_13879);
nand U14463 (N_14463,N_13216,N_13217);
xnor U14464 (N_14464,N_13311,N_13357);
and U14465 (N_14465,N_13028,N_13697);
nor U14466 (N_14466,N_13909,N_13606);
nor U14467 (N_14467,N_13411,N_13429);
xnor U14468 (N_14468,N_13962,N_13610);
or U14469 (N_14469,N_13806,N_13877);
and U14470 (N_14470,N_13374,N_13770);
nor U14471 (N_14471,N_13897,N_13097);
xnor U14472 (N_14472,N_13177,N_13000);
nor U14473 (N_14473,N_13846,N_13358);
nor U14474 (N_14474,N_13237,N_13821);
and U14475 (N_14475,N_13261,N_13698);
or U14476 (N_14476,N_13029,N_13330);
and U14477 (N_14477,N_13582,N_13300);
xnor U14478 (N_14478,N_13091,N_13220);
or U14479 (N_14479,N_13395,N_13771);
and U14480 (N_14480,N_13548,N_13774);
and U14481 (N_14481,N_13010,N_13032);
xor U14482 (N_14482,N_13180,N_13437);
nand U14483 (N_14483,N_13152,N_13946);
or U14484 (N_14484,N_13344,N_13412);
or U14485 (N_14485,N_13313,N_13151);
nor U14486 (N_14486,N_13679,N_13328);
nor U14487 (N_14487,N_13234,N_13184);
nor U14488 (N_14488,N_13665,N_13691);
and U14489 (N_14489,N_13465,N_13587);
nand U14490 (N_14490,N_13420,N_13569);
nor U14491 (N_14491,N_13168,N_13662);
xor U14492 (N_14492,N_13171,N_13111);
and U14493 (N_14493,N_13596,N_13549);
or U14494 (N_14494,N_13303,N_13917);
or U14495 (N_14495,N_13026,N_13370);
and U14496 (N_14496,N_13279,N_13447);
xor U14497 (N_14497,N_13801,N_13652);
and U14498 (N_14498,N_13675,N_13971);
and U14499 (N_14499,N_13038,N_13073);
nor U14500 (N_14500,N_13067,N_13866);
nor U14501 (N_14501,N_13362,N_13554);
xnor U14502 (N_14502,N_13873,N_13488);
and U14503 (N_14503,N_13025,N_13073);
and U14504 (N_14504,N_13009,N_13374);
and U14505 (N_14505,N_13898,N_13162);
nor U14506 (N_14506,N_13814,N_13093);
or U14507 (N_14507,N_13391,N_13789);
or U14508 (N_14508,N_13824,N_13147);
or U14509 (N_14509,N_13105,N_13268);
xnor U14510 (N_14510,N_13513,N_13500);
and U14511 (N_14511,N_13831,N_13090);
xnor U14512 (N_14512,N_13169,N_13208);
xnor U14513 (N_14513,N_13880,N_13895);
and U14514 (N_14514,N_13624,N_13587);
xor U14515 (N_14515,N_13265,N_13030);
or U14516 (N_14516,N_13991,N_13884);
xnor U14517 (N_14517,N_13186,N_13347);
or U14518 (N_14518,N_13591,N_13252);
nor U14519 (N_14519,N_13104,N_13594);
xnor U14520 (N_14520,N_13814,N_13508);
and U14521 (N_14521,N_13817,N_13109);
or U14522 (N_14522,N_13344,N_13247);
and U14523 (N_14523,N_13914,N_13557);
nand U14524 (N_14524,N_13390,N_13258);
and U14525 (N_14525,N_13603,N_13373);
or U14526 (N_14526,N_13144,N_13611);
xor U14527 (N_14527,N_13040,N_13503);
nor U14528 (N_14528,N_13924,N_13612);
and U14529 (N_14529,N_13411,N_13932);
nand U14530 (N_14530,N_13797,N_13353);
and U14531 (N_14531,N_13543,N_13779);
or U14532 (N_14532,N_13430,N_13818);
xnor U14533 (N_14533,N_13100,N_13259);
nand U14534 (N_14534,N_13835,N_13356);
xnor U14535 (N_14535,N_13381,N_13974);
nand U14536 (N_14536,N_13577,N_13113);
or U14537 (N_14537,N_13184,N_13407);
and U14538 (N_14538,N_13640,N_13741);
nand U14539 (N_14539,N_13185,N_13192);
or U14540 (N_14540,N_13321,N_13734);
nor U14541 (N_14541,N_13911,N_13607);
or U14542 (N_14542,N_13170,N_13216);
nor U14543 (N_14543,N_13573,N_13087);
nand U14544 (N_14544,N_13787,N_13893);
xor U14545 (N_14545,N_13842,N_13924);
xor U14546 (N_14546,N_13304,N_13689);
nor U14547 (N_14547,N_13575,N_13189);
xnor U14548 (N_14548,N_13406,N_13801);
or U14549 (N_14549,N_13685,N_13292);
xnor U14550 (N_14550,N_13898,N_13487);
or U14551 (N_14551,N_13591,N_13014);
nor U14552 (N_14552,N_13196,N_13524);
nor U14553 (N_14553,N_13530,N_13548);
nand U14554 (N_14554,N_13799,N_13991);
nand U14555 (N_14555,N_13300,N_13868);
and U14556 (N_14556,N_13169,N_13064);
or U14557 (N_14557,N_13937,N_13347);
nor U14558 (N_14558,N_13023,N_13846);
or U14559 (N_14559,N_13657,N_13862);
nand U14560 (N_14560,N_13713,N_13207);
xor U14561 (N_14561,N_13008,N_13480);
nor U14562 (N_14562,N_13841,N_13216);
nor U14563 (N_14563,N_13628,N_13623);
nor U14564 (N_14564,N_13041,N_13351);
nand U14565 (N_14565,N_13264,N_13706);
nand U14566 (N_14566,N_13184,N_13294);
xor U14567 (N_14567,N_13787,N_13797);
or U14568 (N_14568,N_13107,N_13616);
nand U14569 (N_14569,N_13114,N_13153);
xnor U14570 (N_14570,N_13057,N_13317);
xor U14571 (N_14571,N_13062,N_13881);
or U14572 (N_14572,N_13764,N_13371);
or U14573 (N_14573,N_13650,N_13513);
nor U14574 (N_14574,N_13148,N_13594);
nor U14575 (N_14575,N_13823,N_13566);
nand U14576 (N_14576,N_13945,N_13092);
nor U14577 (N_14577,N_13619,N_13074);
nand U14578 (N_14578,N_13923,N_13762);
nand U14579 (N_14579,N_13994,N_13372);
xor U14580 (N_14580,N_13497,N_13340);
xnor U14581 (N_14581,N_13436,N_13964);
xor U14582 (N_14582,N_13224,N_13709);
nand U14583 (N_14583,N_13533,N_13757);
nand U14584 (N_14584,N_13819,N_13566);
xor U14585 (N_14585,N_13960,N_13463);
xor U14586 (N_14586,N_13862,N_13299);
or U14587 (N_14587,N_13113,N_13214);
and U14588 (N_14588,N_13437,N_13350);
and U14589 (N_14589,N_13297,N_13193);
and U14590 (N_14590,N_13786,N_13695);
nand U14591 (N_14591,N_13325,N_13466);
nand U14592 (N_14592,N_13026,N_13160);
or U14593 (N_14593,N_13226,N_13961);
nand U14594 (N_14594,N_13484,N_13540);
and U14595 (N_14595,N_13860,N_13421);
or U14596 (N_14596,N_13413,N_13698);
nor U14597 (N_14597,N_13125,N_13885);
nand U14598 (N_14598,N_13126,N_13321);
or U14599 (N_14599,N_13203,N_13369);
nand U14600 (N_14600,N_13490,N_13045);
or U14601 (N_14601,N_13643,N_13523);
nor U14602 (N_14602,N_13831,N_13243);
xnor U14603 (N_14603,N_13908,N_13880);
nand U14604 (N_14604,N_13277,N_13581);
or U14605 (N_14605,N_13113,N_13520);
xnor U14606 (N_14606,N_13609,N_13086);
xor U14607 (N_14607,N_13804,N_13823);
and U14608 (N_14608,N_13087,N_13443);
xor U14609 (N_14609,N_13908,N_13087);
or U14610 (N_14610,N_13404,N_13369);
xor U14611 (N_14611,N_13097,N_13533);
nand U14612 (N_14612,N_13583,N_13013);
xor U14613 (N_14613,N_13392,N_13466);
xor U14614 (N_14614,N_13746,N_13471);
or U14615 (N_14615,N_13002,N_13450);
or U14616 (N_14616,N_13654,N_13898);
and U14617 (N_14617,N_13364,N_13723);
nor U14618 (N_14618,N_13745,N_13636);
xnor U14619 (N_14619,N_13402,N_13491);
and U14620 (N_14620,N_13621,N_13093);
xor U14621 (N_14621,N_13306,N_13403);
or U14622 (N_14622,N_13744,N_13856);
nand U14623 (N_14623,N_13948,N_13903);
or U14624 (N_14624,N_13532,N_13033);
nor U14625 (N_14625,N_13966,N_13054);
or U14626 (N_14626,N_13727,N_13988);
nor U14627 (N_14627,N_13094,N_13424);
xor U14628 (N_14628,N_13044,N_13482);
and U14629 (N_14629,N_13845,N_13017);
xor U14630 (N_14630,N_13324,N_13953);
or U14631 (N_14631,N_13797,N_13643);
nand U14632 (N_14632,N_13574,N_13482);
nand U14633 (N_14633,N_13709,N_13337);
or U14634 (N_14634,N_13061,N_13701);
nand U14635 (N_14635,N_13557,N_13348);
nor U14636 (N_14636,N_13038,N_13331);
nand U14637 (N_14637,N_13727,N_13286);
xnor U14638 (N_14638,N_13540,N_13410);
nor U14639 (N_14639,N_13801,N_13595);
and U14640 (N_14640,N_13827,N_13562);
nor U14641 (N_14641,N_13144,N_13737);
nor U14642 (N_14642,N_13661,N_13375);
xor U14643 (N_14643,N_13799,N_13190);
nand U14644 (N_14644,N_13998,N_13215);
or U14645 (N_14645,N_13831,N_13379);
and U14646 (N_14646,N_13550,N_13243);
nor U14647 (N_14647,N_13106,N_13119);
or U14648 (N_14648,N_13128,N_13011);
xor U14649 (N_14649,N_13418,N_13399);
xor U14650 (N_14650,N_13400,N_13877);
and U14651 (N_14651,N_13976,N_13424);
nor U14652 (N_14652,N_13967,N_13823);
nor U14653 (N_14653,N_13719,N_13806);
and U14654 (N_14654,N_13084,N_13898);
and U14655 (N_14655,N_13014,N_13396);
or U14656 (N_14656,N_13960,N_13879);
nand U14657 (N_14657,N_13438,N_13684);
xor U14658 (N_14658,N_13673,N_13193);
nor U14659 (N_14659,N_13025,N_13267);
and U14660 (N_14660,N_13550,N_13643);
or U14661 (N_14661,N_13801,N_13068);
or U14662 (N_14662,N_13179,N_13975);
or U14663 (N_14663,N_13228,N_13499);
and U14664 (N_14664,N_13751,N_13526);
and U14665 (N_14665,N_13202,N_13940);
or U14666 (N_14666,N_13227,N_13257);
xnor U14667 (N_14667,N_13278,N_13763);
nor U14668 (N_14668,N_13854,N_13466);
nand U14669 (N_14669,N_13633,N_13877);
or U14670 (N_14670,N_13266,N_13875);
nor U14671 (N_14671,N_13410,N_13392);
or U14672 (N_14672,N_13499,N_13113);
and U14673 (N_14673,N_13681,N_13207);
xnor U14674 (N_14674,N_13144,N_13355);
and U14675 (N_14675,N_13562,N_13915);
and U14676 (N_14676,N_13752,N_13192);
and U14677 (N_14677,N_13459,N_13352);
xor U14678 (N_14678,N_13374,N_13215);
or U14679 (N_14679,N_13061,N_13936);
xnor U14680 (N_14680,N_13377,N_13335);
and U14681 (N_14681,N_13554,N_13599);
nor U14682 (N_14682,N_13703,N_13739);
or U14683 (N_14683,N_13755,N_13934);
nand U14684 (N_14684,N_13838,N_13771);
nand U14685 (N_14685,N_13647,N_13982);
nor U14686 (N_14686,N_13859,N_13450);
and U14687 (N_14687,N_13866,N_13369);
nor U14688 (N_14688,N_13399,N_13528);
and U14689 (N_14689,N_13694,N_13816);
or U14690 (N_14690,N_13578,N_13986);
xnor U14691 (N_14691,N_13087,N_13777);
or U14692 (N_14692,N_13740,N_13368);
nor U14693 (N_14693,N_13838,N_13166);
xor U14694 (N_14694,N_13605,N_13993);
and U14695 (N_14695,N_13704,N_13171);
and U14696 (N_14696,N_13048,N_13138);
xnor U14697 (N_14697,N_13286,N_13697);
and U14698 (N_14698,N_13531,N_13844);
or U14699 (N_14699,N_13676,N_13068);
or U14700 (N_14700,N_13116,N_13149);
nand U14701 (N_14701,N_13317,N_13391);
or U14702 (N_14702,N_13479,N_13898);
and U14703 (N_14703,N_13807,N_13137);
nand U14704 (N_14704,N_13141,N_13066);
nor U14705 (N_14705,N_13164,N_13355);
or U14706 (N_14706,N_13212,N_13716);
or U14707 (N_14707,N_13636,N_13066);
or U14708 (N_14708,N_13210,N_13264);
and U14709 (N_14709,N_13339,N_13465);
nor U14710 (N_14710,N_13971,N_13892);
or U14711 (N_14711,N_13132,N_13843);
or U14712 (N_14712,N_13230,N_13431);
nor U14713 (N_14713,N_13003,N_13993);
xnor U14714 (N_14714,N_13040,N_13201);
xor U14715 (N_14715,N_13492,N_13927);
and U14716 (N_14716,N_13786,N_13626);
nor U14717 (N_14717,N_13882,N_13608);
and U14718 (N_14718,N_13827,N_13308);
and U14719 (N_14719,N_13469,N_13654);
nand U14720 (N_14720,N_13989,N_13659);
xor U14721 (N_14721,N_13149,N_13499);
or U14722 (N_14722,N_13444,N_13064);
nand U14723 (N_14723,N_13287,N_13386);
and U14724 (N_14724,N_13145,N_13058);
or U14725 (N_14725,N_13245,N_13665);
or U14726 (N_14726,N_13727,N_13810);
nand U14727 (N_14727,N_13549,N_13136);
and U14728 (N_14728,N_13720,N_13937);
nand U14729 (N_14729,N_13429,N_13731);
nor U14730 (N_14730,N_13260,N_13107);
nor U14731 (N_14731,N_13717,N_13921);
or U14732 (N_14732,N_13476,N_13921);
nand U14733 (N_14733,N_13671,N_13188);
nor U14734 (N_14734,N_13626,N_13629);
or U14735 (N_14735,N_13434,N_13895);
and U14736 (N_14736,N_13276,N_13943);
or U14737 (N_14737,N_13423,N_13461);
and U14738 (N_14738,N_13824,N_13635);
nor U14739 (N_14739,N_13609,N_13608);
nand U14740 (N_14740,N_13949,N_13937);
xnor U14741 (N_14741,N_13721,N_13725);
and U14742 (N_14742,N_13587,N_13422);
nor U14743 (N_14743,N_13396,N_13102);
nor U14744 (N_14744,N_13837,N_13831);
nand U14745 (N_14745,N_13019,N_13533);
nor U14746 (N_14746,N_13463,N_13978);
nor U14747 (N_14747,N_13734,N_13876);
or U14748 (N_14748,N_13413,N_13243);
nand U14749 (N_14749,N_13996,N_13127);
nor U14750 (N_14750,N_13702,N_13086);
xnor U14751 (N_14751,N_13668,N_13717);
or U14752 (N_14752,N_13911,N_13024);
nor U14753 (N_14753,N_13631,N_13718);
xnor U14754 (N_14754,N_13769,N_13763);
nand U14755 (N_14755,N_13895,N_13737);
xor U14756 (N_14756,N_13583,N_13839);
nand U14757 (N_14757,N_13112,N_13381);
nand U14758 (N_14758,N_13111,N_13705);
nor U14759 (N_14759,N_13456,N_13009);
and U14760 (N_14760,N_13733,N_13750);
nor U14761 (N_14761,N_13366,N_13997);
and U14762 (N_14762,N_13788,N_13177);
nand U14763 (N_14763,N_13767,N_13728);
nand U14764 (N_14764,N_13504,N_13209);
and U14765 (N_14765,N_13354,N_13041);
xnor U14766 (N_14766,N_13303,N_13035);
and U14767 (N_14767,N_13483,N_13137);
and U14768 (N_14768,N_13039,N_13615);
nor U14769 (N_14769,N_13430,N_13483);
nand U14770 (N_14770,N_13316,N_13094);
xor U14771 (N_14771,N_13437,N_13841);
and U14772 (N_14772,N_13268,N_13416);
nand U14773 (N_14773,N_13343,N_13028);
xnor U14774 (N_14774,N_13889,N_13011);
xor U14775 (N_14775,N_13069,N_13291);
nand U14776 (N_14776,N_13202,N_13736);
or U14777 (N_14777,N_13631,N_13063);
nor U14778 (N_14778,N_13154,N_13721);
nor U14779 (N_14779,N_13321,N_13721);
nand U14780 (N_14780,N_13985,N_13899);
nor U14781 (N_14781,N_13224,N_13145);
nand U14782 (N_14782,N_13915,N_13355);
nor U14783 (N_14783,N_13896,N_13109);
nand U14784 (N_14784,N_13926,N_13066);
and U14785 (N_14785,N_13096,N_13907);
or U14786 (N_14786,N_13915,N_13151);
nor U14787 (N_14787,N_13063,N_13021);
and U14788 (N_14788,N_13556,N_13964);
and U14789 (N_14789,N_13570,N_13721);
nor U14790 (N_14790,N_13126,N_13788);
and U14791 (N_14791,N_13914,N_13037);
or U14792 (N_14792,N_13513,N_13929);
nor U14793 (N_14793,N_13037,N_13794);
and U14794 (N_14794,N_13182,N_13263);
or U14795 (N_14795,N_13862,N_13506);
nor U14796 (N_14796,N_13595,N_13723);
nor U14797 (N_14797,N_13538,N_13860);
and U14798 (N_14798,N_13514,N_13875);
nand U14799 (N_14799,N_13316,N_13783);
and U14800 (N_14800,N_13326,N_13243);
nor U14801 (N_14801,N_13871,N_13610);
nor U14802 (N_14802,N_13052,N_13568);
or U14803 (N_14803,N_13496,N_13239);
xor U14804 (N_14804,N_13206,N_13780);
nor U14805 (N_14805,N_13321,N_13625);
and U14806 (N_14806,N_13347,N_13051);
or U14807 (N_14807,N_13379,N_13364);
nor U14808 (N_14808,N_13114,N_13578);
nand U14809 (N_14809,N_13889,N_13376);
nand U14810 (N_14810,N_13798,N_13630);
xor U14811 (N_14811,N_13116,N_13199);
xor U14812 (N_14812,N_13881,N_13666);
xor U14813 (N_14813,N_13097,N_13186);
nand U14814 (N_14814,N_13325,N_13527);
nor U14815 (N_14815,N_13747,N_13366);
or U14816 (N_14816,N_13057,N_13835);
nand U14817 (N_14817,N_13276,N_13120);
nor U14818 (N_14818,N_13720,N_13104);
nor U14819 (N_14819,N_13731,N_13255);
or U14820 (N_14820,N_13837,N_13121);
nand U14821 (N_14821,N_13457,N_13783);
and U14822 (N_14822,N_13686,N_13394);
or U14823 (N_14823,N_13186,N_13242);
and U14824 (N_14824,N_13666,N_13285);
and U14825 (N_14825,N_13588,N_13725);
xor U14826 (N_14826,N_13308,N_13496);
nand U14827 (N_14827,N_13587,N_13977);
nand U14828 (N_14828,N_13941,N_13416);
nand U14829 (N_14829,N_13984,N_13905);
xnor U14830 (N_14830,N_13288,N_13135);
and U14831 (N_14831,N_13607,N_13410);
or U14832 (N_14832,N_13618,N_13741);
nor U14833 (N_14833,N_13235,N_13497);
nand U14834 (N_14834,N_13850,N_13295);
xor U14835 (N_14835,N_13461,N_13988);
xnor U14836 (N_14836,N_13136,N_13551);
xnor U14837 (N_14837,N_13025,N_13246);
xor U14838 (N_14838,N_13054,N_13788);
nand U14839 (N_14839,N_13004,N_13869);
xor U14840 (N_14840,N_13348,N_13005);
or U14841 (N_14841,N_13306,N_13916);
xnor U14842 (N_14842,N_13432,N_13173);
and U14843 (N_14843,N_13741,N_13405);
and U14844 (N_14844,N_13018,N_13615);
and U14845 (N_14845,N_13765,N_13003);
or U14846 (N_14846,N_13407,N_13063);
xnor U14847 (N_14847,N_13370,N_13560);
and U14848 (N_14848,N_13567,N_13171);
xor U14849 (N_14849,N_13921,N_13931);
nand U14850 (N_14850,N_13252,N_13316);
nand U14851 (N_14851,N_13441,N_13306);
or U14852 (N_14852,N_13049,N_13655);
and U14853 (N_14853,N_13592,N_13335);
nor U14854 (N_14854,N_13934,N_13483);
xor U14855 (N_14855,N_13979,N_13596);
and U14856 (N_14856,N_13745,N_13661);
nor U14857 (N_14857,N_13981,N_13754);
and U14858 (N_14858,N_13017,N_13834);
nor U14859 (N_14859,N_13444,N_13943);
nand U14860 (N_14860,N_13305,N_13496);
or U14861 (N_14861,N_13287,N_13557);
xnor U14862 (N_14862,N_13477,N_13242);
nand U14863 (N_14863,N_13754,N_13107);
nand U14864 (N_14864,N_13953,N_13736);
xor U14865 (N_14865,N_13520,N_13673);
xor U14866 (N_14866,N_13197,N_13519);
xor U14867 (N_14867,N_13644,N_13113);
nand U14868 (N_14868,N_13465,N_13616);
nor U14869 (N_14869,N_13276,N_13936);
xnor U14870 (N_14870,N_13638,N_13507);
and U14871 (N_14871,N_13224,N_13995);
and U14872 (N_14872,N_13766,N_13349);
xor U14873 (N_14873,N_13108,N_13927);
xor U14874 (N_14874,N_13809,N_13622);
nor U14875 (N_14875,N_13149,N_13011);
xor U14876 (N_14876,N_13880,N_13503);
nor U14877 (N_14877,N_13199,N_13372);
and U14878 (N_14878,N_13094,N_13785);
nor U14879 (N_14879,N_13147,N_13523);
nor U14880 (N_14880,N_13562,N_13958);
nand U14881 (N_14881,N_13945,N_13558);
nor U14882 (N_14882,N_13230,N_13754);
nor U14883 (N_14883,N_13679,N_13329);
nand U14884 (N_14884,N_13931,N_13686);
or U14885 (N_14885,N_13610,N_13257);
xnor U14886 (N_14886,N_13103,N_13698);
nor U14887 (N_14887,N_13172,N_13760);
and U14888 (N_14888,N_13998,N_13565);
or U14889 (N_14889,N_13369,N_13808);
nand U14890 (N_14890,N_13355,N_13876);
or U14891 (N_14891,N_13740,N_13597);
and U14892 (N_14892,N_13500,N_13645);
xor U14893 (N_14893,N_13565,N_13165);
nor U14894 (N_14894,N_13924,N_13560);
or U14895 (N_14895,N_13673,N_13761);
nor U14896 (N_14896,N_13836,N_13867);
and U14897 (N_14897,N_13591,N_13098);
nor U14898 (N_14898,N_13385,N_13443);
or U14899 (N_14899,N_13673,N_13628);
xor U14900 (N_14900,N_13907,N_13395);
xnor U14901 (N_14901,N_13857,N_13850);
xor U14902 (N_14902,N_13878,N_13986);
or U14903 (N_14903,N_13208,N_13138);
xnor U14904 (N_14904,N_13559,N_13618);
nor U14905 (N_14905,N_13112,N_13924);
nor U14906 (N_14906,N_13317,N_13962);
nand U14907 (N_14907,N_13707,N_13463);
or U14908 (N_14908,N_13668,N_13510);
nor U14909 (N_14909,N_13300,N_13777);
nor U14910 (N_14910,N_13683,N_13380);
and U14911 (N_14911,N_13483,N_13262);
xor U14912 (N_14912,N_13730,N_13001);
and U14913 (N_14913,N_13500,N_13545);
nor U14914 (N_14914,N_13024,N_13839);
nor U14915 (N_14915,N_13372,N_13037);
nor U14916 (N_14916,N_13039,N_13630);
or U14917 (N_14917,N_13161,N_13224);
nand U14918 (N_14918,N_13738,N_13193);
nand U14919 (N_14919,N_13324,N_13593);
or U14920 (N_14920,N_13254,N_13380);
nor U14921 (N_14921,N_13979,N_13967);
nand U14922 (N_14922,N_13948,N_13536);
nor U14923 (N_14923,N_13202,N_13226);
xnor U14924 (N_14924,N_13432,N_13403);
xnor U14925 (N_14925,N_13051,N_13903);
nor U14926 (N_14926,N_13479,N_13595);
nand U14927 (N_14927,N_13057,N_13869);
nand U14928 (N_14928,N_13435,N_13487);
xnor U14929 (N_14929,N_13661,N_13961);
nor U14930 (N_14930,N_13780,N_13578);
or U14931 (N_14931,N_13386,N_13410);
nor U14932 (N_14932,N_13042,N_13802);
nand U14933 (N_14933,N_13593,N_13114);
xnor U14934 (N_14934,N_13541,N_13502);
or U14935 (N_14935,N_13469,N_13495);
nor U14936 (N_14936,N_13568,N_13806);
and U14937 (N_14937,N_13867,N_13707);
and U14938 (N_14938,N_13895,N_13190);
or U14939 (N_14939,N_13847,N_13614);
xor U14940 (N_14940,N_13619,N_13761);
nor U14941 (N_14941,N_13305,N_13432);
nand U14942 (N_14942,N_13608,N_13363);
nor U14943 (N_14943,N_13509,N_13816);
nand U14944 (N_14944,N_13227,N_13846);
nand U14945 (N_14945,N_13188,N_13507);
xnor U14946 (N_14946,N_13301,N_13811);
nand U14947 (N_14947,N_13407,N_13205);
nand U14948 (N_14948,N_13054,N_13762);
and U14949 (N_14949,N_13655,N_13246);
nand U14950 (N_14950,N_13135,N_13639);
or U14951 (N_14951,N_13213,N_13555);
nand U14952 (N_14952,N_13385,N_13912);
and U14953 (N_14953,N_13091,N_13662);
xnor U14954 (N_14954,N_13591,N_13272);
or U14955 (N_14955,N_13955,N_13849);
nor U14956 (N_14956,N_13401,N_13130);
nand U14957 (N_14957,N_13793,N_13817);
nor U14958 (N_14958,N_13338,N_13230);
and U14959 (N_14959,N_13833,N_13326);
nor U14960 (N_14960,N_13068,N_13553);
or U14961 (N_14961,N_13986,N_13290);
and U14962 (N_14962,N_13522,N_13116);
nand U14963 (N_14963,N_13526,N_13753);
xnor U14964 (N_14964,N_13347,N_13147);
and U14965 (N_14965,N_13894,N_13621);
nor U14966 (N_14966,N_13272,N_13630);
and U14967 (N_14967,N_13432,N_13969);
and U14968 (N_14968,N_13577,N_13796);
and U14969 (N_14969,N_13701,N_13436);
nor U14970 (N_14970,N_13668,N_13050);
nand U14971 (N_14971,N_13518,N_13269);
or U14972 (N_14972,N_13492,N_13981);
and U14973 (N_14973,N_13287,N_13897);
and U14974 (N_14974,N_13006,N_13878);
and U14975 (N_14975,N_13202,N_13553);
and U14976 (N_14976,N_13197,N_13994);
nor U14977 (N_14977,N_13705,N_13043);
nor U14978 (N_14978,N_13014,N_13091);
or U14979 (N_14979,N_13568,N_13807);
xor U14980 (N_14980,N_13688,N_13278);
nand U14981 (N_14981,N_13174,N_13502);
and U14982 (N_14982,N_13598,N_13486);
xnor U14983 (N_14983,N_13334,N_13609);
or U14984 (N_14984,N_13455,N_13108);
and U14985 (N_14985,N_13641,N_13363);
nor U14986 (N_14986,N_13211,N_13261);
xor U14987 (N_14987,N_13086,N_13873);
nand U14988 (N_14988,N_13603,N_13053);
xor U14989 (N_14989,N_13269,N_13557);
nand U14990 (N_14990,N_13250,N_13964);
xnor U14991 (N_14991,N_13579,N_13031);
xnor U14992 (N_14992,N_13100,N_13480);
and U14993 (N_14993,N_13913,N_13783);
nor U14994 (N_14994,N_13476,N_13729);
xnor U14995 (N_14995,N_13928,N_13038);
or U14996 (N_14996,N_13825,N_13237);
or U14997 (N_14997,N_13843,N_13518);
nor U14998 (N_14998,N_13071,N_13815);
xor U14999 (N_14999,N_13433,N_13754);
nor U15000 (N_15000,N_14931,N_14202);
or U15001 (N_15001,N_14616,N_14155);
and U15002 (N_15002,N_14986,N_14469);
and U15003 (N_15003,N_14493,N_14165);
nor U15004 (N_15004,N_14452,N_14848);
or U15005 (N_15005,N_14892,N_14370);
and U15006 (N_15006,N_14478,N_14223);
nor U15007 (N_15007,N_14160,N_14828);
or U15008 (N_15008,N_14689,N_14062);
xnor U15009 (N_15009,N_14523,N_14617);
and U15010 (N_15010,N_14387,N_14188);
xnor U15011 (N_15011,N_14681,N_14106);
nor U15012 (N_15012,N_14210,N_14095);
xnor U15013 (N_15013,N_14415,N_14485);
and U15014 (N_15014,N_14395,N_14167);
nand U15015 (N_15015,N_14000,N_14050);
nand U15016 (N_15016,N_14655,N_14433);
nor U15017 (N_15017,N_14268,N_14683);
xnor U15018 (N_15018,N_14358,N_14653);
and U15019 (N_15019,N_14646,N_14135);
nand U15020 (N_15020,N_14814,N_14938);
and U15021 (N_15021,N_14067,N_14317);
or U15022 (N_15022,N_14075,N_14034);
nor U15023 (N_15023,N_14905,N_14934);
or U15024 (N_15024,N_14988,N_14163);
and U15025 (N_15025,N_14791,N_14593);
or U15026 (N_15026,N_14103,N_14968);
xor U15027 (N_15027,N_14212,N_14325);
nor U15028 (N_15028,N_14482,N_14271);
xor U15029 (N_15029,N_14102,N_14276);
xnor U15030 (N_15030,N_14760,N_14007);
nand U15031 (N_15031,N_14525,N_14498);
xnor U15032 (N_15032,N_14115,N_14782);
xnor U15033 (N_15033,N_14451,N_14394);
or U15034 (N_15034,N_14870,N_14954);
nor U15035 (N_15035,N_14418,N_14648);
nor U15036 (N_15036,N_14408,N_14149);
and U15037 (N_15037,N_14013,N_14471);
nor U15038 (N_15038,N_14804,N_14726);
xor U15039 (N_15039,N_14048,N_14477);
and U15040 (N_15040,N_14383,N_14625);
nor U15041 (N_15041,N_14561,N_14156);
xor U15042 (N_15042,N_14083,N_14239);
nor U15043 (N_15043,N_14707,N_14173);
nand U15044 (N_15044,N_14295,N_14659);
nand U15045 (N_15045,N_14093,N_14704);
and U15046 (N_15046,N_14594,N_14855);
and U15047 (N_15047,N_14565,N_14654);
or U15048 (N_15048,N_14425,N_14518);
and U15049 (N_15049,N_14833,N_14566);
xor U15050 (N_15050,N_14090,N_14049);
nor U15051 (N_15051,N_14448,N_14830);
xor U15052 (N_15052,N_14950,N_14001);
xor U15053 (N_15053,N_14436,N_14789);
nor U15054 (N_15054,N_14227,N_14628);
nor U15055 (N_15055,N_14835,N_14423);
and U15056 (N_15056,N_14132,N_14304);
nand U15057 (N_15057,N_14715,N_14169);
and U15058 (N_15058,N_14308,N_14738);
and U15059 (N_15059,N_14720,N_14144);
nand U15060 (N_15060,N_14601,N_14311);
xnor U15061 (N_15061,N_14912,N_14813);
nand U15062 (N_15062,N_14261,N_14060);
xor U15063 (N_15063,N_14906,N_14230);
nor U15064 (N_15064,N_14410,N_14140);
and U15065 (N_15065,N_14762,N_14357);
and U15066 (N_15066,N_14035,N_14164);
and U15067 (N_15067,N_14059,N_14189);
nor U15068 (N_15068,N_14945,N_14520);
nand U15069 (N_15069,N_14454,N_14296);
or U15070 (N_15070,N_14610,N_14382);
xor U15071 (N_15071,N_14922,N_14618);
xnor U15072 (N_15072,N_14854,N_14107);
and U15073 (N_15073,N_14248,N_14439);
or U15074 (N_15074,N_14320,N_14861);
or U15075 (N_15075,N_14669,N_14850);
nor U15076 (N_15076,N_14853,N_14199);
or U15077 (N_15077,N_14475,N_14897);
or U15078 (N_15078,N_14764,N_14006);
nand U15079 (N_15079,N_14840,N_14122);
nand U15080 (N_15080,N_14399,N_14919);
xor U15081 (N_15081,N_14847,N_14379);
nor U15082 (N_15082,N_14688,N_14576);
or U15083 (N_15083,N_14389,N_14258);
or U15084 (N_15084,N_14825,N_14590);
nor U15085 (N_15085,N_14647,N_14925);
xnor U15086 (N_15086,N_14880,N_14815);
nand U15087 (N_15087,N_14303,N_14005);
xnor U15088 (N_15088,N_14966,N_14392);
nand U15089 (N_15089,N_14717,N_14026);
and U15090 (N_15090,N_14728,N_14204);
or U15091 (N_15091,N_14624,N_14547);
xnor U15092 (N_15092,N_14709,N_14935);
xnor U15093 (N_15093,N_14930,N_14595);
nor U15094 (N_15094,N_14335,N_14371);
nand U15095 (N_15095,N_14578,N_14413);
or U15096 (N_15096,N_14642,N_14974);
xnor U15097 (N_15097,N_14264,N_14043);
and U15098 (N_15098,N_14114,N_14176);
nor U15099 (N_15099,N_14354,N_14290);
xor U15100 (N_15100,N_14228,N_14432);
and U15101 (N_15101,N_14332,N_14197);
nand U15102 (N_15102,N_14723,N_14277);
or U15103 (N_15103,N_14041,N_14077);
or U15104 (N_15104,N_14591,N_14573);
nor U15105 (N_15105,N_14430,N_14645);
or U15106 (N_15106,N_14238,N_14299);
nand U15107 (N_15107,N_14535,N_14839);
or U15108 (N_15108,N_14801,N_14231);
or U15109 (N_15109,N_14592,N_14080);
or U15110 (N_15110,N_14893,N_14891);
nand U15111 (N_15111,N_14722,N_14929);
or U15112 (N_15112,N_14445,N_14622);
and U15113 (N_15113,N_14241,N_14047);
nor U15114 (N_15114,N_14860,N_14606);
nand U15115 (N_15115,N_14372,N_14073);
nor U15116 (N_15116,N_14703,N_14812);
or U15117 (N_15117,N_14509,N_14914);
xnor U15118 (N_15118,N_14033,N_14965);
nand U15119 (N_15119,N_14406,N_14698);
xnor U15120 (N_15120,N_14908,N_14958);
or U15121 (N_15121,N_14031,N_14676);
nand U15122 (N_15122,N_14883,N_14401);
or U15123 (N_15123,N_14548,N_14443);
and U15124 (N_15124,N_14447,N_14611);
xor U15125 (N_15125,N_14602,N_14154);
xor U15126 (N_15126,N_14810,N_14362);
nand U15127 (N_15127,N_14461,N_14262);
nor U15128 (N_15128,N_14240,N_14201);
or U15129 (N_15129,N_14824,N_14838);
and U15130 (N_15130,N_14352,N_14545);
nor U15131 (N_15131,N_14292,N_14657);
xnor U15132 (N_15132,N_14081,N_14397);
and U15133 (N_15133,N_14237,N_14856);
and U15134 (N_15134,N_14822,N_14719);
and U15135 (N_15135,N_14513,N_14976);
and U15136 (N_15136,N_14673,N_14046);
nand U15137 (N_15137,N_14586,N_14374);
nand U15138 (N_15138,N_14867,N_14110);
nor U15139 (N_15139,N_14143,N_14771);
xnor U15140 (N_15140,N_14881,N_14263);
or U15141 (N_15141,N_14318,N_14989);
nand U15142 (N_15142,N_14729,N_14514);
or U15143 (N_15143,N_14570,N_14329);
nor U15144 (N_15144,N_14419,N_14025);
xor U15145 (N_15145,N_14393,N_14817);
nor U15146 (N_15146,N_14342,N_14744);
nor U15147 (N_15147,N_14677,N_14569);
nor U15148 (N_15148,N_14932,N_14457);
nand U15149 (N_15149,N_14100,N_14118);
or U15150 (N_15150,N_14775,N_14137);
or U15151 (N_15151,N_14221,N_14533);
nor U15152 (N_15152,N_14428,N_14607);
or U15153 (N_15153,N_14270,N_14679);
nand U15154 (N_15154,N_14424,N_14711);
xnor U15155 (N_15155,N_14057,N_14288);
or U15156 (N_15156,N_14947,N_14437);
or U15157 (N_15157,N_14404,N_14843);
and U15158 (N_15158,N_14215,N_14269);
xor U15159 (N_15159,N_14038,N_14913);
nor U15160 (N_15160,N_14864,N_14472);
nor U15161 (N_15161,N_14384,N_14032);
nor U15162 (N_15162,N_14562,N_14536);
nand U15163 (N_15163,N_14195,N_14480);
or U15164 (N_15164,N_14126,N_14266);
nor U15165 (N_15165,N_14702,N_14249);
xor U15166 (N_15166,N_14313,N_14405);
and U15167 (N_15167,N_14596,N_14146);
nor U15168 (N_15168,N_14844,N_14846);
and U15169 (N_15169,N_14208,N_14076);
nor U15170 (N_15170,N_14613,N_14306);
or U15171 (N_15171,N_14633,N_14494);
xnor U15172 (N_15172,N_14427,N_14420);
and U15173 (N_15173,N_14141,N_14924);
xor U15174 (N_15174,N_14502,N_14869);
or U15175 (N_15175,N_14829,N_14203);
or U15176 (N_15176,N_14222,N_14984);
xor U15177 (N_15177,N_14367,N_14980);
nor U15178 (N_15178,N_14583,N_14667);
nor U15179 (N_15179,N_14641,N_14978);
nand U15180 (N_15180,N_14558,N_14730);
or U15181 (N_15181,N_14145,N_14663);
or U15182 (N_15182,N_14699,N_14884);
nand U15183 (N_15183,N_14064,N_14849);
nor U15184 (N_15184,N_14515,N_14130);
or U15185 (N_15185,N_14743,N_14429);
or U15186 (N_15186,N_14928,N_14759);
nand U15187 (N_15187,N_14507,N_14449);
xnor U15188 (N_15188,N_14800,N_14148);
or U15189 (N_15189,N_14307,N_14900);
and U15190 (N_15190,N_14585,N_14882);
and U15191 (N_15191,N_14716,N_14862);
or U15192 (N_15192,N_14125,N_14608);
nor U15193 (N_15193,N_14396,N_14435);
nand U15194 (N_15194,N_14024,N_14302);
nand U15195 (N_15195,N_14129,N_14746);
or U15196 (N_15196,N_14030,N_14467);
or U15197 (N_15197,N_14951,N_14944);
nand U15198 (N_15198,N_14766,N_14322);
nand U15199 (N_15199,N_14529,N_14421);
nand U15200 (N_15200,N_14138,N_14065);
and U15201 (N_15201,N_14735,N_14907);
nor U15202 (N_15202,N_14953,N_14124);
xor U15203 (N_15203,N_14002,N_14575);
or U15204 (N_15204,N_14021,N_14180);
xor U15205 (N_15205,N_14623,N_14267);
nor U15206 (N_15206,N_14982,N_14769);
and U15207 (N_15207,N_14708,N_14859);
xnor U15208 (N_15208,N_14301,N_14274);
nand U15209 (N_15209,N_14940,N_14456);
nor U15210 (N_15210,N_14783,N_14453);
xor U15211 (N_15211,N_14278,N_14629);
or U15212 (N_15212,N_14326,N_14084);
and U15213 (N_15213,N_14460,N_14336);
or U15214 (N_15214,N_14631,N_14923);
or U15215 (N_15215,N_14996,N_14211);
nand U15216 (N_15216,N_14273,N_14011);
xnor U15217 (N_15217,N_14732,N_14377);
nand U15218 (N_15218,N_14010,N_14054);
nor U15219 (N_15219,N_14580,N_14310);
or U15220 (N_15220,N_14373,N_14637);
nor U15221 (N_15221,N_14416,N_14793);
xnor U15222 (N_15222,N_14651,N_14555);
or U15223 (N_15223,N_14170,N_14634);
nor U15224 (N_15224,N_14995,N_14027);
or U15225 (N_15225,N_14158,N_14250);
nor U15226 (N_15226,N_14321,N_14538);
and U15227 (N_15227,N_14826,N_14462);
xnor U15228 (N_15228,N_14078,N_14464);
or U15229 (N_15229,N_14476,N_14564);
and U15230 (N_15230,N_14319,N_14243);
xor U15231 (N_15231,N_14577,N_14365);
or U15232 (N_15232,N_14508,N_14082);
nor U15233 (N_15233,N_14630,N_14971);
xor U15234 (N_15234,N_14560,N_14949);
xnor U15235 (N_15235,N_14094,N_14957);
and U15236 (N_15236,N_14487,N_14666);
and U15237 (N_15237,N_14973,N_14380);
nand U15238 (N_15238,N_14857,N_14640);
and U15239 (N_15239,N_14961,N_14582);
nand U15240 (N_15240,N_14684,N_14776);
and U15241 (N_15241,N_14589,N_14751);
and U15242 (N_15242,N_14187,N_14692);
or U15243 (N_15243,N_14123,N_14260);
xor U15244 (N_15244,N_14450,N_14092);
xor U15245 (N_15245,N_14499,N_14942);
and U15246 (N_15246,N_14153,N_14346);
xor U15247 (N_15247,N_14224,N_14470);
nor U15248 (N_15248,N_14386,N_14792);
nor U15249 (N_15249,N_14910,N_14754);
or U15250 (N_15250,N_14312,N_14946);
nand U15251 (N_15251,N_14851,N_14297);
nand U15252 (N_15252,N_14682,N_14511);
and U15253 (N_15253,N_14216,N_14168);
or U15254 (N_15254,N_14287,N_14400);
nand U15255 (N_15255,N_14504,N_14353);
nor U15256 (N_15256,N_14051,N_14740);
and U15257 (N_15257,N_14956,N_14600);
nand U15258 (N_15258,N_14015,N_14279);
nor U15259 (N_15259,N_14983,N_14119);
xor U15260 (N_15260,N_14757,N_14725);
nand U15261 (N_15261,N_14375,N_14805);
nor U15262 (N_15262,N_14434,N_14468);
or U15263 (N_15263,N_14541,N_14975);
or U15264 (N_15264,N_14823,N_14537);
or U15265 (N_15265,N_14294,N_14879);
xnor U15266 (N_15266,N_14876,N_14714);
xnor U15267 (N_15267,N_14012,N_14898);
or U15268 (N_15268,N_14661,N_14904);
nor U15269 (N_15269,N_14816,N_14852);
nor U15270 (N_15270,N_14255,N_14773);
nand U15271 (N_15271,N_14736,N_14172);
xor U15272 (N_15272,N_14438,N_14486);
and U15273 (N_15273,N_14779,N_14842);
xor U15274 (N_15274,N_14112,N_14678);
and U15275 (N_15275,N_14650,N_14972);
nand U15276 (N_15276,N_14915,N_14737);
xnor U15277 (N_15277,N_14497,N_14756);
nand U15278 (N_15278,N_14808,N_14331);
nor U15279 (N_15279,N_14785,N_14023);
nand U15280 (N_15280,N_14232,N_14670);
xnor U15281 (N_15281,N_14778,N_14183);
or U15282 (N_15282,N_14289,N_14970);
or U15283 (N_15283,N_14675,N_14894);
or U15284 (N_15284,N_14116,N_14489);
or U15285 (N_15285,N_14797,N_14712);
xor U15286 (N_15286,N_14016,N_14315);
or U15287 (N_15287,N_14526,N_14191);
nor U15288 (N_15288,N_14385,N_14705);
nand U15289 (N_15289,N_14557,N_14926);
and U15290 (N_15290,N_14841,N_14540);
xnor U15291 (N_15291,N_14798,N_14568);
xor U15292 (N_15292,N_14658,N_14411);
nor U15293 (N_15293,N_14672,N_14052);
or U15294 (N_15294,N_14542,N_14139);
or U15295 (N_15295,N_14086,N_14603);
or U15296 (N_15296,N_14977,N_14008);
nor U15297 (N_15297,N_14786,N_14559);
nor U15298 (N_15298,N_14936,N_14916);
nand U15299 (N_15299,N_14579,N_14638);
or U15300 (N_15300,N_14151,N_14327);
xor U15301 (N_15301,N_14903,N_14162);
and U15302 (N_15302,N_14739,N_14044);
nor U15303 (N_15303,N_14752,N_14175);
nand U15304 (N_15304,N_14398,N_14674);
xor U15305 (N_15305,N_14943,N_14865);
nand U15306 (N_15306,N_14587,N_14004);
and U15307 (N_15307,N_14376,N_14465);
nor U15308 (N_15308,N_14161,N_14710);
nand U15309 (N_15309,N_14442,N_14517);
nor U15310 (N_15310,N_14022,N_14981);
xnor U15311 (N_15311,N_14952,N_14403);
or U15312 (N_15312,N_14693,N_14831);
xnor U15313 (N_15313,N_14368,N_14390);
nor U15314 (N_15314,N_14422,N_14018);
or U15315 (N_15315,N_14117,N_14992);
and U15316 (N_15316,N_14889,N_14040);
and U15317 (N_15317,N_14696,N_14506);
nand U15318 (N_15318,N_14019,N_14334);
xor U15319 (N_15319,N_14567,N_14939);
nor U15320 (N_15320,N_14085,N_14781);
nor U15321 (N_15321,N_14056,N_14272);
or U15322 (N_15322,N_14473,N_14807);
nor U15323 (N_15323,N_14182,N_14099);
and U15324 (N_15324,N_14283,N_14484);
xor U15325 (N_15325,N_14788,N_14770);
and U15326 (N_15326,N_14747,N_14662);
xnor U15327 (N_15327,N_14753,N_14496);
xnor U15328 (N_15328,N_14528,N_14818);
and U15329 (N_15329,N_14369,N_14721);
or U15330 (N_15330,N_14909,N_14742);
nor U15331 (N_15331,N_14553,N_14495);
and U15332 (N_15332,N_14985,N_14694);
and U15333 (N_15333,N_14718,N_14444);
xor U15334 (N_15334,N_14074,N_14347);
nor U15335 (N_15335,N_14619,N_14820);
xnor U15336 (N_15336,N_14878,N_14402);
nand U15337 (N_15337,N_14656,N_14483);
xnor U15338 (N_15338,N_14921,N_14233);
nor U15339 (N_15339,N_14796,N_14556);
or U15340 (N_15340,N_14488,N_14474);
and U15341 (N_15341,N_14069,N_14933);
nand U15342 (N_15342,N_14323,N_14503);
nor U15343 (N_15343,N_14058,N_14522);
nand U15344 (N_15344,N_14868,N_14127);
nor U15345 (N_15345,N_14731,N_14045);
nor U15346 (N_15346,N_14257,N_14501);
and U15347 (N_15347,N_14190,N_14217);
and U15348 (N_15348,N_14068,N_14960);
nor U15349 (N_15349,N_14772,N_14177);
nor U15350 (N_15350,N_14519,N_14256);
or U15351 (N_15351,N_14811,N_14194);
xor U15352 (N_15352,N_14426,N_14079);
or U15353 (N_15353,N_14544,N_14293);
nor U15354 (N_15354,N_14096,N_14089);
xor U15355 (N_15355,N_14790,N_14874);
nand U15356 (N_15356,N_14660,N_14193);
nand U15357 (N_15357,N_14863,N_14282);
nand U15358 (N_15358,N_14604,N_14845);
or U15359 (N_15359,N_14254,N_14516);
xor U15360 (N_15360,N_14899,N_14236);
or U15361 (N_15361,N_14466,N_14340);
or U15362 (N_15362,N_14749,N_14113);
and U15363 (N_15363,N_14245,N_14539);
nor U15364 (N_15364,N_14458,N_14280);
and U15365 (N_15365,N_14361,N_14459);
nor U15366 (N_15366,N_14070,N_14134);
nand U15367 (N_15367,N_14324,N_14333);
or U15368 (N_15368,N_14991,N_14104);
nand U15369 (N_15369,N_14339,N_14955);
xnor U15370 (N_15370,N_14758,N_14407);
nor U15371 (N_15371,N_14774,N_14969);
nand U15372 (N_15372,N_14745,N_14902);
or U15373 (N_15373,N_14834,N_14087);
nor U15374 (N_15374,N_14455,N_14691);
nor U15375 (N_15375,N_14706,N_14777);
or U15376 (N_15376,N_14235,N_14214);
nor U15377 (N_15377,N_14098,N_14226);
nand U15378 (N_15378,N_14291,N_14987);
or U15379 (N_15379,N_14741,N_14755);
xnor U15380 (N_15380,N_14787,N_14341);
nor U15381 (N_15381,N_14351,N_14108);
nand U15382 (N_15382,N_14285,N_14330);
xor U15383 (N_15383,N_14534,N_14225);
and U15384 (N_15384,N_14524,N_14431);
and U15385 (N_15385,N_14120,N_14733);
and U15386 (N_15386,N_14993,N_14492);
nand U15387 (N_15387,N_14948,N_14588);
nand U15388 (N_15388,N_14875,N_14328);
nand U15389 (N_15389,N_14885,N_14171);
or U15390 (N_15390,N_14500,N_14441);
xnor U15391 (N_15391,N_14701,N_14055);
or U15392 (N_15392,N_14184,N_14795);
or U15393 (N_15393,N_14314,N_14364);
and U15394 (N_15394,N_14872,N_14136);
or U15395 (N_15395,N_14131,N_14213);
xor U15396 (N_15396,N_14802,N_14574);
nor U15397 (N_15397,N_14794,N_14609);
or U15398 (N_15398,N_14252,N_14598);
and U15399 (N_15399,N_14806,N_14409);
nor U15400 (N_15400,N_14111,N_14366);
and U15401 (N_15401,N_14552,N_14873);
and U15402 (N_15402,N_14748,N_14803);
nand U15403 (N_15403,N_14286,N_14554);
or U15404 (N_15404,N_14028,N_14999);
xnor U15405 (N_15405,N_14521,N_14166);
or U15406 (N_15406,N_14927,N_14490);
nor U15407 (N_15407,N_14029,N_14017);
and U15408 (N_15408,N_14799,N_14644);
xnor U15409 (N_15409,N_14546,N_14036);
and U15410 (N_15410,N_14381,N_14652);
or U15411 (N_15411,N_14877,N_14819);
xor U15412 (N_15412,N_14157,N_14234);
nand U15413 (N_15413,N_14097,N_14391);
and U15414 (N_15414,N_14837,N_14246);
nand U15415 (N_15415,N_14671,N_14896);
nor U15416 (N_15416,N_14042,N_14599);
and U15417 (N_15417,N_14886,N_14244);
and U15418 (N_15418,N_14152,N_14636);
nor U15419 (N_15419,N_14763,N_14920);
nor U15420 (N_15420,N_14229,N_14061);
or U15421 (N_15421,N_14871,N_14014);
nor U15422 (N_15422,N_14071,N_14680);
or U15423 (N_15423,N_14360,N_14962);
nand U15424 (N_15424,N_14780,N_14687);
or U15425 (N_15425,N_14414,N_14219);
and U15426 (N_15426,N_14697,N_14196);
xnor U15427 (N_15427,N_14531,N_14686);
or U15428 (N_15428,N_14298,N_14150);
nor U15429 (N_15429,N_14761,N_14639);
or U15430 (N_15430,N_14412,N_14388);
or U15431 (N_15431,N_14901,N_14614);
and U15432 (N_15432,N_14363,N_14765);
nor U15433 (N_15433,N_14265,N_14247);
nand U15434 (N_15434,N_14209,N_14344);
nand U15435 (N_15435,N_14020,N_14918);
or U15436 (N_15436,N_14178,N_14128);
or U15437 (N_15437,N_14990,N_14959);
nand U15438 (N_15438,N_14505,N_14997);
and U15439 (N_15439,N_14668,N_14887);
or U15440 (N_15440,N_14836,N_14037);
or U15441 (N_15441,N_14713,N_14481);
or U15442 (N_15442,N_14994,N_14727);
nand U15443 (N_15443,N_14581,N_14937);
nor U15444 (N_15444,N_14463,N_14527);
and U15445 (N_15445,N_14359,N_14890);
xor U15446 (N_15446,N_14192,N_14979);
nand U15447 (N_15447,N_14355,N_14185);
nand U15448 (N_15448,N_14345,N_14911);
xor U15449 (N_15449,N_14550,N_14417);
and U15450 (N_15450,N_14440,N_14300);
nand U15451 (N_15451,N_14147,N_14690);
and U15452 (N_15452,N_14337,N_14809);
nand U15453 (N_15453,N_14446,N_14091);
nor U15454 (N_15454,N_14003,N_14784);
nor U15455 (N_15455,N_14572,N_14009);
xnor U15456 (N_15456,N_14378,N_14917);
nand U15457 (N_15457,N_14597,N_14259);
nand U15458 (N_15458,N_14284,N_14734);
or U15459 (N_15459,N_14316,N_14612);
xor U15460 (N_15460,N_14685,N_14512);
or U15461 (N_15461,N_14088,N_14275);
xor U15462 (N_15462,N_14105,N_14242);
nand U15463 (N_15463,N_14700,N_14767);
nand U15464 (N_15464,N_14066,N_14343);
nor U15465 (N_15465,N_14615,N_14750);
or U15466 (N_15466,N_14253,N_14821);
or U15467 (N_15467,N_14063,N_14159);
nor U15468 (N_15468,N_14571,N_14109);
nor U15469 (N_15469,N_14281,N_14348);
or U15470 (N_15470,N_14998,N_14967);
xnor U15471 (N_15471,N_14626,N_14605);
or U15472 (N_15472,N_14072,N_14827);
and U15473 (N_15473,N_14510,N_14649);
nand U15474 (N_15474,N_14179,N_14479);
nand U15475 (N_15475,N_14866,N_14643);
xnor U15476 (N_15476,N_14620,N_14349);
and U15477 (N_15477,N_14724,N_14635);
or U15478 (N_15478,N_14220,N_14584);
and U15479 (N_15479,N_14858,N_14621);
nor U15480 (N_15480,N_14053,N_14532);
xnor U15481 (N_15481,N_14207,N_14200);
and U15482 (N_15482,N_14549,N_14206);
or U15483 (N_15483,N_14039,N_14174);
or U15484 (N_15484,N_14543,N_14491);
and U15485 (N_15485,N_14133,N_14627);
and U15486 (N_15486,N_14832,N_14205);
xnor U15487 (N_15487,N_14198,N_14695);
or U15488 (N_15488,N_14665,N_14768);
and U15489 (N_15489,N_14941,N_14181);
and U15490 (N_15490,N_14309,N_14551);
nor U15491 (N_15491,N_14186,N_14632);
or U15492 (N_15492,N_14121,N_14563);
nor U15493 (N_15493,N_14664,N_14350);
and U15494 (N_15494,N_14964,N_14888);
xnor U15495 (N_15495,N_14338,N_14895);
nand U15496 (N_15496,N_14356,N_14305);
or U15497 (N_15497,N_14142,N_14101);
nand U15498 (N_15498,N_14218,N_14963);
nor U15499 (N_15499,N_14530,N_14251);
nand U15500 (N_15500,N_14456,N_14084);
nor U15501 (N_15501,N_14767,N_14397);
nor U15502 (N_15502,N_14637,N_14679);
or U15503 (N_15503,N_14511,N_14733);
xnor U15504 (N_15504,N_14313,N_14985);
nor U15505 (N_15505,N_14477,N_14884);
or U15506 (N_15506,N_14961,N_14544);
xnor U15507 (N_15507,N_14892,N_14245);
nand U15508 (N_15508,N_14971,N_14311);
or U15509 (N_15509,N_14491,N_14936);
nand U15510 (N_15510,N_14884,N_14399);
and U15511 (N_15511,N_14870,N_14181);
nor U15512 (N_15512,N_14761,N_14485);
or U15513 (N_15513,N_14445,N_14870);
or U15514 (N_15514,N_14483,N_14281);
or U15515 (N_15515,N_14422,N_14258);
nand U15516 (N_15516,N_14708,N_14637);
and U15517 (N_15517,N_14491,N_14433);
xnor U15518 (N_15518,N_14564,N_14031);
nor U15519 (N_15519,N_14246,N_14963);
nand U15520 (N_15520,N_14594,N_14230);
xor U15521 (N_15521,N_14142,N_14500);
xnor U15522 (N_15522,N_14638,N_14179);
and U15523 (N_15523,N_14827,N_14810);
or U15524 (N_15524,N_14908,N_14941);
nor U15525 (N_15525,N_14420,N_14710);
nor U15526 (N_15526,N_14617,N_14581);
or U15527 (N_15527,N_14884,N_14768);
or U15528 (N_15528,N_14243,N_14375);
nor U15529 (N_15529,N_14536,N_14666);
nand U15530 (N_15530,N_14388,N_14643);
and U15531 (N_15531,N_14579,N_14011);
nand U15532 (N_15532,N_14596,N_14348);
or U15533 (N_15533,N_14831,N_14800);
and U15534 (N_15534,N_14743,N_14615);
nand U15535 (N_15535,N_14298,N_14659);
and U15536 (N_15536,N_14731,N_14950);
nand U15537 (N_15537,N_14838,N_14468);
xnor U15538 (N_15538,N_14729,N_14800);
nand U15539 (N_15539,N_14277,N_14047);
xnor U15540 (N_15540,N_14716,N_14662);
and U15541 (N_15541,N_14285,N_14687);
or U15542 (N_15542,N_14370,N_14688);
nand U15543 (N_15543,N_14740,N_14391);
nand U15544 (N_15544,N_14321,N_14111);
or U15545 (N_15545,N_14587,N_14130);
xnor U15546 (N_15546,N_14829,N_14993);
xnor U15547 (N_15547,N_14808,N_14344);
xor U15548 (N_15548,N_14468,N_14623);
nand U15549 (N_15549,N_14042,N_14959);
nand U15550 (N_15550,N_14157,N_14701);
or U15551 (N_15551,N_14345,N_14770);
xnor U15552 (N_15552,N_14078,N_14154);
nor U15553 (N_15553,N_14903,N_14119);
nor U15554 (N_15554,N_14855,N_14263);
xnor U15555 (N_15555,N_14404,N_14123);
or U15556 (N_15556,N_14069,N_14631);
xnor U15557 (N_15557,N_14132,N_14208);
xor U15558 (N_15558,N_14822,N_14439);
xnor U15559 (N_15559,N_14508,N_14334);
nand U15560 (N_15560,N_14139,N_14006);
nor U15561 (N_15561,N_14008,N_14139);
and U15562 (N_15562,N_14750,N_14628);
or U15563 (N_15563,N_14347,N_14077);
or U15564 (N_15564,N_14071,N_14600);
and U15565 (N_15565,N_14397,N_14236);
or U15566 (N_15566,N_14459,N_14059);
nor U15567 (N_15567,N_14343,N_14835);
or U15568 (N_15568,N_14872,N_14062);
or U15569 (N_15569,N_14410,N_14980);
nand U15570 (N_15570,N_14410,N_14763);
nor U15571 (N_15571,N_14033,N_14906);
and U15572 (N_15572,N_14499,N_14094);
and U15573 (N_15573,N_14020,N_14040);
or U15574 (N_15574,N_14491,N_14944);
nor U15575 (N_15575,N_14043,N_14484);
nand U15576 (N_15576,N_14380,N_14620);
and U15577 (N_15577,N_14999,N_14670);
xnor U15578 (N_15578,N_14698,N_14473);
nand U15579 (N_15579,N_14037,N_14136);
and U15580 (N_15580,N_14421,N_14116);
nand U15581 (N_15581,N_14163,N_14459);
xor U15582 (N_15582,N_14958,N_14791);
and U15583 (N_15583,N_14392,N_14451);
nor U15584 (N_15584,N_14889,N_14731);
or U15585 (N_15585,N_14893,N_14662);
or U15586 (N_15586,N_14694,N_14270);
or U15587 (N_15587,N_14407,N_14620);
xnor U15588 (N_15588,N_14798,N_14639);
or U15589 (N_15589,N_14685,N_14622);
or U15590 (N_15590,N_14666,N_14875);
nor U15591 (N_15591,N_14418,N_14626);
and U15592 (N_15592,N_14636,N_14364);
nand U15593 (N_15593,N_14223,N_14401);
xnor U15594 (N_15594,N_14917,N_14156);
xnor U15595 (N_15595,N_14071,N_14722);
nand U15596 (N_15596,N_14074,N_14738);
and U15597 (N_15597,N_14659,N_14254);
and U15598 (N_15598,N_14856,N_14103);
and U15599 (N_15599,N_14108,N_14271);
nand U15600 (N_15600,N_14781,N_14183);
nor U15601 (N_15601,N_14103,N_14016);
nand U15602 (N_15602,N_14553,N_14705);
xnor U15603 (N_15603,N_14609,N_14875);
and U15604 (N_15604,N_14861,N_14604);
and U15605 (N_15605,N_14324,N_14012);
and U15606 (N_15606,N_14583,N_14236);
or U15607 (N_15607,N_14182,N_14804);
and U15608 (N_15608,N_14033,N_14200);
xnor U15609 (N_15609,N_14850,N_14407);
nor U15610 (N_15610,N_14339,N_14465);
xor U15611 (N_15611,N_14138,N_14935);
and U15612 (N_15612,N_14914,N_14112);
or U15613 (N_15613,N_14688,N_14135);
nand U15614 (N_15614,N_14472,N_14192);
xor U15615 (N_15615,N_14036,N_14552);
xor U15616 (N_15616,N_14158,N_14655);
nand U15617 (N_15617,N_14624,N_14515);
and U15618 (N_15618,N_14821,N_14586);
or U15619 (N_15619,N_14390,N_14898);
nor U15620 (N_15620,N_14081,N_14828);
nor U15621 (N_15621,N_14380,N_14569);
nor U15622 (N_15622,N_14387,N_14424);
and U15623 (N_15623,N_14442,N_14670);
nand U15624 (N_15624,N_14177,N_14450);
nand U15625 (N_15625,N_14428,N_14773);
nand U15626 (N_15626,N_14786,N_14970);
xnor U15627 (N_15627,N_14156,N_14361);
and U15628 (N_15628,N_14500,N_14306);
or U15629 (N_15629,N_14703,N_14903);
and U15630 (N_15630,N_14987,N_14989);
nand U15631 (N_15631,N_14214,N_14807);
xor U15632 (N_15632,N_14037,N_14249);
and U15633 (N_15633,N_14156,N_14386);
or U15634 (N_15634,N_14062,N_14798);
nor U15635 (N_15635,N_14191,N_14960);
and U15636 (N_15636,N_14438,N_14040);
xor U15637 (N_15637,N_14224,N_14210);
nor U15638 (N_15638,N_14107,N_14601);
and U15639 (N_15639,N_14245,N_14133);
or U15640 (N_15640,N_14295,N_14181);
or U15641 (N_15641,N_14829,N_14825);
and U15642 (N_15642,N_14641,N_14752);
or U15643 (N_15643,N_14288,N_14918);
nand U15644 (N_15644,N_14016,N_14722);
or U15645 (N_15645,N_14300,N_14861);
and U15646 (N_15646,N_14060,N_14406);
nor U15647 (N_15647,N_14242,N_14167);
nor U15648 (N_15648,N_14721,N_14267);
xor U15649 (N_15649,N_14319,N_14309);
xnor U15650 (N_15650,N_14153,N_14698);
nand U15651 (N_15651,N_14832,N_14784);
and U15652 (N_15652,N_14660,N_14387);
or U15653 (N_15653,N_14352,N_14595);
nor U15654 (N_15654,N_14841,N_14347);
nor U15655 (N_15655,N_14314,N_14765);
and U15656 (N_15656,N_14404,N_14084);
nand U15657 (N_15657,N_14748,N_14233);
xor U15658 (N_15658,N_14458,N_14579);
or U15659 (N_15659,N_14845,N_14921);
and U15660 (N_15660,N_14359,N_14914);
nor U15661 (N_15661,N_14951,N_14150);
nor U15662 (N_15662,N_14374,N_14417);
nor U15663 (N_15663,N_14435,N_14540);
or U15664 (N_15664,N_14386,N_14405);
and U15665 (N_15665,N_14448,N_14133);
and U15666 (N_15666,N_14233,N_14494);
nor U15667 (N_15667,N_14817,N_14013);
nand U15668 (N_15668,N_14816,N_14349);
nor U15669 (N_15669,N_14541,N_14679);
or U15670 (N_15670,N_14125,N_14133);
and U15671 (N_15671,N_14081,N_14694);
xor U15672 (N_15672,N_14621,N_14480);
nor U15673 (N_15673,N_14319,N_14881);
or U15674 (N_15674,N_14602,N_14577);
nor U15675 (N_15675,N_14411,N_14962);
or U15676 (N_15676,N_14704,N_14364);
nand U15677 (N_15677,N_14296,N_14471);
nor U15678 (N_15678,N_14287,N_14007);
nand U15679 (N_15679,N_14733,N_14068);
or U15680 (N_15680,N_14379,N_14048);
nor U15681 (N_15681,N_14520,N_14131);
nor U15682 (N_15682,N_14127,N_14769);
xnor U15683 (N_15683,N_14420,N_14802);
and U15684 (N_15684,N_14373,N_14349);
or U15685 (N_15685,N_14476,N_14388);
nor U15686 (N_15686,N_14414,N_14595);
nor U15687 (N_15687,N_14869,N_14726);
or U15688 (N_15688,N_14627,N_14213);
or U15689 (N_15689,N_14405,N_14098);
and U15690 (N_15690,N_14285,N_14642);
nand U15691 (N_15691,N_14317,N_14560);
or U15692 (N_15692,N_14575,N_14493);
nor U15693 (N_15693,N_14984,N_14870);
or U15694 (N_15694,N_14903,N_14346);
xor U15695 (N_15695,N_14843,N_14406);
xnor U15696 (N_15696,N_14190,N_14923);
and U15697 (N_15697,N_14154,N_14683);
nand U15698 (N_15698,N_14312,N_14871);
and U15699 (N_15699,N_14383,N_14602);
or U15700 (N_15700,N_14839,N_14784);
and U15701 (N_15701,N_14008,N_14571);
xnor U15702 (N_15702,N_14499,N_14303);
nor U15703 (N_15703,N_14928,N_14817);
xor U15704 (N_15704,N_14688,N_14988);
nor U15705 (N_15705,N_14335,N_14533);
or U15706 (N_15706,N_14296,N_14409);
nand U15707 (N_15707,N_14332,N_14059);
nand U15708 (N_15708,N_14967,N_14776);
and U15709 (N_15709,N_14599,N_14916);
nor U15710 (N_15710,N_14503,N_14453);
xor U15711 (N_15711,N_14539,N_14935);
nand U15712 (N_15712,N_14419,N_14193);
xnor U15713 (N_15713,N_14207,N_14967);
and U15714 (N_15714,N_14801,N_14387);
xor U15715 (N_15715,N_14460,N_14244);
xnor U15716 (N_15716,N_14570,N_14699);
or U15717 (N_15717,N_14576,N_14344);
nor U15718 (N_15718,N_14247,N_14519);
or U15719 (N_15719,N_14767,N_14765);
nand U15720 (N_15720,N_14401,N_14180);
and U15721 (N_15721,N_14977,N_14730);
or U15722 (N_15722,N_14997,N_14448);
and U15723 (N_15723,N_14165,N_14092);
xor U15724 (N_15724,N_14462,N_14504);
or U15725 (N_15725,N_14963,N_14197);
nand U15726 (N_15726,N_14918,N_14843);
nor U15727 (N_15727,N_14926,N_14614);
nor U15728 (N_15728,N_14034,N_14353);
or U15729 (N_15729,N_14384,N_14281);
xor U15730 (N_15730,N_14562,N_14494);
nor U15731 (N_15731,N_14882,N_14267);
or U15732 (N_15732,N_14217,N_14363);
and U15733 (N_15733,N_14479,N_14260);
and U15734 (N_15734,N_14523,N_14720);
xnor U15735 (N_15735,N_14616,N_14350);
and U15736 (N_15736,N_14700,N_14480);
nand U15737 (N_15737,N_14404,N_14065);
nor U15738 (N_15738,N_14886,N_14305);
or U15739 (N_15739,N_14991,N_14512);
or U15740 (N_15740,N_14790,N_14433);
or U15741 (N_15741,N_14954,N_14071);
nor U15742 (N_15742,N_14000,N_14067);
nor U15743 (N_15743,N_14146,N_14482);
or U15744 (N_15744,N_14658,N_14277);
xor U15745 (N_15745,N_14249,N_14461);
nor U15746 (N_15746,N_14296,N_14564);
nand U15747 (N_15747,N_14432,N_14614);
or U15748 (N_15748,N_14970,N_14724);
xnor U15749 (N_15749,N_14027,N_14593);
xnor U15750 (N_15750,N_14340,N_14666);
and U15751 (N_15751,N_14490,N_14371);
or U15752 (N_15752,N_14659,N_14544);
nand U15753 (N_15753,N_14248,N_14243);
or U15754 (N_15754,N_14213,N_14705);
xnor U15755 (N_15755,N_14323,N_14505);
nor U15756 (N_15756,N_14261,N_14477);
nor U15757 (N_15757,N_14060,N_14798);
and U15758 (N_15758,N_14678,N_14541);
or U15759 (N_15759,N_14122,N_14544);
nor U15760 (N_15760,N_14495,N_14815);
nor U15761 (N_15761,N_14054,N_14938);
and U15762 (N_15762,N_14875,N_14808);
xnor U15763 (N_15763,N_14057,N_14903);
nor U15764 (N_15764,N_14610,N_14981);
nor U15765 (N_15765,N_14180,N_14632);
and U15766 (N_15766,N_14468,N_14905);
nor U15767 (N_15767,N_14141,N_14695);
nand U15768 (N_15768,N_14813,N_14983);
xnor U15769 (N_15769,N_14945,N_14959);
nor U15770 (N_15770,N_14394,N_14129);
nand U15771 (N_15771,N_14857,N_14383);
or U15772 (N_15772,N_14169,N_14263);
or U15773 (N_15773,N_14933,N_14574);
xnor U15774 (N_15774,N_14224,N_14602);
and U15775 (N_15775,N_14530,N_14378);
nand U15776 (N_15776,N_14576,N_14978);
nand U15777 (N_15777,N_14626,N_14163);
nand U15778 (N_15778,N_14200,N_14510);
nor U15779 (N_15779,N_14144,N_14520);
nand U15780 (N_15780,N_14826,N_14228);
xor U15781 (N_15781,N_14464,N_14980);
nor U15782 (N_15782,N_14101,N_14467);
or U15783 (N_15783,N_14650,N_14885);
xnor U15784 (N_15784,N_14461,N_14493);
nor U15785 (N_15785,N_14321,N_14080);
or U15786 (N_15786,N_14575,N_14550);
or U15787 (N_15787,N_14032,N_14042);
nor U15788 (N_15788,N_14905,N_14320);
xor U15789 (N_15789,N_14856,N_14815);
and U15790 (N_15790,N_14486,N_14113);
nand U15791 (N_15791,N_14546,N_14581);
nand U15792 (N_15792,N_14183,N_14425);
nand U15793 (N_15793,N_14993,N_14364);
xor U15794 (N_15794,N_14762,N_14270);
nor U15795 (N_15795,N_14306,N_14923);
nor U15796 (N_15796,N_14252,N_14680);
nand U15797 (N_15797,N_14782,N_14735);
xnor U15798 (N_15798,N_14785,N_14708);
and U15799 (N_15799,N_14342,N_14325);
or U15800 (N_15800,N_14932,N_14811);
nor U15801 (N_15801,N_14118,N_14032);
nand U15802 (N_15802,N_14294,N_14620);
xor U15803 (N_15803,N_14775,N_14093);
nor U15804 (N_15804,N_14195,N_14688);
nand U15805 (N_15805,N_14699,N_14285);
and U15806 (N_15806,N_14803,N_14521);
nor U15807 (N_15807,N_14680,N_14896);
xnor U15808 (N_15808,N_14498,N_14160);
or U15809 (N_15809,N_14810,N_14747);
or U15810 (N_15810,N_14338,N_14207);
nor U15811 (N_15811,N_14641,N_14595);
and U15812 (N_15812,N_14280,N_14324);
nor U15813 (N_15813,N_14644,N_14833);
and U15814 (N_15814,N_14504,N_14835);
nand U15815 (N_15815,N_14042,N_14112);
nand U15816 (N_15816,N_14313,N_14445);
nand U15817 (N_15817,N_14250,N_14664);
nand U15818 (N_15818,N_14281,N_14871);
nand U15819 (N_15819,N_14915,N_14326);
nand U15820 (N_15820,N_14754,N_14084);
nand U15821 (N_15821,N_14204,N_14748);
nor U15822 (N_15822,N_14030,N_14800);
xor U15823 (N_15823,N_14122,N_14119);
xnor U15824 (N_15824,N_14876,N_14599);
xnor U15825 (N_15825,N_14668,N_14947);
nor U15826 (N_15826,N_14779,N_14840);
nand U15827 (N_15827,N_14175,N_14077);
nand U15828 (N_15828,N_14079,N_14526);
nand U15829 (N_15829,N_14499,N_14284);
and U15830 (N_15830,N_14423,N_14567);
and U15831 (N_15831,N_14639,N_14082);
nand U15832 (N_15832,N_14559,N_14775);
nor U15833 (N_15833,N_14314,N_14373);
nand U15834 (N_15834,N_14054,N_14978);
nor U15835 (N_15835,N_14538,N_14100);
or U15836 (N_15836,N_14708,N_14447);
and U15837 (N_15837,N_14367,N_14366);
nand U15838 (N_15838,N_14462,N_14392);
or U15839 (N_15839,N_14469,N_14281);
or U15840 (N_15840,N_14124,N_14005);
and U15841 (N_15841,N_14269,N_14022);
and U15842 (N_15842,N_14955,N_14357);
and U15843 (N_15843,N_14071,N_14178);
and U15844 (N_15844,N_14954,N_14232);
and U15845 (N_15845,N_14557,N_14634);
and U15846 (N_15846,N_14102,N_14331);
xor U15847 (N_15847,N_14372,N_14176);
or U15848 (N_15848,N_14982,N_14803);
and U15849 (N_15849,N_14269,N_14132);
or U15850 (N_15850,N_14587,N_14376);
and U15851 (N_15851,N_14347,N_14646);
xnor U15852 (N_15852,N_14148,N_14887);
xnor U15853 (N_15853,N_14837,N_14990);
xor U15854 (N_15854,N_14470,N_14410);
or U15855 (N_15855,N_14484,N_14959);
xor U15856 (N_15856,N_14300,N_14561);
and U15857 (N_15857,N_14149,N_14517);
and U15858 (N_15858,N_14188,N_14554);
xor U15859 (N_15859,N_14072,N_14356);
nor U15860 (N_15860,N_14721,N_14386);
or U15861 (N_15861,N_14633,N_14487);
or U15862 (N_15862,N_14296,N_14498);
and U15863 (N_15863,N_14304,N_14040);
xnor U15864 (N_15864,N_14255,N_14243);
nand U15865 (N_15865,N_14442,N_14931);
and U15866 (N_15866,N_14539,N_14693);
and U15867 (N_15867,N_14797,N_14906);
or U15868 (N_15868,N_14238,N_14690);
and U15869 (N_15869,N_14124,N_14298);
xnor U15870 (N_15870,N_14264,N_14753);
and U15871 (N_15871,N_14153,N_14351);
and U15872 (N_15872,N_14873,N_14900);
and U15873 (N_15873,N_14407,N_14366);
nor U15874 (N_15874,N_14978,N_14929);
nor U15875 (N_15875,N_14836,N_14902);
xnor U15876 (N_15876,N_14623,N_14556);
nor U15877 (N_15877,N_14195,N_14200);
xor U15878 (N_15878,N_14163,N_14916);
nor U15879 (N_15879,N_14538,N_14219);
and U15880 (N_15880,N_14785,N_14354);
and U15881 (N_15881,N_14472,N_14665);
nand U15882 (N_15882,N_14364,N_14017);
nand U15883 (N_15883,N_14598,N_14817);
nor U15884 (N_15884,N_14920,N_14743);
or U15885 (N_15885,N_14432,N_14884);
xor U15886 (N_15886,N_14443,N_14097);
or U15887 (N_15887,N_14115,N_14422);
nand U15888 (N_15888,N_14281,N_14216);
nor U15889 (N_15889,N_14774,N_14975);
xor U15890 (N_15890,N_14875,N_14462);
and U15891 (N_15891,N_14647,N_14726);
xnor U15892 (N_15892,N_14816,N_14067);
nor U15893 (N_15893,N_14041,N_14103);
nor U15894 (N_15894,N_14898,N_14563);
and U15895 (N_15895,N_14575,N_14247);
xor U15896 (N_15896,N_14741,N_14231);
nor U15897 (N_15897,N_14085,N_14788);
or U15898 (N_15898,N_14913,N_14897);
or U15899 (N_15899,N_14720,N_14602);
nor U15900 (N_15900,N_14458,N_14162);
nand U15901 (N_15901,N_14327,N_14936);
nand U15902 (N_15902,N_14961,N_14637);
and U15903 (N_15903,N_14661,N_14019);
nor U15904 (N_15904,N_14690,N_14321);
nor U15905 (N_15905,N_14222,N_14179);
or U15906 (N_15906,N_14975,N_14245);
xor U15907 (N_15907,N_14663,N_14292);
or U15908 (N_15908,N_14896,N_14845);
or U15909 (N_15909,N_14525,N_14555);
and U15910 (N_15910,N_14853,N_14828);
nand U15911 (N_15911,N_14591,N_14193);
or U15912 (N_15912,N_14097,N_14918);
or U15913 (N_15913,N_14215,N_14838);
xor U15914 (N_15914,N_14200,N_14152);
nand U15915 (N_15915,N_14315,N_14607);
and U15916 (N_15916,N_14958,N_14670);
nor U15917 (N_15917,N_14864,N_14924);
or U15918 (N_15918,N_14461,N_14648);
or U15919 (N_15919,N_14533,N_14880);
and U15920 (N_15920,N_14731,N_14909);
nand U15921 (N_15921,N_14523,N_14626);
nor U15922 (N_15922,N_14865,N_14592);
and U15923 (N_15923,N_14767,N_14182);
nor U15924 (N_15924,N_14309,N_14866);
and U15925 (N_15925,N_14569,N_14277);
xnor U15926 (N_15926,N_14149,N_14520);
and U15927 (N_15927,N_14094,N_14039);
and U15928 (N_15928,N_14996,N_14621);
xor U15929 (N_15929,N_14740,N_14790);
or U15930 (N_15930,N_14421,N_14227);
nor U15931 (N_15931,N_14564,N_14902);
nor U15932 (N_15932,N_14211,N_14118);
xnor U15933 (N_15933,N_14733,N_14480);
nor U15934 (N_15934,N_14893,N_14095);
nand U15935 (N_15935,N_14201,N_14188);
xor U15936 (N_15936,N_14545,N_14240);
or U15937 (N_15937,N_14399,N_14445);
nor U15938 (N_15938,N_14281,N_14659);
xor U15939 (N_15939,N_14303,N_14667);
xor U15940 (N_15940,N_14798,N_14973);
nand U15941 (N_15941,N_14655,N_14206);
and U15942 (N_15942,N_14806,N_14095);
and U15943 (N_15943,N_14110,N_14248);
or U15944 (N_15944,N_14610,N_14424);
or U15945 (N_15945,N_14921,N_14936);
and U15946 (N_15946,N_14744,N_14009);
nand U15947 (N_15947,N_14274,N_14908);
xnor U15948 (N_15948,N_14414,N_14050);
nand U15949 (N_15949,N_14106,N_14139);
and U15950 (N_15950,N_14295,N_14991);
and U15951 (N_15951,N_14516,N_14533);
or U15952 (N_15952,N_14722,N_14983);
nor U15953 (N_15953,N_14913,N_14663);
or U15954 (N_15954,N_14709,N_14403);
xnor U15955 (N_15955,N_14291,N_14485);
nand U15956 (N_15956,N_14184,N_14428);
and U15957 (N_15957,N_14589,N_14223);
xnor U15958 (N_15958,N_14449,N_14719);
xor U15959 (N_15959,N_14813,N_14652);
nor U15960 (N_15960,N_14231,N_14611);
nand U15961 (N_15961,N_14280,N_14519);
xor U15962 (N_15962,N_14390,N_14574);
xor U15963 (N_15963,N_14485,N_14738);
nand U15964 (N_15964,N_14941,N_14329);
nand U15965 (N_15965,N_14134,N_14322);
and U15966 (N_15966,N_14806,N_14357);
and U15967 (N_15967,N_14687,N_14929);
and U15968 (N_15968,N_14025,N_14471);
xnor U15969 (N_15969,N_14810,N_14261);
xnor U15970 (N_15970,N_14977,N_14014);
nand U15971 (N_15971,N_14755,N_14108);
nand U15972 (N_15972,N_14029,N_14270);
and U15973 (N_15973,N_14884,N_14304);
or U15974 (N_15974,N_14555,N_14431);
nand U15975 (N_15975,N_14125,N_14520);
nor U15976 (N_15976,N_14327,N_14669);
and U15977 (N_15977,N_14697,N_14733);
xnor U15978 (N_15978,N_14699,N_14745);
xor U15979 (N_15979,N_14862,N_14352);
or U15980 (N_15980,N_14394,N_14061);
nand U15981 (N_15981,N_14245,N_14259);
or U15982 (N_15982,N_14078,N_14447);
xnor U15983 (N_15983,N_14052,N_14134);
nor U15984 (N_15984,N_14722,N_14404);
nand U15985 (N_15985,N_14378,N_14652);
xor U15986 (N_15986,N_14216,N_14798);
xnor U15987 (N_15987,N_14713,N_14284);
nor U15988 (N_15988,N_14637,N_14979);
nor U15989 (N_15989,N_14291,N_14714);
nor U15990 (N_15990,N_14298,N_14945);
and U15991 (N_15991,N_14571,N_14708);
or U15992 (N_15992,N_14728,N_14743);
nand U15993 (N_15993,N_14340,N_14863);
and U15994 (N_15994,N_14420,N_14595);
nor U15995 (N_15995,N_14725,N_14548);
xnor U15996 (N_15996,N_14238,N_14083);
and U15997 (N_15997,N_14530,N_14438);
and U15998 (N_15998,N_14303,N_14698);
or U15999 (N_15999,N_14556,N_14029);
or U16000 (N_16000,N_15331,N_15463);
or U16001 (N_16001,N_15244,N_15202);
nor U16002 (N_16002,N_15896,N_15062);
nor U16003 (N_16003,N_15689,N_15630);
nor U16004 (N_16004,N_15852,N_15232);
or U16005 (N_16005,N_15453,N_15544);
nand U16006 (N_16006,N_15631,N_15478);
xor U16007 (N_16007,N_15441,N_15785);
nand U16008 (N_16008,N_15077,N_15530);
or U16009 (N_16009,N_15097,N_15435);
and U16010 (N_16010,N_15117,N_15508);
xnor U16011 (N_16011,N_15114,N_15138);
nand U16012 (N_16012,N_15765,N_15854);
nand U16013 (N_16013,N_15172,N_15588);
nand U16014 (N_16014,N_15068,N_15764);
or U16015 (N_16015,N_15294,N_15434);
and U16016 (N_16016,N_15247,N_15812);
nor U16017 (N_16017,N_15953,N_15798);
nand U16018 (N_16018,N_15072,N_15430);
nor U16019 (N_16019,N_15086,N_15352);
nor U16020 (N_16020,N_15939,N_15165);
or U16021 (N_16021,N_15404,N_15370);
and U16022 (N_16022,N_15106,N_15877);
nor U16023 (N_16023,N_15504,N_15512);
or U16024 (N_16024,N_15205,N_15959);
nor U16025 (N_16025,N_15449,N_15047);
and U16026 (N_16026,N_15201,N_15026);
and U16027 (N_16027,N_15310,N_15168);
nand U16028 (N_16028,N_15250,N_15350);
nor U16029 (N_16029,N_15087,N_15966);
xor U16030 (N_16030,N_15088,N_15417);
and U16031 (N_16031,N_15917,N_15273);
and U16032 (N_16032,N_15075,N_15558);
nand U16033 (N_16033,N_15412,N_15292);
nand U16034 (N_16034,N_15708,N_15687);
and U16035 (N_16035,N_15634,N_15519);
nand U16036 (N_16036,N_15030,N_15091);
and U16037 (N_16037,N_15345,N_15112);
xor U16038 (N_16038,N_15291,N_15614);
and U16039 (N_16039,N_15079,N_15586);
xor U16040 (N_16040,N_15636,N_15500);
xor U16041 (N_16041,N_15926,N_15699);
nand U16042 (N_16042,N_15318,N_15050);
nand U16043 (N_16043,N_15471,N_15469);
and U16044 (N_16044,N_15141,N_15899);
nor U16045 (N_16045,N_15024,N_15568);
xor U16046 (N_16046,N_15431,N_15730);
or U16047 (N_16047,N_15938,N_15195);
and U16048 (N_16048,N_15637,N_15391);
or U16049 (N_16049,N_15652,N_15304);
xnor U16050 (N_16050,N_15888,N_15272);
nand U16051 (N_16051,N_15628,N_15314);
xor U16052 (N_16052,N_15143,N_15805);
nor U16053 (N_16053,N_15376,N_15120);
and U16054 (N_16054,N_15189,N_15045);
nor U16055 (N_16055,N_15616,N_15243);
nor U16056 (N_16056,N_15155,N_15535);
xor U16057 (N_16057,N_15006,N_15549);
xnor U16058 (N_16058,N_15793,N_15581);
and U16059 (N_16059,N_15306,N_15380);
nand U16060 (N_16060,N_15862,N_15505);
or U16061 (N_16061,N_15332,N_15646);
nor U16062 (N_16062,N_15697,N_15335);
nor U16063 (N_16063,N_15199,N_15761);
or U16064 (N_16064,N_15194,N_15690);
nor U16065 (N_16065,N_15948,N_15661);
nor U16066 (N_16066,N_15161,N_15957);
xnor U16067 (N_16067,N_15437,N_15109);
or U16068 (N_16068,N_15067,N_15758);
nor U16069 (N_16069,N_15947,N_15691);
nand U16070 (N_16070,N_15514,N_15386);
nand U16071 (N_16071,N_15935,N_15280);
xnor U16072 (N_16072,N_15063,N_15105);
and U16073 (N_16073,N_15559,N_15692);
and U16074 (N_16074,N_15988,N_15032);
nand U16075 (N_16075,N_15498,N_15246);
xor U16076 (N_16076,N_15492,N_15647);
or U16077 (N_16077,N_15864,N_15756);
and U16078 (N_16078,N_15290,N_15902);
and U16079 (N_16079,N_15015,N_15179);
and U16080 (N_16080,N_15719,N_15170);
nand U16081 (N_16081,N_15837,N_15010);
and U16082 (N_16082,N_15943,N_15574);
nor U16083 (N_16083,N_15074,N_15260);
nor U16084 (N_16084,N_15287,N_15525);
xor U16085 (N_16085,N_15094,N_15059);
or U16086 (N_16086,N_15499,N_15459);
nor U16087 (N_16087,N_15672,N_15510);
nand U16088 (N_16088,N_15124,N_15983);
nand U16089 (N_16089,N_15562,N_15491);
and U16090 (N_16090,N_15619,N_15592);
and U16091 (N_16091,N_15967,N_15375);
xor U16092 (N_16092,N_15208,N_15455);
nand U16093 (N_16093,N_15893,N_15324);
and U16094 (N_16094,N_15956,N_15134);
and U16095 (N_16095,N_15041,N_15996);
and U16096 (N_16096,N_15819,N_15999);
and U16097 (N_16097,N_15946,N_15178);
xor U16098 (N_16098,N_15762,N_15142);
and U16099 (N_16099,N_15799,N_15266);
xor U16100 (N_16100,N_15958,N_15664);
nand U16101 (N_16101,N_15704,N_15490);
or U16102 (N_16102,N_15796,N_15012);
xnor U16103 (N_16103,N_15278,N_15150);
nor U16104 (N_16104,N_15497,N_15144);
or U16105 (N_16105,N_15728,N_15828);
nor U16106 (N_16106,N_15644,N_15415);
and U16107 (N_16107,N_15995,N_15108);
nor U16108 (N_16108,N_15919,N_15521);
nor U16109 (N_16109,N_15627,N_15301);
or U16110 (N_16110,N_15347,N_15025);
and U16111 (N_16111,N_15356,N_15641);
nand U16112 (N_16112,N_15746,N_15842);
nor U16113 (N_16113,N_15531,N_15334);
xnor U16114 (N_16114,N_15416,N_15556);
and U16115 (N_16115,N_15394,N_15209);
nand U16116 (N_16116,N_15850,N_15901);
xnor U16117 (N_16117,N_15683,N_15659);
and U16118 (N_16118,N_15925,N_15210);
xor U16119 (N_16119,N_15892,N_15387);
or U16120 (N_16120,N_15049,N_15863);
nor U16121 (N_16121,N_15669,N_15311);
nand U16122 (N_16122,N_15501,N_15613);
nand U16123 (N_16123,N_15537,N_15685);
xor U16124 (N_16124,N_15298,N_15033);
xnor U16125 (N_16125,N_15714,N_15251);
xnor U16126 (N_16126,N_15259,N_15022);
and U16127 (N_16127,N_15567,N_15662);
and U16128 (N_16128,N_15240,N_15547);
nand U16129 (N_16129,N_15281,N_15268);
or U16130 (N_16130,N_15060,N_15555);
and U16131 (N_16131,N_15952,N_15136);
nand U16132 (N_16132,N_15233,N_15320);
nor U16133 (N_16133,N_15912,N_15972);
or U16134 (N_16134,N_15526,N_15101);
nand U16135 (N_16135,N_15121,N_15517);
nor U16136 (N_16136,N_15890,N_15548);
xnor U16137 (N_16137,N_15020,N_15763);
and U16138 (N_16138,N_15865,N_15949);
nor U16139 (N_16139,N_15698,N_15879);
xor U16140 (N_16140,N_15781,N_15187);
xnor U16141 (N_16141,N_15932,N_15682);
and U16142 (N_16142,N_15656,N_15225);
xor U16143 (N_16143,N_15388,N_15696);
xnor U16144 (N_16144,N_15721,N_15610);
nand U16145 (N_16145,N_15891,N_15913);
and U16146 (N_16146,N_15566,N_15701);
nand U16147 (N_16147,N_15014,N_15818);
nor U16148 (N_16148,N_15263,N_15667);
nand U16149 (N_16149,N_15889,N_15365);
or U16150 (N_16150,N_15061,N_15909);
or U16151 (N_16151,N_15856,N_15846);
or U16152 (N_16152,N_15339,N_15718);
and U16153 (N_16153,N_15288,N_15680);
or U16154 (N_16154,N_15894,N_15817);
or U16155 (N_16155,N_15978,N_15171);
nor U16156 (N_16156,N_15137,N_15571);
nand U16157 (N_16157,N_15466,N_15078);
nand U16158 (N_16158,N_15295,N_15600);
and U16159 (N_16159,N_15231,N_15176);
xnor U16160 (N_16160,N_15082,N_15220);
and U16161 (N_16161,N_15706,N_15942);
nand U16162 (N_16162,N_15822,N_15729);
and U16163 (N_16163,N_15315,N_15148);
and U16164 (N_16164,N_15465,N_15783);
nor U16165 (N_16165,N_15915,N_15399);
nand U16166 (N_16166,N_15200,N_15974);
xor U16167 (N_16167,N_15584,N_15744);
and U16168 (N_16168,N_15343,N_15612);
nor U16169 (N_16169,N_15065,N_15882);
or U16170 (N_16170,N_15599,N_15057);
xnor U16171 (N_16171,N_15874,N_15971);
xor U16172 (N_16172,N_15895,N_15792);
nand U16173 (N_16173,N_15360,N_15164);
nand U16174 (N_16174,N_15820,N_15325);
and U16175 (N_16175,N_15808,N_15007);
or U16176 (N_16176,N_15257,N_15414);
xor U16177 (N_16177,N_15594,N_15759);
xor U16178 (N_16178,N_15085,N_15342);
nand U16179 (N_16179,N_15480,N_15830);
or U16180 (N_16180,N_15645,N_15810);
or U16181 (N_16181,N_15354,N_15736);
and U16182 (N_16182,N_15866,N_15069);
nor U16183 (N_16183,N_15751,N_15994);
nor U16184 (N_16184,N_15507,N_15277);
and U16185 (N_16185,N_15963,N_15162);
or U16186 (N_16186,N_15363,N_15224);
nand U16187 (N_16187,N_15330,N_15541);
nor U16188 (N_16188,N_15193,N_15760);
nand U16189 (N_16189,N_15169,N_15782);
nand U16190 (N_16190,N_15346,N_15596);
or U16191 (N_16191,N_15139,N_15831);
xor U16192 (N_16192,N_15409,N_15274);
xnor U16193 (N_16193,N_15475,N_15623);
or U16194 (N_16194,N_15906,N_15990);
xor U16195 (N_16195,N_15707,N_15791);
and U16196 (N_16196,N_15089,N_15326);
or U16197 (N_16197,N_15035,N_15255);
nor U16198 (N_16198,N_15769,N_15132);
nand U16199 (N_16199,N_15073,N_15099);
nand U16200 (N_16200,N_15445,N_15369);
and U16201 (N_16201,N_15029,N_15262);
or U16202 (N_16202,N_15472,N_15424);
and U16203 (N_16203,N_15361,N_15931);
nor U16204 (N_16204,N_15486,N_15561);
nand U16205 (N_16205,N_15159,N_15017);
or U16206 (N_16206,N_15423,N_15309);
nor U16207 (N_16207,N_15368,N_15591);
xor U16208 (N_16208,N_15192,N_15040);
xor U16209 (N_16209,N_15384,N_15100);
and U16210 (N_16210,N_15621,N_15235);
or U16211 (N_16211,N_15524,N_15536);
xnor U16212 (N_16212,N_15390,N_15838);
nand U16213 (N_16213,N_15476,N_15910);
nand U16214 (N_16214,N_15496,N_15989);
xnor U16215 (N_16215,N_15219,N_15845);
xnor U16216 (N_16216,N_15945,N_15520);
and U16217 (N_16217,N_15635,N_15396);
and U16218 (N_16218,N_15464,N_15671);
xor U16219 (N_16219,N_15776,N_15495);
nor U16220 (N_16220,N_15538,N_15825);
or U16221 (N_16221,N_15229,N_15844);
or U16222 (N_16222,N_15217,N_15440);
and U16223 (N_16223,N_15784,N_15154);
and U16224 (N_16224,N_15797,N_15296);
and U16225 (N_16225,N_15824,N_15484);
xor U16226 (N_16226,N_15654,N_15980);
xor U16227 (N_16227,N_15857,N_15146);
or U16228 (N_16228,N_15151,N_15651);
xnor U16229 (N_16229,N_15186,N_15611);
and U16230 (N_16230,N_15768,N_15551);
nand U16231 (N_16231,N_15589,N_15239);
and U16232 (N_16232,N_15482,N_15338);
or U16233 (N_16233,N_15420,N_15595);
nor U16234 (N_16234,N_15518,N_15407);
xor U16235 (N_16235,N_15587,N_15447);
or U16236 (N_16236,N_15833,N_15802);
and U16237 (N_16237,N_15234,N_15960);
nand U16238 (N_16238,N_15276,N_15398);
nand U16239 (N_16239,N_15815,N_15640);
nor U16240 (N_16240,N_15726,N_15673);
or U16241 (N_16241,N_15928,N_15546);
nand U16242 (N_16242,N_15305,N_15705);
nand U16243 (N_16243,N_15569,N_15403);
and U16244 (N_16244,N_15657,N_15737);
xor U16245 (N_16245,N_15848,N_15271);
xnor U16246 (N_16246,N_15908,N_15483);
or U16247 (N_16247,N_15603,N_15855);
xor U16248 (N_16248,N_15362,N_15264);
xor U16249 (N_16249,N_15488,N_15145);
nor U16250 (N_16250,N_15395,N_15754);
nand U16251 (N_16251,N_15907,N_15275);
nor U16252 (N_16252,N_15458,N_15355);
xor U16253 (N_16253,N_15577,N_15695);
and U16254 (N_16254,N_15993,N_15190);
and U16255 (N_16255,N_15160,N_15344);
nor U16256 (N_16256,N_15527,N_15900);
nand U16257 (N_16257,N_15175,N_15419);
nand U16258 (N_16258,N_15212,N_15044);
xor U16259 (N_16259,N_15740,N_15432);
or U16260 (N_16260,N_15506,N_15422);
or U16261 (N_16261,N_15557,N_15887);
and U16262 (N_16262,N_15312,N_15904);
xor U16263 (N_16263,N_15303,N_15191);
and U16264 (N_16264,N_15734,N_15027);
nor U16265 (N_16265,N_15583,N_15821);
nand U16266 (N_16266,N_15009,N_15794);
and U16267 (N_16267,N_15757,N_15789);
xor U16268 (N_16268,N_15215,N_15572);
nor U16269 (N_16269,N_15598,N_15515);
and U16270 (N_16270,N_15357,N_15321);
nand U16271 (N_16271,N_15694,N_15502);
or U16272 (N_16272,N_15031,N_15055);
xnor U16273 (N_16273,N_15371,N_15745);
xnor U16274 (N_16274,N_15803,N_15991);
or U16275 (N_16275,N_15269,N_15826);
xor U16276 (N_16276,N_15379,N_15750);
nor U16277 (N_16277,N_15147,N_15579);
and U16278 (N_16278,N_15941,N_15529);
or U16279 (N_16279,N_15649,N_15166);
or U16280 (N_16280,N_15227,N_15564);
or U16281 (N_16281,N_15602,N_15920);
nand U16282 (N_16282,N_15372,N_15878);
nor U16283 (N_16283,N_15732,N_15131);
nand U16284 (N_16284,N_15329,N_15742);
or U16285 (N_16285,N_15313,N_15336);
nand U16286 (N_16286,N_15104,N_15543);
nor U16287 (N_16287,N_15397,N_15738);
and U16288 (N_16288,N_15849,N_15092);
nand U16289 (N_16289,N_15929,N_15270);
and U16290 (N_16290,N_15328,N_15979);
xor U16291 (N_16291,N_15046,N_15934);
and U16292 (N_16292,N_15998,N_15982);
nand U16293 (N_16293,N_15575,N_15364);
nand U16294 (N_16294,N_15702,N_15681);
nand U16295 (N_16295,N_15238,N_15897);
xnor U16296 (N_16296,N_15004,N_15283);
nor U16297 (N_16297,N_15660,N_15992);
nor U16298 (N_16298,N_15113,N_15747);
or U16299 (N_16299,N_15509,N_15358);
nor U16300 (N_16300,N_15735,N_15779);
xnor U16301 (N_16301,N_15316,N_15054);
xor U16302 (N_16302,N_15684,N_15724);
nand U16303 (N_16303,N_15226,N_15157);
xnor U16304 (N_16304,N_15622,N_15237);
or U16305 (N_16305,N_15307,N_15023);
xnor U16306 (N_16306,N_15410,N_15725);
nor U16307 (N_16307,N_15021,N_15460);
nand U16308 (N_16308,N_15213,N_15133);
nor U16309 (N_16309,N_15755,N_15905);
xnor U16310 (N_16310,N_15402,N_15198);
xor U16311 (N_16311,N_15563,N_15279);
nand U16312 (N_16312,N_15840,N_15438);
and U16313 (N_16313,N_15319,N_15858);
nand U16314 (N_16314,N_15493,N_15381);
or U16315 (N_16315,N_15254,N_15038);
and U16316 (N_16316,N_15400,N_15977);
xor U16317 (N_16317,N_15052,N_15716);
nor U16318 (N_16318,N_15058,N_15985);
nor U16319 (N_16319,N_15377,N_15560);
nand U16320 (N_16320,N_15110,N_15016);
xnor U16321 (N_16321,N_15712,N_15373);
and U16322 (N_16322,N_15071,N_15473);
nand U16323 (N_16323,N_15236,N_15405);
xnor U16324 (N_16324,N_15722,N_15411);
nand U16325 (N_16325,N_15847,N_15140);
nor U16326 (N_16326,N_15617,N_15550);
and U16327 (N_16327,N_15429,N_15064);
nor U16328 (N_16328,N_15806,N_15228);
and U16329 (N_16329,N_15426,N_15267);
or U16330 (N_16330,N_15118,N_15503);
or U16331 (N_16331,N_15096,N_15851);
and U16332 (N_16332,N_15011,N_15715);
or U16333 (N_16333,N_15801,N_15090);
xnor U16334 (N_16334,N_15249,N_15048);
or U16335 (N_16335,N_15348,N_15710);
or U16336 (N_16336,N_15774,N_15658);
xnor U16337 (N_16337,N_15177,N_15670);
nor U16338 (N_16338,N_15444,N_15629);
or U16339 (N_16339,N_15965,N_15098);
nor U16340 (N_16340,N_15468,N_15300);
xnor U16341 (N_16341,N_15083,N_15446);
or U16342 (N_16342,N_15204,N_15308);
nand U16343 (N_16343,N_15911,N_15081);
xor U16344 (N_16344,N_15413,N_15688);
or U16345 (N_16345,N_15076,N_15028);
nor U16346 (N_16346,N_15353,N_15513);
and U16347 (N_16347,N_15230,N_15666);
xnor U16348 (N_16348,N_15427,N_15655);
nand U16349 (N_16349,N_15448,N_15573);
and U16350 (N_16350,N_15080,N_15258);
or U16351 (N_16351,N_15000,N_15123);
xnor U16352 (N_16352,N_15481,N_15962);
and U16353 (N_16353,N_15663,N_15727);
xor U16354 (N_16354,N_15322,N_15923);
nand U16355 (N_16355,N_15383,N_15772);
or U16356 (N_16356,N_15470,N_15184);
nor U16357 (N_16357,N_15489,N_15975);
nand U16358 (N_16358,N_15554,N_15359);
and U16359 (N_16359,N_15954,N_15608);
nand U16360 (N_16360,N_15485,N_15607);
or U16361 (N_16361,N_15771,N_15955);
or U16362 (N_16362,N_15853,N_15002);
nand U16363 (N_16363,N_15787,N_15676);
and U16364 (N_16364,N_15289,N_15317);
nor U16365 (N_16365,N_15051,N_15969);
nor U16366 (N_16366,N_15743,N_15814);
or U16367 (N_16367,N_15522,N_15418);
nand U16368 (N_16368,N_15752,N_15582);
xor U16369 (N_16369,N_15018,N_15450);
nor U16370 (N_16370,N_15731,N_15153);
nor U16371 (N_16371,N_15158,N_15927);
xor U16372 (N_16372,N_15119,N_15921);
nand U16373 (N_16373,N_15606,N_15103);
xnor U16374 (N_16374,N_15615,N_15129);
xor U16375 (N_16375,N_15378,N_15436);
xor U16376 (N_16376,N_15216,N_15881);
xnor U16377 (N_16377,N_15107,N_15968);
or U16378 (N_16378,N_15180,N_15933);
xnor U16379 (N_16379,N_15832,N_15807);
and U16380 (N_16380,N_15679,N_15461);
or U16381 (N_16381,N_15678,N_15930);
or U16382 (N_16382,N_15872,N_15540);
nor U16383 (N_16383,N_15474,N_15775);
nand U16384 (N_16384,N_15070,N_15374);
or U16385 (N_16385,N_15095,N_15674);
xor U16386 (N_16386,N_15005,N_15182);
xor U16387 (N_16387,N_15039,N_15723);
nor U16388 (N_16388,N_15811,N_15860);
nor U16389 (N_16389,N_15809,N_15053);
nand U16390 (N_16390,N_15382,N_15618);
or U16391 (N_16391,N_15116,N_15218);
nand U16392 (N_16392,N_15196,N_15570);
or U16393 (N_16393,N_15984,N_15341);
and U16394 (N_16394,N_15836,N_15185);
nand U16395 (N_16395,N_15880,N_15393);
nor U16396 (N_16396,N_15643,N_15741);
or U16397 (N_16397,N_15876,N_15261);
nor U16398 (N_16398,N_15019,N_15997);
nand U16399 (N_16399,N_15827,N_15102);
or U16400 (N_16400,N_15632,N_15425);
xor U16401 (N_16401,N_15884,N_15221);
and U16402 (N_16402,N_15633,N_15457);
nor U16403 (N_16403,N_15780,N_15585);
nor U16404 (N_16404,N_15717,N_15823);
nand U16405 (N_16405,N_15976,N_15293);
xor U16406 (N_16406,N_15340,N_15037);
or U16407 (N_16407,N_15285,N_15916);
nand U16408 (N_16408,N_15443,N_15286);
xnor U16409 (N_16409,N_15428,N_15886);
xor U16410 (N_16410,N_15337,N_15389);
nand U16411 (N_16411,N_15834,N_15392);
or U16412 (N_16412,N_15973,N_15111);
nor U16413 (N_16413,N_15668,N_15149);
nor U16414 (N_16414,N_15883,N_15944);
and U16415 (N_16415,N_15885,N_15650);
xor U16416 (N_16416,N_15003,N_15207);
nor U16417 (N_16417,N_15156,N_15349);
nand U16418 (N_16418,N_15835,N_15868);
nand U16419 (N_16419,N_15282,N_15624);
nor U16420 (N_16420,N_15421,N_15351);
nor U16421 (N_16421,N_15451,N_15511);
and U16422 (N_16422,N_15829,N_15861);
or U16423 (N_16423,N_15638,N_15626);
nand U16424 (N_16424,N_15950,N_15749);
and U16425 (N_16425,N_15914,N_15256);
or U16426 (N_16426,N_15553,N_15940);
and U16427 (N_16427,N_15043,N_15013);
xor U16428 (N_16428,N_15516,N_15008);
or U16429 (N_16429,N_15433,N_15128);
nor U16430 (N_16430,N_15800,N_15211);
nor U16431 (N_16431,N_15539,N_15733);
and U16432 (N_16432,N_15036,N_15188);
and U16433 (N_16433,N_15084,N_15248);
and U16434 (N_16434,N_15578,N_15580);
or U16435 (N_16435,N_15163,N_15001);
nand U16436 (N_16436,N_15790,N_15333);
and U16437 (N_16437,N_15323,N_15859);
and U16438 (N_16438,N_15703,N_15528);
nand U16439 (N_16439,N_15869,N_15284);
nand U16440 (N_16440,N_15675,N_15873);
nor U16441 (N_16441,N_15813,N_15843);
nand U16442 (N_16442,N_15590,N_15183);
and U16443 (N_16443,N_15214,N_15713);
and U16444 (N_16444,N_15462,N_15839);
nor U16445 (N_16445,N_15918,N_15970);
and U16446 (N_16446,N_15795,N_15816);
xnor U16447 (N_16447,N_15265,N_15302);
nand U16448 (N_16448,N_15126,N_15452);
and U16449 (N_16449,N_15456,N_15327);
nor U16450 (N_16450,N_15093,N_15903);
xor U16451 (N_16451,N_15408,N_15986);
and U16452 (N_16452,N_15253,N_15401);
and U16453 (N_16453,N_15770,N_15034);
nor U16454 (N_16454,N_15773,N_15181);
nor U16455 (N_16455,N_15297,N_15937);
nor U16456 (N_16456,N_15665,N_15066);
nand U16457 (N_16457,N_15545,N_15639);
or U16458 (N_16458,N_15597,N_15609);
nand U16459 (N_16459,N_15206,N_15642);
nor U16460 (N_16460,N_15951,N_15693);
or U16461 (N_16461,N_15961,N_15477);
xnor U16462 (N_16462,N_15936,N_15042);
xnor U16463 (N_16463,N_15922,N_15593);
nand U16464 (N_16464,N_15777,N_15924);
xor U16465 (N_16465,N_15981,N_15625);
nand U16466 (N_16466,N_15299,N_15788);
xnor U16467 (N_16467,N_15604,N_15898);
and U16468 (N_16468,N_15766,N_15601);
or U16469 (N_16469,N_15653,N_15875);
xor U16470 (N_16470,N_15174,N_15406);
and U16471 (N_16471,N_15127,N_15479);
nand U16472 (N_16472,N_15252,N_15677);
nand U16473 (N_16473,N_15454,N_15532);
or U16474 (N_16474,N_15173,N_15223);
xor U16475 (N_16475,N_15241,N_15620);
nand U16476 (N_16476,N_15686,N_15576);
nand U16477 (N_16477,N_15467,N_15130);
nand U16478 (N_16478,N_15709,N_15711);
nor U16479 (N_16479,N_15552,N_15739);
xor U16480 (N_16480,N_15542,N_15778);
nand U16481 (N_16481,N_15122,N_15366);
xnor U16482 (N_16482,N_15605,N_15786);
and U16483 (N_16483,N_15841,N_15115);
nor U16484 (N_16484,N_15867,N_15804);
nor U16485 (N_16485,N_15870,N_15767);
xor U16486 (N_16486,N_15533,N_15494);
and U16487 (N_16487,N_15565,N_15753);
nor U16488 (N_16488,N_15203,N_15648);
and U16489 (N_16489,N_15385,N_15964);
nand U16490 (N_16490,N_15720,N_15439);
and U16491 (N_16491,N_15056,N_15167);
xor U16492 (N_16492,N_15700,N_15523);
or U16493 (N_16493,N_15442,N_15534);
or U16494 (N_16494,N_15125,N_15748);
xnor U16495 (N_16495,N_15135,N_15242);
and U16496 (N_16496,N_15222,N_15245);
and U16497 (N_16497,N_15197,N_15487);
nand U16498 (N_16498,N_15367,N_15152);
nand U16499 (N_16499,N_15987,N_15871);
and U16500 (N_16500,N_15286,N_15516);
and U16501 (N_16501,N_15682,N_15522);
nor U16502 (N_16502,N_15172,N_15389);
nand U16503 (N_16503,N_15466,N_15957);
and U16504 (N_16504,N_15657,N_15829);
nand U16505 (N_16505,N_15174,N_15258);
or U16506 (N_16506,N_15570,N_15665);
xnor U16507 (N_16507,N_15326,N_15362);
nand U16508 (N_16508,N_15118,N_15497);
and U16509 (N_16509,N_15726,N_15832);
nor U16510 (N_16510,N_15918,N_15194);
and U16511 (N_16511,N_15800,N_15502);
xor U16512 (N_16512,N_15678,N_15873);
nor U16513 (N_16513,N_15578,N_15643);
nor U16514 (N_16514,N_15896,N_15834);
or U16515 (N_16515,N_15424,N_15066);
nand U16516 (N_16516,N_15693,N_15683);
and U16517 (N_16517,N_15989,N_15103);
xor U16518 (N_16518,N_15386,N_15428);
or U16519 (N_16519,N_15658,N_15765);
and U16520 (N_16520,N_15115,N_15502);
nor U16521 (N_16521,N_15263,N_15562);
and U16522 (N_16522,N_15162,N_15438);
or U16523 (N_16523,N_15750,N_15697);
xor U16524 (N_16524,N_15022,N_15162);
nor U16525 (N_16525,N_15724,N_15275);
or U16526 (N_16526,N_15613,N_15068);
xor U16527 (N_16527,N_15765,N_15246);
xor U16528 (N_16528,N_15010,N_15803);
xnor U16529 (N_16529,N_15360,N_15131);
and U16530 (N_16530,N_15505,N_15925);
nand U16531 (N_16531,N_15265,N_15003);
nand U16532 (N_16532,N_15095,N_15206);
nand U16533 (N_16533,N_15748,N_15911);
nand U16534 (N_16534,N_15752,N_15616);
and U16535 (N_16535,N_15563,N_15589);
and U16536 (N_16536,N_15012,N_15767);
or U16537 (N_16537,N_15247,N_15713);
nand U16538 (N_16538,N_15276,N_15194);
and U16539 (N_16539,N_15946,N_15926);
nand U16540 (N_16540,N_15698,N_15059);
xnor U16541 (N_16541,N_15683,N_15797);
and U16542 (N_16542,N_15109,N_15116);
nand U16543 (N_16543,N_15508,N_15456);
and U16544 (N_16544,N_15574,N_15010);
or U16545 (N_16545,N_15005,N_15520);
nor U16546 (N_16546,N_15457,N_15391);
xor U16547 (N_16547,N_15070,N_15748);
nor U16548 (N_16548,N_15604,N_15061);
and U16549 (N_16549,N_15145,N_15670);
nand U16550 (N_16550,N_15028,N_15228);
and U16551 (N_16551,N_15427,N_15408);
xnor U16552 (N_16552,N_15774,N_15831);
and U16553 (N_16553,N_15495,N_15936);
or U16554 (N_16554,N_15565,N_15650);
xnor U16555 (N_16555,N_15595,N_15384);
nand U16556 (N_16556,N_15726,N_15668);
or U16557 (N_16557,N_15706,N_15005);
or U16558 (N_16558,N_15552,N_15811);
or U16559 (N_16559,N_15926,N_15869);
nand U16560 (N_16560,N_15095,N_15684);
and U16561 (N_16561,N_15098,N_15565);
nand U16562 (N_16562,N_15975,N_15337);
nand U16563 (N_16563,N_15490,N_15887);
xor U16564 (N_16564,N_15358,N_15543);
nand U16565 (N_16565,N_15701,N_15319);
and U16566 (N_16566,N_15259,N_15612);
nand U16567 (N_16567,N_15107,N_15769);
nor U16568 (N_16568,N_15007,N_15259);
xor U16569 (N_16569,N_15225,N_15359);
nor U16570 (N_16570,N_15445,N_15480);
xnor U16571 (N_16571,N_15715,N_15626);
or U16572 (N_16572,N_15425,N_15757);
nor U16573 (N_16573,N_15277,N_15146);
nand U16574 (N_16574,N_15942,N_15818);
and U16575 (N_16575,N_15397,N_15774);
nor U16576 (N_16576,N_15835,N_15961);
xnor U16577 (N_16577,N_15221,N_15503);
nor U16578 (N_16578,N_15911,N_15812);
xnor U16579 (N_16579,N_15316,N_15193);
or U16580 (N_16580,N_15886,N_15610);
nand U16581 (N_16581,N_15867,N_15317);
xnor U16582 (N_16582,N_15003,N_15680);
nand U16583 (N_16583,N_15466,N_15496);
nor U16584 (N_16584,N_15825,N_15402);
xnor U16585 (N_16585,N_15185,N_15911);
nand U16586 (N_16586,N_15100,N_15615);
or U16587 (N_16587,N_15176,N_15521);
or U16588 (N_16588,N_15335,N_15445);
and U16589 (N_16589,N_15893,N_15881);
nor U16590 (N_16590,N_15068,N_15742);
or U16591 (N_16591,N_15192,N_15831);
xor U16592 (N_16592,N_15359,N_15787);
and U16593 (N_16593,N_15129,N_15855);
nand U16594 (N_16594,N_15348,N_15578);
xnor U16595 (N_16595,N_15052,N_15627);
or U16596 (N_16596,N_15274,N_15113);
and U16597 (N_16597,N_15136,N_15148);
xnor U16598 (N_16598,N_15126,N_15642);
or U16599 (N_16599,N_15503,N_15400);
nand U16600 (N_16600,N_15111,N_15414);
and U16601 (N_16601,N_15201,N_15257);
or U16602 (N_16602,N_15785,N_15234);
and U16603 (N_16603,N_15890,N_15956);
nand U16604 (N_16604,N_15332,N_15886);
nor U16605 (N_16605,N_15984,N_15196);
and U16606 (N_16606,N_15128,N_15527);
nand U16607 (N_16607,N_15559,N_15502);
nand U16608 (N_16608,N_15601,N_15660);
or U16609 (N_16609,N_15636,N_15134);
or U16610 (N_16610,N_15346,N_15644);
xnor U16611 (N_16611,N_15856,N_15590);
xnor U16612 (N_16612,N_15580,N_15093);
nor U16613 (N_16613,N_15250,N_15080);
nand U16614 (N_16614,N_15937,N_15687);
xnor U16615 (N_16615,N_15957,N_15078);
nor U16616 (N_16616,N_15198,N_15185);
nand U16617 (N_16617,N_15082,N_15037);
nor U16618 (N_16618,N_15503,N_15647);
xnor U16619 (N_16619,N_15738,N_15769);
xnor U16620 (N_16620,N_15413,N_15809);
xor U16621 (N_16621,N_15104,N_15330);
and U16622 (N_16622,N_15164,N_15795);
nand U16623 (N_16623,N_15345,N_15200);
nand U16624 (N_16624,N_15484,N_15751);
xor U16625 (N_16625,N_15846,N_15811);
xnor U16626 (N_16626,N_15142,N_15597);
xor U16627 (N_16627,N_15931,N_15647);
nor U16628 (N_16628,N_15138,N_15555);
xnor U16629 (N_16629,N_15965,N_15520);
nor U16630 (N_16630,N_15435,N_15511);
xor U16631 (N_16631,N_15913,N_15163);
nor U16632 (N_16632,N_15801,N_15070);
and U16633 (N_16633,N_15447,N_15153);
and U16634 (N_16634,N_15811,N_15702);
and U16635 (N_16635,N_15678,N_15004);
nor U16636 (N_16636,N_15909,N_15846);
nand U16637 (N_16637,N_15224,N_15563);
nand U16638 (N_16638,N_15857,N_15288);
or U16639 (N_16639,N_15160,N_15558);
nor U16640 (N_16640,N_15378,N_15616);
and U16641 (N_16641,N_15380,N_15500);
and U16642 (N_16642,N_15661,N_15077);
nand U16643 (N_16643,N_15769,N_15732);
or U16644 (N_16644,N_15880,N_15510);
or U16645 (N_16645,N_15196,N_15177);
nand U16646 (N_16646,N_15427,N_15996);
and U16647 (N_16647,N_15974,N_15284);
and U16648 (N_16648,N_15614,N_15423);
xnor U16649 (N_16649,N_15718,N_15620);
xor U16650 (N_16650,N_15021,N_15351);
xnor U16651 (N_16651,N_15641,N_15379);
nand U16652 (N_16652,N_15466,N_15226);
nand U16653 (N_16653,N_15682,N_15233);
and U16654 (N_16654,N_15395,N_15309);
xor U16655 (N_16655,N_15372,N_15476);
nand U16656 (N_16656,N_15999,N_15470);
and U16657 (N_16657,N_15993,N_15302);
nor U16658 (N_16658,N_15641,N_15020);
nand U16659 (N_16659,N_15338,N_15561);
or U16660 (N_16660,N_15605,N_15812);
nand U16661 (N_16661,N_15902,N_15597);
or U16662 (N_16662,N_15131,N_15019);
or U16663 (N_16663,N_15699,N_15482);
or U16664 (N_16664,N_15915,N_15948);
xnor U16665 (N_16665,N_15278,N_15476);
xnor U16666 (N_16666,N_15800,N_15463);
and U16667 (N_16667,N_15914,N_15566);
nand U16668 (N_16668,N_15209,N_15992);
or U16669 (N_16669,N_15799,N_15503);
and U16670 (N_16670,N_15045,N_15067);
nor U16671 (N_16671,N_15646,N_15075);
xor U16672 (N_16672,N_15952,N_15085);
and U16673 (N_16673,N_15871,N_15971);
and U16674 (N_16674,N_15669,N_15888);
nand U16675 (N_16675,N_15517,N_15008);
or U16676 (N_16676,N_15737,N_15510);
nor U16677 (N_16677,N_15121,N_15727);
or U16678 (N_16678,N_15655,N_15956);
or U16679 (N_16679,N_15055,N_15135);
and U16680 (N_16680,N_15784,N_15796);
or U16681 (N_16681,N_15315,N_15725);
nand U16682 (N_16682,N_15515,N_15910);
and U16683 (N_16683,N_15755,N_15056);
or U16684 (N_16684,N_15448,N_15677);
nor U16685 (N_16685,N_15789,N_15361);
xnor U16686 (N_16686,N_15610,N_15749);
xor U16687 (N_16687,N_15689,N_15927);
xor U16688 (N_16688,N_15321,N_15491);
and U16689 (N_16689,N_15257,N_15719);
and U16690 (N_16690,N_15520,N_15235);
xnor U16691 (N_16691,N_15266,N_15771);
xor U16692 (N_16692,N_15601,N_15904);
and U16693 (N_16693,N_15281,N_15190);
xor U16694 (N_16694,N_15626,N_15157);
xor U16695 (N_16695,N_15504,N_15855);
nor U16696 (N_16696,N_15178,N_15957);
or U16697 (N_16697,N_15567,N_15807);
and U16698 (N_16698,N_15216,N_15123);
xor U16699 (N_16699,N_15817,N_15790);
nor U16700 (N_16700,N_15528,N_15024);
nor U16701 (N_16701,N_15406,N_15734);
nor U16702 (N_16702,N_15424,N_15611);
nand U16703 (N_16703,N_15070,N_15282);
nand U16704 (N_16704,N_15582,N_15899);
xor U16705 (N_16705,N_15228,N_15210);
nand U16706 (N_16706,N_15617,N_15515);
and U16707 (N_16707,N_15889,N_15438);
and U16708 (N_16708,N_15534,N_15857);
or U16709 (N_16709,N_15716,N_15209);
nor U16710 (N_16710,N_15368,N_15683);
or U16711 (N_16711,N_15212,N_15346);
or U16712 (N_16712,N_15124,N_15604);
nor U16713 (N_16713,N_15482,N_15626);
nor U16714 (N_16714,N_15333,N_15005);
or U16715 (N_16715,N_15034,N_15137);
or U16716 (N_16716,N_15389,N_15286);
or U16717 (N_16717,N_15406,N_15078);
or U16718 (N_16718,N_15586,N_15362);
or U16719 (N_16719,N_15264,N_15415);
or U16720 (N_16720,N_15829,N_15776);
nor U16721 (N_16721,N_15770,N_15558);
nor U16722 (N_16722,N_15801,N_15729);
or U16723 (N_16723,N_15627,N_15862);
and U16724 (N_16724,N_15091,N_15645);
and U16725 (N_16725,N_15903,N_15786);
and U16726 (N_16726,N_15534,N_15964);
nand U16727 (N_16727,N_15665,N_15664);
or U16728 (N_16728,N_15739,N_15376);
nor U16729 (N_16729,N_15414,N_15185);
nor U16730 (N_16730,N_15100,N_15628);
or U16731 (N_16731,N_15640,N_15157);
xor U16732 (N_16732,N_15379,N_15910);
xor U16733 (N_16733,N_15241,N_15429);
xnor U16734 (N_16734,N_15921,N_15279);
nand U16735 (N_16735,N_15626,N_15738);
and U16736 (N_16736,N_15146,N_15639);
xnor U16737 (N_16737,N_15526,N_15316);
nor U16738 (N_16738,N_15616,N_15270);
xor U16739 (N_16739,N_15003,N_15136);
xor U16740 (N_16740,N_15845,N_15859);
nor U16741 (N_16741,N_15513,N_15226);
xnor U16742 (N_16742,N_15940,N_15395);
or U16743 (N_16743,N_15946,N_15293);
and U16744 (N_16744,N_15034,N_15470);
xor U16745 (N_16745,N_15933,N_15375);
nand U16746 (N_16746,N_15186,N_15196);
nand U16747 (N_16747,N_15273,N_15967);
or U16748 (N_16748,N_15066,N_15084);
nor U16749 (N_16749,N_15486,N_15302);
nand U16750 (N_16750,N_15519,N_15230);
xor U16751 (N_16751,N_15962,N_15055);
nand U16752 (N_16752,N_15158,N_15276);
or U16753 (N_16753,N_15417,N_15989);
nor U16754 (N_16754,N_15522,N_15348);
nor U16755 (N_16755,N_15789,N_15197);
nor U16756 (N_16756,N_15273,N_15816);
xor U16757 (N_16757,N_15934,N_15886);
nor U16758 (N_16758,N_15965,N_15203);
nor U16759 (N_16759,N_15309,N_15177);
or U16760 (N_16760,N_15311,N_15587);
nor U16761 (N_16761,N_15486,N_15446);
and U16762 (N_16762,N_15497,N_15405);
or U16763 (N_16763,N_15146,N_15743);
or U16764 (N_16764,N_15881,N_15196);
or U16765 (N_16765,N_15502,N_15964);
nand U16766 (N_16766,N_15099,N_15317);
nand U16767 (N_16767,N_15046,N_15616);
and U16768 (N_16768,N_15406,N_15182);
or U16769 (N_16769,N_15496,N_15654);
and U16770 (N_16770,N_15794,N_15376);
xor U16771 (N_16771,N_15129,N_15887);
xor U16772 (N_16772,N_15964,N_15549);
or U16773 (N_16773,N_15125,N_15071);
xnor U16774 (N_16774,N_15160,N_15787);
and U16775 (N_16775,N_15101,N_15218);
or U16776 (N_16776,N_15401,N_15432);
and U16777 (N_16777,N_15199,N_15714);
nor U16778 (N_16778,N_15648,N_15711);
xnor U16779 (N_16779,N_15131,N_15469);
xor U16780 (N_16780,N_15816,N_15149);
and U16781 (N_16781,N_15814,N_15225);
and U16782 (N_16782,N_15110,N_15827);
and U16783 (N_16783,N_15741,N_15932);
nor U16784 (N_16784,N_15281,N_15186);
xnor U16785 (N_16785,N_15467,N_15013);
nand U16786 (N_16786,N_15346,N_15827);
or U16787 (N_16787,N_15721,N_15107);
and U16788 (N_16788,N_15053,N_15891);
and U16789 (N_16789,N_15576,N_15455);
or U16790 (N_16790,N_15162,N_15073);
or U16791 (N_16791,N_15385,N_15478);
xnor U16792 (N_16792,N_15581,N_15246);
xnor U16793 (N_16793,N_15879,N_15976);
and U16794 (N_16794,N_15658,N_15541);
and U16795 (N_16795,N_15316,N_15237);
and U16796 (N_16796,N_15979,N_15827);
nand U16797 (N_16797,N_15844,N_15102);
xor U16798 (N_16798,N_15427,N_15899);
xor U16799 (N_16799,N_15490,N_15776);
or U16800 (N_16800,N_15947,N_15226);
or U16801 (N_16801,N_15155,N_15269);
or U16802 (N_16802,N_15060,N_15307);
and U16803 (N_16803,N_15491,N_15990);
and U16804 (N_16804,N_15480,N_15208);
or U16805 (N_16805,N_15170,N_15020);
nand U16806 (N_16806,N_15302,N_15389);
and U16807 (N_16807,N_15879,N_15936);
nor U16808 (N_16808,N_15985,N_15956);
nor U16809 (N_16809,N_15191,N_15742);
nand U16810 (N_16810,N_15882,N_15181);
xor U16811 (N_16811,N_15898,N_15951);
nor U16812 (N_16812,N_15335,N_15931);
and U16813 (N_16813,N_15413,N_15443);
and U16814 (N_16814,N_15617,N_15764);
nor U16815 (N_16815,N_15681,N_15592);
and U16816 (N_16816,N_15959,N_15399);
and U16817 (N_16817,N_15579,N_15259);
or U16818 (N_16818,N_15996,N_15391);
nor U16819 (N_16819,N_15256,N_15105);
or U16820 (N_16820,N_15818,N_15896);
and U16821 (N_16821,N_15832,N_15579);
xor U16822 (N_16822,N_15726,N_15579);
and U16823 (N_16823,N_15070,N_15845);
nand U16824 (N_16824,N_15389,N_15912);
or U16825 (N_16825,N_15960,N_15728);
or U16826 (N_16826,N_15324,N_15013);
or U16827 (N_16827,N_15114,N_15403);
or U16828 (N_16828,N_15662,N_15998);
and U16829 (N_16829,N_15806,N_15525);
or U16830 (N_16830,N_15664,N_15456);
or U16831 (N_16831,N_15216,N_15648);
xnor U16832 (N_16832,N_15744,N_15761);
and U16833 (N_16833,N_15123,N_15135);
nand U16834 (N_16834,N_15911,N_15871);
nand U16835 (N_16835,N_15579,N_15975);
or U16836 (N_16836,N_15501,N_15519);
and U16837 (N_16837,N_15750,N_15503);
nand U16838 (N_16838,N_15900,N_15040);
xor U16839 (N_16839,N_15806,N_15135);
xnor U16840 (N_16840,N_15366,N_15985);
nor U16841 (N_16841,N_15658,N_15125);
nor U16842 (N_16842,N_15891,N_15336);
nor U16843 (N_16843,N_15332,N_15193);
xor U16844 (N_16844,N_15847,N_15815);
xor U16845 (N_16845,N_15606,N_15526);
or U16846 (N_16846,N_15007,N_15290);
nor U16847 (N_16847,N_15312,N_15577);
or U16848 (N_16848,N_15047,N_15792);
nor U16849 (N_16849,N_15253,N_15357);
xor U16850 (N_16850,N_15316,N_15445);
nor U16851 (N_16851,N_15471,N_15833);
xor U16852 (N_16852,N_15616,N_15775);
and U16853 (N_16853,N_15318,N_15480);
or U16854 (N_16854,N_15213,N_15076);
or U16855 (N_16855,N_15138,N_15021);
and U16856 (N_16856,N_15651,N_15210);
and U16857 (N_16857,N_15808,N_15543);
nor U16858 (N_16858,N_15332,N_15255);
xnor U16859 (N_16859,N_15924,N_15211);
or U16860 (N_16860,N_15877,N_15495);
xor U16861 (N_16861,N_15380,N_15059);
nor U16862 (N_16862,N_15609,N_15409);
and U16863 (N_16863,N_15611,N_15252);
xnor U16864 (N_16864,N_15586,N_15051);
nand U16865 (N_16865,N_15691,N_15942);
or U16866 (N_16866,N_15784,N_15320);
nand U16867 (N_16867,N_15829,N_15600);
and U16868 (N_16868,N_15279,N_15035);
nor U16869 (N_16869,N_15322,N_15914);
and U16870 (N_16870,N_15457,N_15498);
nor U16871 (N_16871,N_15455,N_15359);
nand U16872 (N_16872,N_15968,N_15706);
or U16873 (N_16873,N_15900,N_15622);
nand U16874 (N_16874,N_15428,N_15336);
xnor U16875 (N_16875,N_15058,N_15627);
or U16876 (N_16876,N_15599,N_15090);
and U16877 (N_16877,N_15065,N_15029);
xnor U16878 (N_16878,N_15692,N_15023);
xnor U16879 (N_16879,N_15637,N_15611);
and U16880 (N_16880,N_15038,N_15994);
nand U16881 (N_16881,N_15965,N_15087);
nand U16882 (N_16882,N_15996,N_15889);
nand U16883 (N_16883,N_15208,N_15046);
or U16884 (N_16884,N_15881,N_15844);
nand U16885 (N_16885,N_15132,N_15397);
nand U16886 (N_16886,N_15553,N_15165);
nand U16887 (N_16887,N_15199,N_15788);
xnor U16888 (N_16888,N_15690,N_15265);
nor U16889 (N_16889,N_15207,N_15820);
or U16890 (N_16890,N_15034,N_15105);
xnor U16891 (N_16891,N_15073,N_15910);
nor U16892 (N_16892,N_15021,N_15633);
and U16893 (N_16893,N_15611,N_15098);
nand U16894 (N_16894,N_15099,N_15218);
xnor U16895 (N_16895,N_15633,N_15400);
nor U16896 (N_16896,N_15955,N_15234);
xor U16897 (N_16897,N_15996,N_15420);
and U16898 (N_16898,N_15809,N_15208);
or U16899 (N_16899,N_15437,N_15653);
or U16900 (N_16900,N_15218,N_15604);
nand U16901 (N_16901,N_15618,N_15989);
xnor U16902 (N_16902,N_15283,N_15961);
nand U16903 (N_16903,N_15829,N_15726);
and U16904 (N_16904,N_15789,N_15441);
or U16905 (N_16905,N_15414,N_15402);
and U16906 (N_16906,N_15729,N_15868);
xor U16907 (N_16907,N_15332,N_15965);
nor U16908 (N_16908,N_15018,N_15573);
and U16909 (N_16909,N_15041,N_15588);
nand U16910 (N_16910,N_15227,N_15403);
and U16911 (N_16911,N_15961,N_15797);
and U16912 (N_16912,N_15749,N_15757);
and U16913 (N_16913,N_15119,N_15270);
or U16914 (N_16914,N_15088,N_15629);
xor U16915 (N_16915,N_15441,N_15591);
or U16916 (N_16916,N_15618,N_15548);
nor U16917 (N_16917,N_15793,N_15184);
or U16918 (N_16918,N_15489,N_15494);
xor U16919 (N_16919,N_15275,N_15098);
and U16920 (N_16920,N_15761,N_15958);
and U16921 (N_16921,N_15014,N_15138);
and U16922 (N_16922,N_15094,N_15198);
and U16923 (N_16923,N_15341,N_15506);
and U16924 (N_16924,N_15059,N_15835);
nand U16925 (N_16925,N_15762,N_15930);
nand U16926 (N_16926,N_15190,N_15888);
or U16927 (N_16927,N_15298,N_15042);
nand U16928 (N_16928,N_15473,N_15744);
xnor U16929 (N_16929,N_15702,N_15318);
xor U16930 (N_16930,N_15672,N_15853);
xor U16931 (N_16931,N_15409,N_15222);
nor U16932 (N_16932,N_15135,N_15870);
xnor U16933 (N_16933,N_15382,N_15987);
xor U16934 (N_16934,N_15404,N_15162);
and U16935 (N_16935,N_15876,N_15490);
nand U16936 (N_16936,N_15264,N_15142);
and U16937 (N_16937,N_15273,N_15207);
and U16938 (N_16938,N_15299,N_15682);
xor U16939 (N_16939,N_15600,N_15724);
nand U16940 (N_16940,N_15610,N_15342);
xnor U16941 (N_16941,N_15727,N_15599);
nor U16942 (N_16942,N_15721,N_15823);
nor U16943 (N_16943,N_15094,N_15778);
nand U16944 (N_16944,N_15471,N_15422);
and U16945 (N_16945,N_15638,N_15192);
or U16946 (N_16946,N_15140,N_15855);
nand U16947 (N_16947,N_15199,N_15557);
xor U16948 (N_16948,N_15306,N_15202);
nor U16949 (N_16949,N_15133,N_15073);
nand U16950 (N_16950,N_15475,N_15717);
xnor U16951 (N_16951,N_15968,N_15320);
xor U16952 (N_16952,N_15070,N_15923);
or U16953 (N_16953,N_15007,N_15151);
nand U16954 (N_16954,N_15773,N_15628);
and U16955 (N_16955,N_15542,N_15230);
or U16956 (N_16956,N_15484,N_15913);
nand U16957 (N_16957,N_15577,N_15863);
and U16958 (N_16958,N_15549,N_15627);
nand U16959 (N_16959,N_15087,N_15185);
nand U16960 (N_16960,N_15789,N_15702);
xnor U16961 (N_16961,N_15318,N_15550);
nand U16962 (N_16962,N_15173,N_15058);
or U16963 (N_16963,N_15251,N_15754);
and U16964 (N_16964,N_15417,N_15219);
or U16965 (N_16965,N_15720,N_15789);
xor U16966 (N_16966,N_15396,N_15231);
and U16967 (N_16967,N_15381,N_15247);
nand U16968 (N_16968,N_15592,N_15370);
and U16969 (N_16969,N_15640,N_15588);
and U16970 (N_16970,N_15173,N_15782);
nand U16971 (N_16971,N_15506,N_15026);
nand U16972 (N_16972,N_15654,N_15450);
nor U16973 (N_16973,N_15211,N_15898);
and U16974 (N_16974,N_15240,N_15878);
or U16975 (N_16975,N_15148,N_15468);
nand U16976 (N_16976,N_15579,N_15487);
and U16977 (N_16977,N_15692,N_15194);
nand U16978 (N_16978,N_15539,N_15848);
nand U16979 (N_16979,N_15750,N_15045);
or U16980 (N_16980,N_15334,N_15045);
nand U16981 (N_16981,N_15806,N_15460);
or U16982 (N_16982,N_15110,N_15000);
nand U16983 (N_16983,N_15935,N_15812);
and U16984 (N_16984,N_15450,N_15318);
and U16985 (N_16985,N_15223,N_15126);
nand U16986 (N_16986,N_15897,N_15600);
xnor U16987 (N_16987,N_15030,N_15579);
and U16988 (N_16988,N_15384,N_15008);
or U16989 (N_16989,N_15980,N_15072);
nor U16990 (N_16990,N_15091,N_15830);
or U16991 (N_16991,N_15258,N_15901);
and U16992 (N_16992,N_15834,N_15625);
and U16993 (N_16993,N_15604,N_15053);
xnor U16994 (N_16994,N_15349,N_15069);
and U16995 (N_16995,N_15093,N_15882);
and U16996 (N_16996,N_15961,N_15026);
nor U16997 (N_16997,N_15529,N_15624);
or U16998 (N_16998,N_15371,N_15484);
nand U16999 (N_16999,N_15211,N_15252);
and U17000 (N_17000,N_16022,N_16459);
and U17001 (N_17001,N_16398,N_16091);
nand U17002 (N_17002,N_16178,N_16656);
or U17003 (N_17003,N_16793,N_16057);
or U17004 (N_17004,N_16208,N_16150);
xor U17005 (N_17005,N_16577,N_16330);
or U17006 (N_17006,N_16152,N_16565);
nand U17007 (N_17007,N_16781,N_16928);
or U17008 (N_17008,N_16002,N_16950);
nand U17009 (N_17009,N_16893,N_16762);
and U17010 (N_17010,N_16641,N_16308);
nand U17011 (N_17011,N_16069,N_16340);
nor U17012 (N_17012,N_16855,N_16881);
nand U17013 (N_17013,N_16320,N_16257);
and U17014 (N_17014,N_16958,N_16275);
or U17015 (N_17015,N_16559,N_16860);
or U17016 (N_17016,N_16366,N_16765);
nor U17017 (N_17017,N_16584,N_16688);
nand U17018 (N_17018,N_16965,N_16934);
xnor U17019 (N_17019,N_16072,N_16725);
nand U17020 (N_17020,N_16792,N_16117);
xor U17021 (N_17021,N_16906,N_16021);
nand U17022 (N_17022,N_16768,N_16795);
xnor U17023 (N_17023,N_16583,N_16966);
and U17024 (N_17024,N_16419,N_16972);
nor U17025 (N_17025,N_16227,N_16301);
or U17026 (N_17026,N_16046,N_16411);
xnor U17027 (N_17027,N_16242,N_16267);
or U17028 (N_17028,N_16809,N_16240);
or U17029 (N_17029,N_16335,N_16367);
xor U17030 (N_17030,N_16035,N_16075);
or U17031 (N_17031,N_16593,N_16438);
nor U17032 (N_17032,N_16226,N_16957);
or U17033 (N_17033,N_16704,N_16735);
nor U17034 (N_17034,N_16286,N_16806);
or U17035 (N_17035,N_16328,N_16917);
or U17036 (N_17036,N_16192,N_16219);
xnor U17037 (N_17037,N_16554,N_16104);
nor U17038 (N_17038,N_16751,N_16200);
or U17039 (N_17039,N_16359,N_16517);
nor U17040 (N_17040,N_16682,N_16107);
or U17041 (N_17041,N_16140,N_16414);
nand U17042 (N_17042,N_16382,N_16142);
and U17043 (N_17043,N_16610,N_16803);
nor U17044 (N_17044,N_16537,N_16757);
and U17045 (N_17045,N_16500,N_16499);
nand U17046 (N_17046,N_16829,N_16456);
or U17047 (N_17047,N_16785,N_16455);
and U17048 (N_17048,N_16428,N_16826);
nor U17049 (N_17049,N_16759,N_16827);
or U17050 (N_17050,N_16348,N_16418);
and U17051 (N_17051,N_16945,N_16217);
xnor U17052 (N_17052,N_16259,N_16523);
nand U17053 (N_17053,N_16319,N_16129);
nand U17054 (N_17054,N_16712,N_16442);
or U17055 (N_17055,N_16939,N_16655);
nor U17056 (N_17056,N_16321,N_16106);
and U17057 (N_17057,N_16221,N_16253);
and U17058 (N_17058,N_16215,N_16049);
nand U17059 (N_17059,N_16872,N_16201);
nand U17060 (N_17060,N_16730,N_16982);
nor U17061 (N_17061,N_16099,N_16944);
or U17062 (N_17062,N_16908,N_16369);
or U17063 (N_17063,N_16051,N_16303);
xor U17064 (N_17064,N_16202,N_16068);
nand U17065 (N_17065,N_16805,N_16334);
or U17066 (N_17066,N_16003,N_16044);
or U17067 (N_17067,N_16963,N_16123);
and U17068 (N_17068,N_16596,N_16941);
and U17069 (N_17069,N_16420,N_16771);
xnor U17070 (N_17070,N_16005,N_16125);
xor U17071 (N_17071,N_16946,N_16225);
nor U17072 (N_17072,N_16643,N_16845);
and U17073 (N_17073,N_16535,N_16862);
xnor U17074 (N_17074,N_16276,N_16155);
xor U17075 (N_17075,N_16479,N_16601);
nor U17076 (N_17076,N_16790,N_16495);
or U17077 (N_17077,N_16362,N_16973);
nor U17078 (N_17078,N_16783,N_16964);
and U17079 (N_17079,N_16191,N_16160);
xnor U17080 (N_17080,N_16011,N_16992);
nand U17081 (N_17081,N_16676,N_16617);
xor U17082 (N_17082,N_16938,N_16065);
nand U17083 (N_17083,N_16530,N_16450);
xor U17084 (N_17084,N_16498,N_16100);
nor U17085 (N_17085,N_16731,N_16912);
xnor U17086 (N_17086,N_16871,N_16029);
nor U17087 (N_17087,N_16415,N_16548);
or U17088 (N_17088,N_16623,N_16087);
nor U17089 (N_17089,N_16451,N_16391);
nand U17090 (N_17090,N_16076,N_16258);
and U17091 (N_17091,N_16262,N_16932);
or U17092 (N_17092,N_16841,N_16284);
nor U17093 (N_17093,N_16167,N_16977);
nor U17094 (N_17094,N_16055,N_16830);
or U17095 (N_17095,N_16914,N_16590);
or U17096 (N_17096,N_16810,N_16098);
xor U17097 (N_17097,N_16338,N_16612);
or U17098 (N_17098,N_16635,N_16361);
xnor U17099 (N_17099,N_16605,N_16477);
or U17100 (N_17100,N_16628,N_16653);
or U17101 (N_17101,N_16396,N_16542);
nand U17102 (N_17102,N_16431,N_16968);
xor U17103 (N_17103,N_16042,N_16880);
nor U17104 (N_17104,N_16313,N_16863);
or U17105 (N_17105,N_16980,N_16251);
xnor U17106 (N_17106,N_16004,N_16329);
xor U17107 (N_17107,N_16758,N_16859);
or U17108 (N_17108,N_16085,N_16324);
nor U17109 (N_17109,N_16948,N_16888);
xnor U17110 (N_17110,N_16408,N_16169);
and U17111 (N_17111,N_16036,N_16198);
nand U17112 (N_17112,N_16525,N_16911);
or U17113 (N_17113,N_16587,N_16344);
nor U17114 (N_17114,N_16170,N_16470);
nor U17115 (N_17115,N_16270,N_16309);
and U17116 (N_17116,N_16481,N_16176);
nand U17117 (N_17117,N_16818,N_16209);
or U17118 (N_17118,N_16831,N_16996);
xnor U17119 (N_17119,N_16607,N_16505);
nand U17120 (N_17120,N_16678,N_16705);
nor U17121 (N_17121,N_16734,N_16307);
nand U17122 (N_17122,N_16311,N_16819);
nand U17123 (N_17123,N_16846,N_16960);
nor U17124 (N_17124,N_16564,N_16484);
or U17125 (N_17125,N_16926,N_16386);
nand U17126 (N_17126,N_16502,N_16063);
xor U17127 (N_17127,N_16814,N_16918);
or U17128 (N_17128,N_16374,N_16626);
nand U17129 (N_17129,N_16794,N_16896);
nand U17130 (N_17130,N_16546,N_16598);
xnor U17131 (N_17131,N_16526,N_16475);
nor U17132 (N_17132,N_16220,N_16280);
xnor U17133 (N_17133,N_16388,N_16037);
xnor U17134 (N_17134,N_16218,N_16715);
nor U17135 (N_17135,N_16951,N_16817);
and U17136 (N_17136,N_16824,N_16649);
nand U17137 (N_17137,N_16812,N_16245);
nor U17138 (N_17138,N_16567,N_16358);
and U17139 (N_17139,N_16317,N_16323);
or U17140 (N_17140,N_16569,N_16058);
xor U17141 (N_17141,N_16522,N_16365);
xor U17142 (N_17142,N_16184,N_16861);
or U17143 (N_17143,N_16562,N_16211);
nand U17144 (N_17144,N_16416,N_16853);
nand U17145 (N_17145,N_16639,N_16447);
or U17146 (N_17146,N_16122,N_16999);
and U17147 (N_17147,N_16385,N_16113);
nand U17148 (N_17148,N_16784,N_16102);
nor U17149 (N_17149,N_16620,N_16297);
nand U17150 (N_17150,N_16978,N_16985);
nor U17151 (N_17151,N_16744,N_16835);
and U17152 (N_17152,N_16677,N_16133);
xnor U17153 (N_17153,N_16417,N_16693);
nand U17154 (N_17154,N_16707,N_16402);
or U17155 (N_17155,N_16264,N_16648);
nor U17156 (N_17156,N_16709,N_16984);
nand U17157 (N_17157,N_16165,N_16609);
nor U17158 (N_17158,N_16356,N_16745);
nand U17159 (N_17159,N_16302,N_16886);
nor U17160 (N_17160,N_16347,N_16663);
nor U17161 (N_17161,N_16574,N_16173);
xor U17162 (N_17162,N_16971,N_16718);
nand U17163 (N_17163,N_16357,N_16599);
xnor U17164 (N_17164,N_16904,N_16064);
xor U17165 (N_17165,N_16190,N_16728);
xnor U17166 (N_17166,N_16540,N_16713);
nor U17167 (N_17167,N_16448,N_16273);
nor U17168 (N_17168,N_16698,N_16746);
and U17169 (N_17169,N_16995,N_16921);
xor U17170 (N_17170,N_16332,N_16719);
xor U17171 (N_17171,N_16060,N_16683);
xor U17172 (N_17172,N_16723,N_16882);
xor U17173 (N_17173,N_16848,N_16364);
and U17174 (N_17174,N_16508,N_16993);
nor U17175 (N_17175,N_16778,N_16796);
nor U17176 (N_17176,N_16486,N_16798);
and U17177 (N_17177,N_16128,N_16674);
or U17178 (N_17178,N_16389,N_16494);
nor U17179 (N_17179,N_16252,N_16149);
xor U17180 (N_17180,N_16487,N_16788);
or U17181 (N_17181,N_16014,N_16851);
xnor U17182 (N_17182,N_16124,N_16062);
and U17183 (N_17183,N_16488,N_16392);
nor U17184 (N_17184,N_16084,N_16134);
or U17185 (N_17185,N_16491,N_16018);
xnor U17186 (N_17186,N_16720,N_16314);
and U17187 (N_17187,N_16711,N_16769);
xor U17188 (N_17188,N_16452,N_16235);
and U17189 (N_17189,N_16175,N_16873);
and U17190 (N_17190,N_16640,N_16103);
xnor U17191 (N_17191,N_16027,N_16791);
or U17192 (N_17192,N_16244,N_16444);
and U17193 (N_17193,N_16237,N_16205);
nand U17194 (N_17194,N_16645,N_16222);
nor U17195 (N_17195,N_16608,N_16151);
nor U17196 (N_17196,N_16157,N_16594);
xor U17197 (N_17197,N_16439,N_16557);
nand U17198 (N_17198,N_16807,N_16092);
xnor U17199 (N_17199,N_16962,N_16660);
nand U17200 (N_17200,N_16028,N_16986);
or U17201 (N_17201,N_16039,N_16801);
nor U17202 (N_17202,N_16346,N_16453);
xor U17203 (N_17203,N_16424,N_16147);
nor U17204 (N_17204,N_16787,N_16413);
nand U17205 (N_17205,N_16239,N_16513);
nand U17206 (N_17206,N_16189,N_16458);
xor U17207 (N_17207,N_16256,N_16714);
xnor U17208 (N_17208,N_16636,N_16421);
and U17209 (N_17209,N_16766,N_16808);
nor U17210 (N_17210,N_16706,N_16379);
xnor U17211 (N_17211,N_16994,N_16233);
nor U17212 (N_17212,N_16139,N_16680);
xor U17213 (N_17213,N_16898,N_16834);
nor U17214 (N_17214,N_16377,N_16738);
nor U17215 (N_17215,N_16490,N_16843);
nand U17216 (N_17216,N_16148,N_16333);
and U17217 (N_17217,N_16897,N_16326);
and U17218 (N_17218,N_16802,N_16959);
or U17219 (N_17219,N_16110,N_16925);
nand U17220 (N_17220,N_16291,N_16696);
nand U17221 (N_17221,N_16729,N_16933);
or U17222 (N_17222,N_16954,N_16007);
nand U17223 (N_17223,N_16168,N_16520);
nor U17224 (N_17224,N_16287,N_16998);
xnor U17225 (N_17225,N_16422,N_16254);
nand U17226 (N_17226,N_16573,N_16195);
or U17227 (N_17227,N_16724,N_16231);
nand U17228 (N_17228,N_16813,N_16216);
nand U17229 (N_17229,N_16449,N_16260);
nor U17230 (N_17230,N_16754,N_16047);
nor U17231 (N_17231,N_16339,N_16250);
nor U17232 (N_17232,N_16852,N_16327);
xnor U17233 (N_17233,N_16025,N_16282);
nor U17234 (N_17234,N_16336,N_16325);
nor U17235 (N_17235,N_16111,N_16089);
nand U17236 (N_17236,N_16070,N_16355);
nand U17237 (N_17237,N_16555,N_16485);
xnor U17238 (N_17238,N_16131,N_16828);
nor U17239 (N_17239,N_16507,N_16694);
xnor U17240 (N_17240,N_16457,N_16351);
nand U17241 (N_17241,N_16836,N_16514);
or U17242 (N_17242,N_16012,N_16578);
and U17243 (N_17243,N_16545,N_16033);
xor U17244 (N_17244,N_16739,N_16164);
nand U17245 (N_17245,N_16476,N_16126);
and U17246 (N_17246,N_16544,N_16529);
nor U17247 (N_17247,N_16825,N_16179);
nor U17248 (N_17248,N_16299,N_16561);
nor U17249 (N_17249,N_16269,N_16159);
nor U17250 (N_17250,N_16699,N_16685);
nand U17251 (N_17251,N_16633,N_16690);
xnor U17252 (N_17252,N_16969,N_16342);
nand U17253 (N_17253,N_16947,N_16265);
and U17254 (N_17254,N_16412,N_16576);
and U17255 (N_17255,N_16294,N_16375);
or U17256 (N_17256,N_16034,N_16844);
or U17257 (N_17257,N_16953,N_16478);
or U17258 (N_17258,N_16558,N_16255);
nor U17259 (N_17259,N_16474,N_16733);
or U17260 (N_17260,N_16644,N_16183);
and U17261 (N_17261,N_16407,N_16890);
nor U17262 (N_17262,N_16445,N_16689);
xor U17263 (N_17263,N_16527,N_16797);
and U17264 (N_17264,N_16721,N_16858);
or U17265 (N_17265,N_16924,N_16371);
and U17266 (N_17266,N_16232,N_16040);
or U17267 (N_17267,N_16041,N_16296);
xnor U17268 (N_17268,N_16534,N_16675);
xor U17269 (N_17269,N_16869,N_16616);
and U17270 (N_17270,N_16017,N_16266);
nor U17271 (N_17271,N_16353,N_16212);
and U17272 (N_17272,N_16592,N_16919);
nand U17273 (N_17273,N_16372,N_16902);
or U17274 (N_17274,N_16073,N_16038);
xor U17275 (N_17275,N_16395,N_16595);
nor U17276 (N_17276,N_16433,N_16988);
or U17277 (N_17277,N_16879,N_16820);
nand U17278 (N_17278,N_16390,N_16097);
nor U17279 (N_17279,N_16315,N_16510);
or U17280 (N_17280,N_16464,N_16405);
xor U17281 (N_17281,N_16318,N_16717);
nor U17282 (N_17282,N_16384,N_16341);
nor U17283 (N_17283,N_16823,N_16363);
nand U17284 (N_17284,N_16095,N_16094);
nand U17285 (N_17285,N_16188,N_16658);
or U17286 (N_17286,N_16763,N_16847);
or U17287 (N_17287,N_16397,N_16849);
nor U17288 (N_17288,N_16409,N_16870);
nand U17289 (N_17289,N_16833,N_16504);
nand U17290 (N_17290,N_16080,N_16249);
nor U17291 (N_17291,N_16376,N_16955);
xor U17292 (N_17292,N_16604,N_16632);
and U17293 (N_17293,N_16659,N_16821);
xnor U17294 (N_17294,N_16120,N_16887);
xnor U17295 (N_17295,N_16096,N_16077);
xnor U17296 (N_17296,N_16983,N_16775);
or U17297 (N_17297,N_16749,N_16492);
xnor U17298 (N_17298,N_16591,N_16753);
nand U17299 (N_17299,N_16570,N_16774);
xnor U17300 (N_17300,N_16185,N_16974);
and U17301 (N_17301,N_16991,N_16748);
and U17302 (N_17302,N_16161,N_16642);
or U17303 (N_17303,N_16153,N_16172);
nor U17304 (N_17304,N_16700,N_16158);
nand U17305 (N_17305,N_16572,N_16703);
nor U17306 (N_17306,N_16054,N_16614);
xnor U17307 (N_17307,N_16619,N_16750);
nor U17308 (N_17308,N_16312,N_16929);
or U17309 (N_17309,N_16114,N_16979);
nor U17310 (N_17310,N_16426,N_16764);
and U17311 (N_17311,N_16144,N_16316);
nand U17312 (N_17312,N_16083,N_16716);
or U17313 (N_17313,N_16987,N_16304);
and U17314 (N_17314,N_16892,N_16135);
nor U17315 (N_17315,N_16597,N_16132);
xor U17316 (N_17316,N_16350,N_16615);
nand U17317 (N_17317,N_16427,N_16467);
or U17318 (N_17318,N_16582,N_16509);
xnor U17319 (N_17319,N_16702,N_16854);
xor U17320 (N_17320,N_16279,N_16695);
nand U17321 (N_17321,N_16920,N_16866);
or U17322 (N_17322,N_16624,N_16000);
nand U17323 (N_17323,N_16547,N_16497);
and U17324 (N_17324,N_16672,N_16079);
and U17325 (N_17325,N_16661,N_16043);
xnor U17326 (N_17326,N_16539,N_16883);
xnor U17327 (N_17327,N_16630,N_16206);
nor U17328 (N_17328,N_16726,N_16441);
and U17329 (N_17329,N_16687,N_16471);
and U17330 (N_17330,N_16552,N_16446);
or U17331 (N_17331,N_16560,N_16343);
xor U17332 (N_17332,N_16586,N_16310);
or U17333 (N_17333,N_16618,N_16381);
nor U17334 (N_17334,N_16621,N_16187);
nor U17335 (N_17335,N_16864,N_16300);
and U17336 (N_17336,N_16967,N_16740);
xor U17337 (N_17337,N_16842,N_16536);
nand U17338 (N_17338,N_16581,N_16922);
nor U17339 (N_17339,N_16602,N_16019);
xor U17340 (N_17340,N_16393,N_16708);
or U17341 (N_17341,N_16290,N_16910);
nor U17342 (N_17342,N_16931,N_16378);
nor U17343 (N_17343,N_16646,N_16213);
nor U17344 (N_17344,N_16121,N_16874);
xnor U17345 (N_17345,N_16940,N_16528);
and U17346 (N_17346,N_16354,N_16143);
and U17347 (N_17347,N_16045,N_16901);
xnor U17348 (N_17348,N_16894,N_16511);
nand U17349 (N_17349,N_16786,N_16454);
or U17350 (N_17350,N_16611,N_16647);
and U17351 (N_17351,N_16306,N_16937);
and U17352 (N_17352,N_16086,N_16370);
nor U17353 (N_17353,N_16186,N_16691);
xnor U17354 (N_17354,N_16146,N_16589);
nand U17355 (N_17355,N_16961,N_16432);
and U17356 (N_17356,N_16877,N_16016);
or U17357 (N_17357,N_16777,N_16629);
or U17358 (N_17358,N_16277,N_16177);
nand U17359 (N_17359,N_16163,N_16368);
xor U17360 (N_17360,N_16466,N_16981);
nand U17361 (N_17361,N_16138,N_16761);
or U17362 (N_17362,N_16247,N_16196);
and U17363 (N_17363,N_16154,N_16236);
nand U17364 (N_17364,N_16283,N_16010);
nand U17365 (N_17365,N_16533,N_16001);
nand U17366 (N_17366,N_16876,N_16105);
and U17367 (N_17367,N_16909,N_16204);
nand U17368 (N_17368,N_16119,N_16600);
nand U17369 (N_17369,N_16773,N_16943);
xnor U17370 (N_17370,N_16048,N_16230);
xnor U17371 (N_17371,N_16900,N_16162);
nor U17372 (N_17372,N_16288,N_16373);
nor U17373 (N_17373,N_16440,N_16657);
xor U17374 (N_17374,N_16352,N_16501);
xnor U17375 (N_17375,N_16811,N_16568);
and U17376 (N_17376,N_16625,N_16903);
nor U17377 (N_17377,N_16637,N_16606);
nor U17378 (N_17378,N_16115,N_16789);
xor U17379 (N_17379,N_16837,N_16930);
nor U17380 (N_17380,N_16112,N_16473);
nor U17381 (N_17381,N_16686,N_16889);
nand U17382 (N_17382,N_16182,N_16246);
xnor U17383 (N_17383,N_16403,N_16975);
xor U17384 (N_17384,N_16868,N_16838);
and U17385 (N_17385,N_16936,N_16780);
nand U17386 (N_17386,N_16697,N_16243);
xnor U17387 (N_17387,N_16180,N_16118);
nor U17388 (N_17388,N_16779,N_16737);
nand U17389 (N_17389,N_16638,N_16238);
and U17390 (N_17390,N_16090,N_16101);
xnor U17391 (N_17391,N_16194,N_16710);
nand U17392 (N_17392,N_16506,N_16430);
nand U17393 (N_17393,N_16496,N_16443);
xor U17394 (N_17394,N_16722,N_16662);
nand U17395 (N_17395,N_16480,N_16515);
xor U17396 (N_17396,N_16268,N_16970);
and U17397 (N_17397,N_16732,N_16627);
nor U17398 (N_17398,N_16331,N_16093);
and U17399 (N_17399,N_16679,N_16741);
nor U17400 (N_17400,N_16130,N_16856);
nand U17401 (N_17401,N_16423,N_16156);
xnor U17402 (N_17402,N_16214,N_16434);
or U17403 (N_17403,N_16631,N_16603);
or U17404 (N_17404,N_16634,N_16952);
and U17405 (N_17405,N_16772,N_16181);
nand U17406 (N_17406,N_16295,N_16274);
xor U17407 (N_17407,N_16436,N_16483);
nor U17408 (N_17408,N_16799,N_16571);
nand U17409 (N_17409,N_16482,N_16278);
nand U17410 (N_17410,N_16907,N_16472);
nand U17411 (N_17411,N_16337,N_16015);
nor U17412 (N_17412,N_16078,N_16293);
nor U17413 (N_17413,N_16360,N_16580);
or U17414 (N_17414,N_16997,N_16210);
and U17415 (N_17415,N_16832,N_16241);
nand U17416 (N_17416,N_16550,N_16816);
or U17417 (N_17417,N_16145,N_16292);
nor U17418 (N_17418,N_16463,N_16915);
xnor U17419 (N_17419,N_16468,N_16305);
or U17420 (N_17420,N_16199,N_16727);
and U17421 (N_17421,N_16551,N_16008);
nand U17422 (N_17422,N_16261,N_16061);
xor U17423 (N_17423,N_16193,N_16171);
xnor U17424 (N_17424,N_16684,N_16031);
nand U17425 (N_17425,N_16942,N_16666);
and U17426 (N_17426,N_16345,N_16141);
xnor U17427 (N_17427,N_16822,N_16671);
nor U17428 (N_17428,N_16782,N_16429);
or U17429 (N_17429,N_16166,N_16857);
and U17430 (N_17430,N_16349,N_16263);
nand U17431 (N_17431,N_16878,N_16752);
nand U17432 (N_17432,N_16030,N_16013);
nor U17433 (N_17433,N_16203,N_16050);
or U17434 (N_17434,N_16664,N_16116);
and U17435 (N_17435,N_16081,N_16024);
nor U17436 (N_17436,N_16667,N_16322);
and U17437 (N_17437,N_16531,N_16673);
nand U17438 (N_17438,N_16538,N_16136);
nand U17439 (N_17439,N_16289,N_16905);
xnor U17440 (N_17440,N_16088,N_16776);
and U17441 (N_17441,N_16521,N_16056);
or U17442 (N_17442,N_16512,N_16949);
or U17443 (N_17443,N_16469,N_16074);
or U17444 (N_17444,N_16742,N_16174);
and U17445 (N_17445,N_16399,N_16383);
nand U17446 (N_17446,N_16563,N_16884);
or U17447 (N_17447,N_16197,N_16503);
nand U17448 (N_17448,N_16271,N_16023);
nor U17449 (N_17449,N_16770,N_16410);
or U17450 (N_17450,N_16815,N_16585);
or U17451 (N_17451,N_16935,N_16556);
or U17452 (N_17452,N_16956,N_16489);
xor U17453 (N_17453,N_16223,N_16394);
or U17454 (N_17454,N_16865,N_16519);
nor U17455 (N_17455,N_16207,N_16380);
or U17456 (N_17456,N_16009,N_16575);
and U17457 (N_17457,N_16404,N_16622);
or U17458 (N_17458,N_16224,N_16228);
xor U17459 (N_17459,N_16387,N_16804);
and U17460 (N_17460,N_16067,N_16566);
and U17461 (N_17461,N_16665,N_16701);
xor U17462 (N_17462,N_16127,N_16756);
nor U17463 (N_17463,N_16032,N_16652);
nand U17464 (N_17464,N_16066,N_16524);
nand U17465 (N_17465,N_16435,N_16518);
xor U17466 (N_17466,N_16875,N_16272);
nand U17467 (N_17467,N_16927,N_16651);
and U17468 (N_17468,N_16923,N_16588);
nand U17469 (N_17469,N_16493,N_16899);
and U17470 (N_17470,N_16020,N_16532);
and U17471 (N_17471,N_16891,N_16579);
and U17472 (N_17472,N_16743,N_16437);
nand U17473 (N_17473,N_16668,N_16281);
nor U17474 (N_17474,N_16298,N_16800);
nand U17475 (N_17475,N_16460,N_16006);
or U17476 (N_17476,N_16755,N_16916);
xor U17477 (N_17477,N_16681,N_16895);
nor U17478 (N_17478,N_16669,N_16913);
and U17479 (N_17479,N_16767,N_16549);
nor U17480 (N_17480,N_16082,N_16248);
xor U17481 (N_17481,N_16401,N_16990);
nand U17482 (N_17482,N_16234,N_16059);
and U17483 (N_17483,N_16613,N_16760);
and U17484 (N_17484,N_16461,N_16840);
and U17485 (N_17485,N_16850,N_16553);
or U17486 (N_17486,N_16425,N_16650);
nand U17487 (N_17487,N_16400,N_16976);
and U17488 (N_17488,N_16885,N_16285);
nand U17489 (N_17489,N_16736,N_16052);
or U17490 (N_17490,N_16137,N_16071);
nand U17491 (N_17491,N_16867,N_16109);
nor U17492 (N_17492,N_16465,N_16692);
nand U17493 (N_17493,N_16543,N_16839);
or U17494 (N_17494,N_16541,N_16462);
nand U17495 (N_17495,N_16053,N_16989);
or U17496 (N_17496,N_16654,N_16026);
nor U17497 (N_17497,N_16229,N_16670);
nand U17498 (N_17498,N_16406,N_16747);
nand U17499 (N_17499,N_16516,N_16108);
or U17500 (N_17500,N_16940,N_16392);
nor U17501 (N_17501,N_16708,N_16931);
nand U17502 (N_17502,N_16527,N_16054);
nor U17503 (N_17503,N_16070,N_16030);
or U17504 (N_17504,N_16566,N_16867);
xnor U17505 (N_17505,N_16135,N_16172);
or U17506 (N_17506,N_16559,N_16361);
or U17507 (N_17507,N_16089,N_16213);
xor U17508 (N_17508,N_16827,N_16823);
or U17509 (N_17509,N_16548,N_16270);
nor U17510 (N_17510,N_16845,N_16213);
xnor U17511 (N_17511,N_16967,N_16879);
nand U17512 (N_17512,N_16554,N_16845);
nor U17513 (N_17513,N_16589,N_16652);
xor U17514 (N_17514,N_16982,N_16963);
nand U17515 (N_17515,N_16434,N_16424);
and U17516 (N_17516,N_16328,N_16929);
nor U17517 (N_17517,N_16419,N_16087);
or U17518 (N_17518,N_16189,N_16559);
xnor U17519 (N_17519,N_16045,N_16303);
xnor U17520 (N_17520,N_16477,N_16035);
nand U17521 (N_17521,N_16094,N_16148);
nor U17522 (N_17522,N_16208,N_16885);
nor U17523 (N_17523,N_16438,N_16500);
nand U17524 (N_17524,N_16072,N_16056);
xnor U17525 (N_17525,N_16264,N_16105);
or U17526 (N_17526,N_16368,N_16775);
nand U17527 (N_17527,N_16889,N_16738);
and U17528 (N_17528,N_16951,N_16814);
nand U17529 (N_17529,N_16250,N_16746);
nand U17530 (N_17530,N_16439,N_16182);
and U17531 (N_17531,N_16477,N_16299);
xor U17532 (N_17532,N_16741,N_16519);
and U17533 (N_17533,N_16890,N_16426);
xnor U17534 (N_17534,N_16341,N_16017);
nor U17535 (N_17535,N_16796,N_16230);
xor U17536 (N_17536,N_16050,N_16620);
nor U17537 (N_17537,N_16938,N_16542);
or U17538 (N_17538,N_16905,N_16434);
nand U17539 (N_17539,N_16907,N_16554);
nor U17540 (N_17540,N_16506,N_16788);
nor U17541 (N_17541,N_16004,N_16756);
and U17542 (N_17542,N_16664,N_16929);
xor U17543 (N_17543,N_16227,N_16456);
xor U17544 (N_17544,N_16613,N_16043);
nand U17545 (N_17545,N_16081,N_16838);
or U17546 (N_17546,N_16873,N_16072);
xor U17547 (N_17547,N_16778,N_16785);
or U17548 (N_17548,N_16726,N_16719);
and U17549 (N_17549,N_16567,N_16297);
or U17550 (N_17550,N_16843,N_16198);
xnor U17551 (N_17551,N_16289,N_16633);
xnor U17552 (N_17552,N_16838,N_16936);
nor U17553 (N_17553,N_16919,N_16448);
nor U17554 (N_17554,N_16277,N_16198);
nand U17555 (N_17555,N_16338,N_16437);
and U17556 (N_17556,N_16616,N_16489);
xnor U17557 (N_17557,N_16547,N_16915);
xor U17558 (N_17558,N_16596,N_16679);
xor U17559 (N_17559,N_16137,N_16523);
nor U17560 (N_17560,N_16682,N_16633);
nand U17561 (N_17561,N_16575,N_16667);
and U17562 (N_17562,N_16529,N_16704);
and U17563 (N_17563,N_16582,N_16189);
and U17564 (N_17564,N_16421,N_16890);
and U17565 (N_17565,N_16003,N_16214);
nor U17566 (N_17566,N_16898,N_16328);
xor U17567 (N_17567,N_16194,N_16200);
and U17568 (N_17568,N_16062,N_16836);
or U17569 (N_17569,N_16706,N_16887);
or U17570 (N_17570,N_16337,N_16280);
xor U17571 (N_17571,N_16739,N_16512);
nor U17572 (N_17572,N_16403,N_16780);
nor U17573 (N_17573,N_16425,N_16171);
and U17574 (N_17574,N_16872,N_16180);
nand U17575 (N_17575,N_16637,N_16110);
nand U17576 (N_17576,N_16652,N_16085);
nor U17577 (N_17577,N_16403,N_16816);
xor U17578 (N_17578,N_16926,N_16495);
nor U17579 (N_17579,N_16382,N_16058);
nand U17580 (N_17580,N_16871,N_16023);
and U17581 (N_17581,N_16157,N_16265);
nor U17582 (N_17582,N_16466,N_16335);
xnor U17583 (N_17583,N_16672,N_16085);
nand U17584 (N_17584,N_16266,N_16892);
or U17585 (N_17585,N_16277,N_16472);
and U17586 (N_17586,N_16149,N_16958);
or U17587 (N_17587,N_16024,N_16994);
nand U17588 (N_17588,N_16274,N_16320);
and U17589 (N_17589,N_16828,N_16951);
xnor U17590 (N_17590,N_16819,N_16869);
and U17591 (N_17591,N_16498,N_16184);
and U17592 (N_17592,N_16815,N_16294);
nand U17593 (N_17593,N_16242,N_16073);
or U17594 (N_17594,N_16274,N_16782);
and U17595 (N_17595,N_16459,N_16340);
and U17596 (N_17596,N_16170,N_16413);
nand U17597 (N_17597,N_16400,N_16980);
nand U17598 (N_17598,N_16490,N_16216);
and U17599 (N_17599,N_16387,N_16137);
or U17600 (N_17600,N_16731,N_16668);
or U17601 (N_17601,N_16923,N_16151);
or U17602 (N_17602,N_16103,N_16413);
and U17603 (N_17603,N_16643,N_16004);
nand U17604 (N_17604,N_16586,N_16776);
xor U17605 (N_17605,N_16934,N_16418);
nor U17606 (N_17606,N_16600,N_16997);
and U17607 (N_17607,N_16780,N_16643);
xor U17608 (N_17608,N_16117,N_16893);
nand U17609 (N_17609,N_16320,N_16913);
nor U17610 (N_17610,N_16829,N_16180);
nor U17611 (N_17611,N_16757,N_16241);
or U17612 (N_17612,N_16773,N_16852);
and U17613 (N_17613,N_16609,N_16366);
and U17614 (N_17614,N_16622,N_16197);
and U17615 (N_17615,N_16060,N_16671);
or U17616 (N_17616,N_16790,N_16793);
and U17617 (N_17617,N_16082,N_16139);
and U17618 (N_17618,N_16346,N_16196);
nand U17619 (N_17619,N_16820,N_16627);
and U17620 (N_17620,N_16433,N_16614);
nor U17621 (N_17621,N_16324,N_16828);
and U17622 (N_17622,N_16169,N_16645);
nand U17623 (N_17623,N_16377,N_16222);
or U17624 (N_17624,N_16280,N_16755);
nand U17625 (N_17625,N_16082,N_16435);
nand U17626 (N_17626,N_16106,N_16318);
xnor U17627 (N_17627,N_16630,N_16945);
or U17628 (N_17628,N_16382,N_16309);
nor U17629 (N_17629,N_16502,N_16489);
and U17630 (N_17630,N_16821,N_16027);
and U17631 (N_17631,N_16121,N_16160);
nand U17632 (N_17632,N_16200,N_16456);
nor U17633 (N_17633,N_16671,N_16929);
or U17634 (N_17634,N_16492,N_16494);
nor U17635 (N_17635,N_16673,N_16984);
and U17636 (N_17636,N_16548,N_16923);
or U17637 (N_17637,N_16038,N_16552);
and U17638 (N_17638,N_16421,N_16308);
nand U17639 (N_17639,N_16701,N_16640);
and U17640 (N_17640,N_16355,N_16299);
or U17641 (N_17641,N_16200,N_16043);
or U17642 (N_17642,N_16472,N_16547);
nand U17643 (N_17643,N_16227,N_16555);
nor U17644 (N_17644,N_16205,N_16514);
xor U17645 (N_17645,N_16039,N_16572);
or U17646 (N_17646,N_16668,N_16064);
nor U17647 (N_17647,N_16362,N_16514);
xor U17648 (N_17648,N_16428,N_16855);
xnor U17649 (N_17649,N_16734,N_16614);
nor U17650 (N_17650,N_16906,N_16294);
nand U17651 (N_17651,N_16032,N_16530);
nand U17652 (N_17652,N_16316,N_16785);
or U17653 (N_17653,N_16788,N_16321);
nor U17654 (N_17654,N_16914,N_16975);
and U17655 (N_17655,N_16801,N_16697);
or U17656 (N_17656,N_16121,N_16031);
xnor U17657 (N_17657,N_16213,N_16257);
xnor U17658 (N_17658,N_16402,N_16335);
and U17659 (N_17659,N_16005,N_16914);
and U17660 (N_17660,N_16801,N_16633);
nor U17661 (N_17661,N_16170,N_16594);
nor U17662 (N_17662,N_16409,N_16937);
xnor U17663 (N_17663,N_16835,N_16950);
nor U17664 (N_17664,N_16475,N_16775);
nand U17665 (N_17665,N_16397,N_16567);
or U17666 (N_17666,N_16217,N_16604);
and U17667 (N_17667,N_16889,N_16714);
nand U17668 (N_17668,N_16327,N_16274);
and U17669 (N_17669,N_16522,N_16601);
nor U17670 (N_17670,N_16574,N_16415);
and U17671 (N_17671,N_16206,N_16858);
or U17672 (N_17672,N_16781,N_16264);
nor U17673 (N_17673,N_16638,N_16143);
and U17674 (N_17674,N_16308,N_16295);
nand U17675 (N_17675,N_16429,N_16249);
or U17676 (N_17676,N_16527,N_16189);
nor U17677 (N_17677,N_16066,N_16537);
or U17678 (N_17678,N_16017,N_16788);
nor U17679 (N_17679,N_16977,N_16551);
xnor U17680 (N_17680,N_16621,N_16473);
and U17681 (N_17681,N_16188,N_16310);
nor U17682 (N_17682,N_16474,N_16327);
or U17683 (N_17683,N_16204,N_16325);
or U17684 (N_17684,N_16220,N_16070);
or U17685 (N_17685,N_16717,N_16481);
nor U17686 (N_17686,N_16644,N_16315);
or U17687 (N_17687,N_16259,N_16850);
or U17688 (N_17688,N_16350,N_16936);
nor U17689 (N_17689,N_16788,N_16937);
or U17690 (N_17690,N_16313,N_16202);
xor U17691 (N_17691,N_16271,N_16047);
and U17692 (N_17692,N_16447,N_16252);
nor U17693 (N_17693,N_16548,N_16027);
or U17694 (N_17694,N_16497,N_16618);
xor U17695 (N_17695,N_16837,N_16437);
or U17696 (N_17696,N_16187,N_16772);
nor U17697 (N_17697,N_16564,N_16785);
nor U17698 (N_17698,N_16404,N_16831);
or U17699 (N_17699,N_16524,N_16820);
nor U17700 (N_17700,N_16783,N_16320);
nand U17701 (N_17701,N_16430,N_16431);
nand U17702 (N_17702,N_16935,N_16220);
nor U17703 (N_17703,N_16216,N_16198);
or U17704 (N_17704,N_16692,N_16966);
nand U17705 (N_17705,N_16710,N_16395);
or U17706 (N_17706,N_16960,N_16845);
and U17707 (N_17707,N_16397,N_16911);
and U17708 (N_17708,N_16235,N_16428);
nand U17709 (N_17709,N_16249,N_16575);
xor U17710 (N_17710,N_16572,N_16968);
nand U17711 (N_17711,N_16079,N_16299);
nand U17712 (N_17712,N_16914,N_16250);
nand U17713 (N_17713,N_16399,N_16659);
or U17714 (N_17714,N_16669,N_16117);
nand U17715 (N_17715,N_16555,N_16193);
nor U17716 (N_17716,N_16997,N_16837);
nand U17717 (N_17717,N_16270,N_16756);
or U17718 (N_17718,N_16432,N_16159);
xor U17719 (N_17719,N_16743,N_16054);
and U17720 (N_17720,N_16777,N_16146);
nor U17721 (N_17721,N_16212,N_16223);
or U17722 (N_17722,N_16024,N_16091);
or U17723 (N_17723,N_16107,N_16415);
nand U17724 (N_17724,N_16891,N_16842);
nand U17725 (N_17725,N_16950,N_16149);
xor U17726 (N_17726,N_16283,N_16401);
and U17727 (N_17727,N_16041,N_16834);
or U17728 (N_17728,N_16738,N_16119);
xnor U17729 (N_17729,N_16012,N_16396);
or U17730 (N_17730,N_16424,N_16856);
and U17731 (N_17731,N_16115,N_16375);
nand U17732 (N_17732,N_16994,N_16799);
nor U17733 (N_17733,N_16128,N_16267);
and U17734 (N_17734,N_16701,N_16945);
and U17735 (N_17735,N_16438,N_16493);
xor U17736 (N_17736,N_16306,N_16619);
nor U17737 (N_17737,N_16559,N_16051);
and U17738 (N_17738,N_16539,N_16270);
nor U17739 (N_17739,N_16578,N_16337);
nor U17740 (N_17740,N_16305,N_16802);
nand U17741 (N_17741,N_16563,N_16058);
xnor U17742 (N_17742,N_16792,N_16519);
nand U17743 (N_17743,N_16065,N_16750);
or U17744 (N_17744,N_16876,N_16990);
xor U17745 (N_17745,N_16462,N_16441);
xnor U17746 (N_17746,N_16106,N_16644);
nor U17747 (N_17747,N_16503,N_16984);
or U17748 (N_17748,N_16470,N_16562);
nand U17749 (N_17749,N_16574,N_16513);
and U17750 (N_17750,N_16644,N_16346);
nor U17751 (N_17751,N_16136,N_16090);
or U17752 (N_17752,N_16783,N_16546);
nor U17753 (N_17753,N_16273,N_16011);
or U17754 (N_17754,N_16287,N_16329);
nand U17755 (N_17755,N_16793,N_16990);
xor U17756 (N_17756,N_16098,N_16894);
or U17757 (N_17757,N_16247,N_16698);
and U17758 (N_17758,N_16992,N_16667);
xor U17759 (N_17759,N_16305,N_16390);
nor U17760 (N_17760,N_16257,N_16109);
and U17761 (N_17761,N_16784,N_16239);
and U17762 (N_17762,N_16757,N_16875);
nor U17763 (N_17763,N_16490,N_16341);
nand U17764 (N_17764,N_16440,N_16555);
or U17765 (N_17765,N_16589,N_16300);
and U17766 (N_17766,N_16231,N_16901);
xor U17767 (N_17767,N_16788,N_16662);
and U17768 (N_17768,N_16109,N_16140);
and U17769 (N_17769,N_16780,N_16313);
and U17770 (N_17770,N_16675,N_16370);
nand U17771 (N_17771,N_16829,N_16135);
or U17772 (N_17772,N_16647,N_16823);
nor U17773 (N_17773,N_16399,N_16563);
nor U17774 (N_17774,N_16814,N_16593);
and U17775 (N_17775,N_16283,N_16028);
nand U17776 (N_17776,N_16071,N_16367);
or U17777 (N_17777,N_16085,N_16975);
nor U17778 (N_17778,N_16419,N_16147);
or U17779 (N_17779,N_16031,N_16439);
xnor U17780 (N_17780,N_16479,N_16572);
or U17781 (N_17781,N_16145,N_16619);
and U17782 (N_17782,N_16101,N_16460);
xor U17783 (N_17783,N_16505,N_16813);
nand U17784 (N_17784,N_16005,N_16077);
nor U17785 (N_17785,N_16045,N_16482);
or U17786 (N_17786,N_16320,N_16387);
xor U17787 (N_17787,N_16866,N_16582);
nand U17788 (N_17788,N_16990,N_16276);
or U17789 (N_17789,N_16387,N_16478);
and U17790 (N_17790,N_16065,N_16914);
and U17791 (N_17791,N_16977,N_16646);
nor U17792 (N_17792,N_16385,N_16057);
nor U17793 (N_17793,N_16428,N_16476);
nor U17794 (N_17794,N_16517,N_16818);
nand U17795 (N_17795,N_16337,N_16990);
nand U17796 (N_17796,N_16275,N_16103);
nor U17797 (N_17797,N_16905,N_16115);
nor U17798 (N_17798,N_16279,N_16990);
and U17799 (N_17799,N_16104,N_16248);
nor U17800 (N_17800,N_16021,N_16383);
xor U17801 (N_17801,N_16880,N_16597);
nor U17802 (N_17802,N_16755,N_16582);
nor U17803 (N_17803,N_16725,N_16750);
xnor U17804 (N_17804,N_16939,N_16806);
or U17805 (N_17805,N_16808,N_16032);
nor U17806 (N_17806,N_16961,N_16822);
nor U17807 (N_17807,N_16262,N_16166);
and U17808 (N_17808,N_16500,N_16525);
and U17809 (N_17809,N_16158,N_16372);
xor U17810 (N_17810,N_16396,N_16256);
nand U17811 (N_17811,N_16224,N_16971);
or U17812 (N_17812,N_16063,N_16948);
and U17813 (N_17813,N_16781,N_16530);
and U17814 (N_17814,N_16608,N_16031);
and U17815 (N_17815,N_16229,N_16358);
or U17816 (N_17816,N_16458,N_16903);
or U17817 (N_17817,N_16395,N_16817);
and U17818 (N_17818,N_16877,N_16992);
nor U17819 (N_17819,N_16414,N_16062);
or U17820 (N_17820,N_16224,N_16411);
xnor U17821 (N_17821,N_16261,N_16534);
xnor U17822 (N_17822,N_16759,N_16138);
nand U17823 (N_17823,N_16363,N_16335);
nand U17824 (N_17824,N_16789,N_16377);
nand U17825 (N_17825,N_16164,N_16199);
and U17826 (N_17826,N_16846,N_16426);
xnor U17827 (N_17827,N_16294,N_16536);
xnor U17828 (N_17828,N_16380,N_16019);
and U17829 (N_17829,N_16176,N_16029);
or U17830 (N_17830,N_16581,N_16420);
nand U17831 (N_17831,N_16543,N_16619);
and U17832 (N_17832,N_16042,N_16534);
and U17833 (N_17833,N_16356,N_16321);
nand U17834 (N_17834,N_16942,N_16109);
xnor U17835 (N_17835,N_16248,N_16310);
or U17836 (N_17836,N_16139,N_16437);
nand U17837 (N_17837,N_16061,N_16169);
nand U17838 (N_17838,N_16786,N_16374);
and U17839 (N_17839,N_16563,N_16281);
nor U17840 (N_17840,N_16416,N_16329);
or U17841 (N_17841,N_16871,N_16887);
or U17842 (N_17842,N_16508,N_16719);
and U17843 (N_17843,N_16421,N_16286);
and U17844 (N_17844,N_16595,N_16834);
nor U17845 (N_17845,N_16394,N_16850);
or U17846 (N_17846,N_16305,N_16761);
nor U17847 (N_17847,N_16884,N_16971);
or U17848 (N_17848,N_16190,N_16386);
or U17849 (N_17849,N_16490,N_16946);
xnor U17850 (N_17850,N_16424,N_16627);
xor U17851 (N_17851,N_16524,N_16426);
xnor U17852 (N_17852,N_16757,N_16765);
and U17853 (N_17853,N_16083,N_16326);
or U17854 (N_17854,N_16350,N_16801);
and U17855 (N_17855,N_16743,N_16137);
and U17856 (N_17856,N_16135,N_16683);
nand U17857 (N_17857,N_16072,N_16260);
nor U17858 (N_17858,N_16908,N_16902);
xnor U17859 (N_17859,N_16398,N_16065);
xor U17860 (N_17860,N_16258,N_16704);
nor U17861 (N_17861,N_16589,N_16649);
nor U17862 (N_17862,N_16461,N_16707);
xor U17863 (N_17863,N_16267,N_16594);
and U17864 (N_17864,N_16124,N_16791);
nor U17865 (N_17865,N_16206,N_16417);
or U17866 (N_17866,N_16374,N_16726);
nand U17867 (N_17867,N_16483,N_16053);
xor U17868 (N_17868,N_16954,N_16051);
xnor U17869 (N_17869,N_16519,N_16518);
or U17870 (N_17870,N_16527,N_16613);
nand U17871 (N_17871,N_16355,N_16251);
xnor U17872 (N_17872,N_16627,N_16620);
nand U17873 (N_17873,N_16755,N_16372);
and U17874 (N_17874,N_16480,N_16504);
or U17875 (N_17875,N_16318,N_16744);
xnor U17876 (N_17876,N_16437,N_16514);
nor U17877 (N_17877,N_16215,N_16414);
or U17878 (N_17878,N_16487,N_16696);
or U17879 (N_17879,N_16614,N_16073);
or U17880 (N_17880,N_16725,N_16387);
xor U17881 (N_17881,N_16009,N_16006);
nor U17882 (N_17882,N_16552,N_16378);
or U17883 (N_17883,N_16088,N_16751);
xor U17884 (N_17884,N_16267,N_16609);
or U17885 (N_17885,N_16736,N_16498);
and U17886 (N_17886,N_16983,N_16187);
nand U17887 (N_17887,N_16749,N_16892);
xor U17888 (N_17888,N_16933,N_16851);
or U17889 (N_17889,N_16937,N_16281);
or U17890 (N_17890,N_16932,N_16199);
nand U17891 (N_17891,N_16237,N_16250);
or U17892 (N_17892,N_16283,N_16487);
nor U17893 (N_17893,N_16233,N_16125);
and U17894 (N_17894,N_16118,N_16099);
and U17895 (N_17895,N_16919,N_16944);
nor U17896 (N_17896,N_16706,N_16117);
and U17897 (N_17897,N_16962,N_16267);
xnor U17898 (N_17898,N_16939,N_16555);
xnor U17899 (N_17899,N_16235,N_16040);
or U17900 (N_17900,N_16124,N_16049);
nor U17901 (N_17901,N_16879,N_16186);
and U17902 (N_17902,N_16421,N_16641);
xor U17903 (N_17903,N_16511,N_16231);
or U17904 (N_17904,N_16918,N_16131);
and U17905 (N_17905,N_16785,N_16021);
xnor U17906 (N_17906,N_16968,N_16840);
nand U17907 (N_17907,N_16863,N_16107);
nor U17908 (N_17908,N_16302,N_16809);
nor U17909 (N_17909,N_16020,N_16822);
nand U17910 (N_17910,N_16907,N_16433);
and U17911 (N_17911,N_16488,N_16723);
or U17912 (N_17912,N_16327,N_16430);
xnor U17913 (N_17913,N_16447,N_16230);
and U17914 (N_17914,N_16267,N_16135);
xnor U17915 (N_17915,N_16988,N_16954);
nand U17916 (N_17916,N_16454,N_16400);
nor U17917 (N_17917,N_16382,N_16224);
xnor U17918 (N_17918,N_16559,N_16468);
xor U17919 (N_17919,N_16016,N_16371);
or U17920 (N_17920,N_16426,N_16330);
xnor U17921 (N_17921,N_16238,N_16487);
nor U17922 (N_17922,N_16054,N_16217);
or U17923 (N_17923,N_16246,N_16611);
or U17924 (N_17924,N_16474,N_16208);
or U17925 (N_17925,N_16305,N_16449);
nor U17926 (N_17926,N_16973,N_16681);
xnor U17927 (N_17927,N_16165,N_16599);
or U17928 (N_17928,N_16592,N_16953);
nand U17929 (N_17929,N_16614,N_16935);
xor U17930 (N_17930,N_16336,N_16863);
nor U17931 (N_17931,N_16002,N_16784);
and U17932 (N_17932,N_16174,N_16847);
xor U17933 (N_17933,N_16805,N_16279);
and U17934 (N_17934,N_16676,N_16137);
nor U17935 (N_17935,N_16068,N_16259);
xor U17936 (N_17936,N_16190,N_16765);
nand U17937 (N_17937,N_16572,N_16684);
and U17938 (N_17938,N_16300,N_16674);
nand U17939 (N_17939,N_16789,N_16682);
xnor U17940 (N_17940,N_16538,N_16740);
nor U17941 (N_17941,N_16709,N_16812);
xor U17942 (N_17942,N_16987,N_16087);
nor U17943 (N_17943,N_16110,N_16302);
and U17944 (N_17944,N_16875,N_16125);
xor U17945 (N_17945,N_16316,N_16656);
and U17946 (N_17946,N_16736,N_16579);
nor U17947 (N_17947,N_16671,N_16807);
xnor U17948 (N_17948,N_16950,N_16812);
and U17949 (N_17949,N_16381,N_16458);
xnor U17950 (N_17950,N_16619,N_16212);
nand U17951 (N_17951,N_16668,N_16857);
xnor U17952 (N_17952,N_16798,N_16936);
and U17953 (N_17953,N_16681,N_16202);
and U17954 (N_17954,N_16098,N_16092);
nand U17955 (N_17955,N_16399,N_16879);
xor U17956 (N_17956,N_16891,N_16117);
or U17957 (N_17957,N_16646,N_16824);
xnor U17958 (N_17958,N_16598,N_16470);
xor U17959 (N_17959,N_16114,N_16747);
nand U17960 (N_17960,N_16329,N_16057);
xor U17961 (N_17961,N_16331,N_16532);
and U17962 (N_17962,N_16110,N_16042);
xor U17963 (N_17963,N_16086,N_16772);
nor U17964 (N_17964,N_16313,N_16965);
nor U17965 (N_17965,N_16896,N_16011);
nand U17966 (N_17966,N_16309,N_16727);
nand U17967 (N_17967,N_16352,N_16393);
nor U17968 (N_17968,N_16302,N_16245);
nand U17969 (N_17969,N_16822,N_16399);
and U17970 (N_17970,N_16371,N_16806);
and U17971 (N_17971,N_16229,N_16742);
and U17972 (N_17972,N_16742,N_16692);
nand U17973 (N_17973,N_16709,N_16135);
or U17974 (N_17974,N_16224,N_16563);
nand U17975 (N_17975,N_16513,N_16224);
or U17976 (N_17976,N_16678,N_16492);
or U17977 (N_17977,N_16497,N_16442);
nand U17978 (N_17978,N_16358,N_16700);
nor U17979 (N_17979,N_16230,N_16445);
or U17980 (N_17980,N_16733,N_16817);
xnor U17981 (N_17981,N_16553,N_16673);
nor U17982 (N_17982,N_16582,N_16925);
or U17983 (N_17983,N_16848,N_16025);
nand U17984 (N_17984,N_16066,N_16649);
xnor U17985 (N_17985,N_16747,N_16674);
xnor U17986 (N_17986,N_16330,N_16382);
xnor U17987 (N_17987,N_16171,N_16936);
nor U17988 (N_17988,N_16303,N_16400);
or U17989 (N_17989,N_16138,N_16047);
nor U17990 (N_17990,N_16696,N_16729);
or U17991 (N_17991,N_16439,N_16720);
or U17992 (N_17992,N_16702,N_16143);
and U17993 (N_17993,N_16221,N_16915);
xor U17994 (N_17994,N_16083,N_16472);
nor U17995 (N_17995,N_16827,N_16844);
nor U17996 (N_17996,N_16351,N_16603);
xnor U17997 (N_17997,N_16736,N_16775);
and U17998 (N_17998,N_16405,N_16171);
xor U17999 (N_17999,N_16133,N_16644);
or U18000 (N_18000,N_17880,N_17593);
xor U18001 (N_18001,N_17500,N_17585);
nor U18002 (N_18002,N_17219,N_17730);
xnor U18003 (N_18003,N_17360,N_17586);
nand U18004 (N_18004,N_17706,N_17042);
or U18005 (N_18005,N_17336,N_17617);
nor U18006 (N_18006,N_17134,N_17418);
or U18007 (N_18007,N_17731,N_17115);
nand U18008 (N_18008,N_17169,N_17697);
nor U18009 (N_18009,N_17061,N_17338);
or U18010 (N_18010,N_17849,N_17653);
nand U18011 (N_18011,N_17898,N_17078);
xor U18012 (N_18012,N_17856,N_17794);
nand U18013 (N_18013,N_17575,N_17105);
xor U18014 (N_18014,N_17170,N_17840);
nand U18015 (N_18015,N_17453,N_17519);
and U18016 (N_18016,N_17168,N_17759);
nand U18017 (N_18017,N_17532,N_17292);
or U18018 (N_18018,N_17309,N_17761);
nor U18019 (N_18019,N_17234,N_17238);
or U18020 (N_18020,N_17518,N_17404);
nor U18021 (N_18021,N_17414,N_17574);
xnor U18022 (N_18022,N_17075,N_17356);
nor U18023 (N_18023,N_17290,N_17311);
nor U18024 (N_18024,N_17273,N_17452);
nand U18025 (N_18025,N_17122,N_17663);
nor U18026 (N_18026,N_17627,N_17304);
nand U18027 (N_18027,N_17968,N_17685);
or U18028 (N_18028,N_17397,N_17364);
nor U18029 (N_18029,N_17215,N_17354);
nand U18030 (N_18030,N_17071,N_17307);
nor U18031 (N_18031,N_17295,N_17337);
or U18032 (N_18032,N_17953,N_17654);
and U18033 (N_18033,N_17989,N_17040);
and U18034 (N_18034,N_17358,N_17068);
nand U18035 (N_18035,N_17264,N_17220);
or U18036 (N_18036,N_17463,N_17941);
xor U18037 (N_18037,N_17276,N_17736);
xor U18038 (N_18038,N_17510,N_17966);
and U18039 (N_18039,N_17462,N_17227);
xnor U18040 (N_18040,N_17063,N_17378);
xnor U18041 (N_18041,N_17286,N_17380);
and U18042 (N_18042,N_17490,N_17249);
nand U18043 (N_18043,N_17480,N_17353);
xnor U18044 (N_18044,N_17515,N_17504);
or U18045 (N_18045,N_17324,N_17280);
nor U18046 (N_18046,N_17434,N_17154);
nor U18047 (N_18047,N_17606,N_17955);
xnor U18048 (N_18048,N_17177,N_17862);
or U18049 (N_18049,N_17657,N_17881);
xor U18050 (N_18050,N_17130,N_17211);
and U18051 (N_18051,N_17031,N_17143);
or U18052 (N_18052,N_17066,N_17098);
or U18053 (N_18053,N_17121,N_17330);
or U18054 (N_18054,N_17164,N_17628);
nor U18055 (N_18055,N_17086,N_17120);
and U18056 (N_18056,N_17402,N_17080);
or U18057 (N_18057,N_17832,N_17316);
nor U18058 (N_18058,N_17808,N_17967);
nand U18059 (N_18059,N_17693,N_17781);
nand U18060 (N_18060,N_17376,N_17952);
xor U18061 (N_18061,N_17251,N_17332);
nand U18062 (N_18062,N_17538,N_17702);
nand U18063 (N_18063,N_17253,N_17159);
and U18064 (N_18064,N_17647,N_17436);
nor U18065 (N_18065,N_17558,N_17509);
and U18066 (N_18066,N_17624,N_17481);
and U18067 (N_18067,N_17934,N_17455);
nor U18068 (N_18068,N_17384,N_17587);
xnor U18069 (N_18069,N_17357,N_17093);
nor U18070 (N_18070,N_17132,N_17118);
and U18071 (N_18071,N_17788,N_17834);
or U18072 (N_18072,N_17493,N_17554);
nor U18073 (N_18073,N_17416,N_17770);
or U18074 (N_18074,N_17431,N_17839);
xor U18075 (N_18075,N_17923,N_17870);
nand U18076 (N_18076,N_17607,N_17858);
nand U18077 (N_18077,N_17799,N_17724);
nor U18078 (N_18078,N_17676,N_17537);
and U18079 (N_18079,N_17508,N_17263);
or U18080 (N_18080,N_17938,N_17331);
nor U18081 (N_18081,N_17056,N_17296);
nand U18082 (N_18082,N_17461,N_17597);
nand U18083 (N_18083,N_17872,N_17076);
or U18084 (N_18084,N_17725,N_17720);
nand U18085 (N_18085,N_17729,N_17100);
and U18086 (N_18086,N_17682,N_17392);
nand U18087 (N_18087,N_17648,N_17454);
or U18088 (N_18088,N_17494,N_17757);
and U18089 (N_18089,N_17630,N_17909);
nand U18090 (N_18090,N_17861,N_17795);
xor U18091 (N_18091,N_17990,N_17008);
xnor U18092 (N_18092,N_17974,N_17689);
or U18093 (N_18093,N_17368,N_17014);
or U18094 (N_18094,N_17235,N_17279);
xnor U18095 (N_18095,N_17813,N_17433);
xnor U18096 (N_18096,N_17541,N_17780);
and U18097 (N_18097,N_17787,N_17301);
xor U18098 (N_18098,N_17440,N_17860);
nand U18099 (N_18099,N_17172,N_17087);
and U18100 (N_18100,N_17944,N_17284);
xor U18101 (N_18101,N_17717,N_17456);
and U18102 (N_18102,N_17678,N_17176);
nor U18103 (N_18103,N_17171,N_17252);
xor U18104 (N_18104,N_17435,N_17668);
and U18105 (N_18105,N_17970,N_17800);
or U18106 (N_18106,N_17831,N_17728);
nor U18107 (N_18107,N_17529,N_17988);
xnor U18108 (N_18108,N_17660,N_17527);
and U18109 (N_18109,N_17517,N_17469);
xor U18110 (N_18110,N_17041,N_17045);
nor U18111 (N_18111,N_17244,N_17283);
or U18112 (N_18112,N_17820,N_17672);
and U18113 (N_18113,N_17409,N_17233);
xnor U18114 (N_18114,N_17084,N_17686);
nor U18115 (N_18115,N_17015,N_17741);
nor U18116 (N_18116,N_17260,N_17393);
nor U18117 (N_18117,N_17323,N_17700);
or U18118 (N_18118,N_17748,N_17466);
nor U18119 (N_18119,N_17767,N_17889);
or U18120 (N_18120,N_17305,N_17407);
nor U18121 (N_18121,N_17327,N_17012);
xnor U18122 (N_18122,N_17605,N_17719);
xnor U18123 (N_18123,N_17072,N_17125);
nand U18124 (N_18124,N_17894,N_17218);
or U18125 (N_18125,N_17557,N_17603);
nand U18126 (N_18126,N_17536,N_17108);
or U18127 (N_18127,N_17773,N_17312);
xor U18128 (N_18128,N_17194,N_17888);
and U18129 (N_18129,N_17341,N_17282);
or U18130 (N_18130,N_17184,N_17670);
or U18131 (N_18131,N_17225,N_17101);
xor U18132 (N_18132,N_17733,N_17265);
and U18133 (N_18133,N_17289,N_17037);
nor U18134 (N_18134,N_17425,N_17851);
xor U18135 (N_18135,N_17957,N_17188);
nand U18136 (N_18136,N_17954,N_17921);
xnor U18137 (N_18137,N_17222,N_17548);
nand U18138 (N_18138,N_17885,N_17326);
nor U18139 (N_18139,N_17698,N_17403);
or U18140 (N_18140,N_17577,N_17415);
or U18141 (N_18141,N_17900,N_17027);
and U18142 (N_18142,N_17762,N_17530);
xor U18143 (N_18143,N_17544,N_17300);
xor U18144 (N_18144,N_17531,N_17285);
nor U18145 (N_18145,N_17314,N_17918);
nor U18146 (N_18146,N_17993,N_17691);
nand U18147 (N_18147,N_17514,N_17058);
nor U18148 (N_18148,N_17444,N_17542);
and U18149 (N_18149,N_17334,N_17578);
or U18150 (N_18150,N_17250,N_17569);
nand U18151 (N_18151,N_17568,N_17951);
or U18152 (N_18152,N_17038,N_17180);
nand U18153 (N_18153,N_17204,N_17810);
nand U18154 (N_18154,N_17620,N_17343);
nand U18155 (N_18155,N_17398,N_17916);
xnor U18156 (N_18156,N_17147,N_17319);
xnor U18157 (N_18157,N_17223,N_17271);
xnor U18158 (N_18158,N_17566,N_17303);
and U18159 (N_18159,N_17915,N_17884);
and U18160 (N_18160,N_17011,N_17024);
and U18161 (N_18161,N_17774,N_17026);
nand U18162 (N_18162,N_17209,N_17644);
nor U18163 (N_18163,N_17502,N_17248);
nand U18164 (N_18164,N_17842,N_17294);
nor U18165 (N_18165,N_17136,N_17789);
nor U18166 (N_18166,N_17556,N_17550);
and U18167 (N_18167,N_17727,N_17083);
and U18168 (N_18168,N_17838,N_17847);
and U18169 (N_18169,N_17895,N_17595);
xor U18170 (N_18170,N_17474,N_17412);
nor U18171 (N_18171,N_17257,N_17359);
nor U18172 (N_18172,N_17287,N_17346);
nor U18173 (N_18173,N_17023,N_17032);
nand U18174 (N_18174,N_17449,N_17546);
or U18175 (N_18175,N_17675,N_17158);
and U18176 (N_18176,N_17344,N_17123);
nand U18177 (N_18177,N_17389,N_17124);
and U18178 (N_18178,N_17588,N_17961);
nor U18179 (N_18179,N_17755,N_17793);
and U18180 (N_18180,N_17166,N_17138);
and U18181 (N_18181,N_17293,N_17520);
nand U18182 (N_18182,N_17598,N_17854);
and U18183 (N_18183,N_17362,N_17299);
xor U18184 (N_18184,N_17109,N_17210);
nand U18185 (N_18185,N_17723,N_17448);
and U18186 (N_18186,N_17665,N_17708);
or U18187 (N_18187,N_17768,N_17740);
xor U18188 (N_18188,N_17491,N_17367);
nor U18189 (N_18189,N_17812,N_17406);
nand U18190 (N_18190,N_17703,N_17712);
nor U18191 (N_18191,N_17459,N_17096);
or U18192 (N_18192,N_17313,N_17460);
nand U18193 (N_18193,N_17877,N_17528);
and U18194 (N_18194,N_17131,N_17796);
nor U18195 (N_18195,N_17734,N_17874);
and U18196 (N_18196,N_17201,N_17361);
and U18197 (N_18197,N_17427,N_17973);
nand U18198 (N_18198,N_17772,N_17377);
xor U18199 (N_18199,N_17472,N_17417);
or U18200 (N_18200,N_17226,N_17410);
nor U18201 (N_18201,N_17266,N_17447);
nand U18202 (N_18202,N_17906,N_17196);
or U18203 (N_18203,N_17278,N_17174);
xor U18204 (N_18204,N_17875,N_17231);
xor U18205 (N_18205,N_17713,N_17828);
nor U18206 (N_18206,N_17864,N_17545);
or U18207 (N_18207,N_17516,N_17352);
nand U18208 (N_18208,N_17609,N_17479);
nor U18209 (N_18209,N_17625,N_17614);
or U18210 (N_18210,N_17661,N_17621);
nor U18211 (N_18211,N_17571,N_17564);
and U18212 (N_18212,N_17029,N_17200);
nand U18213 (N_18213,N_17555,N_17043);
nand U18214 (N_18214,N_17333,N_17738);
xnor U18215 (N_18215,N_17424,N_17651);
xor U18216 (N_18216,N_17565,N_17189);
nand U18217 (N_18217,N_17743,N_17411);
or U18218 (N_18218,N_17107,N_17601);
nor U18219 (N_18219,N_17010,N_17423);
nand U18220 (N_18220,N_17945,N_17985);
nand U18221 (N_18221,N_17638,N_17369);
nor U18222 (N_18222,N_17099,N_17744);
and U18223 (N_18223,N_17203,N_17005);
nor U18224 (N_18224,N_17937,N_17929);
and U18225 (N_18225,N_17792,N_17582);
or U18226 (N_18226,N_17814,N_17821);
nand U18227 (N_18227,N_17212,N_17674);
xnor U18228 (N_18228,N_17751,N_17395);
and U18229 (N_18229,N_17382,N_17205);
xor U18230 (N_18230,N_17195,N_17737);
xnor U18231 (N_18231,N_17892,N_17901);
nand U18232 (N_18232,N_17347,N_17385);
and U18233 (N_18233,N_17155,N_17866);
and U18234 (N_18234,N_17245,N_17470);
nor U18235 (N_18235,N_17464,N_17948);
or U18236 (N_18236,N_17057,N_17394);
xor U18237 (N_18237,N_17028,N_17467);
and U18238 (N_18238,N_17683,N_17830);
and U18239 (N_18239,N_17752,N_17476);
and U18240 (N_18240,N_17776,N_17562);
nor U18241 (N_18241,N_17735,N_17206);
and U18242 (N_18242,N_17230,N_17050);
nor U18243 (N_18243,N_17443,N_17513);
and U18244 (N_18244,N_17034,N_17855);
or U18245 (N_18245,N_17650,N_17659);
or U18246 (N_18246,N_17002,N_17498);
or U18247 (N_18247,N_17863,N_17694);
nand U18248 (N_18248,N_17329,N_17576);
xnor U18249 (N_18249,N_17458,N_17869);
or U18250 (N_18250,N_17190,N_17355);
nor U18251 (N_18251,N_17186,N_17950);
nand U18252 (N_18252,N_17859,N_17615);
or U18253 (N_18253,N_17589,N_17254);
or U18254 (N_18254,N_17742,N_17580);
xnor U18255 (N_18255,N_17065,N_17696);
or U18256 (N_18256,N_17949,N_17039);
nor U18257 (N_18257,N_17972,N_17386);
nor U18258 (N_18258,N_17996,N_17485);
and U18259 (N_18259,N_17766,N_17999);
nor U18260 (N_18260,N_17635,N_17927);
nor U18261 (N_18261,N_17809,N_17350);
nor U18262 (N_18262,N_17306,N_17687);
or U18263 (N_18263,N_17786,N_17649);
nand U18264 (N_18264,N_17262,N_17202);
and U18265 (N_18265,N_17963,N_17471);
and U18266 (N_18266,N_17383,N_17247);
or U18267 (N_18267,N_17317,N_17797);
and U18268 (N_18268,N_17511,N_17871);
nand U18269 (N_18269,N_17632,N_17910);
xnor U18270 (N_18270,N_17399,N_17618);
nor U18271 (N_18271,N_17887,N_17714);
and U18272 (N_18272,N_17473,N_17976);
nand U18273 (N_18273,N_17497,N_17771);
xor U18274 (N_18274,N_17995,N_17718);
xor U18275 (N_18275,N_17704,N_17825);
and U18276 (N_18276,N_17298,N_17432);
or U18277 (N_18277,N_17259,N_17006);
or U18278 (N_18278,N_17321,N_17335);
xor U18279 (N_18279,N_17082,N_17126);
xnor U18280 (N_18280,N_17805,N_17827);
nand U18281 (N_18281,N_17419,N_17631);
xnor U18282 (N_18282,N_17882,N_17522);
and U18283 (N_18283,N_17465,N_17960);
nor U18284 (N_18284,N_17077,N_17000);
nand U18285 (N_18285,N_17505,N_17549);
and U18286 (N_18286,N_17173,N_17629);
nand U18287 (N_18287,N_17913,N_17818);
xor U18288 (N_18288,N_17388,N_17604);
xnor U18289 (N_18289,N_17030,N_17156);
nor U18290 (N_18290,N_17085,N_17020);
nor U18291 (N_18291,N_17987,N_17157);
nor U18292 (N_18292,N_17148,N_17701);
nor U18293 (N_18293,N_17381,N_17833);
nand U18294 (N_18294,N_17681,N_17645);
or U18295 (N_18295,N_17763,N_17179);
nor U18296 (N_18296,N_17599,N_17823);
and U18297 (N_18297,N_17062,N_17992);
or U18298 (N_18298,N_17193,N_17239);
nand U18299 (N_18299,N_17070,N_17097);
or U18300 (N_18300,N_17667,N_17496);
or U18301 (N_18301,N_17373,N_17001);
nand U18302 (N_18302,N_17745,N_17591);
nor U18303 (N_18303,N_17052,N_17268);
xor U18304 (N_18304,N_17561,N_17836);
nor U18305 (N_18305,N_17750,N_17739);
and U18306 (N_18306,N_17845,N_17016);
or U18307 (N_18307,N_17930,N_17711);
nor U18308 (N_18308,N_17602,N_17904);
nand U18309 (N_18309,N_17939,N_17181);
and U18310 (N_18310,N_17563,N_17981);
nor U18311 (N_18311,N_17983,N_17060);
and U18312 (N_18312,N_17804,N_17710);
nand U18313 (N_18313,N_17004,N_17634);
and U18314 (N_18314,N_17413,N_17903);
xnor U18315 (N_18315,N_17371,N_17666);
and U18316 (N_18316,N_17664,N_17408);
nand U18317 (N_18317,N_17009,N_17446);
and U18318 (N_18318,N_17662,N_17328);
nor U18319 (N_18319,N_17348,N_17658);
or U18320 (N_18320,N_17611,N_17053);
and U18321 (N_18321,N_17499,N_17198);
nor U18322 (N_18322,N_17274,N_17868);
nand U18323 (N_18323,N_17920,N_17161);
xor U18324 (N_18324,N_17288,N_17133);
nand U18325 (N_18325,N_17197,N_17089);
xnor U18326 (N_18326,N_17102,N_17837);
and U18327 (N_18327,N_17322,N_17090);
xor U18328 (N_18328,N_17583,N_17256);
nand U18329 (N_18329,N_17092,N_17552);
or U18330 (N_18330,N_17094,N_17081);
and U18331 (N_18331,N_17401,N_17656);
and U18332 (N_18332,N_17936,N_17022);
and U18333 (N_18333,N_17119,N_17139);
nand U18334 (N_18334,N_17917,N_17110);
xnor U18335 (N_18335,N_17162,N_17521);
and U18336 (N_18336,N_17325,N_17732);
nor U18337 (N_18337,N_17764,N_17104);
or U18338 (N_18338,N_17572,N_17844);
xnor U18339 (N_18339,N_17044,N_17946);
and U18340 (N_18340,N_17815,N_17997);
or U18341 (N_18341,N_17457,N_17149);
xnor U18342 (N_18342,N_17857,N_17495);
nor U18343 (N_18343,N_17451,N_17979);
xor U18344 (N_18344,N_17145,N_17958);
and U18345 (N_18345,N_17229,N_17214);
nand U18346 (N_18346,N_17551,N_17379);
or U18347 (N_18347,N_17940,N_17146);
xor U18348 (N_18348,N_17144,N_17971);
xor U18349 (N_18349,N_17486,N_17051);
nor U18350 (N_18350,N_17852,N_17956);
and U18351 (N_18351,N_17965,N_17873);
or U18352 (N_18352,N_17641,N_17308);
nor U18353 (N_18353,N_17524,N_17567);
or U18354 (N_18354,N_17366,N_17978);
and U18355 (N_18355,N_17726,N_17779);
and U18356 (N_18356,N_17592,N_17281);
nor U18357 (N_18357,N_17420,N_17243);
nor U18358 (N_18358,N_17912,N_17964);
nand U18359 (N_18359,N_17943,N_17112);
or U18360 (N_18360,N_17754,N_17269);
or U18361 (N_18361,N_17579,N_17207);
nand U18362 (N_18362,N_17896,N_17816);
and U18363 (N_18363,N_17919,N_17539);
and U18364 (N_18364,N_17320,N_17152);
nand U18365 (N_18365,N_17374,N_17370);
nor U18366 (N_18366,N_17931,N_17709);
or U18367 (N_18367,N_17492,N_17533);
nor U18368 (N_18368,N_17807,N_17817);
xnor U18369 (N_18369,N_17643,N_17275);
or U18370 (N_18370,N_17035,N_17850);
nor U18371 (N_18371,N_17942,N_17526);
xor U18372 (N_18372,N_17560,N_17705);
or U18373 (N_18373,N_17342,N_17778);
and U18374 (N_18374,N_17506,N_17475);
or U18375 (N_18375,N_17396,N_17707);
or U18376 (N_18376,N_17258,N_17986);
xnor U18377 (N_18377,N_17876,N_17907);
nand U18378 (N_18378,N_17540,N_17242);
or U18379 (N_18379,N_17153,N_17192);
xnor U18380 (N_18380,N_17843,N_17074);
and U18381 (N_18381,N_17932,N_17722);
nor U18382 (N_18382,N_17372,N_17902);
nor U18383 (N_18383,N_17600,N_17477);
nand U18384 (N_18384,N_17246,N_17046);
xor U18385 (N_18385,N_17947,N_17749);
or U18386 (N_18386,N_17255,N_17160);
nand U18387 (N_18387,N_17426,N_17982);
nand U18388 (N_18388,N_17114,N_17962);
or U18389 (N_18389,N_17117,N_17182);
xor U18390 (N_18390,N_17191,N_17547);
or U18391 (N_18391,N_17622,N_17135);
xnor U18392 (N_18392,N_17669,N_17049);
and U18393 (N_18393,N_17232,N_17073);
xnor U18394 (N_18394,N_17984,N_17018);
or U18395 (N_18395,N_17261,N_17482);
nor U18396 (N_18396,N_17975,N_17777);
nor U18397 (N_18397,N_17183,N_17679);
xnor U18398 (N_18398,N_17891,N_17914);
or U18399 (N_18399,N_17178,N_17573);
nand U18400 (N_18400,N_17784,N_17695);
xor U18401 (N_18401,N_17503,N_17439);
nand U18402 (N_18402,N_17908,N_17747);
and U18403 (N_18403,N_17835,N_17637);
nor U18404 (N_18404,N_17802,N_17584);
or U18405 (N_18405,N_17775,N_17596);
nor U18406 (N_18406,N_17512,N_17400);
nand U18407 (N_18407,N_17199,N_17428);
or U18408 (N_18408,N_17095,N_17626);
xnor U18409 (N_18409,N_17213,N_17187);
xor U18410 (N_18410,N_17865,N_17345);
nand U18411 (N_18411,N_17017,N_17003);
nor U18412 (N_18412,N_17692,N_17430);
or U18413 (N_18413,N_17619,N_17534);
nand U18414 (N_18414,N_17523,N_17570);
xor U18415 (N_18415,N_17899,N_17608);
and U18416 (N_18416,N_17760,N_17765);
xnor U18417 (N_18417,N_17853,N_17228);
or U18418 (N_18418,N_17445,N_17142);
or U18419 (N_18419,N_17277,N_17911);
nor U18420 (N_18420,N_17067,N_17994);
nand U18421 (N_18421,N_17824,N_17151);
xnor U18422 (N_18422,N_17310,N_17021);
and U18423 (N_18423,N_17088,N_17237);
nor U18424 (N_18424,N_17033,N_17848);
and U18425 (N_18425,N_17867,N_17064);
xor U18426 (N_18426,N_17025,N_17878);
and U18427 (N_18427,N_17216,N_17886);
or U18428 (N_18428,N_17442,N_17240);
and U18429 (N_18429,N_17801,N_17141);
xnor U18430 (N_18430,N_17128,N_17349);
and U18431 (N_18431,N_17208,N_17150);
nor U18432 (N_18432,N_17048,N_17127);
or U18433 (N_18433,N_17488,N_17340);
xnor U18434 (N_18434,N_17935,N_17113);
nor U18435 (N_18435,N_17391,N_17036);
xor U18436 (N_18436,N_17924,N_17933);
xor U18437 (N_18437,N_17829,N_17925);
xnor U18438 (N_18438,N_17291,N_17613);
nand U18439 (N_18439,N_17525,N_17175);
nand U18440 (N_18440,N_17217,N_17928);
and U18441 (N_18441,N_17103,N_17811);
nor U18442 (N_18442,N_17688,N_17959);
nor U18443 (N_18443,N_17363,N_17047);
nand U18444 (N_18444,N_17581,N_17421);
nand U18445 (N_18445,N_17422,N_17055);
or U18446 (N_18446,N_17441,N_17069);
nand U18447 (N_18447,N_17543,N_17819);
nor U18448 (N_18448,N_17616,N_17883);
or U18449 (N_18449,N_17980,N_17339);
and U18450 (N_18450,N_17302,N_17922);
xnor U18451 (N_18451,N_17140,N_17826);
or U18452 (N_18452,N_17137,N_17437);
nor U18453 (N_18453,N_17351,N_17646);
nor U18454 (N_18454,N_17267,N_17535);
or U18455 (N_18455,N_17106,N_17716);
or U18456 (N_18456,N_17639,N_17977);
and U18457 (N_18457,N_17315,N_17468);
nor U18458 (N_18458,N_17803,N_17905);
and U18459 (N_18459,N_17926,N_17297);
nor U18460 (N_18460,N_17487,N_17841);
and U18461 (N_18461,N_17756,N_17438);
nor U18462 (N_18462,N_17721,N_17270);
and U18463 (N_18463,N_17623,N_17241);
nor U18464 (N_18464,N_17507,N_17553);
or U18465 (N_18465,N_17501,N_17483);
and U18466 (N_18466,N_17387,N_17590);
and U18467 (N_18467,N_17633,N_17079);
xnor U18468 (N_18468,N_17013,N_17059);
and U18469 (N_18469,N_17769,N_17165);
nor U18470 (N_18470,N_17129,N_17091);
and U18471 (N_18471,N_17405,N_17111);
nand U18472 (N_18472,N_17690,N_17272);
xnor U18473 (N_18473,N_17655,N_17782);
nor U18474 (N_18474,N_17318,N_17365);
nand U18475 (N_18475,N_17484,N_17007);
and U18476 (N_18476,N_17116,N_17758);
nand U18477 (N_18477,N_17785,N_17879);
and U18478 (N_18478,N_17893,N_17680);
and U18479 (N_18479,N_17897,N_17684);
and U18480 (N_18480,N_17636,N_17822);
nor U18481 (N_18481,N_17594,N_17489);
and U18482 (N_18482,N_17652,N_17673);
or U18483 (N_18483,N_17640,N_17699);
nor U18484 (N_18484,N_17791,N_17798);
and U18485 (N_18485,N_17969,N_17610);
nor U18486 (N_18486,N_17612,N_17019);
xnor U18487 (N_18487,N_17163,N_17890);
or U18488 (N_18488,N_17450,N_17671);
nand U18489 (N_18489,N_17224,N_17429);
nor U18490 (N_18490,N_17998,N_17236);
nand U18491 (N_18491,N_17991,N_17746);
and U18492 (N_18492,N_17753,N_17677);
and U18493 (N_18493,N_17221,N_17478);
and U18494 (N_18494,N_17790,N_17559);
xor U18495 (N_18495,N_17806,N_17054);
nand U18496 (N_18496,N_17642,N_17846);
or U18497 (N_18497,N_17167,N_17783);
or U18498 (N_18498,N_17375,N_17390);
nand U18499 (N_18499,N_17715,N_17185);
xor U18500 (N_18500,N_17968,N_17795);
nor U18501 (N_18501,N_17993,N_17099);
nor U18502 (N_18502,N_17360,N_17872);
or U18503 (N_18503,N_17456,N_17887);
nor U18504 (N_18504,N_17318,N_17633);
nand U18505 (N_18505,N_17640,N_17911);
or U18506 (N_18506,N_17415,N_17334);
and U18507 (N_18507,N_17515,N_17176);
nor U18508 (N_18508,N_17627,N_17188);
nor U18509 (N_18509,N_17789,N_17423);
and U18510 (N_18510,N_17871,N_17717);
nor U18511 (N_18511,N_17517,N_17153);
and U18512 (N_18512,N_17040,N_17966);
nor U18513 (N_18513,N_17200,N_17689);
nand U18514 (N_18514,N_17729,N_17905);
nor U18515 (N_18515,N_17814,N_17512);
xnor U18516 (N_18516,N_17375,N_17154);
and U18517 (N_18517,N_17664,N_17085);
xor U18518 (N_18518,N_17175,N_17615);
and U18519 (N_18519,N_17234,N_17382);
xor U18520 (N_18520,N_17246,N_17125);
nor U18521 (N_18521,N_17698,N_17067);
xnor U18522 (N_18522,N_17642,N_17166);
or U18523 (N_18523,N_17547,N_17916);
or U18524 (N_18524,N_17621,N_17671);
xor U18525 (N_18525,N_17856,N_17178);
nand U18526 (N_18526,N_17353,N_17540);
nand U18527 (N_18527,N_17106,N_17885);
nand U18528 (N_18528,N_17280,N_17711);
and U18529 (N_18529,N_17280,N_17618);
xor U18530 (N_18530,N_17318,N_17388);
nor U18531 (N_18531,N_17355,N_17670);
nor U18532 (N_18532,N_17856,N_17394);
and U18533 (N_18533,N_17879,N_17983);
or U18534 (N_18534,N_17252,N_17587);
nand U18535 (N_18535,N_17358,N_17300);
or U18536 (N_18536,N_17667,N_17236);
and U18537 (N_18537,N_17732,N_17885);
xnor U18538 (N_18538,N_17741,N_17328);
nand U18539 (N_18539,N_17126,N_17248);
nor U18540 (N_18540,N_17414,N_17733);
and U18541 (N_18541,N_17223,N_17689);
nor U18542 (N_18542,N_17127,N_17496);
xnor U18543 (N_18543,N_17501,N_17806);
xor U18544 (N_18544,N_17953,N_17348);
nor U18545 (N_18545,N_17347,N_17415);
nand U18546 (N_18546,N_17005,N_17488);
nand U18547 (N_18547,N_17988,N_17900);
nor U18548 (N_18548,N_17615,N_17298);
and U18549 (N_18549,N_17401,N_17648);
or U18550 (N_18550,N_17940,N_17629);
or U18551 (N_18551,N_17714,N_17348);
and U18552 (N_18552,N_17015,N_17384);
nand U18553 (N_18553,N_17400,N_17359);
or U18554 (N_18554,N_17979,N_17142);
xor U18555 (N_18555,N_17790,N_17461);
nand U18556 (N_18556,N_17910,N_17906);
nand U18557 (N_18557,N_17083,N_17331);
or U18558 (N_18558,N_17018,N_17130);
or U18559 (N_18559,N_17150,N_17151);
or U18560 (N_18560,N_17121,N_17983);
xnor U18561 (N_18561,N_17400,N_17392);
xor U18562 (N_18562,N_17834,N_17322);
and U18563 (N_18563,N_17155,N_17790);
nor U18564 (N_18564,N_17216,N_17938);
xnor U18565 (N_18565,N_17388,N_17450);
nand U18566 (N_18566,N_17675,N_17998);
nor U18567 (N_18567,N_17684,N_17756);
nand U18568 (N_18568,N_17099,N_17415);
xnor U18569 (N_18569,N_17291,N_17844);
nand U18570 (N_18570,N_17289,N_17963);
xnor U18571 (N_18571,N_17868,N_17470);
nor U18572 (N_18572,N_17024,N_17241);
or U18573 (N_18573,N_17754,N_17755);
xor U18574 (N_18574,N_17090,N_17473);
or U18575 (N_18575,N_17750,N_17170);
and U18576 (N_18576,N_17875,N_17610);
nand U18577 (N_18577,N_17993,N_17814);
nor U18578 (N_18578,N_17990,N_17794);
and U18579 (N_18579,N_17286,N_17405);
nor U18580 (N_18580,N_17226,N_17928);
or U18581 (N_18581,N_17922,N_17560);
xor U18582 (N_18582,N_17872,N_17764);
or U18583 (N_18583,N_17985,N_17987);
nand U18584 (N_18584,N_17830,N_17770);
and U18585 (N_18585,N_17546,N_17342);
or U18586 (N_18586,N_17282,N_17673);
or U18587 (N_18587,N_17029,N_17736);
and U18588 (N_18588,N_17983,N_17331);
xor U18589 (N_18589,N_17318,N_17237);
nor U18590 (N_18590,N_17698,N_17701);
xor U18591 (N_18591,N_17306,N_17147);
xor U18592 (N_18592,N_17188,N_17739);
and U18593 (N_18593,N_17258,N_17233);
nor U18594 (N_18594,N_17566,N_17252);
nor U18595 (N_18595,N_17085,N_17357);
and U18596 (N_18596,N_17352,N_17885);
and U18597 (N_18597,N_17169,N_17266);
or U18598 (N_18598,N_17801,N_17542);
nor U18599 (N_18599,N_17453,N_17306);
nor U18600 (N_18600,N_17176,N_17424);
xnor U18601 (N_18601,N_17568,N_17417);
nand U18602 (N_18602,N_17320,N_17749);
and U18603 (N_18603,N_17954,N_17389);
and U18604 (N_18604,N_17956,N_17902);
and U18605 (N_18605,N_17827,N_17632);
nor U18606 (N_18606,N_17394,N_17874);
nand U18607 (N_18607,N_17587,N_17443);
and U18608 (N_18608,N_17143,N_17065);
xor U18609 (N_18609,N_17655,N_17717);
xor U18610 (N_18610,N_17878,N_17694);
nor U18611 (N_18611,N_17642,N_17051);
or U18612 (N_18612,N_17527,N_17624);
nand U18613 (N_18613,N_17078,N_17120);
nor U18614 (N_18614,N_17249,N_17628);
or U18615 (N_18615,N_17613,N_17381);
nor U18616 (N_18616,N_17525,N_17559);
nor U18617 (N_18617,N_17623,N_17277);
and U18618 (N_18618,N_17354,N_17636);
nand U18619 (N_18619,N_17708,N_17448);
nor U18620 (N_18620,N_17822,N_17441);
or U18621 (N_18621,N_17763,N_17623);
or U18622 (N_18622,N_17973,N_17204);
nor U18623 (N_18623,N_17260,N_17408);
xnor U18624 (N_18624,N_17879,N_17298);
xor U18625 (N_18625,N_17086,N_17170);
or U18626 (N_18626,N_17345,N_17516);
xor U18627 (N_18627,N_17479,N_17011);
xnor U18628 (N_18628,N_17215,N_17864);
or U18629 (N_18629,N_17311,N_17524);
nand U18630 (N_18630,N_17840,N_17953);
nor U18631 (N_18631,N_17814,N_17910);
and U18632 (N_18632,N_17098,N_17474);
or U18633 (N_18633,N_17751,N_17328);
xnor U18634 (N_18634,N_17327,N_17888);
nor U18635 (N_18635,N_17799,N_17590);
and U18636 (N_18636,N_17716,N_17907);
xor U18637 (N_18637,N_17194,N_17763);
xnor U18638 (N_18638,N_17989,N_17708);
nor U18639 (N_18639,N_17212,N_17975);
nor U18640 (N_18640,N_17201,N_17609);
nand U18641 (N_18641,N_17169,N_17575);
and U18642 (N_18642,N_17056,N_17759);
xnor U18643 (N_18643,N_17001,N_17147);
nand U18644 (N_18644,N_17592,N_17775);
and U18645 (N_18645,N_17083,N_17427);
or U18646 (N_18646,N_17934,N_17575);
and U18647 (N_18647,N_17247,N_17753);
xnor U18648 (N_18648,N_17623,N_17025);
xnor U18649 (N_18649,N_17527,N_17060);
xor U18650 (N_18650,N_17421,N_17201);
and U18651 (N_18651,N_17838,N_17343);
and U18652 (N_18652,N_17966,N_17677);
or U18653 (N_18653,N_17588,N_17636);
nor U18654 (N_18654,N_17213,N_17347);
nor U18655 (N_18655,N_17847,N_17095);
or U18656 (N_18656,N_17315,N_17553);
and U18657 (N_18657,N_17347,N_17292);
nor U18658 (N_18658,N_17374,N_17087);
and U18659 (N_18659,N_17536,N_17709);
xor U18660 (N_18660,N_17993,N_17024);
nand U18661 (N_18661,N_17634,N_17128);
and U18662 (N_18662,N_17817,N_17537);
nand U18663 (N_18663,N_17820,N_17867);
nand U18664 (N_18664,N_17694,N_17116);
nor U18665 (N_18665,N_17958,N_17835);
xnor U18666 (N_18666,N_17983,N_17377);
and U18667 (N_18667,N_17722,N_17554);
nand U18668 (N_18668,N_17744,N_17778);
or U18669 (N_18669,N_17016,N_17735);
xor U18670 (N_18670,N_17431,N_17208);
nor U18671 (N_18671,N_17627,N_17189);
xor U18672 (N_18672,N_17855,N_17075);
xor U18673 (N_18673,N_17752,N_17067);
nor U18674 (N_18674,N_17447,N_17604);
and U18675 (N_18675,N_17684,N_17755);
or U18676 (N_18676,N_17113,N_17875);
xnor U18677 (N_18677,N_17910,N_17802);
nor U18678 (N_18678,N_17042,N_17695);
or U18679 (N_18679,N_17739,N_17523);
nor U18680 (N_18680,N_17708,N_17429);
nor U18681 (N_18681,N_17897,N_17207);
and U18682 (N_18682,N_17370,N_17970);
or U18683 (N_18683,N_17663,N_17444);
nor U18684 (N_18684,N_17706,N_17197);
nand U18685 (N_18685,N_17551,N_17416);
xor U18686 (N_18686,N_17382,N_17583);
nor U18687 (N_18687,N_17580,N_17804);
and U18688 (N_18688,N_17147,N_17722);
or U18689 (N_18689,N_17305,N_17126);
nand U18690 (N_18690,N_17212,N_17814);
and U18691 (N_18691,N_17348,N_17330);
nor U18692 (N_18692,N_17356,N_17353);
nor U18693 (N_18693,N_17663,N_17081);
and U18694 (N_18694,N_17968,N_17202);
and U18695 (N_18695,N_17255,N_17329);
xor U18696 (N_18696,N_17477,N_17008);
and U18697 (N_18697,N_17500,N_17451);
and U18698 (N_18698,N_17960,N_17356);
nand U18699 (N_18699,N_17411,N_17110);
nor U18700 (N_18700,N_17486,N_17745);
nor U18701 (N_18701,N_17405,N_17618);
nor U18702 (N_18702,N_17778,N_17154);
or U18703 (N_18703,N_17922,N_17487);
nand U18704 (N_18704,N_17481,N_17427);
nand U18705 (N_18705,N_17199,N_17936);
or U18706 (N_18706,N_17100,N_17814);
nand U18707 (N_18707,N_17273,N_17503);
or U18708 (N_18708,N_17590,N_17039);
xor U18709 (N_18709,N_17095,N_17089);
nand U18710 (N_18710,N_17518,N_17868);
and U18711 (N_18711,N_17435,N_17206);
nor U18712 (N_18712,N_17084,N_17995);
xor U18713 (N_18713,N_17072,N_17233);
nor U18714 (N_18714,N_17055,N_17908);
or U18715 (N_18715,N_17490,N_17806);
or U18716 (N_18716,N_17039,N_17861);
nor U18717 (N_18717,N_17801,N_17097);
nand U18718 (N_18718,N_17653,N_17577);
nor U18719 (N_18719,N_17789,N_17574);
and U18720 (N_18720,N_17931,N_17968);
xor U18721 (N_18721,N_17649,N_17195);
and U18722 (N_18722,N_17238,N_17243);
nor U18723 (N_18723,N_17650,N_17348);
nor U18724 (N_18724,N_17920,N_17784);
xnor U18725 (N_18725,N_17520,N_17715);
xnor U18726 (N_18726,N_17048,N_17333);
or U18727 (N_18727,N_17779,N_17836);
or U18728 (N_18728,N_17808,N_17844);
nor U18729 (N_18729,N_17082,N_17495);
and U18730 (N_18730,N_17410,N_17211);
nand U18731 (N_18731,N_17133,N_17165);
and U18732 (N_18732,N_17125,N_17039);
nand U18733 (N_18733,N_17641,N_17711);
nand U18734 (N_18734,N_17725,N_17807);
nor U18735 (N_18735,N_17302,N_17693);
xor U18736 (N_18736,N_17784,N_17430);
nand U18737 (N_18737,N_17974,N_17031);
nand U18738 (N_18738,N_17437,N_17187);
or U18739 (N_18739,N_17841,N_17723);
nand U18740 (N_18740,N_17560,N_17337);
xor U18741 (N_18741,N_17087,N_17893);
nand U18742 (N_18742,N_17401,N_17664);
nor U18743 (N_18743,N_17472,N_17337);
and U18744 (N_18744,N_17420,N_17884);
and U18745 (N_18745,N_17093,N_17409);
xnor U18746 (N_18746,N_17137,N_17842);
nand U18747 (N_18747,N_17133,N_17212);
or U18748 (N_18748,N_17482,N_17207);
xnor U18749 (N_18749,N_17020,N_17564);
xor U18750 (N_18750,N_17738,N_17258);
and U18751 (N_18751,N_17577,N_17003);
and U18752 (N_18752,N_17881,N_17433);
nor U18753 (N_18753,N_17783,N_17252);
and U18754 (N_18754,N_17097,N_17174);
nand U18755 (N_18755,N_17978,N_17936);
nor U18756 (N_18756,N_17120,N_17566);
nand U18757 (N_18757,N_17968,N_17373);
nand U18758 (N_18758,N_17846,N_17321);
nor U18759 (N_18759,N_17579,N_17211);
and U18760 (N_18760,N_17572,N_17103);
or U18761 (N_18761,N_17010,N_17402);
xor U18762 (N_18762,N_17220,N_17762);
and U18763 (N_18763,N_17755,N_17855);
or U18764 (N_18764,N_17365,N_17038);
nand U18765 (N_18765,N_17290,N_17525);
nor U18766 (N_18766,N_17348,N_17453);
and U18767 (N_18767,N_17421,N_17764);
nand U18768 (N_18768,N_17630,N_17556);
nand U18769 (N_18769,N_17253,N_17072);
xnor U18770 (N_18770,N_17674,N_17821);
xnor U18771 (N_18771,N_17130,N_17869);
xnor U18772 (N_18772,N_17497,N_17489);
nand U18773 (N_18773,N_17310,N_17608);
xor U18774 (N_18774,N_17644,N_17027);
nand U18775 (N_18775,N_17693,N_17859);
nand U18776 (N_18776,N_17457,N_17840);
nor U18777 (N_18777,N_17020,N_17373);
xnor U18778 (N_18778,N_17382,N_17797);
and U18779 (N_18779,N_17281,N_17870);
nor U18780 (N_18780,N_17729,N_17478);
xor U18781 (N_18781,N_17003,N_17897);
nand U18782 (N_18782,N_17122,N_17484);
xor U18783 (N_18783,N_17829,N_17157);
xor U18784 (N_18784,N_17549,N_17048);
nor U18785 (N_18785,N_17834,N_17069);
xnor U18786 (N_18786,N_17998,N_17004);
nand U18787 (N_18787,N_17778,N_17647);
and U18788 (N_18788,N_17693,N_17840);
or U18789 (N_18789,N_17810,N_17093);
nand U18790 (N_18790,N_17155,N_17572);
nand U18791 (N_18791,N_17035,N_17514);
nor U18792 (N_18792,N_17881,N_17530);
xor U18793 (N_18793,N_17629,N_17016);
xnor U18794 (N_18794,N_17189,N_17216);
xnor U18795 (N_18795,N_17055,N_17096);
xor U18796 (N_18796,N_17683,N_17028);
and U18797 (N_18797,N_17100,N_17796);
and U18798 (N_18798,N_17498,N_17818);
nor U18799 (N_18799,N_17653,N_17572);
xnor U18800 (N_18800,N_17766,N_17806);
nand U18801 (N_18801,N_17477,N_17680);
or U18802 (N_18802,N_17759,N_17108);
and U18803 (N_18803,N_17368,N_17118);
or U18804 (N_18804,N_17236,N_17685);
nor U18805 (N_18805,N_17222,N_17351);
or U18806 (N_18806,N_17639,N_17377);
nand U18807 (N_18807,N_17241,N_17756);
nor U18808 (N_18808,N_17423,N_17257);
nor U18809 (N_18809,N_17856,N_17116);
xnor U18810 (N_18810,N_17631,N_17208);
or U18811 (N_18811,N_17501,N_17355);
xor U18812 (N_18812,N_17247,N_17482);
xor U18813 (N_18813,N_17914,N_17681);
nor U18814 (N_18814,N_17412,N_17481);
xnor U18815 (N_18815,N_17298,N_17481);
or U18816 (N_18816,N_17666,N_17016);
and U18817 (N_18817,N_17856,N_17177);
and U18818 (N_18818,N_17494,N_17964);
nand U18819 (N_18819,N_17546,N_17999);
xor U18820 (N_18820,N_17325,N_17439);
xnor U18821 (N_18821,N_17607,N_17980);
and U18822 (N_18822,N_17283,N_17887);
nand U18823 (N_18823,N_17444,N_17577);
and U18824 (N_18824,N_17420,N_17710);
or U18825 (N_18825,N_17147,N_17801);
or U18826 (N_18826,N_17659,N_17513);
xnor U18827 (N_18827,N_17635,N_17535);
xnor U18828 (N_18828,N_17889,N_17044);
or U18829 (N_18829,N_17562,N_17627);
and U18830 (N_18830,N_17509,N_17823);
nor U18831 (N_18831,N_17370,N_17648);
nor U18832 (N_18832,N_17750,N_17403);
nor U18833 (N_18833,N_17812,N_17294);
and U18834 (N_18834,N_17619,N_17737);
nor U18835 (N_18835,N_17745,N_17528);
nand U18836 (N_18836,N_17354,N_17384);
nand U18837 (N_18837,N_17935,N_17680);
nor U18838 (N_18838,N_17312,N_17790);
xor U18839 (N_18839,N_17845,N_17035);
nor U18840 (N_18840,N_17985,N_17868);
or U18841 (N_18841,N_17878,N_17157);
or U18842 (N_18842,N_17250,N_17679);
nor U18843 (N_18843,N_17346,N_17724);
nand U18844 (N_18844,N_17142,N_17243);
xnor U18845 (N_18845,N_17875,N_17621);
and U18846 (N_18846,N_17476,N_17512);
nand U18847 (N_18847,N_17412,N_17266);
nand U18848 (N_18848,N_17562,N_17603);
xnor U18849 (N_18849,N_17998,N_17764);
nand U18850 (N_18850,N_17850,N_17441);
nand U18851 (N_18851,N_17595,N_17724);
or U18852 (N_18852,N_17727,N_17894);
and U18853 (N_18853,N_17687,N_17315);
nor U18854 (N_18854,N_17387,N_17983);
xnor U18855 (N_18855,N_17456,N_17698);
nand U18856 (N_18856,N_17012,N_17380);
or U18857 (N_18857,N_17004,N_17336);
nand U18858 (N_18858,N_17705,N_17919);
and U18859 (N_18859,N_17857,N_17901);
or U18860 (N_18860,N_17962,N_17155);
xnor U18861 (N_18861,N_17208,N_17212);
nor U18862 (N_18862,N_17848,N_17292);
and U18863 (N_18863,N_17350,N_17983);
and U18864 (N_18864,N_17306,N_17846);
and U18865 (N_18865,N_17217,N_17961);
and U18866 (N_18866,N_17762,N_17735);
nor U18867 (N_18867,N_17310,N_17366);
xor U18868 (N_18868,N_17812,N_17548);
nor U18869 (N_18869,N_17507,N_17052);
or U18870 (N_18870,N_17145,N_17708);
or U18871 (N_18871,N_17134,N_17514);
nor U18872 (N_18872,N_17722,N_17531);
and U18873 (N_18873,N_17987,N_17546);
nor U18874 (N_18874,N_17369,N_17581);
and U18875 (N_18875,N_17039,N_17944);
nor U18876 (N_18876,N_17698,N_17219);
or U18877 (N_18877,N_17537,N_17456);
xnor U18878 (N_18878,N_17132,N_17072);
and U18879 (N_18879,N_17646,N_17389);
xor U18880 (N_18880,N_17947,N_17247);
nand U18881 (N_18881,N_17100,N_17077);
nor U18882 (N_18882,N_17545,N_17249);
and U18883 (N_18883,N_17648,N_17046);
nand U18884 (N_18884,N_17713,N_17800);
xnor U18885 (N_18885,N_17555,N_17326);
xor U18886 (N_18886,N_17634,N_17773);
or U18887 (N_18887,N_17672,N_17019);
and U18888 (N_18888,N_17451,N_17419);
xor U18889 (N_18889,N_17954,N_17160);
nand U18890 (N_18890,N_17856,N_17587);
and U18891 (N_18891,N_17944,N_17962);
nand U18892 (N_18892,N_17381,N_17391);
and U18893 (N_18893,N_17469,N_17899);
xor U18894 (N_18894,N_17334,N_17282);
or U18895 (N_18895,N_17228,N_17108);
and U18896 (N_18896,N_17024,N_17175);
nand U18897 (N_18897,N_17677,N_17269);
nand U18898 (N_18898,N_17169,N_17210);
and U18899 (N_18899,N_17855,N_17825);
or U18900 (N_18900,N_17093,N_17904);
or U18901 (N_18901,N_17822,N_17891);
nor U18902 (N_18902,N_17532,N_17002);
nand U18903 (N_18903,N_17576,N_17770);
xnor U18904 (N_18904,N_17004,N_17598);
and U18905 (N_18905,N_17944,N_17580);
nor U18906 (N_18906,N_17527,N_17361);
or U18907 (N_18907,N_17811,N_17680);
or U18908 (N_18908,N_17318,N_17647);
nand U18909 (N_18909,N_17049,N_17955);
xnor U18910 (N_18910,N_17152,N_17816);
xnor U18911 (N_18911,N_17434,N_17457);
nand U18912 (N_18912,N_17044,N_17735);
xnor U18913 (N_18913,N_17136,N_17234);
nor U18914 (N_18914,N_17483,N_17632);
nor U18915 (N_18915,N_17755,N_17496);
nand U18916 (N_18916,N_17161,N_17256);
and U18917 (N_18917,N_17575,N_17953);
nand U18918 (N_18918,N_17567,N_17003);
xnor U18919 (N_18919,N_17706,N_17400);
and U18920 (N_18920,N_17117,N_17507);
nor U18921 (N_18921,N_17080,N_17974);
or U18922 (N_18922,N_17629,N_17529);
and U18923 (N_18923,N_17958,N_17519);
xor U18924 (N_18924,N_17680,N_17587);
nand U18925 (N_18925,N_17069,N_17434);
or U18926 (N_18926,N_17251,N_17113);
or U18927 (N_18927,N_17919,N_17807);
or U18928 (N_18928,N_17594,N_17139);
xor U18929 (N_18929,N_17644,N_17964);
nor U18930 (N_18930,N_17124,N_17108);
xnor U18931 (N_18931,N_17951,N_17270);
nand U18932 (N_18932,N_17294,N_17431);
and U18933 (N_18933,N_17250,N_17344);
or U18934 (N_18934,N_17616,N_17056);
xnor U18935 (N_18935,N_17880,N_17302);
or U18936 (N_18936,N_17202,N_17527);
nor U18937 (N_18937,N_17789,N_17131);
xor U18938 (N_18938,N_17130,N_17663);
and U18939 (N_18939,N_17891,N_17198);
or U18940 (N_18940,N_17301,N_17730);
or U18941 (N_18941,N_17025,N_17069);
nor U18942 (N_18942,N_17932,N_17003);
nor U18943 (N_18943,N_17660,N_17951);
xor U18944 (N_18944,N_17392,N_17442);
or U18945 (N_18945,N_17231,N_17053);
and U18946 (N_18946,N_17654,N_17668);
nand U18947 (N_18947,N_17096,N_17409);
nor U18948 (N_18948,N_17924,N_17869);
xnor U18949 (N_18949,N_17430,N_17137);
or U18950 (N_18950,N_17356,N_17792);
xnor U18951 (N_18951,N_17282,N_17523);
nor U18952 (N_18952,N_17791,N_17994);
nor U18953 (N_18953,N_17314,N_17231);
nand U18954 (N_18954,N_17506,N_17754);
nand U18955 (N_18955,N_17079,N_17312);
nor U18956 (N_18956,N_17231,N_17168);
xnor U18957 (N_18957,N_17117,N_17207);
xnor U18958 (N_18958,N_17601,N_17479);
or U18959 (N_18959,N_17704,N_17862);
or U18960 (N_18960,N_17192,N_17395);
nand U18961 (N_18961,N_17661,N_17921);
nor U18962 (N_18962,N_17922,N_17142);
xor U18963 (N_18963,N_17505,N_17013);
nor U18964 (N_18964,N_17683,N_17527);
nand U18965 (N_18965,N_17548,N_17220);
and U18966 (N_18966,N_17362,N_17937);
xor U18967 (N_18967,N_17123,N_17969);
or U18968 (N_18968,N_17144,N_17072);
and U18969 (N_18969,N_17081,N_17091);
xnor U18970 (N_18970,N_17514,N_17204);
or U18971 (N_18971,N_17897,N_17020);
nand U18972 (N_18972,N_17006,N_17537);
nor U18973 (N_18973,N_17569,N_17321);
xnor U18974 (N_18974,N_17940,N_17724);
xor U18975 (N_18975,N_17831,N_17981);
nand U18976 (N_18976,N_17823,N_17972);
or U18977 (N_18977,N_17840,N_17640);
or U18978 (N_18978,N_17222,N_17809);
nand U18979 (N_18979,N_17760,N_17714);
nand U18980 (N_18980,N_17650,N_17158);
or U18981 (N_18981,N_17128,N_17302);
xnor U18982 (N_18982,N_17325,N_17551);
xor U18983 (N_18983,N_17001,N_17876);
xor U18984 (N_18984,N_17592,N_17586);
or U18985 (N_18985,N_17438,N_17509);
xor U18986 (N_18986,N_17656,N_17339);
nand U18987 (N_18987,N_17956,N_17915);
nand U18988 (N_18988,N_17430,N_17669);
and U18989 (N_18989,N_17727,N_17327);
nand U18990 (N_18990,N_17574,N_17726);
xor U18991 (N_18991,N_17412,N_17511);
nor U18992 (N_18992,N_17909,N_17369);
xor U18993 (N_18993,N_17285,N_17387);
nor U18994 (N_18994,N_17384,N_17331);
and U18995 (N_18995,N_17661,N_17810);
xor U18996 (N_18996,N_17223,N_17267);
nand U18997 (N_18997,N_17681,N_17282);
and U18998 (N_18998,N_17265,N_17834);
nor U18999 (N_18999,N_17203,N_17503);
nor U19000 (N_19000,N_18000,N_18972);
and U19001 (N_19001,N_18984,N_18467);
xnor U19002 (N_19002,N_18922,N_18331);
nor U19003 (N_19003,N_18745,N_18706);
xnor U19004 (N_19004,N_18412,N_18202);
and U19005 (N_19005,N_18968,N_18668);
or U19006 (N_19006,N_18554,N_18468);
nand U19007 (N_19007,N_18937,N_18788);
nor U19008 (N_19008,N_18075,N_18849);
and U19009 (N_19009,N_18276,N_18287);
nand U19010 (N_19010,N_18621,N_18566);
and U19011 (N_19011,N_18047,N_18766);
and U19012 (N_19012,N_18198,N_18014);
or U19013 (N_19013,N_18609,N_18522);
or U19014 (N_19014,N_18455,N_18438);
nor U19015 (N_19015,N_18956,N_18881);
nor U19016 (N_19016,N_18016,N_18628);
nor U19017 (N_19017,N_18065,N_18663);
nor U19018 (N_19018,N_18058,N_18481);
nand U19019 (N_19019,N_18967,N_18188);
nand U19020 (N_19020,N_18282,N_18400);
or U19021 (N_19021,N_18524,N_18393);
xnor U19022 (N_19022,N_18698,N_18187);
and U19023 (N_19023,N_18818,N_18925);
and U19024 (N_19024,N_18041,N_18503);
nor U19025 (N_19025,N_18839,N_18970);
nor U19026 (N_19026,N_18985,N_18596);
xnor U19027 (N_19027,N_18223,N_18192);
nor U19028 (N_19028,N_18394,N_18551);
nor U19029 (N_19029,N_18595,N_18212);
nand U19030 (N_19030,N_18244,N_18778);
and U19031 (N_19031,N_18130,N_18900);
and U19032 (N_19032,N_18576,N_18491);
xnor U19033 (N_19033,N_18093,N_18804);
and U19034 (N_19034,N_18279,N_18517);
nor U19035 (N_19035,N_18666,N_18251);
xnor U19036 (N_19036,N_18068,N_18339);
xnor U19037 (N_19037,N_18611,N_18946);
xnor U19038 (N_19038,N_18345,N_18141);
nand U19039 (N_19039,N_18962,N_18147);
nand U19040 (N_19040,N_18323,N_18957);
nand U19041 (N_19041,N_18555,N_18919);
or U19042 (N_19042,N_18459,N_18765);
nand U19043 (N_19043,N_18351,N_18040);
nand U19044 (N_19044,N_18843,N_18098);
and U19045 (N_19045,N_18623,N_18873);
xnor U19046 (N_19046,N_18172,N_18820);
or U19047 (N_19047,N_18190,N_18777);
or U19048 (N_19048,N_18505,N_18964);
and U19049 (N_19049,N_18879,N_18631);
nor U19050 (N_19050,N_18506,N_18743);
nor U19051 (N_19051,N_18565,N_18292);
nand U19052 (N_19052,N_18726,N_18911);
nand U19053 (N_19053,N_18164,N_18975);
nor U19054 (N_19054,N_18377,N_18015);
nor U19055 (N_19055,N_18654,N_18070);
and U19056 (N_19056,N_18858,N_18391);
or U19057 (N_19057,N_18862,N_18562);
xor U19058 (N_19058,N_18480,N_18739);
nand U19059 (N_19059,N_18362,N_18694);
or U19060 (N_19060,N_18785,N_18604);
or U19061 (N_19061,N_18906,N_18882);
or U19062 (N_19062,N_18143,N_18240);
nor U19063 (N_19063,N_18994,N_18891);
nor U19064 (N_19064,N_18368,N_18606);
and U19065 (N_19065,N_18886,N_18681);
nand U19066 (N_19066,N_18514,N_18473);
and U19067 (N_19067,N_18857,N_18090);
and U19068 (N_19068,N_18645,N_18527);
and U19069 (N_19069,N_18952,N_18578);
xor U19070 (N_19070,N_18056,N_18178);
nor U19071 (N_19071,N_18655,N_18885);
nand U19072 (N_19072,N_18341,N_18736);
and U19073 (N_19073,N_18215,N_18912);
nor U19074 (N_19074,N_18883,N_18704);
nand U19075 (N_19075,N_18246,N_18308);
nor U19076 (N_19076,N_18544,N_18941);
or U19077 (N_19077,N_18581,N_18415);
or U19078 (N_19078,N_18652,N_18144);
xor U19079 (N_19079,N_18784,N_18594);
nor U19080 (N_19080,N_18634,N_18060);
nand U19081 (N_19081,N_18314,N_18299);
or U19082 (N_19082,N_18929,N_18660);
or U19083 (N_19083,N_18313,N_18507);
or U19084 (N_19084,N_18096,N_18315);
nor U19085 (N_19085,N_18210,N_18475);
xnor U19086 (N_19086,N_18914,N_18490);
nor U19087 (N_19087,N_18974,N_18332);
and U19088 (N_19088,N_18811,N_18186);
nand U19089 (N_19089,N_18081,N_18369);
nor U19090 (N_19090,N_18955,N_18294);
nand U19091 (N_19091,N_18048,N_18763);
or U19092 (N_19092,N_18440,N_18267);
and U19093 (N_19093,N_18028,N_18860);
xnor U19094 (N_19094,N_18918,N_18781);
or U19095 (N_19095,N_18709,N_18958);
nand U19096 (N_19096,N_18521,N_18474);
nor U19097 (N_19097,N_18902,N_18378);
nand U19098 (N_19098,N_18169,N_18328);
nand U19099 (N_19099,N_18568,N_18727);
and U19100 (N_19100,N_18477,N_18520);
and U19101 (N_19101,N_18125,N_18484);
nand U19102 (N_19102,N_18133,N_18277);
or U19103 (N_19103,N_18478,N_18615);
xor U19104 (N_19104,N_18852,N_18034);
xor U19105 (N_19105,N_18350,N_18747);
or U19106 (N_19106,N_18492,N_18532);
or U19107 (N_19107,N_18951,N_18306);
xnor U19108 (N_19108,N_18355,N_18586);
and U19109 (N_19109,N_18176,N_18808);
or U19110 (N_19110,N_18829,N_18095);
xnor U19111 (N_19111,N_18786,N_18538);
nand U19112 (N_19112,N_18513,N_18358);
nor U19113 (N_19113,N_18453,N_18731);
nor U19114 (N_19114,N_18526,N_18079);
nor U19115 (N_19115,N_18884,N_18846);
xnor U19116 (N_19116,N_18089,N_18220);
nor U19117 (N_19117,N_18998,N_18605);
nor U19118 (N_19118,N_18387,N_18120);
nor U19119 (N_19119,N_18838,N_18138);
xnor U19120 (N_19120,N_18311,N_18942);
and U19121 (N_19121,N_18398,N_18775);
nand U19122 (N_19122,N_18441,N_18013);
nor U19123 (N_19123,N_18012,N_18052);
xor U19124 (N_19124,N_18336,N_18653);
xor U19125 (N_19125,N_18003,N_18298);
xnor U19126 (N_19126,N_18278,N_18274);
and U19127 (N_19127,N_18427,N_18257);
and U19128 (N_19128,N_18370,N_18430);
xor U19129 (N_19129,N_18423,N_18866);
and U19130 (N_19130,N_18676,N_18795);
nand U19131 (N_19131,N_18807,N_18979);
xor U19132 (N_19132,N_18115,N_18699);
or U19133 (N_19133,N_18556,N_18221);
or U19134 (N_19134,N_18167,N_18734);
and U19135 (N_19135,N_18559,N_18097);
nor U19136 (N_19136,N_18887,N_18110);
xnor U19137 (N_19137,N_18867,N_18131);
nand U19138 (N_19138,N_18217,N_18191);
nor U19139 (N_19139,N_18717,N_18529);
nor U19140 (N_19140,N_18211,N_18069);
or U19141 (N_19141,N_18247,N_18626);
and U19142 (N_19142,N_18280,N_18632);
xnor U19143 (N_19143,N_18462,N_18153);
nor U19144 (N_19144,N_18017,N_18502);
or U19145 (N_19145,N_18193,N_18563);
nand U19146 (N_19146,N_18949,N_18386);
or U19147 (N_19147,N_18757,N_18152);
or U19148 (N_19148,N_18254,N_18317);
nand U19149 (N_19149,N_18327,N_18738);
nor U19150 (N_19150,N_18755,N_18094);
nand U19151 (N_19151,N_18713,N_18061);
nor U19152 (N_19152,N_18269,N_18037);
or U19153 (N_19153,N_18610,N_18909);
nor U19154 (N_19154,N_18549,N_18410);
and U19155 (N_19155,N_18658,N_18732);
nand U19156 (N_19156,N_18293,N_18241);
and U19157 (N_19157,N_18744,N_18344);
xnor U19158 (N_19158,N_18403,N_18616);
nor U19159 (N_19159,N_18197,N_18696);
nor U19160 (N_19160,N_18402,N_18580);
and U19161 (N_19161,N_18018,N_18712);
and U19162 (N_19162,N_18284,N_18792);
and U19163 (N_19163,N_18534,N_18510);
or U19164 (N_19164,N_18724,N_18817);
or U19165 (N_19165,N_18154,N_18650);
xor U19166 (N_19166,N_18647,N_18026);
and U19167 (N_19167,N_18295,N_18161);
or U19168 (N_19168,N_18206,N_18272);
nand U19169 (N_19169,N_18043,N_18776);
xor U19170 (N_19170,N_18112,N_18685);
and U19171 (N_19171,N_18679,N_18434);
xor U19172 (N_19172,N_18579,N_18286);
and U19173 (N_19173,N_18216,N_18901);
or U19174 (N_19174,N_18961,N_18446);
xnor U19175 (N_19175,N_18536,N_18691);
nor U19176 (N_19176,N_18519,N_18119);
nand U19177 (N_19177,N_18312,N_18102);
xor U19178 (N_19178,N_18950,N_18497);
nand U19179 (N_19179,N_18780,N_18258);
or U19180 (N_19180,N_18155,N_18470);
nand U19181 (N_19181,N_18250,N_18767);
or U19182 (N_19182,N_18714,N_18285);
or U19183 (N_19183,N_18445,N_18460);
xor U19184 (N_19184,N_18450,N_18993);
and U19185 (N_19185,N_18237,N_18051);
or U19186 (N_19186,N_18944,N_18486);
nor U19187 (N_19187,N_18913,N_18334);
and U19188 (N_19188,N_18770,N_18371);
or U19189 (N_19189,N_18988,N_18031);
or U19190 (N_19190,N_18406,N_18960);
nor U19191 (N_19191,N_18592,N_18487);
or U19192 (N_19192,N_18225,N_18337);
or U19193 (N_19193,N_18768,N_18796);
xnor U19194 (N_19194,N_18335,N_18905);
xnor U19195 (N_19195,N_18444,N_18542);
or U19196 (N_19196,N_18598,N_18408);
nor U19197 (N_19197,N_18567,N_18349);
or U19198 (N_19198,N_18092,N_18401);
nor U19199 (N_19199,N_18546,N_18149);
xnor U19200 (N_19200,N_18457,N_18404);
nor U19201 (N_19201,N_18981,N_18124);
and U19202 (N_19202,N_18674,N_18173);
xnor U19203 (N_19203,N_18531,N_18471);
xnor U19204 (N_19204,N_18841,N_18664);
xnor U19205 (N_19205,N_18088,N_18307);
and U19206 (N_19206,N_18528,N_18383);
and U19207 (N_19207,N_18289,N_18201);
xnor U19208 (N_19208,N_18425,N_18813);
or U19209 (N_19209,N_18758,N_18452);
or U19210 (N_19210,N_18232,N_18516);
nor U19211 (N_19211,N_18607,N_18963);
or U19212 (N_19212,N_18413,N_18669);
nor U19213 (N_19213,N_18454,N_18608);
nand U19214 (N_19214,N_18931,N_18570);
or U19215 (N_19215,N_18417,N_18997);
nor U19216 (N_19216,N_18035,N_18023);
nor U19217 (N_19217,N_18910,N_18374);
nand U19218 (N_19218,N_18360,N_18751);
nand U19219 (N_19219,N_18105,N_18865);
nand U19220 (N_19220,N_18501,N_18875);
nor U19221 (N_19221,N_18148,N_18939);
xor U19222 (N_19222,N_18001,N_18690);
nand U19223 (N_19223,N_18924,N_18346);
or U19224 (N_19224,N_18156,N_18890);
nand U19225 (N_19225,N_18903,N_18010);
xnor U19226 (N_19226,N_18118,N_18973);
nand U19227 (N_19227,N_18431,N_18971);
or U19228 (N_19228,N_18730,N_18702);
nand U19229 (N_19229,N_18033,N_18518);
or U19230 (N_19230,N_18671,N_18326);
nand U19231 (N_19231,N_18140,N_18987);
nor U19232 (N_19232,N_18305,N_18500);
nand U19233 (N_19233,N_18723,N_18091);
or U19234 (N_19234,N_18139,N_18597);
nand U19235 (N_19235,N_18659,N_18742);
xnor U19236 (N_19236,N_18195,N_18129);
and U19237 (N_19237,N_18451,N_18205);
and U19238 (N_19238,N_18469,N_18255);
nand U19239 (N_19239,N_18687,N_18179);
or U19240 (N_19240,N_18136,N_18049);
nand U19241 (N_19241,N_18847,N_18703);
or U19242 (N_19242,N_18057,N_18199);
nand U19243 (N_19243,N_18525,N_18101);
or U19244 (N_19244,N_18411,N_18572);
nor U19245 (N_19245,N_18162,N_18259);
xnor U19246 (N_19246,N_18686,N_18587);
and U19247 (N_19247,N_18024,N_18853);
or U19248 (N_19248,N_18100,N_18680);
or U19249 (N_19249,N_18800,N_18376);
and U19250 (N_19250,N_18322,N_18779);
nand U19251 (N_19251,N_18157,N_18230);
nor U19252 (N_19252,N_18617,N_18837);
nand U19253 (N_19253,N_18348,N_18116);
and U19254 (N_19254,N_18835,N_18508);
nand U19255 (N_19255,N_18356,N_18548);
nor U19256 (N_19256,N_18038,N_18045);
nand U19257 (N_19257,N_18256,N_18651);
and U19258 (N_19258,N_18823,N_18281);
and U19259 (N_19259,N_18643,N_18200);
and U19260 (N_19260,N_18810,N_18420);
and U19261 (N_19261,N_18814,N_18801);
and U19262 (N_19262,N_18675,N_18022);
or U19263 (N_19263,N_18488,N_18845);
nand U19264 (N_19264,N_18318,N_18809);
and U19265 (N_19265,N_18086,N_18103);
nor U19266 (N_19266,N_18373,N_18725);
and U19267 (N_19267,N_18329,N_18833);
and U19268 (N_19268,N_18208,N_18228);
nor U19269 (N_19269,N_18999,N_18442);
nand U19270 (N_19270,N_18848,N_18407);
nand U19271 (N_19271,N_18146,N_18002);
nor U19272 (N_19272,N_18564,N_18893);
and U19273 (N_19273,N_18135,N_18389);
xnor U19274 (N_19274,N_18177,N_18443);
or U19275 (N_19275,N_18347,N_18180);
xnor U19276 (N_19276,N_18657,N_18812);
nand U19277 (N_19277,N_18824,N_18803);
or U19278 (N_19278,N_18614,N_18271);
or U19279 (N_19279,N_18983,N_18359);
xnor U19280 (N_19280,N_18137,N_18573);
nand U19281 (N_19281,N_18343,N_18877);
and U19282 (N_19282,N_18978,N_18831);
nor U19283 (N_19283,N_18209,N_18575);
or U19284 (N_19284,N_18082,N_18711);
xor U19285 (N_19285,N_18871,N_18080);
xor U19286 (N_19286,N_18384,N_18071);
xnor U19287 (N_19287,N_18769,N_18266);
nor U19288 (N_19288,N_18923,N_18150);
xor U19289 (N_19289,N_18435,N_18753);
and U19290 (N_19290,N_18249,N_18752);
and U19291 (N_19291,N_18476,N_18930);
nand U19292 (N_19292,N_18027,N_18264);
xor U19293 (N_19293,N_18721,N_18793);
nor U19294 (N_19294,N_18619,N_18301);
nor U19295 (N_19295,N_18077,N_18283);
nor U19296 (N_19296,N_18625,N_18053);
or U19297 (N_19297,N_18561,N_18718);
nand U19298 (N_19298,N_18541,N_18330);
or U19299 (N_19299,N_18361,N_18005);
nor U19300 (N_19300,N_18908,N_18342);
or U19301 (N_19301,N_18512,N_18722);
xnor U19302 (N_19302,N_18449,N_18990);
nor U19303 (N_19303,N_18836,N_18036);
nand U19304 (N_19304,N_18482,N_18165);
xor U19305 (N_19305,N_18122,N_18969);
nor U19306 (N_19306,N_18636,N_18772);
xnor U19307 (N_19307,N_18218,N_18224);
nand U19308 (N_19308,N_18708,N_18754);
or U19309 (N_19309,N_18108,N_18692);
xnor U19310 (N_19310,N_18644,N_18134);
or U19311 (N_19311,N_18265,N_18109);
nor U19312 (N_19312,N_18290,N_18850);
nor U19313 (N_19313,N_18456,N_18380);
or U19314 (N_19314,N_18158,N_18543);
xor U19315 (N_19315,N_18021,N_18828);
nor U19316 (N_19316,N_18499,N_18683);
or U19317 (N_19317,N_18637,N_18799);
and U19318 (N_19318,N_18791,N_18953);
and U19319 (N_19319,N_18114,N_18733);
or U19320 (N_19320,N_18688,N_18085);
or U19321 (N_19321,N_18288,N_18340);
nor U19322 (N_19322,N_18006,N_18854);
nand U19323 (N_19323,N_18054,N_18421);
and U19324 (N_19324,N_18750,N_18011);
xnor U19325 (N_19325,N_18270,N_18855);
nor U19326 (N_19326,N_18707,N_18117);
or U19327 (N_19327,N_18934,N_18560);
and U19328 (N_19328,N_18511,N_18163);
nand U19329 (N_19329,N_18868,N_18620);
nand U19330 (N_19330,N_18365,N_18840);
nor U19331 (N_19331,N_18458,N_18557);
and U19332 (N_19332,N_18325,N_18989);
xnor U19333 (N_19333,N_18126,N_18066);
xor U19334 (N_19334,N_18748,N_18214);
xor U19335 (N_19335,N_18509,N_18170);
nor U19336 (N_19336,N_18142,N_18826);
or U19337 (N_19337,N_18168,N_18789);
nand U19338 (N_19338,N_18219,N_18261);
nor U19339 (N_19339,N_18782,N_18976);
xor U19340 (N_19340,N_18494,N_18864);
nand U19341 (N_19341,N_18405,N_18710);
nor U19342 (N_19342,N_18062,N_18007);
nor U19343 (N_19343,N_18869,N_18805);
or U19344 (N_19344,N_18695,N_18189);
and U19345 (N_19345,N_18333,N_18907);
nor U19346 (N_19346,N_18665,N_18539);
xnor U19347 (N_19347,N_18309,N_18055);
or U19348 (N_19348,N_18667,N_18310);
nor U19349 (N_19349,N_18959,N_18720);
and U19350 (N_19350,N_18992,N_18464);
xor U19351 (N_19351,N_18547,N_18029);
and U19352 (N_19352,N_18275,N_18545);
nor U19353 (N_19353,N_18390,N_18078);
nor U19354 (N_19354,N_18773,N_18633);
nand U19355 (N_19355,N_18926,N_18856);
xor U19356 (N_19356,N_18428,N_18316);
and U19357 (N_19357,N_18947,N_18716);
or U19358 (N_19358,N_18363,N_18977);
nand U19359 (N_19359,N_18297,N_18104);
nor U19360 (N_19360,N_18830,N_18461);
and U19361 (N_19361,N_18815,N_18059);
or U19362 (N_19362,N_18050,N_18612);
nand U19363 (N_19363,N_18904,N_18042);
and U19364 (N_19364,N_18426,N_18945);
and U19365 (N_19365,N_18338,N_18008);
nor U19366 (N_19366,N_18375,N_18319);
or U19367 (N_19367,N_18182,N_18046);
xnor U19368 (N_19368,N_18185,N_18489);
nor U19369 (N_19369,N_18196,N_18762);
and U19370 (N_19370,N_18399,N_18472);
xnor U19371 (N_19371,N_18746,N_18515);
nand U19372 (N_19372,N_18876,N_18954);
or U19373 (N_19373,N_18072,N_18844);
xnor U19374 (N_19374,N_18759,N_18263);
xnor U19375 (N_19375,N_18966,N_18927);
nor U19376 (N_19376,N_18030,N_18203);
and U19377 (N_19377,N_18737,N_18673);
nand U19378 (N_19378,N_18076,N_18935);
or U19379 (N_19379,N_18385,N_18728);
xnor U19380 (N_19380,N_18656,N_18463);
nand U19381 (N_19381,N_18729,N_18273);
xor U19382 (N_19382,N_18419,N_18429);
xnor U19383 (N_19383,N_18802,N_18790);
xnor U19384 (N_19384,N_18895,N_18174);
nand U19385 (N_19385,N_18917,N_18677);
nor U19386 (N_19386,N_18019,N_18638);
or U19387 (N_19387,N_18253,N_18825);
xnor U19388 (N_19388,N_18236,N_18583);
and U19389 (N_19389,N_18422,N_18416);
and U19390 (N_19390,N_18083,N_18107);
xnor U19391 (N_19391,N_18321,N_18819);
nand U19392 (N_19392,N_18291,N_18433);
and U19393 (N_19393,N_18151,N_18550);
nand U19394 (N_19394,N_18248,N_18466);
nand U19395 (N_19395,N_18889,N_18483);
nand U19396 (N_19396,N_18268,N_18649);
xnor U19397 (N_19397,N_18320,N_18588);
or U19398 (N_19398,N_18396,N_18213);
nand U19399 (N_19399,N_18584,N_18372);
and U19400 (N_19400,N_18670,N_18872);
and U19401 (N_19401,N_18700,N_18235);
nand U19402 (N_19402,N_18798,N_18234);
xor U19403 (N_19403,N_18558,N_18175);
nand U19404 (N_19404,N_18437,N_18648);
and U19405 (N_19405,N_18227,N_18447);
xnor U19406 (N_19406,N_18245,N_18569);
nand U19407 (N_19407,N_18063,N_18127);
or U19408 (N_19408,N_18222,N_18366);
or U19409 (N_19409,N_18231,N_18204);
or U19410 (N_19410,N_18894,N_18646);
or U19411 (N_19411,N_18132,N_18303);
nand U19412 (N_19412,N_18599,N_18498);
or U19413 (N_19413,N_18834,N_18921);
or U19414 (N_19414,N_18601,N_18540);
or U19415 (N_19415,N_18300,N_18641);
and U19416 (N_19416,N_18020,N_18113);
and U19417 (N_19417,N_18920,N_18530);
nor U19418 (N_19418,N_18392,N_18689);
nor U19419 (N_19419,N_18899,N_18642);
nand U19420 (N_19420,N_18980,N_18128);
and U19421 (N_19421,N_18493,N_18896);
or U19422 (N_19422,N_18794,N_18194);
or U19423 (N_19423,N_18705,N_18160);
xnor U19424 (N_19424,N_18627,N_18701);
or U19425 (N_19425,N_18639,N_18874);
nand U19426 (N_19426,N_18936,N_18661);
xor U19427 (N_19427,N_18603,N_18354);
and U19428 (N_19428,N_18774,N_18229);
xor U19429 (N_19429,N_18171,N_18044);
nand U19430 (N_19430,N_18262,N_18418);
and U19431 (N_19431,N_18986,N_18948);
nand U19432 (N_19432,N_18892,N_18682);
nor U19433 (N_19433,N_18982,N_18485);
and U19434 (N_19434,N_18496,N_18409);
or U19435 (N_19435,N_18898,N_18740);
or U19436 (N_19436,N_18996,N_18537);
nor U19437 (N_19437,N_18448,N_18302);
or U19438 (N_19438,N_18367,N_18870);
nand U19439 (N_19439,N_18395,N_18861);
or U19440 (N_19440,N_18571,N_18039);
nor U19441 (N_19441,N_18357,N_18123);
and U19442 (N_19442,N_18574,N_18940);
xnor U19443 (N_19443,N_18760,N_18741);
and U19444 (N_19444,N_18073,N_18589);
nor U19445 (N_19445,N_18239,N_18859);
and U19446 (N_19446,N_18381,N_18535);
xnor U19447 (N_19447,N_18851,N_18629);
xnor U19448 (N_19448,N_18121,N_18414);
or U19449 (N_19449,N_18379,N_18106);
nor U19450 (N_19450,N_18624,N_18943);
or U19451 (N_19451,N_18916,N_18684);
and U19452 (N_19452,N_18938,N_18087);
nor U19453 (N_19453,N_18523,N_18252);
nor U19454 (N_19454,N_18397,N_18697);
nor U19455 (N_19455,N_18099,N_18436);
nand U19456 (N_19456,N_18915,N_18324);
or U19457 (N_19457,N_18243,N_18928);
xnor U19458 (N_19458,N_18166,N_18424);
nand U19459 (N_19459,N_18635,N_18897);
nor U19460 (N_19460,N_18593,N_18353);
or U19461 (N_19461,N_18630,N_18756);
or U19462 (N_19462,N_18577,N_18145);
or U19463 (N_19463,N_18111,N_18465);
or U19464 (N_19464,N_18552,N_18821);
xnor U19465 (N_19465,N_18184,N_18304);
nor U19466 (N_19466,N_18600,N_18591);
and U19467 (N_19467,N_18025,N_18832);
nor U19468 (N_19468,N_18064,N_18827);
nor U19469 (N_19469,N_18074,N_18032);
or U19470 (N_19470,N_18888,N_18806);
nand U19471 (N_19471,N_18764,N_18693);
nor U19472 (N_19472,N_18933,N_18432);
nand U19473 (N_19473,N_18602,N_18504);
nand U19474 (N_19474,N_18797,N_18715);
or U19475 (N_19475,N_18816,N_18352);
or U19476 (N_19476,N_18965,N_18613);
or U19477 (N_19477,N_18735,N_18880);
xor U19478 (N_19478,N_18585,N_18238);
or U19479 (N_19479,N_18260,N_18479);
and U19480 (N_19480,N_18207,N_18233);
nor U19481 (N_19481,N_18364,N_18822);
or U19482 (N_19482,N_18382,N_18084);
or U19483 (N_19483,N_18783,N_18878);
and U19484 (N_19484,N_18582,N_18662);
nor U19485 (N_19485,N_18067,N_18761);
or U19486 (N_19486,N_18181,N_18590);
and U19487 (N_19487,N_18771,N_18553);
xnor U19488 (N_19488,N_18226,N_18863);
xnor U19489 (N_19489,N_18622,N_18618);
nor U19490 (N_19490,N_18678,N_18495);
or U19491 (N_19491,N_18842,N_18749);
nor U19492 (N_19492,N_18183,N_18242);
xnor U19493 (N_19493,N_18533,N_18009);
and U19494 (N_19494,N_18932,N_18296);
xnor U19495 (N_19495,N_18719,N_18388);
nor U19496 (N_19496,N_18640,N_18787);
xnor U19497 (N_19497,N_18991,N_18159);
xnor U19498 (N_19498,N_18672,N_18439);
or U19499 (N_19499,N_18004,N_18995);
nor U19500 (N_19500,N_18814,N_18670);
xnor U19501 (N_19501,N_18250,N_18359);
nor U19502 (N_19502,N_18018,N_18582);
nand U19503 (N_19503,N_18952,N_18257);
nand U19504 (N_19504,N_18477,N_18892);
nor U19505 (N_19505,N_18279,N_18459);
and U19506 (N_19506,N_18161,N_18263);
xnor U19507 (N_19507,N_18356,N_18785);
nand U19508 (N_19508,N_18211,N_18941);
and U19509 (N_19509,N_18271,N_18321);
and U19510 (N_19510,N_18525,N_18126);
nor U19511 (N_19511,N_18796,N_18606);
nand U19512 (N_19512,N_18160,N_18784);
and U19513 (N_19513,N_18587,N_18221);
and U19514 (N_19514,N_18833,N_18692);
nand U19515 (N_19515,N_18209,N_18655);
nor U19516 (N_19516,N_18611,N_18092);
and U19517 (N_19517,N_18982,N_18527);
nor U19518 (N_19518,N_18625,N_18634);
xnor U19519 (N_19519,N_18134,N_18131);
or U19520 (N_19520,N_18158,N_18723);
nand U19521 (N_19521,N_18105,N_18641);
nand U19522 (N_19522,N_18719,N_18034);
nor U19523 (N_19523,N_18903,N_18260);
or U19524 (N_19524,N_18341,N_18794);
xor U19525 (N_19525,N_18883,N_18456);
xor U19526 (N_19526,N_18828,N_18197);
or U19527 (N_19527,N_18742,N_18771);
xnor U19528 (N_19528,N_18047,N_18050);
xor U19529 (N_19529,N_18220,N_18087);
nor U19530 (N_19530,N_18987,N_18622);
xnor U19531 (N_19531,N_18144,N_18001);
and U19532 (N_19532,N_18791,N_18902);
or U19533 (N_19533,N_18719,N_18844);
or U19534 (N_19534,N_18141,N_18752);
or U19535 (N_19535,N_18135,N_18378);
and U19536 (N_19536,N_18119,N_18419);
xor U19537 (N_19537,N_18314,N_18768);
nand U19538 (N_19538,N_18550,N_18852);
xnor U19539 (N_19539,N_18605,N_18258);
or U19540 (N_19540,N_18993,N_18731);
nor U19541 (N_19541,N_18063,N_18326);
or U19542 (N_19542,N_18897,N_18032);
and U19543 (N_19543,N_18084,N_18110);
and U19544 (N_19544,N_18909,N_18961);
nand U19545 (N_19545,N_18790,N_18230);
nor U19546 (N_19546,N_18951,N_18751);
and U19547 (N_19547,N_18472,N_18594);
or U19548 (N_19548,N_18138,N_18135);
or U19549 (N_19549,N_18046,N_18555);
xor U19550 (N_19550,N_18424,N_18961);
nor U19551 (N_19551,N_18503,N_18904);
nand U19552 (N_19552,N_18434,N_18061);
nand U19553 (N_19553,N_18594,N_18877);
nor U19554 (N_19554,N_18684,N_18319);
nand U19555 (N_19555,N_18923,N_18838);
nand U19556 (N_19556,N_18647,N_18770);
and U19557 (N_19557,N_18280,N_18069);
nand U19558 (N_19558,N_18722,N_18522);
xnor U19559 (N_19559,N_18125,N_18230);
xor U19560 (N_19560,N_18604,N_18141);
nor U19561 (N_19561,N_18371,N_18897);
xor U19562 (N_19562,N_18867,N_18680);
xnor U19563 (N_19563,N_18093,N_18160);
and U19564 (N_19564,N_18014,N_18329);
nor U19565 (N_19565,N_18976,N_18023);
xnor U19566 (N_19566,N_18121,N_18367);
nor U19567 (N_19567,N_18888,N_18554);
xor U19568 (N_19568,N_18502,N_18471);
nand U19569 (N_19569,N_18323,N_18601);
nand U19570 (N_19570,N_18150,N_18388);
nand U19571 (N_19571,N_18305,N_18215);
nand U19572 (N_19572,N_18650,N_18477);
nor U19573 (N_19573,N_18906,N_18113);
nand U19574 (N_19574,N_18333,N_18115);
xnor U19575 (N_19575,N_18442,N_18567);
xor U19576 (N_19576,N_18681,N_18633);
nor U19577 (N_19577,N_18022,N_18411);
xor U19578 (N_19578,N_18467,N_18337);
or U19579 (N_19579,N_18476,N_18456);
or U19580 (N_19580,N_18799,N_18628);
and U19581 (N_19581,N_18514,N_18764);
and U19582 (N_19582,N_18505,N_18710);
nand U19583 (N_19583,N_18940,N_18384);
and U19584 (N_19584,N_18044,N_18639);
nand U19585 (N_19585,N_18034,N_18077);
nand U19586 (N_19586,N_18242,N_18682);
or U19587 (N_19587,N_18914,N_18091);
and U19588 (N_19588,N_18497,N_18032);
xnor U19589 (N_19589,N_18982,N_18736);
nand U19590 (N_19590,N_18081,N_18888);
or U19591 (N_19591,N_18489,N_18220);
and U19592 (N_19592,N_18682,N_18503);
nor U19593 (N_19593,N_18748,N_18589);
and U19594 (N_19594,N_18410,N_18936);
nand U19595 (N_19595,N_18524,N_18313);
nand U19596 (N_19596,N_18998,N_18844);
and U19597 (N_19597,N_18970,N_18406);
nand U19598 (N_19598,N_18841,N_18200);
nor U19599 (N_19599,N_18665,N_18814);
nor U19600 (N_19600,N_18448,N_18541);
nor U19601 (N_19601,N_18612,N_18487);
nor U19602 (N_19602,N_18987,N_18938);
and U19603 (N_19603,N_18119,N_18897);
nand U19604 (N_19604,N_18716,N_18394);
or U19605 (N_19605,N_18924,N_18269);
nor U19606 (N_19606,N_18940,N_18761);
nand U19607 (N_19607,N_18196,N_18217);
xnor U19608 (N_19608,N_18598,N_18782);
or U19609 (N_19609,N_18640,N_18639);
or U19610 (N_19610,N_18377,N_18523);
nor U19611 (N_19611,N_18338,N_18855);
xor U19612 (N_19612,N_18733,N_18983);
and U19613 (N_19613,N_18086,N_18455);
xnor U19614 (N_19614,N_18779,N_18931);
nand U19615 (N_19615,N_18377,N_18271);
or U19616 (N_19616,N_18006,N_18962);
or U19617 (N_19617,N_18894,N_18326);
and U19618 (N_19618,N_18181,N_18842);
xor U19619 (N_19619,N_18738,N_18645);
nor U19620 (N_19620,N_18489,N_18819);
xnor U19621 (N_19621,N_18893,N_18973);
and U19622 (N_19622,N_18368,N_18646);
nand U19623 (N_19623,N_18513,N_18636);
nor U19624 (N_19624,N_18045,N_18471);
xor U19625 (N_19625,N_18410,N_18827);
or U19626 (N_19626,N_18514,N_18986);
and U19627 (N_19627,N_18872,N_18947);
xor U19628 (N_19628,N_18830,N_18584);
nand U19629 (N_19629,N_18733,N_18195);
or U19630 (N_19630,N_18967,N_18576);
or U19631 (N_19631,N_18858,N_18290);
nor U19632 (N_19632,N_18906,N_18533);
nor U19633 (N_19633,N_18482,N_18285);
and U19634 (N_19634,N_18937,N_18302);
nor U19635 (N_19635,N_18336,N_18527);
and U19636 (N_19636,N_18480,N_18592);
nand U19637 (N_19637,N_18158,N_18573);
or U19638 (N_19638,N_18736,N_18675);
or U19639 (N_19639,N_18295,N_18701);
xor U19640 (N_19640,N_18403,N_18854);
or U19641 (N_19641,N_18996,N_18603);
nand U19642 (N_19642,N_18232,N_18605);
nor U19643 (N_19643,N_18663,N_18368);
or U19644 (N_19644,N_18583,N_18832);
nor U19645 (N_19645,N_18691,N_18235);
xnor U19646 (N_19646,N_18178,N_18550);
nand U19647 (N_19647,N_18547,N_18104);
nor U19648 (N_19648,N_18605,N_18618);
nand U19649 (N_19649,N_18220,N_18966);
xnor U19650 (N_19650,N_18246,N_18437);
nand U19651 (N_19651,N_18261,N_18046);
xor U19652 (N_19652,N_18913,N_18627);
nand U19653 (N_19653,N_18460,N_18842);
or U19654 (N_19654,N_18996,N_18107);
or U19655 (N_19655,N_18296,N_18788);
nor U19656 (N_19656,N_18205,N_18063);
and U19657 (N_19657,N_18441,N_18140);
nand U19658 (N_19658,N_18150,N_18417);
or U19659 (N_19659,N_18776,N_18508);
or U19660 (N_19660,N_18525,N_18790);
or U19661 (N_19661,N_18834,N_18039);
nor U19662 (N_19662,N_18888,N_18279);
xor U19663 (N_19663,N_18900,N_18405);
xor U19664 (N_19664,N_18887,N_18913);
xnor U19665 (N_19665,N_18301,N_18001);
nand U19666 (N_19666,N_18589,N_18763);
nor U19667 (N_19667,N_18344,N_18709);
or U19668 (N_19668,N_18983,N_18071);
or U19669 (N_19669,N_18662,N_18317);
nor U19670 (N_19670,N_18280,N_18845);
nor U19671 (N_19671,N_18957,N_18518);
or U19672 (N_19672,N_18738,N_18723);
and U19673 (N_19673,N_18501,N_18717);
nor U19674 (N_19674,N_18325,N_18209);
nand U19675 (N_19675,N_18442,N_18441);
or U19676 (N_19676,N_18382,N_18194);
xnor U19677 (N_19677,N_18816,N_18249);
or U19678 (N_19678,N_18599,N_18794);
and U19679 (N_19679,N_18890,N_18007);
nand U19680 (N_19680,N_18790,N_18680);
or U19681 (N_19681,N_18370,N_18712);
and U19682 (N_19682,N_18836,N_18096);
nor U19683 (N_19683,N_18246,N_18374);
nor U19684 (N_19684,N_18871,N_18786);
and U19685 (N_19685,N_18876,N_18953);
nor U19686 (N_19686,N_18441,N_18312);
nor U19687 (N_19687,N_18164,N_18432);
xor U19688 (N_19688,N_18734,N_18556);
or U19689 (N_19689,N_18042,N_18440);
or U19690 (N_19690,N_18055,N_18840);
or U19691 (N_19691,N_18655,N_18182);
nand U19692 (N_19692,N_18053,N_18476);
or U19693 (N_19693,N_18278,N_18026);
nor U19694 (N_19694,N_18428,N_18932);
xnor U19695 (N_19695,N_18318,N_18508);
nand U19696 (N_19696,N_18632,N_18381);
and U19697 (N_19697,N_18023,N_18911);
nand U19698 (N_19698,N_18619,N_18815);
nand U19699 (N_19699,N_18682,N_18215);
nor U19700 (N_19700,N_18723,N_18803);
and U19701 (N_19701,N_18387,N_18777);
nor U19702 (N_19702,N_18524,N_18101);
or U19703 (N_19703,N_18832,N_18193);
nor U19704 (N_19704,N_18629,N_18759);
or U19705 (N_19705,N_18221,N_18263);
nand U19706 (N_19706,N_18400,N_18395);
nor U19707 (N_19707,N_18502,N_18926);
nand U19708 (N_19708,N_18836,N_18411);
xor U19709 (N_19709,N_18069,N_18170);
and U19710 (N_19710,N_18896,N_18966);
nor U19711 (N_19711,N_18072,N_18857);
xor U19712 (N_19712,N_18401,N_18271);
or U19713 (N_19713,N_18146,N_18648);
xnor U19714 (N_19714,N_18051,N_18263);
and U19715 (N_19715,N_18440,N_18113);
nor U19716 (N_19716,N_18854,N_18499);
or U19717 (N_19717,N_18608,N_18558);
nor U19718 (N_19718,N_18182,N_18349);
nor U19719 (N_19719,N_18283,N_18781);
and U19720 (N_19720,N_18336,N_18141);
nor U19721 (N_19721,N_18982,N_18508);
nand U19722 (N_19722,N_18651,N_18599);
xor U19723 (N_19723,N_18590,N_18853);
and U19724 (N_19724,N_18193,N_18210);
nand U19725 (N_19725,N_18689,N_18028);
nor U19726 (N_19726,N_18316,N_18775);
nor U19727 (N_19727,N_18658,N_18652);
nor U19728 (N_19728,N_18923,N_18718);
nor U19729 (N_19729,N_18859,N_18763);
xnor U19730 (N_19730,N_18886,N_18585);
and U19731 (N_19731,N_18856,N_18567);
xnor U19732 (N_19732,N_18600,N_18771);
nand U19733 (N_19733,N_18864,N_18621);
xor U19734 (N_19734,N_18076,N_18890);
nor U19735 (N_19735,N_18600,N_18413);
nand U19736 (N_19736,N_18756,N_18475);
nor U19737 (N_19737,N_18299,N_18220);
nand U19738 (N_19738,N_18542,N_18056);
or U19739 (N_19739,N_18949,N_18260);
nor U19740 (N_19740,N_18305,N_18882);
nand U19741 (N_19741,N_18908,N_18460);
xor U19742 (N_19742,N_18816,N_18231);
xor U19743 (N_19743,N_18272,N_18201);
xnor U19744 (N_19744,N_18796,N_18586);
or U19745 (N_19745,N_18732,N_18847);
nor U19746 (N_19746,N_18763,N_18390);
nor U19747 (N_19747,N_18928,N_18930);
and U19748 (N_19748,N_18726,N_18495);
nor U19749 (N_19749,N_18956,N_18404);
xor U19750 (N_19750,N_18173,N_18410);
nand U19751 (N_19751,N_18295,N_18885);
nand U19752 (N_19752,N_18689,N_18787);
nor U19753 (N_19753,N_18655,N_18878);
xnor U19754 (N_19754,N_18460,N_18151);
nand U19755 (N_19755,N_18555,N_18022);
or U19756 (N_19756,N_18815,N_18553);
and U19757 (N_19757,N_18020,N_18341);
and U19758 (N_19758,N_18786,N_18898);
and U19759 (N_19759,N_18473,N_18095);
nor U19760 (N_19760,N_18612,N_18155);
xor U19761 (N_19761,N_18194,N_18811);
xor U19762 (N_19762,N_18074,N_18360);
or U19763 (N_19763,N_18450,N_18841);
and U19764 (N_19764,N_18889,N_18071);
nand U19765 (N_19765,N_18612,N_18280);
or U19766 (N_19766,N_18075,N_18258);
xnor U19767 (N_19767,N_18950,N_18085);
and U19768 (N_19768,N_18377,N_18155);
nand U19769 (N_19769,N_18291,N_18995);
and U19770 (N_19770,N_18664,N_18503);
and U19771 (N_19771,N_18558,N_18647);
and U19772 (N_19772,N_18057,N_18854);
nand U19773 (N_19773,N_18629,N_18588);
nand U19774 (N_19774,N_18479,N_18389);
or U19775 (N_19775,N_18686,N_18898);
nand U19776 (N_19776,N_18872,N_18605);
xor U19777 (N_19777,N_18215,N_18210);
nand U19778 (N_19778,N_18991,N_18196);
and U19779 (N_19779,N_18749,N_18832);
nor U19780 (N_19780,N_18805,N_18725);
xor U19781 (N_19781,N_18650,N_18248);
xnor U19782 (N_19782,N_18196,N_18192);
xnor U19783 (N_19783,N_18686,N_18940);
and U19784 (N_19784,N_18892,N_18709);
nand U19785 (N_19785,N_18957,N_18234);
xnor U19786 (N_19786,N_18488,N_18045);
xor U19787 (N_19787,N_18236,N_18981);
nor U19788 (N_19788,N_18884,N_18892);
xor U19789 (N_19789,N_18407,N_18350);
and U19790 (N_19790,N_18363,N_18527);
nor U19791 (N_19791,N_18069,N_18155);
nor U19792 (N_19792,N_18844,N_18101);
and U19793 (N_19793,N_18515,N_18308);
xnor U19794 (N_19794,N_18191,N_18117);
and U19795 (N_19795,N_18975,N_18671);
nor U19796 (N_19796,N_18869,N_18686);
xor U19797 (N_19797,N_18856,N_18399);
or U19798 (N_19798,N_18949,N_18667);
nand U19799 (N_19799,N_18201,N_18479);
xor U19800 (N_19800,N_18743,N_18349);
and U19801 (N_19801,N_18307,N_18989);
xnor U19802 (N_19802,N_18870,N_18827);
nor U19803 (N_19803,N_18789,N_18849);
and U19804 (N_19804,N_18983,N_18047);
nand U19805 (N_19805,N_18021,N_18294);
xnor U19806 (N_19806,N_18446,N_18409);
and U19807 (N_19807,N_18242,N_18099);
nand U19808 (N_19808,N_18023,N_18076);
nor U19809 (N_19809,N_18474,N_18703);
xor U19810 (N_19810,N_18366,N_18937);
nor U19811 (N_19811,N_18926,N_18111);
nor U19812 (N_19812,N_18595,N_18244);
xor U19813 (N_19813,N_18039,N_18920);
nor U19814 (N_19814,N_18129,N_18440);
and U19815 (N_19815,N_18300,N_18621);
nor U19816 (N_19816,N_18510,N_18907);
or U19817 (N_19817,N_18876,N_18355);
or U19818 (N_19818,N_18888,N_18836);
nor U19819 (N_19819,N_18311,N_18566);
and U19820 (N_19820,N_18862,N_18864);
xnor U19821 (N_19821,N_18779,N_18352);
nor U19822 (N_19822,N_18025,N_18603);
or U19823 (N_19823,N_18204,N_18924);
and U19824 (N_19824,N_18777,N_18048);
nor U19825 (N_19825,N_18389,N_18301);
nand U19826 (N_19826,N_18965,N_18129);
or U19827 (N_19827,N_18853,N_18689);
xnor U19828 (N_19828,N_18750,N_18106);
xor U19829 (N_19829,N_18075,N_18370);
and U19830 (N_19830,N_18486,N_18143);
or U19831 (N_19831,N_18608,N_18613);
nand U19832 (N_19832,N_18534,N_18200);
or U19833 (N_19833,N_18740,N_18141);
or U19834 (N_19834,N_18901,N_18255);
xor U19835 (N_19835,N_18188,N_18070);
nor U19836 (N_19836,N_18934,N_18321);
and U19837 (N_19837,N_18058,N_18625);
or U19838 (N_19838,N_18727,N_18163);
or U19839 (N_19839,N_18127,N_18506);
and U19840 (N_19840,N_18559,N_18252);
and U19841 (N_19841,N_18233,N_18177);
nor U19842 (N_19842,N_18583,N_18295);
nand U19843 (N_19843,N_18452,N_18787);
nor U19844 (N_19844,N_18947,N_18370);
and U19845 (N_19845,N_18710,N_18230);
xor U19846 (N_19846,N_18543,N_18652);
xor U19847 (N_19847,N_18584,N_18349);
xor U19848 (N_19848,N_18830,N_18565);
or U19849 (N_19849,N_18076,N_18769);
xnor U19850 (N_19850,N_18110,N_18947);
and U19851 (N_19851,N_18111,N_18368);
and U19852 (N_19852,N_18172,N_18879);
and U19853 (N_19853,N_18864,N_18922);
and U19854 (N_19854,N_18229,N_18816);
or U19855 (N_19855,N_18482,N_18976);
nand U19856 (N_19856,N_18716,N_18853);
or U19857 (N_19857,N_18771,N_18666);
nand U19858 (N_19858,N_18597,N_18456);
nand U19859 (N_19859,N_18627,N_18526);
nor U19860 (N_19860,N_18008,N_18767);
xnor U19861 (N_19861,N_18594,N_18268);
nand U19862 (N_19862,N_18194,N_18845);
and U19863 (N_19863,N_18771,N_18622);
nor U19864 (N_19864,N_18107,N_18298);
or U19865 (N_19865,N_18633,N_18306);
xor U19866 (N_19866,N_18634,N_18309);
and U19867 (N_19867,N_18860,N_18530);
or U19868 (N_19868,N_18951,N_18351);
xnor U19869 (N_19869,N_18141,N_18805);
nor U19870 (N_19870,N_18206,N_18685);
nand U19871 (N_19871,N_18260,N_18716);
nand U19872 (N_19872,N_18183,N_18520);
and U19873 (N_19873,N_18359,N_18979);
nand U19874 (N_19874,N_18424,N_18058);
and U19875 (N_19875,N_18973,N_18006);
nand U19876 (N_19876,N_18941,N_18285);
and U19877 (N_19877,N_18912,N_18879);
nand U19878 (N_19878,N_18222,N_18162);
or U19879 (N_19879,N_18890,N_18336);
nor U19880 (N_19880,N_18130,N_18763);
or U19881 (N_19881,N_18628,N_18910);
and U19882 (N_19882,N_18726,N_18810);
and U19883 (N_19883,N_18424,N_18934);
and U19884 (N_19884,N_18164,N_18182);
xor U19885 (N_19885,N_18643,N_18889);
and U19886 (N_19886,N_18711,N_18274);
nor U19887 (N_19887,N_18086,N_18640);
or U19888 (N_19888,N_18879,N_18384);
xor U19889 (N_19889,N_18560,N_18389);
xor U19890 (N_19890,N_18079,N_18705);
xor U19891 (N_19891,N_18309,N_18667);
and U19892 (N_19892,N_18098,N_18575);
nand U19893 (N_19893,N_18233,N_18442);
xnor U19894 (N_19894,N_18455,N_18377);
nand U19895 (N_19895,N_18017,N_18216);
xor U19896 (N_19896,N_18527,N_18420);
nor U19897 (N_19897,N_18556,N_18836);
nor U19898 (N_19898,N_18027,N_18271);
or U19899 (N_19899,N_18808,N_18265);
nand U19900 (N_19900,N_18938,N_18285);
xor U19901 (N_19901,N_18381,N_18344);
nor U19902 (N_19902,N_18014,N_18953);
xnor U19903 (N_19903,N_18826,N_18114);
xnor U19904 (N_19904,N_18888,N_18807);
and U19905 (N_19905,N_18735,N_18785);
nor U19906 (N_19906,N_18867,N_18745);
nand U19907 (N_19907,N_18175,N_18802);
or U19908 (N_19908,N_18559,N_18560);
xnor U19909 (N_19909,N_18692,N_18890);
nor U19910 (N_19910,N_18013,N_18925);
nand U19911 (N_19911,N_18250,N_18216);
or U19912 (N_19912,N_18338,N_18604);
and U19913 (N_19913,N_18982,N_18111);
nand U19914 (N_19914,N_18836,N_18431);
nand U19915 (N_19915,N_18723,N_18042);
or U19916 (N_19916,N_18927,N_18579);
xnor U19917 (N_19917,N_18408,N_18832);
nand U19918 (N_19918,N_18285,N_18881);
nor U19919 (N_19919,N_18668,N_18586);
xnor U19920 (N_19920,N_18610,N_18222);
xnor U19921 (N_19921,N_18962,N_18224);
xor U19922 (N_19922,N_18548,N_18602);
xnor U19923 (N_19923,N_18063,N_18573);
and U19924 (N_19924,N_18002,N_18542);
and U19925 (N_19925,N_18876,N_18576);
nor U19926 (N_19926,N_18849,N_18341);
xnor U19927 (N_19927,N_18413,N_18068);
and U19928 (N_19928,N_18512,N_18170);
nor U19929 (N_19929,N_18385,N_18907);
xnor U19930 (N_19930,N_18616,N_18755);
and U19931 (N_19931,N_18649,N_18404);
nor U19932 (N_19932,N_18133,N_18394);
xnor U19933 (N_19933,N_18015,N_18126);
xor U19934 (N_19934,N_18486,N_18763);
and U19935 (N_19935,N_18965,N_18517);
xnor U19936 (N_19936,N_18730,N_18791);
or U19937 (N_19937,N_18668,N_18410);
nand U19938 (N_19938,N_18785,N_18610);
nand U19939 (N_19939,N_18396,N_18822);
nand U19940 (N_19940,N_18851,N_18156);
xor U19941 (N_19941,N_18741,N_18624);
and U19942 (N_19942,N_18721,N_18881);
nand U19943 (N_19943,N_18066,N_18884);
or U19944 (N_19944,N_18477,N_18777);
xnor U19945 (N_19945,N_18809,N_18306);
xnor U19946 (N_19946,N_18500,N_18414);
or U19947 (N_19947,N_18326,N_18886);
xor U19948 (N_19948,N_18240,N_18070);
xnor U19949 (N_19949,N_18538,N_18139);
and U19950 (N_19950,N_18951,N_18279);
xor U19951 (N_19951,N_18785,N_18049);
xor U19952 (N_19952,N_18351,N_18191);
nor U19953 (N_19953,N_18563,N_18588);
and U19954 (N_19954,N_18774,N_18721);
nand U19955 (N_19955,N_18223,N_18803);
and U19956 (N_19956,N_18026,N_18760);
and U19957 (N_19957,N_18690,N_18144);
nor U19958 (N_19958,N_18729,N_18850);
xnor U19959 (N_19959,N_18068,N_18257);
nor U19960 (N_19960,N_18415,N_18305);
and U19961 (N_19961,N_18827,N_18998);
nand U19962 (N_19962,N_18335,N_18307);
or U19963 (N_19963,N_18247,N_18586);
nor U19964 (N_19964,N_18143,N_18650);
nor U19965 (N_19965,N_18193,N_18746);
or U19966 (N_19966,N_18765,N_18470);
nand U19967 (N_19967,N_18789,N_18661);
xor U19968 (N_19968,N_18543,N_18868);
nand U19969 (N_19969,N_18786,N_18740);
nor U19970 (N_19970,N_18045,N_18799);
nand U19971 (N_19971,N_18398,N_18312);
and U19972 (N_19972,N_18437,N_18403);
and U19973 (N_19973,N_18626,N_18171);
and U19974 (N_19974,N_18784,N_18017);
xnor U19975 (N_19975,N_18865,N_18595);
nand U19976 (N_19976,N_18582,N_18685);
nor U19977 (N_19977,N_18960,N_18249);
or U19978 (N_19978,N_18464,N_18693);
or U19979 (N_19979,N_18184,N_18236);
nor U19980 (N_19980,N_18418,N_18357);
nor U19981 (N_19981,N_18166,N_18021);
and U19982 (N_19982,N_18284,N_18172);
or U19983 (N_19983,N_18737,N_18837);
nor U19984 (N_19984,N_18188,N_18795);
or U19985 (N_19985,N_18676,N_18346);
and U19986 (N_19986,N_18185,N_18043);
nor U19987 (N_19987,N_18956,N_18497);
or U19988 (N_19988,N_18682,N_18062);
or U19989 (N_19989,N_18312,N_18634);
or U19990 (N_19990,N_18224,N_18535);
and U19991 (N_19991,N_18969,N_18981);
nor U19992 (N_19992,N_18761,N_18337);
nand U19993 (N_19993,N_18569,N_18686);
or U19994 (N_19994,N_18514,N_18325);
nand U19995 (N_19995,N_18359,N_18590);
nor U19996 (N_19996,N_18992,N_18495);
nor U19997 (N_19997,N_18803,N_18742);
or U19998 (N_19998,N_18904,N_18740);
nor U19999 (N_19999,N_18695,N_18583);
xor U20000 (N_20000,N_19933,N_19205);
nor U20001 (N_20001,N_19815,N_19245);
or U20002 (N_20002,N_19882,N_19171);
or U20003 (N_20003,N_19988,N_19047);
and U20004 (N_20004,N_19089,N_19691);
and U20005 (N_20005,N_19616,N_19301);
nor U20006 (N_20006,N_19352,N_19437);
or U20007 (N_20007,N_19235,N_19258);
and U20008 (N_20008,N_19878,N_19214);
or U20009 (N_20009,N_19754,N_19650);
nor U20010 (N_20010,N_19901,N_19541);
and U20011 (N_20011,N_19561,N_19978);
or U20012 (N_20012,N_19240,N_19073);
xnor U20013 (N_20013,N_19493,N_19805);
xnor U20014 (N_20014,N_19323,N_19838);
or U20015 (N_20015,N_19522,N_19197);
and U20016 (N_20016,N_19779,N_19040);
or U20017 (N_20017,N_19244,N_19989);
or U20018 (N_20018,N_19856,N_19028);
nor U20019 (N_20019,N_19926,N_19219);
xor U20020 (N_20020,N_19870,N_19496);
and U20021 (N_20021,N_19431,N_19302);
or U20022 (N_20022,N_19123,N_19160);
xnor U20023 (N_20023,N_19532,N_19286);
and U20024 (N_20024,N_19339,N_19506);
or U20025 (N_20025,N_19742,N_19417);
and U20026 (N_20026,N_19565,N_19480);
or U20027 (N_20027,N_19865,N_19049);
nor U20028 (N_20028,N_19043,N_19939);
nand U20029 (N_20029,N_19179,N_19334);
nand U20030 (N_20030,N_19918,N_19587);
or U20031 (N_20031,N_19169,N_19422);
nand U20032 (N_20032,N_19038,N_19743);
nor U20033 (N_20033,N_19002,N_19198);
xor U20034 (N_20034,N_19460,N_19615);
nor U20035 (N_20035,N_19257,N_19226);
nand U20036 (N_20036,N_19030,N_19003);
and U20037 (N_20037,N_19741,N_19381);
nor U20038 (N_20038,N_19461,N_19632);
nand U20039 (N_20039,N_19213,N_19344);
or U20040 (N_20040,N_19181,N_19410);
or U20041 (N_20041,N_19370,N_19507);
nor U20042 (N_20042,N_19780,N_19800);
and U20043 (N_20043,N_19494,N_19308);
and U20044 (N_20044,N_19877,N_19156);
and U20045 (N_20045,N_19278,N_19412);
nor U20046 (N_20046,N_19332,N_19673);
nand U20047 (N_20047,N_19702,N_19440);
or U20048 (N_20048,N_19150,N_19611);
or U20049 (N_20049,N_19623,N_19117);
nand U20050 (N_20050,N_19919,N_19145);
or U20051 (N_20051,N_19424,N_19873);
nor U20052 (N_20052,N_19377,N_19465);
xnor U20053 (N_20053,N_19822,N_19275);
nor U20054 (N_20054,N_19523,N_19902);
and U20055 (N_20055,N_19737,N_19788);
or U20056 (N_20056,N_19844,N_19980);
nand U20057 (N_20057,N_19559,N_19233);
nor U20058 (N_20058,N_19158,N_19659);
nor U20059 (N_20059,N_19828,N_19132);
xnor U20060 (N_20060,N_19393,N_19327);
and U20061 (N_20061,N_19354,N_19879);
nand U20062 (N_20062,N_19817,N_19984);
xor U20063 (N_20063,N_19639,N_19148);
nand U20064 (N_20064,N_19897,N_19135);
xor U20065 (N_20065,N_19225,N_19854);
and U20066 (N_20066,N_19391,N_19544);
nand U20067 (N_20067,N_19704,N_19651);
or U20068 (N_20068,N_19312,N_19051);
and U20069 (N_20069,N_19464,N_19316);
nand U20070 (N_20070,N_19062,N_19674);
and U20071 (N_20071,N_19239,N_19435);
or U20072 (N_20072,N_19095,N_19320);
and U20073 (N_20073,N_19201,N_19972);
or U20074 (N_20074,N_19859,N_19098);
and U20075 (N_20075,N_19328,N_19745);
nand U20076 (N_20076,N_19887,N_19299);
and U20077 (N_20077,N_19725,N_19868);
nand U20078 (N_20078,N_19773,N_19272);
or U20079 (N_20079,N_19036,N_19037);
and U20080 (N_20080,N_19599,N_19362);
nand U20081 (N_20081,N_19029,N_19941);
xor U20082 (N_20082,N_19284,N_19729);
nor U20083 (N_20083,N_19505,N_19686);
xnor U20084 (N_20084,N_19841,N_19684);
nor U20085 (N_20085,N_19768,N_19648);
and U20086 (N_20086,N_19970,N_19161);
and U20087 (N_20087,N_19900,N_19005);
and U20088 (N_20088,N_19373,N_19113);
nor U20089 (N_20089,N_19141,N_19472);
xnor U20090 (N_20090,N_19259,N_19818);
nor U20091 (N_20091,N_19336,N_19490);
nand U20092 (N_20092,N_19577,N_19318);
or U20093 (N_20093,N_19767,N_19666);
and U20094 (N_20094,N_19041,N_19994);
and U20095 (N_20095,N_19738,N_19291);
xor U20096 (N_20096,N_19597,N_19238);
and U20097 (N_20097,N_19755,N_19039);
nor U20098 (N_20098,N_19944,N_19215);
and U20099 (N_20099,N_19531,N_19916);
nor U20100 (N_20100,N_19542,N_19836);
nor U20101 (N_20101,N_19133,N_19612);
and U20102 (N_20102,N_19094,N_19649);
and U20103 (N_20103,N_19968,N_19309);
xor U20104 (N_20104,N_19142,N_19605);
or U20105 (N_20105,N_19000,N_19190);
nor U20106 (N_20106,N_19170,N_19657);
nand U20107 (N_20107,N_19384,N_19629);
nand U20108 (N_20108,N_19357,N_19671);
or U20109 (N_20109,N_19626,N_19937);
nand U20110 (N_20110,N_19798,N_19064);
and U20111 (N_20111,N_19645,N_19503);
xnor U20112 (N_20112,N_19851,N_19683);
xor U20113 (N_20113,N_19924,N_19285);
xor U20114 (N_20114,N_19837,N_19614);
or U20115 (N_20115,N_19950,N_19004);
xor U20116 (N_20116,N_19557,N_19016);
or U20117 (N_20117,N_19338,N_19891);
or U20118 (N_20118,N_19760,N_19956);
nor U20119 (N_20119,N_19409,N_19153);
xor U20120 (N_20120,N_19007,N_19564);
or U20121 (N_20121,N_19826,N_19931);
xnor U20122 (N_20122,N_19399,N_19720);
nand U20123 (N_20123,N_19356,N_19621);
and U20124 (N_20124,N_19045,N_19467);
nand U20125 (N_20125,N_19630,N_19736);
or U20126 (N_20126,N_19595,N_19162);
nand U20127 (N_20127,N_19688,N_19310);
nor U20128 (N_20128,N_19250,N_19191);
and U20129 (N_20129,N_19230,N_19146);
nor U20130 (N_20130,N_19761,N_19078);
nand U20131 (N_20131,N_19646,N_19820);
nand U20132 (N_20132,N_19242,N_19385);
xnor U20133 (N_20133,N_19023,N_19395);
xor U20134 (N_20134,N_19387,N_19508);
or U20135 (N_20135,N_19166,N_19426);
nand U20136 (N_20136,N_19392,N_19462);
nor U20137 (N_20137,N_19692,N_19194);
nor U20138 (N_20138,N_19343,N_19090);
nand U20139 (N_20139,N_19775,N_19609);
and U20140 (N_20140,N_19669,N_19488);
or U20141 (N_20141,N_19346,N_19317);
or U20142 (N_20142,N_19155,N_19174);
and U20143 (N_20143,N_19884,N_19946);
and U20144 (N_20144,N_19986,N_19330);
or U20145 (N_20145,N_19167,N_19847);
nand U20146 (N_20146,N_19396,N_19707);
xnor U20147 (N_20147,N_19789,N_19954);
nand U20148 (N_20148,N_19450,N_19102);
nor U20149 (N_20149,N_19640,N_19675);
xnor U20150 (N_20150,N_19175,N_19787);
nand U20151 (N_20151,N_19287,N_19183);
or U20152 (N_20152,N_19074,N_19189);
and U20153 (N_20153,N_19811,N_19315);
xor U20154 (N_20154,N_19898,N_19529);
nor U20155 (N_20155,N_19081,N_19716);
or U20156 (N_20156,N_19568,N_19379);
nand U20157 (N_20157,N_19177,N_19546);
or U20158 (N_20158,N_19072,N_19052);
nand U20159 (N_20159,N_19006,N_19011);
nand U20160 (N_20160,N_19375,N_19961);
or U20161 (N_20161,N_19653,N_19273);
nand U20162 (N_20162,N_19592,N_19846);
nand U20163 (N_20163,N_19187,N_19050);
or U20164 (N_20164,N_19696,N_19468);
nor U20165 (N_20165,N_19567,N_19861);
nand U20166 (N_20166,N_19790,N_19080);
or U20167 (N_20167,N_19679,N_19816);
nand U20168 (N_20168,N_19283,N_19420);
or U20169 (N_20169,N_19964,N_19063);
nand U20170 (N_20170,N_19703,N_19990);
and U20171 (N_20171,N_19104,N_19699);
nand U20172 (N_20172,N_19927,N_19015);
and U20173 (N_20173,N_19173,N_19010);
nor U20174 (N_20174,N_19517,N_19804);
nor U20175 (N_20175,N_19813,N_19252);
xnor U20176 (N_20176,N_19752,N_19721);
nand U20177 (N_20177,N_19061,N_19554);
and U20178 (N_20178,N_19509,N_19116);
and U20179 (N_20179,N_19504,N_19710);
nand U20180 (N_20180,N_19575,N_19853);
xor U20181 (N_20181,N_19724,N_19405);
nor U20182 (N_20182,N_19203,N_19447);
nand U20183 (N_20183,N_19733,N_19658);
or U20184 (N_20184,N_19572,N_19753);
and U20185 (N_20185,N_19065,N_19935);
or U20186 (N_20186,N_19976,N_19008);
xnor U20187 (N_20187,N_19758,N_19613);
xor U20188 (N_20188,N_19383,N_19122);
nor U20189 (N_20189,N_19711,N_19032);
nand U20190 (N_20190,N_19484,N_19478);
nand U20191 (N_20191,N_19670,N_19543);
nor U20192 (N_20192,N_19325,N_19152);
and U20193 (N_20193,N_19067,N_19368);
xnor U20194 (N_20194,N_19627,N_19389);
nor U20195 (N_20195,N_19911,N_19608);
or U20196 (N_20196,N_19634,N_19551);
xnor U20197 (N_20197,N_19139,N_19473);
or U20198 (N_20198,N_19289,N_19552);
nor U20199 (N_20199,N_19959,N_19101);
xnor U20200 (N_20200,N_19580,N_19021);
and U20201 (N_20201,N_19364,N_19188);
and U20202 (N_20202,N_19031,N_19553);
and U20203 (N_20203,N_19223,N_19382);
xnor U20204 (N_20204,N_19677,N_19734);
xor U20205 (N_20205,N_19034,N_19014);
and U20206 (N_20206,N_19111,N_19894);
nor U20207 (N_20207,N_19769,N_19678);
and U20208 (N_20208,N_19012,N_19855);
nand U20209 (N_20209,N_19705,N_19321);
and U20210 (N_20210,N_19211,N_19642);
xor U20211 (N_20211,N_19965,N_19566);
and U20212 (N_20212,N_19009,N_19498);
xnor U20213 (N_20213,N_19969,N_19469);
nand U20214 (N_20214,N_19172,N_19376);
xor U20215 (N_20215,N_19411,N_19921);
xnor U20216 (N_20216,N_19985,N_19936);
xnor U20217 (N_20217,N_19269,N_19774);
xnor U20218 (N_20218,N_19718,N_19366);
or U20219 (N_20219,N_19114,N_19647);
xor U20220 (N_20220,N_19660,N_19355);
or U20221 (N_20221,N_19456,N_19681);
nand U20222 (N_20222,N_19463,N_19687);
and U20223 (N_20223,N_19999,N_19351);
xor U20224 (N_20224,N_19654,N_19831);
xnor U20225 (N_20225,N_19157,N_19335);
nor U20226 (N_20226,N_19581,N_19695);
or U20227 (N_20227,N_19256,N_19513);
nand U20228 (N_20228,N_19664,N_19125);
or U20229 (N_20229,N_19727,N_19394);
xor U20230 (N_20230,N_19193,N_19501);
nand U20231 (N_20231,N_19421,N_19538);
nand U20232 (N_20232,N_19319,N_19843);
xnor U20233 (N_20233,N_19582,N_19539);
or U20234 (N_20234,N_19829,N_19076);
or U20235 (N_20235,N_19848,N_19739);
and U20236 (N_20236,N_19347,N_19255);
and U20237 (N_20237,N_19088,N_19821);
and U20238 (N_20238,N_19998,N_19908);
and U20239 (N_20239,N_19726,N_19057);
xnor U20240 (N_20240,N_19112,N_19652);
and U20241 (N_20241,N_19401,N_19680);
xnor U20242 (N_20242,N_19097,N_19303);
or U20243 (N_20243,N_19708,N_19620);
xor U20244 (N_20244,N_19860,N_19962);
nor U20245 (N_20245,N_19667,N_19583);
xnor U20246 (N_20246,N_19747,N_19129);
nor U20247 (N_20247,N_19863,N_19305);
nor U20248 (N_20248,N_19163,N_19020);
or U20249 (N_20249,N_19601,N_19408);
xor U20250 (N_20250,N_19528,N_19518);
nor U20251 (N_20251,N_19361,N_19459);
and U20252 (N_20252,N_19340,N_19665);
or U20253 (N_20253,N_19326,N_19295);
or U20254 (N_20254,N_19558,N_19949);
or U20255 (N_20255,N_19598,N_19912);
nor U20256 (N_20256,N_19812,N_19455);
or U20257 (N_20257,N_19479,N_19147);
and U20258 (N_20258,N_19083,N_19249);
xor U20259 (N_20259,N_19209,N_19143);
and U20260 (N_20260,N_19092,N_19514);
and U20261 (N_20261,N_19358,N_19140);
and U20262 (N_20262,N_19087,N_19407);
or U20263 (N_20263,N_19093,N_19271);
xor U20264 (N_20264,N_19434,N_19121);
or U20265 (N_20265,N_19866,N_19204);
nand U20266 (N_20266,N_19525,N_19261);
nor U20267 (N_20267,N_19717,N_19796);
or U20268 (N_20268,N_19397,N_19403);
nand U20269 (N_20269,N_19991,N_19292);
and U20270 (N_20270,N_19633,N_19026);
xor U20271 (N_20271,N_19224,N_19709);
and U20272 (N_20272,N_19858,N_19109);
xor U20273 (N_20273,N_19594,N_19625);
or U20274 (N_20274,N_19697,N_19110);
nand U20275 (N_20275,N_19512,N_19270);
nor U20276 (N_20276,N_19869,N_19452);
or U20277 (N_20277,N_19519,N_19850);
nand U20278 (N_20278,N_19685,N_19433);
or U20279 (N_20279,N_19719,N_19369);
and U20280 (N_20280,N_19164,N_19096);
nand U20281 (N_20281,N_19091,N_19151);
nand U20282 (N_20282,N_19212,N_19059);
nand U20283 (N_20283,N_19932,N_19547);
nand U20284 (N_20284,N_19485,N_19220);
and U20285 (N_20285,N_19159,N_19917);
or U20286 (N_20286,N_19341,N_19825);
or U20287 (N_20287,N_19953,N_19706);
xor U20288 (N_20288,N_19281,N_19910);
and U20289 (N_20289,N_19035,N_19243);
nand U20290 (N_20290,N_19521,N_19372);
nand U20291 (N_20291,N_19348,N_19909);
nor U20292 (N_20292,N_19886,N_19342);
xor U20293 (N_20293,N_19386,N_19442);
nor U20294 (N_20294,N_19839,N_19714);
xor U20295 (N_20295,N_19066,N_19550);
or U20296 (N_20296,N_19483,N_19108);
nand U20297 (N_20297,N_19195,N_19631);
nand U20298 (N_20298,N_19723,N_19746);
xor U20299 (N_20299,N_19118,N_19904);
nand U20300 (N_20300,N_19536,N_19771);
and U20301 (N_20301,N_19262,N_19444);
nor U20302 (N_20302,N_19127,N_19624);
nor U20303 (N_20303,N_19237,N_19307);
and U20304 (N_20304,N_19845,N_19981);
xor U20305 (N_20305,N_19987,N_19349);
and U20306 (N_20306,N_19929,N_19967);
xor U20307 (N_20307,N_19524,N_19712);
and U20308 (N_20308,N_19418,N_19100);
nor U20309 (N_20309,N_19236,N_19797);
and U20310 (N_20310,N_19231,N_19070);
or U20311 (N_20311,N_19644,N_19294);
nand U20312 (N_20312,N_19834,N_19446);
nor U20313 (N_20313,N_19276,N_19589);
nor U20314 (N_20314,N_19947,N_19400);
or U20315 (N_20315,N_19251,N_19574);
or U20316 (N_20316,N_19492,N_19803);
or U20317 (N_20317,N_19477,N_19265);
nor U20318 (N_20318,N_19196,N_19874);
nand U20319 (N_20319,N_19992,N_19906);
nand U20320 (N_20320,N_19951,N_19791);
xnor U20321 (N_20321,N_19562,N_19776);
or U20322 (N_20322,N_19656,N_19001);
and U20323 (N_20323,N_19533,N_19136);
or U20324 (N_20324,N_19585,N_19277);
or U20325 (N_20325,N_19690,N_19017);
xnor U20326 (N_20326,N_19495,N_19983);
nand U20327 (N_20327,N_19527,N_19331);
nor U20328 (N_20328,N_19731,N_19054);
and U20329 (N_20329,N_19573,N_19466);
and U20330 (N_20330,N_19055,N_19103);
nor U20331 (N_20331,N_19735,N_19862);
or U20332 (N_20332,N_19248,N_19306);
or U20333 (N_20333,N_19622,N_19033);
xnor U20334 (N_20334,N_19638,N_19819);
nand U20335 (N_20335,N_19290,N_19602);
and U20336 (N_20336,N_19311,N_19274);
nand U20337 (N_20337,N_19928,N_19086);
xor U20338 (N_20338,N_19732,N_19178);
xnor U20339 (N_20339,N_19963,N_19458);
and U20340 (N_20340,N_19893,N_19439);
and U20341 (N_20341,N_19329,N_19077);
nand U20342 (N_20342,N_19471,N_19606);
nor U20343 (N_20343,N_19618,N_19371);
or U20344 (N_20344,N_19835,N_19540);
or U20345 (N_20345,N_19499,N_19728);
nor U20346 (N_20346,N_19880,N_19930);
xor U20347 (N_20347,N_19892,N_19176);
and U20348 (N_20348,N_19810,N_19748);
and U20349 (N_20349,N_19068,N_19857);
nor U20350 (N_20350,N_19872,N_19635);
or U20351 (N_20351,N_19304,N_19415);
xor U20352 (N_20352,N_19751,N_19128);
xnor U20353 (N_20353,N_19764,N_19428);
or U20354 (N_20354,N_19920,N_19713);
nor U20355 (N_20355,N_19792,N_19516);
nor U20356 (N_20356,N_19526,N_19333);
and U20357 (N_20357,N_19475,N_19545);
and U20358 (N_20358,N_19266,N_19022);
or U20359 (N_20359,N_19974,N_19537);
and U20360 (N_20360,N_19107,N_19470);
and U20361 (N_20361,N_19571,N_19889);
xor U20362 (N_20362,N_19628,N_19852);
xor U20363 (N_20363,N_19324,N_19555);
and U20364 (N_20364,N_19263,N_19823);
nor U20365 (N_20365,N_19165,N_19560);
or U20366 (N_20366,N_19227,N_19130);
and U20367 (N_20367,N_19184,N_19530);
xor U20368 (N_20368,N_19216,N_19682);
and U20369 (N_20369,N_19925,N_19757);
and U20370 (N_20370,N_19693,N_19617);
or U20371 (N_20371,N_19794,N_19474);
nor U20372 (N_20372,N_19402,N_19406);
or U20373 (N_20373,N_19958,N_19661);
nand U20374 (N_20374,N_19907,N_19260);
or U20375 (N_20375,N_19228,N_19264);
nand U20376 (N_20376,N_19849,N_19481);
nand U20377 (N_20377,N_19268,N_19390);
nand U20378 (N_20378,N_19192,N_19025);
nor U20379 (N_20379,N_19378,N_19832);
xnor U20380 (N_20380,N_19247,N_19229);
or U20381 (N_20381,N_19802,N_19202);
and U20382 (N_20382,N_19979,N_19515);
or U20383 (N_20383,N_19099,N_19783);
and U20384 (N_20384,N_19942,N_19591);
nand U20385 (N_20385,N_19350,N_19782);
or U20386 (N_20386,N_19922,N_19762);
nor U20387 (N_20387,N_19085,N_19888);
nand U20388 (N_20388,N_19079,N_19876);
xnor U20389 (N_20389,N_19432,N_19363);
xnor U20390 (N_20390,N_19124,N_19182);
or U20391 (N_20391,N_19966,N_19636);
nor U20392 (N_20392,N_19715,N_19668);
xor U20393 (N_20393,N_19590,N_19772);
nor U20394 (N_20394,N_19778,N_19071);
and U20395 (N_20395,N_19842,N_19663);
nand U20396 (N_20396,N_19940,N_19476);
nor U20397 (N_20397,N_19934,N_19048);
or U20398 (N_20398,N_19084,N_19785);
or U20399 (N_20399,N_19436,N_19069);
nand U20400 (N_20400,N_19570,N_19053);
or U20401 (N_20401,N_19423,N_19082);
xor U20402 (N_20402,N_19425,N_19443);
xnor U20403 (N_20403,N_19296,N_19607);
and U20404 (N_20404,N_19763,N_19044);
or U20405 (N_20405,N_19416,N_19722);
xnor U20406 (N_20406,N_19806,N_19997);
and U20407 (N_20407,N_19042,N_19793);
xnor U20408 (N_20408,N_19267,N_19438);
nor U20409 (N_20409,N_19814,N_19883);
and U20410 (N_20410,N_19895,N_19578);
xor U20411 (N_20411,N_19106,N_19896);
nor U20412 (N_20412,N_19995,N_19337);
xor U20413 (N_20413,N_19905,N_19701);
nand U20414 (N_20414,N_19795,N_19548);
xnor U20415 (N_20415,N_19619,N_19672);
nor U20416 (N_20416,N_19777,N_19300);
and U20417 (N_20417,N_19730,N_19414);
and U20418 (N_20418,N_19218,N_19427);
or U20419 (N_20419,N_19154,N_19207);
or U20420 (N_20420,N_19801,N_19380);
nor U20421 (N_20421,N_19298,N_19134);
nor U20422 (N_20422,N_19808,N_19448);
or U20423 (N_20423,N_19871,N_19429);
nand U20424 (N_20424,N_19535,N_19960);
and U20425 (N_20425,N_19288,N_19486);
and U20426 (N_20426,N_19534,N_19971);
nor U20427 (N_20427,N_19058,N_19945);
nand U20428 (N_20428,N_19948,N_19232);
or U20429 (N_20429,N_19119,N_19497);
xnor U20430 (N_20430,N_19511,N_19584);
or U20431 (N_20431,N_19641,N_19313);
nor U20432 (N_20432,N_19867,N_19120);
xnor U20433 (N_20433,N_19643,N_19807);
or U20434 (N_20434,N_19018,N_19221);
nor U20435 (N_20435,N_19875,N_19637);
nor U20436 (N_20436,N_19914,N_19457);
xor U20437 (N_20437,N_19833,N_19293);
and U20438 (N_20438,N_19500,N_19359);
nor U20439 (N_20439,N_19445,N_19840);
or U20440 (N_20440,N_19913,N_19885);
xor U20441 (N_20441,N_19149,N_19137);
and U20442 (N_20442,N_19604,N_19596);
and U20443 (N_20443,N_19353,N_19200);
nor U20444 (N_20444,N_19280,N_19993);
and U20445 (N_20445,N_19579,N_19698);
and U20446 (N_20446,N_19689,N_19864);
or U20447 (N_20447,N_19770,N_19180);
and U20448 (N_20448,N_19046,N_19210);
nand U20449 (N_20449,N_19700,N_19482);
nand U20450 (N_20450,N_19279,N_19915);
xor U20451 (N_20451,N_19824,N_19246);
and U20452 (N_20452,N_19510,N_19019);
or U20453 (N_20453,N_19563,N_19075);
or U20454 (N_20454,N_19168,N_19588);
xnor U20455 (N_20455,N_19056,N_19199);
and U20456 (N_20456,N_19977,N_19923);
xnor U20457 (N_20457,N_19676,N_19890);
or U20458 (N_20458,N_19208,N_19185);
nor U20459 (N_20459,N_19360,N_19502);
nand U20460 (N_20460,N_19593,N_19600);
or U20461 (N_20461,N_19781,N_19144);
or U20462 (N_20462,N_19487,N_19241);
or U20463 (N_20463,N_19060,N_19784);
and U20464 (N_20464,N_19603,N_19453);
nand U20465 (N_20465,N_19955,N_19827);
nand U20466 (N_20466,N_19314,N_19206);
and U20467 (N_20467,N_19786,N_19254);
or U20468 (N_20468,N_19234,N_19186);
or U20469 (N_20469,N_19126,N_19830);
xnor U20470 (N_20470,N_19957,N_19655);
nor U20471 (N_20471,N_19549,N_19138);
xnor U20472 (N_20472,N_19374,N_19105);
xnor U20473 (N_20473,N_19610,N_19222);
nand U20474 (N_20474,N_19765,N_19973);
nor U20475 (N_20475,N_19115,N_19441);
nand U20476 (N_20476,N_19430,N_19899);
and U20477 (N_20477,N_19938,N_19024);
xor U20478 (N_20478,N_19975,N_19586);
nor U20479 (N_20479,N_19217,N_19756);
or U20480 (N_20480,N_19419,N_19451);
and U20481 (N_20481,N_19322,N_19520);
nand U20482 (N_20482,N_19398,N_19766);
and U20483 (N_20483,N_19367,N_19694);
nand U20484 (N_20484,N_19809,N_19027);
or U20485 (N_20485,N_19365,N_19952);
xnor U20486 (N_20486,N_19297,N_19345);
or U20487 (N_20487,N_19404,N_19903);
or U20488 (N_20488,N_19996,N_19799);
and U20489 (N_20489,N_19489,N_19388);
or U20490 (N_20490,N_19982,N_19491);
or U20491 (N_20491,N_19013,N_19759);
nor U20492 (N_20492,N_19740,N_19131);
xnor U20493 (N_20493,N_19576,N_19449);
nand U20494 (N_20494,N_19556,N_19569);
and U20495 (N_20495,N_19282,N_19750);
nand U20496 (N_20496,N_19943,N_19662);
and U20497 (N_20497,N_19454,N_19749);
nor U20498 (N_20498,N_19413,N_19253);
nand U20499 (N_20499,N_19881,N_19744);
xnor U20500 (N_20500,N_19193,N_19565);
nor U20501 (N_20501,N_19653,N_19246);
nand U20502 (N_20502,N_19707,N_19935);
nor U20503 (N_20503,N_19747,N_19578);
nand U20504 (N_20504,N_19719,N_19382);
and U20505 (N_20505,N_19431,N_19765);
xnor U20506 (N_20506,N_19691,N_19156);
or U20507 (N_20507,N_19040,N_19202);
and U20508 (N_20508,N_19252,N_19898);
nor U20509 (N_20509,N_19971,N_19555);
nor U20510 (N_20510,N_19591,N_19415);
or U20511 (N_20511,N_19349,N_19923);
and U20512 (N_20512,N_19558,N_19744);
and U20513 (N_20513,N_19430,N_19882);
and U20514 (N_20514,N_19619,N_19237);
nand U20515 (N_20515,N_19820,N_19322);
nor U20516 (N_20516,N_19389,N_19439);
nor U20517 (N_20517,N_19962,N_19358);
or U20518 (N_20518,N_19336,N_19329);
nor U20519 (N_20519,N_19440,N_19042);
and U20520 (N_20520,N_19308,N_19894);
nor U20521 (N_20521,N_19320,N_19774);
xnor U20522 (N_20522,N_19551,N_19823);
nand U20523 (N_20523,N_19766,N_19699);
nor U20524 (N_20524,N_19430,N_19994);
nand U20525 (N_20525,N_19863,N_19150);
or U20526 (N_20526,N_19113,N_19466);
or U20527 (N_20527,N_19139,N_19637);
or U20528 (N_20528,N_19237,N_19073);
and U20529 (N_20529,N_19800,N_19783);
and U20530 (N_20530,N_19457,N_19385);
nand U20531 (N_20531,N_19617,N_19932);
nor U20532 (N_20532,N_19372,N_19286);
or U20533 (N_20533,N_19869,N_19434);
nor U20534 (N_20534,N_19427,N_19071);
or U20535 (N_20535,N_19614,N_19121);
nor U20536 (N_20536,N_19243,N_19313);
nand U20537 (N_20537,N_19289,N_19164);
nand U20538 (N_20538,N_19995,N_19772);
nand U20539 (N_20539,N_19657,N_19505);
nor U20540 (N_20540,N_19014,N_19042);
and U20541 (N_20541,N_19902,N_19277);
or U20542 (N_20542,N_19546,N_19748);
or U20543 (N_20543,N_19798,N_19379);
and U20544 (N_20544,N_19792,N_19282);
and U20545 (N_20545,N_19054,N_19337);
nor U20546 (N_20546,N_19745,N_19937);
xor U20547 (N_20547,N_19930,N_19602);
nand U20548 (N_20548,N_19183,N_19422);
nand U20549 (N_20549,N_19985,N_19879);
nand U20550 (N_20550,N_19626,N_19976);
nand U20551 (N_20551,N_19872,N_19211);
xnor U20552 (N_20552,N_19872,N_19562);
nor U20553 (N_20553,N_19752,N_19307);
nand U20554 (N_20554,N_19179,N_19005);
nand U20555 (N_20555,N_19086,N_19655);
and U20556 (N_20556,N_19256,N_19962);
nand U20557 (N_20557,N_19341,N_19782);
nor U20558 (N_20558,N_19447,N_19192);
nor U20559 (N_20559,N_19735,N_19373);
nand U20560 (N_20560,N_19874,N_19395);
nor U20561 (N_20561,N_19114,N_19543);
xnor U20562 (N_20562,N_19562,N_19824);
and U20563 (N_20563,N_19821,N_19444);
and U20564 (N_20564,N_19533,N_19275);
xnor U20565 (N_20565,N_19615,N_19069);
or U20566 (N_20566,N_19884,N_19459);
xnor U20567 (N_20567,N_19640,N_19990);
nor U20568 (N_20568,N_19537,N_19703);
and U20569 (N_20569,N_19869,N_19458);
and U20570 (N_20570,N_19960,N_19899);
and U20571 (N_20571,N_19704,N_19201);
or U20572 (N_20572,N_19819,N_19611);
or U20573 (N_20573,N_19062,N_19150);
xnor U20574 (N_20574,N_19450,N_19108);
and U20575 (N_20575,N_19581,N_19006);
xnor U20576 (N_20576,N_19465,N_19871);
xnor U20577 (N_20577,N_19492,N_19440);
nor U20578 (N_20578,N_19267,N_19740);
and U20579 (N_20579,N_19881,N_19320);
xnor U20580 (N_20580,N_19054,N_19032);
or U20581 (N_20581,N_19367,N_19363);
and U20582 (N_20582,N_19353,N_19197);
and U20583 (N_20583,N_19092,N_19138);
nand U20584 (N_20584,N_19238,N_19545);
or U20585 (N_20585,N_19949,N_19639);
nand U20586 (N_20586,N_19109,N_19076);
and U20587 (N_20587,N_19186,N_19133);
and U20588 (N_20588,N_19550,N_19241);
xor U20589 (N_20589,N_19624,N_19028);
or U20590 (N_20590,N_19484,N_19329);
nand U20591 (N_20591,N_19361,N_19096);
or U20592 (N_20592,N_19354,N_19973);
nand U20593 (N_20593,N_19639,N_19665);
nor U20594 (N_20594,N_19541,N_19331);
and U20595 (N_20595,N_19212,N_19063);
nand U20596 (N_20596,N_19996,N_19518);
nand U20597 (N_20597,N_19066,N_19073);
or U20598 (N_20598,N_19185,N_19284);
xor U20599 (N_20599,N_19736,N_19150);
xor U20600 (N_20600,N_19930,N_19687);
nand U20601 (N_20601,N_19074,N_19066);
nor U20602 (N_20602,N_19119,N_19227);
and U20603 (N_20603,N_19561,N_19132);
and U20604 (N_20604,N_19160,N_19425);
or U20605 (N_20605,N_19831,N_19768);
nor U20606 (N_20606,N_19913,N_19533);
and U20607 (N_20607,N_19606,N_19438);
xnor U20608 (N_20608,N_19405,N_19256);
or U20609 (N_20609,N_19551,N_19755);
and U20610 (N_20610,N_19350,N_19612);
and U20611 (N_20611,N_19240,N_19545);
nor U20612 (N_20612,N_19100,N_19404);
nand U20613 (N_20613,N_19601,N_19841);
nor U20614 (N_20614,N_19848,N_19966);
or U20615 (N_20615,N_19549,N_19776);
and U20616 (N_20616,N_19457,N_19066);
or U20617 (N_20617,N_19293,N_19420);
or U20618 (N_20618,N_19808,N_19512);
nor U20619 (N_20619,N_19209,N_19682);
and U20620 (N_20620,N_19391,N_19733);
or U20621 (N_20621,N_19692,N_19949);
nand U20622 (N_20622,N_19979,N_19387);
or U20623 (N_20623,N_19250,N_19555);
and U20624 (N_20624,N_19951,N_19237);
xnor U20625 (N_20625,N_19437,N_19451);
or U20626 (N_20626,N_19393,N_19360);
or U20627 (N_20627,N_19752,N_19345);
and U20628 (N_20628,N_19794,N_19599);
nor U20629 (N_20629,N_19913,N_19691);
nand U20630 (N_20630,N_19393,N_19339);
and U20631 (N_20631,N_19186,N_19677);
nand U20632 (N_20632,N_19093,N_19471);
nand U20633 (N_20633,N_19094,N_19745);
and U20634 (N_20634,N_19986,N_19068);
nand U20635 (N_20635,N_19066,N_19520);
xnor U20636 (N_20636,N_19074,N_19183);
or U20637 (N_20637,N_19790,N_19049);
and U20638 (N_20638,N_19751,N_19382);
nor U20639 (N_20639,N_19695,N_19892);
or U20640 (N_20640,N_19816,N_19132);
nand U20641 (N_20641,N_19351,N_19125);
nor U20642 (N_20642,N_19248,N_19779);
xnor U20643 (N_20643,N_19950,N_19095);
xor U20644 (N_20644,N_19168,N_19226);
or U20645 (N_20645,N_19886,N_19060);
or U20646 (N_20646,N_19357,N_19461);
and U20647 (N_20647,N_19953,N_19194);
nand U20648 (N_20648,N_19234,N_19836);
xor U20649 (N_20649,N_19947,N_19639);
xnor U20650 (N_20650,N_19835,N_19437);
xnor U20651 (N_20651,N_19133,N_19269);
and U20652 (N_20652,N_19465,N_19515);
nand U20653 (N_20653,N_19953,N_19261);
xnor U20654 (N_20654,N_19765,N_19165);
nor U20655 (N_20655,N_19243,N_19354);
xor U20656 (N_20656,N_19462,N_19864);
xnor U20657 (N_20657,N_19565,N_19530);
xnor U20658 (N_20658,N_19699,N_19989);
nor U20659 (N_20659,N_19698,N_19852);
nor U20660 (N_20660,N_19050,N_19782);
or U20661 (N_20661,N_19053,N_19561);
xor U20662 (N_20662,N_19680,N_19940);
xor U20663 (N_20663,N_19836,N_19703);
nand U20664 (N_20664,N_19500,N_19944);
xnor U20665 (N_20665,N_19903,N_19188);
or U20666 (N_20666,N_19897,N_19240);
nand U20667 (N_20667,N_19913,N_19659);
or U20668 (N_20668,N_19674,N_19388);
or U20669 (N_20669,N_19399,N_19055);
nor U20670 (N_20670,N_19274,N_19710);
nor U20671 (N_20671,N_19193,N_19075);
xnor U20672 (N_20672,N_19774,N_19676);
xnor U20673 (N_20673,N_19277,N_19698);
nand U20674 (N_20674,N_19993,N_19301);
nor U20675 (N_20675,N_19629,N_19364);
xnor U20676 (N_20676,N_19668,N_19130);
nand U20677 (N_20677,N_19382,N_19546);
or U20678 (N_20678,N_19487,N_19814);
and U20679 (N_20679,N_19371,N_19969);
nand U20680 (N_20680,N_19239,N_19595);
nand U20681 (N_20681,N_19473,N_19733);
nand U20682 (N_20682,N_19886,N_19438);
or U20683 (N_20683,N_19925,N_19471);
xor U20684 (N_20684,N_19139,N_19746);
or U20685 (N_20685,N_19463,N_19421);
xor U20686 (N_20686,N_19673,N_19511);
and U20687 (N_20687,N_19792,N_19984);
xor U20688 (N_20688,N_19730,N_19288);
nor U20689 (N_20689,N_19700,N_19087);
nand U20690 (N_20690,N_19256,N_19541);
or U20691 (N_20691,N_19626,N_19416);
and U20692 (N_20692,N_19192,N_19475);
xnor U20693 (N_20693,N_19000,N_19563);
nand U20694 (N_20694,N_19587,N_19506);
nand U20695 (N_20695,N_19645,N_19537);
xnor U20696 (N_20696,N_19281,N_19863);
xnor U20697 (N_20697,N_19475,N_19250);
or U20698 (N_20698,N_19952,N_19050);
nor U20699 (N_20699,N_19438,N_19343);
or U20700 (N_20700,N_19876,N_19223);
xor U20701 (N_20701,N_19641,N_19768);
xor U20702 (N_20702,N_19114,N_19346);
and U20703 (N_20703,N_19205,N_19190);
or U20704 (N_20704,N_19598,N_19039);
nor U20705 (N_20705,N_19797,N_19759);
or U20706 (N_20706,N_19517,N_19441);
nor U20707 (N_20707,N_19717,N_19228);
xnor U20708 (N_20708,N_19585,N_19017);
xor U20709 (N_20709,N_19142,N_19464);
xnor U20710 (N_20710,N_19523,N_19544);
xor U20711 (N_20711,N_19223,N_19169);
and U20712 (N_20712,N_19575,N_19385);
and U20713 (N_20713,N_19661,N_19796);
nor U20714 (N_20714,N_19429,N_19094);
nand U20715 (N_20715,N_19066,N_19294);
xnor U20716 (N_20716,N_19081,N_19065);
xnor U20717 (N_20717,N_19709,N_19689);
nor U20718 (N_20718,N_19914,N_19594);
and U20719 (N_20719,N_19107,N_19380);
and U20720 (N_20720,N_19214,N_19519);
and U20721 (N_20721,N_19994,N_19867);
or U20722 (N_20722,N_19031,N_19262);
or U20723 (N_20723,N_19001,N_19745);
nand U20724 (N_20724,N_19456,N_19733);
nand U20725 (N_20725,N_19919,N_19431);
and U20726 (N_20726,N_19649,N_19677);
or U20727 (N_20727,N_19992,N_19688);
and U20728 (N_20728,N_19926,N_19937);
or U20729 (N_20729,N_19107,N_19659);
or U20730 (N_20730,N_19446,N_19180);
and U20731 (N_20731,N_19206,N_19706);
and U20732 (N_20732,N_19181,N_19124);
or U20733 (N_20733,N_19368,N_19333);
nand U20734 (N_20734,N_19530,N_19956);
nand U20735 (N_20735,N_19290,N_19150);
nor U20736 (N_20736,N_19732,N_19697);
nor U20737 (N_20737,N_19187,N_19309);
and U20738 (N_20738,N_19836,N_19374);
nand U20739 (N_20739,N_19935,N_19418);
and U20740 (N_20740,N_19691,N_19272);
xor U20741 (N_20741,N_19913,N_19840);
and U20742 (N_20742,N_19572,N_19024);
or U20743 (N_20743,N_19569,N_19231);
and U20744 (N_20744,N_19687,N_19325);
nor U20745 (N_20745,N_19070,N_19357);
xnor U20746 (N_20746,N_19278,N_19741);
and U20747 (N_20747,N_19427,N_19944);
and U20748 (N_20748,N_19061,N_19618);
or U20749 (N_20749,N_19157,N_19696);
and U20750 (N_20750,N_19860,N_19380);
xor U20751 (N_20751,N_19288,N_19692);
nor U20752 (N_20752,N_19991,N_19808);
or U20753 (N_20753,N_19863,N_19624);
or U20754 (N_20754,N_19757,N_19317);
nand U20755 (N_20755,N_19138,N_19556);
and U20756 (N_20756,N_19761,N_19506);
or U20757 (N_20757,N_19537,N_19434);
or U20758 (N_20758,N_19396,N_19321);
and U20759 (N_20759,N_19217,N_19827);
and U20760 (N_20760,N_19487,N_19110);
nand U20761 (N_20761,N_19002,N_19875);
nor U20762 (N_20762,N_19905,N_19539);
and U20763 (N_20763,N_19983,N_19015);
and U20764 (N_20764,N_19108,N_19646);
or U20765 (N_20765,N_19292,N_19993);
or U20766 (N_20766,N_19821,N_19918);
or U20767 (N_20767,N_19056,N_19423);
xor U20768 (N_20768,N_19959,N_19574);
and U20769 (N_20769,N_19632,N_19614);
nor U20770 (N_20770,N_19165,N_19798);
nand U20771 (N_20771,N_19615,N_19973);
nand U20772 (N_20772,N_19693,N_19663);
nand U20773 (N_20773,N_19474,N_19774);
nand U20774 (N_20774,N_19936,N_19952);
and U20775 (N_20775,N_19444,N_19328);
nor U20776 (N_20776,N_19944,N_19898);
and U20777 (N_20777,N_19873,N_19206);
or U20778 (N_20778,N_19184,N_19241);
nor U20779 (N_20779,N_19205,N_19181);
xnor U20780 (N_20780,N_19997,N_19262);
nor U20781 (N_20781,N_19568,N_19833);
nor U20782 (N_20782,N_19454,N_19849);
xnor U20783 (N_20783,N_19133,N_19965);
nor U20784 (N_20784,N_19861,N_19381);
and U20785 (N_20785,N_19751,N_19801);
and U20786 (N_20786,N_19876,N_19624);
or U20787 (N_20787,N_19920,N_19130);
nor U20788 (N_20788,N_19156,N_19312);
or U20789 (N_20789,N_19480,N_19698);
xnor U20790 (N_20790,N_19430,N_19893);
nor U20791 (N_20791,N_19367,N_19979);
xnor U20792 (N_20792,N_19792,N_19945);
nand U20793 (N_20793,N_19971,N_19609);
or U20794 (N_20794,N_19062,N_19995);
nor U20795 (N_20795,N_19433,N_19398);
nor U20796 (N_20796,N_19588,N_19067);
nor U20797 (N_20797,N_19179,N_19302);
and U20798 (N_20798,N_19618,N_19079);
nor U20799 (N_20799,N_19891,N_19897);
or U20800 (N_20800,N_19937,N_19776);
and U20801 (N_20801,N_19356,N_19429);
nor U20802 (N_20802,N_19758,N_19457);
or U20803 (N_20803,N_19422,N_19529);
or U20804 (N_20804,N_19408,N_19053);
nor U20805 (N_20805,N_19515,N_19145);
and U20806 (N_20806,N_19116,N_19204);
xnor U20807 (N_20807,N_19451,N_19607);
nand U20808 (N_20808,N_19324,N_19055);
xnor U20809 (N_20809,N_19003,N_19957);
xnor U20810 (N_20810,N_19052,N_19571);
and U20811 (N_20811,N_19878,N_19621);
or U20812 (N_20812,N_19824,N_19827);
or U20813 (N_20813,N_19857,N_19901);
nand U20814 (N_20814,N_19547,N_19580);
nand U20815 (N_20815,N_19572,N_19412);
nand U20816 (N_20816,N_19767,N_19001);
nor U20817 (N_20817,N_19155,N_19936);
nor U20818 (N_20818,N_19776,N_19657);
and U20819 (N_20819,N_19654,N_19363);
nand U20820 (N_20820,N_19799,N_19644);
nand U20821 (N_20821,N_19972,N_19493);
or U20822 (N_20822,N_19568,N_19344);
and U20823 (N_20823,N_19816,N_19222);
and U20824 (N_20824,N_19013,N_19773);
nor U20825 (N_20825,N_19802,N_19475);
nand U20826 (N_20826,N_19557,N_19463);
nor U20827 (N_20827,N_19334,N_19636);
nor U20828 (N_20828,N_19678,N_19528);
nand U20829 (N_20829,N_19483,N_19515);
and U20830 (N_20830,N_19588,N_19957);
nand U20831 (N_20831,N_19859,N_19791);
nand U20832 (N_20832,N_19045,N_19937);
nand U20833 (N_20833,N_19574,N_19072);
and U20834 (N_20834,N_19505,N_19976);
nand U20835 (N_20835,N_19479,N_19177);
or U20836 (N_20836,N_19489,N_19995);
or U20837 (N_20837,N_19452,N_19474);
xnor U20838 (N_20838,N_19621,N_19796);
xor U20839 (N_20839,N_19910,N_19593);
and U20840 (N_20840,N_19908,N_19252);
or U20841 (N_20841,N_19103,N_19025);
nand U20842 (N_20842,N_19922,N_19410);
or U20843 (N_20843,N_19939,N_19436);
nand U20844 (N_20844,N_19821,N_19491);
and U20845 (N_20845,N_19344,N_19177);
nor U20846 (N_20846,N_19170,N_19640);
nand U20847 (N_20847,N_19100,N_19771);
and U20848 (N_20848,N_19260,N_19150);
or U20849 (N_20849,N_19093,N_19729);
and U20850 (N_20850,N_19969,N_19273);
nand U20851 (N_20851,N_19918,N_19483);
and U20852 (N_20852,N_19538,N_19607);
nor U20853 (N_20853,N_19782,N_19279);
xnor U20854 (N_20854,N_19493,N_19198);
and U20855 (N_20855,N_19168,N_19420);
and U20856 (N_20856,N_19305,N_19716);
xnor U20857 (N_20857,N_19104,N_19034);
nand U20858 (N_20858,N_19498,N_19932);
xnor U20859 (N_20859,N_19894,N_19732);
nor U20860 (N_20860,N_19827,N_19362);
xnor U20861 (N_20861,N_19091,N_19491);
and U20862 (N_20862,N_19195,N_19490);
nand U20863 (N_20863,N_19285,N_19125);
nand U20864 (N_20864,N_19335,N_19851);
or U20865 (N_20865,N_19648,N_19671);
and U20866 (N_20866,N_19336,N_19433);
nand U20867 (N_20867,N_19088,N_19677);
or U20868 (N_20868,N_19852,N_19462);
or U20869 (N_20869,N_19747,N_19089);
nand U20870 (N_20870,N_19714,N_19366);
or U20871 (N_20871,N_19208,N_19702);
nand U20872 (N_20872,N_19785,N_19476);
and U20873 (N_20873,N_19010,N_19333);
nor U20874 (N_20874,N_19879,N_19260);
and U20875 (N_20875,N_19951,N_19185);
nand U20876 (N_20876,N_19331,N_19688);
nand U20877 (N_20877,N_19921,N_19432);
nand U20878 (N_20878,N_19624,N_19766);
xnor U20879 (N_20879,N_19885,N_19199);
and U20880 (N_20880,N_19446,N_19393);
or U20881 (N_20881,N_19384,N_19860);
xnor U20882 (N_20882,N_19806,N_19744);
or U20883 (N_20883,N_19154,N_19293);
or U20884 (N_20884,N_19400,N_19811);
xor U20885 (N_20885,N_19768,N_19776);
and U20886 (N_20886,N_19147,N_19161);
and U20887 (N_20887,N_19763,N_19905);
nand U20888 (N_20888,N_19804,N_19064);
nor U20889 (N_20889,N_19707,N_19056);
xor U20890 (N_20890,N_19052,N_19681);
nor U20891 (N_20891,N_19524,N_19978);
nand U20892 (N_20892,N_19330,N_19422);
nand U20893 (N_20893,N_19041,N_19990);
xnor U20894 (N_20894,N_19012,N_19471);
nand U20895 (N_20895,N_19462,N_19024);
xnor U20896 (N_20896,N_19566,N_19765);
or U20897 (N_20897,N_19763,N_19870);
or U20898 (N_20898,N_19964,N_19573);
nor U20899 (N_20899,N_19989,N_19991);
nand U20900 (N_20900,N_19670,N_19452);
nand U20901 (N_20901,N_19120,N_19884);
or U20902 (N_20902,N_19608,N_19361);
or U20903 (N_20903,N_19304,N_19255);
or U20904 (N_20904,N_19974,N_19346);
or U20905 (N_20905,N_19156,N_19666);
or U20906 (N_20906,N_19082,N_19245);
and U20907 (N_20907,N_19304,N_19430);
nor U20908 (N_20908,N_19748,N_19754);
or U20909 (N_20909,N_19785,N_19935);
nor U20910 (N_20910,N_19696,N_19999);
and U20911 (N_20911,N_19406,N_19181);
xor U20912 (N_20912,N_19602,N_19403);
or U20913 (N_20913,N_19603,N_19913);
and U20914 (N_20914,N_19632,N_19756);
nand U20915 (N_20915,N_19150,N_19245);
nor U20916 (N_20916,N_19963,N_19374);
nand U20917 (N_20917,N_19038,N_19402);
nor U20918 (N_20918,N_19112,N_19382);
and U20919 (N_20919,N_19305,N_19475);
or U20920 (N_20920,N_19291,N_19094);
nor U20921 (N_20921,N_19939,N_19847);
nand U20922 (N_20922,N_19723,N_19286);
xnor U20923 (N_20923,N_19779,N_19333);
xnor U20924 (N_20924,N_19276,N_19254);
nand U20925 (N_20925,N_19777,N_19013);
xnor U20926 (N_20926,N_19568,N_19445);
or U20927 (N_20927,N_19054,N_19387);
nor U20928 (N_20928,N_19098,N_19587);
xor U20929 (N_20929,N_19715,N_19580);
nor U20930 (N_20930,N_19664,N_19657);
and U20931 (N_20931,N_19035,N_19600);
nor U20932 (N_20932,N_19594,N_19329);
and U20933 (N_20933,N_19952,N_19853);
xnor U20934 (N_20934,N_19081,N_19924);
nor U20935 (N_20935,N_19518,N_19117);
or U20936 (N_20936,N_19658,N_19054);
nand U20937 (N_20937,N_19419,N_19654);
nor U20938 (N_20938,N_19092,N_19455);
xor U20939 (N_20939,N_19270,N_19861);
nand U20940 (N_20940,N_19750,N_19273);
xnor U20941 (N_20941,N_19399,N_19680);
nor U20942 (N_20942,N_19968,N_19287);
nand U20943 (N_20943,N_19032,N_19566);
xor U20944 (N_20944,N_19712,N_19026);
nand U20945 (N_20945,N_19389,N_19748);
xnor U20946 (N_20946,N_19874,N_19175);
nand U20947 (N_20947,N_19416,N_19699);
nor U20948 (N_20948,N_19690,N_19145);
xor U20949 (N_20949,N_19495,N_19619);
and U20950 (N_20950,N_19389,N_19947);
or U20951 (N_20951,N_19082,N_19662);
or U20952 (N_20952,N_19916,N_19702);
xor U20953 (N_20953,N_19386,N_19548);
and U20954 (N_20954,N_19740,N_19985);
and U20955 (N_20955,N_19185,N_19402);
nand U20956 (N_20956,N_19226,N_19600);
nor U20957 (N_20957,N_19759,N_19457);
and U20958 (N_20958,N_19795,N_19773);
and U20959 (N_20959,N_19068,N_19341);
xor U20960 (N_20960,N_19863,N_19596);
or U20961 (N_20961,N_19804,N_19079);
and U20962 (N_20962,N_19012,N_19680);
xor U20963 (N_20963,N_19267,N_19891);
nor U20964 (N_20964,N_19239,N_19335);
or U20965 (N_20965,N_19786,N_19140);
or U20966 (N_20966,N_19044,N_19955);
xnor U20967 (N_20967,N_19801,N_19046);
nand U20968 (N_20968,N_19296,N_19501);
xnor U20969 (N_20969,N_19645,N_19817);
and U20970 (N_20970,N_19897,N_19968);
and U20971 (N_20971,N_19289,N_19480);
or U20972 (N_20972,N_19989,N_19652);
or U20973 (N_20973,N_19063,N_19426);
nor U20974 (N_20974,N_19552,N_19708);
and U20975 (N_20975,N_19514,N_19347);
nor U20976 (N_20976,N_19898,N_19808);
nor U20977 (N_20977,N_19460,N_19617);
nor U20978 (N_20978,N_19021,N_19494);
xnor U20979 (N_20979,N_19293,N_19958);
and U20980 (N_20980,N_19305,N_19189);
and U20981 (N_20981,N_19183,N_19106);
nor U20982 (N_20982,N_19214,N_19477);
nand U20983 (N_20983,N_19590,N_19255);
xor U20984 (N_20984,N_19452,N_19013);
nand U20985 (N_20985,N_19384,N_19974);
or U20986 (N_20986,N_19648,N_19219);
xnor U20987 (N_20987,N_19603,N_19985);
xor U20988 (N_20988,N_19754,N_19371);
and U20989 (N_20989,N_19965,N_19975);
and U20990 (N_20990,N_19143,N_19607);
nand U20991 (N_20991,N_19242,N_19005);
and U20992 (N_20992,N_19398,N_19175);
xor U20993 (N_20993,N_19759,N_19407);
xnor U20994 (N_20994,N_19903,N_19196);
and U20995 (N_20995,N_19260,N_19428);
xor U20996 (N_20996,N_19066,N_19350);
and U20997 (N_20997,N_19326,N_19330);
or U20998 (N_20998,N_19399,N_19936);
nor U20999 (N_20999,N_19407,N_19431);
and U21000 (N_21000,N_20524,N_20844);
or U21001 (N_21001,N_20744,N_20275);
xor U21002 (N_21002,N_20779,N_20915);
nor U21003 (N_21003,N_20563,N_20062);
xnor U21004 (N_21004,N_20700,N_20196);
nand U21005 (N_21005,N_20813,N_20268);
nor U21006 (N_21006,N_20038,N_20909);
and U21007 (N_21007,N_20978,N_20167);
xor U21008 (N_21008,N_20967,N_20458);
xnor U21009 (N_21009,N_20519,N_20316);
and U21010 (N_21010,N_20745,N_20867);
xor U21011 (N_21011,N_20684,N_20827);
xnor U21012 (N_21012,N_20231,N_20694);
nor U21013 (N_21013,N_20259,N_20993);
nor U21014 (N_21014,N_20082,N_20509);
nor U21015 (N_21015,N_20195,N_20849);
xnor U21016 (N_21016,N_20617,N_20816);
or U21017 (N_21017,N_20024,N_20814);
and U21018 (N_21018,N_20720,N_20863);
nor U21019 (N_21019,N_20707,N_20203);
or U21020 (N_21020,N_20468,N_20857);
and U21021 (N_21021,N_20184,N_20030);
and U21022 (N_21022,N_20363,N_20091);
and U21023 (N_21023,N_20862,N_20318);
nor U21024 (N_21024,N_20800,N_20242);
and U21025 (N_21025,N_20096,N_20898);
nand U21026 (N_21026,N_20561,N_20313);
or U21027 (N_21027,N_20523,N_20326);
nand U21028 (N_21028,N_20350,N_20801);
and U21029 (N_21029,N_20003,N_20330);
nor U21030 (N_21030,N_20197,N_20864);
or U21031 (N_21031,N_20160,N_20175);
or U21032 (N_21032,N_20402,N_20940);
and U21033 (N_21033,N_20878,N_20409);
and U21034 (N_21034,N_20151,N_20532);
nand U21035 (N_21035,N_20772,N_20150);
xnor U21036 (N_21036,N_20164,N_20792);
xnor U21037 (N_21037,N_20022,N_20450);
or U21038 (N_21038,N_20361,N_20202);
xnor U21039 (N_21039,N_20434,N_20504);
nand U21040 (N_21040,N_20911,N_20227);
or U21041 (N_21041,N_20838,N_20455);
nor U21042 (N_21042,N_20728,N_20642);
nand U21043 (N_21043,N_20241,N_20820);
nand U21044 (N_21044,N_20056,N_20299);
nand U21045 (N_21045,N_20896,N_20696);
xor U21046 (N_21046,N_20127,N_20329);
nor U21047 (N_21047,N_20077,N_20636);
xor U21048 (N_21048,N_20635,N_20602);
nor U21049 (N_21049,N_20295,N_20992);
and U21050 (N_21050,N_20346,N_20185);
or U21051 (N_21051,N_20803,N_20607);
xor U21052 (N_21052,N_20163,N_20530);
or U21053 (N_21053,N_20328,N_20702);
nand U21054 (N_21054,N_20173,N_20836);
or U21055 (N_21055,N_20616,N_20638);
nand U21056 (N_21056,N_20076,N_20614);
nor U21057 (N_21057,N_20209,N_20172);
or U21058 (N_21058,N_20390,N_20970);
nor U21059 (N_21059,N_20860,N_20947);
nand U21060 (N_21060,N_20748,N_20976);
and U21061 (N_21061,N_20325,N_20569);
or U21062 (N_21062,N_20348,N_20232);
nand U21063 (N_21063,N_20550,N_20264);
or U21064 (N_21064,N_20655,N_20539);
and U21065 (N_21065,N_20144,N_20681);
xnor U21066 (N_21066,N_20333,N_20510);
nor U21067 (N_21067,N_20287,N_20025);
or U21068 (N_21068,N_20634,N_20305);
nand U21069 (N_21069,N_20930,N_20987);
xnor U21070 (N_21070,N_20985,N_20027);
or U21071 (N_21071,N_20042,N_20907);
nor U21072 (N_21072,N_20078,N_20537);
and U21073 (N_21073,N_20087,N_20861);
xor U21074 (N_21074,N_20248,N_20183);
and U21075 (N_21075,N_20875,N_20274);
xor U21076 (N_21076,N_20579,N_20641);
nor U21077 (N_21077,N_20417,N_20522);
nand U21078 (N_21078,N_20729,N_20063);
nor U21079 (N_21079,N_20604,N_20050);
nand U21080 (N_21080,N_20893,N_20156);
or U21081 (N_21081,N_20223,N_20923);
or U21082 (N_21082,N_20805,N_20775);
nor U21083 (N_21083,N_20971,N_20252);
nor U21084 (N_21084,N_20126,N_20407);
nor U21085 (N_21085,N_20317,N_20491);
xor U21086 (N_21086,N_20406,N_20640);
and U21087 (N_21087,N_20719,N_20016);
nor U21088 (N_21088,N_20324,N_20136);
nor U21089 (N_21089,N_20486,N_20538);
nor U21090 (N_21090,N_20286,N_20675);
or U21091 (N_21091,N_20633,N_20422);
nand U21092 (N_21092,N_20131,N_20632);
xnor U21093 (N_21093,N_20307,N_20322);
nor U21094 (N_21094,N_20986,N_20804);
xor U21095 (N_21095,N_20843,N_20228);
xor U21096 (N_21096,N_20605,N_20595);
nor U21097 (N_21097,N_20858,N_20431);
and U21098 (N_21098,N_20370,N_20656);
nor U21099 (N_21099,N_20041,N_20683);
xnor U21100 (N_21100,N_20193,N_20213);
nand U21101 (N_21101,N_20693,N_20599);
or U21102 (N_21102,N_20574,N_20997);
nor U21103 (N_21103,N_20780,N_20446);
nand U21104 (N_21104,N_20709,N_20397);
and U21105 (N_21105,N_20437,N_20393);
or U21106 (N_21106,N_20277,N_20447);
xnor U21107 (N_21107,N_20420,N_20722);
nand U21108 (N_21108,N_20122,N_20756);
nor U21109 (N_21109,N_20036,N_20888);
and U21110 (N_21110,N_20984,N_20680);
nor U21111 (N_21111,N_20462,N_20754);
and U21112 (N_21112,N_20066,N_20960);
and U21113 (N_21113,N_20289,N_20250);
xnor U21114 (N_21114,N_20181,N_20104);
nand U21115 (N_21115,N_20883,N_20587);
and U21116 (N_21116,N_20483,N_20865);
and U21117 (N_21117,N_20375,N_20549);
nand U21118 (N_21118,N_20668,N_20618);
nor U21119 (N_21119,N_20005,N_20601);
and U21120 (N_21120,N_20663,N_20021);
nor U21121 (N_21121,N_20753,N_20777);
nor U21122 (N_21122,N_20321,N_20059);
or U21123 (N_21123,N_20552,N_20244);
nand U21124 (N_21124,N_20531,N_20314);
or U21125 (N_21125,N_20536,N_20302);
nand U21126 (N_21126,N_20651,N_20047);
or U21127 (N_21127,N_20678,N_20502);
and U21128 (N_21128,N_20917,N_20500);
xnor U21129 (N_21129,N_20735,N_20107);
nor U21130 (N_21130,N_20399,N_20750);
and U21131 (N_21131,N_20235,N_20829);
or U21132 (N_21132,N_20981,N_20269);
or U21133 (N_21133,N_20479,N_20237);
or U21134 (N_21134,N_20043,N_20726);
or U21135 (N_21135,N_20225,N_20263);
xor U21136 (N_21136,N_20906,N_20764);
and U21137 (N_21137,N_20095,N_20508);
xor U21138 (N_21138,N_20391,N_20189);
xnor U21139 (N_21139,N_20426,N_20889);
xor U21140 (N_21140,N_20413,N_20588);
nor U21141 (N_21141,N_20033,N_20824);
nand U21142 (N_21142,N_20414,N_20841);
or U21143 (N_21143,N_20100,N_20471);
nand U21144 (N_21144,N_20188,N_20020);
nand U21145 (N_21145,N_20855,N_20380);
and U21146 (N_21146,N_20137,N_20541);
xor U21147 (N_21147,N_20443,N_20123);
xor U21148 (N_21148,N_20125,N_20254);
and U21149 (N_21149,N_20247,N_20396);
nand U21150 (N_21150,N_20647,N_20400);
or U21151 (N_21151,N_20395,N_20384);
or U21152 (N_21152,N_20288,N_20236);
nor U21153 (N_21153,N_20449,N_20210);
nand U21154 (N_21154,N_20945,N_20989);
and U21155 (N_21155,N_20742,N_20854);
or U21156 (N_21156,N_20685,N_20498);
nand U21157 (N_21157,N_20902,N_20276);
nor U21158 (N_21158,N_20723,N_20146);
or U21159 (N_21159,N_20578,N_20162);
nor U21160 (N_21160,N_20028,N_20597);
or U21161 (N_21161,N_20545,N_20895);
or U21162 (N_21162,N_20686,N_20124);
nor U21163 (N_21163,N_20881,N_20874);
nor U21164 (N_21164,N_20461,N_20948);
or U21165 (N_21165,N_20535,N_20529);
xor U21166 (N_21166,N_20734,N_20799);
or U21167 (N_21167,N_20416,N_20782);
nand U21168 (N_21168,N_20703,N_20645);
xnor U21169 (N_21169,N_20925,N_20736);
and U21170 (N_21170,N_20637,N_20831);
xnor U21171 (N_21171,N_20489,N_20919);
and U21172 (N_21172,N_20044,N_20267);
xnor U21173 (N_21173,N_20731,N_20963);
and U21174 (N_21174,N_20432,N_20639);
xnor U21175 (N_21175,N_20961,N_20011);
nor U21176 (N_21176,N_20293,N_20904);
or U21177 (N_21177,N_20732,N_20755);
nand U21178 (N_21178,N_20004,N_20323);
and U21179 (N_21179,N_20015,N_20628);
nand U21180 (N_21180,N_20029,N_20715);
nand U21181 (N_21181,N_20965,N_20320);
xor U21182 (N_21182,N_20939,N_20619);
nand U21183 (N_21183,N_20751,N_20879);
nor U21184 (N_21184,N_20679,N_20953);
xor U21185 (N_21185,N_20944,N_20442);
and U21186 (N_21186,N_20376,N_20856);
xnor U21187 (N_21187,N_20784,N_20743);
and U21188 (N_21188,N_20566,N_20718);
and U21189 (N_21189,N_20064,N_20142);
nor U21190 (N_21190,N_20075,N_20596);
nand U21191 (N_21191,N_20952,N_20518);
or U21192 (N_21192,N_20847,N_20996);
nor U21193 (N_21193,N_20187,N_20284);
nand U21194 (N_21194,N_20215,N_20897);
or U21195 (N_21195,N_20892,N_20469);
and U21196 (N_21196,N_20759,N_20337);
nor U21197 (N_21197,N_20752,N_20212);
nor U21198 (N_21198,N_20155,N_20999);
xor U21199 (N_21199,N_20418,N_20783);
or U21200 (N_21200,N_20311,N_20593);
or U21201 (N_21201,N_20079,N_20112);
nor U21202 (N_21202,N_20866,N_20891);
xnor U21203 (N_21203,N_20620,N_20916);
and U21204 (N_21204,N_20084,N_20834);
xnor U21205 (N_21205,N_20154,N_20933);
xor U21206 (N_21206,N_20503,N_20762);
and U21207 (N_21207,N_20010,N_20186);
nor U21208 (N_21208,N_20401,N_20922);
or U21209 (N_21209,N_20977,N_20873);
xnor U21210 (N_21210,N_20631,N_20201);
nand U21211 (N_21211,N_20367,N_20962);
nand U21212 (N_21212,N_20886,N_20382);
xnor U21213 (N_21213,N_20558,N_20546);
and U21214 (N_21214,N_20830,N_20665);
xor U21215 (N_21215,N_20791,N_20257);
or U21216 (N_21216,N_20515,N_20262);
xor U21217 (N_21217,N_20551,N_20332);
xor U21218 (N_21218,N_20472,N_20219);
or U21219 (N_21219,N_20994,N_20053);
nor U21220 (N_21220,N_20170,N_20802);
or U21221 (N_21221,N_20493,N_20528);
or U21222 (N_21222,N_20589,N_20365);
xor U21223 (N_21223,N_20613,N_20222);
nand U21224 (N_21224,N_20023,N_20852);
or U21225 (N_21225,N_20476,N_20704);
and U21226 (N_21226,N_20141,N_20340);
nor U21227 (N_21227,N_20386,N_20007);
xor U21228 (N_21228,N_20290,N_20433);
or U21229 (N_21229,N_20435,N_20738);
and U21230 (N_21230,N_20226,N_20001);
and U21231 (N_21231,N_20934,N_20068);
xor U21232 (N_21232,N_20501,N_20224);
nand U21233 (N_21233,N_20627,N_20440);
nand U21234 (N_21234,N_20478,N_20760);
nor U21235 (N_21235,N_20770,N_20427);
nor U21236 (N_21236,N_20110,N_20559);
and U21237 (N_21237,N_20851,N_20882);
xnor U21238 (N_21238,N_20763,N_20360);
or U21239 (N_21239,N_20039,N_20327);
nor U21240 (N_21240,N_20344,N_20474);
xor U21241 (N_21241,N_20794,N_20667);
nor U21242 (N_21242,N_20877,N_20698);
or U21243 (N_21243,N_20354,N_20793);
and U21244 (N_21244,N_20761,N_20377);
xor U21245 (N_21245,N_20525,N_20372);
xnor U21246 (N_21246,N_20415,N_20105);
xnor U21247 (N_21247,N_20809,N_20585);
nor U21248 (N_21248,N_20494,N_20935);
xnor U21249 (N_21249,N_20387,N_20757);
xnor U21250 (N_21250,N_20527,N_20065);
and U21251 (N_21251,N_20218,N_20009);
or U21252 (N_21252,N_20034,N_20699);
nand U21253 (N_21253,N_20785,N_20454);
nor U21254 (N_21254,N_20002,N_20672);
and U21255 (N_21255,N_20921,N_20347);
xor U21256 (N_21256,N_20610,N_20629);
and U21257 (N_21257,N_20526,N_20482);
nor U21258 (N_21258,N_20941,N_20810);
nor U21259 (N_21259,N_20833,N_20018);
and U21260 (N_21260,N_20359,N_20089);
nor U21261 (N_21261,N_20725,N_20341);
nor U21262 (N_21262,N_20499,N_20148);
xor U21263 (N_21263,N_20876,N_20428);
nand U21264 (N_21264,N_20179,N_20130);
and U21265 (N_21265,N_20533,N_20576);
or U21266 (N_21266,N_20106,N_20216);
nand U21267 (N_21267,N_20331,N_20198);
and U21268 (N_21268,N_20026,N_20439);
and U21269 (N_21269,N_20918,N_20711);
or U21270 (N_21270,N_20787,N_20872);
xnor U21271 (N_21271,N_20055,N_20562);
and U21272 (N_21272,N_20147,N_20575);
or U21273 (N_21273,N_20606,N_20355);
and U21274 (N_21274,N_20658,N_20334);
and U21275 (N_21275,N_20773,N_20343);
xnor U21276 (N_21276,N_20927,N_20306);
xor U21277 (N_21277,N_20969,N_20979);
or U21278 (N_21278,N_20998,N_20453);
or U21279 (N_21279,N_20300,N_20070);
xnor U21280 (N_21280,N_20600,N_20520);
xnor U21281 (N_21281,N_20312,N_20408);
xnor U21282 (N_21282,N_20900,N_20914);
nor U21283 (N_21283,N_20133,N_20283);
xor U21284 (N_21284,N_20817,N_20964);
and U21285 (N_21285,N_20052,N_20776);
xor U21286 (N_21286,N_20630,N_20871);
nor U21287 (N_21287,N_20088,N_20837);
xnor U21288 (N_21288,N_20669,N_20788);
nor U21289 (N_21289,N_20828,N_20339);
or U21290 (N_21290,N_20470,N_20705);
xor U21291 (N_21291,N_20583,N_20128);
xnor U21292 (N_21292,N_20205,N_20812);
nand U21293 (N_21293,N_20165,N_20362);
nand U21294 (N_21294,N_20135,N_20958);
and U21295 (N_21295,N_20995,N_20572);
nor U21296 (N_21296,N_20206,N_20929);
nand U21297 (N_21297,N_20721,N_20514);
and U21298 (N_21298,N_20771,N_20338);
nand U21299 (N_21299,N_20369,N_20204);
xnor U21300 (N_21300,N_20990,N_20229);
or U21301 (N_21301,N_20868,N_20345);
and U21302 (N_21302,N_20093,N_20710);
and U21303 (N_21303,N_20701,N_20176);
or U21304 (N_21304,N_20521,N_20716);
nand U21305 (N_21305,N_20294,N_20543);
or U21306 (N_21306,N_20603,N_20966);
xor U21307 (N_21307,N_20336,N_20942);
nand U21308 (N_21308,N_20594,N_20111);
nor U21309 (N_21309,N_20733,N_20790);
xor U21310 (N_21310,N_20848,N_20405);
nand U21311 (N_21311,N_20724,N_20485);
and U21312 (N_21312,N_20840,N_20664);
nand U21313 (N_21313,N_20513,N_20310);
or U21314 (N_21314,N_20903,N_20436);
xor U21315 (N_21315,N_20281,N_20116);
nor U21316 (N_21316,N_20657,N_20292);
or U21317 (N_21317,N_20279,N_20611);
or U21318 (N_21318,N_20480,N_20560);
or U21319 (N_21319,N_20548,N_20012);
or U21320 (N_21320,N_20308,N_20090);
and U21321 (N_21321,N_20643,N_20194);
nor U21322 (N_21322,N_20781,N_20074);
xor U21323 (N_21323,N_20404,N_20239);
nand U21324 (N_21324,N_20910,N_20319);
nand U21325 (N_21325,N_20061,N_20608);
nand U21326 (N_21326,N_20571,N_20835);
and U21327 (N_21327,N_20000,N_20577);
and U21328 (N_21328,N_20797,N_20517);
or U21329 (N_21329,N_20954,N_20676);
xor U21330 (N_21330,N_20646,N_20497);
nor U21331 (N_21331,N_20425,N_20568);
or U21332 (N_21332,N_20484,N_20598);
or U21333 (N_21333,N_20272,N_20980);
and U21334 (N_21334,N_20211,N_20463);
and U21335 (N_21335,N_20258,N_20815);
nand U21336 (N_21336,N_20553,N_20652);
nand U21337 (N_21337,N_20689,N_20905);
xor U21338 (N_21338,N_20475,N_20246);
nand U21339 (N_21339,N_20988,N_20045);
nor U21340 (N_21340,N_20261,N_20688);
and U21341 (N_21341,N_20832,N_20612);
xor U21342 (N_21342,N_20495,N_20768);
or U21343 (N_21343,N_20101,N_20171);
or U21344 (N_21344,N_20644,N_20581);
nor U21345 (N_21345,N_20846,N_20920);
nand U21346 (N_21346,N_20955,N_20490);
and U21347 (N_21347,N_20567,N_20256);
and U21348 (N_21348,N_20880,N_20058);
nand U21349 (N_21349,N_20556,N_20429);
or U21350 (N_21350,N_20251,N_20177);
or U21351 (N_21351,N_20342,N_20032);
nand U21352 (N_21352,N_20488,N_20795);
and U21353 (N_21353,N_20625,N_20238);
xor U21354 (N_21354,N_20371,N_20394);
nand U21355 (N_21355,N_20924,N_20512);
nor U21356 (N_21356,N_20057,N_20073);
and U21357 (N_21357,N_20808,N_20621);
xnor U21358 (N_21358,N_20412,N_20959);
and U21359 (N_21359,N_20496,N_20438);
nand U21360 (N_21360,N_20730,N_20388);
nand U21361 (N_21361,N_20653,N_20280);
xnor U21362 (N_21362,N_20691,N_20582);
xnor U21363 (N_21363,N_20200,N_20249);
nor U21364 (N_21364,N_20648,N_20765);
and U21365 (N_21365,N_20071,N_20951);
nor U21366 (N_21366,N_20233,N_20353);
nand U21367 (N_21367,N_20378,N_20221);
xnor U21368 (N_21368,N_20385,N_20913);
and U21369 (N_21369,N_20040,N_20051);
nand U21370 (N_21370,N_20853,N_20444);
nor U21371 (N_21371,N_20767,N_20708);
and U21372 (N_21372,N_20885,N_20291);
and U21373 (N_21373,N_20168,N_20448);
nor U21374 (N_21374,N_20516,N_20740);
xor U21375 (N_21375,N_20411,N_20072);
nor U21376 (N_21376,N_20477,N_20956);
nor U21377 (N_21377,N_20870,N_20682);
nand U21378 (N_21378,N_20430,N_20622);
nor U21379 (N_21379,N_20356,N_20786);
nand U21380 (N_21380,N_20859,N_20465);
and U21381 (N_21381,N_20014,N_20932);
nand U21382 (N_21382,N_20234,N_20373);
nand U21383 (N_21383,N_20749,N_20094);
and U21384 (N_21384,N_20114,N_20931);
xnor U21385 (N_21385,N_20991,N_20457);
and U21386 (N_21386,N_20230,N_20120);
nand U21387 (N_21387,N_20690,N_20623);
nor U21388 (N_21388,N_20191,N_20938);
nand U21389 (N_21389,N_20481,N_20208);
nand U21390 (N_21390,N_20747,N_20121);
nor U21391 (N_21391,N_20973,N_20118);
xnor U21392 (N_21392,N_20169,N_20789);
nand U21393 (N_21393,N_20296,N_20467);
and U21394 (N_21394,N_20717,N_20928);
or U21395 (N_21395,N_20017,N_20139);
or U21396 (N_21396,N_20466,N_20968);
or U21397 (N_21397,N_20615,N_20145);
and U21398 (N_21398,N_20049,N_20737);
nor U21399 (N_21399,N_20161,N_20129);
xnor U21400 (N_21400,N_20182,N_20887);
xor U21401 (N_21401,N_20271,N_20149);
and U21402 (N_21402,N_20069,N_20554);
or U21403 (N_21403,N_20534,N_20117);
nand U21404 (N_21404,N_20303,N_20464);
xor U21405 (N_21405,N_20487,N_20822);
or U21406 (N_21406,N_20008,N_20048);
or U21407 (N_21407,N_20649,N_20739);
xnor U21408 (N_21408,N_20687,N_20174);
and U21409 (N_21409,N_20441,N_20946);
or U21410 (N_21410,N_20083,N_20661);
or U21411 (N_21411,N_20309,N_20214);
or U21412 (N_21412,N_20807,N_20626);
nor U21413 (N_21413,N_20243,N_20908);
or U21414 (N_21414,N_20143,N_20159);
nor U21415 (N_21415,N_20046,N_20421);
nor U21416 (N_21416,N_20890,N_20366);
or U21417 (N_21417,N_20806,N_20060);
or U21418 (N_21418,N_20565,N_20671);
nand U21419 (N_21419,N_20769,N_20253);
nor U21420 (N_21420,N_20166,N_20845);
nand U21421 (N_21421,N_20884,N_20937);
nor U21422 (N_21422,N_20712,N_20403);
nand U21423 (N_21423,N_20975,N_20778);
and U21424 (N_21424,N_20273,N_20086);
nor U21425 (N_21425,N_20943,N_20957);
xor U21426 (N_21426,N_20573,N_20037);
or U21427 (N_21427,N_20392,N_20564);
and U21428 (N_21428,N_20108,N_20591);
nand U21429 (N_21429,N_20266,N_20349);
or U21430 (N_21430,N_20507,N_20796);
xnor U21431 (N_21431,N_20298,N_20054);
nor U21432 (N_21432,N_20654,N_20452);
and U21433 (N_21433,N_20609,N_20217);
and U21434 (N_21434,N_20423,N_20660);
nor U21435 (N_21435,N_20138,N_20798);
and U21436 (N_21436,N_20983,N_20972);
and U21437 (N_21437,N_20659,N_20379);
xnor U21438 (N_21438,N_20674,N_20677);
nor U21439 (N_21439,N_20506,N_20358);
or U21440 (N_21440,N_20153,N_20035);
or U21441 (N_21441,N_20282,N_20673);
and U21442 (N_21442,N_20424,N_20492);
and U21443 (N_21443,N_20926,N_20285);
or U21444 (N_21444,N_20109,N_20357);
and U21445 (N_21445,N_20220,N_20505);
nand U21446 (N_21446,N_20140,N_20666);
or U21447 (N_21447,N_20451,N_20758);
and U21448 (N_21448,N_20850,N_20381);
or U21449 (N_21449,N_20584,N_20019);
and U21450 (N_21450,N_20662,N_20670);
nor U21451 (N_21451,N_20706,N_20650);
nor U21452 (N_21452,N_20624,N_20982);
and U21453 (N_21453,N_20901,N_20842);
nor U21454 (N_21454,N_20297,N_20540);
and U21455 (N_21455,N_20270,N_20974);
and U21456 (N_21456,N_20713,N_20586);
nor U21457 (N_21457,N_20199,N_20555);
nor U21458 (N_21458,N_20115,N_20590);
xor U21459 (N_21459,N_20899,N_20697);
and U21460 (N_21460,N_20157,N_20335);
xnor U21461 (N_21461,N_20132,N_20158);
or U21462 (N_21462,N_20727,N_20383);
and U21463 (N_21463,N_20826,N_20374);
nand U21464 (N_21464,N_20818,N_20746);
and U21465 (N_21465,N_20825,N_20459);
and U21466 (N_21466,N_20190,N_20255);
or U21467 (N_21467,N_20013,N_20445);
xor U21468 (N_21468,N_20419,N_20811);
nor U21469 (N_21469,N_20265,N_20819);
and U21470 (N_21470,N_20180,N_20547);
nand U21471 (N_21471,N_20580,N_20695);
nand U21472 (N_21472,N_20315,N_20894);
nand U21473 (N_21473,N_20557,N_20364);
xor U21474 (N_21474,N_20152,N_20102);
nor U21475 (N_21475,N_20006,N_20544);
nor U21476 (N_21476,N_20192,N_20099);
and U21477 (N_21477,N_20692,N_20542);
and U21478 (N_21478,N_20398,N_20085);
and U21479 (N_21479,N_20410,N_20473);
xor U21480 (N_21480,N_20092,N_20456);
xnor U21481 (N_21481,N_20869,N_20592);
nor U21482 (N_21482,N_20080,N_20823);
xor U21483 (N_21483,N_20260,N_20511);
nor U21484 (N_21484,N_20081,N_20774);
and U21485 (N_21485,N_20113,N_20240);
nor U21486 (N_21486,N_20821,N_20134);
or U21487 (N_21487,N_20301,N_20936);
nand U21488 (N_21488,N_20714,N_20207);
nand U21489 (N_21489,N_20097,N_20570);
or U21490 (N_21490,N_20460,N_20098);
or U21491 (N_21491,N_20351,N_20031);
xnor U21492 (N_21492,N_20278,N_20389);
nand U21493 (N_21493,N_20245,N_20119);
xnor U21494 (N_21494,N_20741,N_20839);
nor U21495 (N_21495,N_20949,N_20067);
xnor U21496 (N_21496,N_20950,N_20352);
xor U21497 (N_21497,N_20304,N_20912);
or U21498 (N_21498,N_20178,N_20368);
nor U21499 (N_21499,N_20103,N_20766);
nor U21500 (N_21500,N_20971,N_20138);
or U21501 (N_21501,N_20520,N_20708);
or U21502 (N_21502,N_20344,N_20069);
nor U21503 (N_21503,N_20832,N_20071);
or U21504 (N_21504,N_20208,N_20927);
nand U21505 (N_21505,N_20208,N_20913);
xnor U21506 (N_21506,N_20590,N_20999);
and U21507 (N_21507,N_20528,N_20507);
nor U21508 (N_21508,N_20064,N_20799);
nand U21509 (N_21509,N_20993,N_20996);
xor U21510 (N_21510,N_20349,N_20372);
and U21511 (N_21511,N_20144,N_20524);
nand U21512 (N_21512,N_20036,N_20925);
nand U21513 (N_21513,N_20504,N_20754);
nor U21514 (N_21514,N_20742,N_20593);
and U21515 (N_21515,N_20739,N_20316);
or U21516 (N_21516,N_20723,N_20804);
or U21517 (N_21517,N_20173,N_20390);
nor U21518 (N_21518,N_20218,N_20811);
xnor U21519 (N_21519,N_20449,N_20420);
or U21520 (N_21520,N_20160,N_20032);
and U21521 (N_21521,N_20725,N_20072);
or U21522 (N_21522,N_20170,N_20267);
nor U21523 (N_21523,N_20359,N_20714);
or U21524 (N_21524,N_20088,N_20537);
xnor U21525 (N_21525,N_20019,N_20388);
nand U21526 (N_21526,N_20418,N_20107);
and U21527 (N_21527,N_20881,N_20876);
and U21528 (N_21528,N_20182,N_20230);
nor U21529 (N_21529,N_20786,N_20832);
nand U21530 (N_21530,N_20223,N_20206);
and U21531 (N_21531,N_20235,N_20956);
nor U21532 (N_21532,N_20120,N_20319);
nor U21533 (N_21533,N_20677,N_20435);
and U21534 (N_21534,N_20446,N_20394);
nand U21535 (N_21535,N_20179,N_20510);
xnor U21536 (N_21536,N_20019,N_20358);
nor U21537 (N_21537,N_20604,N_20833);
nor U21538 (N_21538,N_20078,N_20488);
and U21539 (N_21539,N_20037,N_20123);
and U21540 (N_21540,N_20031,N_20842);
xnor U21541 (N_21541,N_20135,N_20166);
nor U21542 (N_21542,N_20753,N_20121);
xor U21543 (N_21543,N_20901,N_20297);
nand U21544 (N_21544,N_20319,N_20460);
nor U21545 (N_21545,N_20920,N_20405);
nand U21546 (N_21546,N_20415,N_20446);
xor U21547 (N_21547,N_20728,N_20119);
xnor U21548 (N_21548,N_20756,N_20147);
and U21549 (N_21549,N_20344,N_20303);
and U21550 (N_21550,N_20089,N_20038);
nand U21551 (N_21551,N_20185,N_20134);
or U21552 (N_21552,N_20356,N_20809);
xnor U21553 (N_21553,N_20188,N_20700);
or U21554 (N_21554,N_20437,N_20110);
or U21555 (N_21555,N_20520,N_20093);
or U21556 (N_21556,N_20917,N_20739);
nor U21557 (N_21557,N_20977,N_20554);
xor U21558 (N_21558,N_20153,N_20156);
and U21559 (N_21559,N_20917,N_20984);
nor U21560 (N_21560,N_20920,N_20456);
nor U21561 (N_21561,N_20652,N_20945);
or U21562 (N_21562,N_20779,N_20498);
xor U21563 (N_21563,N_20925,N_20874);
nand U21564 (N_21564,N_20965,N_20610);
xor U21565 (N_21565,N_20309,N_20510);
and U21566 (N_21566,N_20830,N_20825);
and U21567 (N_21567,N_20347,N_20700);
or U21568 (N_21568,N_20003,N_20557);
or U21569 (N_21569,N_20092,N_20779);
and U21570 (N_21570,N_20564,N_20537);
nand U21571 (N_21571,N_20739,N_20378);
or U21572 (N_21572,N_20298,N_20377);
or U21573 (N_21573,N_20821,N_20143);
xor U21574 (N_21574,N_20098,N_20626);
xor U21575 (N_21575,N_20919,N_20698);
xor U21576 (N_21576,N_20993,N_20792);
xor U21577 (N_21577,N_20669,N_20854);
nand U21578 (N_21578,N_20403,N_20676);
nor U21579 (N_21579,N_20878,N_20127);
xnor U21580 (N_21580,N_20696,N_20499);
xnor U21581 (N_21581,N_20033,N_20157);
and U21582 (N_21582,N_20900,N_20183);
nand U21583 (N_21583,N_20297,N_20607);
nor U21584 (N_21584,N_20747,N_20778);
nand U21585 (N_21585,N_20042,N_20917);
nand U21586 (N_21586,N_20412,N_20154);
or U21587 (N_21587,N_20549,N_20664);
xor U21588 (N_21588,N_20284,N_20243);
nand U21589 (N_21589,N_20362,N_20487);
or U21590 (N_21590,N_20572,N_20405);
xor U21591 (N_21591,N_20199,N_20119);
xor U21592 (N_21592,N_20855,N_20545);
nand U21593 (N_21593,N_20631,N_20010);
nor U21594 (N_21594,N_20063,N_20290);
xor U21595 (N_21595,N_20237,N_20249);
and U21596 (N_21596,N_20455,N_20258);
nor U21597 (N_21597,N_20726,N_20909);
or U21598 (N_21598,N_20100,N_20110);
nor U21599 (N_21599,N_20223,N_20093);
and U21600 (N_21600,N_20400,N_20260);
and U21601 (N_21601,N_20348,N_20174);
and U21602 (N_21602,N_20748,N_20856);
and U21603 (N_21603,N_20034,N_20655);
and U21604 (N_21604,N_20349,N_20883);
or U21605 (N_21605,N_20755,N_20550);
xnor U21606 (N_21606,N_20313,N_20460);
nor U21607 (N_21607,N_20114,N_20555);
or U21608 (N_21608,N_20962,N_20920);
nor U21609 (N_21609,N_20194,N_20610);
nand U21610 (N_21610,N_20042,N_20419);
nor U21611 (N_21611,N_20747,N_20786);
xor U21612 (N_21612,N_20323,N_20458);
nor U21613 (N_21613,N_20205,N_20102);
xor U21614 (N_21614,N_20758,N_20237);
nor U21615 (N_21615,N_20111,N_20336);
or U21616 (N_21616,N_20467,N_20982);
or U21617 (N_21617,N_20321,N_20706);
nor U21618 (N_21618,N_20729,N_20366);
nor U21619 (N_21619,N_20787,N_20571);
nor U21620 (N_21620,N_20025,N_20112);
and U21621 (N_21621,N_20196,N_20727);
or U21622 (N_21622,N_20809,N_20906);
or U21623 (N_21623,N_20055,N_20519);
or U21624 (N_21624,N_20930,N_20985);
nand U21625 (N_21625,N_20749,N_20765);
or U21626 (N_21626,N_20999,N_20668);
nor U21627 (N_21627,N_20153,N_20524);
or U21628 (N_21628,N_20696,N_20448);
nand U21629 (N_21629,N_20604,N_20900);
and U21630 (N_21630,N_20224,N_20133);
nand U21631 (N_21631,N_20764,N_20791);
or U21632 (N_21632,N_20178,N_20093);
nor U21633 (N_21633,N_20434,N_20064);
xor U21634 (N_21634,N_20401,N_20846);
nor U21635 (N_21635,N_20390,N_20759);
nand U21636 (N_21636,N_20406,N_20622);
and U21637 (N_21637,N_20337,N_20580);
or U21638 (N_21638,N_20175,N_20065);
xor U21639 (N_21639,N_20493,N_20134);
and U21640 (N_21640,N_20880,N_20197);
or U21641 (N_21641,N_20790,N_20173);
or U21642 (N_21642,N_20774,N_20737);
nor U21643 (N_21643,N_20663,N_20830);
nor U21644 (N_21644,N_20683,N_20614);
and U21645 (N_21645,N_20302,N_20555);
or U21646 (N_21646,N_20870,N_20538);
xnor U21647 (N_21647,N_20096,N_20774);
xor U21648 (N_21648,N_20478,N_20972);
and U21649 (N_21649,N_20249,N_20836);
nor U21650 (N_21650,N_20023,N_20691);
xor U21651 (N_21651,N_20284,N_20682);
and U21652 (N_21652,N_20159,N_20511);
nand U21653 (N_21653,N_20741,N_20426);
xor U21654 (N_21654,N_20471,N_20727);
xnor U21655 (N_21655,N_20358,N_20490);
nand U21656 (N_21656,N_20537,N_20647);
xor U21657 (N_21657,N_20752,N_20323);
and U21658 (N_21658,N_20459,N_20349);
or U21659 (N_21659,N_20975,N_20421);
nor U21660 (N_21660,N_20082,N_20959);
xor U21661 (N_21661,N_20772,N_20477);
xor U21662 (N_21662,N_20241,N_20674);
and U21663 (N_21663,N_20292,N_20922);
and U21664 (N_21664,N_20098,N_20527);
nand U21665 (N_21665,N_20396,N_20253);
and U21666 (N_21666,N_20495,N_20507);
nor U21667 (N_21667,N_20047,N_20056);
or U21668 (N_21668,N_20611,N_20987);
nor U21669 (N_21669,N_20063,N_20467);
xnor U21670 (N_21670,N_20622,N_20377);
and U21671 (N_21671,N_20318,N_20361);
xor U21672 (N_21672,N_20585,N_20477);
nor U21673 (N_21673,N_20003,N_20501);
nor U21674 (N_21674,N_20649,N_20947);
xnor U21675 (N_21675,N_20759,N_20910);
nor U21676 (N_21676,N_20044,N_20486);
nor U21677 (N_21677,N_20501,N_20712);
and U21678 (N_21678,N_20651,N_20196);
and U21679 (N_21679,N_20465,N_20726);
and U21680 (N_21680,N_20652,N_20136);
or U21681 (N_21681,N_20256,N_20058);
xnor U21682 (N_21682,N_20995,N_20567);
or U21683 (N_21683,N_20473,N_20621);
xor U21684 (N_21684,N_20329,N_20487);
nand U21685 (N_21685,N_20811,N_20061);
and U21686 (N_21686,N_20796,N_20475);
xnor U21687 (N_21687,N_20320,N_20670);
nand U21688 (N_21688,N_20608,N_20607);
or U21689 (N_21689,N_20443,N_20243);
xor U21690 (N_21690,N_20860,N_20014);
nand U21691 (N_21691,N_20960,N_20417);
or U21692 (N_21692,N_20212,N_20367);
nand U21693 (N_21693,N_20470,N_20329);
xor U21694 (N_21694,N_20893,N_20263);
nand U21695 (N_21695,N_20117,N_20207);
and U21696 (N_21696,N_20523,N_20553);
or U21697 (N_21697,N_20255,N_20217);
or U21698 (N_21698,N_20238,N_20313);
and U21699 (N_21699,N_20751,N_20366);
nor U21700 (N_21700,N_20820,N_20011);
nor U21701 (N_21701,N_20695,N_20039);
xnor U21702 (N_21702,N_20097,N_20952);
nand U21703 (N_21703,N_20764,N_20695);
or U21704 (N_21704,N_20584,N_20919);
nand U21705 (N_21705,N_20434,N_20021);
or U21706 (N_21706,N_20263,N_20528);
xnor U21707 (N_21707,N_20584,N_20382);
xor U21708 (N_21708,N_20765,N_20266);
xor U21709 (N_21709,N_20910,N_20133);
or U21710 (N_21710,N_20880,N_20865);
nand U21711 (N_21711,N_20492,N_20775);
and U21712 (N_21712,N_20381,N_20375);
and U21713 (N_21713,N_20007,N_20403);
xor U21714 (N_21714,N_20182,N_20544);
or U21715 (N_21715,N_20919,N_20097);
xnor U21716 (N_21716,N_20508,N_20926);
and U21717 (N_21717,N_20489,N_20402);
xnor U21718 (N_21718,N_20640,N_20985);
nand U21719 (N_21719,N_20440,N_20544);
or U21720 (N_21720,N_20305,N_20797);
nor U21721 (N_21721,N_20902,N_20784);
or U21722 (N_21722,N_20252,N_20526);
nor U21723 (N_21723,N_20718,N_20169);
nor U21724 (N_21724,N_20675,N_20683);
nand U21725 (N_21725,N_20689,N_20046);
xor U21726 (N_21726,N_20615,N_20348);
nor U21727 (N_21727,N_20049,N_20406);
nor U21728 (N_21728,N_20870,N_20305);
nor U21729 (N_21729,N_20842,N_20832);
or U21730 (N_21730,N_20861,N_20770);
nand U21731 (N_21731,N_20187,N_20290);
nor U21732 (N_21732,N_20924,N_20859);
xor U21733 (N_21733,N_20295,N_20338);
nand U21734 (N_21734,N_20773,N_20893);
nor U21735 (N_21735,N_20971,N_20150);
xor U21736 (N_21736,N_20972,N_20057);
xor U21737 (N_21737,N_20314,N_20324);
or U21738 (N_21738,N_20753,N_20327);
or U21739 (N_21739,N_20952,N_20445);
or U21740 (N_21740,N_20063,N_20660);
and U21741 (N_21741,N_20812,N_20894);
nor U21742 (N_21742,N_20410,N_20317);
nand U21743 (N_21743,N_20408,N_20908);
nor U21744 (N_21744,N_20989,N_20161);
or U21745 (N_21745,N_20054,N_20880);
and U21746 (N_21746,N_20771,N_20141);
xor U21747 (N_21747,N_20418,N_20563);
nand U21748 (N_21748,N_20529,N_20407);
or U21749 (N_21749,N_20930,N_20221);
nand U21750 (N_21750,N_20384,N_20858);
xnor U21751 (N_21751,N_20645,N_20549);
or U21752 (N_21752,N_20981,N_20773);
xor U21753 (N_21753,N_20516,N_20131);
and U21754 (N_21754,N_20637,N_20614);
or U21755 (N_21755,N_20111,N_20256);
nor U21756 (N_21756,N_20597,N_20632);
nand U21757 (N_21757,N_20600,N_20815);
or U21758 (N_21758,N_20850,N_20872);
and U21759 (N_21759,N_20237,N_20659);
and U21760 (N_21760,N_20794,N_20399);
and U21761 (N_21761,N_20976,N_20449);
and U21762 (N_21762,N_20348,N_20082);
nand U21763 (N_21763,N_20692,N_20599);
and U21764 (N_21764,N_20835,N_20041);
and U21765 (N_21765,N_20791,N_20130);
and U21766 (N_21766,N_20987,N_20565);
and U21767 (N_21767,N_20297,N_20328);
and U21768 (N_21768,N_20237,N_20352);
nor U21769 (N_21769,N_20069,N_20867);
nand U21770 (N_21770,N_20597,N_20553);
and U21771 (N_21771,N_20232,N_20006);
and U21772 (N_21772,N_20613,N_20991);
and U21773 (N_21773,N_20724,N_20848);
and U21774 (N_21774,N_20993,N_20147);
nand U21775 (N_21775,N_20037,N_20859);
nor U21776 (N_21776,N_20361,N_20314);
nor U21777 (N_21777,N_20098,N_20173);
nor U21778 (N_21778,N_20515,N_20365);
xor U21779 (N_21779,N_20048,N_20734);
and U21780 (N_21780,N_20626,N_20148);
or U21781 (N_21781,N_20640,N_20518);
nand U21782 (N_21782,N_20036,N_20548);
xor U21783 (N_21783,N_20811,N_20808);
and U21784 (N_21784,N_20460,N_20627);
nor U21785 (N_21785,N_20283,N_20452);
or U21786 (N_21786,N_20838,N_20306);
or U21787 (N_21787,N_20497,N_20996);
nand U21788 (N_21788,N_20452,N_20345);
nor U21789 (N_21789,N_20912,N_20868);
xnor U21790 (N_21790,N_20898,N_20948);
nand U21791 (N_21791,N_20875,N_20149);
nor U21792 (N_21792,N_20209,N_20929);
xor U21793 (N_21793,N_20670,N_20932);
or U21794 (N_21794,N_20745,N_20118);
or U21795 (N_21795,N_20486,N_20869);
and U21796 (N_21796,N_20231,N_20936);
nor U21797 (N_21797,N_20400,N_20531);
xor U21798 (N_21798,N_20884,N_20742);
or U21799 (N_21799,N_20272,N_20421);
nor U21800 (N_21800,N_20318,N_20933);
or U21801 (N_21801,N_20633,N_20587);
nor U21802 (N_21802,N_20196,N_20895);
and U21803 (N_21803,N_20354,N_20678);
nand U21804 (N_21804,N_20467,N_20358);
and U21805 (N_21805,N_20678,N_20484);
xnor U21806 (N_21806,N_20370,N_20514);
and U21807 (N_21807,N_20502,N_20121);
or U21808 (N_21808,N_20160,N_20308);
or U21809 (N_21809,N_20711,N_20317);
and U21810 (N_21810,N_20928,N_20609);
nand U21811 (N_21811,N_20965,N_20452);
nand U21812 (N_21812,N_20903,N_20684);
or U21813 (N_21813,N_20877,N_20276);
or U21814 (N_21814,N_20895,N_20202);
and U21815 (N_21815,N_20825,N_20866);
and U21816 (N_21816,N_20819,N_20171);
nor U21817 (N_21817,N_20714,N_20462);
nor U21818 (N_21818,N_20024,N_20736);
nand U21819 (N_21819,N_20858,N_20141);
or U21820 (N_21820,N_20628,N_20347);
nor U21821 (N_21821,N_20640,N_20792);
nand U21822 (N_21822,N_20708,N_20063);
nand U21823 (N_21823,N_20785,N_20692);
xor U21824 (N_21824,N_20766,N_20278);
or U21825 (N_21825,N_20129,N_20753);
or U21826 (N_21826,N_20009,N_20108);
xor U21827 (N_21827,N_20466,N_20629);
xor U21828 (N_21828,N_20941,N_20767);
xnor U21829 (N_21829,N_20950,N_20429);
xor U21830 (N_21830,N_20615,N_20622);
or U21831 (N_21831,N_20324,N_20628);
or U21832 (N_21832,N_20282,N_20362);
or U21833 (N_21833,N_20417,N_20843);
or U21834 (N_21834,N_20597,N_20195);
nor U21835 (N_21835,N_20363,N_20968);
and U21836 (N_21836,N_20421,N_20590);
and U21837 (N_21837,N_20550,N_20800);
nand U21838 (N_21838,N_20366,N_20300);
and U21839 (N_21839,N_20444,N_20974);
and U21840 (N_21840,N_20391,N_20249);
or U21841 (N_21841,N_20220,N_20018);
nor U21842 (N_21842,N_20196,N_20340);
nand U21843 (N_21843,N_20614,N_20700);
nor U21844 (N_21844,N_20177,N_20910);
nand U21845 (N_21845,N_20511,N_20657);
or U21846 (N_21846,N_20920,N_20805);
nand U21847 (N_21847,N_20185,N_20018);
or U21848 (N_21848,N_20796,N_20580);
or U21849 (N_21849,N_20936,N_20487);
and U21850 (N_21850,N_20288,N_20942);
and U21851 (N_21851,N_20910,N_20080);
and U21852 (N_21852,N_20336,N_20541);
and U21853 (N_21853,N_20763,N_20856);
nand U21854 (N_21854,N_20968,N_20650);
or U21855 (N_21855,N_20570,N_20825);
and U21856 (N_21856,N_20498,N_20921);
or U21857 (N_21857,N_20432,N_20526);
xor U21858 (N_21858,N_20737,N_20197);
xnor U21859 (N_21859,N_20054,N_20099);
or U21860 (N_21860,N_20309,N_20988);
xnor U21861 (N_21861,N_20978,N_20028);
or U21862 (N_21862,N_20831,N_20674);
xnor U21863 (N_21863,N_20770,N_20668);
nor U21864 (N_21864,N_20694,N_20738);
nand U21865 (N_21865,N_20051,N_20457);
and U21866 (N_21866,N_20940,N_20173);
and U21867 (N_21867,N_20257,N_20441);
or U21868 (N_21868,N_20532,N_20023);
and U21869 (N_21869,N_20640,N_20149);
or U21870 (N_21870,N_20775,N_20972);
nand U21871 (N_21871,N_20972,N_20861);
nand U21872 (N_21872,N_20914,N_20832);
or U21873 (N_21873,N_20690,N_20988);
and U21874 (N_21874,N_20628,N_20888);
or U21875 (N_21875,N_20932,N_20377);
and U21876 (N_21876,N_20305,N_20540);
xnor U21877 (N_21877,N_20745,N_20949);
or U21878 (N_21878,N_20919,N_20594);
nand U21879 (N_21879,N_20930,N_20385);
and U21880 (N_21880,N_20555,N_20962);
or U21881 (N_21881,N_20762,N_20114);
or U21882 (N_21882,N_20556,N_20609);
nor U21883 (N_21883,N_20027,N_20891);
nand U21884 (N_21884,N_20278,N_20659);
or U21885 (N_21885,N_20211,N_20453);
or U21886 (N_21886,N_20690,N_20003);
nand U21887 (N_21887,N_20673,N_20067);
nand U21888 (N_21888,N_20052,N_20715);
or U21889 (N_21889,N_20204,N_20277);
or U21890 (N_21890,N_20971,N_20887);
nor U21891 (N_21891,N_20180,N_20380);
xor U21892 (N_21892,N_20324,N_20589);
nor U21893 (N_21893,N_20557,N_20127);
or U21894 (N_21894,N_20483,N_20950);
xor U21895 (N_21895,N_20255,N_20668);
nor U21896 (N_21896,N_20342,N_20175);
nand U21897 (N_21897,N_20773,N_20674);
and U21898 (N_21898,N_20328,N_20716);
xnor U21899 (N_21899,N_20320,N_20187);
and U21900 (N_21900,N_20320,N_20961);
or U21901 (N_21901,N_20422,N_20631);
nor U21902 (N_21902,N_20011,N_20611);
xor U21903 (N_21903,N_20474,N_20705);
and U21904 (N_21904,N_20825,N_20370);
nor U21905 (N_21905,N_20896,N_20929);
nor U21906 (N_21906,N_20979,N_20030);
and U21907 (N_21907,N_20895,N_20190);
nand U21908 (N_21908,N_20140,N_20677);
nor U21909 (N_21909,N_20586,N_20839);
xor U21910 (N_21910,N_20105,N_20823);
and U21911 (N_21911,N_20245,N_20410);
xnor U21912 (N_21912,N_20707,N_20090);
nand U21913 (N_21913,N_20696,N_20618);
nor U21914 (N_21914,N_20883,N_20385);
nand U21915 (N_21915,N_20738,N_20157);
nor U21916 (N_21916,N_20116,N_20804);
or U21917 (N_21917,N_20929,N_20567);
or U21918 (N_21918,N_20625,N_20717);
or U21919 (N_21919,N_20873,N_20806);
or U21920 (N_21920,N_20187,N_20830);
nand U21921 (N_21921,N_20325,N_20476);
nand U21922 (N_21922,N_20552,N_20441);
nor U21923 (N_21923,N_20036,N_20002);
or U21924 (N_21924,N_20794,N_20122);
nor U21925 (N_21925,N_20664,N_20346);
or U21926 (N_21926,N_20245,N_20587);
or U21927 (N_21927,N_20611,N_20844);
and U21928 (N_21928,N_20465,N_20851);
and U21929 (N_21929,N_20925,N_20276);
nand U21930 (N_21930,N_20793,N_20357);
or U21931 (N_21931,N_20905,N_20949);
or U21932 (N_21932,N_20721,N_20648);
and U21933 (N_21933,N_20723,N_20883);
nand U21934 (N_21934,N_20885,N_20770);
nor U21935 (N_21935,N_20064,N_20890);
and U21936 (N_21936,N_20747,N_20197);
or U21937 (N_21937,N_20664,N_20810);
or U21938 (N_21938,N_20246,N_20867);
nand U21939 (N_21939,N_20206,N_20572);
or U21940 (N_21940,N_20628,N_20499);
xor U21941 (N_21941,N_20713,N_20363);
nand U21942 (N_21942,N_20432,N_20081);
nand U21943 (N_21943,N_20640,N_20438);
nand U21944 (N_21944,N_20852,N_20499);
xor U21945 (N_21945,N_20039,N_20821);
and U21946 (N_21946,N_20323,N_20884);
and U21947 (N_21947,N_20112,N_20861);
nand U21948 (N_21948,N_20587,N_20469);
or U21949 (N_21949,N_20976,N_20352);
nor U21950 (N_21950,N_20108,N_20177);
nand U21951 (N_21951,N_20549,N_20994);
and U21952 (N_21952,N_20883,N_20801);
nor U21953 (N_21953,N_20096,N_20291);
nand U21954 (N_21954,N_20377,N_20398);
nor U21955 (N_21955,N_20470,N_20256);
nand U21956 (N_21956,N_20699,N_20980);
nor U21957 (N_21957,N_20789,N_20242);
and U21958 (N_21958,N_20969,N_20082);
or U21959 (N_21959,N_20550,N_20925);
nand U21960 (N_21960,N_20220,N_20894);
and U21961 (N_21961,N_20845,N_20408);
and U21962 (N_21962,N_20031,N_20893);
nand U21963 (N_21963,N_20149,N_20449);
nand U21964 (N_21964,N_20400,N_20752);
nand U21965 (N_21965,N_20924,N_20720);
or U21966 (N_21966,N_20020,N_20995);
nand U21967 (N_21967,N_20732,N_20421);
and U21968 (N_21968,N_20457,N_20925);
xnor U21969 (N_21969,N_20020,N_20287);
nor U21970 (N_21970,N_20580,N_20811);
or U21971 (N_21971,N_20638,N_20750);
and U21972 (N_21972,N_20779,N_20763);
nor U21973 (N_21973,N_20810,N_20491);
nand U21974 (N_21974,N_20219,N_20142);
or U21975 (N_21975,N_20119,N_20925);
or U21976 (N_21976,N_20558,N_20029);
nand U21977 (N_21977,N_20245,N_20762);
or U21978 (N_21978,N_20557,N_20322);
and U21979 (N_21979,N_20278,N_20944);
xnor U21980 (N_21980,N_20562,N_20643);
nor U21981 (N_21981,N_20848,N_20942);
and U21982 (N_21982,N_20244,N_20615);
xor U21983 (N_21983,N_20836,N_20380);
nor U21984 (N_21984,N_20863,N_20029);
or U21985 (N_21985,N_20871,N_20345);
nand U21986 (N_21986,N_20483,N_20461);
nor U21987 (N_21987,N_20701,N_20636);
nand U21988 (N_21988,N_20299,N_20715);
or U21989 (N_21989,N_20548,N_20255);
and U21990 (N_21990,N_20516,N_20708);
nor U21991 (N_21991,N_20887,N_20777);
nor U21992 (N_21992,N_20365,N_20190);
xor U21993 (N_21993,N_20669,N_20248);
nor U21994 (N_21994,N_20830,N_20222);
xnor U21995 (N_21995,N_20733,N_20277);
xor U21996 (N_21996,N_20304,N_20981);
and U21997 (N_21997,N_20136,N_20503);
xor U21998 (N_21998,N_20678,N_20145);
nand U21999 (N_21999,N_20300,N_20535);
xor U22000 (N_22000,N_21039,N_21422);
xnor U22001 (N_22001,N_21128,N_21226);
nand U22002 (N_22002,N_21471,N_21972);
or U22003 (N_22003,N_21136,N_21732);
or U22004 (N_22004,N_21088,N_21264);
and U22005 (N_22005,N_21238,N_21971);
and U22006 (N_22006,N_21416,N_21617);
nor U22007 (N_22007,N_21431,N_21442);
nand U22008 (N_22008,N_21190,N_21270);
xor U22009 (N_22009,N_21690,N_21480);
xor U22010 (N_22010,N_21433,N_21596);
xor U22011 (N_22011,N_21888,N_21944);
nor U22012 (N_22012,N_21445,N_21710);
nor U22013 (N_22013,N_21294,N_21542);
nand U22014 (N_22014,N_21257,N_21929);
and U22015 (N_22015,N_21462,N_21071);
xnor U22016 (N_22016,N_21811,N_21603);
and U22017 (N_22017,N_21218,N_21319);
or U22018 (N_22018,N_21403,N_21568);
xnor U22019 (N_22019,N_21530,N_21861);
nand U22020 (N_22020,N_21073,N_21463);
xor U22021 (N_22021,N_21395,N_21535);
and U22022 (N_22022,N_21460,N_21636);
nand U22023 (N_22023,N_21826,N_21897);
nand U22024 (N_22024,N_21814,N_21590);
nor U22025 (N_22025,N_21778,N_21178);
xnor U22026 (N_22026,N_21388,N_21056);
nor U22027 (N_22027,N_21261,N_21909);
nand U22028 (N_22028,N_21864,N_21585);
nand U22029 (N_22029,N_21827,N_21420);
xnor U22030 (N_22030,N_21657,N_21326);
nand U22031 (N_22031,N_21867,N_21127);
nor U22032 (N_22032,N_21608,N_21459);
nand U22033 (N_22033,N_21780,N_21225);
xnor U22034 (N_22034,N_21419,N_21993);
xnor U22035 (N_22035,N_21749,N_21974);
nand U22036 (N_22036,N_21032,N_21936);
nand U22037 (N_22037,N_21824,N_21072);
and U22038 (N_22038,N_21510,N_21671);
nand U22039 (N_22039,N_21878,N_21094);
nand U22040 (N_22040,N_21455,N_21833);
and U22041 (N_22041,N_21910,N_21432);
and U22042 (N_22042,N_21819,N_21044);
nand U22043 (N_22043,N_21777,N_21576);
nand U22044 (N_22044,N_21160,N_21231);
nor U22045 (N_22045,N_21076,N_21591);
or U22046 (N_22046,N_21805,N_21251);
xnor U22047 (N_22047,N_21447,N_21115);
nor U22048 (N_22048,N_21210,N_21499);
and U22049 (N_22049,N_21725,N_21075);
nor U22050 (N_22050,N_21383,N_21009);
and U22051 (N_22051,N_21120,N_21318);
nand U22052 (N_22052,N_21640,N_21730);
or U22053 (N_22053,N_21604,N_21900);
nor U22054 (N_22054,N_21047,N_21247);
xnor U22055 (N_22055,N_21742,N_21779);
nand U22056 (N_22056,N_21797,N_21293);
nor U22057 (N_22057,N_21611,N_21391);
nor U22058 (N_22058,N_21062,N_21298);
or U22059 (N_22059,N_21942,N_21299);
and U22060 (N_22060,N_21467,N_21731);
nand U22061 (N_22061,N_21052,N_21717);
xor U22062 (N_22062,N_21135,N_21667);
nand U22063 (N_22063,N_21557,N_21322);
or U22064 (N_22064,N_21818,N_21286);
nor U22065 (N_22065,N_21505,N_21172);
nor U22066 (N_22066,N_21143,N_21165);
nand U22067 (N_22067,N_21303,N_21453);
nor U22068 (N_22068,N_21110,N_21891);
nand U22069 (N_22069,N_21332,N_21243);
xnor U22070 (N_22070,N_21262,N_21368);
nor U22071 (N_22071,N_21567,N_21623);
xnor U22072 (N_22072,N_21968,N_21102);
or U22073 (N_22073,N_21022,N_21470);
or U22074 (N_22074,N_21171,N_21037);
and U22075 (N_22075,N_21830,N_21776);
nor U22076 (N_22076,N_21738,N_21089);
nand U22077 (N_22077,N_21950,N_21061);
or U22078 (N_22078,N_21847,N_21845);
xor U22079 (N_22079,N_21249,N_21650);
or U22080 (N_22080,N_21750,N_21028);
nand U22081 (N_22081,N_21869,N_21130);
and U22082 (N_22082,N_21843,N_21144);
xor U22083 (N_22083,N_21848,N_21441);
nor U22084 (N_22084,N_21131,N_21543);
nand U22085 (N_22085,N_21838,N_21464);
and U22086 (N_22086,N_21615,N_21158);
xor U22087 (N_22087,N_21578,N_21983);
or U22088 (N_22088,N_21343,N_21125);
and U22089 (N_22089,N_21469,N_21563);
or U22090 (N_22090,N_21266,N_21227);
xor U22091 (N_22091,N_21141,N_21182);
xnor U22092 (N_22092,N_21114,N_21381);
and U22093 (N_22093,N_21524,N_21870);
xnor U22094 (N_22094,N_21164,N_21356);
xnor U22095 (N_22095,N_21129,N_21877);
and U22096 (N_22096,N_21759,N_21862);
or U22097 (N_22097,N_21003,N_21452);
or U22098 (N_22098,N_21451,N_21450);
and U22099 (N_22099,N_21767,N_21336);
xor U22100 (N_22100,N_21309,N_21969);
and U22101 (N_22101,N_21021,N_21768);
nand U22102 (N_22102,N_21561,N_21612);
nand U22103 (N_22103,N_21979,N_21670);
nand U22104 (N_22104,N_21191,N_21770);
nand U22105 (N_22105,N_21137,N_21902);
xor U22106 (N_22106,N_21915,N_21526);
or U22107 (N_22107,N_21652,N_21747);
xnor U22108 (N_22108,N_21355,N_21019);
or U22109 (N_22109,N_21975,N_21173);
xor U22110 (N_22110,N_21560,N_21290);
nor U22111 (N_22111,N_21565,N_21562);
or U22112 (N_22112,N_21223,N_21256);
or U22113 (N_22113,N_21219,N_21651);
or U22114 (N_22114,N_21134,N_21523);
nor U22115 (N_22115,N_21539,N_21889);
and U22116 (N_22116,N_21289,N_21872);
or U22117 (N_22117,N_21001,N_21775);
nor U22118 (N_22118,N_21084,N_21895);
or U22119 (N_22119,N_21883,N_21914);
or U22120 (N_22120,N_21335,N_21438);
and U22121 (N_22121,N_21211,N_21609);
xnor U22122 (N_22122,N_21829,N_21534);
nand U22123 (N_22123,N_21796,N_21268);
xor U22124 (N_22124,N_21051,N_21554);
nand U22125 (N_22125,N_21132,N_21248);
xnor U22126 (N_22126,N_21588,N_21679);
nor U22127 (N_22127,N_21235,N_21366);
or U22128 (N_22128,N_21150,N_21834);
nand U22129 (N_22129,N_21879,N_21406);
nor U22130 (N_22130,N_21321,N_21116);
nand U22131 (N_22131,N_21372,N_21209);
xnor U22132 (N_22132,N_21297,N_21674);
xnor U22133 (N_22133,N_21720,N_21367);
xnor U22134 (N_22134,N_21040,N_21916);
nor U22135 (N_22135,N_21769,N_21295);
nand U22136 (N_22136,N_21077,N_21698);
and U22137 (N_22137,N_21569,N_21733);
and U22138 (N_22138,N_21746,N_21546);
nand U22139 (N_22139,N_21217,N_21798);
and U22140 (N_22140,N_21943,N_21186);
nor U22141 (N_22141,N_21736,N_21648);
or U22142 (N_22142,N_21058,N_21481);
or U22143 (N_22143,N_21204,N_21175);
xor U22144 (N_22144,N_21229,N_21232);
nand U22145 (N_22145,N_21146,N_21498);
xnor U22146 (N_22146,N_21390,N_21821);
xor U22147 (N_22147,N_21740,N_21709);
xor U22148 (N_22148,N_21766,N_21913);
nor U22149 (N_22149,N_21379,N_21506);
nand U22150 (N_22150,N_21296,N_21111);
nor U22151 (N_22151,N_21280,N_21387);
and U22152 (N_22152,N_21645,N_21624);
and U22153 (N_22153,N_21606,N_21091);
nor U22154 (N_22154,N_21068,N_21363);
or U22155 (N_22155,N_21788,N_21066);
xnor U22156 (N_22156,N_21435,N_21458);
and U22157 (N_22157,N_21378,N_21873);
and U22158 (N_22158,N_21189,N_21718);
nor U22159 (N_22159,N_21761,N_21728);
xor U22160 (N_22160,N_21820,N_21937);
and U22161 (N_22161,N_21904,N_21119);
nor U22162 (N_22162,N_21203,N_21347);
or U22163 (N_22163,N_21556,N_21785);
or U22164 (N_22164,N_21308,N_21491);
nor U22165 (N_22165,N_21493,N_21839);
and U22166 (N_22166,N_21465,N_21197);
and U22167 (N_22167,N_21985,N_21836);
nor U22168 (N_22168,N_21512,N_21919);
or U22169 (N_22169,N_21547,N_21933);
nand U22170 (N_22170,N_21553,N_21351);
and U22171 (N_22171,N_21448,N_21643);
nand U22172 (N_22172,N_21668,N_21314);
nor U22173 (N_22173,N_21274,N_21704);
nor U22174 (N_22174,N_21754,N_21349);
xnor U22175 (N_22175,N_21370,N_21016);
or U22176 (N_22176,N_21188,N_21622);
and U22177 (N_22177,N_21691,N_21067);
nor U22178 (N_22178,N_21927,N_21517);
or U22179 (N_22179,N_21564,N_21457);
and U22180 (N_22180,N_21685,N_21054);
nor U22181 (N_22181,N_21783,N_21147);
and U22182 (N_22182,N_21287,N_21267);
nand U22183 (N_22183,N_21017,N_21528);
nor U22184 (N_22184,N_21429,N_21315);
xor U22185 (N_22185,N_21988,N_21922);
nor U22186 (N_22186,N_21570,N_21206);
and U22187 (N_22187,N_21133,N_21398);
nor U22188 (N_22188,N_21959,N_21887);
nand U22189 (N_22189,N_21581,N_21311);
xor U22190 (N_22190,N_21680,N_21193);
nand U22191 (N_22191,N_21616,N_21896);
xor U22192 (N_22192,N_21036,N_21572);
xnor U22193 (N_22193,N_21678,N_21857);
and U22194 (N_22194,N_21817,N_21509);
xor U22195 (N_22195,N_21377,N_21781);
nor U22196 (N_22196,N_21940,N_21216);
xnor U22197 (N_22197,N_21882,N_21810);
xor U22198 (N_22198,N_21236,N_21245);
xor U22199 (N_22199,N_21283,N_21664);
nor U22200 (N_22200,N_21350,N_21105);
and U22201 (N_22201,N_21330,N_21487);
and U22202 (N_22202,N_21239,N_21333);
and U22203 (N_22203,N_21756,N_21014);
xnor U22204 (N_22204,N_21962,N_21874);
or U22205 (N_22205,N_21418,N_21276);
nor U22206 (N_22206,N_21537,N_21584);
or U22207 (N_22207,N_21174,N_21694);
nand U22208 (N_22208,N_21575,N_21104);
nand U22209 (N_22209,N_21697,N_21577);
nor U22210 (N_22210,N_21007,N_21400);
and U22211 (N_22211,N_21426,N_21010);
xor U22212 (N_22212,N_21832,N_21026);
nor U22213 (N_22213,N_21707,N_21855);
and U22214 (N_22214,N_21923,N_21573);
and U22215 (N_22215,N_21373,N_21894);
or U22216 (N_22216,N_21515,N_21346);
nand U22217 (N_22217,N_21637,N_21275);
or U22218 (N_22218,N_21514,N_21414);
nor U22219 (N_22219,N_21307,N_21109);
or U22220 (N_22220,N_21835,N_21170);
or U22221 (N_22221,N_21316,N_21151);
nand U22222 (N_22222,N_21952,N_21719);
nor U22223 (N_22223,N_21748,N_21233);
nor U22224 (N_22224,N_21853,N_21662);
or U22225 (N_22225,N_21486,N_21508);
nand U22226 (N_22226,N_21804,N_21163);
nor U22227 (N_22227,N_21503,N_21729);
nand U22228 (N_22228,N_21686,N_21153);
nand U22229 (N_22229,N_21329,N_21661);
and U22230 (N_22230,N_21434,N_21574);
xnor U22231 (N_22231,N_21908,N_21083);
or U22232 (N_22232,N_21986,N_21989);
nor U22233 (N_22233,N_21866,N_21477);
nor U22234 (N_22234,N_21790,N_21361);
xor U22235 (N_22235,N_21284,N_21237);
nor U22236 (N_22236,N_21187,N_21034);
and U22237 (N_22237,N_21483,N_21000);
and U22238 (N_22238,N_21589,N_21166);
and U22239 (N_22239,N_21113,N_21982);
and U22240 (N_22240,N_21757,N_21774);
nor U22241 (N_22241,N_21744,N_21389);
nand U22242 (N_22242,N_21080,N_21841);
and U22243 (N_22243,N_21254,N_21948);
or U22244 (N_22244,N_21846,N_21430);
nor U22245 (N_22245,N_21706,N_21352);
and U22246 (N_22246,N_21202,N_21328);
and U22247 (N_22247,N_21583,N_21384);
and U22248 (N_22248,N_21006,N_21939);
nand U22249 (N_22249,N_21946,N_21427);
and U22250 (N_22250,N_21550,N_21341);
xor U22251 (N_22251,N_21712,N_21890);
nand U22252 (N_22252,N_21721,N_21594);
and U22253 (N_22253,N_21148,N_21375);
nor U22254 (N_22254,N_21626,N_21123);
and U22255 (N_22255,N_21941,N_21527);
nand U22256 (N_22256,N_21259,N_21376);
and U22257 (N_22257,N_21302,N_21292);
nor U22258 (N_22258,N_21682,N_21644);
nor U22259 (N_22259,N_21100,N_21934);
nand U22260 (N_22260,N_21555,N_21997);
nand U22261 (N_22261,N_21152,N_21050);
and U22262 (N_22262,N_21029,N_21212);
and U22263 (N_22263,N_21789,N_21340);
and U22264 (N_22264,N_21437,N_21641);
and U22265 (N_22265,N_21250,N_21466);
nand U22266 (N_22266,N_21488,N_21758);
nand U22267 (N_22267,N_21126,N_21155);
and U22268 (N_22268,N_21064,N_21924);
nor U22269 (N_22269,N_21393,N_21911);
nor U22270 (N_22270,N_21639,N_21149);
nor U22271 (N_22271,N_21497,N_21207);
and U22272 (N_22272,N_21177,N_21899);
nor U22273 (N_22273,N_21802,N_21168);
xnor U22274 (N_22274,N_21522,N_21646);
and U22275 (N_22275,N_21038,N_21823);
nand U22276 (N_22276,N_21580,N_21921);
or U22277 (N_22277,N_21489,N_21693);
xnor U22278 (N_22278,N_21300,N_21199);
nor U22279 (N_22279,N_21753,N_21240);
and U22280 (N_22280,N_21404,N_21222);
and U22281 (N_22281,N_21004,N_21214);
xor U22282 (N_22282,N_21385,N_21196);
nand U22283 (N_22283,N_21593,N_21683);
nor U22284 (N_22284,N_21665,N_21525);
and U22285 (N_22285,N_21070,N_21765);
nor U22286 (N_22286,N_21042,N_21601);
nor U22287 (N_22287,N_21096,N_21192);
nand U22288 (N_22288,N_21184,N_21317);
and U22289 (N_22289,N_21912,N_21965);
or U22290 (N_22290,N_21041,N_21801);
nand U22291 (N_22291,N_21074,N_21030);
nor U22292 (N_22292,N_21673,N_21484);
and U22293 (N_22293,N_21439,N_21791);
and U22294 (N_22294,N_21529,N_21868);
nand U22295 (N_22295,N_21394,N_21279);
nor U22296 (N_22296,N_21195,N_21632);
nand U22297 (N_22297,N_21695,N_21500);
nor U22298 (N_22298,N_21666,N_21551);
or U22299 (N_22299,N_21476,N_21692);
and U22300 (N_22300,N_21099,N_21246);
or U22301 (N_22301,N_21025,N_21844);
or U22302 (N_22302,N_21945,N_21475);
xnor U22303 (N_22303,N_21610,N_21842);
and U22304 (N_22304,N_21806,N_21456);
or U22305 (N_22305,N_21424,N_21947);
nor U22306 (N_22306,N_21544,N_21715);
xnor U22307 (N_22307,N_21139,N_21359);
or U22308 (N_22308,N_21087,N_21627);
or U22309 (N_22309,N_21415,N_21230);
and U22310 (N_22310,N_21884,N_21122);
nor U22311 (N_22311,N_21677,N_21063);
nand U22312 (N_22312,N_21630,N_21023);
nand U22313 (N_22313,N_21957,N_21011);
or U22314 (N_22314,N_21002,N_21607);
or U22315 (N_22315,N_21600,N_21595);
nor U22316 (N_22316,N_21386,N_21371);
and U22317 (N_22317,N_21221,N_21271);
xnor U22318 (N_22318,N_21956,N_21048);
nand U22319 (N_22319,N_21306,N_21614);
nand U22320 (N_22320,N_21597,N_21005);
or U22321 (N_22321,N_21012,N_21468);
xnor U22322 (N_22322,N_21031,N_21713);
nand U22323 (N_22323,N_21324,N_21358);
xor U22324 (N_22324,N_21176,N_21540);
nor U22325 (N_22325,N_21278,N_21334);
xor U22326 (N_22326,N_21955,N_21440);
or U22327 (N_22327,N_21625,N_21331);
xnor U22328 (N_22328,N_21724,N_21490);
or U22329 (N_22329,N_21852,N_21812);
or U22330 (N_22330,N_21549,N_21885);
and U22331 (N_22331,N_21399,N_21185);
nor U22332 (N_22332,N_21531,N_21978);
xor U22333 (N_22333,N_21124,N_21980);
or U22334 (N_22334,N_21474,N_21635);
xnor U22335 (N_22335,N_21169,N_21320);
and U22336 (N_22336,N_21559,N_21984);
and U22337 (N_22337,N_21949,N_21587);
or U22338 (N_22338,N_21092,N_21545);
nor U22339 (N_22339,N_21208,N_21815);
nand U22340 (N_22340,N_21903,N_21473);
or U22341 (N_22341,N_21976,N_21252);
or U22342 (N_22342,N_21224,N_21504);
nor U22343 (N_22343,N_21716,N_21828);
or U22344 (N_22344,N_21773,N_21402);
and U22345 (N_22345,N_21881,N_21374);
nand U22346 (N_22346,N_21059,N_21620);
xnor U22347 (N_22347,N_21705,N_21858);
or U22348 (N_22348,N_21397,N_21258);
nor U22349 (N_22349,N_21215,N_21342);
nor U22350 (N_22350,N_21901,N_21495);
nor U22351 (N_22351,N_21755,N_21850);
xor U22352 (N_22352,N_21541,N_21327);
nand U22353 (N_22353,N_21931,N_21737);
nand U22354 (N_22354,N_21880,N_21837);
and U22355 (N_22355,N_21619,N_21689);
xnor U22356 (N_22356,N_21964,N_21069);
nand U22357 (N_22357,N_21288,N_21027);
nor U22358 (N_22358,N_21739,N_21521);
xor U22359 (N_22359,N_21145,N_21991);
or U22360 (N_22360,N_21323,N_21970);
nor U22361 (N_22361,N_21905,N_21095);
nor U22362 (N_22362,N_21702,N_21700);
or U22363 (N_22363,N_21886,N_21687);
nor U22364 (N_22364,N_21977,N_21813);
and U22365 (N_22365,N_21953,N_21408);
xnor U22366 (N_22366,N_21304,N_21472);
nand U22367 (N_22367,N_21461,N_21157);
xor U22368 (N_22368,N_21482,N_21772);
and U22369 (N_22369,N_21365,N_21660);
nor U22370 (N_22370,N_21325,N_21362);
and U22371 (N_22371,N_21856,N_21161);
nor U22372 (N_22372,N_21312,N_21180);
and U22373 (N_22373,N_21793,N_21140);
and U22374 (N_22374,N_21357,N_21795);
or U22375 (N_22375,N_21822,N_21263);
xnor U22376 (N_22376,N_21082,N_21995);
nor U22377 (N_22377,N_21935,N_21055);
nand U22378 (N_22378,N_21538,N_21436);
and U22379 (N_22379,N_21981,N_21876);
nor U22380 (N_22380,N_21078,N_21344);
nor U22381 (N_22381,N_21108,N_21727);
xnor U22382 (N_22382,N_21396,N_21380);
nor U22383 (N_22383,N_21851,N_21642);
nor U22384 (N_22384,N_21425,N_21726);
nand U22385 (N_22385,N_21338,N_21013);
or U22386 (N_22386,N_21998,N_21053);
nor U22387 (N_22387,N_21421,N_21183);
or U22388 (N_22388,N_21807,N_21518);
xnor U22389 (N_22389,N_21973,N_21684);
nand U22390 (N_22390,N_21444,N_21121);
and U22391 (N_22391,N_21631,N_21752);
or U22392 (N_22392,N_21443,N_21552);
xor U22393 (N_22393,N_21265,N_21722);
nand U22394 (N_22394,N_21057,N_21241);
and U22395 (N_22395,N_21782,N_21906);
and U22396 (N_22396,N_21519,N_21784);
nand U22397 (N_22397,N_21696,N_21808);
or U22398 (N_22398,N_21951,N_21269);
nor U22399 (N_22399,N_21106,N_21582);
nand U22400 (N_22400,N_21800,N_21162);
nor U22401 (N_22401,N_21961,N_21825);
nor U22402 (N_22402,N_21065,N_21649);
nor U22403 (N_22403,N_21198,N_21928);
nor U22404 (N_22404,N_21085,N_21741);
nor U22405 (N_22405,N_21272,N_21990);
nor U22406 (N_22406,N_21098,N_21138);
nor U22407 (N_22407,N_21656,N_21954);
xnor U22408 (N_22408,N_21996,N_21015);
nand U22409 (N_22409,N_21840,N_21967);
nand U22410 (N_22410,N_21167,N_21875);
or U22411 (N_22411,N_21413,N_21213);
xnor U22412 (N_22412,N_21994,N_21963);
nor U22413 (N_22413,N_21762,N_21405);
nor U22414 (N_22414,N_21865,N_21655);
or U22415 (N_22415,N_21502,N_21285);
or U22416 (N_22416,N_21485,N_21478);
nand U22417 (N_22417,N_21792,N_21745);
xor U22418 (N_22418,N_21479,N_21020);
nand U22419 (N_22419,N_21277,N_21703);
xnor U22420 (N_22420,N_21255,N_21107);
nor U22421 (N_22421,N_21764,N_21079);
and U22422 (N_22422,N_21658,N_21179);
or U22423 (N_22423,N_21310,N_21410);
and U22424 (N_22424,N_21699,N_21273);
nand U22425 (N_22425,N_21918,N_21253);
nand U22426 (N_22426,N_21787,N_21364);
or U22427 (N_22427,N_21220,N_21917);
and U22428 (N_22428,N_21926,N_21194);
and U22429 (N_22429,N_21494,N_21507);
xor U22430 (N_22430,N_21723,N_21060);
nor U22431 (N_22431,N_21409,N_21205);
and U22432 (N_22432,N_21859,N_21533);
nand U22433 (N_22433,N_21958,N_21743);
nor U22434 (N_22434,N_21401,N_21708);
xnor U22435 (N_22435,N_21392,N_21548);
xnor U22436 (N_22436,N_21860,N_21228);
xnor U22437 (N_22437,N_21676,N_21181);
nor U22438 (N_22438,N_21045,N_21907);
and U22439 (N_22439,N_21992,N_21628);
or U22440 (N_22440,N_21086,N_21669);
nor U22441 (N_22441,N_21871,N_21043);
nand U22442 (N_22442,N_21301,N_21313);
xor U22443 (N_22443,N_21681,N_21966);
nand U22444 (N_22444,N_21898,N_21751);
xor U22445 (N_22445,N_21033,N_21035);
xnor U22446 (N_22446,N_21663,N_21513);
nand U22447 (N_22447,N_21008,N_21282);
nor U22448 (N_22448,N_21339,N_21892);
nand U22449 (N_22449,N_21369,N_21714);
or U22450 (N_22450,N_21159,N_21849);
nor U22451 (N_22451,N_21605,N_21156);
or U22452 (N_22452,N_21960,N_21097);
nor U22453 (N_22453,N_21654,N_21496);
xor U22454 (N_22454,N_21794,N_21618);
and U22455 (N_22455,N_21659,N_21734);
xnor U22456 (N_22456,N_21647,N_21501);
nand U22457 (N_22457,N_21201,N_21348);
xor U22458 (N_22458,N_21999,N_21893);
xnor U22459 (N_22459,N_21532,N_21103);
xor U22460 (N_22460,N_21018,N_21200);
nand U22461 (N_22461,N_21799,N_21112);
nand U22462 (N_22462,N_21602,N_21423);
xnor U22463 (N_22463,N_21407,N_21154);
nand U22464 (N_22464,N_21621,N_21592);
nand U22465 (N_22465,N_21688,N_21599);
nand U22466 (N_22466,N_21516,N_21803);
nand U22467 (N_22467,N_21260,N_21711);
and U22468 (N_22468,N_21629,N_21354);
nor U22469 (N_22469,N_21417,N_21024);
xnor U22470 (N_22470,N_21831,N_21735);
and U22471 (N_22471,N_21816,N_21520);
xor U22472 (N_22472,N_21142,N_21586);
or U22473 (N_22473,N_21511,N_21987);
or U22474 (N_22474,N_21613,N_21566);
nand U22475 (N_22475,N_21454,N_21925);
nor U22476 (N_22476,N_21932,N_21049);
and U22477 (N_22477,N_21760,N_21633);
nor U22478 (N_22478,N_21492,N_21536);
nand U22479 (N_22479,N_21090,N_21337);
or U22480 (N_22480,N_21809,N_21411);
and U22481 (N_22481,N_21771,N_21345);
xnor U22482 (N_22482,N_21428,N_21446);
nor U22483 (N_22483,N_21938,N_21382);
xor U22484 (N_22484,N_21046,N_21242);
nor U22485 (N_22485,N_21786,N_21101);
nor U22486 (N_22486,N_21854,N_21675);
nor U22487 (N_22487,N_21360,N_21638);
or U22488 (N_22488,N_21672,N_21305);
and U22489 (N_22489,N_21863,N_21118);
or U22490 (N_22490,N_21117,N_21449);
or U22491 (N_22491,N_21634,N_21291);
or U22492 (N_22492,N_21093,N_21653);
nor U22493 (N_22493,N_21412,N_21930);
xor U22494 (N_22494,N_21558,N_21234);
xor U22495 (N_22495,N_21701,N_21920);
and U22496 (N_22496,N_21579,N_21081);
and U22497 (N_22497,N_21353,N_21763);
and U22498 (N_22498,N_21598,N_21281);
or U22499 (N_22499,N_21244,N_21571);
and U22500 (N_22500,N_21240,N_21707);
and U22501 (N_22501,N_21476,N_21469);
and U22502 (N_22502,N_21359,N_21434);
nand U22503 (N_22503,N_21503,N_21777);
xor U22504 (N_22504,N_21598,N_21296);
xor U22505 (N_22505,N_21031,N_21705);
xnor U22506 (N_22506,N_21860,N_21597);
nand U22507 (N_22507,N_21705,N_21677);
nor U22508 (N_22508,N_21691,N_21420);
and U22509 (N_22509,N_21068,N_21062);
nand U22510 (N_22510,N_21813,N_21237);
xnor U22511 (N_22511,N_21545,N_21340);
nand U22512 (N_22512,N_21700,N_21972);
nor U22513 (N_22513,N_21535,N_21460);
xor U22514 (N_22514,N_21327,N_21084);
nor U22515 (N_22515,N_21188,N_21509);
nor U22516 (N_22516,N_21786,N_21466);
and U22517 (N_22517,N_21977,N_21658);
xor U22518 (N_22518,N_21464,N_21772);
and U22519 (N_22519,N_21214,N_21242);
nand U22520 (N_22520,N_21585,N_21806);
xnor U22521 (N_22521,N_21363,N_21508);
xnor U22522 (N_22522,N_21423,N_21988);
nor U22523 (N_22523,N_21823,N_21327);
and U22524 (N_22524,N_21875,N_21649);
and U22525 (N_22525,N_21003,N_21033);
nor U22526 (N_22526,N_21931,N_21754);
or U22527 (N_22527,N_21769,N_21993);
nand U22528 (N_22528,N_21128,N_21985);
and U22529 (N_22529,N_21168,N_21908);
or U22530 (N_22530,N_21328,N_21376);
nand U22531 (N_22531,N_21589,N_21007);
nand U22532 (N_22532,N_21310,N_21368);
nand U22533 (N_22533,N_21759,N_21388);
xnor U22534 (N_22534,N_21426,N_21944);
or U22535 (N_22535,N_21395,N_21722);
or U22536 (N_22536,N_21613,N_21324);
nand U22537 (N_22537,N_21452,N_21875);
or U22538 (N_22538,N_21148,N_21220);
nand U22539 (N_22539,N_21516,N_21841);
nand U22540 (N_22540,N_21921,N_21119);
or U22541 (N_22541,N_21140,N_21825);
xor U22542 (N_22542,N_21665,N_21239);
and U22543 (N_22543,N_21495,N_21644);
xor U22544 (N_22544,N_21801,N_21763);
xnor U22545 (N_22545,N_21488,N_21688);
xor U22546 (N_22546,N_21626,N_21859);
or U22547 (N_22547,N_21135,N_21228);
or U22548 (N_22548,N_21206,N_21037);
xor U22549 (N_22549,N_21787,N_21576);
xnor U22550 (N_22550,N_21038,N_21882);
nor U22551 (N_22551,N_21559,N_21790);
and U22552 (N_22552,N_21464,N_21021);
nor U22553 (N_22553,N_21918,N_21498);
nand U22554 (N_22554,N_21506,N_21320);
xnor U22555 (N_22555,N_21562,N_21694);
nand U22556 (N_22556,N_21242,N_21112);
or U22557 (N_22557,N_21035,N_21011);
nand U22558 (N_22558,N_21852,N_21664);
and U22559 (N_22559,N_21490,N_21892);
and U22560 (N_22560,N_21292,N_21719);
nor U22561 (N_22561,N_21169,N_21560);
nand U22562 (N_22562,N_21399,N_21049);
and U22563 (N_22563,N_21011,N_21405);
xor U22564 (N_22564,N_21802,N_21155);
nand U22565 (N_22565,N_21934,N_21172);
or U22566 (N_22566,N_21539,N_21400);
nand U22567 (N_22567,N_21662,N_21430);
xor U22568 (N_22568,N_21707,N_21946);
nor U22569 (N_22569,N_21804,N_21783);
nor U22570 (N_22570,N_21243,N_21524);
and U22571 (N_22571,N_21775,N_21977);
nand U22572 (N_22572,N_21308,N_21530);
or U22573 (N_22573,N_21619,N_21734);
or U22574 (N_22574,N_21454,N_21430);
and U22575 (N_22575,N_21240,N_21935);
xor U22576 (N_22576,N_21307,N_21207);
and U22577 (N_22577,N_21284,N_21200);
or U22578 (N_22578,N_21426,N_21835);
xnor U22579 (N_22579,N_21572,N_21879);
xnor U22580 (N_22580,N_21554,N_21724);
nand U22581 (N_22581,N_21843,N_21706);
nor U22582 (N_22582,N_21035,N_21058);
xnor U22583 (N_22583,N_21700,N_21885);
xnor U22584 (N_22584,N_21977,N_21905);
xor U22585 (N_22585,N_21750,N_21865);
nand U22586 (N_22586,N_21344,N_21250);
and U22587 (N_22587,N_21553,N_21486);
nor U22588 (N_22588,N_21096,N_21727);
nand U22589 (N_22589,N_21507,N_21672);
nor U22590 (N_22590,N_21983,N_21255);
xnor U22591 (N_22591,N_21028,N_21538);
nand U22592 (N_22592,N_21913,N_21016);
and U22593 (N_22593,N_21074,N_21325);
nor U22594 (N_22594,N_21652,N_21539);
and U22595 (N_22595,N_21780,N_21682);
nor U22596 (N_22596,N_21350,N_21467);
nor U22597 (N_22597,N_21677,N_21289);
or U22598 (N_22598,N_21315,N_21489);
and U22599 (N_22599,N_21153,N_21339);
xnor U22600 (N_22600,N_21052,N_21480);
and U22601 (N_22601,N_21008,N_21451);
nand U22602 (N_22602,N_21640,N_21414);
or U22603 (N_22603,N_21298,N_21760);
or U22604 (N_22604,N_21811,N_21203);
or U22605 (N_22605,N_21228,N_21098);
nand U22606 (N_22606,N_21110,N_21908);
xor U22607 (N_22607,N_21157,N_21059);
xor U22608 (N_22608,N_21788,N_21362);
and U22609 (N_22609,N_21229,N_21112);
nor U22610 (N_22610,N_21692,N_21606);
or U22611 (N_22611,N_21917,N_21076);
and U22612 (N_22612,N_21708,N_21928);
and U22613 (N_22613,N_21451,N_21916);
and U22614 (N_22614,N_21082,N_21599);
and U22615 (N_22615,N_21219,N_21325);
nand U22616 (N_22616,N_21132,N_21819);
and U22617 (N_22617,N_21343,N_21094);
xor U22618 (N_22618,N_21065,N_21001);
xnor U22619 (N_22619,N_21015,N_21383);
nor U22620 (N_22620,N_21022,N_21162);
nor U22621 (N_22621,N_21577,N_21928);
and U22622 (N_22622,N_21859,N_21643);
and U22623 (N_22623,N_21630,N_21692);
xnor U22624 (N_22624,N_21796,N_21167);
or U22625 (N_22625,N_21453,N_21695);
nand U22626 (N_22626,N_21348,N_21619);
and U22627 (N_22627,N_21768,N_21851);
xnor U22628 (N_22628,N_21970,N_21881);
or U22629 (N_22629,N_21020,N_21220);
xor U22630 (N_22630,N_21310,N_21077);
or U22631 (N_22631,N_21408,N_21156);
nor U22632 (N_22632,N_21090,N_21195);
and U22633 (N_22633,N_21405,N_21771);
nand U22634 (N_22634,N_21984,N_21166);
and U22635 (N_22635,N_21801,N_21630);
xnor U22636 (N_22636,N_21358,N_21279);
xor U22637 (N_22637,N_21836,N_21167);
or U22638 (N_22638,N_21601,N_21384);
xor U22639 (N_22639,N_21052,N_21096);
nor U22640 (N_22640,N_21357,N_21452);
xor U22641 (N_22641,N_21998,N_21251);
xor U22642 (N_22642,N_21694,N_21840);
nor U22643 (N_22643,N_21794,N_21498);
or U22644 (N_22644,N_21809,N_21387);
or U22645 (N_22645,N_21344,N_21029);
nor U22646 (N_22646,N_21682,N_21081);
xnor U22647 (N_22647,N_21414,N_21673);
or U22648 (N_22648,N_21633,N_21673);
xor U22649 (N_22649,N_21698,N_21058);
or U22650 (N_22650,N_21371,N_21639);
or U22651 (N_22651,N_21631,N_21647);
and U22652 (N_22652,N_21355,N_21172);
and U22653 (N_22653,N_21078,N_21232);
or U22654 (N_22654,N_21727,N_21654);
nand U22655 (N_22655,N_21680,N_21851);
nor U22656 (N_22656,N_21278,N_21865);
nor U22657 (N_22657,N_21151,N_21932);
or U22658 (N_22658,N_21732,N_21101);
and U22659 (N_22659,N_21070,N_21120);
and U22660 (N_22660,N_21706,N_21336);
and U22661 (N_22661,N_21604,N_21601);
nor U22662 (N_22662,N_21967,N_21538);
nor U22663 (N_22663,N_21897,N_21409);
or U22664 (N_22664,N_21375,N_21423);
and U22665 (N_22665,N_21185,N_21652);
or U22666 (N_22666,N_21538,N_21876);
nand U22667 (N_22667,N_21892,N_21207);
nand U22668 (N_22668,N_21816,N_21993);
nor U22669 (N_22669,N_21677,N_21374);
nor U22670 (N_22670,N_21763,N_21761);
nor U22671 (N_22671,N_21260,N_21241);
and U22672 (N_22672,N_21607,N_21230);
nor U22673 (N_22673,N_21547,N_21192);
nor U22674 (N_22674,N_21527,N_21816);
nor U22675 (N_22675,N_21257,N_21478);
and U22676 (N_22676,N_21770,N_21653);
nand U22677 (N_22677,N_21442,N_21096);
or U22678 (N_22678,N_21081,N_21449);
xnor U22679 (N_22679,N_21544,N_21430);
nand U22680 (N_22680,N_21496,N_21902);
xnor U22681 (N_22681,N_21957,N_21483);
xor U22682 (N_22682,N_21996,N_21866);
nor U22683 (N_22683,N_21596,N_21896);
nor U22684 (N_22684,N_21194,N_21909);
xnor U22685 (N_22685,N_21797,N_21303);
and U22686 (N_22686,N_21906,N_21295);
nor U22687 (N_22687,N_21096,N_21483);
nor U22688 (N_22688,N_21702,N_21844);
or U22689 (N_22689,N_21745,N_21352);
or U22690 (N_22690,N_21203,N_21091);
nand U22691 (N_22691,N_21419,N_21056);
nand U22692 (N_22692,N_21734,N_21063);
nand U22693 (N_22693,N_21166,N_21445);
and U22694 (N_22694,N_21549,N_21535);
or U22695 (N_22695,N_21111,N_21364);
nand U22696 (N_22696,N_21239,N_21480);
xor U22697 (N_22697,N_21241,N_21973);
or U22698 (N_22698,N_21144,N_21920);
or U22699 (N_22699,N_21740,N_21752);
nor U22700 (N_22700,N_21032,N_21849);
nand U22701 (N_22701,N_21261,N_21928);
and U22702 (N_22702,N_21301,N_21962);
nor U22703 (N_22703,N_21542,N_21970);
xor U22704 (N_22704,N_21638,N_21831);
and U22705 (N_22705,N_21199,N_21862);
xor U22706 (N_22706,N_21210,N_21120);
nor U22707 (N_22707,N_21228,N_21745);
xnor U22708 (N_22708,N_21194,N_21972);
and U22709 (N_22709,N_21348,N_21015);
nand U22710 (N_22710,N_21040,N_21492);
nand U22711 (N_22711,N_21614,N_21097);
nor U22712 (N_22712,N_21846,N_21833);
nand U22713 (N_22713,N_21859,N_21552);
and U22714 (N_22714,N_21825,N_21986);
nor U22715 (N_22715,N_21404,N_21513);
and U22716 (N_22716,N_21589,N_21800);
nand U22717 (N_22717,N_21070,N_21507);
xor U22718 (N_22718,N_21569,N_21801);
nor U22719 (N_22719,N_21401,N_21515);
nand U22720 (N_22720,N_21105,N_21893);
nand U22721 (N_22721,N_21876,N_21140);
or U22722 (N_22722,N_21325,N_21576);
or U22723 (N_22723,N_21872,N_21963);
and U22724 (N_22724,N_21345,N_21654);
nand U22725 (N_22725,N_21203,N_21821);
or U22726 (N_22726,N_21077,N_21344);
nor U22727 (N_22727,N_21867,N_21474);
nor U22728 (N_22728,N_21632,N_21210);
nor U22729 (N_22729,N_21526,N_21283);
and U22730 (N_22730,N_21717,N_21073);
or U22731 (N_22731,N_21060,N_21844);
and U22732 (N_22732,N_21130,N_21650);
nand U22733 (N_22733,N_21331,N_21736);
nor U22734 (N_22734,N_21503,N_21167);
xnor U22735 (N_22735,N_21814,N_21303);
xnor U22736 (N_22736,N_21231,N_21755);
and U22737 (N_22737,N_21502,N_21068);
nor U22738 (N_22738,N_21843,N_21707);
nor U22739 (N_22739,N_21844,N_21189);
xnor U22740 (N_22740,N_21401,N_21868);
and U22741 (N_22741,N_21216,N_21011);
and U22742 (N_22742,N_21405,N_21475);
xnor U22743 (N_22743,N_21624,N_21935);
or U22744 (N_22744,N_21452,N_21064);
xnor U22745 (N_22745,N_21231,N_21827);
nor U22746 (N_22746,N_21658,N_21751);
nor U22747 (N_22747,N_21740,N_21014);
and U22748 (N_22748,N_21700,N_21971);
xor U22749 (N_22749,N_21894,N_21454);
xor U22750 (N_22750,N_21872,N_21501);
xor U22751 (N_22751,N_21737,N_21672);
or U22752 (N_22752,N_21988,N_21207);
xnor U22753 (N_22753,N_21066,N_21348);
or U22754 (N_22754,N_21553,N_21538);
and U22755 (N_22755,N_21775,N_21413);
nand U22756 (N_22756,N_21438,N_21422);
or U22757 (N_22757,N_21494,N_21828);
or U22758 (N_22758,N_21422,N_21226);
and U22759 (N_22759,N_21840,N_21731);
and U22760 (N_22760,N_21105,N_21486);
or U22761 (N_22761,N_21721,N_21946);
or U22762 (N_22762,N_21831,N_21635);
or U22763 (N_22763,N_21435,N_21085);
nand U22764 (N_22764,N_21463,N_21858);
nand U22765 (N_22765,N_21436,N_21312);
nor U22766 (N_22766,N_21601,N_21964);
and U22767 (N_22767,N_21977,N_21705);
nand U22768 (N_22768,N_21913,N_21306);
xor U22769 (N_22769,N_21252,N_21655);
and U22770 (N_22770,N_21541,N_21559);
or U22771 (N_22771,N_21137,N_21706);
nor U22772 (N_22772,N_21837,N_21252);
and U22773 (N_22773,N_21131,N_21542);
and U22774 (N_22774,N_21490,N_21037);
xor U22775 (N_22775,N_21680,N_21070);
nor U22776 (N_22776,N_21770,N_21348);
or U22777 (N_22777,N_21471,N_21809);
nand U22778 (N_22778,N_21758,N_21751);
nor U22779 (N_22779,N_21901,N_21443);
or U22780 (N_22780,N_21433,N_21749);
or U22781 (N_22781,N_21127,N_21594);
nor U22782 (N_22782,N_21292,N_21444);
nand U22783 (N_22783,N_21026,N_21092);
and U22784 (N_22784,N_21339,N_21771);
xnor U22785 (N_22785,N_21783,N_21677);
xnor U22786 (N_22786,N_21094,N_21573);
xor U22787 (N_22787,N_21530,N_21596);
xor U22788 (N_22788,N_21971,N_21764);
xor U22789 (N_22789,N_21398,N_21064);
or U22790 (N_22790,N_21383,N_21451);
xor U22791 (N_22791,N_21327,N_21179);
or U22792 (N_22792,N_21207,N_21201);
or U22793 (N_22793,N_21068,N_21731);
nor U22794 (N_22794,N_21764,N_21932);
xor U22795 (N_22795,N_21364,N_21324);
or U22796 (N_22796,N_21547,N_21733);
xor U22797 (N_22797,N_21139,N_21437);
or U22798 (N_22798,N_21591,N_21778);
xor U22799 (N_22799,N_21724,N_21199);
and U22800 (N_22800,N_21619,N_21121);
or U22801 (N_22801,N_21515,N_21463);
and U22802 (N_22802,N_21081,N_21239);
nor U22803 (N_22803,N_21210,N_21005);
or U22804 (N_22804,N_21032,N_21845);
or U22805 (N_22805,N_21874,N_21300);
nor U22806 (N_22806,N_21183,N_21736);
xnor U22807 (N_22807,N_21233,N_21373);
nor U22808 (N_22808,N_21952,N_21863);
nand U22809 (N_22809,N_21815,N_21067);
nand U22810 (N_22810,N_21120,N_21422);
nor U22811 (N_22811,N_21932,N_21749);
xor U22812 (N_22812,N_21238,N_21961);
and U22813 (N_22813,N_21000,N_21750);
xnor U22814 (N_22814,N_21107,N_21613);
and U22815 (N_22815,N_21931,N_21638);
nor U22816 (N_22816,N_21730,N_21341);
and U22817 (N_22817,N_21534,N_21687);
and U22818 (N_22818,N_21521,N_21113);
and U22819 (N_22819,N_21961,N_21882);
or U22820 (N_22820,N_21466,N_21649);
xnor U22821 (N_22821,N_21749,N_21622);
nor U22822 (N_22822,N_21076,N_21368);
nand U22823 (N_22823,N_21374,N_21884);
and U22824 (N_22824,N_21375,N_21608);
nor U22825 (N_22825,N_21825,N_21608);
or U22826 (N_22826,N_21496,N_21964);
and U22827 (N_22827,N_21057,N_21761);
nor U22828 (N_22828,N_21043,N_21645);
xnor U22829 (N_22829,N_21224,N_21002);
or U22830 (N_22830,N_21957,N_21959);
xor U22831 (N_22831,N_21363,N_21740);
nor U22832 (N_22832,N_21505,N_21850);
xnor U22833 (N_22833,N_21817,N_21383);
nor U22834 (N_22834,N_21830,N_21365);
nor U22835 (N_22835,N_21724,N_21851);
xor U22836 (N_22836,N_21344,N_21989);
and U22837 (N_22837,N_21617,N_21116);
nand U22838 (N_22838,N_21573,N_21207);
or U22839 (N_22839,N_21174,N_21953);
xnor U22840 (N_22840,N_21845,N_21519);
xor U22841 (N_22841,N_21442,N_21518);
xnor U22842 (N_22842,N_21795,N_21676);
or U22843 (N_22843,N_21630,N_21010);
nand U22844 (N_22844,N_21526,N_21404);
and U22845 (N_22845,N_21177,N_21122);
and U22846 (N_22846,N_21843,N_21427);
and U22847 (N_22847,N_21081,N_21177);
nand U22848 (N_22848,N_21390,N_21522);
and U22849 (N_22849,N_21457,N_21816);
or U22850 (N_22850,N_21838,N_21357);
xnor U22851 (N_22851,N_21456,N_21098);
and U22852 (N_22852,N_21033,N_21975);
nand U22853 (N_22853,N_21259,N_21372);
nor U22854 (N_22854,N_21048,N_21316);
nor U22855 (N_22855,N_21617,N_21997);
nor U22856 (N_22856,N_21500,N_21477);
nor U22857 (N_22857,N_21925,N_21817);
xor U22858 (N_22858,N_21605,N_21135);
nand U22859 (N_22859,N_21520,N_21910);
nor U22860 (N_22860,N_21571,N_21161);
or U22861 (N_22861,N_21518,N_21963);
nor U22862 (N_22862,N_21374,N_21028);
and U22863 (N_22863,N_21018,N_21674);
xor U22864 (N_22864,N_21059,N_21640);
or U22865 (N_22865,N_21171,N_21939);
nand U22866 (N_22866,N_21060,N_21966);
or U22867 (N_22867,N_21518,N_21995);
xnor U22868 (N_22868,N_21519,N_21844);
xor U22869 (N_22869,N_21173,N_21185);
and U22870 (N_22870,N_21138,N_21717);
nand U22871 (N_22871,N_21434,N_21655);
xor U22872 (N_22872,N_21804,N_21937);
xor U22873 (N_22873,N_21865,N_21696);
nor U22874 (N_22874,N_21233,N_21600);
or U22875 (N_22875,N_21292,N_21894);
or U22876 (N_22876,N_21874,N_21837);
nor U22877 (N_22877,N_21802,N_21097);
xor U22878 (N_22878,N_21952,N_21828);
and U22879 (N_22879,N_21486,N_21526);
and U22880 (N_22880,N_21198,N_21575);
or U22881 (N_22881,N_21075,N_21295);
nand U22882 (N_22882,N_21129,N_21928);
xnor U22883 (N_22883,N_21844,N_21421);
or U22884 (N_22884,N_21219,N_21829);
or U22885 (N_22885,N_21722,N_21351);
xnor U22886 (N_22886,N_21387,N_21694);
nor U22887 (N_22887,N_21724,N_21745);
or U22888 (N_22888,N_21987,N_21440);
nand U22889 (N_22889,N_21016,N_21995);
and U22890 (N_22890,N_21407,N_21123);
nor U22891 (N_22891,N_21429,N_21973);
xnor U22892 (N_22892,N_21640,N_21931);
nand U22893 (N_22893,N_21429,N_21642);
nor U22894 (N_22894,N_21530,N_21606);
nor U22895 (N_22895,N_21718,N_21172);
xor U22896 (N_22896,N_21847,N_21800);
and U22897 (N_22897,N_21394,N_21172);
and U22898 (N_22898,N_21897,N_21449);
and U22899 (N_22899,N_21688,N_21754);
and U22900 (N_22900,N_21645,N_21033);
and U22901 (N_22901,N_21075,N_21079);
nor U22902 (N_22902,N_21405,N_21788);
and U22903 (N_22903,N_21385,N_21227);
xor U22904 (N_22904,N_21724,N_21078);
xor U22905 (N_22905,N_21604,N_21405);
and U22906 (N_22906,N_21762,N_21686);
xor U22907 (N_22907,N_21719,N_21298);
and U22908 (N_22908,N_21678,N_21513);
and U22909 (N_22909,N_21581,N_21891);
and U22910 (N_22910,N_21390,N_21676);
xor U22911 (N_22911,N_21625,N_21857);
xnor U22912 (N_22912,N_21355,N_21392);
nor U22913 (N_22913,N_21789,N_21373);
or U22914 (N_22914,N_21672,N_21347);
and U22915 (N_22915,N_21571,N_21378);
and U22916 (N_22916,N_21991,N_21867);
or U22917 (N_22917,N_21773,N_21514);
xnor U22918 (N_22918,N_21082,N_21141);
nor U22919 (N_22919,N_21434,N_21442);
and U22920 (N_22920,N_21532,N_21601);
or U22921 (N_22921,N_21573,N_21308);
nor U22922 (N_22922,N_21718,N_21146);
and U22923 (N_22923,N_21385,N_21991);
and U22924 (N_22924,N_21384,N_21054);
xor U22925 (N_22925,N_21931,N_21922);
nor U22926 (N_22926,N_21096,N_21015);
and U22927 (N_22927,N_21495,N_21024);
or U22928 (N_22928,N_21790,N_21442);
or U22929 (N_22929,N_21368,N_21107);
and U22930 (N_22930,N_21765,N_21155);
nor U22931 (N_22931,N_21064,N_21363);
or U22932 (N_22932,N_21220,N_21416);
or U22933 (N_22933,N_21568,N_21075);
nand U22934 (N_22934,N_21436,N_21752);
nand U22935 (N_22935,N_21571,N_21430);
nor U22936 (N_22936,N_21079,N_21565);
nor U22937 (N_22937,N_21551,N_21501);
and U22938 (N_22938,N_21430,N_21278);
or U22939 (N_22939,N_21728,N_21322);
nor U22940 (N_22940,N_21270,N_21880);
nand U22941 (N_22941,N_21464,N_21634);
and U22942 (N_22942,N_21659,N_21936);
nor U22943 (N_22943,N_21551,N_21042);
nor U22944 (N_22944,N_21564,N_21892);
nor U22945 (N_22945,N_21614,N_21762);
nor U22946 (N_22946,N_21654,N_21957);
nor U22947 (N_22947,N_21962,N_21437);
nand U22948 (N_22948,N_21596,N_21132);
nor U22949 (N_22949,N_21525,N_21297);
and U22950 (N_22950,N_21238,N_21178);
nor U22951 (N_22951,N_21098,N_21751);
xnor U22952 (N_22952,N_21695,N_21824);
nor U22953 (N_22953,N_21555,N_21487);
or U22954 (N_22954,N_21993,N_21373);
and U22955 (N_22955,N_21353,N_21856);
or U22956 (N_22956,N_21042,N_21452);
nor U22957 (N_22957,N_21548,N_21604);
nand U22958 (N_22958,N_21882,N_21613);
nand U22959 (N_22959,N_21756,N_21073);
or U22960 (N_22960,N_21738,N_21907);
nand U22961 (N_22961,N_21576,N_21946);
or U22962 (N_22962,N_21241,N_21436);
nor U22963 (N_22963,N_21040,N_21256);
and U22964 (N_22964,N_21370,N_21622);
or U22965 (N_22965,N_21747,N_21880);
nand U22966 (N_22966,N_21994,N_21270);
or U22967 (N_22967,N_21186,N_21168);
nand U22968 (N_22968,N_21375,N_21369);
or U22969 (N_22969,N_21239,N_21134);
nand U22970 (N_22970,N_21275,N_21124);
nand U22971 (N_22971,N_21779,N_21371);
xor U22972 (N_22972,N_21947,N_21311);
or U22973 (N_22973,N_21227,N_21923);
and U22974 (N_22974,N_21777,N_21208);
nor U22975 (N_22975,N_21659,N_21636);
nand U22976 (N_22976,N_21189,N_21536);
nand U22977 (N_22977,N_21736,N_21968);
and U22978 (N_22978,N_21228,N_21823);
xnor U22979 (N_22979,N_21657,N_21885);
nor U22980 (N_22980,N_21399,N_21413);
nand U22981 (N_22981,N_21911,N_21065);
xor U22982 (N_22982,N_21334,N_21644);
nand U22983 (N_22983,N_21903,N_21815);
or U22984 (N_22984,N_21947,N_21521);
nand U22985 (N_22985,N_21571,N_21099);
xnor U22986 (N_22986,N_21412,N_21126);
or U22987 (N_22987,N_21350,N_21270);
nor U22988 (N_22988,N_21076,N_21777);
nor U22989 (N_22989,N_21211,N_21403);
or U22990 (N_22990,N_21105,N_21991);
and U22991 (N_22991,N_21629,N_21395);
or U22992 (N_22992,N_21805,N_21960);
or U22993 (N_22993,N_21326,N_21878);
nor U22994 (N_22994,N_21969,N_21749);
nand U22995 (N_22995,N_21287,N_21375);
and U22996 (N_22996,N_21538,N_21026);
and U22997 (N_22997,N_21831,N_21174);
and U22998 (N_22998,N_21570,N_21120);
xnor U22999 (N_22999,N_21184,N_21356);
nand U23000 (N_23000,N_22791,N_22547);
xor U23001 (N_23001,N_22830,N_22598);
xor U23002 (N_23002,N_22856,N_22885);
or U23003 (N_23003,N_22499,N_22198);
nand U23004 (N_23004,N_22979,N_22223);
or U23005 (N_23005,N_22265,N_22799);
or U23006 (N_23006,N_22392,N_22860);
and U23007 (N_23007,N_22011,N_22735);
or U23008 (N_23008,N_22784,N_22273);
or U23009 (N_23009,N_22955,N_22588);
or U23010 (N_23010,N_22074,N_22601);
nand U23011 (N_23011,N_22787,N_22161);
and U23012 (N_23012,N_22460,N_22705);
xor U23013 (N_23013,N_22980,N_22441);
nand U23014 (N_23014,N_22016,N_22530);
nor U23015 (N_23015,N_22818,N_22476);
and U23016 (N_23016,N_22987,N_22536);
or U23017 (N_23017,N_22880,N_22896);
and U23018 (N_23018,N_22754,N_22356);
and U23019 (N_23019,N_22910,N_22683);
nor U23020 (N_23020,N_22914,N_22719);
nor U23021 (N_23021,N_22557,N_22444);
or U23022 (N_23022,N_22883,N_22768);
and U23023 (N_23023,N_22626,N_22450);
nand U23024 (N_23024,N_22636,N_22809);
nand U23025 (N_23025,N_22470,N_22751);
nand U23026 (N_23026,N_22371,N_22121);
or U23027 (N_23027,N_22587,N_22898);
or U23028 (N_23028,N_22948,N_22328);
xnor U23029 (N_23029,N_22301,N_22419);
xnor U23030 (N_23030,N_22343,N_22015);
nand U23031 (N_23031,N_22713,N_22580);
or U23032 (N_23032,N_22489,N_22733);
and U23033 (N_23033,N_22072,N_22855);
or U23034 (N_23034,N_22316,N_22999);
or U23035 (N_23035,N_22272,N_22229);
and U23036 (N_23036,N_22826,N_22796);
nor U23037 (N_23037,N_22442,N_22668);
nor U23038 (N_23038,N_22817,N_22188);
nor U23039 (N_23039,N_22413,N_22279);
nor U23040 (N_23040,N_22964,N_22061);
or U23041 (N_23041,N_22632,N_22710);
nor U23042 (N_23042,N_22977,N_22829);
xor U23043 (N_23043,N_22618,N_22305);
xnor U23044 (N_23044,N_22675,N_22421);
and U23045 (N_23045,N_22216,N_22583);
xor U23046 (N_23046,N_22227,N_22113);
or U23047 (N_23047,N_22220,N_22050);
or U23048 (N_23048,N_22084,N_22008);
and U23049 (N_23049,N_22471,N_22953);
or U23050 (N_23050,N_22394,N_22067);
nand U23051 (N_23051,N_22221,N_22317);
nand U23052 (N_23052,N_22628,N_22769);
and U23053 (N_23053,N_22531,N_22092);
nor U23054 (N_23054,N_22767,N_22226);
and U23055 (N_23055,N_22969,N_22892);
or U23056 (N_23056,N_22621,N_22385);
nand U23057 (N_23057,N_22204,N_22065);
and U23058 (N_23058,N_22040,N_22650);
xnor U23059 (N_23059,N_22303,N_22047);
nor U23060 (N_23060,N_22129,N_22157);
nand U23061 (N_23061,N_22319,N_22868);
nand U23062 (N_23062,N_22039,N_22009);
xor U23063 (N_23063,N_22622,N_22036);
or U23064 (N_23064,N_22431,N_22136);
and U23065 (N_23065,N_22562,N_22326);
nand U23066 (N_23066,N_22352,N_22783);
nand U23067 (N_23067,N_22452,N_22174);
and U23068 (N_23068,N_22058,N_22024);
nor U23069 (N_23069,N_22234,N_22678);
xnor U23070 (N_23070,N_22137,N_22607);
nand U23071 (N_23071,N_22921,N_22887);
nor U23072 (N_23072,N_22456,N_22222);
nand U23073 (N_23073,N_22734,N_22781);
nand U23074 (N_23074,N_22417,N_22045);
nor U23075 (N_23075,N_22753,N_22776);
nand U23076 (N_23076,N_22110,N_22746);
or U23077 (N_23077,N_22182,N_22014);
nand U23078 (N_23078,N_22000,N_22582);
and U23079 (N_23079,N_22913,N_22816);
or U23080 (N_23080,N_22379,N_22187);
xnor U23081 (N_23081,N_22595,N_22637);
nand U23082 (N_23082,N_22355,N_22331);
xnor U23083 (N_23083,N_22515,N_22365);
xor U23084 (N_23084,N_22145,N_22037);
nor U23085 (N_23085,N_22771,N_22491);
and U23086 (N_23086,N_22730,N_22199);
nor U23087 (N_23087,N_22917,N_22759);
nand U23088 (N_23088,N_22728,N_22832);
xnor U23089 (N_23089,N_22603,N_22873);
nor U23090 (N_23090,N_22647,N_22612);
and U23091 (N_23091,N_22520,N_22461);
nand U23092 (N_23092,N_22160,N_22928);
nand U23093 (N_23093,N_22423,N_22027);
nand U23094 (N_23094,N_22044,N_22333);
nor U23095 (N_23095,N_22882,N_22790);
xor U23096 (N_23096,N_22646,N_22414);
nand U23097 (N_23097,N_22100,N_22402);
xnor U23098 (N_23098,N_22230,N_22965);
and U23099 (N_23099,N_22060,N_22820);
and U23100 (N_23100,N_22858,N_22154);
nand U23101 (N_23101,N_22398,N_22558);
nor U23102 (N_23102,N_22006,N_22950);
xnor U23103 (N_23103,N_22410,N_22656);
xor U23104 (N_23104,N_22670,N_22958);
nor U23105 (N_23105,N_22158,N_22228);
and U23106 (N_23106,N_22091,N_22908);
and U23107 (N_23107,N_22561,N_22353);
or U23108 (N_23108,N_22082,N_22718);
and U23109 (N_23109,N_22287,N_22259);
nor U23110 (N_23110,N_22897,N_22043);
nand U23111 (N_23111,N_22652,N_22159);
xnor U23112 (N_23112,N_22853,N_22609);
and U23113 (N_23113,N_22116,N_22555);
or U23114 (N_23114,N_22335,N_22173);
xor U23115 (N_23115,N_22737,N_22823);
or U23116 (N_23116,N_22256,N_22378);
xnor U23117 (N_23117,N_22803,N_22695);
nand U23118 (N_23118,N_22981,N_22849);
xor U23119 (N_23119,N_22361,N_22923);
and U23120 (N_23120,N_22134,N_22930);
nor U23121 (N_23121,N_22929,N_22945);
or U23122 (N_23122,N_22155,N_22978);
or U23123 (N_23123,N_22195,N_22590);
or U23124 (N_23124,N_22519,N_22828);
and U23125 (N_23125,N_22164,N_22971);
and U23126 (N_23126,N_22351,N_22942);
and U23127 (N_23127,N_22453,N_22786);
xor U23128 (N_23128,N_22697,N_22801);
nand U23129 (N_23129,N_22821,N_22564);
or U23130 (N_23130,N_22667,N_22684);
or U23131 (N_23131,N_22949,N_22773);
or U23132 (N_23132,N_22020,N_22521);
nor U23133 (N_23133,N_22982,N_22878);
nor U23134 (N_23134,N_22481,N_22834);
nor U23135 (N_23135,N_22542,N_22390);
xor U23136 (N_23136,N_22800,N_22277);
or U23137 (N_23137,N_22545,N_22480);
xnor U23138 (N_23138,N_22947,N_22577);
nand U23139 (N_23139,N_22189,N_22619);
xor U23140 (N_23140,N_22602,N_22132);
or U23141 (N_23141,N_22574,N_22035);
xor U23142 (N_23142,N_22623,N_22032);
xor U23143 (N_23143,N_22117,N_22680);
and U23144 (N_23144,N_22096,N_22935);
nand U23145 (N_23145,N_22957,N_22765);
and U23146 (N_23146,N_22611,N_22151);
nand U23147 (N_23147,N_22862,N_22991);
or U23148 (N_23148,N_22393,N_22313);
xor U23149 (N_23149,N_22167,N_22986);
nand U23150 (N_23150,N_22599,N_22090);
or U23151 (N_23151,N_22320,N_22556);
or U23152 (N_23152,N_22815,N_22696);
or U23153 (N_23153,N_22712,N_22966);
or U23154 (N_23154,N_22563,N_22893);
or U23155 (N_23155,N_22681,N_22387);
nor U23156 (N_23156,N_22870,N_22141);
nor U23157 (N_23157,N_22679,N_22183);
xor U23158 (N_23158,N_22727,N_22989);
nand U23159 (N_23159,N_22150,N_22107);
xor U23160 (N_23160,N_22495,N_22932);
or U23161 (N_23161,N_22926,N_22613);
xnor U23162 (N_23162,N_22049,N_22951);
xnor U23163 (N_23163,N_22645,N_22788);
xor U23164 (N_23164,N_22943,N_22937);
nand U23165 (N_23165,N_22889,N_22886);
nand U23166 (N_23166,N_22498,N_22846);
and U23167 (N_23167,N_22996,N_22692);
nand U23168 (N_23168,N_22997,N_22366);
nor U23169 (N_23169,N_22232,N_22118);
nand U23170 (N_23170,N_22732,N_22505);
and U23171 (N_23171,N_22237,N_22057);
xor U23172 (N_23172,N_22546,N_22290);
xnor U23173 (N_23173,N_22778,N_22254);
nand U23174 (N_23174,N_22248,N_22494);
xnor U23175 (N_23175,N_22907,N_22475);
xnor U23176 (N_23176,N_22706,N_22002);
nand U23177 (N_23177,N_22785,N_22376);
nor U23178 (N_23178,N_22029,N_22124);
nor U23179 (N_23179,N_22252,N_22946);
nor U23180 (N_23180,N_22411,N_22034);
and U23181 (N_23181,N_22446,N_22956);
nor U23182 (N_23182,N_22349,N_22640);
xnor U23183 (N_23183,N_22876,N_22224);
or U23184 (N_23184,N_22813,N_22007);
nand U23185 (N_23185,N_22202,N_22443);
or U23186 (N_23186,N_22852,N_22716);
and U23187 (N_23187,N_22406,N_22916);
nor U23188 (N_23188,N_22630,N_22347);
nand U23189 (N_23189,N_22323,N_22792);
xor U23190 (N_23190,N_22021,N_22837);
xnor U23191 (N_23191,N_22915,N_22496);
and U23192 (N_23192,N_22615,N_22472);
xor U23193 (N_23193,N_22133,N_22066);
xnor U23194 (N_23194,N_22418,N_22642);
nor U23195 (N_23195,N_22258,N_22604);
nand U23196 (N_23196,N_22748,N_22899);
and U23197 (N_23197,N_22725,N_22938);
nor U23198 (N_23198,N_22827,N_22140);
xor U23199 (N_23199,N_22686,N_22435);
and U23200 (N_23200,N_22825,N_22225);
or U23201 (N_23201,N_22983,N_22108);
or U23202 (N_23202,N_22432,N_22631);
nor U23203 (N_23203,N_22685,N_22804);
and U23204 (N_23204,N_22522,N_22927);
or U23205 (N_23205,N_22726,N_22436);
or U23206 (N_23206,N_22972,N_22835);
nor U23207 (N_23207,N_22283,N_22963);
nand U23208 (N_23208,N_22135,N_22608);
nor U23209 (N_23209,N_22597,N_22080);
and U23210 (N_23210,N_22936,N_22616);
nor U23211 (N_23211,N_22163,N_22798);
or U23212 (N_23212,N_22872,N_22478);
xnor U23213 (N_23213,N_22428,N_22993);
nor U23214 (N_23214,N_22038,N_22111);
or U23215 (N_23215,N_22425,N_22445);
nand U23216 (N_23216,N_22644,N_22660);
xnor U23217 (N_23217,N_22750,N_22268);
nor U23218 (N_23218,N_22389,N_22156);
nor U23219 (N_23219,N_22115,N_22180);
nor U23220 (N_23220,N_22664,N_22747);
nand U23221 (N_23221,N_22062,N_22627);
nand U23222 (N_23222,N_22723,N_22346);
or U23223 (N_23223,N_22031,N_22203);
nand U23224 (N_23224,N_22152,N_22700);
and U23225 (N_23225,N_22477,N_22780);
or U23226 (N_23226,N_22633,N_22434);
and U23227 (N_23227,N_22181,N_22854);
or U23228 (N_23228,N_22438,N_22077);
or U23229 (N_23229,N_22171,N_22426);
and U23230 (N_23230,N_22805,N_22219);
xnor U23231 (N_23231,N_22560,N_22168);
nand U23232 (N_23232,N_22247,N_22833);
nand U23233 (N_23233,N_22620,N_22375);
xnor U23234 (N_23234,N_22127,N_22324);
nor U23235 (N_23235,N_22779,N_22462);
nor U23236 (N_23236,N_22302,N_22755);
xor U23237 (N_23237,N_22552,N_22403);
nor U23238 (N_23238,N_22424,N_22304);
and U23239 (N_23239,N_22209,N_22524);
or U23240 (N_23240,N_22708,N_22641);
nand U23241 (N_23241,N_22968,N_22760);
nand U23242 (N_23242,N_22253,N_22401);
or U23243 (N_23243,N_22380,N_22172);
and U23244 (N_23244,N_22698,N_22871);
or U23245 (N_23245,N_22079,N_22336);
xnor U23246 (N_23246,N_22210,N_22756);
nand U23247 (N_23247,N_22177,N_22201);
nand U23248 (N_23248,N_22053,N_22857);
nor U23249 (N_23249,N_22493,N_22842);
xor U23250 (N_23250,N_22448,N_22720);
and U23251 (N_23251,N_22125,N_22538);
nor U23252 (N_23252,N_22890,N_22689);
nor U23253 (N_23253,N_22255,N_22528);
and U23254 (N_23254,N_22322,N_22251);
nor U23255 (N_23255,N_22407,N_22506);
nand U23256 (N_23256,N_22592,N_22539);
nor U23257 (N_23257,N_22575,N_22075);
nand U23258 (N_23258,N_22391,N_22193);
nor U23259 (N_23259,N_22373,N_22381);
nand U23260 (N_23260,N_22397,N_22906);
nand U23261 (N_23261,N_22330,N_22533);
nor U23262 (N_23262,N_22439,N_22138);
xor U23263 (N_23263,N_22440,N_22427);
nor U23264 (N_23264,N_22147,N_22447);
nor U23265 (N_23265,N_22299,N_22501);
xor U23266 (N_23266,N_22018,N_22739);
nand U23267 (N_23267,N_22023,N_22148);
and U23268 (N_23268,N_22659,N_22794);
nand U23269 (N_23269,N_22275,N_22812);
xor U23270 (N_23270,N_22578,N_22239);
or U23271 (N_23271,N_22625,N_22408);
or U23272 (N_23272,N_22934,N_22745);
or U23273 (N_23273,N_22022,N_22042);
nand U23274 (N_23274,N_22128,N_22503);
xor U23275 (N_23275,N_22162,N_22344);
xor U23276 (N_23276,N_22257,N_22264);
nor U23277 (N_23277,N_22758,N_22206);
nand U23278 (N_23278,N_22070,N_22338);
nand U23279 (N_23279,N_22088,N_22666);
nand U23280 (N_23280,N_22648,N_22208);
nand U23281 (N_23281,N_22178,N_22102);
and U23282 (N_23282,N_22722,N_22298);
and U23283 (N_23283,N_22565,N_22076);
and U23284 (N_23284,N_22192,N_22166);
nand U23285 (N_23285,N_22924,N_22775);
nor U23286 (N_23286,N_22274,N_22674);
xnor U23287 (N_23287,N_22383,N_22836);
nand U23288 (N_23288,N_22474,N_22242);
xor U23289 (N_23289,N_22231,N_22342);
xor U23290 (N_23290,N_22877,N_22510);
nor U23291 (N_23291,N_22238,N_22988);
nor U23292 (N_23292,N_22153,N_22581);
and U23293 (N_23293,N_22639,N_22850);
nand U23294 (N_23294,N_22990,N_22551);
and U23295 (N_23295,N_22098,N_22415);
nand U23296 (N_23296,N_22869,N_22296);
xor U23297 (N_23297,N_22586,N_22311);
and U23298 (N_23298,N_22691,N_22055);
or U23299 (N_23299,N_22358,N_22715);
xor U23300 (N_23300,N_22717,N_22511);
nand U23301 (N_23301,N_22245,N_22954);
nand U23302 (N_23302,N_22197,N_22702);
or U23303 (N_23303,N_22537,N_22688);
or U23304 (N_23304,N_22321,N_22281);
and U23305 (N_23305,N_22743,N_22831);
xnor U23306 (N_23306,N_22433,N_22984);
or U23307 (N_23307,N_22120,N_22962);
xnor U23308 (N_23308,N_22593,N_22329);
or U23309 (N_23309,N_22742,N_22454);
and U23310 (N_23310,N_22654,N_22286);
and U23311 (N_23311,N_22518,N_22041);
or U23312 (N_23312,N_22861,N_22992);
xnor U23313 (N_23313,N_22711,N_22341);
or U23314 (N_23314,N_22740,N_22584);
nand U23315 (N_23315,N_22741,N_22490);
or U23316 (N_23316,N_22467,N_22701);
nand U23317 (N_23317,N_22811,N_22396);
nor U23318 (N_23318,N_22059,N_22502);
nor U23319 (N_23319,N_22793,N_22738);
nor U23320 (N_23320,N_22658,N_22875);
nor U23321 (N_23321,N_22762,N_22808);
or U23322 (N_23322,N_22819,N_22900);
xnor U23323 (N_23323,N_22360,N_22430);
nor U23324 (N_23324,N_22634,N_22694);
nand U23325 (N_23325,N_22165,N_22271);
xnor U23326 (N_23326,N_22559,N_22844);
nor U23327 (N_23327,N_22569,N_22516);
or U23328 (N_23328,N_22653,N_22196);
or U23329 (N_23329,N_22013,N_22895);
nand U23330 (N_23330,N_22655,N_22149);
nor U23331 (N_23331,N_22269,N_22464);
xor U23332 (N_23332,N_22030,N_22736);
and U23333 (N_23333,N_22540,N_22961);
or U23334 (N_23334,N_22661,N_22369);
and U23335 (N_23335,N_22184,N_22672);
nor U23336 (N_23336,N_22416,N_22384);
nand U23337 (N_23337,N_22614,N_22922);
and U23338 (N_23338,N_22881,N_22789);
nand U23339 (N_23339,N_22863,N_22544);
nor U23340 (N_23340,N_22840,N_22918);
xnor U23341 (N_23341,N_22437,N_22960);
and U23342 (N_23342,N_22367,N_22714);
xnor U23343 (N_23343,N_22554,N_22814);
nand U23344 (N_23344,N_22568,N_22549);
xnor U23345 (N_23345,N_22761,N_22309);
nand U23346 (N_23346,N_22967,N_22282);
xnor U23347 (N_23347,N_22214,N_22651);
xor U23348 (N_23348,N_22482,N_22099);
nand U23349 (N_23349,N_22212,N_22463);
nand U23350 (N_23350,N_22903,N_22843);
and U23351 (N_23351,N_22112,N_22010);
and U23352 (N_23352,N_22068,N_22244);
and U23353 (N_23353,N_22970,N_22497);
xor U23354 (N_23354,N_22486,N_22797);
or U23355 (N_23355,N_22676,N_22795);
and U23356 (N_23356,N_22284,N_22399);
nor U23357 (N_23357,N_22131,N_22422);
nor U23358 (N_23358,N_22867,N_22465);
nand U23359 (N_23359,N_22851,N_22101);
nor U23360 (N_23360,N_22643,N_22483);
nor U23361 (N_23361,N_22845,N_22859);
and U23362 (N_23362,N_22919,N_22280);
nand U23363 (N_23363,N_22105,N_22624);
or U23364 (N_23364,N_22429,N_22291);
nand U23365 (N_23365,N_22451,N_22205);
or U23366 (N_23366,N_22449,N_22529);
or U23367 (N_23367,N_22327,N_22669);
and U23368 (N_23368,N_22362,N_22570);
xnor U23369 (N_23369,N_22334,N_22276);
xnor U23370 (N_23370,N_22412,N_22931);
or U23371 (N_23371,N_22139,N_22606);
nor U23372 (N_23372,N_22218,N_22468);
or U23373 (N_23373,N_22455,N_22146);
nor U23374 (N_23374,N_22806,N_22508);
and U23375 (N_23375,N_22025,N_22270);
nand U23376 (N_23376,N_22553,N_22142);
nor U23377 (N_23377,N_22169,N_22589);
or U23378 (N_23378,N_22363,N_22995);
xnor U23379 (N_23379,N_22388,N_22534);
and U23380 (N_23380,N_22763,N_22894);
xnor U23381 (N_23381,N_22267,N_22236);
xor U23382 (N_23382,N_22841,N_22026);
nand U23383 (N_23383,N_22704,N_22998);
xor U23384 (N_23384,N_22617,N_22864);
xor U23385 (N_23385,N_22063,N_22939);
nand U23386 (N_23386,N_22318,N_22975);
xnor U23387 (N_23387,N_22097,N_22865);
and U23388 (N_23388,N_22485,N_22909);
nand U23389 (N_23389,N_22033,N_22249);
and U23390 (N_23390,N_22404,N_22512);
or U23391 (N_23391,N_22048,N_22517);
and U23392 (N_23392,N_22777,N_22071);
and U23393 (N_23393,N_22004,N_22364);
or U23394 (N_23394,N_22191,N_22523);
and U23395 (N_23395,N_22782,N_22976);
nand U23396 (N_23396,N_22350,N_22901);
nand U23397 (N_23397,N_22332,N_22017);
nand U23398 (N_23398,N_22687,N_22143);
or U23399 (N_23399,N_22089,N_22119);
nand U23400 (N_23400,N_22677,N_22211);
or U23401 (N_23401,N_22484,N_22473);
and U23402 (N_23402,N_22293,N_22001);
nor U23403 (N_23403,N_22054,N_22368);
nand U23404 (N_23404,N_22207,N_22217);
or U23405 (N_23405,N_22504,N_22822);
or U23406 (N_23406,N_22543,N_22952);
xor U23407 (N_23407,N_22469,N_22752);
and U23408 (N_23408,N_22081,N_22576);
or U23409 (N_23409,N_22847,N_22573);
nor U23410 (N_23410,N_22104,N_22003);
nor U23411 (N_23411,N_22629,N_22395);
and U23412 (N_23412,N_22243,N_22525);
nand U23413 (N_23413,N_22535,N_22514);
and U23414 (N_23414,N_22087,N_22064);
xnor U23415 (N_23415,N_22176,N_22459);
nor U23416 (N_23416,N_22749,N_22420);
and U23417 (N_23417,N_22073,N_22250);
or U23418 (N_23418,N_22095,N_22591);
and U23419 (N_23419,N_22126,N_22170);
nand U23420 (N_23420,N_22370,N_22078);
xnor U23421 (N_23421,N_22310,N_22807);
and U23422 (N_23422,N_22213,N_22764);
xnor U23423 (N_23423,N_22888,N_22409);
and U23424 (N_23424,N_22665,N_22377);
and U23425 (N_23425,N_22262,N_22374);
and U23426 (N_23426,N_22579,N_22028);
xor U23427 (N_23427,N_22810,N_22904);
nor U23428 (N_23428,N_22526,N_22292);
nand U23429 (N_23429,N_22487,N_22925);
xor U23430 (N_23430,N_22838,N_22005);
nand U23431 (N_23431,N_22911,N_22289);
or U23432 (N_23432,N_22920,N_22693);
and U23433 (N_23433,N_22114,N_22266);
or U23434 (N_23434,N_22466,N_22610);
nor U23435 (N_23435,N_22673,N_22571);
nand U23436 (N_23436,N_22566,N_22527);
nor U23437 (N_23437,N_22190,N_22359);
and U23438 (N_23438,N_22594,N_22122);
and U23439 (N_23439,N_22635,N_22848);
or U23440 (N_23440,N_22479,N_22772);
nor U23441 (N_23441,N_22260,N_22532);
nor U23442 (N_23442,N_22357,N_22690);
nor U23443 (N_23443,N_22959,N_22703);
nand U23444 (N_23444,N_22405,N_22974);
nor U23445 (N_23445,N_22509,N_22596);
nor U23446 (N_23446,N_22671,N_22314);
or U23447 (N_23447,N_22235,N_22707);
xor U23448 (N_23448,N_22985,N_22884);
nand U23449 (N_23449,N_22548,N_22550);
and U23450 (N_23450,N_22094,N_22766);
or U23451 (N_23451,N_22649,N_22315);
nand U23452 (N_23452,N_22802,N_22354);
or U23453 (N_23453,N_22106,N_22185);
xor U23454 (N_23454,N_22085,N_22400);
nor U23455 (N_23455,N_22109,N_22339);
and U23456 (N_23456,N_22662,N_22724);
and U23457 (N_23457,N_22051,N_22308);
nor U23458 (N_23458,N_22994,N_22731);
nor U23459 (N_23459,N_22744,N_22312);
nor U23460 (N_23460,N_22839,N_22194);
nand U23461 (N_23461,N_22973,N_22103);
nand U23462 (N_23462,N_22012,N_22500);
xnor U23463 (N_23463,N_22069,N_22307);
nor U23464 (N_23464,N_22306,N_22729);
nand U23465 (N_23465,N_22709,N_22585);
or U23466 (N_23466,N_22572,N_22757);
xnor U23467 (N_23467,N_22175,N_22046);
or U23468 (N_23468,N_22297,N_22288);
and U23469 (N_23469,N_22513,N_22507);
xor U23470 (N_23470,N_22294,N_22261);
xnor U23471 (N_23471,N_22052,N_22144);
and U23472 (N_23472,N_22458,N_22774);
or U23473 (N_23473,N_22682,N_22824);
xnor U23474 (N_23474,N_22278,N_22083);
nor U23475 (N_23475,N_22348,N_22492);
nor U23476 (N_23476,N_22770,N_22941);
nor U23477 (N_23477,N_22891,N_22056);
nand U23478 (N_23478,N_22186,N_22541);
and U23479 (N_23479,N_22019,N_22866);
and U23480 (N_23480,N_22300,N_22699);
nand U23481 (N_23481,N_22325,N_22940);
xor U23482 (N_23482,N_22638,N_22457);
or U23483 (N_23483,N_22130,N_22721);
nor U23484 (N_23484,N_22663,N_22902);
xnor U23485 (N_23485,N_22912,N_22263);
or U23486 (N_23486,N_22933,N_22605);
nor U23487 (N_23487,N_22944,N_22123);
and U23488 (N_23488,N_22600,N_22567);
and U23489 (N_23489,N_22657,N_22086);
xor U23490 (N_23490,N_22874,N_22295);
xor U23491 (N_23491,N_22285,N_22372);
and U23492 (N_23492,N_22240,N_22386);
nand U23493 (N_23493,N_22233,N_22488);
xor U23494 (N_23494,N_22879,N_22337);
nor U23495 (N_23495,N_22093,N_22382);
nor U23496 (N_23496,N_22241,N_22905);
and U23497 (N_23497,N_22200,N_22179);
nor U23498 (N_23498,N_22345,N_22215);
nand U23499 (N_23499,N_22246,N_22340);
nand U23500 (N_23500,N_22076,N_22359);
or U23501 (N_23501,N_22242,N_22826);
or U23502 (N_23502,N_22031,N_22802);
or U23503 (N_23503,N_22339,N_22183);
xor U23504 (N_23504,N_22573,N_22809);
or U23505 (N_23505,N_22956,N_22989);
or U23506 (N_23506,N_22150,N_22011);
nand U23507 (N_23507,N_22306,N_22812);
nor U23508 (N_23508,N_22082,N_22517);
xor U23509 (N_23509,N_22708,N_22841);
and U23510 (N_23510,N_22355,N_22041);
nor U23511 (N_23511,N_22081,N_22903);
nand U23512 (N_23512,N_22537,N_22351);
or U23513 (N_23513,N_22163,N_22242);
nor U23514 (N_23514,N_22775,N_22176);
nor U23515 (N_23515,N_22670,N_22680);
xor U23516 (N_23516,N_22685,N_22555);
and U23517 (N_23517,N_22699,N_22585);
nor U23518 (N_23518,N_22264,N_22671);
xor U23519 (N_23519,N_22743,N_22414);
xnor U23520 (N_23520,N_22403,N_22631);
nand U23521 (N_23521,N_22587,N_22031);
nor U23522 (N_23522,N_22635,N_22817);
and U23523 (N_23523,N_22317,N_22970);
nor U23524 (N_23524,N_22110,N_22629);
or U23525 (N_23525,N_22089,N_22181);
nor U23526 (N_23526,N_22702,N_22644);
nand U23527 (N_23527,N_22034,N_22226);
or U23528 (N_23528,N_22557,N_22842);
nand U23529 (N_23529,N_22057,N_22367);
xnor U23530 (N_23530,N_22650,N_22621);
nor U23531 (N_23531,N_22949,N_22515);
nor U23532 (N_23532,N_22302,N_22634);
nor U23533 (N_23533,N_22184,N_22902);
nand U23534 (N_23534,N_22194,N_22965);
and U23535 (N_23535,N_22723,N_22909);
or U23536 (N_23536,N_22094,N_22791);
nor U23537 (N_23537,N_22075,N_22742);
xor U23538 (N_23538,N_22347,N_22780);
nor U23539 (N_23539,N_22845,N_22420);
nand U23540 (N_23540,N_22658,N_22042);
and U23541 (N_23541,N_22236,N_22145);
nand U23542 (N_23542,N_22400,N_22805);
nand U23543 (N_23543,N_22600,N_22279);
and U23544 (N_23544,N_22406,N_22190);
xor U23545 (N_23545,N_22191,N_22569);
xor U23546 (N_23546,N_22591,N_22516);
or U23547 (N_23547,N_22581,N_22191);
nand U23548 (N_23548,N_22942,N_22431);
nor U23549 (N_23549,N_22975,N_22557);
and U23550 (N_23550,N_22290,N_22146);
nor U23551 (N_23551,N_22530,N_22968);
and U23552 (N_23552,N_22508,N_22062);
or U23553 (N_23553,N_22170,N_22633);
xor U23554 (N_23554,N_22491,N_22875);
nand U23555 (N_23555,N_22308,N_22746);
and U23556 (N_23556,N_22903,N_22218);
nor U23557 (N_23557,N_22122,N_22178);
nor U23558 (N_23558,N_22630,N_22678);
or U23559 (N_23559,N_22432,N_22226);
nand U23560 (N_23560,N_22767,N_22802);
nor U23561 (N_23561,N_22295,N_22817);
nand U23562 (N_23562,N_22273,N_22419);
and U23563 (N_23563,N_22863,N_22369);
and U23564 (N_23564,N_22566,N_22365);
nand U23565 (N_23565,N_22478,N_22381);
and U23566 (N_23566,N_22148,N_22368);
nand U23567 (N_23567,N_22924,N_22539);
or U23568 (N_23568,N_22677,N_22380);
and U23569 (N_23569,N_22970,N_22611);
nor U23570 (N_23570,N_22459,N_22648);
nand U23571 (N_23571,N_22827,N_22046);
xor U23572 (N_23572,N_22840,N_22850);
nor U23573 (N_23573,N_22399,N_22028);
nor U23574 (N_23574,N_22095,N_22784);
nand U23575 (N_23575,N_22563,N_22906);
and U23576 (N_23576,N_22699,N_22709);
nand U23577 (N_23577,N_22481,N_22660);
nor U23578 (N_23578,N_22969,N_22248);
xnor U23579 (N_23579,N_22391,N_22370);
xor U23580 (N_23580,N_22678,N_22347);
nor U23581 (N_23581,N_22322,N_22454);
and U23582 (N_23582,N_22688,N_22625);
or U23583 (N_23583,N_22866,N_22211);
nor U23584 (N_23584,N_22757,N_22005);
and U23585 (N_23585,N_22965,N_22810);
and U23586 (N_23586,N_22225,N_22227);
nor U23587 (N_23587,N_22431,N_22911);
or U23588 (N_23588,N_22391,N_22461);
and U23589 (N_23589,N_22471,N_22869);
and U23590 (N_23590,N_22154,N_22897);
nand U23591 (N_23591,N_22515,N_22523);
nand U23592 (N_23592,N_22093,N_22561);
or U23593 (N_23593,N_22154,N_22839);
xnor U23594 (N_23594,N_22883,N_22763);
nand U23595 (N_23595,N_22987,N_22865);
and U23596 (N_23596,N_22156,N_22696);
xnor U23597 (N_23597,N_22921,N_22244);
xor U23598 (N_23598,N_22797,N_22667);
xnor U23599 (N_23599,N_22649,N_22306);
or U23600 (N_23600,N_22230,N_22873);
or U23601 (N_23601,N_22271,N_22025);
nand U23602 (N_23602,N_22500,N_22139);
and U23603 (N_23603,N_22563,N_22821);
nor U23604 (N_23604,N_22896,N_22625);
nand U23605 (N_23605,N_22545,N_22452);
xnor U23606 (N_23606,N_22812,N_22779);
and U23607 (N_23607,N_22572,N_22833);
nor U23608 (N_23608,N_22104,N_22412);
nand U23609 (N_23609,N_22031,N_22515);
and U23610 (N_23610,N_22952,N_22901);
nor U23611 (N_23611,N_22593,N_22167);
and U23612 (N_23612,N_22283,N_22126);
and U23613 (N_23613,N_22175,N_22555);
xor U23614 (N_23614,N_22267,N_22427);
nor U23615 (N_23615,N_22910,N_22307);
nand U23616 (N_23616,N_22134,N_22211);
nor U23617 (N_23617,N_22899,N_22014);
nand U23618 (N_23618,N_22525,N_22277);
and U23619 (N_23619,N_22077,N_22029);
nand U23620 (N_23620,N_22935,N_22061);
nor U23621 (N_23621,N_22420,N_22537);
or U23622 (N_23622,N_22094,N_22162);
nor U23623 (N_23623,N_22676,N_22029);
nor U23624 (N_23624,N_22176,N_22773);
nor U23625 (N_23625,N_22211,N_22607);
xor U23626 (N_23626,N_22354,N_22601);
nor U23627 (N_23627,N_22546,N_22561);
and U23628 (N_23628,N_22956,N_22339);
or U23629 (N_23629,N_22189,N_22791);
and U23630 (N_23630,N_22716,N_22967);
nor U23631 (N_23631,N_22595,N_22807);
xnor U23632 (N_23632,N_22794,N_22273);
or U23633 (N_23633,N_22384,N_22334);
nand U23634 (N_23634,N_22271,N_22157);
nand U23635 (N_23635,N_22845,N_22322);
nand U23636 (N_23636,N_22602,N_22413);
nand U23637 (N_23637,N_22237,N_22045);
and U23638 (N_23638,N_22716,N_22121);
xnor U23639 (N_23639,N_22156,N_22789);
and U23640 (N_23640,N_22842,N_22325);
nand U23641 (N_23641,N_22128,N_22997);
or U23642 (N_23642,N_22836,N_22616);
and U23643 (N_23643,N_22817,N_22769);
nor U23644 (N_23644,N_22303,N_22832);
nand U23645 (N_23645,N_22330,N_22847);
nor U23646 (N_23646,N_22083,N_22215);
xnor U23647 (N_23647,N_22199,N_22552);
nor U23648 (N_23648,N_22921,N_22073);
nand U23649 (N_23649,N_22360,N_22875);
xor U23650 (N_23650,N_22379,N_22700);
and U23651 (N_23651,N_22532,N_22796);
xnor U23652 (N_23652,N_22286,N_22294);
nor U23653 (N_23653,N_22878,N_22622);
xor U23654 (N_23654,N_22625,N_22603);
xor U23655 (N_23655,N_22312,N_22566);
nand U23656 (N_23656,N_22742,N_22272);
nor U23657 (N_23657,N_22602,N_22187);
or U23658 (N_23658,N_22797,N_22231);
nor U23659 (N_23659,N_22123,N_22986);
and U23660 (N_23660,N_22327,N_22533);
xor U23661 (N_23661,N_22572,N_22698);
nand U23662 (N_23662,N_22472,N_22703);
and U23663 (N_23663,N_22735,N_22847);
or U23664 (N_23664,N_22523,N_22101);
nand U23665 (N_23665,N_22767,N_22691);
nor U23666 (N_23666,N_22964,N_22385);
or U23667 (N_23667,N_22935,N_22111);
or U23668 (N_23668,N_22138,N_22277);
nand U23669 (N_23669,N_22190,N_22421);
nand U23670 (N_23670,N_22574,N_22412);
and U23671 (N_23671,N_22722,N_22874);
or U23672 (N_23672,N_22021,N_22968);
and U23673 (N_23673,N_22281,N_22070);
nand U23674 (N_23674,N_22234,N_22863);
nand U23675 (N_23675,N_22977,N_22592);
xor U23676 (N_23676,N_22475,N_22317);
and U23677 (N_23677,N_22690,N_22347);
or U23678 (N_23678,N_22285,N_22413);
and U23679 (N_23679,N_22422,N_22671);
xnor U23680 (N_23680,N_22457,N_22651);
xor U23681 (N_23681,N_22246,N_22341);
and U23682 (N_23682,N_22240,N_22256);
or U23683 (N_23683,N_22417,N_22367);
or U23684 (N_23684,N_22256,N_22025);
nor U23685 (N_23685,N_22204,N_22200);
nor U23686 (N_23686,N_22314,N_22809);
xor U23687 (N_23687,N_22378,N_22968);
nand U23688 (N_23688,N_22374,N_22605);
xnor U23689 (N_23689,N_22004,N_22078);
xor U23690 (N_23690,N_22063,N_22945);
nor U23691 (N_23691,N_22465,N_22489);
nand U23692 (N_23692,N_22680,N_22828);
or U23693 (N_23693,N_22348,N_22690);
or U23694 (N_23694,N_22249,N_22320);
nand U23695 (N_23695,N_22639,N_22785);
and U23696 (N_23696,N_22743,N_22628);
nor U23697 (N_23697,N_22799,N_22165);
xor U23698 (N_23698,N_22631,N_22814);
and U23699 (N_23699,N_22924,N_22463);
or U23700 (N_23700,N_22837,N_22738);
and U23701 (N_23701,N_22584,N_22913);
or U23702 (N_23702,N_22257,N_22988);
and U23703 (N_23703,N_22014,N_22546);
xor U23704 (N_23704,N_22212,N_22729);
nor U23705 (N_23705,N_22880,N_22804);
nor U23706 (N_23706,N_22795,N_22541);
nor U23707 (N_23707,N_22722,N_22545);
xnor U23708 (N_23708,N_22675,N_22882);
or U23709 (N_23709,N_22278,N_22354);
nand U23710 (N_23710,N_22028,N_22879);
nor U23711 (N_23711,N_22634,N_22757);
or U23712 (N_23712,N_22902,N_22352);
xnor U23713 (N_23713,N_22862,N_22057);
nor U23714 (N_23714,N_22746,N_22770);
and U23715 (N_23715,N_22726,N_22604);
and U23716 (N_23716,N_22110,N_22476);
nor U23717 (N_23717,N_22861,N_22209);
xnor U23718 (N_23718,N_22549,N_22999);
nor U23719 (N_23719,N_22146,N_22610);
xnor U23720 (N_23720,N_22316,N_22435);
nor U23721 (N_23721,N_22138,N_22705);
nor U23722 (N_23722,N_22742,N_22444);
or U23723 (N_23723,N_22948,N_22564);
nor U23724 (N_23724,N_22593,N_22536);
nand U23725 (N_23725,N_22920,N_22412);
nand U23726 (N_23726,N_22032,N_22802);
or U23727 (N_23727,N_22255,N_22023);
and U23728 (N_23728,N_22328,N_22332);
xnor U23729 (N_23729,N_22722,N_22651);
xnor U23730 (N_23730,N_22514,N_22051);
xor U23731 (N_23731,N_22125,N_22333);
nor U23732 (N_23732,N_22064,N_22841);
xor U23733 (N_23733,N_22120,N_22904);
or U23734 (N_23734,N_22613,N_22932);
or U23735 (N_23735,N_22242,N_22930);
nand U23736 (N_23736,N_22523,N_22722);
or U23737 (N_23737,N_22493,N_22453);
xor U23738 (N_23738,N_22850,N_22051);
or U23739 (N_23739,N_22348,N_22419);
or U23740 (N_23740,N_22716,N_22382);
nand U23741 (N_23741,N_22734,N_22621);
or U23742 (N_23742,N_22056,N_22492);
and U23743 (N_23743,N_22757,N_22479);
nor U23744 (N_23744,N_22625,N_22662);
nor U23745 (N_23745,N_22154,N_22264);
nand U23746 (N_23746,N_22233,N_22606);
or U23747 (N_23747,N_22396,N_22333);
or U23748 (N_23748,N_22476,N_22696);
and U23749 (N_23749,N_22798,N_22224);
or U23750 (N_23750,N_22156,N_22203);
xor U23751 (N_23751,N_22670,N_22003);
nor U23752 (N_23752,N_22235,N_22876);
nor U23753 (N_23753,N_22330,N_22041);
nor U23754 (N_23754,N_22465,N_22072);
xor U23755 (N_23755,N_22702,N_22528);
xor U23756 (N_23756,N_22879,N_22553);
and U23757 (N_23757,N_22905,N_22137);
nor U23758 (N_23758,N_22792,N_22780);
nand U23759 (N_23759,N_22642,N_22753);
or U23760 (N_23760,N_22393,N_22791);
or U23761 (N_23761,N_22872,N_22137);
nor U23762 (N_23762,N_22079,N_22466);
or U23763 (N_23763,N_22897,N_22460);
and U23764 (N_23764,N_22683,N_22048);
and U23765 (N_23765,N_22405,N_22257);
and U23766 (N_23766,N_22580,N_22166);
xnor U23767 (N_23767,N_22765,N_22503);
or U23768 (N_23768,N_22253,N_22646);
xnor U23769 (N_23769,N_22109,N_22558);
nand U23770 (N_23770,N_22861,N_22980);
or U23771 (N_23771,N_22608,N_22408);
nand U23772 (N_23772,N_22315,N_22532);
and U23773 (N_23773,N_22182,N_22090);
and U23774 (N_23774,N_22198,N_22482);
or U23775 (N_23775,N_22540,N_22643);
and U23776 (N_23776,N_22047,N_22192);
xor U23777 (N_23777,N_22132,N_22083);
xnor U23778 (N_23778,N_22237,N_22839);
or U23779 (N_23779,N_22860,N_22710);
or U23780 (N_23780,N_22200,N_22578);
and U23781 (N_23781,N_22674,N_22854);
and U23782 (N_23782,N_22835,N_22887);
nor U23783 (N_23783,N_22589,N_22136);
nor U23784 (N_23784,N_22047,N_22210);
and U23785 (N_23785,N_22128,N_22752);
nor U23786 (N_23786,N_22332,N_22661);
nand U23787 (N_23787,N_22511,N_22507);
or U23788 (N_23788,N_22673,N_22625);
nand U23789 (N_23789,N_22362,N_22786);
nor U23790 (N_23790,N_22868,N_22287);
xor U23791 (N_23791,N_22144,N_22352);
nor U23792 (N_23792,N_22076,N_22517);
xor U23793 (N_23793,N_22703,N_22992);
xnor U23794 (N_23794,N_22081,N_22342);
nor U23795 (N_23795,N_22177,N_22373);
xor U23796 (N_23796,N_22809,N_22168);
nand U23797 (N_23797,N_22796,N_22340);
nand U23798 (N_23798,N_22398,N_22270);
or U23799 (N_23799,N_22647,N_22170);
xnor U23800 (N_23800,N_22978,N_22415);
nor U23801 (N_23801,N_22861,N_22773);
nor U23802 (N_23802,N_22908,N_22186);
xnor U23803 (N_23803,N_22478,N_22637);
xnor U23804 (N_23804,N_22644,N_22814);
and U23805 (N_23805,N_22119,N_22553);
nand U23806 (N_23806,N_22147,N_22345);
nor U23807 (N_23807,N_22869,N_22352);
xnor U23808 (N_23808,N_22296,N_22983);
xnor U23809 (N_23809,N_22390,N_22580);
nand U23810 (N_23810,N_22831,N_22196);
nand U23811 (N_23811,N_22223,N_22087);
or U23812 (N_23812,N_22627,N_22455);
and U23813 (N_23813,N_22919,N_22661);
nand U23814 (N_23814,N_22819,N_22374);
xnor U23815 (N_23815,N_22602,N_22225);
and U23816 (N_23816,N_22084,N_22552);
nor U23817 (N_23817,N_22386,N_22460);
xnor U23818 (N_23818,N_22458,N_22771);
or U23819 (N_23819,N_22509,N_22407);
or U23820 (N_23820,N_22824,N_22663);
xnor U23821 (N_23821,N_22743,N_22386);
and U23822 (N_23822,N_22565,N_22742);
and U23823 (N_23823,N_22412,N_22722);
nand U23824 (N_23824,N_22635,N_22210);
or U23825 (N_23825,N_22680,N_22379);
and U23826 (N_23826,N_22217,N_22434);
and U23827 (N_23827,N_22008,N_22072);
nor U23828 (N_23828,N_22137,N_22127);
xnor U23829 (N_23829,N_22289,N_22958);
and U23830 (N_23830,N_22407,N_22210);
nand U23831 (N_23831,N_22458,N_22532);
and U23832 (N_23832,N_22480,N_22849);
xnor U23833 (N_23833,N_22898,N_22501);
nand U23834 (N_23834,N_22316,N_22217);
nand U23835 (N_23835,N_22093,N_22104);
nor U23836 (N_23836,N_22677,N_22503);
xnor U23837 (N_23837,N_22052,N_22584);
or U23838 (N_23838,N_22780,N_22445);
and U23839 (N_23839,N_22884,N_22797);
or U23840 (N_23840,N_22713,N_22031);
or U23841 (N_23841,N_22248,N_22872);
xnor U23842 (N_23842,N_22924,N_22960);
or U23843 (N_23843,N_22166,N_22175);
nor U23844 (N_23844,N_22647,N_22652);
or U23845 (N_23845,N_22582,N_22768);
and U23846 (N_23846,N_22607,N_22531);
nor U23847 (N_23847,N_22536,N_22012);
and U23848 (N_23848,N_22716,N_22168);
xnor U23849 (N_23849,N_22764,N_22879);
nand U23850 (N_23850,N_22625,N_22884);
nor U23851 (N_23851,N_22168,N_22164);
nor U23852 (N_23852,N_22150,N_22667);
xor U23853 (N_23853,N_22775,N_22632);
nor U23854 (N_23854,N_22826,N_22856);
or U23855 (N_23855,N_22222,N_22656);
or U23856 (N_23856,N_22623,N_22662);
or U23857 (N_23857,N_22666,N_22573);
and U23858 (N_23858,N_22123,N_22920);
or U23859 (N_23859,N_22138,N_22163);
nand U23860 (N_23860,N_22553,N_22245);
nand U23861 (N_23861,N_22643,N_22302);
or U23862 (N_23862,N_22735,N_22684);
nor U23863 (N_23863,N_22006,N_22023);
nor U23864 (N_23864,N_22930,N_22660);
nand U23865 (N_23865,N_22458,N_22892);
nor U23866 (N_23866,N_22262,N_22580);
or U23867 (N_23867,N_22510,N_22164);
or U23868 (N_23868,N_22545,N_22640);
nor U23869 (N_23869,N_22847,N_22777);
or U23870 (N_23870,N_22239,N_22084);
xnor U23871 (N_23871,N_22604,N_22716);
xor U23872 (N_23872,N_22993,N_22978);
xor U23873 (N_23873,N_22180,N_22715);
or U23874 (N_23874,N_22252,N_22982);
xnor U23875 (N_23875,N_22126,N_22656);
xnor U23876 (N_23876,N_22702,N_22949);
nor U23877 (N_23877,N_22843,N_22810);
nand U23878 (N_23878,N_22279,N_22820);
and U23879 (N_23879,N_22834,N_22635);
xnor U23880 (N_23880,N_22785,N_22448);
nand U23881 (N_23881,N_22299,N_22265);
nor U23882 (N_23882,N_22589,N_22703);
xor U23883 (N_23883,N_22590,N_22775);
and U23884 (N_23884,N_22481,N_22455);
xnor U23885 (N_23885,N_22414,N_22954);
nand U23886 (N_23886,N_22390,N_22762);
xnor U23887 (N_23887,N_22051,N_22964);
or U23888 (N_23888,N_22500,N_22531);
or U23889 (N_23889,N_22618,N_22569);
nand U23890 (N_23890,N_22129,N_22792);
nand U23891 (N_23891,N_22254,N_22865);
or U23892 (N_23892,N_22809,N_22321);
nor U23893 (N_23893,N_22341,N_22298);
nand U23894 (N_23894,N_22808,N_22265);
and U23895 (N_23895,N_22287,N_22348);
or U23896 (N_23896,N_22610,N_22881);
xor U23897 (N_23897,N_22090,N_22022);
nor U23898 (N_23898,N_22089,N_22924);
or U23899 (N_23899,N_22922,N_22738);
or U23900 (N_23900,N_22718,N_22454);
and U23901 (N_23901,N_22760,N_22848);
nor U23902 (N_23902,N_22516,N_22313);
nand U23903 (N_23903,N_22997,N_22268);
nor U23904 (N_23904,N_22185,N_22465);
and U23905 (N_23905,N_22494,N_22499);
or U23906 (N_23906,N_22417,N_22858);
or U23907 (N_23907,N_22988,N_22106);
nand U23908 (N_23908,N_22632,N_22451);
xnor U23909 (N_23909,N_22647,N_22022);
and U23910 (N_23910,N_22513,N_22368);
and U23911 (N_23911,N_22028,N_22647);
xor U23912 (N_23912,N_22039,N_22088);
nor U23913 (N_23913,N_22406,N_22258);
or U23914 (N_23914,N_22894,N_22509);
nand U23915 (N_23915,N_22451,N_22176);
or U23916 (N_23916,N_22638,N_22460);
or U23917 (N_23917,N_22053,N_22434);
xor U23918 (N_23918,N_22515,N_22342);
xnor U23919 (N_23919,N_22803,N_22683);
or U23920 (N_23920,N_22230,N_22860);
nor U23921 (N_23921,N_22406,N_22221);
and U23922 (N_23922,N_22788,N_22918);
nand U23923 (N_23923,N_22724,N_22781);
nor U23924 (N_23924,N_22209,N_22309);
nor U23925 (N_23925,N_22409,N_22180);
nor U23926 (N_23926,N_22295,N_22209);
or U23927 (N_23927,N_22502,N_22404);
xor U23928 (N_23928,N_22031,N_22273);
and U23929 (N_23929,N_22703,N_22431);
nand U23930 (N_23930,N_22296,N_22679);
xnor U23931 (N_23931,N_22184,N_22086);
nand U23932 (N_23932,N_22601,N_22554);
xnor U23933 (N_23933,N_22763,N_22450);
nor U23934 (N_23934,N_22282,N_22235);
or U23935 (N_23935,N_22670,N_22739);
xor U23936 (N_23936,N_22400,N_22079);
and U23937 (N_23937,N_22897,N_22078);
xor U23938 (N_23938,N_22603,N_22883);
or U23939 (N_23939,N_22101,N_22635);
xor U23940 (N_23940,N_22570,N_22633);
nor U23941 (N_23941,N_22145,N_22454);
and U23942 (N_23942,N_22530,N_22049);
nor U23943 (N_23943,N_22003,N_22353);
xnor U23944 (N_23944,N_22600,N_22728);
nor U23945 (N_23945,N_22648,N_22499);
nor U23946 (N_23946,N_22639,N_22130);
nor U23947 (N_23947,N_22526,N_22153);
and U23948 (N_23948,N_22870,N_22749);
nand U23949 (N_23949,N_22142,N_22590);
xor U23950 (N_23950,N_22308,N_22320);
and U23951 (N_23951,N_22797,N_22134);
xnor U23952 (N_23952,N_22548,N_22817);
nor U23953 (N_23953,N_22608,N_22896);
or U23954 (N_23954,N_22412,N_22817);
nor U23955 (N_23955,N_22918,N_22461);
nor U23956 (N_23956,N_22330,N_22606);
xor U23957 (N_23957,N_22902,N_22618);
nand U23958 (N_23958,N_22165,N_22973);
nor U23959 (N_23959,N_22966,N_22326);
or U23960 (N_23960,N_22318,N_22408);
xnor U23961 (N_23961,N_22269,N_22180);
nand U23962 (N_23962,N_22935,N_22176);
nand U23963 (N_23963,N_22582,N_22833);
nand U23964 (N_23964,N_22674,N_22925);
xor U23965 (N_23965,N_22743,N_22108);
nand U23966 (N_23966,N_22592,N_22295);
nand U23967 (N_23967,N_22994,N_22005);
xnor U23968 (N_23968,N_22508,N_22447);
nor U23969 (N_23969,N_22943,N_22640);
nand U23970 (N_23970,N_22911,N_22595);
nor U23971 (N_23971,N_22939,N_22205);
xor U23972 (N_23972,N_22322,N_22616);
and U23973 (N_23973,N_22219,N_22472);
or U23974 (N_23974,N_22007,N_22514);
and U23975 (N_23975,N_22635,N_22993);
or U23976 (N_23976,N_22974,N_22482);
or U23977 (N_23977,N_22145,N_22541);
nor U23978 (N_23978,N_22298,N_22022);
nor U23979 (N_23979,N_22466,N_22838);
nand U23980 (N_23980,N_22115,N_22763);
or U23981 (N_23981,N_22858,N_22555);
or U23982 (N_23982,N_22014,N_22590);
xnor U23983 (N_23983,N_22922,N_22694);
nor U23984 (N_23984,N_22166,N_22261);
or U23985 (N_23985,N_22233,N_22726);
or U23986 (N_23986,N_22248,N_22930);
and U23987 (N_23987,N_22058,N_22130);
nand U23988 (N_23988,N_22110,N_22217);
xnor U23989 (N_23989,N_22703,N_22746);
xor U23990 (N_23990,N_22518,N_22947);
or U23991 (N_23991,N_22443,N_22538);
nand U23992 (N_23992,N_22016,N_22311);
nor U23993 (N_23993,N_22995,N_22670);
nor U23994 (N_23994,N_22311,N_22724);
nand U23995 (N_23995,N_22370,N_22209);
or U23996 (N_23996,N_22932,N_22649);
xnor U23997 (N_23997,N_22542,N_22177);
xor U23998 (N_23998,N_22523,N_22775);
nand U23999 (N_23999,N_22374,N_22290);
nor U24000 (N_24000,N_23093,N_23267);
xnor U24001 (N_24001,N_23935,N_23137);
xnor U24002 (N_24002,N_23508,N_23556);
nand U24003 (N_24003,N_23627,N_23078);
nand U24004 (N_24004,N_23184,N_23472);
xor U24005 (N_24005,N_23357,N_23776);
and U24006 (N_24006,N_23804,N_23528);
xor U24007 (N_24007,N_23883,N_23660);
or U24008 (N_24008,N_23655,N_23286);
and U24009 (N_24009,N_23852,N_23542);
and U24010 (N_24010,N_23320,N_23530);
and U24011 (N_24011,N_23182,N_23207);
nand U24012 (N_24012,N_23754,N_23964);
and U24013 (N_24013,N_23767,N_23661);
and U24014 (N_24014,N_23584,N_23930);
xor U24015 (N_24015,N_23006,N_23509);
xor U24016 (N_24016,N_23225,N_23511);
nand U24017 (N_24017,N_23107,N_23733);
xor U24018 (N_24018,N_23665,N_23546);
and U24019 (N_24019,N_23725,N_23663);
nor U24020 (N_24020,N_23963,N_23626);
and U24021 (N_24021,N_23987,N_23489);
nor U24022 (N_24022,N_23213,N_23903);
and U24023 (N_24023,N_23868,N_23143);
nand U24024 (N_24024,N_23798,N_23040);
or U24025 (N_24025,N_23527,N_23075);
nor U24026 (N_24026,N_23965,N_23693);
nand U24027 (N_24027,N_23447,N_23988);
xnor U24028 (N_24028,N_23768,N_23594);
nor U24029 (N_24029,N_23432,N_23023);
and U24030 (N_24030,N_23314,N_23881);
xnor U24031 (N_24031,N_23013,N_23215);
nor U24032 (N_24032,N_23344,N_23893);
and U24033 (N_24033,N_23356,N_23406);
xor U24034 (N_24034,N_23774,N_23354);
nand U24035 (N_24035,N_23108,N_23667);
nor U24036 (N_24036,N_23050,N_23424);
nor U24037 (N_24037,N_23278,N_23195);
xor U24038 (N_24038,N_23756,N_23970);
or U24039 (N_24039,N_23832,N_23150);
nor U24040 (N_24040,N_23192,N_23346);
and U24041 (N_24041,N_23545,N_23156);
or U24042 (N_24042,N_23334,N_23824);
xor U24043 (N_24043,N_23117,N_23308);
xor U24044 (N_24044,N_23291,N_23414);
nor U24045 (N_24045,N_23098,N_23088);
nand U24046 (N_24046,N_23484,N_23752);
nand U24047 (N_24047,N_23715,N_23951);
xnor U24048 (N_24048,N_23747,N_23980);
nand U24049 (N_24049,N_23766,N_23731);
xnor U24050 (N_24050,N_23142,N_23807);
and U24051 (N_24051,N_23407,N_23989);
nand U24052 (N_24052,N_23934,N_23140);
nor U24053 (N_24053,N_23697,N_23004);
and U24054 (N_24054,N_23639,N_23158);
or U24055 (N_24055,N_23638,N_23479);
nor U24056 (N_24056,N_23478,N_23986);
xnor U24057 (N_24057,N_23403,N_23872);
nor U24058 (N_24058,N_23822,N_23596);
nand U24059 (N_24059,N_23941,N_23429);
and U24060 (N_24060,N_23246,N_23214);
or U24061 (N_24061,N_23276,N_23735);
or U24062 (N_24062,N_23915,N_23421);
nand U24063 (N_24063,N_23871,N_23381);
nor U24064 (N_24064,N_23717,N_23452);
or U24065 (N_24065,N_23387,N_23180);
nand U24066 (N_24066,N_23914,N_23526);
nor U24067 (N_24067,N_23695,N_23514);
and U24068 (N_24068,N_23097,N_23659);
nor U24069 (N_24069,N_23401,N_23703);
and U24070 (N_24070,N_23692,N_23065);
or U24071 (N_24071,N_23255,N_23198);
nand U24072 (N_24072,N_23055,N_23592);
nand U24073 (N_24073,N_23653,N_23073);
nand U24074 (N_24074,N_23814,N_23034);
and U24075 (N_24075,N_23400,N_23386);
or U24076 (N_24076,N_23938,N_23818);
nor U24077 (N_24077,N_23242,N_23196);
nor U24078 (N_24078,N_23590,N_23100);
and U24079 (N_24079,N_23573,N_23337);
and U24080 (N_24080,N_23059,N_23457);
or U24081 (N_24081,N_23516,N_23601);
and U24082 (N_24082,N_23578,N_23032);
or U24083 (N_24083,N_23809,N_23764);
xnor U24084 (N_24084,N_23190,N_23277);
nand U24085 (N_24085,N_23293,N_23686);
nand U24086 (N_24086,N_23624,N_23373);
and U24087 (N_24087,N_23275,N_23550);
and U24088 (N_24088,N_23285,N_23981);
nor U24089 (N_24089,N_23228,N_23569);
xnor U24090 (N_24090,N_23673,N_23537);
nand U24091 (N_24091,N_23269,N_23147);
and U24092 (N_24092,N_23873,N_23253);
nand U24093 (N_24093,N_23751,N_23669);
nand U24094 (N_24094,N_23805,N_23940);
or U24095 (N_24095,N_23786,N_23323);
and U24096 (N_24096,N_23899,N_23666);
xnor U24097 (N_24097,N_23755,N_23904);
and U24098 (N_24098,N_23271,N_23737);
and U24099 (N_24099,N_23002,N_23794);
nor U24100 (N_24100,N_23051,N_23119);
and U24101 (N_24101,N_23290,N_23456);
xnor U24102 (N_24102,N_23652,N_23947);
xnor U24103 (N_24103,N_23770,N_23929);
xnor U24104 (N_24104,N_23124,N_23700);
and U24105 (N_24105,N_23926,N_23463);
nand U24106 (N_24106,N_23576,N_23070);
nand U24107 (N_24107,N_23232,N_23847);
nor U24108 (N_24108,N_23945,N_23816);
xor U24109 (N_24109,N_23466,N_23363);
and U24110 (N_24110,N_23349,N_23920);
nand U24111 (N_24111,N_23483,N_23713);
or U24112 (N_24112,N_23165,N_23561);
xnor U24113 (N_24113,N_23942,N_23061);
xnor U24114 (N_24114,N_23122,N_23038);
nor U24115 (N_24115,N_23110,N_23258);
or U24116 (N_24116,N_23238,N_23604);
nor U24117 (N_24117,N_23315,N_23605);
and U24118 (N_24118,N_23475,N_23729);
nand U24119 (N_24119,N_23758,N_23897);
and U24120 (N_24120,N_23205,N_23895);
xor U24121 (N_24121,N_23145,N_23558);
xnor U24122 (N_24122,N_23112,N_23017);
or U24123 (N_24123,N_23138,N_23919);
or U24124 (N_24124,N_23916,N_23698);
xor U24125 (N_24125,N_23155,N_23706);
nor U24126 (N_24126,N_23887,N_23699);
and U24127 (N_24127,N_23282,N_23829);
nor U24128 (N_24128,N_23338,N_23619);
or U24129 (N_24129,N_23736,N_23091);
or U24130 (N_24130,N_23911,N_23239);
nand U24131 (N_24131,N_23115,N_23801);
and U24132 (N_24132,N_23557,N_23772);
nand U24133 (N_24133,N_23996,N_23146);
nor U24134 (N_24134,N_23379,N_23782);
or U24135 (N_24135,N_23812,N_23311);
xnor U24136 (N_24136,N_23010,N_23992);
and U24137 (N_24137,N_23762,N_23796);
nor U24138 (N_24138,N_23808,N_23902);
or U24139 (N_24139,N_23853,N_23613);
or U24140 (N_24140,N_23876,N_23515);
and U24141 (N_24141,N_23218,N_23200);
and U24142 (N_24142,N_23304,N_23364);
nand U24143 (N_24143,N_23591,N_23330);
nor U24144 (N_24144,N_23481,N_23845);
and U24145 (N_24145,N_23079,N_23614);
xor U24146 (N_24146,N_23744,N_23380);
or U24147 (N_24147,N_23983,N_23679);
or U24148 (N_24148,N_23329,N_23309);
or U24149 (N_24149,N_23047,N_23532);
xnor U24150 (N_24150,N_23046,N_23237);
or U24151 (N_24151,N_23030,N_23132);
and U24152 (N_24152,N_23523,N_23496);
xnor U24153 (N_24153,N_23519,N_23779);
nor U24154 (N_24154,N_23103,N_23450);
and U24155 (N_24155,N_23795,N_23303);
nor U24156 (N_24156,N_23505,N_23102);
nand U24157 (N_24157,N_23843,N_23890);
and U24158 (N_24158,N_23734,N_23946);
xnor U24159 (N_24159,N_23392,N_23628);
nor U24160 (N_24160,N_23943,N_23007);
and U24161 (N_24161,N_23933,N_23748);
or U24162 (N_24162,N_23683,N_23092);
xnor U24163 (N_24163,N_23780,N_23118);
nand U24164 (N_24164,N_23212,N_23813);
nand U24165 (N_24165,N_23281,N_23841);
nand U24166 (N_24166,N_23788,N_23647);
and U24167 (N_24167,N_23470,N_23377);
nor U24168 (N_24168,N_23979,N_23823);
and U24169 (N_24169,N_23325,N_23106);
nor U24170 (N_24170,N_23476,N_23520);
nor U24171 (N_24171,N_23273,N_23567);
and U24172 (N_24172,N_23086,N_23622);
xnor U24173 (N_24173,N_23778,N_23153);
nor U24174 (N_24174,N_23949,N_23008);
or U24175 (N_24175,N_23727,N_23547);
xor U24176 (N_24176,N_23799,N_23444);
xnor U24177 (N_24177,N_23759,N_23825);
xnor U24178 (N_24178,N_23927,N_23080);
or U24179 (N_24179,N_23015,N_23211);
or U24180 (N_24180,N_23244,N_23707);
nand U24181 (N_24181,N_23595,N_23454);
nor U24182 (N_24182,N_23366,N_23410);
nand U24183 (N_24183,N_23838,N_23169);
nor U24184 (N_24184,N_23564,N_23197);
nand U24185 (N_24185,N_23300,N_23861);
and U24186 (N_24186,N_23536,N_23399);
nand U24187 (N_24187,N_23085,N_23966);
nand U24188 (N_24188,N_23453,N_23923);
and U24189 (N_24189,N_23039,N_23127);
nand U24190 (N_24190,N_23284,N_23036);
nand U24191 (N_24191,N_23888,N_23687);
or U24192 (N_24192,N_23264,N_23521);
and U24193 (N_24193,N_23328,N_23602);
xnor U24194 (N_24194,N_23235,N_23283);
nor U24195 (N_24195,N_23869,N_23201);
nand U24196 (N_24196,N_23568,N_23321);
xnor U24197 (N_24197,N_23775,N_23343);
nand U24198 (N_24198,N_23361,N_23402);
nor U24199 (N_24199,N_23125,N_23833);
nor U24200 (N_24200,N_23016,N_23087);
and U24201 (N_24201,N_23741,N_23459);
and U24202 (N_24202,N_23384,N_23723);
nand U24203 (N_24203,N_23451,N_23898);
nor U24204 (N_24204,N_23997,N_23152);
and U24205 (N_24205,N_23765,N_23139);
xnor U24206 (N_24206,N_23307,N_23062);
xnor U24207 (N_24207,N_23784,N_23993);
nand U24208 (N_24208,N_23425,N_23222);
and U24209 (N_24209,N_23850,N_23575);
nand U24210 (N_24210,N_23571,N_23405);
nand U24211 (N_24211,N_23298,N_23045);
or U24212 (N_24212,N_23114,N_23159);
xor U24213 (N_24213,N_23608,N_23135);
xnor U24214 (N_24214,N_23292,N_23531);
xnor U24215 (N_24215,N_23793,N_23969);
or U24216 (N_24216,N_23493,N_23099);
xor U24217 (N_24217,N_23705,N_23418);
and U24218 (N_24218,N_23958,N_23299);
nor U24219 (N_24219,N_23428,N_23412);
and U24220 (N_24220,N_23579,N_23183);
or U24221 (N_24221,N_23581,N_23440);
xor U24222 (N_24222,N_23404,N_23249);
or U24223 (N_24223,N_23461,N_23932);
or U24224 (N_24224,N_23543,N_23477);
xnor U24225 (N_24225,N_23773,N_23552);
xnor U24226 (N_24226,N_23858,N_23005);
xnor U24227 (N_24227,N_23181,N_23306);
xor U24228 (N_24228,N_23830,N_23011);
and U24229 (N_24229,N_23296,N_23014);
nand U24230 (N_24230,N_23629,N_23854);
nand U24231 (N_24231,N_23057,N_23998);
or U24232 (N_24232,N_23339,N_23064);
nor U24233 (N_24233,N_23416,N_23178);
and U24234 (N_24234,N_23396,N_23191);
nand U24235 (N_24235,N_23708,N_23730);
or U24236 (N_24236,N_23123,N_23395);
or U24237 (N_24237,N_23297,N_23719);
xnor U24238 (N_24238,N_23990,N_23690);
nand U24239 (N_24239,N_23113,N_23971);
or U24240 (N_24240,N_23257,N_23921);
or U24241 (N_24241,N_23783,N_23210);
nand U24242 (N_24242,N_23732,N_23513);
and U24243 (N_24243,N_23718,N_23318);
nor U24244 (N_24244,N_23024,N_23577);
nand U24245 (N_24245,N_23021,N_23240);
xor U24246 (N_24246,N_23710,N_23130);
nor U24247 (N_24247,N_23000,N_23574);
and U24248 (N_24248,N_23335,N_23260);
and U24249 (N_24249,N_23445,N_23651);
xor U24250 (N_24250,N_23785,N_23362);
nor U24251 (N_24251,N_23288,N_23041);
nand U24252 (N_24252,N_23160,N_23168);
nor U24253 (N_24253,N_23985,N_23524);
nand U24254 (N_24254,N_23846,N_23711);
or U24255 (N_24255,N_23819,N_23658);
and U24256 (N_24256,N_23676,N_23714);
or U24257 (N_24257,N_23991,N_23185);
nor U24258 (N_24258,N_23555,N_23044);
and U24259 (N_24259,N_23607,N_23900);
and U24260 (N_24260,N_23109,N_23442);
nor U24261 (N_24261,N_23680,N_23372);
and U24262 (N_24262,N_23603,N_23261);
and U24263 (N_24263,N_23488,N_23226);
nand U24264 (N_24264,N_23167,N_23230);
or U24265 (N_24265,N_23559,N_23136);
nor U24266 (N_24266,N_23637,N_23826);
or U24267 (N_24267,N_23355,N_23077);
and U24268 (N_24268,N_23252,N_23394);
nand U24269 (N_24269,N_23797,N_23151);
nor U24270 (N_24270,N_23312,N_23740);
xnor U24271 (N_24271,N_23962,N_23241);
nor U24272 (N_24272,N_23009,N_23166);
nor U24273 (N_24273,N_23533,N_23615);
and U24274 (N_24274,N_23209,N_23874);
xor U24275 (N_24275,N_23095,N_23974);
nor U24276 (N_24276,N_23398,N_23068);
and U24277 (N_24277,N_23501,N_23909);
nand U24278 (N_24278,N_23984,N_23391);
or U24279 (N_24279,N_23671,N_23161);
xor U24280 (N_24280,N_23517,N_23365);
nor U24281 (N_24281,N_23860,N_23769);
and U24282 (N_24282,N_23265,N_23322);
nor U24283 (N_24283,N_23753,N_23074);
nor U24284 (N_24284,N_23562,N_23593);
or U24285 (N_24285,N_23625,N_23623);
nand U24286 (N_24286,N_23722,N_23560);
or U24287 (N_24287,N_23367,N_23674);
xor U24288 (N_24288,N_23173,N_23018);
and U24289 (N_24289,N_23083,N_23957);
nor U24290 (N_24290,N_23487,N_23341);
and U24291 (N_24291,N_23060,N_23891);
and U24292 (N_24292,N_23612,N_23053);
or U24293 (N_24293,N_23208,N_23879);
nor U24294 (N_24294,N_23111,N_23052);
and U24295 (N_24295,N_23928,N_23411);
nor U24296 (N_24296,N_23465,N_23417);
nand U24297 (N_24297,N_23864,N_23423);
xor U24298 (N_24298,N_23179,N_23433);
nand U24299 (N_24299,N_23999,N_23462);
xor U24300 (N_24300,N_23684,N_23875);
xnor U24301 (N_24301,N_23378,N_23128);
nand U24302 (N_24302,N_23154,N_23781);
nand U24303 (N_24303,N_23675,N_23712);
nand U24304 (N_24304,N_23360,N_23548);
xnor U24305 (N_24305,N_23867,N_23069);
nand U24306 (N_24306,N_23022,N_23096);
nand U24307 (N_24307,N_23486,N_23716);
or U24308 (N_24308,N_23172,N_23482);
xor U24309 (N_24309,N_23177,N_23750);
and U24310 (N_24310,N_23954,N_23289);
nand U24311 (N_24311,N_23464,N_23640);
nor U24312 (N_24312,N_23757,N_23174);
and U24313 (N_24313,N_23792,N_23924);
and U24314 (N_24314,N_23617,N_23565);
nand U24315 (N_24315,N_23570,N_23702);
or U24316 (N_24316,N_23701,N_23811);
nor U24317 (N_24317,N_23031,N_23802);
or U24318 (N_24318,N_23742,N_23968);
nand U24319 (N_24319,N_23905,N_23657);
or U24320 (N_24320,N_23071,N_23840);
xnor U24321 (N_24321,N_23485,N_23316);
or U24322 (N_24322,N_23620,N_23089);
xor U24323 (N_24323,N_23352,N_23383);
and U24324 (N_24324,N_23019,N_23886);
xor U24325 (N_24325,N_23681,N_23333);
xnor U24326 (N_24326,N_23650,N_23977);
and U24327 (N_24327,N_23630,N_23609);
nand U24328 (N_24328,N_23437,N_23371);
nor U24329 (N_24329,N_23787,N_23606);
xnor U24330 (N_24330,N_23302,N_23319);
or U24331 (N_24331,N_23141,N_23390);
nor U24332 (N_24332,N_23540,N_23611);
xnor U24333 (N_24333,N_23908,N_23345);
xnor U24334 (N_24334,N_23885,N_23668);
or U24335 (N_24335,N_23430,N_23912);
nor U24336 (N_24336,N_23834,N_23171);
nand U24337 (N_24337,N_23922,N_23842);
and U24338 (N_24338,N_23507,N_23810);
or U24339 (N_24339,N_23549,N_23350);
and U24340 (N_24340,N_23682,N_23917);
or U24341 (N_24341,N_23641,N_23163);
and U24342 (N_24342,N_23295,N_23294);
nor U24343 (N_24343,N_23262,N_23033);
nand U24344 (N_24344,N_23616,N_23896);
xor U24345 (N_24345,N_23491,N_23953);
nand U24346 (N_24346,N_23133,N_23206);
nor U24347 (N_24347,N_23121,N_23189);
nor U24348 (N_24348,N_23862,N_23082);
or U24349 (N_24349,N_23771,N_23572);
nor U24350 (N_24350,N_23104,N_23455);
nand U24351 (N_24351,N_23301,N_23243);
nand U24352 (N_24352,N_23254,N_23251);
and U24353 (N_24353,N_23469,N_23199);
nand U24354 (N_24354,N_23670,N_23855);
nor U24355 (N_24355,N_23721,N_23274);
nor U24356 (N_24356,N_23170,N_23857);
or U24357 (N_24357,N_23101,N_23551);
xor U24358 (N_24358,N_23490,N_23877);
nor U24359 (N_24359,N_23586,N_23203);
nor U24360 (N_24360,N_23599,N_23446);
and U24361 (N_24361,N_23270,N_23026);
xnor U24362 (N_24362,N_23910,N_23848);
nor U24363 (N_24363,N_23506,N_23664);
nor U24364 (N_24364,N_23633,N_23906);
and U24365 (N_24365,N_23157,N_23761);
nand U24366 (N_24366,N_23634,N_23918);
xor U24367 (N_24367,N_23791,N_23054);
or U24368 (N_24368,N_23600,N_23458);
or U24369 (N_24369,N_23336,N_23368);
and U24370 (N_24370,N_23216,N_23956);
xor U24371 (N_24371,N_23844,N_23678);
nor U24372 (N_24372,N_23043,N_23995);
xor U24373 (N_24373,N_23743,N_23076);
or U24374 (N_24374,N_23149,N_23631);
nor U24375 (N_24375,N_23646,N_23831);
xnor U24376 (N_24376,N_23878,N_23534);
nand U24377 (N_24377,N_23925,N_23704);
nor U24378 (N_24378,N_23397,N_23305);
nand U24379 (N_24379,N_23585,N_23512);
and U24380 (N_24380,N_23468,N_23467);
and U24381 (N_24381,N_23313,N_23229);
or U24382 (N_24382,N_23677,N_23806);
xnor U24383 (N_24383,N_23126,N_23495);
or U24384 (N_24384,N_23827,N_23347);
nand U24385 (N_24385,N_23851,N_23648);
xnor U24386 (N_24386,N_23094,N_23374);
nand U24387 (N_24387,N_23116,N_23223);
or U24388 (N_24388,N_23120,N_23863);
or U24389 (N_24389,N_23502,N_23480);
xnor U24390 (N_24390,N_23449,N_23369);
and U24391 (N_24391,N_23866,N_23544);
or U24392 (N_24392,N_23994,N_23382);
or U24393 (N_24393,N_23056,N_23081);
nor U24394 (N_24394,N_23067,N_23975);
nor U24395 (N_24395,N_23849,N_23500);
or U24396 (N_24396,N_23696,N_23803);
xor U24397 (N_24397,N_23760,N_23413);
and U24398 (N_24398,N_23492,N_23131);
and U24399 (N_24399,N_23327,N_23892);
nor U24400 (N_24400,N_23931,N_23164);
nand U24401 (N_24401,N_23777,N_23982);
or U24402 (N_24402,N_23566,N_23800);
nand U24403 (N_24403,N_23589,N_23250);
and U24404 (N_24404,N_23870,N_23415);
xor U24405 (N_24405,N_23385,N_23376);
and U24406 (N_24406,N_23789,N_23066);
nand U24407 (N_24407,N_23880,N_23645);
or U24408 (N_24408,N_23434,N_23029);
and U24409 (N_24409,N_23541,N_23193);
or U24410 (N_24410,N_23259,N_23324);
nor U24411 (N_24411,N_23256,N_23351);
and U24412 (N_24412,N_23538,N_23027);
and U24413 (N_24413,N_23272,N_23090);
or U24414 (N_24414,N_23554,N_23894);
xor U24415 (N_24415,N_23642,N_23865);
and U24416 (N_24416,N_23175,N_23580);
nand U24417 (N_24417,N_23236,N_23221);
xnor U24418 (N_24418,N_23247,N_23419);
nand U24419 (N_24419,N_23370,N_23510);
or U24420 (N_24420,N_23003,N_23287);
or U24421 (N_24421,N_23939,N_23375);
and U24422 (N_24422,N_23204,N_23389);
and U24423 (N_24423,N_23936,N_23331);
or U24424 (N_24424,N_23263,N_23959);
nand U24425 (N_24425,N_23186,N_23728);
xor U24426 (N_24426,N_23907,N_23937);
and U24427 (N_24427,N_23280,N_23738);
and U24428 (N_24428,N_23072,N_23635);
and U24429 (N_24429,N_23884,N_23944);
and U24430 (N_24430,N_23961,N_23162);
and U24431 (N_24431,N_23972,N_23426);
nor U24432 (N_24432,N_23408,N_23420);
and U24433 (N_24433,N_23644,N_23358);
or U24434 (N_24434,N_23474,N_23028);
nand U24435 (N_24435,N_23815,N_23820);
nand U24436 (N_24436,N_23709,N_23950);
or U24437 (N_24437,N_23129,N_23835);
nor U24438 (N_24438,N_23248,N_23340);
and U24439 (N_24439,N_23649,N_23726);
or U24440 (N_24440,N_23105,N_23431);
nor U24441 (N_24441,N_23035,N_23268);
nand U24442 (N_24442,N_23134,N_23393);
nand U24443 (N_24443,N_23234,N_23220);
nand U24444 (N_24444,N_23058,N_23448);
or U24445 (N_24445,N_23348,N_23889);
or U24446 (N_24446,N_23817,N_23438);
or U24447 (N_24447,N_23499,N_23694);
or U24448 (N_24448,N_23525,N_23588);
nor U24449 (N_24449,N_23967,N_23245);
nor U24450 (N_24450,N_23443,N_23498);
xor U24451 (N_24451,N_23749,N_23144);
and U24452 (N_24452,N_23227,N_23224);
xor U24453 (N_24453,N_23084,N_23435);
or U24454 (N_24454,N_23856,N_23471);
or U24455 (N_24455,N_23636,N_23563);
and U24456 (N_24456,N_23194,N_23978);
or U24457 (N_24457,N_23494,N_23233);
or U24458 (N_24458,N_23353,N_23422);
nand U24459 (N_24459,N_23960,N_23739);
nor U24460 (N_24460,N_23643,N_23828);
nor U24461 (N_24461,N_23049,N_23231);
nor U24462 (N_24462,N_23202,N_23187);
or U24463 (N_24463,N_23529,N_23436);
or U24464 (N_24464,N_23317,N_23763);
nor U24465 (N_24465,N_23176,N_23583);
nand U24466 (N_24466,N_23518,N_23662);
and U24467 (N_24467,N_23063,N_23837);
or U24468 (N_24468,N_23689,N_23821);
and U24469 (N_24469,N_23597,N_23553);
and U24470 (N_24470,N_23037,N_23901);
xor U24471 (N_24471,N_23976,N_23497);
nor U24472 (N_24472,N_23882,N_23388);
or U24473 (N_24473,N_23439,N_23952);
xor U24474 (N_24474,N_23656,N_23441);
xor U24475 (N_24475,N_23913,N_23582);
xnor U24476 (N_24476,N_23342,N_23427);
nand U24477 (N_24477,N_23610,N_23839);
xnor U24478 (N_24478,N_23587,N_23460);
nand U24479 (N_24479,N_23621,N_23048);
and U24480 (N_24480,N_23025,N_23503);
or U24481 (N_24481,N_23504,N_23724);
or U24482 (N_24482,N_23522,N_23042);
nand U24483 (N_24483,N_23332,N_23148);
nand U24484 (N_24484,N_23020,N_23217);
xor U24485 (N_24485,N_23219,N_23955);
xnor U24486 (N_24486,N_23266,N_23279);
nand U24487 (N_24487,N_23473,N_23598);
and U24488 (N_24488,N_23310,N_23691);
and U24489 (N_24489,N_23535,N_23188);
nor U24490 (N_24490,N_23672,N_23654);
nand U24491 (N_24491,N_23745,N_23688);
xor U24492 (N_24492,N_23618,N_23012);
and U24493 (N_24493,N_23859,N_23409);
and U24494 (N_24494,N_23720,N_23359);
nor U24495 (N_24495,N_23685,N_23973);
or U24496 (N_24496,N_23790,N_23836);
and U24497 (N_24497,N_23001,N_23746);
or U24498 (N_24498,N_23948,N_23539);
nand U24499 (N_24499,N_23326,N_23632);
nor U24500 (N_24500,N_23241,N_23100);
nand U24501 (N_24501,N_23984,N_23776);
nor U24502 (N_24502,N_23026,N_23598);
nand U24503 (N_24503,N_23960,N_23703);
or U24504 (N_24504,N_23395,N_23646);
nand U24505 (N_24505,N_23025,N_23747);
and U24506 (N_24506,N_23180,N_23136);
xnor U24507 (N_24507,N_23700,N_23856);
and U24508 (N_24508,N_23998,N_23059);
or U24509 (N_24509,N_23226,N_23873);
nor U24510 (N_24510,N_23125,N_23522);
and U24511 (N_24511,N_23652,N_23611);
nor U24512 (N_24512,N_23839,N_23280);
and U24513 (N_24513,N_23794,N_23908);
and U24514 (N_24514,N_23356,N_23682);
or U24515 (N_24515,N_23196,N_23739);
nor U24516 (N_24516,N_23250,N_23591);
nand U24517 (N_24517,N_23868,N_23760);
xor U24518 (N_24518,N_23501,N_23408);
nor U24519 (N_24519,N_23030,N_23597);
xnor U24520 (N_24520,N_23323,N_23870);
nand U24521 (N_24521,N_23245,N_23495);
nand U24522 (N_24522,N_23902,N_23216);
and U24523 (N_24523,N_23207,N_23862);
and U24524 (N_24524,N_23830,N_23260);
or U24525 (N_24525,N_23053,N_23146);
nor U24526 (N_24526,N_23159,N_23985);
or U24527 (N_24527,N_23568,N_23072);
xnor U24528 (N_24528,N_23135,N_23628);
or U24529 (N_24529,N_23809,N_23203);
nor U24530 (N_24530,N_23623,N_23247);
nand U24531 (N_24531,N_23897,N_23987);
nor U24532 (N_24532,N_23798,N_23753);
and U24533 (N_24533,N_23806,N_23917);
nand U24534 (N_24534,N_23159,N_23513);
and U24535 (N_24535,N_23806,N_23629);
nor U24536 (N_24536,N_23586,N_23697);
and U24537 (N_24537,N_23501,N_23379);
xnor U24538 (N_24538,N_23709,N_23919);
nor U24539 (N_24539,N_23002,N_23975);
xnor U24540 (N_24540,N_23374,N_23789);
or U24541 (N_24541,N_23235,N_23515);
or U24542 (N_24542,N_23146,N_23609);
and U24543 (N_24543,N_23109,N_23341);
nand U24544 (N_24544,N_23628,N_23849);
and U24545 (N_24545,N_23326,N_23376);
and U24546 (N_24546,N_23756,N_23128);
xor U24547 (N_24547,N_23933,N_23458);
nor U24548 (N_24548,N_23675,N_23554);
nand U24549 (N_24549,N_23531,N_23870);
nor U24550 (N_24550,N_23919,N_23715);
nand U24551 (N_24551,N_23943,N_23660);
nand U24552 (N_24552,N_23748,N_23828);
and U24553 (N_24553,N_23714,N_23041);
or U24554 (N_24554,N_23661,N_23531);
xor U24555 (N_24555,N_23906,N_23697);
and U24556 (N_24556,N_23742,N_23414);
or U24557 (N_24557,N_23542,N_23072);
xor U24558 (N_24558,N_23825,N_23722);
nand U24559 (N_24559,N_23649,N_23239);
nand U24560 (N_24560,N_23471,N_23862);
or U24561 (N_24561,N_23898,N_23516);
nand U24562 (N_24562,N_23117,N_23063);
xor U24563 (N_24563,N_23170,N_23900);
and U24564 (N_24564,N_23817,N_23146);
xor U24565 (N_24565,N_23477,N_23639);
and U24566 (N_24566,N_23407,N_23357);
or U24567 (N_24567,N_23510,N_23291);
xnor U24568 (N_24568,N_23295,N_23053);
nor U24569 (N_24569,N_23818,N_23655);
and U24570 (N_24570,N_23033,N_23604);
nand U24571 (N_24571,N_23085,N_23826);
nand U24572 (N_24572,N_23202,N_23331);
or U24573 (N_24573,N_23604,N_23045);
nand U24574 (N_24574,N_23098,N_23061);
nand U24575 (N_24575,N_23997,N_23322);
xor U24576 (N_24576,N_23815,N_23929);
or U24577 (N_24577,N_23824,N_23314);
or U24578 (N_24578,N_23461,N_23651);
nor U24579 (N_24579,N_23749,N_23665);
nand U24580 (N_24580,N_23102,N_23201);
and U24581 (N_24581,N_23674,N_23357);
and U24582 (N_24582,N_23380,N_23159);
xor U24583 (N_24583,N_23121,N_23655);
and U24584 (N_24584,N_23093,N_23675);
xor U24585 (N_24585,N_23790,N_23663);
and U24586 (N_24586,N_23625,N_23936);
nand U24587 (N_24587,N_23192,N_23964);
nor U24588 (N_24588,N_23932,N_23049);
or U24589 (N_24589,N_23519,N_23385);
nand U24590 (N_24590,N_23748,N_23094);
nor U24591 (N_24591,N_23855,N_23933);
or U24592 (N_24592,N_23135,N_23488);
nor U24593 (N_24593,N_23768,N_23634);
and U24594 (N_24594,N_23211,N_23066);
nand U24595 (N_24595,N_23565,N_23131);
nand U24596 (N_24596,N_23010,N_23560);
or U24597 (N_24597,N_23966,N_23034);
nand U24598 (N_24598,N_23086,N_23093);
or U24599 (N_24599,N_23182,N_23794);
nand U24600 (N_24600,N_23693,N_23991);
nand U24601 (N_24601,N_23293,N_23983);
or U24602 (N_24602,N_23894,N_23710);
and U24603 (N_24603,N_23058,N_23458);
nor U24604 (N_24604,N_23538,N_23775);
nand U24605 (N_24605,N_23771,N_23076);
nor U24606 (N_24606,N_23259,N_23038);
or U24607 (N_24607,N_23581,N_23404);
nand U24608 (N_24608,N_23943,N_23541);
nand U24609 (N_24609,N_23730,N_23158);
nand U24610 (N_24610,N_23419,N_23873);
xnor U24611 (N_24611,N_23359,N_23853);
xor U24612 (N_24612,N_23378,N_23492);
nor U24613 (N_24613,N_23910,N_23134);
and U24614 (N_24614,N_23901,N_23934);
nand U24615 (N_24615,N_23767,N_23181);
nor U24616 (N_24616,N_23252,N_23558);
nor U24617 (N_24617,N_23748,N_23790);
xor U24618 (N_24618,N_23224,N_23241);
or U24619 (N_24619,N_23825,N_23322);
or U24620 (N_24620,N_23534,N_23095);
and U24621 (N_24621,N_23843,N_23132);
nand U24622 (N_24622,N_23211,N_23987);
nor U24623 (N_24623,N_23282,N_23767);
or U24624 (N_24624,N_23920,N_23701);
and U24625 (N_24625,N_23140,N_23429);
and U24626 (N_24626,N_23367,N_23277);
nor U24627 (N_24627,N_23715,N_23599);
nor U24628 (N_24628,N_23135,N_23978);
xnor U24629 (N_24629,N_23785,N_23738);
xor U24630 (N_24630,N_23167,N_23676);
nor U24631 (N_24631,N_23530,N_23166);
xor U24632 (N_24632,N_23876,N_23610);
and U24633 (N_24633,N_23143,N_23837);
nand U24634 (N_24634,N_23839,N_23563);
xnor U24635 (N_24635,N_23428,N_23664);
nor U24636 (N_24636,N_23105,N_23992);
or U24637 (N_24637,N_23012,N_23930);
nand U24638 (N_24638,N_23077,N_23377);
and U24639 (N_24639,N_23055,N_23198);
or U24640 (N_24640,N_23427,N_23603);
xor U24641 (N_24641,N_23963,N_23095);
nor U24642 (N_24642,N_23913,N_23228);
nand U24643 (N_24643,N_23604,N_23003);
xnor U24644 (N_24644,N_23768,N_23313);
xor U24645 (N_24645,N_23341,N_23046);
and U24646 (N_24646,N_23812,N_23674);
xnor U24647 (N_24647,N_23740,N_23423);
or U24648 (N_24648,N_23815,N_23857);
nor U24649 (N_24649,N_23423,N_23121);
nor U24650 (N_24650,N_23356,N_23885);
xnor U24651 (N_24651,N_23975,N_23183);
nor U24652 (N_24652,N_23829,N_23755);
nor U24653 (N_24653,N_23971,N_23238);
and U24654 (N_24654,N_23347,N_23134);
and U24655 (N_24655,N_23578,N_23410);
and U24656 (N_24656,N_23294,N_23198);
and U24657 (N_24657,N_23900,N_23996);
nand U24658 (N_24658,N_23371,N_23564);
nor U24659 (N_24659,N_23234,N_23542);
and U24660 (N_24660,N_23013,N_23965);
xnor U24661 (N_24661,N_23785,N_23894);
nand U24662 (N_24662,N_23726,N_23220);
xor U24663 (N_24663,N_23066,N_23277);
or U24664 (N_24664,N_23006,N_23895);
nand U24665 (N_24665,N_23476,N_23719);
nor U24666 (N_24666,N_23716,N_23399);
nor U24667 (N_24667,N_23315,N_23703);
or U24668 (N_24668,N_23109,N_23042);
nor U24669 (N_24669,N_23609,N_23590);
and U24670 (N_24670,N_23448,N_23700);
and U24671 (N_24671,N_23777,N_23621);
or U24672 (N_24672,N_23128,N_23436);
or U24673 (N_24673,N_23767,N_23235);
and U24674 (N_24674,N_23394,N_23122);
nor U24675 (N_24675,N_23936,N_23883);
nand U24676 (N_24676,N_23257,N_23755);
and U24677 (N_24677,N_23730,N_23005);
nor U24678 (N_24678,N_23468,N_23261);
and U24679 (N_24679,N_23287,N_23173);
nand U24680 (N_24680,N_23361,N_23439);
xnor U24681 (N_24681,N_23345,N_23497);
xnor U24682 (N_24682,N_23556,N_23510);
nand U24683 (N_24683,N_23635,N_23043);
nand U24684 (N_24684,N_23861,N_23125);
xnor U24685 (N_24685,N_23965,N_23039);
or U24686 (N_24686,N_23230,N_23030);
and U24687 (N_24687,N_23406,N_23980);
nor U24688 (N_24688,N_23147,N_23791);
nand U24689 (N_24689,N_23276,N_23325);
nand U24690 (N_24690,N_23028,N_23166);
nor U24691 (N_24691,N_23893,N_23986);
or U24692 (N_24692,N_23234,N_23847);
nand U24693 (N_24693,N_23747,N_23194);
nor U24694 (N_24694,N_23462,N_23495);
nand U24695 (N_24695,N_23322,N_23601);
nand U24696 (N_24696,N_23479,N_23874);
or U24697 (N_24697,N_23692,N_23115);
and U24698 (N_24698,N_23288,N_23695);
nor U24699 (N_24699,N_23562,N_23446);
or U24700 (N_24700,N_23685,N_23844);
or U24701 (N_24701,N_23051,N_23596);
and U24702 (N_24702,N_23323,N_23528);
or U24703 (N_24703,N_23496,N_23591);
nand U24704 (N_24704,N_23110,N_23068);
nor U24705 (N_24705,N_23540,N_23857);
and U24706 (N_24706,N_23373,N_23822);
nor U24707 (N_24707,N_23747,N_23582);
xnor U24708 (N_24708,N_23775,N_23073);
nor U24709 (N_24709,N_23413,N_23310);
and U24710 (N_24710,N_23990,N_23587);
nor U24711 (N_24711,N_23816,N_23599);
nor U24712 (N_24712,N_23380,N_23770);
nand U24713 (N_24713,N_23703,N_23202);
and U24714 (N_24714,N_23506,N_23836);
xor U24715 (N_24715,N_23239,N_23206);
nor U24716 (N_24716,N_23125,N_23034);
nand U24717 (N_24717,N_23788,N_23981);
nor U24718 (N_24718,N_23008,N_23903);
nand U24719 (N_24719,N_23866,N_23699);
nand U24720 (N_24720,N_23658,N_23641);
and U24721 (N_24721,N_23473,N_23090);
and U24722 (N_24722,N_23373,N_23887);
xor U24723 (N_24723,N_23796,N_23975);
xor U24724 (N_24724,N_23565,N_23404);
nor U24725 (N_24725,N_23653,N_23176);
nand U24726 (N_24726,N_23719,N_23972);
xnor U24727 (N_24727,N_23861,N_23645);
nand U24728 (N_24728,N_23881,N_23976);
nand U24729 (N_24729,N_23917,N_23430);
nor U24730 (N_24730,N_23277,N_23207);
or U24731 (N_24731,N_23900,N_23017);
or U24732 (N_24732,N_23786,N_23886);
and U24733 (N_24733,N_23590,N_23639);
or U24734 (N_24734,N_23991,N_23012);
and U24735 (N_24735,N_23486,N_23663);
or U24736 (N_24736,N_23581,N_23963);
nand U24737 (N_24737,N_23220,N_23167);
nand U24738 (N_24738,N_23105,N_23215);
nand U24739 (N_24739,N_23388,N_23292);
nor U24740 (N_24740,N_23688,N_23149);
or U24741 (N_24741,N_23969,N_23203);
xnor U24742 (N_24742,N_23313,N_23202);
and U24743 (N_24743,N_23395,N_23961);
nor U24744 (N_24744,N_23406,N_23894);
and U24745 (N_24745,N_23154,N_23719);
xnor U24746 (N_24746,N_23155,N_23997);
nor U24747 (N_24747,N_23532,N_23687);
xnor U24748 (N_24748,N_23366,N_23808);
xnor U24749 (N_24749,N_23512,N_23255);
nor U24750 (N_24750,N_23477,N_23584);
and U24751 (N_24751,N_23651,N_23374);
nor U24752 (N_24752,N_23371,N_23350);
xnor U24753 (N_24753,N_23549,N_23610);
nand U24754 (N_24754,N_23419,N_23762);
xor U24755 (N_24755,N_23198,N_23589);
nand U24756 (N_24756,N_23895,N_23421);
and U24757 (N_24757,N_23308,N_23867);
and U24758 (N_24758,N_23540,N_23494);
or U24759 (N_24759,N_23004,N_23208);
nand U24760 (N_24760,N_23346,N_23333);
and U24761 (N_24761,N_23031,N_23966);
nor U24762 (N_24762,N_23994,N_23696);
nor U24763 (N_24763,N_23267,N_23134);
or U24764 (N_24764,N_23230,N_23596);
or U24765 (N_24765,N_23682,N_23085);
or U24766 (N_24766,N_23845,N_23974);
nand U24767 (N_24767,N_23007,N_23849);
nand U24768 (N_24768,N_23797,N_23985);
or U24769 (N_24769,N_23250,N_23802);
or U24770 (N_24770,N_23646,N_23126);
xnor U24771 (N_24771,N_23182,N_23898);
nand U24772 (N_24772,N_23383,N_23258);
nor U24773 (N_24773,N_23660,N_23433);
nand U24774 (N_24774,N_23500,N_23128);
and U24775 (N_24775,N_23887,N_23194);
nor U24776 (N_24776,N_23616,N_23253);
xnor U24777 (N_24777,N_23146,N_23268);
and U24778 (N_24778,N_23808,N_23865);
nor U24779 (N_24779,N_23193,N_23539);
or U24780 (N_24780,N_23027,N_23807);
nor U24781 (N_24781,N_23587,N_23155);
nand U24782 (N_24782,N_23003,N_23787);
xor U24783 (N_24783,N_23301,N_23817);
or U24784 (N_24784,N_23140,N_23210);
nand U24785 (N_24785,N_23994,N_23448);
or U24786 (N_24786,N_23808,N_23199);
or U24787 (N_24787,N_23880,N_23401);
nand U24788 (N_24788,N_23367,N_23508);
and U24789 (N_24789,N_23914,N_23513);
nor U24790 (N_24790,N_23047,N_23193);
nand U24791 (N_24791,N_23593,N_23697);
or U24792 (N_24792,N_23275,N_23658);
nand U24793 (N_24793,N_23495,N_23027);
and U24794 (N_24794,N_23299,N_23748);
nand U24795 (N_24795,N_23583,N_23533);
nor U24796 (N_24796,N_23279,N_23271);
and U24797 (N_24797,N_23082,N_23487);
and U24798 (N_24798,N_23745,N_23491);
and U24799 (N_24799,N_23044,N_23882);
or U24800 (N_24800,N_23827,N_23879);
and U24801 (N_24801,N_23484,N_23917);
nor U24802 (N_24802,N_23469,N_23846);
xor U24803 (N_24803,N_23463,N_23804);
or U24804 (N_24804,N_23768,N_23012);
nor U24805 (N_24805,N_23384,N_23174);
nor U24806 (N_24806,N_23310,N_23563);
or U24807 (N_24807,N_23914,N_23564);
nor U24808 (N_24808,N_23358,N_23305);
nand U24809 (N_24809,N_23342,N_23294);
nor U24810 (N_24810,N_23900,N_23850);
xor U24811 (N_24811,N_23932,N_23751);
and U24812 (N_24812,N_23645,N_23674);
nor U24813 (N_24813,N_23815,N_23948);
nand U24814 (N_24814,N_23969,N_23714);
or U24815 (N_24815,N_23183,N_23068);
or U24816 (N_24816,N_23257,N_23620);
nand U24817 (N_24817,N_23116,N_23900);
or U24818 (N_24818,N_23907,N_23347);
and U24819 (N_24819,N_23577,N_23655);
and U24820 (N_24820,N_23604,N_23035);
and U24821 (N_24821,N_23421,N_23407);
xnor U24822 (N_24822,N_23479,N_23614);
and U24823 (N_24823,N_23131,N_23700);
nor U24824 (N_24824,N_23050,N_23294);
nand U24825 (N_24825,N_23449,N_23558);
nand U24826 (N_24826,N_23666,N_23235);
or U24827 (N_24827,N_23537,N_23846);
xnor U24828 (N_24828,N_23631,N_23971);
or U24829 (N_24829,N_23308,N_23088);
nand U24830 (N_24830,N_23786,N_23377);
xnor U24831 (N_24831,N_23474,N_23872);
nor U24832 (N_24832,N_23085,N_23726);
or U24833 (N_24833,N_23508,N_23925);
xor U24834 (N_24834,N_23485,N_23947);
nand U24835 (N_24835,N_23108,N_23005);
xnor U24836 (N_24836,N_23377,N_23923);
or U24837 (N_24837,N_23033,N_23574);
and U24838 (N_24838,N_23509,N_23023);
or U24839 (N_24839,N_23162,N_23931);
xor U24840 (N_24840,N_23407,N_23717);
and U24841 (N_24841,N_23599,N_23315);
nand U24842 (N_24842,N_23473,N_23299);
and U24843 (N_24843,N_23621,N_23345);
and U24844 (N_24844,N_23103,N_23594);
and U24845 (N_24845,N_23961,N_23825);
and U24846 (N_24846,N_23994,N_23868);
or U24847 (N_24847,N_23839,N_23049);
xor U24848 (N_24848,N_23728,N_23822);
and U24849 (N_24849,N_23555,N_23730);
nand U24850 (N_24850,N_23999,N_23905);
and U24851 (N_24851,N_23607,N_23198);
or U24852 (N_24852,N_23616,N_23731);
nor U24853 (N_24853,N_23762,N_23487);
and U24854 (N_24854,N_23056,N_23576);
nor U24855 (N_24855,N_23935,N_23343);
and U24856 (N_24856,N_23264,N_23181);
nor U24857 (N_24857,N_23763,N_23229);
and U24858 (N_24858,N_23589,N_23149);
or U24859 (N_24859,N_23290,N_23018);
xor U24860 (N_24860,N_23420,N_23993);
xnor U24861 (N_24861,N_23691,N_23721);
or U24862 (N_24862,N_23391,N_23729);
nand U24863 (N_24863,N_23113,N_23458);
xnor U24864 (N_24864,N_23679,N_23006);
nor U24865 (N_24865,N_23323,N_23668);
nand U24866 (N_24866,N_23661,N_23798);
nor U24867 (N_24867,N_23432,N_23935);
nand U24868 (N_24868,N_23612,N_23949);
or U24869 (N_24869,N_23212,N_23306);
or U24870 (N_24870,N_23238,N_23490);
nand U24871 (N_24871,N_23112,N_23204);
nor U24872 (N_24872,N_23167,N_23913);
xor U24873 (N_24873,N_23049,N_23342);
nor U24874 (N_24874,N_23112,N_23536);
or U24875 (N_24875,N_23810,N_23655);
nand U24876 (N_24876,N_23733,N_23277);
nor U24877 (N_24877,N_23669,N_23303);
nand U24878 (N_24878,N_23591,N_23878);
nor U24879 (N_24879,N_23525,N_23797);
or U24880 (N_24880,N_23622,N_23604);
nor U24881 (N_24881,N_23221,N_23109);
or U24882 (N_24882,N_23868,N_23012);
or U24883 (N_24883,N_23547,N_23882);
nor U24884 (N_24884,N_23865,N_23607);
and U24885 (N_24885,N_23911,N_23121);
nand U24886 (N_24886,N_23851,N_23650);
nand U24887 (N_24887,N_23015,N_23224);
nor U24888 (N_24888,N_23719,N_23307);
nor U24889 (N_24889,N_23915,N_23181);
nand U24890 (N_24890,N_23597,N_23642);
or U24891 (N_24891,N_23430,N_23894);
and U24892 (N_24892,N_23278,N_23770);
nor U24893 (N_24893,N_23156,N_23320);
or U24894 (N_24894,N_23175,N_23402);
and U24895 (N_24895,N_23837,N_23845);
nand U24896 (N_24896,N_23481,N_23042);
nor U24897 (N_24897,N_23501,N_23227);
or U24898 (N_24898,N_23692,N_23358);
or U24899 (N_24899,N_23743,N_23376);
and U24900 (N_24900,N_23948,N_23965);
nand U24901 (N_24901,N_23400,N_23417);
xor U24902 (N_24902,N_23786,N_23854);
and U24903 (N_24903,N_23806,N_23937);
xnor U24904 (N_24904,N_23540,N_23853);
xnor U24905 (N_24905,N_23956,N_23026);
nor U24906 (N_24906,N_23668,N_23687);
xor U24907 (N_24907,N_23318,N_23338);
and U24908 (N_24908,N_23168,N_23654);
or U24909 (N_24909,N_23983,N_23193);
and U24910 (N_24910,N_23788,N_23149);
nand U24911 (N_24911,N_23381,N_23356);
xor U24912 (N_24912,N_23978,N_23769);
nand U24913 (N_24913,N_23699,N_23334);
nor U24914 (N_24914,N_23088,N_23612);
nor U24915 (N_24915,N_23124,N_23990);
nand U24916 (N_24916,N_23864,N_23798);
and U24917 (N_24917,N_23531,N_23532);
nand U24918 (N_24918,N_23228,N_23200);
nand U24919 (N_24919,N_23441,N_23031);
nor U24920 (N_24920,N_23938,N_23786);
nor U24921 (N_24921,N_23943,N_23141);
xnor U24922 (N_24922,N_23072,N_23359);
or U24923 (N_24923,N_23169,N_23015);
xnor U24924 (N_24924,N_23729,N_23207);
nor U24925 (N_24925,N_23630,N_23775);
nand U24926 (N_24926,N_23874,N_23007);
xnor U24927 (N_24927,N_23256,N_23314);
or U24928 (N_24928,N_23403,N_23181);
nor U24929 (N_24929,N_23373,N_23398);
xor U24930 (N_24930,N_23335,N_23998);
and U24931 (N_24931,N_23795,N_23005);
nand U24932 (N_24932,N_23099,N_23920);
nand U24933 (N_24933,N_23267,N_23471);
or U24934 (N_24934,N_23063,N_23652);
and U24935 (N_24935,N_23033,N_23473);
or U24936 (N_24936,N_23095,N_23632);
xnor U24937 (N_24937,N_23593,N_23719);
nor U24938 (N_24938,N_23181,N_23473);
and U24939 (N_24939,N_23880,N_23192);
nand U24940 (N_24940,N_23830,N_23570);
and U24941 (N_24941,N_23886,N_23565);
nor U24942 (N_24942,N_23602,N_23361);
or U24943 (N_24943,N_23147,N_23797);
nor U24944 (N_24944,N_23324,N_23197);
xor U24945 (N_24945,N_23262,N_23154);
nand U24946 (N_24946,N_23693,N_23042);
or U24947 (N_24947,N_23086,N_23921);
xor U24948 (N_24948,N_23751,N_23655);
and U24949 (N_24949,N_23203,N_23487);
or U24950 (N_24950,N_23862,N_23545);
nand U24951 (N_24951,N_23213,N_23248);
nor U24952 (N_24952,N_23437,N_23612);
nand U24953 (N_24953,N_23619,N_23057);
nor U24954 (N_24954,N_23494,N_23385);
and U24955 (N_24955,N_23954,N_23945);
or U24956 (N_24956,N_23986,N_23363);
nand U24957 (N_24957,N_23808,N_23941);
and U24958 (N_24958,N_23803,N_23716);
nor U24959 (N_24959,N_23807,N_23087);
nor U24960 (N_24960,N_23601,N_23812);
or U24961 (N_24961,N_23893,N_23020);
and U24962 (N_24962,N_23710,N_23631);
and U24963 (N_24963,N_23063,N_23521);
and U24964 (N_24964,N_23658,N_23485);
and U24965 (N_24965,N_23474,N_23821);
nor U24966 (N_24966,N_23365,N_23661);
nand U24967 (N_24967,N_23699,N_23815);
xor U24968 (N_24968,N_23972,N_23069);
or U24969 (N_24969,N_23043,N_23959);
nand U24970 (N_24970,N_23942,N_23335);
and U24971 (N_24971,N_23011,N_23117);
nor U24972 (N_24972,N_23909,N_23258);
nor U24973 (N_24973,N_23407,N_23820);
and U24974 (N_24974,N_23147,N_23296);
xor U24975 (N_24975,N_23312,N_23289);
and U24976 (N_24976,N_23926,N_23740);
and U24977 (N_24977,N_23414,N_23571);
and U24978 (N_24978,N_23340,N_23686);
and U24979 (N_24979,N_23572,N_23915);
and U24980 (N_24980,N_23009,N_23852);
or U24981 (N_24981,N_23211,N_23069);
nor U24982 (N_24982,N_23818,N_23517);
nand U24983 (N_24983,N_23406,N_23000);
nand U24984 (N_24984,N_23860,N_23549);
xnor U24985 (N_24985,N_23362,N_23177);
nand U24986 (N_24986,N_23446,N_23125);
or U24987 (N_24987,N_23533,N_23211);
nand U24988 (N_24988,N_23418,N_23799);
nand U24989 (N_24989,N_23297,N_23737);
nand U24990 (N_24990,N_23081,N_23901);
xnor U24991 (N_24991,N_23343,N_23641);
and U24992 (N_24992,N_23637,N_23945);
xor U24993 (N_24993,N_23402,N_23025);
nor U24994 (N_24994,N_23040,N_23730);
and U24995 (N_24995,N_23057,N_23858);
and U24996 (N_24996,N_23555,N_23428);
nor U24997 (N_24997,N_23986,N_23740);
or U24998 (N_24998,N_23401,N_23122);
nand U24999 (N_24999,N_23417,N_23424);
nand U25000 (N_25000,N_24219,N_24297);
nand U25001 (N_25001,N_24870,N_24972);
and U25002 (N_25002,N_24812,N_24880);
or U25003 (N_25003,N_24342,N_24910);
nand U25004 (N_25004,N_24209,N_24857);
xnor U25005 (N_25005,N_24763,N_24958);
xor U25006 (N_25006,N_24143,N_24486);
and U25007 (N_25007,N_24771,N_24788);
or U25008 (N_25008,N_24807,N_24122);
nor U25009 (N_25009,N_24742,N_24821);
and U25010 (N_25010,N_24507,N_24890);
nand U25011 (N_25011,N_24450,N_24304);
or U25012 (N_25012,N_24709,N_24469);
or U25013 (N_25013,N_24389,N_24438);
and U25014 (N_25014,N_24093,N_24137);
nor U25015 (N_25015,N_24886,N_24409);
nand U25016 (N_25016,N_24524,N_24430);
nor U25017 (N_25017,N_24236,N_24207);
and U25018 (N_25018,N_24501,N_24801);
or U25019 (N_25019,N_24326,N_24674);
xnor U25020 (N_25020,N_24902,N_24925);
xnor U25021 (N_25021,N_24655,N_24212);
xor U25022 (N_25022,N_24301,N_24615);
nand U25023 (N_25023,N_24035,N_24961);
xnor U25024 (N_25024,N_24878,N_24495);
and U25025 (N_25025,N_24244,N_24052);
xor U25026 (N_25026,N_24999,N_24962);
xnor U25027 (N_25027,N_24444,N_24867);
nand U25028 (N_25028,N_24242,N_24171);
nor U25029 (N_25029,N_24702,N_24249);
nand U25030 (N_25030,N_24017,N_24943);
and U25031 (N_25031,N_24005,N_24467);
nand U25032 (N_25032,N_24422,N_24408);
and U25033 (N_25033,N_24598,N_24809);
nand U25034 (N_25034,N_24105,N_24375);
or U25035 (N_25035,N_24104,N_24038);
or U25036 (N_25036,N_24205,N_24619);
nand U25037 (N_25037,N_24159,N_24838);
nand U25038 (N_25038,N_24359,N_24834);
nand U25039 (N_25039,N_24512,N_24665);
xor U25040 (N_25040,N_24931,N_24976);
and U25041 (N_25041,N_24339,N_24186);
or U25042 (N_25042,N_24117,N_24675);
nor U25043 (N_25043,N_24952,N_24991);
nand U25044 (N_25044,N_24008,N_24449);
nor U25045 (N_25045,N_24168,N_24154);
or U25046 (N_25046,N_24307,N_24669);
and U25047 (N_25047,N_24406,N_24814);
and U25048 (N_25048,N_24403,N_24026);
and U25049 (N_25049,N_24909,N_24893);
nor U25050 (N_25050,N_24975,N_24944);
and U25051 (N_25051,N_24440,N_24077);
or U25052 (N_25052,N_24458,N_24305);
and U25053 (N_25053,N_24491,N_24504);
xnor U25054 (N_25054,N_24855,N_24681);
or U25055 (N_25055,N_24753,N_24348);
or U25056 (N_25056,N_24657,N_24594);
nor U25057 (N_25057,N_24152,N_24290);
nand U25058 (N_25058,N_24576,N_24937);
xnor U25059 (N_25059,N_24575,N_24451);
xnor U25060 (N_25060,N_24213,N_24097);
xor U25061 (N_25061,N_24148,N_24633);
or U25062 (N_25062,N_24025,N_24636);
and U25063 (N_25063,N_24588,N_24695);
nand U25064 (N_25064,N_24523,N_24787);
and U25065 (N_25065,N_24423,N_24885);
nor U25066 (N_25066,N_24531,N_24157);
nor U25067 (N_25067,N_24556,N_24789);
xnor U25068 (N_25068,N_24638,N_24493);
xor U25069 (N_25069,N_24691,N_24019);
xor U25070 (N_25070,N_24622,N_24002);
xnor U25071 (N_25071,N_24955,N_24599);
xnor U25072 (N_25072,N_24484,N_24540);
or U25073 (N_25073,N_24603,N_24377);
nand U25074 (N_25074,N_24967,N_24996);
and U25075 (N_25075,N_24520,N_24061);
or U25076 (N_25076,N_24846,N_24731);
nor U25077 (N_25077,N_24194,N_24490);
and U25078 (N_25078,N_24736,N_24963);
or U25079 (N_25079,N_24472,N_24368);
nand U25080 (N_25080,N_24101,N_24932);
nor U25081 (N_25081,N_24873,N_24965);
or U25082 (N_25082,N_24947,N_24225);
and U25083 (N_25083,N_24732,N_24237);
xor U25084 (N_25084,N_24187,N_24234);
nand U25085 (N_25085,N_24230,N_24116);
or U25086 (N_25086,N_24919,N_24679);
nor U25087 (N_25087,N_24441,N_24687);
or U25088 (N_25088,N_24189,N_24217);
xnor U25089 (N_25089,N_24156,N_24971);
or U25090 (N_25090,N_24069,N_24075);
nor U25091 (N_25091,N_24085,N_24380);
nor U25092 (N_25092,N_24536,N_24772);
and U25093 (N_25093,N_24957,N_24003);
nor U25094 (N_25094,N_24555,N_24593);
and U25095 (N_25095,N_24226,N_24664);
xnor U25096 (N_25096,N_24912,N_24840);
xor U25097 (N_25097,N_24642,N_24605);
nand U25098 (N_25098,N_24037,N_24119);
nand U25099 (N_25099,N_24206,N_24660);
nand U25100 (N_25100,N_24111,N_24724);
nor U25101 (N_25101,N_24843,N_24357);
nor U25102 (N_25102,N_24728,N_24607);
xnor U25103 (N_25103,N_24845,N_24757);
xnor U25104 (N_25104,N_24794,N_24416);
nand U25105 (N_25105,N_24624,N_24903);
xor U25106 (N_25106,N_24269,N_24185);
nand U25107 (N_25107,N_24517,N_24762);
or U25108 (N_25108,N_24898,N_24956);
nor U25109 (N_25109,N_24146,N_24016);
nor U25110 (N_25110,N_24471,N_24969);
or U25111 (N_25111,N_24796,N_24648);
or U25112 (N_25112,N_24365,N_24435);
xor U25113 (N_25113,N_24779,N_24243);
nand U25114 (N_25114,N_24024,N_24783);
and U25115 (N_25115,N_24627,N_24376);
or U25116 (N_25116,N_24927,N_24527);
nor U25117 (N_25117,N_24647,N_24920);
or U25118 (N_25118,N_24267,N_24197);
and U25119 (N_25119,N_24689,N_24806);
and U25120 (N_25120,N_24557,N_24333);
nand U25121 (N_25121,N_24273,N_24711);
or U25122 (N_25122,N_24935,N_24716);
xor U25123 (N_25123,N_24908,N_24871);
or U25124 (N_25124,N_24280,N_24453);
nand U25125 (N_25125,N_24443,N_24699);
nor U25126 (N_25126,N_24247,N_24338);
xor U25127 (N_25127,N_24799,N_24413);
nor U25128 (N_25128,N_24717,N_24892);
and U25129 (N_25129,N_24204,N_24833);
and U25130 (N_25130,N_24046,N_24245);
or U25131 (N_25131,N_24554,N_24150);
or U25132 (N_25132,N_24130,N_24477);
nand U25133 (N_25133,N_24917,N_24573);
and U25134 (N_25134,N_24172,N_24215);
xnor U25135 (N_25135,N_24447,N_24387);
nand U25136 (N_25136,N_24059,N_24337);
xnor U25137 (N_25137,N_24815,N_24850);
nand U25138 (N_25138,N_24361,N_24317);
or U25139 (N_25139,N_24804,N_24545);
nand U25140 (N_25140,N_24620,N_24398);
xnor U25141 (N_25141,N_24921,N_24564);
nand U25142 (N_25142,N_24597,N_24940);
xor U25143 (N_25143,N_24993,N_24670);
xnor U25144 (N_25144,N_24630,N_24228);
nand U25145 (N_25145,N_24210,N_24718);
nor U25146 (N_25146,N_24532,N_24436);
and U25147 (N_25147,N_24916,N_24856);
and U25148 (N_25148,N_24938,N_24064);
nand U25149 (N_25149,N_24175,N_24259);
and U25150 (N_25150,N_24199,N_24045);
nor U25151 (N_25151,N_24417,N_24765);
xnor U25152 (N_25152,N_24211,N_24819);
or U25153 (N_25153,N_24634,N_24579);
nand U25154 (N_25154,N_24822,N_24107);
nand U25155 (N_25155,N_24465,N_24652);
xnor U25156 (N_25156,N_24028,N_24899);
nand U25157 (N_25157,N_24303,N_24754);
nand U25158 (N_25158,N_24776,N_24663);
nand U25159 (N_25159,N_24256,N_24127);
xor U25160 (N_25160,N_24900,N_24138);
nand U25161 (N_25161,N_24509,N_24565);
and U25162 (N_25162,N_24662,N_24513);
and U25163 (N_25163,N_24577,N_24321);
nand U25164 (N_25164,N_24519,N_24004);
nand U25165 (N_25165,N_24705,N_24553);
nand U25166 (N_25166,N_24808,N_24178);
or U25167 (N_25167,N_24281,N_24538);
xor U25168 (N_25168,N_24549,N_24235);
nor U25169 (N_25169,N_24793,N_24781);
or U25170 (N_25170,N_24446,N_24238);
or U25171 (N_25171,N_24404,N_24327);
or U25172 (N_25172,N_24820,N_24515);
xnor U25173 (N_25173,N_24000,N_24087);
nand U25174 (N_25174,N_24322,N_24367);
xnor U25175 (N_25175,N_24637,N_24537);
xor U25176 (N_25176,N_24714,N_24542);
nand U25177 (N_25177,N_24571,N_24852);
nor U25178 (N_25178,N_24986,N_24264);
or U25179 (N_25179,N_24797,N_24525);
or U25180 (N_25180,N_24155,N_24591);
and U25181 (N_25181,N_24853,N_24666);
nand U25182 (N_25182,N_24054,N_24700);
or U25183 (N_25183,N_24109,N_24511);
xor U25184 (N_25184,N_24849,N_24095);
and U25185 (N_25185,N_24907,N_24514);
or U25186 (N_25186,N_24382,N_24391);
xnor U25187 (N_25187,N_24034,N_24680);
nor U25188 (N_25188,N_24192,N_24492);
nor U25189 (N_25189,N_24027,N_24710);
nor U25190 (N_25190,N_24074,N_24534);
and U25191 (N_25191,N_24750,N_24253);
nand U25192 (N_25192,N_24489,N_24419);
and U25193 (N_25193,N_24190,N_24214);
nand U25194 (N_25194,N_24123,N_24865);
and U25195 (N_25195,N_24528,N_24827);
nand U25196 (N_25196,N_24227,N_24713);
nand U25197 (N_25197,N_24078,N_24274);
nor U25198 (N_25198,N_24174,N_24418);
nand U25199 (N_25199,N_24047,N_24924);
xor U25200 (N_25200,N_24191,N_24229);
nor U25201 (N_25201,N_24544,N_24623);
nor U25202 (N_25202,N_24433,N_24690);
and U25203 (N_25203,N_24758,N_24173);
nand U25204 (N_25204,N_24761,N_24183);
nor U25205 (N_25205,N_24319,N_24948);
and U25206 (N_25206,N_24431,N_24402);
and U25207 (N_25207,N_24454,N_24073);
and U25208 (N_25208,N_24769,N_24094);
nor U25209 (N_25209,N_24448,N_24823);
nand U25210 (N_25210,N_24485,N_24659);
nand U25211 (N_25211,N_24697,N_24708);
nand U25212 (N_25212,N_24445,N_24040);
nand U25213 (N_25213,N_24790,N_24086);
nand U25214 (N_25214,N_24306,N_24875);
xor U25215 (N_25215,N_24552,N_24780);
xor U25216 (N_25216,N_24802,N_24158);
nand U25217 (N_25217,N_24121,N_24629);
xor U25218 (N_25218,N_24982,N_24582);
nand U25219 (N_25219,N_24715,N_24463);
xor U25220 (N_25220,N_24058,N_24559);
or U25221 (N_25221,N_24625,N_24455);
and U25222 (N_25222,N_24782,N_24930);
or U25223 (N_25223,N_24500,N_24007);
and U25224 (N_25224,N_24218,N_24600);
xnor U25225 (N_25225,N_24894,N_24847);
or U25226 (N_25226,N_24278,N_24617);
xnor U25227 (N_25227,N_24990,N_24650);
nand U25228 (N_25228,N_24998,N_24378);
xor U25229 (N_25229,N_24096,N_24112);
or U25230 (N_25230,N_24712,N_24727);
and U25231 (N_25231,N_24295,N_24764);
nand U25232 (N_25232,N_24277,N_24195);
nor U25233 (N_25233,N_24639,N_24476);
nor U25234 (N_25234,N_24678,N_24048);
nor U25235 (N_25235,N_24133,N_24103);
and U25236 (N_25236,N_24730,N_24881);
or U25237 (N_25237,N_24261,N_24784);
or U25238 (N_25238,N_24876,N_24496);
nand U25239 (N_25239,N_24198,N_24318);
and U25240 (N_25240,N_24498,N_24241);
xor U25241 (N_25241,N_24795,N_24181);
nand U25242 (N_25242,N_24018,N_24488);
nand U25243 (N_25243,N_24347,N_24602);
or U25244 (N_25244,N_24836,N_24460);
xnor U25245 (N_25245,N_24062,N_24913);
nand U25246 (N_25246,N_24257,N_24631);
and U25247 (N_25247,N_24706,N_24748);
xnor U25248 (N_25248,N_24981,N_24882);
or U25249 (N_25249,N_24977,N_24851);
or U25250 (N_25250,N_24070,N_24254);
or U25251 (N_25251,N_24379,N_24384);
xnor U25252 (N_25252,N_24426,N_24901);
and U25253 (N_25253,N_24221,N_24562);
and U25254 (N_25254,N_24945,N_24401);
nor U25255 (N_25255,N_24124,N_24407);
xor U25256 (N_25256,N_24405,N_24328);
and U25257 (N_25257,N_24934,N_24543);
and U25258 (N_25258,N_24014,N_24421);
nor U25259 (N_25259,N_24785,N_24539);
and U25260 (N_25260,N_24090,N_24381);
or U25261 (N_25261,N_24839,N_24860);
and U25262 (N_25262,N_24151,N_24291);
and U25263 (N_25263,N_24370,N_24928);
nor U25264 (N_25264,N_24824,N_24071);
nand U25265 (N_25265,N_24315,N_24628);
xor U25266 (N_25266,N_24896,N_24114);
and U25267 (N_25267,N_24287,N_24740);
nor U25268 (N_25268,N_24131,N_24915);
xnor U25269 (N_25269,N_24621,N_24248);
xor U25270 (N_25270,N_24583,N_24614);
or U25271 (N_25271,N_24646,N_24997);
nor U25272 (N_25272,N_24468,N_24029);
xnor U25273 (N_25273,N_24558,N_24580);
or U25274 (N_25274,N_24118,N_24153);
nand U25275 (N_25275,N_24080,N_24547);
nand U25276 (N_25276,N_24766,N_24698);
nand U25277 (N_25277,N_24351,N_24701);
xnor U25278 (N_25278,N_24649,N_24271);
or U25279 (N_25279,N_24721,N_24036);
nor U25280 (N_25280,N_24522,N_24092);
nor U25281 (N_25281,N_24009,N_24825);
nand U25282 (N_25282,N_24798,N_24966);
and U25283 (N_25283,N_24129,N_24533);
xnor U25284 (N_25284,N_24661,N_24053);
or U25285 (N_25285,N_24883,N_24428);
nand U25286 (N_25286,N_24632,N_24499);
and U25287 (N_25287,N_24120,N_24336);
or U25288 (N_25288,N_24672,N_24818);
nand U25289 (N_25289,N_24240,N_24176);
or U25290 (N_25290,N_24099,N_24601);
or U25291 (N_25291,N_24412,N_24115);
nor U25292 (N_25292,N_24320,N_24208);
xor U25293 (N_25293,N_24373,N_24560);
nor U25294 (N_25294,N_24222,N_24992);
and U25295 (N_25295,N_24831,N_24682);
xor U25296 (N_25296,N_24858,N_24743);
nor U25297 (N_25297,N_24006,N_24082);
and U25298 (N_25298,N_24561,N_24369);
nand U25299 (N_25299,N_24313,N_24859);
and U25300 (N_25300,N_24610,N_24033);
and U25301 (N_25301,N_24904,N_24911);
nor U25302 (N_25302,N_24106,N_24371);
nor U25303 (N_25303,N_24311,N_24461);
xnor U25304 (N_25304,N_24887,N_24263);
xnor U25305 (N_25305,N_24363,N_24751);
or U25306 (N_25306,N_24031,N_24044);
or U25307 (N_25307,N_24147,N_24266);
nand U25308 (N_25308,N_24478,N_24049);
nand U25309 (N_25309,N_24848,N_24011);
nor U25310 (N_25310,N_24388,N_24964);
and U25311 (N_25311,N_24126,N_24464);
and U25312 (N_25312,N_24693,N_24592);
xor U25313 (N_25313,N_24079,N_24427);
or U25314 (N_25314,N_24884,N_24113);
or U25315 (N_25315,N_24224,N_24300);
xnor U25316 (N_25316,N_24510,N_24144);
xor U25317 (N_25317,N_24250,N_24725);
and U25318 (N_25318,N_24355,N_24747);
nor U25319 (N_25319,N_24656,N_24541);
xor U25320 (N_25320,N_24001,N_24989);
nor U25321 (N_25321,N_24979,N_24868);
and U25322 (N_25322,N_24959,N_24279);
nand U25323 (N_25323,N_24733,N_24994);
nor U25324 (N_25324,N_24020,N_24922);
and U25325 (N_25325,N_24595,N_24995);
or U25326 (N_25326,N_24506,N_24828);
or U25327 (N_25327,N_24844,N_24739);
xor U25328 (N_25328,N_24518,N_24309);
and U25329 (N_25329,N_24390,N_24569);
xor U25330 (N_25330,N_24563,N_24324);
and U25331 (N_25331,N_24149,N_24584);
or U25332 (N_25332,N_24645,N_24010);
or U25333 (N_25333,N_24604,N_24362);
and U25334 (N_25334,N_24720,N_24658);
nor U25335 (N_25335,N_24497,N_24268);
and U25336 (N_25336,N_24810,N_24756);
nor U25337 (N_25337,N_24165,N_24792);
xor U25338 (N_25338,N_24906,N_24284);
and U25339 (N_25339,N_24612,N_24974);
nor U25340 (N_25340,N_24677,N_24043);
xor U25341 (N_25341,N_24574,N_24550);
and U25342 (N_25342,N_24707,N_24673);
xor U25343 (N_25343,N_24233,N_24864);
nor U25344 (N_25344,N_24169,N_24635);
xor U25345 (N_25345,N_24767,N_24626);
and U25346 (N_25346,N_24012,N_24232);
nand U25347 (N_25347,N_24285,N_24414);
nand U25348 (N_25348,N_24360,N_24466);
or U25349 (N_25349,N_24694,N_24644);
nand U25350 (N_25350,N_24826,N_24667);
and U25351 (N_25351,N_24350,N_24968);
and U25352 (N_25352,N_24276,N_24640);
or U25353 (N_25353,N_24572,N_24960);
nor U25354 (N_25354,N_24570,N_24611);
nand U25355 (N_25355,N_24288,N_24744);
and U25356 (N_25356,N_24778,N_24770);
xor U25357 (N_25357,N_24188,N_24918);
nand U25358 (N_25358,N_24773,N_24255);
or U25359 (N_25359,N_24735,N_24722);
nor U25360 (N_25360,N_24429,N_24272);
and U25361 (N_25361,N_24942,N_24067);
and U25362 (N_25362,N_24482,N_24521);
nor U25363 (N_25363,N_24479,N_24946);
or U25364 (N_25364,N_24193,N_24953);
and U25365 (N_25365,N_24973,N_24415);
nand U25366 (N_25366,N_24393,N_24686);
and U25367 (N_25367,N_24729,N_24400);
and U25368 (N_25368,N_24132,N_24895);
and U25369 (N_25369,N_24581,N_24481);
or U25370 (N_25370,N_24142,N_24590);
xor U25371 (N_25371,N_24530,N_24015);
nand U25372 (N_25372,N_24980,N_24805);
nor U25373 (N_25373,N_24223,N_24813);
and U25374 (N_25374,N_24546,N_24032);
or U25375 (N_25375,N_24654,N_24055);
xor U25376 (N_25376,N_24526,N_24888);
xnor U25377 (N_25377,N_24609,N_24889);
nor U25378 (N_25378,N_24329,N_24316);
xor U25379 (N_25379,N_24726,N_24349);
nor U25380 (N_25380,N_24653,N_24723);
and U25381 (N_25381,N_24586,N_24179);
nand U25382 (N_25382,N_24668,N_24102);
and U25383 (N_25383,N_24296,N_24282);
or U25384 (N_25384,N_24335,N_24988);
and U25385 (N_25385,N_24651,N_24098);
nand U25386 (N_25386,N_24984,N_24140);
xnor U25387 (N_25387,N_24741,N_24251);
xor U25388 (N_25388,N_24738,N_24800);
or U25389 (N_25389,N_24551,N_24475);
nand U25390 (N_25390,N_24231,N_24246);
and U25391 (N_25391,N_24494,N_24480);
nor U25392 (N_25392,N_24861,N_24358);
xor U25393 (N_25393,N_24830,N_24180);
xnor U25394 (N_25394,N_24752,N_24299);
and U25395 (N_25395,N_24160,N_24863);
nand U25396 (N_25396,N_24060,N_24719);
and U25397 (N_25397,N_24089,N_24474);
and U25398 (N_25398,N_24897,N_24292);
nor U25399 (N_25399,N_24139,N_24505);
nor U25400 (N_25400,N_24950,N_24110);
nor U25401 (N_25401,N_24987,N_24162);
nand U25402 (N_25402,N_24356,N_24442);
nand U25403 (N_25403,N_24613,N_24083);
xor U25404 (N_25404,N_24734,N_24643);
xnor U25405 (N_25405,N_24817,N_24265);
and U25406 (N_25406,N_24487,N_24410);
or U25407 (N_25407,N_24352,N_24013);
nand U25408 (N_25408,N_24869,N_24196);
or U25409 (N_25409,N_24161,N_24872);
nor U25410 (N_25410,N_24891,N_24587);
nand U25411 (N_25411,N_24366,N_24343);
and U25412 (N_25412,N_24135,N_24688);
and U25413 (N_25413,N_24759,N_24926);
xor U25414 (N_25414,N_24832,N_24791);
or U25415 (N_25415,N_24323,N_24134);
or U25416 (N_25416,N_24022,N_24692);
xor U25417 (N_25417,N_24167,N_24434);
xnor U25418 (N_25418,N_24685,N_24616);
or U25419 (N_25419,N_24310,N_24516);
xnor U25420 (N_25420,N_24050,N_24483);
nand U25421 (N_25421,N_24239,N_24874);
nand U25422 (N_25422,N_24184,N_24372);
nand U25423 (N_25423,N_24425,N_24745);
nor U25424 (N_25424,N_24177,N_24170);
or U25425 (N_25425,N_24042,N_24879);
or U25426 (N_25426,N_24081,N_24939);
nor U25427 (N_25427,N_24374,N_24399);
or U25428 (N_25428,N_24923,N_24385);
nor U25429 (N_25429,N_24746,N_24330);
or U25430 (N_25430,N_24803,N_24051);
or U25431 (N_25431,N_24203,N_24201);
xor U25432 (N_25432,N_24076,N_24877);
and U25433 (N_25433,N_24202,N_24502);
and U25434 (N_25434,N_24816,N_24462);
nand U25435 (N_25435,N_24411,N_24136);
xnor U25436 (N_25436,N_24749,N_24164);
and U25437 (N_25437,N_24866,N_24394);
nand U25438 (N_25438,N_24954,N_24293);
nand U25439 (N_25439,N_24294,N_24439);
or U25440 (N_25440,N_24608,N_24331);
and U25441 (N_25441,N_24618,N_24503);
nand U25442 (N_25442,N_24325,N_24286);
and U25443 (N_25443,N_24432,N_24936);
and U25444 (N_25444,N_24392,N_24914);
xor U25445 (N_25445,N_24084,N_24145);
nand U25446 (N_25446,N_24951,N_24760);
nor U25447 (N_25447,N_24088,N_24262);
nor U25448 (N_25448,N_24683,N_24755);
and U25449 (N_25449,N_24508,N_24332);
nand U25450 (N_25450,N_24023,N_24308);
nor U25451 (N_25451,N_24108,N_24578);
and U25452 (N_25452,N_24841,N_24854);
nor U25453 (N_25453,N_24941,N_24353);
nand U25454 (N_25454,N_24364,N_24260);
or U25455 (N_25455,N_24283,N_24340);
and U25456 (N_25456,N_24704,N_24567);
xnor U25457 (N_25457,N_24216,N_24777);
or U25458 (N_25458,N_24302,N_24641);
nor U25459 (N_25459,N_24345,N_24057);
nand U25460 (N_25460,N_24341,N_24056);
or U25461 (N_25461,N_24983,N_24548);
xnor U25462 (N_25462,N_24837,N_24737);
or U25463 (N_25463,N_24671,N_24566);
nand U25464 (N_25464,N_24842,N_24383);
or U25465 (N_25465,N_24696,N_24021);
or U25466 (N_25466,N_24141,N_24786);
nand U25467 (N_25467,N_24457,N_24424);
or U25468 (N_25468,N_24585,N_24258);
nor U25469 (N_25469,N_24066,N_24068);
xnor U25470 (N_25470,N_24811,N_24063);
nand U25471 (N_25471,N_24929,N_24312);
nand U25472 (N_25472,N_24437,N_24200);
xnor U25473 (N_25473,N_24774,N_24298);
and U25474 (N_25474,N_24568,N_24862);
nand U25475 (N_25475,N_24314,N_24970);
nor U25476 (N_25476,N_24933,N_24606);
nor U25477 (N_25477,N_24535,N_24386);
or U25478 (N_25478,N_24072,N_24473);
xor U25479 (N_25479,N_24334,N_24985);
or U25480 (N_25480,N_24905,N_24768);
nand U25481 (N_25481,N_24041,N_24100);
xor U25482 (N_25482,N_24166,N_24125);
xor U25483 (N_25483,N_24065,N_24030);
xor U25484 (N_25484,N_24220,N_24252);
xor U25485 (N_25485,N_24163,N_24354);
nand U25486 (N_25486,N_24289,N_24459);
or U25487 (N_25487,N_24270,N_24396);
nand U25488 (N_25488,N_24775,N_24703);
or U25489 (N_25489,N_24684,N_24091);
and U25490 (N_25490,N_24420,N_24596);
nand U25491 (N_25491,N_24395,N_24589);
or U25492 (N_25492,N_24346,N_24949);
and U25493 (N_25493,N_24128,N_24529);
and U25494 (N_25494,N_24344,N_24835);
and U25495 (N_25495,N_24456,N_24829);
nand U25496 (N_25496,N_24470,N_24182);
nand U25497 (N_25497,N_24039,N_24978);
nor U25498 (N_25498,N_24275,N_24397);
nor U25499 (N_25499,N_24452,N_24676);
nor U25500 (N_25500,N_24317,N_24423);
or U25501 (N_25501,N_24415,N_24025);
or U25502 (N_25502,N_24591,N_24261);
and U25503 (N_25503,N_24436,N_24865);
nand U25504 (N_25504,N_24047,N_24113);
or U25505 (N_25505,N_24055,N_24452);
and U25506 (N_25506,N_24331,N_24513);
xor U25507 (N_25507,N_24408,N_24954);
nor U25508 (N_25508,N_24905,N_24416);
and U25509 (N_25509,N_24340,N_24429);
nor U25510 (N_25510,N_24925,N_24122);
or U25511 (N_25511,N_24431,N_24159);
xnor U25512 (N_25512,N_24749,N_24633);
xnor U25513 (N_25513,N_24124,N_24834);
xnor U25514 (N_25514,N_24456,N_24268);
nand U25515 (N_25515,N_24733,N_24074);
xor U25516 (N_25516,N_24980,N_24962);
and U25517 (N_25517,N_24344,N_24536);
and U25518 (N_25518,N_24776,N_24803);
nor U25519 (N_25519,N_24498,N_24412);
nand U25520 (N_25520,N_24494,N_24879);
nor U25521 (N_25521,N_24187,N_24132);
nor U25522 (N_25522,N_24823,N_24089);
or U25523 (N_25523,N_24942,N_24085);
nor U25524 (N_25524,N_24814,N_24196);
xor U25525 (N_25525,N_24078,N_24022);
and U25526 (N_25526,N_24846,N_24302);
nand U25527 (N_25527,N_24106,N_24662);
and U25528 (N_25528,N_24545,N_24821);
nand U25529 (N_25529,N_24568,N_24971);
and U25530 (N_25530,N_24404,N_24938);
nor U25531 (N_25531,N_24467,N_24476);
and U25532 (N_25532,N_24649,N_24882);
or U25533 (N_25533,N_24550,N_24321);
nand U25534 (N_25534,N_24964,N_24732);
or U25535 (N_25535,N_24232,N_24512);
and U25536 (N_25536,N_24409,N_24899);
or U25537 (N_25537,N_24703,N_24004);
nor U25538 (N_25538,N_24888,N_24979);
and U25539 (N_25539,N_24876,N_24601);
and U25540 (N_25540,N_24121,N_24355);
nor U25541 (N_25541,N_24694,N_24825);
nand U25542 (N_25542,N_24398,N_24252);
xnor U25543 (N_25543,N_24616,N_24200);
nand U25544 (N_25544,N_24264,N_24109);
and U25545 (N_25545,N_24171,N_24148);
or U25546 (N_25546,N_24711,N_24277);
and U25547 (N_25547,N_24565,N_24640);
or U25548 (N_25548,N_24520,N_24239);
or U25549 (N_25549,N_24475,N_24520);
nor U25550 (N_25550,N_24221,N_24917);
and U25551 (N_25551,N_24891,N_24174);
nor U25552 (N_25552,N_24468,N_24731);
nor U25553 (N_25553,N_24447,N_24723);
xor U25554 (N_25554,N_24299,N_24424);
or U25555 (N_25555,N_24758,N_24303);
and U25556 (N_25556,N_24963,N_24106);
or U25557 (N_25557,N_24545,N_24678);
nand U25558 (N_25558,N_24614,N_24140);
xnor U25559 (N_25559,N_24941,N_24524);
and U25560 (N_25560,N_24582,N_24488);
or U25561 (N_25561,N_24476,N_24647);
xnor U25562 (N_25562,N_24160,N_24839);
nand U25563 (N_25563,N_24467,N_24652);
or U25564 (N_25564,N_24650,N_24942);
or U25565 (N_25565,N_24273,N_24846);
nand U25566 (N_25566,N_24740,N_24998);
nand U25567 (N_25567,N_24282,N_24851);
or U25568 (N_25568,N_24091,N_24675);
xor U25569 (N_25569,N_24988,N_24830);
nand U25570 (N_25570,N_24257,N_24144);
or U25571 (N_25571,N_24000,N_24067);
nor U25572 (N_25572,N_24013,N_24318);
nor U25573 (N_25573,N_24200,N_24835);
xnor U25574 (N_25574,N_24988,N_24833);
nor U25575 (N_25575,N_24522,N_24450);
and U25576 (N_25576,N_24143,N_24553);
nor U25577 (N_25577,N_24740,N_24102);
nor U25578 (N_25578,N_24622,N_24116);
nand U25579 (N_25579,N_24678,N_24433);
nor U25580 (N_25580,N_24778,N_24552);
nand U25581 (N_25581,N_24384,N_24291);
nand U25582 (N_25582,N_24928,N_24264);
nand U25583 (N_25583,N_24122,N_24130);
nor U25584 (N_25584,N_24839,N_24904);
nand U25585 (N_25585,N_24033,N_24276);
nand U25586 (N_25586,N_24291,N_24620);
xor U25587 (N_25587,N_24231,N_24754);
and U25588 (N_25588,N_24566,N_24376);
or U25589 (N_25589,N_24035,N_24304);
and U25590 (N_25590,N_24694,N_24129);
and U25591 (N_25591,N_24905,N_24641);
nor U25592 (N_25592,N_24119,N_24995);
and U25593 (N_25593,N_24051,N_24758);
nor U25594 (N_25594,N_24162,N_24790);
xor U25595 (N_25595,N_24857,N_24014);
xnor U25596 (N_25596,N_24849,N_24070);
xnor U25597 (N_25597,N_24542,N_24119);
nand U25598 (N_25598,N_24144,N_24414);
nand U25599 (N_25599,N_24641,N_24243);
nor U25600 (N_25600,N_24350,N_24858);
or U25601 (N_25601,N_24629,N_24652);
xnor U25602 (N_25602,N_24363,N_24108);
xnor U25603 (N_25603,N_24948,N_24363);
and U25604 (N_25604,N_24933,N_24616);
or U25605 (N_25605,N_24735,N_24368);
and U25606 (N_25606,N_24424,N_24837);
nor U25607 (N_25607,N_24326,N_24913);
nor U25608 (N_25608,N_24356,N_24825);
nand U25609 (N_25609,N_24082,N_24283);
xnor U25610 (N_25610,N_24213,N_24546);
and U25611 (N_25611,N_24170,N_24338);
nor U25612 (N_25612,N_24643,N_24567);
nor U25613 (N_25613,N_24790,N_24912);
or U25614 (N_25614,N_24367,N_24010);
nand U25615 (N_25615,N_24121,N_24246);
or U25616 (N_25616,N_24648,N_24323);
or U25617 (N_25617,N_24175,N_24690);
and U25618 (N_25618,N_24273,N_24448);
and U25619 (N_25619,N_24515,N_24318);
or U25620 (N_25620,N_24490,N_24886);
nand U25621 (N_25621,N_24192,N_24684);
xnor U25622 (N_25622,N_24529,N_24235);
xor U25623 (N_25623,N_24603,N_24319);
and U25624 (N_25624,N_24720,N_24393);
nor U25625 (N_25625,N_24273,N_24364);
and U25626 (N_25626,N_24300,N_24786);
nor U25627 (N_25627,N_24238,N_24333);
and U25628 (N_25628,N_24513,N_24436);
nand U25629 (N_25629,N_24565,N_24892);
nor U25630 (N_25630,N_24669,N_24086);
xnor U25631 (N_25631,N_24697,N_24983);
nor U25632 (N_25632,N_24637,N_24422);
xor U25633 (N_25633,N_24145,N_24890);
nand U25634 (N_25634,N_24762,N_24719);
and U25635 (N_25635,N_24188,N_24798);
nand U25636 (N_25636,N_24748,N_24716);
and U25637 (N_25637,N_24050,N_24691);
and U25638 (N_25638,N_24580,N_24910);
nor U25639 (N_25639,N_24879,N_24361);
nor U25640 (N_25640,N_24458,N_24721);
or U25641 (N_25641,N_24906,N_24465);
nand U25642 (N_25642,N_24817,N_24778);
nand U25643 (N_25643,N_24767,N_24399);
xor U25644 (N_25644,N_24496,N_24849);
nor U25645 (N_25645,N_24791,N_24349);
and U25646 (N_25646,N_24471,N_24313);
nor U25647 (N_25647,N_24002,N_24551);
and U25648 (N_25648,N_24807,N_24348);
nor U25649 (N_25649,N_24316,N_24934);
or U25650 (N_25650,N_24100,N_24610);
nand U25651 (N_25651,N_24957,N_24224);
nand U25652 (N_25652,N_24465,N_24641);
nand U25653 (N_25653,N_24976,N_24220);
nor U25654 (N_25654,N_24131,N_24496);
or U25655 (N_25655,N_24131,N_24440);
or U25656 (N_25656,N_24946,N_24033);
nand U25657 (N_25657,N_24195,N_24597);
nand U25658 (N_25658,N_24908,N_24368);
or U25659 (N_25659,N_24730,N_24444);
or U25660 (N_25660,N_24617,N_24264);
or U25661 (N_25661,N_24868,N_24153);
xnor U25662 (N_25662,N_24828,N_24350);
or U25663 (N_25663,N_24777,N_24138);
nand U25664 (N_25664,N_24819,N_24156);
xor U25665 (N_25665,N_24608,N_24697);
xor U25666 (N_25666,N_24799,N_24209);
nor U25667 (N_25667,N_24747,N_24933);
xnor U25668 (N_25668,N_24359,N_24511);
and U25669 (N_25669,N_24794,N_24879);
nand U25670 (N_25670,N_24771,N_24917);
or U25671 (N_25671,N_24075,N_24678);
nand U25672 (N_25672,N_24157,N_24259);
and U25673 (N_25673,N_24971,N_24282);
xor U25674 (N_25674,N_24827,N_24295);
and U25675 (N_25675,N_24777,N_24023);
nor U25676 (N_25676,N_24535,N_24758);
nor U25677 (N_25677,N_24438,N_24405);
and U25678 (N_25678,N_24240,N_24971);
and U25679 (N_25679,N_24133,N_24997);
and U25680 (N_25680,N_24667,N_24347);
nand U25681 (N_25681,N_24119,N_24741);
or U25682 (N_25682,N_24397,N_24058);
or U25683 (N_25683,N_24583,N_24433);
and U25684 (N_25684,N_24018,N_24836);
nand U25685 (N_25685,N_24298,N_24698);
xor U25686 (N_25686,N_24756,N_24652);
nor U25687 (N_25687,N_24633,N_24447);
xnor U25688 (N_25688,N_24712,N_24449);
and U25689 (N_25689,N_24159,N_24291);
or U25690 (N_25690,N_24653,N_24157);
nor U25691 (N_25691,N_24941,N_24243);
and U25692 (N_25692,N_24606,N_24031);
or U25693 (N_25693,N_24467,N_24993);
and U25694 (N_25694,N_24070,N_24903);
nor U25695 (N_25695,N_24478,N_24302);
and U25696 (N_25696,N_24301,N_24723);
nor U25697 (N_25697,N_24462,N_24738);
and U25698 (N_25698,N_24573,N_24328);
or U25699 (N_25699,N_24234,N_24736);
and U25700 (N_25700,N_24394,N_24957);
nand U25701 (N_25701,N_24908,N_24856);
xor U25702 (N_25702,N_24373,N_24446);
nor U25703 (N_25703,N_24331,N_24058);
xor U25704 (N_25704,N_24309,N_24535);
xnor U25705 (N_25705,N_24291,N_24279);
nor U25706 (N_25706,N_24580,N_24005);
nor U25707 (N_25707,N_24748,N_24580);
xor U25708 (N_25708,N_24611,N_24559);
nand U25709 (N_25709,N_24474,N_24524);
nand U25710 (N_25710,N_24914,N_24668);
or U25711 (N_25711,N_24294,N_24653);
or U25712 (N_25712,N_24669,N_24604);
xnor U25713 (N_25713,N_24856,N_24250);
or U25714 (N_25714,N_24280,N_24512);
nor U25715 (N_25715,N_24924,N_24038);
nand U25716 (N_25716,N_24238,N_24628);
and U25717 (N_25717,N_24113,N_24027);
nor U25718 (N_25718,N_24326,N_24587);
and U25719 (N_25719,N_24430,N_24437);
nand U25720 (N_25720,N_24165,N_24617);
and U25721 (N_25721,N_24818,N_24802);
xor U25722 (N_25722,N_24528,N_24526);
nand U25723 (N_25723,N_24449,N_24111);
and U25724 (N_25724,N_24168,N_24564);
nand U25725 (N_25725,N_24672,N_24325);
and U25726 (N_25726,N_24812,N_24661);
nand U25727 (N_25727,N_24298,N_24362);
xor U25728 (N_25728,N_24578,N_24501);
nor U25729 (N_25729,N_24539,N_24344);
or U25730 (N_25730,N_24657,N_24105);
xor U25731 (N_25731,N_24730,N_24114);
nand U25732 (N_25732,N_24677,N_24945);
nor U25733 (N_25733,N_24681,N_24953);
and U25734 (N_25734,N_24569,N_24568);
nor U25735 (N_25735,N_24534,N_24485);
nor U25736 (N_25736,N_24908,N_24793);
xor U25737 (N_25737,N_24989,N_24844);
nor U25738 (N_25738,N_24578,N_24541);
xor U25739 (N_25739,N_24151,N_24280);
xor U25740 (N_25740,N_24981,N_24473);
and U25741 (N_25741,N_24652,N_24037);
xor U25742 (N_25742,N_24858,N_24787);
and U25743 (N_25743,N_24788,N_24156);
or U25744 (N_25744,N_24713,N_24799);
xnor U25745 (N_25745,N_24258,N_24236);
or U25746 (N_25746,N_24188,N_24782);
nand U25747 (N_25747,N_24003,N_24461);
nor U25748 (N_25748,N_24043,N_24386);
or U25749 (N_25749,N_24656,N_24097);
nand U25750 (N_25750,N_24692,N_24118);
nor U25751 (N_25751,N_24447,N_24668);
nor U25752 (N_25752,N_24407,N_24457);
xor U25753 (N_25753,N_24460,N_24432);
xor U25754 (N_25754,N_24369,N_24325);
or U25755 (N_25755,N_24049,N_24215);
nand U25756 (N_25756,N_24097,N_24720);
nand U25757 (N_25757,N_24646,N_24518);
xnor U25758 (N_25758,N_24383,N_24316);
xnor U25759 (N_25759,N_24126,N_24583);
or U25760 (N_25760,N_24366,N_24697);
nand U25761 (N_25761,N_24014,N_24846);
xnor U25762 (N_25762,N_24416,N_24941);
nand U25763 (N_25763,N_24695,N_24984);
and U25764 (N_25764,N_24172,N_24293);
xor U25765 (N_25765,N_24590,N_24931);
nor U25766 (N_25766,N_24923,N_24672);
nor U25767 (N_25767,N_24090,N_24011);
or U25768 (N_25768,N_24661,N_24854);
xor U25769 (N_25769,N_24937,N_24858);
and U25770 (N_25770,N_24916,N_24643);
or U25771 (N_25771,N_24691,N_24675);
or U25772 (N_25772,N_24585,N_24212);
and U25773 (N_25773,N_24924,N_24676);
xor U25774 (N_25774,N_24912,N_24832);
nand U25775 (N_25775,N_24480,N_24595);
and U25776 (N_25776,N_24641,N_24691);
and U25777 (N_25777,N_24547,N_24128);
or U25778 (N_25778,N_24931,N_24673);
nor U25779 (N_25779,N_24808,N_24626);
and U25780 (N_25780,N_24129,N_24094);
xor U25781 (N_25781,N_24131,N_24274);
nand U25782 (N_25782,N_24198,N_24713);
xnor U25783 (N_25783,N_24504,N_24519);
and U25784 (N_25784,N_24417,N_24075);
xnor U25785 (N_25785,N_24672,N_24367);
nor U25786 (N_25786,N_24638,N_24979);
and U25787 (N_25787,N_24941,N_24141);
xor U25788 (N_25788,N_24371,N_24102);
nand U25789 (N_25789,N_24098,N_24878);
and U25790 (N_25790,N_24768,N_24732);
nor U25791 (N_25791,N_24503,N_24239);
and U25792 (N_25792,N_24957,N_24805);
nand U25793 (N_25793,N_24184,N_24046);
xnor U25794 (N_25794,N_24154,N_24877);
xnor U25795 (N_25795,N_24791,N_24089);
xor U25796 (N_25796,N_24122,N_24118);
xor U25797 (N_25797,N_24045,N_24687);
xor U25798 (N_25798,N_24186,N_24344);
or U25799 (N_25799,N_24679,N_24733);
or U25800 (N_25800,N_24094,N_24611);
or U25801 (N_25801,N_24843,N_24739);
nand U25802 (N_25802,N_24067,N_24906);
nor U25803 (N_25803,N_24178,N_24626);
or U25804 (N_25804,N_24378,N_24182);
xnor U25805 (N_25805,N_24216,N_24234);
xor U25806 (N_25806,N_24470,N_24758);
xnor U25807 (N_25807,N_24065,N_24676);
nor U25808 (N_25808,N_24122,N_24649);
and U25809 (N_25809,N_24746,N_24349);
and U25810 (N_25810,N_24370,N_24316);
or U25811 (N_25811,N_24206,N_24755);
xnor U25812 (N_25812,N_24201,N_24045);
xor U25813 (N_25813,N_24061,N_24966);
and U25814 (N_25814,N_24296,N_24766);
and U25815 (N_25815,N_24930,N_24268);
and U25816 (N_25816,N_24129,N_24838);
and U25817 (N_25817,N_24367,N_24768);
nand U25818 (N_25818,N_24720,N_24460);
xnor U25819 (N_25819,N_24750,N_24518);
nand U25820 (N_25820,N_24301,N_24928);
nor U25821 (N_25821,N_24275,N_24689);
nor U25822 (N_25822,N_24304,N_24521);
nor U25823 (N_25823,N_24297,N_24911);
nor U25824 (N_25824,N_24970,N_24951);
xor U25825 (N_25825,N_24694,N_24180);
nor U25826 (N_25826,N_24309,N_24443);
xor U25827 (N_25827,N_24637,N_24269);
nand U25828 (N_25828,N_24024,N_24799);
or U25829 (N_25829,N_24386,N_24021);
or U25830 (N_25830,N_24086,N_24353);
xnor U25831 (N_25831,N_24317,N_24792);
or U25832 (N_25832,N_24466,N_24097);
and U25833 (N_25833,N_24696,N_24182);
xor U25834 (N_25834,N_24260,N_24408);
and U25835 (N_25835,N_24615,N_24218);
nor U25836 (N_25836,N_24817,N_24264);
nand U25837 (N_25837,N_24844,N_24515);
or U25838 (N_25838,N_24544,N_24297);
nand U25839 (N_25839,N_24098,N_24565);
and U25840 (N_25840,N_24388,N_24727);
xnor U25841 (N_25841,N_24485,N_24846);
xnor U25842 (N_25842,N_24329,N_24649);
and U25843 (N_25843,N_24862,N_24593);
nor U25844 (N_25844,N_24365,N_24559);
or U25845 (N_25845,N_24897,N_24016);
or U25846 (N_25846,N_24063,N_24509);
nor U25847 (N_25847,N_24250,N_24560);
or U25848 (N_25848,N_24385,N_24201);
nor U25849 (N_25849,N_24268,N_24779);
and U25850 (N_25850,N_24949,N_24552);
nor U25851 (N_25851,N_24883,N_24838);
and U25852 (N_25852,N_24110,N_24881);
xnor U25853 (N_25853,N_24413,N_24109);
and U25854 (N_25854,N_24333,N_24031);
xnor U25855 (N_25855,N_24331,N_24987);
or U25856 (N_25856,N_24465,N_24675);
and U25857 (N_25857,N_24125,N_24151);
or U25858 (N_25858,N_24968,N_24951);
xor U25859 (N_25859,N_24347,N_24959);
xnor U25860 (N_25860,N_24487,N_24318);
and U25861 (N_25861,N_24911,N_24164);
or U25862 (N_25862,N_24192,N_24807);
or U25863 (N_25863,N_24573,N_24644);
nand U25864 (N_25864,N_24110,N_24279);
or U25865 (N_25865,N_24503,N_24608);
nand U25866 (N_25866,N_24156,N_24287);
xor U25867 (N_25867,N_24266,N_24071);
and U25868 (N_25868,N_24815,N_24341);
nand U25869 (N_25869,N_24406,N_24518);
and U25870 (N_25870,N_24813,N_24351);
and U25871 (N_25871,N_24141,N_24857);
and U25872 (N_25872,N_24626,N_24002);
or U25873 (N_25873,N_24971,N_24013);
and U25874 (N_25874,N_24904,N_24734);
xnor U25875 (N_25875,N_24149,N_24525);
or U25876 (N_25876,N_24113,N_24898);
nand U25877 (N_25877,N_24805,N_24375);
xnor U25878 (N_25878,N_24200,N_24453);
or U25879 (N_25879,N_24910,N_24962);
or U25880 (N_25880,N_24159,N_24651);
or U25881 (N_25881,N_24703,N_24961);
nand U25882 (N_25882,N_24905,N_24563);
and U25883 (N_25883,N_24504,N_24267);
nor U25884 (N_25884,N_24621,N_24768);
nor U25885 (N_25885,N_24290,N_24313);
xor U25886 (N_25886,N_24934,N_24799);
xnor U25887 (N_25887,N_24654,N_24578);
xor U25888 (N_25888,N_24985,N_24687);
nor U25889 (N_25889,N_24444,N_24623);
xnor U25890 (N_25890,N_24902,N_24758);
nor U25891 (N_25891,N_24036,N_24636);
nor U25892 (N_25892,N_24584,N_24006);
nand U25893 (N_25893,N_24272,N_24619);
xnor U25894 (N_25894,N_24348,N_24504);
xor U25895 (N_25895,N_24789,N_24262);
nand U25896 (N_25896,N_24047,N_24888);
nand U25897 (N_25897,N_24484,N_24749);
and U25898 (N_25898,N_24582,N_24315);
or U25899 (N_25899,N_24141,N_24768);
and U25900 (N_25900,N_24069,N_24118);
and U25901 (N_25901,N_24397,N_24416);
xor U25902 (N_25902,N_24911,N_24774);
and U25903 (N_25903,N_24719,N_24230);
nand U25904 (N_25904,N_24033,N_24153);
nand U25905 (N_25905,N_24883,N_24517);
xor U25906 (N_25906,N_24504,N_24242);
xnor U25907 (N_25907,N_24381,N_24466);
or U25908 (N_25908,N_24920,N_24448);
nand U25909 (N_25909,N_24995,N_24251);
and U25910 (N_25910,N_24830,N_24521);
and U25911 (N_25911,N_24759,N_24967);
and U25912 (N_25912,N_24258,N_24018);
nor U25913 (N_25913,N_24898,N_24048);
nand U25914 (N_25914,N_24280,N_24921);
nand U25915 (N_25915,N_24485,N_24218);
or U25916 (N_25916,N_24046,N_24922);
nand U25917 (N_25917,N_24940,N_24404);
and U25918 (N_25918,N_24666,N_24664);
xnor U25919 (N_25919,N_24513,N_24231);
xor U25920 (N_25920,N_24452,N_24376);
and U25921 (N_25921,N_24370,N_24206);
or U25922 (N_25922,N_24971,N_24199);
nand U25923 (N_25923,N_24102,N_24261);
nand U25924 (N_25924,N_24426,N_24594);
nor U25925 (N_25925,N_24805,N_24746);
or U25926 (N_25926,N_24712,N_24586);
or U25927 (N_25927,N_24050,N_24861);
or U25928 (N_25928,N_24479,N_24675);
xor U25929 (N_25929,N_24544,N_24158);
nand U25930 (N_25930,N_24725,N_24847);
or U25931 (N_25931,N_24098,N_24595);
xnor U25932 (N_25932,N_24794,N_24931);
and U25933 (N_25933,N_24131,N_24540);
or U25934 (N_25934,N_24304,N_24123);
nand U25935 (N_25935,N_24149,N_24216);
or U25936 (N_25936,N_24979,N_24407);
nor U25937 (N_25937,N_24132,N_24007);
xor U25938 (N_25938,N_24973,N_24681);
or U25939 (N_25939,N_24578,N_24923);
and U25940 (N_25940,N_24862,N_24528);
or U25941 (N_25941,N_24044,N_24060);
nand U25942 (N_25942,N_24962,N_24322);
xnor U25943 (N_25943,N_24232,N_24093);
and U25944 (N_25944,N_24725,N_24525);
or U25945 (N_25945,N_24151,N_24956);
and U25946 (N_25946,N_24339,N_24481);
xor U25947 (N_25947,N_24280,N_24433);
nor U25948 (N_25948,N_24662,N_24017);
nand U25949 (N_25949,N_24020,N_24458);
nand U25950 (N_25950,N_24960,N_24300);
nor U25951 (N_25951,N_24776,N_24556);
xor U25952 (N_25952,N_24564,N_24587);
nand U25953 (N_25953,N_24833,N_24749);
and U25954 (N_25954,N_24211,N_24722);
xnor U25955 (N_25955,N_24075,N_24566);
xor U25956 (N_25956,N_24106,N_24118);
and U25957 (N_25957,N_24823,N_24537);
and U25958 (N_25958,N_24635,N_24102);
or U25959 (N_25959,N_24837,N_24670);
nor U25960 (N_25960,N_24377,N_24214);
xor U25961 (N_25961,N_24740,N_24317);
xor U25962 (N_25962,N_24728,N_24770);
nand U25963 (N_25963,N_24965,N_24250);
nor U25964 (N_25964,N_24870,N_24643);
and U25965 (N_25965,N_24004,N_24194);
and U25966 (N_25966,N_24129,N_24275);
nor U25967 (N_25967,N_24369,N_24885);
or U25968 (N_25968,N_24073,N_24896);
xnor U25969 (N_25969,N_24912,N_24525);
nor U25970 (N_25970,N_24992,N_24549);
or U25971 (N_25971,N_24906,N_24917);
nor U25972 (N_25972,N_24664,N_24262);
and U25973 (N_25973,N_24213,N_24935);
xor U25974 (N_25974,N_24741,N_24231);
nor U25975 (N_25975,N_24662,N_24589);
nand U25976 (N_25976,N_24622,N_24479);
nor U25977 (N_25977,N_24986,N_24270);
or U25978 (N_25978,N_24138,N_24652);
or U25979 (N_25979,N_24394,N_24992);
or U25980 (N_25980,N_24881,N_24303);
and U25981 (N_25981,N_24726,N_24252);
and U25982 (N_25982,N_24340,N_24500);
nand U25983 (N_25983,N_24228,N_24351);
nor U25984 (N_25984,N_24828,N_24056);
and U25985 (N_25985,N_24701,N_24817);
xnor U25986 (N_25986,N_24985,N_24387);
xnor U25987 (N_25987,N_24143,N_24803);
xnor U25988 (N_25988,N_24555,N_24422);
nor U25989 (N_25989,N_24956,N_24369);
nand U25990 (N_25990,N_24345,N_24661);
nor U25991 (N_25991,N_24383,N_24696);
or U25992 (N_25992,N_24329,N_24381);
or U25993 (N_25993,N_24227,N_24368);
nor U25994 (N_25994,N_24549,N_24914);
or U25995 (N_25995,N_24247,N_24935);
nand U25996 (N_25996,N_24437,N_24632);
nand U25997 (N_25997,N_24050,N_24757);
nand U25998 (N_25998,N_24334,N_24388);
nor U25999 (N_25999,N_24523,N_24434);
and U26000 (N_26000,N_25754,N_25435);
xor U26001 (N_26001,N_25115,N_25133);
and U26002 (N_26002,N_25048,N_25781);
nand U26003 (N_26003,N_25071,N_25042);
and U26004 (N_26004,N_25338,N_25403);
and U26005 (N_26005,N_25441,N_25278);
nand U26006 (N_26006,N_25503,N_25907);
nor U26007 (N_26007,N_25470,N_25149);
and U26008 (N_26008,N_25995,N_25455);
xor U26009 (N_26009,N_25808,N_25564);
or U26010 (N_26010,N_25237,N_25127);
or U26011 (N_26011,N_25467,N_25955);
and U26012 (N_26012,N_25529,N_25140);
xor U26013 (N_26013,N_25980,N_25898);
nand U26014 (N_26014,N_25689,N_25328);
nor U26015 (N_26015,N_25705,N_25628);
nand U26016 (N_26016,N_25335,N_25703);
or U26017 (N_26017,N_25276,N_25421);
nand U26018 (N_26018,N_25804,N_25119);
nand U26019 (N_26019,N_25256,N_25638);
nor U26020 (N_26020,N_25642,N_25893);
and U26021 (N_26021,N_25481,N_25442);
xor U26022 (N_26022,N_25682,N_25318);
nand U26023 (N_26023,N_25162,N_25692);
nand U26024 (N_26024,N_25685,N_25411);
xnor U26025 (N_26025,N_25444,N_25533);
nand U26026 (N_26026,N_25041,N_25590);
nand U26027 (N_26027,N_25148,N_25539);
nand U26028 (N_26028,N_25005,N_25413);
xor U26029 (N_26029,N_25227,N_25132);
nand U26030 (N_26030,N_25687,N_25963);
or U26031 (N_26031,N_25293,N_25017);
and U26032 (N_26032,N_25561,N_25185);
xnor U26033 (N_26033,N_25888,N_25816);
nor U26034 (N_26034,N_25698,N_25832);
xor U26035 (N_26035,N_25544,N_25345);
nand U26036 (N_26036,N_25262,N_25172);
nand U26037 (N_26037,N_25348,N_25106);
and U26038 (N_26038,N_25131,N_25962);
and U26039 (N_26039,N_25226,N_25667);
nand U26040 (N_26040,N_25213,N_25061);
xnor U26041 (N_26041,N_25908,N_25329);
nor U26042 (N_26042,N_25958,N_25505);
and U26043 (N_26043,N_25849,N_25571);
xnor U26044 (N_26044,N_25979,N_25721);
or U26045 (N_26045,N_25379,N_25299);
or U26046 (N_26046,N_25502,N_25233);
and U26047 (N_26047,N_25507,N_25916);
and U26048 (N_26048,N_25179,N_25271);
or U26049 (N_26049,N_25091,N_25279);
nand U26050 (N_26050,N_25759,N_25225);
nor U26051 (N_26051,N_25538,N_25404);
and U26052 (N_26052,N_25641,N_25987);
xor U26053 (N_26053,N_25825,N_25102);
nand U26054 (N_26054,N_25289,N_25426);
or U26055 (N_26055,N_25531,N_25863);
and U26056 (N_26056,N_25474,N_25866);
xor U26057 (N_26057,N_25229,N_25750);
and U26058 (N_26058,N_25438,N_25761);
and U26059 (N_26059,N_25418,N_25811);
nand U26060 (N_26060,N_25722,N_25889);
nor U26061 (N_26061,N_25113,N_25559);
nand U26062 (N_26062,N_25783,N_25038);
nor U26063 (N_26063,N_25184,N_25944);
nor U26064 (N_26064,N_25314,N_25466);
or U26065 (N_26065,N_25532,N_25392);
nand U26066 (N_26066,N_25308,N_25223);
and U26067 (N_26067,N_25633,N_25190);
nor U26068 (N_26068,N_25188,N_25522);
nand U26069 (N_26069,N_25546,N_25729);
or U26070 (N_26070,N_25087,N_25499);
and U26071 (N_26071,N_25860,N_25463);
or U26072 (N_26072,N_25327,N_25152);
nor U26073 (N_26073,N_25254,N_25145);
xor U26074 (N_26074,N_25934,N_25795);
nand U26075 (N_26075,N_25769,N_25300);
xor U26076 (N_26076,N_25007,N_25550);
nor U26077 (N_26077,N_25696,N_25918);
and U26078 (N_26078,N_25187,N_25224);
or U26079 (N_26079,N_25049,N_25711);
or U26080 (N_26080,N_25373,N_25791);
or U26081 (N_26081,N_25374,N_25552);
or U26082 (N_26082,N_25519,N_25322);
xnor U26083 (N_26083,N_25647,N_25253);
and U26084 (N_26084,N_25855,N_25822);
and U26085 (N_26085,N_25746,N_25242);
nand U26086 (N_26086,N_25417,N_25974);
xor U26087 (N_26087,N_25767,N_25753);
and U26088 (N_26088,N_25891,N_25988);
or U26089 (N_26089,N_25585,N_25983);
xnor U26090 (N_26090,N_25578,N_25197);
nand U26091 (N_26091,N_25842,N_25457);
nor U26092 (N_26092,N_25240,N_25462);
and U26093 (N_26093,N_25994,N_25877);
xnor U26094 (N_26094,N_25221,N_25199);
nor U26095 (N_26095,N_25697,N_25615);
or U26096 (N_26096,N_25880,N_25527);
or U26097 (N_26097,N_25365,N_25812);
nand U26098 (N_26098,N_25357,N_25380);
or U26099 (N_26099,N_25930,N_25016);
or U26100 (N_26100,N_25259,N_25472);
xnor U26101 (N_26101,N_25015,N_25706);
nand U26102 (N_26102,N_25656,N_25551);
or U26103 (N_26103,N_25011,N_25144);
xor U26104 (N_26104,N_25086,N_25033);
nand U26105 (N_26105,N_25219,N_25266);
or U26106 (N_26106,N_25669,N_25824);
nor U26107 (N_26107,N_25116,N_25051);
xor U26108 (N_26108,N_25976,N_25101);
nor U26109 (N_26109,N_25100,N_25580);
or U26110 (N_26110,N_25699,N_25610);
xor U26111 (N_26111,N_25420,N_25449);
nor U26112 (N_26112,N_25526,N_25990);
xor U26113 (N_26113,N_25941,N_25258);
or U26114 (N_26114,N_25997,N_25122);
nor U26115 (N_26115,N_25514,N_25819);
xor U26116 (N_26116,N_25473,N_25440);
nor U26117 (N_26117,N_25634,N_25785);
nand U26118 (N_26118,N_25046,N_25768);
xor U26119 (N_26119,N_25324,N_25107);
xnor U26120 (N_26120,N_25737,N_25541);
and U26121 (N_26121,N_25375,N_25681);
or U26122 (N_26122,N_25024,N_25360);
and U26123 (N_26123,N_25347,N_25575);
or U26124 (N_26124,N_25731,N_25410);
or U26125 (N_26125,N_25920,N_25651);
nor U26126 (N_26126,N_25235,N_25913);
xnor U26127 (N_26127,N_25702,N_25872);
xnor U26128 (N_26128,N_25246,N_25215);
nor U26129 (N_26129,N_25353,N_25873);
xnor U26130 (N_26130,N_25239,N_25579);
nor U26131 (N_26131,N_25194,N_25216);
nand U26132 (N_26132,N_25813,N_25940);
and U26133 (N_26133,N_25170,N_25631);
or U26134 (N_26134,N_25728,N_25874);
xor U26135 (N_26135,N_25139,N_25727);
and U26136 (N_26136,N_25838,N_25105);
or U26137 (N_26137,N_25674,N_25283);
nor U26138 (N_26138,N_25846,N_25247);
nor U26139 (N_26139,N_25542,N_25789);
and U26140 (N_26140,N_25008,N_25182);
and U26141 (N_26141,N_25383,N_25909);
xor U26142 (N_26142,N_25910,N_25310);
or U26143 (N_26143,N_25796,N_25582);
and U26144 (N_26144,N_25207,N_25723);
or U26145 (N_26145,N_25655,N_25611);
nand U26146 (N_26146,N_25359,N_25263);
and U26147 (N_26147,N_25776,N_25097);
xnor U26148 (N_26148,N_25762,N_25884);
nor U26149 (N_26149,N_25050,N_25953);
or U26150 (N_26150,N_25361,N_25181);
and U26151 (N_26151,N_25903,N_25264);
nand U26152 (N_26152,N_25643,N_25952);
nand U26153 (N_26153,N_25053,N_25400);
and U26154 (N_26154,N_25516,N_25482);
or U26155 (N_26155,N_25065,N_25451);
nor U26156 (N_26156,N_25340,N_25217);
xor U26157 (N_26157,N_25282,N_25961);
and U26158 (N_26158,N_25810,N_25871);
xor U26159 (N_26159,N_25892,N_25174);
xor U26160 (N_26160,N_25445,N_25311);
or U26161 (N_26161,N_25999,N_25035);
and U26162 (N_26162,N_25158,N_25637);
nand U26163 (N_26163,N_25709,N_25700);
and U26164 (N_26164,N_25921,N_25675);
xor U26165 (N_26165,N_25012,N_25165);
nand U26166 (N_26166,N_25894,N_25660);
nor U26167 (N_26167,N_25972,N_25288);
or U26168 (N_26168,N_25740,N_25716);
or U26169 (N_26169,N_25592,N_25295);
or U26170 (N_26170,N_25738,N_25806);
and U26171 (N_26171,N_25415,N_25708);
and U26172 (N_26172,N_25805,N_25452);
or U26173 (N_26173,N_25000,N_25901);
nand U26174 (N_26174,N_25870,N_25704);
or U26175 (N_26175,N_25180,N_25661);
nand U26176 (N_26176,N_25847,N_25220);
xor U26177 (N_26177,N_25760,N_25336);
nand U26178 (N_26178,N_25865,N_25914);
nor U26179 (N_26179,N_25414,N_25488);
nand U26180 (N_26180,N_25298,N_25751);
nor U26181 (N_26181,N_25080,N_25946);
nor U26182 (N_26182,N_25862,N_25155);
and U26183 (N_26183,N_25784,N_25268);
and U26184 (N_26184,N_25198,N_25294);
xor U26185 (N_26185,N_25549,N_25807);
and U26186 (N_26186,N_25686,N_25437);
xor U26187 (N_26187,N_25109,N_25362);
or U26188 (N_26188,N_25124,N_25354);
or U26189 (N_26189,N_25809,N_25617);
and U26190 (N_26190,N_25334,N_25562);
xnor U26191 (N_26191,N_25817,N_25009);
xor U26192 (N_26192,N_25927,N_25161);
and U26193 (N_26193,N_25376,N_25117);
and U26194 (N_26194,N_25613,N_25234);
and U26195 (N_26195,N_25883,N_25664);
and U26196 (N_26196,N_25013,N_25540);
nor U26197 (N_26197,N_25911,N_25431);
nor U26198 (N_26198,N_25476,N_25208);
and U26199 (N_26199,N_25079,N_25545);
or U26200 (N_26200,N_25479,N_25175);
nor U26201 (N_26201,N_25222,N_25739);
or U26202 (N_26202,N_25966,N_25093);
nand U26203 (N_26203,N_25596,N_25406);
xor U26204 (N_26204,N_25570,N_25292);
nand U26205 (N_26205,N_25486,N_25287);
nor U26206 (N_26206,N_25189,N_25495);
nand U26207 (N_26207,N_25513,N_25491);
and U26208 (N_26208,N_25548,N_25301);
xnor U26209 (N_26209,N_25654,N_25019);
nand U26210 (N_26210,N_25228,N_25747);
nor U26211 (N_26211,N_25645,N_25386);
xor U26212 (N_26212,N_25153,N_25730);
xnor U26213 (N_26213,N_25173,N_25072);
nor U26214 (N_26214,N_25371,N_25304);
nand U26215 (N_26215,N_25147,N_25468);
nor U26216 (N_26216,N_25399,N_25627);
nor U26217 (N_26217,N_25430,N_25178);
xor U26218 (N_26218,N_25690,N_25986);
xor U26219 (N_26219,N_25799,N_25848);
nor U26220 (N_26220,N_25897,N_25489);
or U26221 (N_26221,N_25679,N_25853);
and U26222 (N_26222,N_25250,N_25577);
nand U26223 (N_26223,N_25625,N_25820);
nand U26224 (N_26224,N_25773,N_25114);
or U26225 (N_26225,N_25480,N_25850);
xor U26226 (N_26226,N_25028,N_25843);
or U26227 (N_26227,N_25936,N_25666);
nand U26228 (N_26228,N_25956,N_25844);
nor U26229 (N_26229,N_25066,N_25523);
and U26230 (N_26230,N_25742,N_25159);
or U26231 (N_26231,N_25981,N_25741);
xor U26232 (N_26232,N_25885,N_25942);
and U26233 (N_26233,N_25350,N_25384);
or U26234 (N_26234,N_25492,N_25830);
or U26235 (N_26235,N_25616,N_25059);
and U26236 (N_26236,N_25121,N_25394);
nand U26237 (N_26237,N_25339,N_25970);
nand U26238 (N_26238,N_25405,N_25733);
nand U26239 (N_26239,N_25663,N_25572);
and U26240 (N_26240,N_25518,N_25261);
nor U26241 (N_26241,N_25484,N_25290);
xnor U26242 (N_26242,N_25443,N_25193);
nor U26243 (N_26243,N_25764,N_25275);
xor U26244 (N_26244,N_25352,N_25211);
xor U26245 (N_26245,N_25302,N_25209);
nor U26246 (N_26246,N_25286,N_25084);
nand U26247 (N_26247,N_25230,N_25141);
or U26248 (N_26248,N_25715,N_25387);
nand U26249 (N_26249,N_25833,N_25297);
and U26250 (N_26250,N_25402,N_25475);
or U26251 (N_26251,N_25978,N_25917);
or U26252 (N_26252,N_25099,N_25867);
nor U26253 (N_26253,N_25605,N_25284);
or U26254 (N_26254,N_25555,N_25662);
nand U26255 (N_26255,N_25875,N_25382);
nand U26256 (N_26256,N_25236,N_25459);
xnor U26257 (N_26257,N_25763,N_25095);
nand U26258 (N_26258,N_25273,N_25037);
nand U26259 (N_26259,N_25834,N_25965);
xor U26260 (N_26260,N_25511,N_25325);
xnor U26261 (N_26261,N_25547,N_25945);
xor U26262 (N_26262,N_25534,N_25201);
xor U26263 (N_26263,N_25925,N_25671);
nand U26264 (N_26264,N_25063,N_25128);
nor U26265 (N_26265,N_25023,N_25563);
and U26266 (N_26266,N_25693,N_25369);
nand U26267 (N_26267,N_25932,N_25391);
and U26268 (N_26268,N_25828,N_25396);
and U26269 (N_26269,N_25589,N_25123);
nand U26270 (N_26270,N_25857,N_25358);
nor U26271 (N_26271,N_25241,N_25790);
nor U26272 (N_26272,N_25553,N_25678);
xnor U26273 (N_26273,N_25291,N_25774);
xnor U26274 (N_26274,N_25757,N_25081);
or U26275 (N_26275,N_25714,N_25797);
and U26276 (N_26276,N_25777,N_25111);
nand U26277 (N_26277,N_25659,N_25274);
xor U26278 (N_26278,N_25070,N_25969);
or U26279 (N_26279,N_25509,N_25951);
and U26280 (N_26280,N_25319,N_25416);
nand U26281 (N_26281,N_25749,N_25409);
xnor U26282 (N_26282,N_25465,N_25422);
or U26283 (N_26283,N_25136,N_25887);
or U26284 (N_26284,N_25154,N_25801);
or U26285 (N_26285,N_25082,N_25604);
nor U26286 (N_26286,N_25971,N_25881);
and U26287 (N_26287,N_25869,N_25618);
nor U26288 (N_26288,N_25321,N_25798);
xnor U26289 (N_26289,N_25535,N_25658);
and U26290 (N_26290,N_25606,N_25895);
xor U26291 (N_26291,N_25793,N_25398);
and U26292 (N_26292,N_25135,N_25342);
or U26293 (N_26293,N_25717,N_25630);
nor U26294 (N_26294,N_25831,N_25991);
and U26295 (N_26295,N_25423,N_25267);
xor U26296 (N_26296,N_25876,N_25904);
nor U26297 (N_26297,N_25501,N_25014);
or U26298 (N_26298,N_25390,N_25653);
nor U26299 (N_26299,N_25829,N_25031);
xor U26300 (N_26300,N_25040,N_25151);
nor U26301 (N_26301,N_25636,N_25203);
nor U26302 (N_26302,N_25576,N_25719);
xor U26303 (N_26303,N_25096,N_25861);
xor U26304 (N_26304,N_25525,N_25346);
xnor U26305 (N_26305,N_25926,N_25372);
nand U26306 (N_26306,N_25163,N_25609);
or U26307 (N_26307,N_25092,N_25772);
and U26308 (N_26308,N_25620,N_25977);
nand U26309 (N_26309,N_25560,N_25039);
nor U26310 (N_26310,N_25388,N_25770);
xnor U26311 (N_26311,N_25464,N_25177);
or U26312 (N_26312,N_25401,N_25214);
and U26313 (N_26313,N_25868,N_25064);
xor U26314 (N_26314,N_25982,N_25556);
and U26315 (N_26315,N_25517,N_25010);
and U26316 (N_26316,N_25103,N_25018);
and U26317 (N_26317,N_25090,N_25967);
xor U26318 (N_26318,N_25668,N_25827);
nor U26319 (N_26319,N_25270,N_25098);
and U26320 (N_26320,N_25640,N_25447);
nor U26321 (N_26321,N_25307,N_25419);
or U26322 (N_26322,N_25156,N_25998);
xnor U26323 (N_26323,N_25088,N_25677);
nor U26324 (N_26324,N_25602,N_25393);
xor U26325 (N_26325,N_25436,N_25778);
xnor U26326 (N_26326,N_25074,N_25558);
and U26327 (N_26327,N_25836,N_25608);
xor U26328 (N_26328,N_25433,N_25249);
and U26329 (N_26329,N_25500,N_25332);
and U26330 (N_26330,N_25315,N_25591);
nand U26331 (N_26331,N_25504,N_25142);
xor U26332 (N_26332,N_25672,N_25929);
nor U26333 (N_26333,N_25890,N_25823);
nand U26334 (N_26334,N_25923,N_25581);
and U26335 (N_26335,N_25412,N_25707);
nor U26336 (N_26336,N_25320,N_25766);
or U26337 (N_26337,N_25792,N_25524);
nand U26338 (N_26338,N_25204,N_25125);
and U26339 (N_26339,N_25684,N_25078);
xnor U26340 (N_26340,N_25748,N_25277);
nand U26341 (N_26341,N_25931,N_25176);
xor U26342 (N_26342,N_25954,N_25619);
and U26343 (N_26343,N_25385,N_25935);
and U26344 (N_26344,N_25231,N_25756);
and U26345 (N_26345,N_25167,N_25607);
nand U26346 (N_26346,N_25614,N_25212);
and U26347 (N_26347,N_25296,N_25164);
or U26348 (N_26348,N_25899,N_25629);
nor U26349 (N_26349,N_25782,N_25543);
and U26350 (N_26350,N_25192,N_25938);
or U26351 (N_26351,N_25368,N_25837);
or U26352 (N_26352,N_25036,N_25802);
nor U26353 (N_26353,N_25110,N_25851);
or U26354 (N_26354,N_25800,N_25052);
xnor U26355 (N_26355,N_25120,N_25303);
nand U26356 (N_26356,N_25326,N_25520);
xor U26357 (N_26357,N_25626,N_25735);
nand U26358 (N_26358,N_25134,N_25202);
nor U26359 (N_26359,N_25924,N_25725);
and U26360 (N_26360,N_25623,N_25062);
nor U26361 (N_26361,N_25157,N_25021);
nand U26362 (N_26362,N_25166,N_25530);
and U26363 (N_26363,N_25316,N_25130);
nand U26364 (N_26364,N_25752,N_25022);
and U26365 (N_26365,N_25252,N_25424);
and U26366 (N_26366,N_25205,N_25900);
and U26367 (N_26367,N_25032,N_25650);
xnor U26368 (N_26368,N_25313,N_25989);
xnor U26369 (N_26369,N_25594,N_25453);
nor U26370 (N_26370,N_25191,N_25330);
or U26371 (N_26371,N_25494,N_25960);
xnor U26372 (N_26372,N_25984,N_25788);
nand U26373 (N_26373,N_25146,N_25724);
or U26374 (N_26374,N_25691,N_25886);
or U26375 (N_26375,N_25996,N_25126);
nand U26376 (N_26376,N_25370,N_25736);
xor U26377 (N_26377,N_25355,N_25665);
nand U26378 (N_26378,N_25232,N_25478);
xnor U26379 (N_26379,N_25508,N_25928);
and U26380 (N_26380,N_25341,N_25044);
or U26381 (N_26381,N_25775,N_25281);
xnor U26382 (N_26382,N_25939,N_25429);
and U26383 (N_26383,N_25515,N_25073);
nand U26384 (N_26384,N_25493,N_25573);
and U26385 (N_26385,N_25557,N_25814);
and U26386 (N_26386,N_25600,N_25448);
and U26387 (N_26387,N_25243,N_25446);
and U26388 (N_26388,N_25461,N_25612);
nor U26389 (N_26389,N_25786,N_25821);
and U26390 (N_26390,N_25758,N_25450);
and U26391 (N_26391,N_25780,N_25160);
and U26392 (N_26392,N_25587,N_25566);
or U26393 (N_26393,N_25726,N_25859);
and U26394 (N_26394,N_25085,N_25001);
nor U26395 (N_26395,N_25057,N_25964);
and U26396 (N_26396,N_25094,N_25902);
nand U26397 (N_26397,N_25456,N_25536);
and U26398 (N_26398,N_25537,N_25569);
and U26399 (N_26399,N_25427,N_25915);
nand U26400 (N_26400,N_25129,N_25574);
or U26401 (N_26401,N_25912,N_25584);
nand U26402 (N_26402,N_25649,N_25839);
nand U26403 (N_26403,N_25644,N_25635);
and U26404 (N_26404,N_25896,N_25458);
nand U26405 (N_26405,N_25150,N_25734);
nor U26406 (N_26406,N_25510,N_25497);
xor U26407 (N_26407,N_25255,N_25864);
nand U26408 (N_26408,N_25858,N_25744);
and U26409 (N_26409,N_25947,N_25068);
and U26410 (N_26410,N_25077,N_25317);
nor U26411 (N_26411,N_25695,N_25108);
xnor U26412 (N_26412,N_25206,N_25676);
xnor U26413 (N_26413,N_25195,N_25280);
nand U26414 (N_26414,N_25251,N_25076);
nor U26415 (N_26415,N_25688,N_25260);
and U26416 (N_26416,N_25593,N_25565);
xor U26417 (N_26417,N_25683,N_25905);
and U26418 (N_26418,N_25646,N_25710);
nor U26419 (N_26419,N_25118,N_25434);
xnor U26420 (N_26420,N_25943,N_25471);
xor U26421 (N_26421,N_25029,N_25632);
xnor U26422 (N_26422,N_25349,N_25743);
or U26423 (N_26423,N_25680,N_25060);
xnor U26424 (N_26424,N_25595,N_25367);
nor U26425 (N_26425,N_25047,N_25701);
nand U26426 (N_26426,N_25337,N_25949);
or U26427 (N_26427,N_25143,N_25248);
nand U26428 (N_26428,N_25378,N_25168);
nor U26429 (N_26429,N_25171,N_25351);
nor U26430 (N_26430,N_25993,N_25713);
and U26431 (N_26431,N_25959,N_25112);
nand U26432 (N_26432,N_25218,N_25603);
nand U26433 (N_26433,N_25043,N_25622);
or U26434 (N_26434,N_25439,N_25512);
xnor U26435 (N_26435,N_25588,N_25878);
nor U26436 (N_26436,N_25356,N_25389);
nand U26437 (N_26437,N_25056,N_25002);
xnor U26438 (N_26438,N_25621,N_25104);
or U26439 (N_26439,N_25265,N_25755);
nor U26440 (N_26440,N_25554,N_25648);
xor U26441 (N_26441,N_25487,N_25408);
or U26442 (N_26442,N_25845,N_25657);
nor U26443 (N_26443,N_25840,N_25957);
nor U26444 (N_26444,N_25395,N_25034);
nand U26445 (N_26445,N_25498,N_25483);
or U26446 (N_26446,N_25407,N_25200);
xnor U26447 (N_26447,N_25835,N_25003);
xor U26448 (N_26448,N_25933,N_25477);
xnor U26449 (N_26449,N_25083,N_25333);
and U26450 (N_26450,N_25652,N_25312);
xnor U26451 (N_26451,N_25323,N_25787);
xnor U26452 (N_26452,N_25026,N_25732);
or U26453 (N_26453,N_25089,N_25027);
nand U26454 (N_26454,N_25196,N_25852);
or U26455 (N_26455,N_25639,N_25973);
or U26456 (N_26456,N_25720,N_25528);
and U26457 (N_26457,N_25485,N_25425);
xor U26458 (N_26458,N_25377,N_25496);
xor U26459 (N_26459,N_25004,N_25765);
and U26460 (N_26460,N_25490,N_25454);
xor U26461 (N_26461,N_25771,N_25257);
xor U26462 (N_26462,N_25624,N_25985);
and U26463 (N_26463,N_25210,N_25815);
or U26464 (N_26464,N_25803,N_25841);
nand U26465 (N_26465,N_25186,N_25331);
nand U26466 (N_26466,N_25506,N_25397);
xor U26467 (N_26467,N_25583,N_25272);
xor U26468 (N_26468,N_25344,N_25712);
or U26469 (N_26469,N_25670,N_25363);
xor U26470 (N_26470,N_25568,N_25968);
or U26471 (N_26471,N_25794,N_25137);
nor U26472 (N_26472,N_25975,N_25075);
and U26473 (N_26473,N_25937,N_25343);
nor U26474 (N_26474,N_25432,N_25694);
nor U26475 (N_26475,N_25826,N_25521);
and U26476 (N_26476,N_25045,N_25469);
nor U26477 (N_26477,N_25138,N_25948);
or U26478 (N_26478,N_25597,N_25718);
nor U26479 (N_26479,N_25601,N_25169);
and U26480 (N_26480,N_25055,N_25006);
nor U26481 (N_26481,N_25567,N_25245);
and U26482 (N_26482,N_25364,N_25950);
or U26483 (N_26483,N_25054,N_25906);
nor U26484 (N_26484,N_25366,N_25381);
nand U26485 (N_26485,N_25460,N_25673);
or U26486 (N_26486,N_25779,N_25183);
nor U26487 (N_26487,N_25919,N_25598);
and U26488 (N_26488,N_25309,N_25856);
or U26489 (N_26489,N_25922,N_25745);
or U26490 (N_26490,N_25030,N_25269);
xnor U26491 (N_26491,N_25020,N_25879);
nand U26492 (N_26492,N_25818,N_25244);
and U26493 (N_26493,N_25599,N_25067);
and U26494 (N_26494,N_25992,N_25882);
and U26495 (N_26495,N_25238,N_25058);
and U26496 (N_26496,N_25025,N_25069);
and U26497 (N_26497,N_25586,N_25854);
or U26498 (N_26498,N_25306,N_25305);
and U26499 (N_26499,N_25428,N_25285);
or U26500 (N_26500,N_25093,N_25379);
xor U26501 (N_26501,N_25882,N_25251);
or U26502 (N_26502,N_25485,N_25688);
or U26503 (N_26503,N_25589,N_25073);
nand U26504 (N_26504,N_25403,N_25869);
nand U26505 (N_26505,N_25490,N_25401);
or U26506 (N_26506,N_25131,N_25246);
or U26507 (N_26507,N_25585,N_25524);
nor U26508 (N_26508,N_25207,N_25124);
or U26509 (N_26509,N_25422,N_25326);
nand U26510 (N_26510,N_25359,N_25131);
and U26511 (N_26511,N_25421,N_25175);
nor U26512 (N_26512,N_25222,N_25410);
xnor U26513 (N_26513,N_25362,N_25084);
xor U26514 (N_26514,N_25596,N_25121);
or U26515 (N_26515,N_25284,N_25600);
xnor U26516 (N_26516,N_25938,N_25185);
or U26517 (N_26517,N_25556,N_25033);
xnor U26518 (N_26518,N_25098,N_25135);
nor U26519 (N_26519,N_25257,N_25385);
nand U26520 (N_26520,N_25501,N_25502);
xor U26521 (N_26521,N_25236,N_25522);
nand U26522 (N_26522,N_25017,N_25091);
and U26523 (N_26523,N_25902,N_25782);
xnor U26524 (N_26524,N_25788,N_25382);
and U26525 (N_26525,N_25008,N_25531);
nor U26526 (N_26526,N_25748,N_25298);
and U26527 (N_26527,N_25835,N_25439);
xnor U26528 (N_26528,N_25644,N_25960);
nor U26529 (N_26529,N_25689,N_25738);
nor U26530 (N_26530,N_25033,N_25845);
or U26531 (N_26531,N_25159,N_25147);
nor U26532 (N_26532,N_25227,N_25808);
nor U26533 (N_26533,N_25240,N_25853);
xor U26534 (N_26534,N_25912,N_25121);
nor U26535 (N_26535,N_25045,N_25577);
nor U26536 (N_26536,N_25170,N_25347);
and U26537 (N_26537,N_25508,N_25273);
xor U26538 (N_26538,N_25881,N_25625);
xnor U26539 (N_26539,N_25961,N_25812);
or U26540 (N_26540,N_25389,N_25134);
and U26541 (N_26541,N_25988,N_25495);
nor U26542 (N_26542,N_25718,N_25050);
and U26543 (N_26543,N_25615,N_25274);
or U26544 (N_26544,N_25960,N_25066);
nor U26545 (N_26545,N_25232,N_25887);
and U26546 (N_26546,N_25985,N_25831);
nor U26547 (N_26547,N_25590,N_25073);
or U26548 (N_26548,N_25025,N_25223);
nand U26549 (N_26549,N_25612,N_25048);
or U26550 (N_26550,N_25987,N_25790);
xor U26551 (N_26551,N_25715,N_25737);
nand U26552 (N_26552,N_25071,N_25209);
xnor U26553 (N_26553,N_25682,N_25723);
or U26554 (N_26554,N_25654,N_25319);
and U26555 (N_26555,N_25586,N_25622);
nand U26556 (N_26556,N_25939,N_25306);
and U26557 (N_26557,N_25394,N_25280);
nor U26558 (N_26558,N_25265,N_25478);
and U26559 (N_26559,N_25635,N_25728);
nor U26560 (N_26560,N_25050,N_25334);
or U26561 (N_26561,N_25083,N_25468);
or U26562 (N_26562,N_25240,N_25331);
nand U26563 (N_26563,N_25158,N_25446);
xnor U26564 (N_26564,N_25405,N_25533);
xor U26565 (N_26565,N_25065,N_25103);
and U26566 (N_26566,N_25757,N_25420);
nand U26567 (N_26567,N_25130,N_25139);
and U26568 (N_26568,N_25944,N_25902);
and U26569 (N_26569,N_25600,N_25455);
xnor U26570 (N_26570,N_25876,N_25943);
nor U26571 (N_26571,N_25788,N_25585);
xor U26572 (N_26572,N_25309,N_25293);
xor U26573 (N_26573,N_25671,N_25830);
nor U26574 (N_26574,N_25515,N_25609);
xor U26575 (N_26575,N_25237,N_25546);
or U26576 (N_26576,N_25536,N_25355);
nand U26577 (N_26577,N_25299,N_25419);
nand U26578 (N_26578,N_25535,N_25927);
nor U26579 (N_26579,N_25604,N_25404);
xor U26580 (N_26580,N_25480,N_25152);
nand U26581 (N_26581,N_25082,N_25321);
nand U26582 (N_26582,N_25262,N_25439);
or U26583 (N_26583,N_25423,N_25098);
and U26584 (N_26584,N_25139,N_25377);
or U26585 (N_26585,N_25918,N_25158);
nor U26586 (N_26586,N_25586,N_25692);
nand U26587 (N_26587,N_25726,N_25915);
nand U26588 (N_26588,N_25234,N_25821);
or U26589 (N_26589,N_25320,N_25615);
or U26590 (N_26590,N_25739,N_25996);
or U26591 (N_26591,N_25865,N_25369);
and U26592 (N_26592,N_25895,N_25448);
nand U26593 (N_26593,N_25937,N_25491);
nor U26594 (N_26594,N_25005,N_25836);
or U26595 (N_26595,N_25155,N_25557);
or U26596 (N_26596,N_25872,N_25373);
xor U26597 (N_26597,N_25834,N_25706);
xor U26598 (N_26598,N_25270,N_25741);
nand U26599 (N_26599,N_25016,N_25584);
and U26600 (N_26600,N_25736,N_25411);
or U26601 (N_26601,N_25369,N_25463);
nor U26602 (N_26602,N_25584,N_25894);
or U26603 (N_26603,N_25618,N_25066);
nand U26604 (N_26604,N_25579,N_25275);
xor U26605 (N_26605,N_25537,N_25658);
xnor U26606 (N_26606,N_25110,N_25743);
nand U26607 (N_26607,N_25878,N_25413);
xor U26608 (N_26608,N_25902,N_25619);
nor U26609 (N_26609,N_25483,N_25376);
xor U26610 (N_26610,N_25157,N_25746);
nand U26611 (N_26611,N_25318,N_25058);
and U26612 (N_26612,N_25116,N_25409);
nand U26613 (N_26613,N_25083,N_25274);
or U26614 (N_26614,N_25957,N_25459);
nand U26615 (N_26615,N_25079,N_25101);
and U26616 (N_26616,N_25927,N_25944);
or U26617 (N_26617,N_25286,N_25990);
nand U26618 (N_26618,N_25537,N_25683);
xnor U26619 (N_26619,N_25115,N_25257);
and U26620 (N_26620,N_25283,N_25641);
and U26621 (N_26621,N_25809,N_25996);
xor U26622 (N_26622,N_25215,N_25820);
nor U26623 (N_26623,N_25744,N_25007);
nor U26624 (N_26624,N_25326,N_25038);
xor U26625 (N_26625,N_25915,N_25349);
nand U26626 (N_26626,N_25487,N_25024);
or U26627 (N_26627,N_25799,N_25489);
and U26628 (N_26628,N_25542,N_25090);
nand U26629 (N_26629,N_25862,N_25376);
xnor U26630 (N_26630,N_25370,N_25342);
nand U26631 (N_26631,N_25300,N_25864);
and U26632 (N_26632,N_25766,N_25219);
xnor U26633 (N_26633,N_25445,N_25510);
xnor U26634 (N_26634,N_25418,N_25303);
nor U26635 (N_26635,N_25793,N_25876);
nor U26636 (N_26636,N_25678,N_25320);
or U26637 (N_26637,N_25382,N_25062);
xor U26638 (N_26638,N_25224,N_25268);
and U26639 (N_26639,N_25532,N_25426);
nand U26640 (N_26640,N_25898,N_25283);
and U26641 (N_26641,N_25101,N_25306);
nor U26642 (N_26642,N_25615,N_25508);
and U26643 (N_26643,N_25856,N_25054);
nor U26644 (N_26644,N_25452,N_25027);
nand U26645 (N_26645,N_25855,N_25182);
nor U26646 (N_26646,N_25111,N_25190);
nand U26647 (N_26647,N_25846,N_25599);
xnor U26648 (N_26648,N_25178,N_25359);
xor U26649 (N_26649,N_25392,N_25541);
and U26650 (N_26650,N_25593,N_25254);
or U26651 (N_26651,N_25161,N_25687);
and U26652 (N_26652,N_25206,N_25376);
xor U26653 (N_26653,N_25292,N_25274);
nand U26654 (N_26654,N_25918,N_25548);
nor U26655 (N_26655,N_25970,N_25131);
nor U26656 (N_26656,N_25986,N_25510);
nand U26657 (N_26657,N_25276,N_25468);
xor U26658 (N_26658,N_25971,N_25547);
nor U26659 (N_26659,N_25867,N_25702);
xor U26660 (N_26660,N_25617,N_25319);
or U26661 (N_26661,N_25455,N_25499);
or U26662 (N_26662,N_25825,N_25568);
xor U26663 (N_26663,N_25411,N_25385);
or U26664 (N_26664,N_25570,N_25243);
nand U26665 (N_26665,N_25966,N_25534);
or U26666 (N_26666,N_25592,N_25011);
or U26667 (N_26667,N_25187,N_25118);
or U26668 (N_26668,N_25484,N_25324);
xnor U26669 (N_26669,N_25583,N_25750);
or U26670 (N_26670,N_25529,N_25758);
or U26671 (N_26671,N_25935,N_25713);
and U26672 (N_26672,N_25385,N_25288);
xor U26673 (N_26673,N_25400,N_25098);
and U26674 (N_26674,N_25914,N_25394);
nor U26675 (N_26675,N_25505,N_25728);
nand U26676 (N_26676,N_25834,N_25194);
or U26677 (N_26677,N_25690,N_25292);
nand U26678 (N_26678,N_25431,N_25458);
nor U26679 (N_26679,N_25737,N_25866);
nor U26680 (N_26680,N_25536,N_25831);
xnor U26681 (N_26681,N_25444,N_25427);
or U26682 (N_26682,N_25421,N_25231);
nor U26683 (N_26683,N_25022,N_25861);
or U26684 (N_26684,N_25438,N_25377);
or U26685 (N_26685,N_25433,N_25872);
xnor U26686 (N_26686,N_25013,N_25525);
and U26687 (N_26687,N_25480,N_25289);
or U26688 (N_26688,N_25381,N_25300);
nor U26689 (N_26689,N_25451,N_25508);
and U26690 (N_26690,N_25707,N_25904);
or U26691 (N_26691,N_25793,N_25728);
and U26692 (N_26692,N_25764,N_25042);
or U26693 (N_26693,N_25102,N_25549);
nor U26694 (N_26694,N_25242,N_25315);
and U26695 (N_26695,N_25768,N_25568);
or U26696 (N_26696,N_25480,N_25789);
xor U26697 (N_26697,N_25316,N_25800);
xor U26698 (N_26698,N_25442,N_25178);
nor U26699 (N_26699,N_25873,N_25256);
nor U26700 (N_26700,N_25962,N_25250);
nand U26701 (N_26701,N_25542,N_25294);
nor U26702 (N_26702,N_25283,N_25307);
and U26703 (N_26703,N_25800,N_25191);
nand U26704 (N_26704,N_25191,N_25344);
nor U26705 (N_26705,N_25453,N_25069);
nor U26706 (N_26706,N_25189,N_25651);
and U26707 (N_26707,N_25543,N_25104);
nor U26708 (N_26708,N_25093,N_25556);
xnor U26709 (N_26709,N_25594,N_25513);
or U26710 (N_26710,N_25925,N_25090);
nand U26711 (N_26711,N_25309,N_25588);
or U26712 (N_26712,N_25311,N_25827);
xor U26713 (N_26713,N_25557,N_25585);
xor U26714 (N_26714,N_25860,N_25055);
or U26715 (N_26715,N_25787,N_25711);
xor U26716 (N_26716,N_25511,N_25607);
nor U26717 (N_26717,N_25177,N_25946);
and U26718 (N_26718,N_25789,N_25095);
and U26719 (N_26719,N_25338,N_25505);
and U26720 (N_26720,N_25192,N_25437);
or U26721 (N_26721,N_25189,N_25650);
xnor U26722 (N_26722,N_25142,N_25061);
xor U26723 (N_26723,N_25570,N_25405);
nand U26724 (N_26724,N_25912,N_25086);
and U26725 (N_26725,N_25481,N_25112);
nor U26726 (N_26726,N_25969,N_25929);
nand U26727 (N_26727,N_25644,N_25776);
and U26728 (N_26728,N_25489,N_25393);
xnor U26729 (N_26729,N_25603,N_25354);
and U26730 (N_26730,N_25932,N_25749);
and U26731 (N_26731,N_25559,N_25384);
nand U26732 (N_26732,N_25385,N_25392);
xnor U26733 (N_26733,N_25937,N_25490);
nand U26734 (N_26734,N_25696,N_25400);
nor U26735 (N_26735,N_25814,N_25740);
nor U26736 (N_26736,N_25143,N_25316);
or U26737 (N_26737,N_25909,N_25197);
nor U26738 (N_26738,N_25699,N_25182);
nand U26739 (N_26739,N_25082,N_25460);
and U26740 (N_26740,N_25590,N_25970);
and U26741 (N_26741,N_25977,N_25245);
nand U26742 (N_26742,N_25520,N_25336);
nand U26743 (N_26743,N_25806,N_25175);
or U26744 (N_26744,N_25529,N_25954);
and U26745 (N_26745,N_25510,N_25128);
xor U26746 (N_26746,N_25278,N_25130);
or U26747 (N_26747,N_25723,N_25199);
nand U26748 (N_26748,N_25286,N_25312);
nand U26749 (N_26749,N_25911,N_25139);
xor U26750 (N_26750,N_25662,N_25449);
xor U26751 (N_26751,N_25657,N_25510);
and U26752 (N_26752,N_25092,N_25425);
nand U26753 (N_26753,N_25069,N_25169);
or U26754 (N_26754,N_25604,N_25680);
or U26755 (N_26755,N_25632,N_25547);
nor U26756 (N_26756,N_25790,N_25227);
xor U26757 (N_26757,N_25982,N_25827);
or U26758 (N_26758,N_25955,N_25301);
or U26759 (N_26759,N_25492,N_25971);
nand U26760 (N_26760,N_25860,N_25136);
xor U26761 (N_26761,N_25899,N_25365);
nor U26762 (N_26762,N_25239,N_25286);
and U26763 (N_26763,N_25945,N_25473);
nand U26764 (N_26764,N_25054,N_25900);
and U26765 (N_26765,N_25447,N_25550);
nor U26766 (N_26766,N_25288,N_25600);
nor U26767 (N_26767,N_25162,N_25502);
nor U26768 (N_26768,N_25952,N_25400);
nand U26769 (N_26769,N_25171,N_25314);
or U26770 (N_26770,N_25051,N_25677);
nor U26771 (N_26771,N_25532,N_25749);
or U26772 (N_26772,N_25485,N_25729);
nor U26773 (N_26773,N_25334,N_25695);
xnor U26774 (N_26774,N_25311,N_25465);
xor U26775 (N_26775,N_25556,N_25577);
or U26776 (N_26776,N_25081,N_25475);
and U26777 (N_26777,N_25931,N_25092);
or U26778 (N_26778,N_25266,N_25579);
nor U26779 (N_26779,N_25107,N_25476);
xnor U26780 (N_26780,N_25546,N_25291);
and U26781 (N_26781,N_25316,N_25289);
nand U26782 (N_26782,N_25414,N_25673);
and U26783 (N_26783,N_25634,N_25851);
nor U26784 (N_26784,N_25471,N_25579);
nor U26785 (N_26785,N_25766,N_25094);
or U26786 (N_26786,N_25041,N_25072);
xor U26787 (N_26787,N_25344,N_25132);
and U26788 (N_26788,N_25554,N_25497);
and U26789 (N_26789,N_25373,N_25360);
and U26790 (N_26790,N_25244,N_25293);
and U26791 (N_26791,N_25155,N_25036);
and U26792 (N_26792,N_25367,N_25044);
and U26793 (N_26793,N_25759,N_25256);
or U26794 (N_26794,N_25904,N_25445);
or U26795 (N_26795,N_25579,N_25469);
or U26796 (N_26796,N_25603,N_25334);
nand U26797 (N_26797,N_25658,N_25076);
and U26798 (N_26798,N_25675,N_25846);
and U26799 (N_26799,N_25386,N_25005);
and U26800 (N_26800,N_25239,N_25802);
and U26801 (N_26801,N_25601,N_25963);
xor U26802 (N_26802,N_25169,N_25967);
and U26803 (N_26803,N_25748,N_25889);
nor U26804 (N_26804,N_25231,N_25159);
nand U26805 (N_26805,N_25390,N_25945);
nor U26806 (N_26806,N_25880,N_25652);
xor U26807 (N_26807,N_25041,N_25172);
or U26808 (N_26808,N_25879,N_25959);
nor U26809 (N_26809,N_25370,N_25004);
nor U26810 (N_26810,N_25745,N_25856);
xnor U26811 (N_26811,N_25660,N_25903);
or U26812 (N_26812,N_25840,N_25551);
nand U26813 (N_26813,N_25534,N_25562);
and U26814 (N_26814,N_25483,N_25815);
xor U26815 (N_26815,N_25405,N_25754);
xor U26816 (N_26816,N_25822,N_25215);
nor U26817 (N_26817,N_25304,N_25991);
xnor U26818 (N_26818,N_25365,N_25062);
and U26819 (N_26819,N_25078,N_25703);
or U26820 (N_26820,N_25626,N_25144);
and U26821 (N_26821,N_25550,N_25870);
and U26822 (N_26822,N_25696,N_25683);
xor U26823 (N_26823,N_25931,N_25924);
nor U26824 (N_26824,N_25594,N_25657);
and U26825 (N_26825,N_25761,N_25270);
and U26826 (N_26826,N_25859,N_25122);
and U26827 (N_26827,N_25962,N_25616);
nand U26828 (N_26828,N_25185,N_25181);
nand U26829 (N_26829,N_25298,N_25186);
nand U26830 (N_26830,N_25491,N_25495);
nor U26831 (N_26831,N_25652,N_25675);
and U26832 (N_26832,N_25251,N_25903);
and U26833 (N_26833,N_25207,N_25290);
nand U26834 (N_26834,N_25773,N_25865);
nor U26835 (N_26835,N_25723,N_25419);
nand U26836 (N_26836,N_25614,N_25763);
or U26837 (N_26837,N_25743,N_25043);
nor U26838 (N_26838,N_25741,N_25640);
and U26839 (N_26839,N_25734,N_25453);
xor U26840 (N_26840,N_25066,N_25896);
and U26841 (N_26841,N_25535,N_25698);
nor U26842 (N_26842,N_25336,N_25594);
xor U26843 (N_26843,N_25109,N_25334);
nor U26844 (N_26844,N_25741,N_25844);
xnor U26845 (N_26845,N_25644,N_25798);
and U26846 (N_26846,N_25821,N_25804);
nor U26847 (N_26847,N_25674,N_25148);
and U26848 (N_26848,N_25991,N_25635);
nor U26849 (N_26849,N_25988,N_25547);
nor U26850 (N_26850,N_25492,N_25375);
or U26851 (N_26851,N_25918,N_25221);
nor U26852 (N_26852,N_25926,N_25948);
or U26853 (N_26853,N_25908,N_25587);
nor U26854 (N_26854,N_25691,N_25003);
nor U26855 (N_26855,N_25621,N_25663);
nor U26856 (N_26856,N_25325,N_25319);
nor U26857 (N_26857,N_25193,N_25883);
nor U26858 (N_26858,N_25843,N_25578);
nand U26859 (N_26859,N_25564,N_25929);
xnor U26860 (N_26860,N_25150,N_25500);
xor U26861 (N_26861,N_25900,N_25606);
nor U26862 (N_26862,N_25234,N_25108);
and U26863 (N_26863,N_25311,N_25846);
and U26864 (N_26864,N_25419,N_25179);
xor U26865 (N_26865,N_25907,N_25083);
or U26866 (N_26866,N_25093,N_25030);
and U26867 (N_26867,N_25466,N_25202);
nand U26868 (N_26868,N_25803,N_25457);
xor U26869 (N_26869,N_25747,N_25529);
or U26870 (N_26870,N_25057,N_25095);
xnor U26871 (N_26871,N_25951,N_25810);
or U26872 (N_26872,N_25304,N_25019);
or U26873 (N_26873,N_25216,N_25608);
nor U26874 (N_26874,N_25079,N_25290);
nor U26875 (N_26875,N_25284,N_25343);
nor U26876 (N_26876,N_25150,N_25876);
nor U26877 (N_26877,N_25732,N_25408);
nand U26878 (N_26878,N_25015,N_25423);
or U26879 (N_26879,N_25972,N_25821);
or U26880 (N_26880,N_25679,N_25134);
and U26881 (N_26881,N_25025,N_25110);
xnor U26882 (N_26882,N_25962,N_25550);
xnor U26883 (N_26883,N_25770,N_25982);
nor U26884 (N_26884,N_25844,N_25293);
xnor U26885 (N_26885,N_25033,N_25115);
or U26886 (N_26886,N_25035,N_25827);
nand U26887 (N_26887,N_25210,N_25591);
or U26888 (N_26888,N_25217,N_25977);
xnor U26889 (N_26889,N_25896,N_25432);
nor U26890 (N_26890,N_25711,N_25765);
xnor U26891 (N_26891,N_25777,N_25600);
or U26892 (N_26892,N_25469,N_25038);
nor U26893 (N_26893,N_25535,N_25352);
nor U26894 (N_26894,N_25786,N_25101);
and U26895 (N_26895,N_25031,N_25569);
nand U26896 (N_26896,N_25457,N_25536);
nand U26897 (N_26897,N_25951,N_25305);
or U26898 (N_26898,N_25329,N_25759);
or U26899 (N_26899,N_25336,N_25854);
xnor U26900 (N_26900,N_25649,N_25603);
nor U26901 (N_26901,N_25394,N_25702);
nand U26902 (N_26902,N_25383,N_25243);
nor U26903 (N_26903,N_25661,N_25834);
and U26904 (N_26904,N_25676,N_25738);
or U26905 (N_26905,N_25518,N_25922);
and U26906 (N_26906,N_25697,N_25146);
xor U26907 (N_26907,N_25059,N_25594);
and U26908 (N_26908,N_25128,N_25429);
and U26909 (N_26909,N_25476,N_25010);
and U26910 (N_26910,N_25087,N_25748);
nor U26911 (N_26911,N_25030,N_25541);
or U26912 (N_26912,N_25978,N_25564);
xnor U26913 (N_26913,N_25298,N_25174);
nand U26914 (N_26914,N_25948,N_25572);
or U26915 (N_26915,N_25180,N_25964);
or U26916 (N_26916,N_25493,N_25477);
nand U26917 (N_26917,N_25085,N_25580);
and U26918 (N_26918,N_25923,N_25323);
xnor U26919 (N_26919,N_25259,N_25580);
nand U26920 (N_26920,N_25157,N_25477);
nor U26921 (N_26921,N_25594,N_25629);
or U26922 (N_26922,N_25991,N_25327);
or U26923 (N_26923,N_25370,N_25108);
or U26924 (N_26924,N_25975,N_25903);
nand U26925 (N_26925,N_25674,N_25554);
or U26926 (N_26926,N_25295,N_25777);
nor U26927 (N_26927,N_25682,N_25480);
xor U26928 (N_26928,N_25463,N_25032);
nand U26929 (N_26929,N_25786,N_25087);
xnor U26930 (N_26930,N_25110,N_25392);
nand U26931 (N_26931,N_25855,N_25986);
xnor U26932 (N_26932,N_25442,N_25208);
or U26933 (N_26933,N_25012,N_25474);
and U26934 (N_26934,N_25395,N_25163);
nor U26935 (N_26935,N_25732,N_25461);
and U26936 (N_26936,N_25358,N_25487);
nor U26937 (N_26937,N_25569,N_25523);
xnor U26938 (N_26938,N_25596,N_25260);
or U26939 (N_26939,N_25065,N_25885);
or U26940 (N_26940,N_25135,N_25495);
or U26941 (N_26941,N_25903,N_25643);
and U26942 (N_26942,N_25956,N_25039);
and U26943 (N_26943,N_25224,N_25338);
xor U26944 (N_26944,N_25442,N_25021);
xor U26945 (N_26945,N_25167,N_25925);
or U26946 (N_26946,N_25045,N_25274);
xor U26947 (N_26947,N_25721,N_25281);
or U26948 (N_26948,N_25344,N_25877);
or U26949 (N_26949,N_25446,N_25147);
nor U26950 (N_26950,N_25675,N_25796);
or U26951 (N_26951,N_25355,N_25918);
nor U26952 (N_26952,N_25867,N_25943);
xor U26953 (N_26953,N_25232,N_25182);
and U26954 (N_26954,N_25823,N_25480);
or U26955 (N_26955,N_25616,N_25865);
xnor U26956 (N_26956,N_25404,N_25293);
xnor U26957 (N_26957,N_25901,N_25352);
or U26958 (N_26958,N_25697,N_25500);
xnor U26959 (N_26959,N_25789,N_25720);
and U26960 (N_26960,N_25528,N_25343);
xnor U26961 (N_26961,N_25685,N_25177);
and U26962 (N_26962,N_25505,N_25053);
nand U26963 (N_26963,N_25381,N_25946);
and U26964 (N_26964,N_25517,N_25107);
nand U26965 (N_26965,N_25004,N_25691);
or U26966 (N_26966,N_25917,N_25007);
nand U26967 (N_26967,N_25102,N_25279);
or U26968 (N_26968,N_25637,N_25349);
and U26969 (N_26969,N_25635,N_25136);
nor U26970 (N_26970,N_25769,N_25493);
and U26971 (N_26971,N_25712,N_25614);
nor U26972 (N_26972,N_25731,N_25088);
or U26973 (N_26973,N_25380,N_25322);
nand U26974 (N_26974,N_25269,N_25807);
and U26975 (N_26975,N_25116,N_25606);
nand U26976 (N_26976,N_25104,N_25083);
nor U26977 (N_26977,N_25205,N_25730);
or U26978 (N_26978,N_25803,N_25986);
and U26979 (N_26979,N_25772,N_25744);
nand U26980 (N_26980,N_25034,N_25406);
nand U26981 (N_26981,N_25153,N_25736);
and U26982 (N_26982,N_25388,N_25411);
nor U26983 (N_26983,N_25669,N_25887);
nor U26984 (N_26984,N_25185,N_25490);
nor U26985 (N_26985,N_25742,N_25187);
nor U26986 (N_26986,N_25472,N_25891);
xor U26987 (N_26987,N_25014,N_25058);
or U26988 (N_26988,N_25196,N_25619);
or U26989 (N_26989,N_25580,N_25357);
xnor U26990 (N_26990,N_25237,N_25019);
xor U26991 (N_26991,N_25306,N_25105);
nand U26992 (N_26992,N_25164,N_25064);
nand U26993 (N_26993,N_25245,N_25438);
nand U26994 (N_26994,N_25013,N_25289);
xnor U26995 (N_26995,N_25780,N_25805);
and U26996 (N_26996,N_25703,N_25805);
and U26997 (N_26997,N_25791,N_25099);
xor U26998 (N_26998,N_25844,N_25512);
nor U26999 (N_26999,N_25219,N_25725);
and U27000 (N_27000,N_26009,N_26321);
xnor U27001 (N_27001,N_26720,N_26690);
nor U27002 (N_27002,N_26116,N_26161);
nand U27003 (N_27003,N_26825,N_26264);
and U27004 (N_27004,N_26565,N_26668);
nand U27005 (N_27005,N_26079,N_26258);
xnor U27006 (N_27006,N_26412,N_26142);
xor U27007 (N_27007,N_26569,N_26910);
and U27008 (N_27008,N_26734,N_26317);
and U27009 (N_27009,N_26121,N_26632);
xnor U27010 (N_27010,N_26562,N_26631);
nand U27011 (N_27011,N_26297,N_26883);
nand U27012 (N_27012,N_26558,N_26556);
nand U27013 (N_27013,N_26078,N_26605);
nand U27014 (N_27014,N_26822,N_26314);
nor U27015 (N_27015,N_26439,N_26359);
or U27016 (N_27016,N_26505,N_26405);
and U27017 (N_27017,N_26953,N_26552);
nor U27018 (N_27018,N_26188,N_26323);
nand U27019 (N_27019,N_26335,N_26561);
nand U27020 (N_27020,N_26383,N_26364);
and U27021 (N_27021,N_26222,N_26463);
nand U27022 (N_27022,N_26326,N_26267);
or U27023 (N_27023,N_26378,N_26217);
and U27024 (N_27024,N_26170,N_26986);
or U27025 (N_27025,N_26376,N_26890);
or U27026 (N_27026,N_26528,N_26905);
and U27027 (N_27027,N_26177,N_26346);
nand U27028 (N_27028,N_26773,N_26752);
xor U27029 (N_27029,N_26760,N_26785);
or U27030 (N_27030,N_26058,N_26714);
or U27031 (N_27031,N_26237,N_26725);
and U27032 (N_27032,N_26347,N_26820);
nand U27033 (N_27033,N_26497,N_26526);
or U27034 (N_27034,N_26319,N_26848);
nand U27035 (N_27035,N_26574,N_26134);
nand U27036 (N_27036,N_26782,N_26304);
or U27037 (N_27037,N_26454,N_26792);
and U27038 (N_27038,N_26841,N_26763);
xnor U27039 (N_27039,N_26008,N_26533);
xnor U27040 (N_27040,N_26824,N_26738);
nor U27041 (N_27041,N_26028,N_26973);
and U27042 (N_27042,N_26193,N_26387);
or U27043 (N_27043,N_26292,N_26580);
and U27044 (N_27044,N_26621,N_26508);
nand U27045 (N_27045,N_26473,N_26642);
nand U27046 (N_27046,N_26732,N_26559);
xnor U27047 (N_27047,N_26160,N_26288);
or U27048 (N_27048,N_26955,N_26420);
nand U27049 (N_27049,N_26514,N_26354);
and U27050 (N_27050,N_26850,N_26675);
or U27051 (N_27051,N_26012,N_26369);
nand U27052 (N_27052,N_26649,N_26827);
nand U27053 (N_27053,N_26650,N_26742);
or U27054 (N_27054,N_26608,N_26902);
nand U27055 (N_27055,N_26694,N_26224);
or U27056 (N_27056,N_26370,N_26909);
nand U27057 (N_27057,N_26598,N_26262);
nor U27058 (N_27058,N_26402,N_26298);
xor U27059 (N_27059,N_26882,N_26316);
xnor U27060 (N_27060,N_26372,N_26894);
xor U27061 (N_27061,N_26733,N_26399);
and U27062 (N_27062,N_26787,N_26933);
nor U27063 (N_27063,N_26010,N_26845);
and U27064 (N_27064,N_26639,N_26547);
nand U27065 (N_27065,N_26174,N_26931);
or U27066 (N_27066,N_26736,N_26455);
or U27067 (N_27067,N_26748,N_26667);
and U27068 (N_27068,N_26087,N_26837);
nor U27069 (N_27069,N_26230,N_26684);
nand U27070 (N_27070,N_26591,N_26430);
or U27071 (N_27071,N_26476,N_26281);
nor U27072 (N_27072,N_26500,N_26685);
and U27073 (N_27073,N_26940,N_26949);
nor U27074 (N_27074,N_26807,N_26524);
nor U27075 (N_27075,N_26770,N_26974);
and U27076 (N_27076,N_26089,N_26941);
nor U27077 (N_27077,N_26020,N_26828);
or U27078 (N_27078,N_26203,N_26265);
or U27079 (N_27079,N_26998,N_26209);
or U27080 (N_27080,N_26799,N_26254);
and U27081 (N_27081,N_26120,N_26227);
nor U27082 (N_27082,N_26112,N_26554);
nor U27083 (N_27083,N_26865,N_26466);
xor U27084 (N_27084,N_26155,N_26576);
nand U27085 (N_27085,N_26681,N_26417);
or U27086 (N_27086,N_26641,N_26067);
xor U27087 (N_27087,N_26935,N_26852);
nand U27088 (N_27088,N_26153,N_26891);
xnor U27089 (N_27089,N_26895,N_26475);
nor U27090 (N_27090,N_26717,N_26866);
nand U27091 (N_27091,N_26447,N_26494);
xnor U27092 (N_27092,N_26654,N_26702);
nor U27093 (N_27093,N_26181,N_26912);
xnor U27094 (N_27094,N_26779,N_26186);
nor U27095 (N_27095,N_26234,N_26406);
xor U27096 (N_27096,N_26031,N_26017);
and U27097 (N_27097,N_26421,N_26219);
and U27098 (N_27098,N_26629,N_26783);
xnor U27099 (N_27099,N_26429,N_26056);
and U27100 (N_27100,N_26626,N_26126);
or U27101 (N_27101,N_26744,N_26542);
xor U27102 (N_27102,N_26696,N_26386);
nand U27103 (N_27103,N_26854,N_26979);
xor U27104 (N_27104,N_26583,N_26794);
nand U27105 (N_27105,N_26983,N_26469);
xor U27106 (N_27106,N_26778,N_26464);
and U27107 (N_27107,N_26391,N_26585);
and U27108 (N_27108,N_26726,N_26210);
and U27109 (N_27109,N_26957,N_26024);
or U27110 (N_27110,N_26432,N_26970);
xnor U27111 (N_27111,N_26047,N_26567);
nand U27112 (N_27112,N_26964,N_26903);
nor U27113 (N_27113,N_26228,N_26414);
xnor U27114 (N_27114,N_26252,N_26590);
or U27115 (N_27115,N_26327,N_26568);
xnor U27116 (N_27116,N_26039,N_26698);
and U27117 (N_27117,N_26269,N_26946);
nor U27118 (N_27118,N_26603,N_26754);
nand U27119 (N_27119,N_26384,N_26498);
or U27120 (N_27120,N_26158,N_26448);
or U27121 (N_27121,N_26647,N_26353);
and U27122 (N_27122,N_26867,N_26460);
xnor U27123 (N_27123,N_26148,N_26208);
xnor U27124 (N_27124,N_26456,N_26990);
nor U27125 (N_27125,N_26495,N_26259);
and U27126 (N_27126,N_26939,N_26016);
or U27127 (N_27127,N_26637,N_26652);
nor U27128 (N_27128,N_26994,N_26442);
nor U27129 (N_27129,N_26881,N_26572);
and U27130 (N_27130,N_26768,N_26861);
nand U27131 (N_27131,N_26747,N_26722);
and U27132 (N_27132,N_26833,N_26176);
xor U27133 (N_27133,N_26507,N_26504);
xor U27134 (N_27134,N_26844,N_26634);
and U27135 (N_27135,N_26408,N_26049);
and U27136 (N_27136,N_26436,N_26446);
and U27137 (N_27137,N_26821,N_26988);
nand U27138 (N_27138,N_26481,N_26543);
or U27139 (N_27139,N_26285,N_26184);
nor U27140 (N_27140,N_26503,N_26266);
nand U27141 (N_27141,N_26200,N_26474);
xor U27142 (N_27142,N_26048,N_26309);
nand U27143 (N_27143,N_26109,N_26706);
nand U27144 (N_27144,N_26589,N_26401);
xnor U27145 (N_27145,N_26615,N_26145);
and U27146 (N_27146,N_26814,N_26862);
nor U27147 (N_27147,N_26606,N_26943);
and U27148 (N_27148,N_26357,N_26594);
nand U27149 (N_27149,N_26462,N_26633);
and U27150 (N_27150,N_26362,N_26512);
and U27151 (N_27151,N_26759,N_26137);
nand U27152 (N_27152,N_26331,N_26766);
or U27153 (N_27153,N_26965,N_26172);
nand U27154 (N_27154,N_26597,N_26315);
nand U27155 (N_27155,N_26651,N_26645);
xor U27156 (N_27156,N_26046,N_26179);
or U27157 (N_27157,N_26437,N_26914);
xnor U27158 (N_27158,N_26936,N_26804);
nor U27159 (N_27159,N_26966,N_26884);
and U27160 (N_27160,N_26846,N_26496);
or U27161 (N_27161,N_26805,N_26104);
xnor U27162 (N_27162,N_26586,N_26027);
or U27163 (N_27163,N_26084,N_26727);
and U27164 (N_27164,N_26545,N_26578);
nand U27165 (N_27165,N_26418,N_26088);
and U27166 (N_27166,N_26484,N_26344);
nor U27167 (N_27167,N_26246,N_26431);
nor U27168 (N_27168,N_26416,N_26777);
or U27169 (N_27169,N_26043,N_26789);
and U27170 (N_27170,N_26810,N_26919);
nand U27171 (N_27171,N_26922,N_26893);
xnor U27172 (N_27172,N_26857,N_26610);
xnor U27173 (N_27173,N_26006,N_26013);
nor U27174 (N_27174,N_26907,N_26878);
and U27175 (N_27175,N_26870,N_26037);
nand U27176 (N_27176,N_26600,N_26993);
and U27177 (N_27177,N_26581,N_26616);
nor U27178 (N_27178,N_26715,N_26124);
nor U27179 (N_27179,N_26368,N_26026);
or U27180 (N_27180,N_26959,N_26187);
nor U27181 (N_27181,N_26938,N_26075);
nand U27182 (N_27182,N_26493,N_26539);
nand U27183 (N_27183,N_26934,N_26519);
and U27184 (N_27184,N_26040,N_26366);
and U27185 (N_27185,N_26871,N_26635);
or U27186 (N_27186,N_26716,N_26280);
nor U27187 (N_27187,N_26025,N_26180);
or U27188 (N_27188,N_26521,N_26233);
nor U27189 (N_27189,N_26450,N_26070);
nand U27190 (N_27190,N_26544,N_26095);
nand U27191 (N_27191,N_26275,N_26441);
or U27192 (N_27192,N_26995,N_26711);
nand U27193 (N_27193,N_26348,N_26057);
nand U27194 (N_27194,N_26197,N_26588);
xnor U27195 (N_27195,N_26488,N_26900);
xor U27196 (N_27196,N_26394,N_26425);
xnor U27197 (N_27197,N_26196,N_26643);
nand U27198 (N_27198,N_26092,N_26669);
or U27199 (N_27199,N_26303,N_26113);
xnor U27200 (N_27200,N_26735,N_26549);
or U27201 (N_27201,N_26007,N_26619);
and U27202 (N_27202,N_26532,N_26125);
nand U27203 (N_27203,N_26864,N_26751);
nand U27204 (N_27204,N_26205,N_26676);
xnor U27205 (N_27205,N_26819,N_26860);
xor U27206 (N_27206,N_26243,N_26816);
nor U27207 (N_27207,N_26062,N_26198);
or U27208 (N_27208,N_26687,N_26413);
or U27209 (N_27209,N_26299,N_26511);
xnor U27210 (N_27210,N_26700,N_26740);
xnor U27211 (N_27211,N_26628,N_26035);
and U27212 (N_27212,N_26163,N_26847);
nor U27213 (N_27213,N_26226,N_26108);
and U27214 (N_27214,N_26086,N_26482);
nor U27215 (N_27215,N_26168,N_26843);
nand U27216 (N_27216,N_26999,N_26015);
nor U27217 (N_27217,N_26081,N_26548);
nor U27218 (N_27218,N_26958,N_26245);
or U27219 (N_27219,N_26036,N_26072);
nor U27220 (N_27220,N_26885,N_26232);
nor U27221 (N_27221,N_26529,N_26167);
and U27222 (N_27222,N_26815,N_26584);
or U27223 (N_27223,N_26294,N_26123);
nand U27224 (N_27224,N_26718,N_26987);
nor U27225 (N_27225,N_26131,N_26422);
and U27226 (N_27226,N_26874,N_26771);
nor U27227 (N_27227,N_26730,N_26756);
or U27228 (N_27228,N_26518,N_26927);
xnor U27229 (N_27229,N_26468,N_26665);
xnor U27230 (N_27230,N_26011,N_26060);
or U27231 (N_27231,N_26896,N_26138);
nor U27232 (N_27232,N_26330,N_26282);
nand U27233 (N_27233,N_26945,N_26229);
nand U27234 (N_27234,N_26788,N_26969);
nor U27235 (N_27235,N_26587,N_26832);
or U27236 (N_27236,N_26930,N_26546);
nand U27237 (N_27237,N_26065,N_26272);
and U27238 (N_27238,N_26293,N_26873);
nand U27239 (N_27239,N_26215,N_26459);
and U27240 (N_27240,N_26212,N_26477);
nand U27241 (N_27241,N_26944,N_26300);
nand U27242 (N_27242,N_26664,N_26090);
or U27243 (N_27243,N_26061,N_26679);
xnor U27244 (N_27244,N_26674,N_26954);
nor U27245 (N_27245,N_26886,N_26758);
or U27246 (N_27246,N_26424,N_26244);
xor U27247 (N_27247,N_26165,N_26762);
or U27248 (N_27248,N_26968,N_26403);
or U27249 (N_27249,N_26753,N_26991);
nand U27250 (N_27250,N_26271,N_26522);
nand U27251 (N_27251,N_26169,N_26178);
xor U27252 (N_27252,N_26284,N_26786);
nor U27253 (N_27253,N_26797,N_26162);
nor U27254 (N_27254,N_26680,N_26053);
xor U27255 (N_27255,N_26301,N_26618);
or U27256 (N_27256,N_26076,N_26579);
nand U27257 (N_27257,N_26851,N_26573);
xor U27258 (N_27258,N_26948,N_26472);
or U27259 (N_27259,N_26918,N_26305);
or U27260 (N_27260,N_26333,N_26361);
nand U27261 (N_27261,N_26336,N_26152);
xnor U27262 (N_27262,N_26739,N_26743);
nand U27263 (N_27263,N_26666,N_26063);
and U27264 (N_27264,N_26071,N_26921);
or U27265 (N_27265,N_26302,N_26980);
xor U27266 (N_27266,N_26901,N_26709);
or U27267 (N_27267,N_26367,N_26154);
nand U27268 (N_27268,N_26373,N_26707);
nor U27269 (N_27269,N_26889,N_26708);
nor U27270 (N_27270,N_26055,N_26656);
and U27271 (N_27271,N_26192,N_26150);
or U27272 (N_27272,N_26310,N_26638);
and U27273 (N_27273,N_26728,N_26555);
and U27274 (N_27274,N_26961,N_26239);
and U27275 (N_27275,N_26478,N_26798);
nand U27276 (N_27276,N_26139,N_26712);
nand U27277 (N_27277,N_26531,N_26924);
and U27278 (N_27278,N_26166,N_26623);
or U27279 (N_27279,N_26206,N_26906);
nand U27280 (N_27280,N_26465,N_26276);
nand U27281 (N_27281,N_26640,N_26801);
nor U27282 (N_27282,N_26451,N_26863);
and U27283 (N_27283,N_26657,N_26840);
nor U27284 (N_27284,N_26951,N_26390);
nor U27285 (N_27285,N_26932,N_26345);
nand U27286 (N_27286,N_26273,N_26073);
nor U27287 (N_27287,N_26617,N_26741);
or U27288 (N_27288,N_26171,N_26577);
or U27289 (N_27289,N_26677,N_26682);
and U27290 (N_27290,N_26207,N_26263);
or U27291 (N_27291,N_26869,N_26050);
and U27292 (N_27292,N_26253,N_26520);
nor U27293 (N_27293,N_26256,N_26411);
nand U27294 (N_27294,N_26795,N_26082);
nor U27295 (N_27295,N_26202,N_26622);
and U27296 (N_27296,N_26975,N_26996);
and U27297 (N_27297,N_26343,N_26080);
or U27298 (N_27298,N_26328,N_26978);
nor U27299 (N_27299,N_26612,N_26018);
nor U27300 (N_27300,N_26251,N_26913);
or U27301 (N_27301,N_26277,N_26388);
or U27302 (N_27302,N_26693,N_26382);
xor U27303 (N_27303,N_26704,N_26000);
or U27304 (N_27304,N_26829,N_26705);
xor U27305 (N_27305,N_26400,N_26839);
xnor U27306 (N_27306,N_26102,N_26904);
xnor U27307 (N_27307,N_26673,N_26099);
nor U27308 (N_27308,N_26757,N_26611);
and U27309 (N_27309,N_26019,N_26005);
and U27310 (N_27310,N_26755,N_26159);
or U27311 (N_27311,N_26793,N_26540);
nor U27312 (N_27312,N_26775,N_26492);
and U27313 (N_27313,N_26190,N_26501);
or U27314 (N_27314,N_26689,N_26032);
and U27315 (N_27315,N_26774,N_26853);
xor U27316 (N_27316,N_26950,N_26128);
nor U27317 (N_27317,N_26340,N_26054);
or U27318 (N_27318,N_26452,N_26404);
nand U27319 (N_27319,N_26042,N_26997);
or U27320 (N_27320,N_26658,N_26613);
or U27321 (N_27321,N_26593,N_26185);
nor U27322 (N_27322,N_26033,N_26453);
nand U27323 (N_27323,N_26249,N_26467);
xnor U27324 (N_27324,N_26211,N_26296);
nand U27325 (N_27325,N_26068,N_26686);
or U27326 (N_27326,N_26776,N_26097);
xnor U27327 (N_27327,N_26074,N_26745);
nor U27328 (N_27328,N_26146,N_26238);
or U27329 (N_27329,N_26445,N_26575);
or U27330 (N_27330,N_26051,N_26103);
xnor U27331 (N_27331,N_26337,N_26213);
nor U27332 (N_27332,N_26371,N_26536);
nand U27333 (N_27333,N_26570,N_26014);
and U27334 (N_27334,N_26858,N_26509);
and U27335 (N_27335,N_26261,N_26077);
and U27336 (N_27336,N_26250,N_26127);
xor U27337 (N_27337,N_26241,N_26044);
nor U27338 (N_27338,N_26338,N_26942);
and U27339 (N_27339,N_26115,N_26678);
or U27340 (N_27340,N_26802,N_26719);
nand U27341 (N_27341,N_26699,N_26479);
xnor U27342 (N_27342,N_26085,N_26352);
and U27343 (N_27343,N_26566,N_26393);
or U27344 (N_27344,N_26899,N_26490);
nor U27345 (N_27345,N_26183,N_26517);
and U27346 (N_27346,N_26737,N_26887);
nor U27347 (N_27347,N_26397,N_26435);
and U27348 (N_27348,N_26510,N_26780);
nand U27349 (N_27349,N_26892,N_26984);
and U27350 (N_27350,N_26438,N_26796);
nand U27351 (N_27351,N_26363,N_26662);
nor U27352 (N_27352,N_26423,N_26981);
nand U27353 (N_27353,N_26697,N_26557);
and U27354 (N_27354,N_26872,N_26398);
and U27355 (N_27355,N_26750,N_26114);
nor U27356 (N_27356,N_26790,N_26977);
nand U27357 (N_27357,N_26917,N_26307);
nor U27358 (N_27358,N_26879,N_26415);
and U27359 (N_27359,N_26132,N_26855);
nor U27360 (N_27360,N_26655,N_26800);
or U27361 (N_27361,N_26604,N_26749);
xnor U27362 (N_27362,N_26449,N_26989);
and U27363 (N_27363,N_26897,N_26784);
and U27364 (N_27364,N_26537,N_26247);
nand U27365 (N_27365,N_26444,N_26880);
nor U27366 (N_27366,N_26646,N_26486);
xor U27367 (N_27367,N_26868,N_26260);
nand U27368 (N_27368,N_26443,N_26332);
xnor U27369 (N_27369,N_26278,N_26295);
nor U27370 (N_27370,N_26830,N_26908);
and U27371 (N_27371,N_26311,N_26916);
and U27372 (N_27372,N_26620,N_26004);
and U27373 (N_27373,N_26808,N_26236);
and U27374 (N_27374,N_26157,N_26066);
and U27375 (N_27375,N_26859,N_26201);
nor U27376 (N_27376,N_26440,N_26257);
xor U27377 (N_27377,N_26002,N_26389);
nand U27378 (N_27378,N_26279,N_26683);
or U27379 (N_27379,N_26041,N_26480);
or U27380 (N_27380,N_26220,N_26194);
and U27381 (N_27381,N_26069,N_26096);
nor U27382 (N_27382,N_26107,N_26483);
nor U27383 (N_27383,N_26289,N_26724);
xnor U27384 (N_27384,N_26287,N_26499);
nand U27385 (N_27385,N_26765,N_26325);
or U27386 (N_27386,N_26491,N_26195);
nor U27387 (N_27387,N_26691,N_26064);
xnor U27388 (N_27388,N_26283,N_26110);
and U27389 (N_27389,N_26199,N_26653);
or U27390 (N_27390,N_26960,N_26118);
nor U27391 (N_27391,N_26947,N_26688);
nand U27392 (N_27392,N_26395,N_26141);
nor U27393 (N_27393,N_26582,N_26769);
nor U27394 (N_27394,N_26322,N_26920);
and U27395 (N_27395,N_26982,N_26703);
xor U27396 (N_27396,N_26614,N_26660);
or U27397 (N_27397,N_26731,N_26764);
nor U27398 (N_27398,N_26175,N_26535);
nor U27399 (N_27399,N_26052,N_26407);
nor U27400 (N_27400,N_26140,N_26147);
xnor U27401 (N_27401,N_26525,N_26875);
and U27402 (N_27402,N_26823,N_26001);
nand U27403 (N_27403,N_26105,N_26876);
nand U27404 (N_27404,N_26596,N_26380);
nor U27405 (N_27405,N_26094,N_26956);
and U27406 (N_27406,N_26392,N_26692);
xnor U27407 (N_27407,N_26255,N_26410);
and U27408 (N_27408,N_26022,N_26836);
and U27409 (N_27409,N_26426,N_26937);
xnor U27410 (N_27410,N_26231,N_26530);
and U27411 (N_27411,N_26136,N_26218);
xnor U27412 (N_27412,N_26029,N_26318);
and U27413 (N_27413,N_26149,N_26550);
nand U27414 (N_27414,N_26268,N_26135);
xnor U27415 (N_27415,N_26242,N_26630);
or U27416 (N_27416,N_26214,N_26551);
or U27417 (N_27417,N_26130,N_26003);
nor U27418 (N_27418,N_26985,N_26428);
nor U27419 (N_27419,N_26571,N_26772);
nand U27420 (N_27420,N_26156,N_26270);
nor U27421 (N_27421,N_26888,N_26513);
or U27422 (N_27422,N_26204,N_26291);
or U27423 (N_27423,N_26396,N_26377);
or U27424 (N_27424,N_26564,N_26877);
nand U27425 (N_27425,N_26929,N_26306);
nand U27426 (N_27426,N_26106,N_26812);
and U27427 (N_27427,N_26923,N_26659);
and U27428 (N_27428,N_26992,N_26502);
nand U27429 (N_27429,N_26216,N_26515);
or U27430 (N_27430,N_26341,N_26563);
nor U27431 (N_27431,N_26767,N_26856);
or U27432 (N_27432,N_26059,N_26021);
or U27433 (N_27433,N_26320,N_26560);
nand U27434 (N_27434,N_26286,N_26607);
and U27435 (N_27435,N_26458,N_26030);
or U27436 (N_27436,N_26928,N_26971);
and U27437 (N_27437,N_26625,N_26723);
nand U27438 (N_27438,N_26312,N_26925);
and U27439 (N_27439,N_26419,N_26835);
nor U27440 (N_27440,N_26670,N_26713);
xnor U27441 (N_27441,N_26695,N_26534);
nor U27442 (N_27442,N_26470,N_26129);
and U27443 (N_27443,N_26385,N_26091);
or U27444 (N_27444,N_26308,N_26433);
and U27445 (N_27445,N_26672,N_26809);
or U27446 (N_27446,N_26826,N_26811);
nand U27447 (N_27447,N_26781,N_26952);
nor U27448 (N_27448,N_26101,N_26471);
or U27449 (N_27449,N_26506,N_26434);
or U27450 (N_27450,N_26379,N_26342);
nor U27451 (N_27451,N_26803,N_26661);
nand U27452 (N_27452,N_26350,N_26746);
nor U27453 (N_27453,N_26599,N_26355);
or U27454 (N_27454,N_26963,N_26290);
and U27455 (N_27455,N_26817,N_26375);
and U27456 (N_27456,N_26093,N_26538);
nand U27457 (N_27457,N_26541,N_26358);
or U27458 (N_27458,N_26915,N_26045);
or U27459 (N_27459,N_26274,N_26365);
nand U27460 (N_27460,N_26911,N_26592);
and U27461 (N_27461,N_26164,N_26360);
nor U27462 (N_27462,N_26461,N_26173);
and U27463 (N_27463,N_26729,N_26485);
or U27464 (N_27464,N_26527,N_26034);
nor U27465 (N_27465,N_26489,N_26818);
nor U27466 (N_27466,N_26324,N_26111);
or U27467 (N_27467,N_26100,N_26223);
and U27468 (N_27468,N_26636,N_26083);
and U27469 (N_27469,N_26849,N_26898);
xnor U27470 (N_27470,N_26144,N_26806);
or U27471 (N_27471,N_26831,N_26842);
and U27472 (N_27472,N_26967,N_26119);
nand U27473 (N_27473,N_26523,N_26122);
xor U27474 (N_27474,N_26609,N_26595);
or U27475 (N_27475,N_26381,N_26374);
or U27476 (N_27476,N_26834,N_26143);
xnor U27477 (N_27477,N_26189,N_26329);
and U27478 (N_27478,N_26151,N_26663);
or U27479 (N_27479,N_26457,N_26813);
and U27480 (N_27480,N_26235,N_26516);
nor U27481 (N_27481,N_26427,N_26339);
or U27482 (N_27482,N_26627,N_26487);
nand U27483 (N_27483,N_26349,N_26962);
nor U27484 (N_27484,N_26761,N_26038);
and U27485 (N_27485,N_26225,N_26221);
nor U27486 (N_27486,N_26701,N_26624);
nor U27487 (N_27487,N_26838,N_26602);
or U27488 (N_27488,N_26671,N_26351);
nand U27489 (N_27489,N_26240,N_26356);
nand U27490 (N_27490,N_26601,N_26334);
or U27491 (N_27491,N_26721,N_26117);
or U27492 (N_27492,N_26791,N_26409);
or U27493 (N_27493,N_26023,N_26926);
nand U27494 (N_27494,N_26972,N_26644);
nor U27495 (N_27495,N_26648,N_26182);
nand U27496 (N_27496,N_26710,N_26098);
nor U27497 (N_27497,N_26133,N_26248);
nand U27498 (N_27498,N_26976,N_26191);
or U27499 (N_27499,N_26553,N_26313);
xnor U27500 (N_27500,N_26981,N_26023);
or U27501 (N_27501,N_26377,N_26806);
and U27502 (N_27502,N_26886,N_26155);
xor U27503 (N_27503,N_26797,N_26331);
nor U27504 (N_27504,N_26152,N_26867);
nor U27505 (N_27505,N_26268,N_26225);
or U27506 (N_27506,N_26129,N_26500);
nor U27507 (N_27507,N_26391,N_26537);
or U27508 (N_27508,N_26425,N_26424);
or U27509 (N_27509,N_26670,N_26494);
xor U27510 (N_27510,N_26791,N_26929);
or U27511 (N_27511,N_26606,N_26150);
xnor U27512 (N_27512,N_26540,N_26575);
nand U27513 (N_27513,N_26267,N_26727);
or U27514 (N_27514,N_26322,N_26340);
or U27515 (N_27515,N_26537,N_26373);
or U27516 (N_27516,N_26415,N_26565);
xnor U27517 (N_27517,N_26614,N_26460);
xor U27518 (N_27518,N_26331,N_26760);
nor U27519 (N_27519,N_26344,N_26683);
or U27520 (N_27520,N_26804,N_26793);
xnor U27521 (N_27521,N_26484,N_26435);
xnor U27522 (N_27522,N_26421,N_26714);
nor U27523 (N_27523,N_26521,N_26931);
xor U27524 (N_27524,N_26589,N_26466);
xor U27525 (N_27525,N_26414,N_26573);
and U27526 (N_27526,N_26127,N_26447);
and U27527 (N_27527,N_26115,N_26011);
nand U27528 (N_27528,N_26113,N_26283);
xor U27529 (N_27529,N_26413,N_26710);
xor U27530 (N_27530,N_26841,N_26594);
or U27531 (N_27531,N_26985,N_26120);
nand U27532 (N_27532,N_26007,N_26876);
or U27533 (N_27533,N_26823,N_26836);
xnor U27534 (N_27534,N_26471,N_26527);
xnor U27535 (N_27535,N_26704,N_26632);
nor U27536 (N_27536,N_26007,N_26505);
xnor U27537 (N_27537,N_26183,N_26069);
and U27538 (N_27538,N_26661,N_26668);
nand U27539 (N_27539,N_26608,N_26189);
nand U27540 (N_27540,N_26033,N_26862);
nand U27541 (N_27541,N_26599,N_26863);
nor U27542 (N_27542,N_26118,N_26852);
xnor U27543 (N_27543,N_26898,N_26872);
and U27544 (N_27544,N_26785,N_26511);
and U27545 (N_27545,N_26927,N_26928);
xnor U27546 (N_27546,N_26853,N_26659);
nor U27547 (N_27547,N_26601,N_26234);
xor U27548 (N_27548,N_26373,N_26016);
nand U27549 (N_27549,N_26334,N_26248);
and U27550 (N_27550,N_26370,N_26886);
nand U27551 (N_27551,N_26713,N_26292);
and U27552 (N_27552,N_26392,N_26584);
nand U27553 (N_27553,N_26618,N_26679);
or U27554 (N_27554,N_26979,N_26093);
xor U27555 (N_27555,N_26398,N_26457);
nand U27556 (N_27556,N_26431,N_26803);
nor U27557 (N_27557,N_26780,N_26386);
nand U27558 (N_27558,N_26364,N_26265);
nand U27559 (N_27559,N_26361,N_26188);
and U27560 (N_27560,N_26083,N_26456);
or U27561 (N_27561,N_26568,N_26408);
or U27562 (N_27562,N_26473,N_26766);
xnor U27563 (N_27563,N_26237,N_26980);
or U27564 (N_27564,N_26754,N_26832);
xor U27565 (N_27565,N_26442,N_26784);
or U27566 (N_27566,N_26088,N_26623);
nand U27567 (N_27567,N_26992,N_26076);
xor U27568 (N_27568,N_26474,N_26292);
or U27569 (N_27569,N_26396,N_26027);
or U27570 (N_27570,N_26427,N_26522);
nand U27571 (N_27571,N_26436,N_26791);
xor U27572 (N_27572,N_26120,N_26158);
nor U27573 (N_27573,N_26296,N_26270);
xor U27574 (N_27574,N_26769,N_26408);
nand U27575 (N_27575,N_26183,N_26902);
nor U27576 (N_27576,N_26783,N_26766);
xor U27577 (N_27577,N_26881,N_26926);
nor U27578 (N_27578,N_26404,N_26843);
or U27579 (N_27579,N_26769,N_26513);
nand U27580 (N_27580,N_26658,N_26188);
nor U27581 (N_27581,N_26445,N_26777);
xor U27582 (N_27582,N_26862,N_26073);
and U27583 (N_27583,N_26340,N_26975);
nor U27584 (N_27584,N_26418,N_26307);
nor U27585 (N_27585,N_26452,N_26580);
xnor U27586 (N_27586,N_26129,N_26987);
nor U27587 (N_27587,N_26018,N_26487);
nand U27588 (N_27588,N_26151,N_26560);
or U27589 (N_27589,N_26497,N_26654);
and U27590 (N_27590,N_26102,N_26877);
nor U27591 (N_27591,N_26385,N_26715);
or U27592 (N_27592,N_26976,N_26564);
nor U27593 (N_27593,N_26401,N_26784);
nand U27594 (N_27594,N_26668,N_26959);
and U27595 (N_27595,N_26451,N_26055);
or U27596 (N_27596,N_26575,N_26512);
nand U27597 (N_27597,N_26009,N_26567);
nor U27598 (N_27598,N_26808,N_26426);
nand U27599 (N_27599,N_26402,N_26406);
or U27600 (N_27600,N_26409,N_26728);
nand U27601 (N_27601,N_26169,N_26708);
or U27602 (N_27602,N_26968,N_26845);
or U27603 (N_27603,N_26439,N_26747);
and U27604 (N_27604,N_26852,N_26609);
nand U27605 (N_27605,N_26682,N_26600);
or U27606 (N_27606,N_26326,N_26377);
xnor U27607 (N_27607,N_26486,N_26112);
or U27608 (N_27608,N_26459,N_26502);
nor U27609 (N_27609,N_26282,N_26114);
xor U27610 (N_27610,N_26408,N_26158);
or U27611 (N_27611,N_26843,N_26957);
nor U27612 (N_27612,N_26229,N_26087);
and U27613 (N_27613,N_26550,N_26499);
xnor U27614 (N_27614,N_26538,N_26704);
or U27615 (N_27615,N_26258,N_26035);
nand U27616 (N_27616,N_26133,N_26180);
nor U27617 (N_27617,N_26839,N_26166);
xor U27618 (N_27618,N_26222,N_26810);
nor U27619 (N_27619,N_26315,N_26318);
and U27620 (N_27620,N_26768,N_26118);
and U27621 (N_27621,N_26895,N_26818);
nand U27622 (N_27622,N_26744,N_26616);
and U27623 (N_27623,N_26357,N_26911);
xor U27624 (N_27624,N_26837,N_26365);
nand U27625 (N_27625,N_26151,N_26626);
and U27626 (N_27626,N_26483,N_26521);
nor U27627 (N_27627,N_26029,N_26131);
and U27628 (N_27628,N_26705,N_26194);
and U27629 (N_27629,N_26465,N_26808);
or U27630 (N_27630,N_26511,N_26627);
and U27631 (N_27631,N_26844,N_26425);
or U27632 (N_27632,N_26261,N_26861);
xnor U27633 (N_27633,N_26542,N_26232);
or U27634 (N_27634,N_26178,N_26899);
or U27635 (N_27635,N_26033,N_26442);
nand U27636 (N_27636,N_26783,N_26145);
or U27637 (N_27637,N_26611,N_26265);
xor U27638 (N_27638,N_26140,N_26602);
nor U27639 (N_27639,N_26045,N_26934);
or U27640 (N_27640,N_26425,N_26744);
and U27641 (N_27641,N_26489,N_26377);
and U27642 (N_27642,N_26530,N_26062);
nor U27643 (N_27643,N_26034,N_26952);
xor U27644 (N_27644,N_26516,N_26815);
nand U27645 (N_27645,N_26065,N_26961);
nand U27646 (N_27646,N_26972,N_26178);
nand U27647 (N_27647,N_26534,N_26602);
xnor U27648 (N_27648,N_26627,N_26795);
and U27649 (N_27649,N_26057,N_26535);
xor U27650 (N_27650,N_26117,N_26870);
or U27651 (N_27651,N_26838,N_26715);
xor U27652 (N_27652,N_26660,N_26265);
or U27653 (N_27653,N_26608,N_26179);
nand U27654 (N_27654,N_26288,N_26984);
or U27655 (N_27655,N_26957,N_26332);
or U27656 (N_27656,N_26439,N_26052);
or U27657 (N_27657,N_26849,N_26834);
and U27658 (N_27658,N_26481,N_26245);
and U27659 (N_27659,N_26661,N_26722);
nor U27660 (N_27660,N_26878,N_26950);
or U27661 (N_27661,N_26553,N_26050);
xnor U27662 (N_27662,N_26443,N_26000);
nand U27663 (N_27663,N_26342,N_26001);
or U27664 (N_27664,N_26353,N_26061);
or U27665 (N_27665,N_26793,N_26225);
and U27666 (N_27666,N_26314,N_26539);
nor U27667 (N_27667,N_26306,N_26432);
or U27668 (N_27668,N_26267,N_26573);
xor U27669 (N_27669,N_26092,N_26520);
nor U27670 (N_27670,N_26575,N_26263);
nand U27671 (N_27671,N_26764,N_26100);
nor U27672 (N_27672,N_26830,N_26851);
nor U27673 (N_27673,N_26880,N_26169);
xnor U27674 (N_27674,N_26715,N_26724);
and U27675 (N_27675,N_26305,N_26857);
nand U27676 (N_27676,N_26863,N_26372);
nand U27677 (N_27677,N_26460,N_26610);
or U27678 (N_27678,N_26725,N_26702);
and U27679 (N_27679,N_26317,N_26128);
or U27680 (N_27680,N_26303,N_26291);
xnor U27681 (N_27681,N_26970,N_26547);
nor U27682 (N_27682,N_26903,N_26290);
nand U27683 (N_27683,N_26211,N_26782);
nand U27684 (N_27684,N_26311,N_26076);
nand U27685 (N_27685,N_26852,N_26821);
or U27686 (N_27686,N_26206,N_26021);
nand U27687 (N_27687,N_26485,N_26131);
and U27688 (N_27688,N_26100,N_26003);
xor U27689 (N_27689,N_26486,N_26956);
or U27690 (N_27690,N_26011,N_26064);
or U27691 (N_27691,N_26056,N_26969);
and U27692 (N_27692,N_26967,N_26277);
nand U27693 (N_27693,N_26193,N_26231);
nor U27694 (N_27694,N_26189,N_26050);
and U27695 (N_27695,N_26265,N_26391);
xor U27696 (N_27696,N_26480,N_26336);
nand U27697 (N_27697,N_26867,N_26813);
xnor U27698 (N_27698,N_26471,N_26463);
xor U27699 (N_27699,N_26002,N_26667);
nor U27700 (N_27700,N_26823,N_26942);
or U27701 (N_27701,N_26028,N_26168);
nor U27702 (N_27702,N_26805,N_26340);
nand U27703 (N_27703,N_26211,N_26668);
and U27704 (N_27704,N_26669,N_26384);
nor U27705 (N_27705,N_26521,N_26601);
and U27706 (N_27706,N_26731,N_26080);
nand U27707 (N_27707,N_26381,N_26176);
and U27708 (N_27708,N_26993,N_26037);
and U27709 (N_27709,N_26989,N_26170);
nand U27710 (N_27710,N_26519,N_26103);
nor U27711 (N_27711,N_26355,N_26284);
nor U27712 (N_27712,N_26571,N_26813);
nor U27713 (N_27713,N_26448,N_26542);
and U27714 (N_27714,N_26486,N_26797);
and U27715 (N_27715,N_26766,N_26886);
xor U27716 (N_27716,N_26664,N_26474);
or U27717 (N_27717,N_26900,N_26511);
or U27718 (N_27718,N_26629,N_26250);
and U27719 (N_27719,N_26522,N_26004);
or U27720 (N_27720,N_26650,N_26554);
xnor U27721 (N_27721,N_26503,N_26967);
or U27722 (N_27722,N_26668,N_26612);
nand U27723 (N_27723,N_26089,N_26879);
and U27724 (N_27724,N_26073,N_26621);
and U27725 (N_27725,N_26476,N_26283);
and U27726 (N_27726,N_26269,N_26472);
xnor U27727 (N_27727,N_26387,N_26454);
and U27728 (N_27728,N_26741,N_26249);
or U27729 (N_27729,N_26937,N_26372);
and U27730 (N_27730,N_26223,N_26936);
xor U27731 (N_27731,N_26618,N_26588);
nor U27732 (N_27732,N_26319,N_26508);
nand U27733 (N_27733,N_26740,N_26975);
and U27734 (N_27734,N_26574,N_26573);
nor U27735 (N_27735,N_26451,N_26364);
nor U27736 (N_27736,N_26336,N_26510);
nor U27737 (N_27737,N_26310,N_26982);
and U27738 (N_27738,N_26124,N_26091);
nand U27739 (N_27739,N_26941,N_26998);
nand U27740 (N_27740,N_26451,N_26896);
nand U27741 (N_27741,N_26641,N_26553);
and U27742 (N_27742,N_26804,N_26178);
and U27743 (N_27743,N_26192,N_26766);
xor U27744 (N_27744,N_26169,N_26739);
nand U27745 (N_27745,N_26852,N_26225);
nor U27746 (N_27746,N_26714,N_26064);
nand U27747 (N_27747,N_26955,N_26930);
or U27748 (N_27748,N_26488,N_26360);
and U27749 (N_27749,N_26888,N_26107);
or U27750 (N_27750,N_26329,N_26193);
or U27751 (N_27751,N_26790,N_26990);
and U27752 (N_27752,N_26881,N_26087);
and U27753 (N_27753,N_26562,N_26888);
and U27754 (N_27754,N_26364,N_26170);
and U27755 (N_27755,N_26349,N_26720);
and U27756 (N_27756,N_26529,N_26894);
and U27757 (N_27757,N_26984,N_26465);
nor U27758 (N_27758,N_26206,N_26955);
or U27759 (N_27759,N_26438,N_26097);
nor U27760 (N_27760,N_26656,N_26568);
and U27761 (N_27761,N_26047,N_26135);
or U27762 (N_27762,N_26913,N_26801);
nand U27763 (N_27763,N_26124,N_26451);
or U27764 (N_27764,N_26889,N_26242);
xor U27765 (N_27765,N_26807,N_26039);
nor U27766 (N_27766,N_26462,N_26539);
and U27767 (N_27767,N_26725,N_26817);
nor U27768 (N_27768,N_26056,N_26414);
or U27769 (N_27769,N_26169,N_26583);
nand U27770 (N_27770,N_26254,N_26314);
nor U27771 (N_27771,N_26225,N_26846);
nand U27772 (N_27772,N_26075,N_26386);
nor U27773 (N_27773,N_26689,N_26572);
or U27774 (N_27774,N_26072,N_26117);
or U27775 (N_27775,N_26535,N_26626);
or U27776 (N_27776,N_26263,N_26185);
xnor U27777 (N_27777,N_26230,N_26683);
nor U27778 (N_27778,N_26033,N_26649);
or U27779 (N_27779,N_26727,N_26047);
and U27780 (N_27780,N_26336,N_26235);
xnor U27781 (N_27781,N_26834,N_26280);
and U27782 (N_27782,N_26253,N_26266);
nor U27783 (N_27783,N_26700,N_26117);
nor U27784 (N_27784,N_26028,N_26318);
xnor U27785 (N_27785,N_26967,N_26835);
and U27786 (N_27786,N_26398,N_26112);
xor U27787 (N_27787,N_26408,N_26588);
or U27788 (N_27788,N_26065,N_26834);
and U27789 (N_27789,N_26410,N_26160);
and U27790 (N_27790,N_26039,N_26561);
and U27791 (N_27791,N_26761,N_26516);
and U27792 (N_27792,N_26796,N_26743);
and U27793 (N_27793,N_26805,N_26758);
and U27794 (N_27794,N_26638,N_26862);
nand U27795 (N_27795,N_26133,N_26760);
xor U27796 (N_27796,N_26633,N_26683);
and U27797 (N_27797,N_26121,N_26582);
or U27798 (N_27798,N_26217,N_26630);
nand U27799 (N_27799,N_26778,N_26013);
or U27800 (N_27800,N_26131,N_26774);
nand U27801 (N_27801,N_26332,N_26579);
nor U27802 (N_27802,N_26853,N_26081);
or U27803 (N_27803,N_26928,N_26655);
nor U27804 (N_27804,N_26181,N_26163);
and U27805 (N_27805,N_26527,N_26055);
xor U27806 (N_27806,N_26273,N_26946);
and U27807 (N_27807,N_26798,N_26846);
xnor U27808 (N_27808,N_26591,N_26864);
nor U27809 (N_27809,N_26901,N_26385);
nor U27810 (N_27810,N_26670,N_26525);
nand U27811 (N_27811,N_26877,N_26769);
xnor U27812 (N_27812,N_26225,N_26881);
or U27813 (N_27813,N_26619,N_26373);
xor U27814 (N_27814,N_26130,N_26307);
xnor U27815 (N_27815,N_26835,N_26762);
and U27816 (N_27816,N_26950,N_26306);
nand U27817 (N_27817,N_26553,N_26255);
nor U27818 (N_27818,N_26531,N_26487);
xnor U27819 (N_27819,N_26486,N_26714);
and U27820 (N_27820,N_26718,N_26755);
xnor U27821 (N_27821,N_26914,N_26096);
or U27822 (N_27822,N_26311,N_26548);
nand U27823 (N_27823,N_26035,N_26802);
xor U27824 (N_27824,N_26675,N_26211);
and U27825 (N_27825,N_26566,N_26028);
and U27826 (N_27826,N_26675,N_26881);
or U27827 (N_27827,N_26442,N_26990);
nand U27828 (N_27828,N_26851,N_26659);
and U27829 (N_27829,N_26892,N_26474);
xor U27830 (N_27830,N_26522,N_26634);
xnor U27831 (N_27831,N_26224,N_26779);
xnor U27832 (N_27832,N_26563,N_26716);
xnor U27833 (N_27833,N_26682,N_26618);
and U27834 (N_27834,N_26514,N_26869);
xnor U27835 (N_27835,N_26316,N_26653);
nor U27836 (N_27836,N_26498,N_26958);
and U27837 (N_27837,N_26700,N_26079);
xnor U27838 (N_27838,N_26064,N_26670);
and U27839 (N_27839,N_26270,N_26931);
xnor U27840 (N_27840,N_26861,N_26544);
or U27841 (N_27841,N_26525,N_26667);
nand U27842 (N_27842,N_26347,N_26726);
xor U27843 (N_27843,N_26808,N_26314);
nor U27844 (N_27844,N_26396,N_26439);
nand U27845 (N_27845,N_26086,N_26983);
or U27846 (N_27846,N_26303,N_26209);
xnor U27847 (N_27847,N_26536,N_26810);
xnor U27848 (N_27848,N_26661,N_26252);
nor U27849 (N_27849,N_26961,N_26287);
and U27850 (N_27850,N_26827,N_26478);
and U27851 (N_27851,N_26929,N_26512);
xnor U27852 (N_27852,N_26105,N_26305);
nor U27853 (N_27853,N_26495,N_26363);
xnor U27854 (N_27854,N_26454,N_26288);
nor U27855 (N_27855,N_26769,N_26476);
xor U27856 (N_27856,N_26954,N_26389);
nor U27857 (N_27857,N_26379,N_26437);
nor U27858 (N_27858,N_26891,N_26618);
xor U27859 (N_27859,N_26894,N_26521);
nor U27860 (N_27860,N_26034,N_26241);
or U27861 (N_27861,N_26275,N_26766);
or U27862 (N_27862,N_26705,N_26385);
nand U27863 (N_27863,N_26942,N_26102);
or U27864 (N_27864,N_26951,N_26282);
or U27865 (N_27865,N_26755,N_26694);
nand U27866 (N_27866,N_26722,N_26674);
or U27867 (N_27867,N_26346,N_26788);
or U27868 (N_27868,N_26015,N_26685);
nor U27869 (N_27869,N_26647,N_26430);
xor U27870 (N_27870,N_26845,N_26596);
or U27871 (N_27871,N_26392,N_26438);
xnor U27872 (N_27872,N_26596,N_26546);
nand U27873 (N_27873,N_26636,N_26355);
xor U27874 (N_27874,N_26637,N_26147);
or U27875 (N_27875,N_26821,N_26159);
and U27876 (N_27876,N_26746,N_26770);
or U27877 (N_27877,N_26757,N_26831);
nand U27878 (N_27878,N_26302,N_26030);
or U27879 (N_27879,N_26981,N_26877);
nand U27880 (N_27880,N_26446,N_26119);
xor U27881 (N_27881,N_26115,N_26701);
xnor U27882 (N_27882,N_26250,N_26709);
or U27883 (N_27883,N_26700,N_26691);
or U27884 (N_27884,N_26169,N_26258);
and U27885 (N_27885,N_26695,N_26543);
xor U27886 (N_27886,N_26926,N_26816);
nor U27887 (N_27887,N_26406,N_26505);
and U27888 (N_27888,N_26067,N_26639);
or U27889 (N_27889,N_26277,N_26832);
nand U27890 (N_27890,N_26815,N_26334);
nand U27891 (N_27891,N_26128,N_26471);
nor U27892 (N_27892,N_26280,N_26099);
nand U27893 (N_27893,N_26998,N_26283);
nor U27894 (N_27894,N_26522,N_26069);
and U27895 (N_27895,N_26890,N_26099);
nand U27896 (N_27896,N_26973,N_26919);
and U27897 (N_27897,N_26412,N_26858);
and U27898 (N_27898,N_26389,N_26929);
nand U27899 (N_27899,N_26839,N_26017);
and U27900 (N_27900,N_26913,N_26455);
and U27901 (N_27901,N_26823,N_26272);
or U27902 (N_27902,N_26346,N_26644);
nand U27903 (N_27903,N_26373,N_26659);
xnor U27904 (N_27904,N_26296,N_26835);
nor U27905 (N_27905,N_26783,N_26595);
nor U27906 (N_27906,N_26202,N_26867);
xnor U27907 (N_27907,N_26380,N_26460);
xnor U27908 (N_27908,N_26494,N_26434);
xor U27909 (N_27909,N_26368,N_26297);
and U27910 (N_27910,N_26513,N_26872);
nor U27911 (N_27911,N_26448,N_26990);
nand U27912 (N_27912,N_26394,N_26744);
and U27913 (N_27913,N_26853,N_26788);
and U27914 (N_27914,N_26042,N_26073);
xnor U27915 (N_27915,N_26059,N_26809);
nand U27916 (N_27916,N_26252,N_26453);
nor U27917 (N_27917,N_26963,N_26505);
and U27918 (N_27918,N_26015,N_26090);
or U27919 (N_27919,N_26642,N_26707);
nor U27920 (N_27920,N_26344,N_26877);
xnor U27921 (N_27921,N_26749,N_26907);
nor U27922 (N_27922,N_26122,N_26342);
and U27923 (N_27923,N_26004,N_26271);
or U27924 (N_27924,N_26291,N_26219);
xor U27925 (N_27925,N_26839,N_26822);
nand U27926 (N_27926,N_26814,N_26411);
nand U27927 (N_27927,N_26380,N_26398);
and U27928 (N_27928,N_26716,N_26658);
nand U27929 (N_27929,N_26127,N_26481);
and U27930 (N_27930,N_26804,N_26107);
xor U27931 (N_27931,N_26963,N_26897);
nand U27932 (N_27932,N_26370,N_26645);
or U27933 (N_27933,N_26919,N_26171);
nor U27934 (N_27934,N_26597,N_26205);
nand U27935 (N_27935,N_26078,N_26255);
or U27936 (N_27936,N_26359,N_26318);
nand U27937 (N_27937,N_26864,N_26096);
and U27938 (N_27938,N_26143,N_26890);
and U27939 (N_27939,N_26991,N_26855);
nand U27940 (N_27940,N_26357,N_26371);
and U27941 (N_27941,N_26595,N_26152);
nand U27942 (N_27942,N_26479,N_26810);
or U27943 (N_27943,N_26272,N_26363);
and U27944 (N_27944,N_26944,N_26199);
nor U27945 (N_27945,N_26282,N_26906);
nor U27946 (N_27946,N_26042,N_26121);
nor U27947 (N_27947,N_26646,N_26573);
nor U27948 (N_27948,N_26337,N_26635);
and U27949 (N_27949,N_26384,N_26320);
xnor U27950 (N_27950,N_26002,N_26243);
xor U27951 (N_27951,N_26603,N_26088);
xnor U27952 (N_27952,N_26584,N_26900);
and U27953 (N_27953,N_26245,N_26990);
and U27954 (N_27954,N_26036,N_26357);
or U27955 (N_27955,N_26754,N_26377);
and U27956 (N_27956,N_26796,N_26783);
nor U27957 (N_27957,N_26434,N_26919);
nand U27958 (N_27958,N_26450,N_26887);
nor U27959 (N_27959,N_26850,N_26538);
and U27960 (N_27960,N_26729,N_26065);
nand U27961 (N_27961,N_26586,N_26353);
nand U27962 (N_27962,N_26318,N_26925);
and U27963 (N_27963,N_26987,N_26045);
xnor U27964 (N_27964,N_26529,N_26518);
xor U27965 (N_27965,N_26901,N_26601);
xnor U27966 (N_27966,N_26192,N_26234);
xor U27967 (N_27967,N_26170,N_26482);
and U27968 (N_27968,N_26060,N_26100);
xor U27969 (N_27969,N_26306,N_26653);
nand U27970 (N_27970,N_26970,N_26549);
nor U27971 (N_27971,N_26671,N_26449);
nor U27972 (N_27972,N_26370,N_26817);
xnor U27973 (N_27973,N_26370,N_26567);
xnor U27974 (N_27974,N_26510,N_26583);
xor U27975 (N_27975,N_26210,N_26316);
or U27976 (N_27976,N_26238,N_26935);
nor U27977 (N_27977,N_26134,N_26301);
nor U27978 (N_27978,N_26931,N_26342);
and U27979 (N_27979,N_26893,N_26902);
and U27980 (N_27980,N_26776,N_26503);
or U27981 (N_27981,N_26856,N_26526);
nand U27982 (N_27982,N_26553,N_26134);
or U27983 (N_27983,N_26150,N_26555);
and U27984 (N_27984,N_26918,N_26638);
or U27985 (N_27985,N_26709,N_26898);
nand U27986 (N_27986,N_26966,N_26696);
or U27987 (N_27987,N_26134,N_26265);
nor U27988 (N_27988,N_26099,N_26835);
nand U27989 (N_27989,N_26455,N_26151);
nor U27990 (N_27990,N_26519,N_26575);
xor U27991 (N_27991,N_26031,N_26602);
or U27992 (N_27992,N_26551,N_26035);
and U27993 (N_27993,N_26499,N_26372);
xor U27994 (N_27994,N_26352,N_26598);
xor U27995 (N_27995,N_26467,N_26775);
and U27996 (N_27996,N_26849,N_26371);
xor U27997 (N_27997,N_26165,N_26639);
and U27998 (N_27998,N_26214,N_26215);
and U27999 (N_27999,N_26362,N_26328);
or U28000 (N_28000,N_27672,N_27514);
or U28001 (N_28001,N_27253,N_27243);
and U28002 (N_28002,N_27978,N_27247);
nand U28003 (N_28003,N_27115,N_27378);
and U28004 (N_28004,N_27915,N_27536);
nor U28005 (N_28005,N_27974,N_27999);
and U28006 (N_28006,N_27187,N_27393);
nand U28007 (N_28007,N_27129,N_27729);
or U28008 (N_28008,N_27359,N_27568);
nand U28009 (N_28009,N_27364,N_27071);
xor U28010 (N_28010,N_27964,N_27108);
nand U28011 (N_28011,N_27264,N_27728);
nand U28012 (N_28012,N_27913,N_27366);
xor U28013 (N_28013,N_27020,N_27120);
nand U28014 (N_28014,N_27440,N_27846);
nor U28015 (N_28015,N_27311,N_27621);
nand U28016 (N_28016,N_27177,N_27347);
nand U28017 (N_28017,N_27124,N_27906);
and U28018 (N_28018,N_27350,N_27426);
and U28019 (N_28019,N_27060,N_27268);
nor U28020 (N_28020,N_27746,N_27315);
or U28021 (N_28021,N_27967,N_27692);
and U28022 (N_28022,N_27618,N_27307);
nor U28023 (N_28023,N_27611,N_27442);
or U28024 (N_28024,N_27153,N_27374);
or U28025 (N_28025,N_27794,N_27168);
and U28026 (N_28026,N_27972,N_27832);
and U28027 (N_28027,N_27863,N_27866);
nand U28028 (N_28028,N_27021,N_27560);
nor U28029 (N_28029,N_27284,N_27154);
nand U28030 (N_28030,N_27919,N_27767);
and U28031 (N_28031,N_27626,N_27569);
xnor U28032 (N_28032,N_27041,N_27281);
and U28033 (N_28033,N_27218,N_27445);
xnor U28034 (N_28034,N_27305,N_27556);
nand U28035 (N_28035,N_27877,N_27959);
nand U28036 (N_28036,N_27766,N_27555);
xnor U28037 (N_28037,N_27046,N_27743);
nor U28038 (N_28038,N_27322,N_27839);
xor U28039 (N_28039,N_27603,N_27163);
or U28040 (N_28040,N_27969,N_27221);
and U28041 (N_28041,N_27271,N_27927);
or U28042 (N_28042,N_27971,N_27418);
or U28043 (N_28043,N_27771,N_27585);
and U28044 (N_28044,N_27539,N_27173);
and U28045 (N_28045,N_27326,N_27921);
xnor U28046 (N_28046,N_27903,N_27107);
or U28047 (N_28047,N_27130,N_27044);
nand U28048 (N_28048,N_27151,N_27096);
nand U28049 (N_28049,N_27605,N_27095);
nor U28050 (N_28050,N_27270,N_27048);
nand U28051 (N_28051,N_27865,N_27678);
and U28052 (N_28052,N_27697,N_27349);
nor U28053 (N_28053,N_27714,N_27637);
xor U28054 (N_28054,N_27127,N_27362);
xor U28055 (N_28055,N_27966,N_27586);
xnor U28056 (N_28056,N_27646,N_27227);
and U28057 (N_28057,N_27195,N_27700);
or U28058 (N_28058,N_27848,N_27008);
nand U28059 (N_28059,N_27564,N_27749);
nor U28060 (N_28060,N_27702,N_27273);
nor U28061 (N_28061,N_27795,N_27880);
nand U28062 (N_28062,N_27402,N_27878);
xnor U28063 (N_28063,N_27252,N_27417);
xnor U28064 (N_28064,N_27067,N_27689);
or U28065 (N_28065,N_27790,N_27787);
xnor U28066 (N_28066,N_27132,N_27354);
or U28067 (N_28067,N_27782,N_27197);
nor U28068 (N_28068,N_27982,N_27502);
and U28069 (N_28069,N_27612,N_27780);
xnor U28070 (N_28070,N_27504,N_27939);
nor U28071 (N_28071,N_27506,N_27294);
xnor U28072 (N_28072,N_27406,N_27431);
nand U28073 (N_28073,N_27109,N_27024);
or U28074 (N_28074,N_27070,N_27463);
or U28075 (N_28075,N_27570,N_27002);
and U28076 (N_28076,N_27357,N_27731);
nor U28077 (N_28077,N_27777,N_27471);
xnor U28078 (N_28078,N_27818,N_27340);
nand U28079 (N_28079,N_27031,N_27664);
nor U28080 (N_28080,N_27812,N_27114);
and U28081 (N_28081,N_27503,N_27673);
and U28082 (N_28082,N_27118,N_27543);
and U28083 (N_28083,N_27867,N_27607);
nor U28084 (N_28084,N_27005,N_27996);
nor U28085 (N_28085,N_27352,N_27019);
and U28086 (N_28086,N_27758,N_27303);
and U28087 (N_28087,N_27926,N_27206);
and U28088 (N_28088,N_27995,N_27458);
and U28089 (N_28089,N_27285,N_27488);
nand U28090 (N_28090,N_27047,N_27407);
or U28091 (N_28091,N_27188,N_27744);
or U28092 (N_28092,N_27475,N_27219);
and U28093 (N_28093,N_27824,N_27935);
xnor U28094 (N_28094,N_27876,N_27547);
nand U28095 (N_28095,N_27314,N_27075);
nand U28096 (N_28096,N_27499,N_27479);
xor U28097 (N_28097,N_27051,N_27335);
nor U28098 (N_28098,N_27566,N_27437);
or U28099 (N_28099,N_27583,N_27461);
xnor U28100 (N_28100,N_27466,N_27822);
xor U28101 (N_28101,N_27868,N_27477);
xor U28102 (N_28102,N_27806,N_27596);
nand U28103 (N_28103,N_27616,N_27713);
nor U28104 (N_28104,N_27233,N_27639);
xnor U28105 (N_28105,N_27941,N_27738);
nand U28106 (N_28106,N_27811,N_27396);
nor U28107 (N_28107,N_27676,N_27801);
nor U28108 (N_28108,N_27199,N_27057);
xnor U28109 (N_28109,N_27111,N_27981);
nor U28110 (N_28110,N_27094,N_27994);
and U28111 (N_28111,N_27361,N_27537);
xor U28112 (N_28112,N_27797,N_27453);
nand U28113 (N_28113,N_27269,N_27381);
nand U28114 (N_28114,N_27950,N_27201);
and U28115 (N_28115,N_27662,N_27561);
nand U28116 (N_28116,N_27302,N_27126);
and U28117 (N_28117,N_27222,N_27148);
and U28118 (N_28118,N_27166,N_27186);
xnor U28119 (N_28119,N_27313,N_27419);
or U28120 (N_28120,N_27263,N_27558);
xor U28121 (N_28121,N_27617,N_27602);
nand U28122 (N_28122,N_27376,N_27256);
nor U28123 (N_28123,N_27844,N_27892);
nor U28124 (N_28124,N_27571,N_27367);
and U28125 (N_28125,N_27933,N_27891);
or U28126 (N_28126,N_27368,N_27146);
and U28127 (N_28127,N_27527,N_27589);
nor U28128 (N_28128,N_27432,N_27784);
nand U28129 (N_28129,N_27698,N_27338);
nor U28130 (N_28130,N_27141,N_27429);
or U28131 (N_28131,N_27510,N_27295);
or U28132 (N_28132,N_27992,N_27321);
nor U28133 (N_28133,N_27371,N_27103);
xnor U28134 (N_28134,N_27144,N_27392);
and U28135 (N_28135,N_27920,N_27924);
and U28136 (N_28136,N_27879,N_27807);
nand U28137 (N_28137,N_27137,N_27989);
and U28138 (N_28138,N_27379,N_27316);
xnor U28139 (N_28139,N_27369,N_27128);
nor U28140 (N_28140,N_27375,N_27291);
and U28141 (N_28141,N_27881,N_27834);
and U28142 (N_28142,N_27736,N_27957);
nand U28143 (N_28143,N_27632,N_27727);
xor U28144 (N_28144,N_27754,N_27423);
and U28145 (N_28145,N_27685,N_27870);
xor U28146 (N_28146,N_27803,N_27712);
nand U28147 (N_28147,N_27883,N_27521);
xor U28148 (N_28148,N_27980,N_27557);
and U28149 (N_28149,N_27175,N_27296);
nor U28150 (N_28150,N_27851,N_27424);
nor U28151 (N_28151,N_27360,N_27099);
or U28152 (N_28152,N_27204,N_27745);
nand U28153 (N_28153,N_27582,N_27280);
or U28154 (N_28154,N_27319,N_27748);
nand U28155 (N_28155,N_27753,N_27363);
xor U28156 (N_28156,N_27170,N_27182);
nand U28157 (N_28157,N_27793,N_27854);
nor U28158 (N_28158,N_27733,N_27654);
nand U28159 (N_28159,N_27925,N_27224);
xor U28160 (N_28160,N_27155,N_27191);
nor U28161 (N_28161,N_27715,N_27985);
and U28162 (N_28162,N_27434,N_27436);
nand U28163 (N_28163,N_27703,N_27087);
and U28164 (N_28164,N_27277,N_27472);
and U28165 (N_28165,N_27056,N_27819);
nor U28166 (N_28166,N_27604,N_27174);
xnor U28167 (N_28167,N_27549,N_27055);
xor U28168 (N_28168,N_27304,N_27559);
xnor U28169 (N_28169,N_27414,N_27827);
xor U28170 (N_28170,N_27526,N_27874);
nor U28171 (N_28171,N_27420,N_27653);
or U28172 (N_28172,N_27231,N_27165);
nand U28173 (N_28173,N_27501,N_27332);
or U28174 (N_28174,N_27635,N_27783);
xor U28175 (N_28175,N_27934,N_27306);
nor U28176 (N_28176,N_27600,N_27886);
and U28177 (N_28177,N_27449,N_27988);
xnor U28178 (N_28178,N_27760,N_27283);
xnor U28179 (N_28179,N_27389,N_27872);
nor U28180 (N_28180,N_27433,N_27553);
xnor U28181 (N_28181,N_27750,N_27532);
xnor U28182 (N_28182,N_27235,N_27644);
and U28183 (N_28183,N_27149,N_27772);
nor U28184 (N_28184,N_27741,N_27929);
or U28185 (N_28185,N_27648,N_27388);
or U28186 (N_28186,N_27318,N_27975);
xnor U28187 (N_28187,N_27911,N_27462);
nand U28188 (N_28188,N_27608,N_27976);
nor U28189 (N_28189,N_27542,N_27403);
nor U28190 (N_28190,N_27507,N_27497);
nand U28191 (N_28191,N_27010,N_27049);
and U28192 (N_28192,N_27932,N_27356);
xnor U28193 (N_28193,N_27524,N_27039);
and U28194 (N_28194,N_27486,N_27439);
xnor U28195 (N_28195,N_27266,N_27732);
xor U28196 (N_28196,N_27718,N_27251);
xor U28197 (N_28197,N_27342,N_27123);
and U28198 (N_28198,N_27970,N_27106);
xor U28199 (N_28199,N_27457,N_27694);
and U28200 (N_28200,N_27482,N_27198);
and U28201 (N_28201,N_27261,N_27387);
or U28202 (N_28202,N_27825,N_27073);
or U28203 (N_28203,N_27837,N_27757);
nor U28204 (N_28204,N_27216,N_27341);
nor U28205 (N_28205,N_27565,N_27343);
xor U28206 (N_28206,N_27829,N_27373);
or U28207 (N_28207,N_27917,N_27152);
xnor U28208 (N_28208,N_27724,N_27956);
nor U28209 (N_28209,N_27642,N_27677);
xnor U28210 (N_28210,N_27215,N_27668);
xnor U28211 (N_28211,N_27563,N_27905);
and U28212 (N_28212,N_27998,N_27276);
xor U28213 (N_28213,N_27993,N_27258);
nor U28214 (N_28214,N_27135,N_27140);
and U28215 (N_28215,N_27657,N_27562);
xnor U28216 (N_28216,N_27548,N_27297);
or U28217 (N_28217,N_27113,N_27147);
or U28218 (N_28218,N_27701,N_27820);
nand U28219 (N_28219,N_27828,N_27489);
xor U28220 (N_28220,N_27228,N_27534);
nor U28221 (N_28221,N_27282,N_27320);
and U28222 (N_28222,N_27640,N_27699);
nor U28223 (N_28223,N_27117,N_27210);
nand U28224 (N_28224,N_27172,N_27598);
xnor U28225 (N_28225,N_27018,N_27546);
and U28226 (N_28226,N_27068,N_27826);
and U28227 (N_28227,N_27591,N_27882);
and U28228 (N_28228,N_27412,N_27916);
xor U28229 (N_28229,N_27451,N_27441);
xnor U28230 (N_28230,N_27237,N_27962);
nand U28231 (N_28231,N_27674,N_27695);
and U28232 (N_28232,N_27945,N_27841);
nor U28233 (N_28233,N_27597,N_27914);
nand U28234 (N_28234,N_27336,N_27234);
xnor U28235 (N_28235,N_27930,N_27290);
nor U28236 (N_28236,N_27409,N_27456);
nand U28237 (N_28237,N_27923,N_27977);
or U28238 (N_28238,N_27652,N_27178);
nor U28239 (N_28239,N_27181,N_27908);
nor U28240 (N_28240,N_27082,N_27208);
or U28241 (N_28241,N_27333,N_27249);
and U28242 (N_28242,N_27791,N_27734);
xor U28243 (N_28243,N_27059,N_27323);
xor U28244 (N_28244,N_27833,N_27014);
xor U28245 (N_28245,N_27544,N_27943);
nor U28246 (N_28246,N_27669,N_27858);
nand U28247 (N_28247,N_27798,N_27465);
and U28248 (N_28248,N_27800,N_27383);
nor U28249 (N_28249,N_27480,N_27004);
and U28250 (N_28250,N_27751,N_27464);
xor U28251 (N_28251,N_27317,N_27370);
nor U28252 (N_28252,N_27158,N_27520);
nand U28253 (N_28253,N_27029,N_27896);
and U28254 (N_28254,N_27830,N_27551);
and U28255 (N_28255,N_27606,N_27267);
nand U28256 (N_28256,N_27609,N_27345);
or U28257 (N_28257,N_27042,N_27469);
xor U28258 (N_28258,N_27481,N_27080);
nor U28259 (N_28259,N_27889,N_27740);
xor U28260 (N_28260,N_27590,N_27428);
and U28261 (N_28261,N_27601,N_27159);
and U28262 (N_28262,N_27448,N_27491);
nand U28263 (N_28263,N_27952,N_27078);
nor U28264 (N_28264,N_27203,N_27622);
nand U28265 (N_28265,N_27006,N_27245);
nor U28266 (N_28266,N_27443,N_27190);
and U28267 (N_28267,N_27627,N_27131);
nor U28268 (N_28268,N_27398,N_27438);
nand U28269 (N_28269,N_27847,N_27660);
and U28270 (N_28270,N_27963,N_27898);
nand U28271 (N_28271,N_27003,N_27397);
nand U28272 (N_28272,N_27885,N_27211);
nand U28273 (N_28273,N_27965,N_27272);
xor U28274 (N_28274,N_27647,N_27064);
xnor U28275 (N_28275,N_27244,N_27902);
xor U28276 (N_28276,N_27893,N_27142);
nor U28277 (N_28277,N_27789,N_27408);
or U28278 (N_28278,N_27391,N_27192);
xor U28279 (N_28279,N_27721,N_27579);
nand U28280 (N_28280,N_27884,N_27139);
or U28281 (N_28281,N_27675,N_27085);
or U28282 (N_28282,N_27116,N_27101);
or U28283 (N_28283,N_27084,N_27027);
nor U28284 (N_28284,N_27455,N_27540);
xnor U28285 (N_28285,N_27167,N_27016);
nand U28286 (N_28286,N_27577,N_27250);
nand U28287 (N_28287,N_27949,N_27991);
nand U28288 (N_28288,N_27940,N_27688);
nand U28289 (N_28289,N_27217,N_27092);
or U28290 (N_28290,N_27979,N_27776);
xnor U28291 (N_28291,N_27200,N_27704);
nor U28292 (N_28292,N_27452,N_27805);
xnor U28293 (N_28293,N_27768,N_27459);
nor U28294 (N_28294,N_27658,N_27567);
or U28295 (N_28295,N_27292,N_27293);
and U28296 (N_28296,N_27063,N_27160);
or U28297 (N_28297,N_27013,N_27756);
nand U28298 (N_28298,N_27860,N_27337);
and U28299 (N_28299,N_27852,N_27009);
xnor U28300 (N_28300,N_27380,N_27512);
and U28301 (N_28301,N_27535,N_27220);
or U28302 (N_28302,N_27100,N_27960);
and U28303 (N_28303,N_27835,N_27705);
xor U28304 (N_28304,N_27817,N_27573);
nand U28305 (N_28305,N_27871,N_27638);
or U28306 (N_28306,N_27894,N_27679);
nand U28307 (N_28307,N_27665,N_27125);
nand U28308 (N_28308,N_27595,N_27083);
nor U28309 (N_28309,N_27522,N_27136);
nand U28310 (N_28310,N_27809,N_27015);
nand U28311 (N_28311,N_27184,N_27089);
nor U28312 (N_28312,N_27509,N_27786);
and U28313 (N_28313,N_27859,N_27873);
or U28314 (N_28314,N_27254,N_27575);
xor U28315 (N_28315,N_27299,N_27189);
and U28316 (N_28316,N_27017,N_27619);
xor U28317 (N_28317,N_27467,N_27840);
or U28318 (N_28318,N_27990,N_27102);
or U28319 (N_28319,N_27620,N_27659);
and U28320 (N_28320,N_27810,N_27265);
and U28321 (N_28321,N_27377,N_27650);
nor U28322 (N_28322,N_27492,N_27470);
nor U28323 (N_28323,N_27761,N_27328);
and U28324 (N_28324,N_27802,N_27987);
nor U28325 (N_28325,N_27788,N_27196);
or U28326 (N_28326,N_27580,N_27661);
xnor U28327 (N_28327,N_27836,N_27578);
nor U28328 (N_28328,N_27325,N_27358);
xnor U28329 (N_28329,N_27246,N_27496);
nor U28330 (N_28330,N_27112,N_27682);
nor U28331 (N_28331,N_27339,N_27156);
nand U28332 (N_28332,N_27110,N_27773);
or U28333 (N_28333,N_27843,N_27735);
xor U28334 (N_28334,N_27842,N_27717);
nor U28335 (N_28335,N_27645,N_27907);
and U28336 (N_28336,N_27900,N_27236);
nor U28337 (N_28337,N_27447,N_27001);
or U28338 (N_28338,N_27856,N_27747);
nand U28339 (N_28339,N_27726,N_27023);
xnor U28340 (N_28340,N_27242,N_27091);
or U28341 (N_28341,N_27026,N_27636);
or U28342 (N_28342,N_27515,N_27038);
nand U28343 (N_28343,N_27683,N_27594);
nand U28344 (N_28344,N_27212,N_27799);
xnor U28345 (N_28345,N_27072,N_27631);
xor U28346 (N_28346,N_27719,N_27725);
nand U28347 (N_28347,N_27054,N_27690);
xnor U28348 (N_28348,N_27308,N_27531);
and U28349 (N_28349,N_27416,N_27922);
or U28350 (N_28350,N_27400,N_27473);
or U28351 (N_28351,N_27936,N_27034);
nand U28352 (N_28352,N_27530,N_27385);
and U28353 (N_28353,N_27427,N_27176);
nand U28354 (N_28354,N_27098,N_27150);
or U28355 (N_28355,N_27498,N_27888);
nand U28356 (N_28356,N_27209,N_27331);
nand U28357 (N_28357,N_27225,N_27525);
nand U28358 (N_28358,N_27671,N_27779);
or U28359 (N_28359,N_27710,N_27194);
nor U28360 (N_28360,N_27122,N_27739);
nand U28361 (N_28361,N_27223,N_27000);
nand U28362 (N_28362,N_27804,N_27552);
nand U28363 (N_28363,N_27239,N_27649);
or U28364 (N_28364,N_27425,N_27062);
nand U28365 (N_28365,N_27484,N_27415);
or U28366 (N_28366,N_27850,N_27505);
or U28367 (N_28367,N_27327,N_27355);
xor U28368 (N_28368,N_27781,N_27937);
nand U28369 (N_28369,N_27968,N_27730);
nand U28370 (N_28370,N_27613,N_27887);
and U28371 (N_28371,N_27869,N_27610);
nor U28372 (N_28372,N_27651,N_27997);
and U28373 (N_28373,N_27032,N_27025);
and U28374 (N_28374,N_27759,N_27275);
nand U28375 (N_28375,N_27478,N_27955);
nand U28376 (N_28376,N_27289,N_27667);
and U28377 (N_28377,N_27814,N_27298);
xor U28378 (N_28378,N_27404,N_27944);
xnor U28379 (N_28379,N_27686,N_27614);
xnor U28380 (N_28380,N_27823,N_27588);
or U28381 (N_28381,N_27052,N_27214);
or U28382 (N_28382,N_27708,N_27769);
and U28383 (N_28383,N_27058,N_27716);
or U28384 (N_28384,N_27845,N_27774);
or U28385 (N_28385,N_27696,N_27951);
and U28386 (N_28386,N_27193,N_27468);
nor U28387 (N_28387,N_27770,N_27365);
nand U28388 (N_28388,N_27711,N_27986);
or U28389 (N_28389,N_27931,N_27630);
nand U28390 (N_28390,N_27641,N_27435);
xnor U28391 (N_28391,N_27813,N_27351);
nor U28392 (N_28392,N_27069,N_27121);
nand U28393 (N_28393,N_27500,N_27928);
or U28394 (N_28394,N_27904,N_27162);
or U28395 (N_28395,N_27909,N_27778);
nand U28396 (N_28396,N_27061,N_27035);
xor U28397 (N_28397,N_27628,N_27693);
nor U28398 (N_28398,N_27330,N_27161);
xnor U28399 (N_28399,N_27036,N_27495);
nor U28400 (N_28400,N_27324,N_27581);
or U28401 (N_28401,N_27076,N_27576);
nor U28402 (N_28402,N_27045,N_27384);
xor U28403 (N_28403,N_27528,N_27516);
xor U28404 (N_28404,N_27584,N_27623);
xor U28405 (N_28405,N_27763,N_27742);
xor U28406 (N_28406,N_27947,N_27229);
or U28407 (N_28407,N_27104,N_27572);
nand U28408 (N_28408,N_27494,N_27709);
nor U28409 (N_28409,N_27309,N_27513);
nand U28410 (N_28410,N_27259,N_27226);
nor U28411 (N_28411,N_27446,N_27086);
nor U28412 (N_28412,N_27954,N_27460);
or U28413 (N_28413,N_27853,N_27663);
or U28414 (N_28414,N_27961,N_27138);
and U28415 (N_28415,N_27279,N_27401);
and U28416 (N_28416,N_27353,N_27119);
or U28417 (N_28417,N_27529,N_27179);
nor U28418 (N_28418,N_27205,N_27762);
nor U28419 (N_28419,N_27680,N_27946);
and U28420 (N_28420,N_27490,N_27240);
nand U28421 (N_28421,N_27030,N_27574);
nand U28422 (N_28422,N_27775,N_27262);
xor U28423 (N_28423,N_27808,N_27861);
and U28424 (N_28424,N_27897,N_27053);
and U28425 (N_28425,N_27953,N_27533);
nor U28426 (N_28426,N_27074,N_27984);
nand U28427 (N_28427,N_27684,N_27344);
nor U28428 (N_28428,N_27634,N_27599);
nand U28429 (N_28429,N_27183,N_27656);
nand U28430 (N_28430,N_27410,N_27079);
nand U28431 (N_28431,N_27065,N_27043);
or U28432 (N_28432,N_27592,N_27755);
xor U28433 (N_28433,N_27517,N_27164);
xor U28434 (N_28434,N_27476,N_27624);
xnor U28435 (N_28435,N_27519,N_27720);
or U28436 (N_28436,N_27145,N_27394);
and U28437 (N_28437,N_27238,N_27033);
xnor U28438 (N_28438,N_27372,N_27105);
xnor U28439 (N_28439,N_27862,N_27765);
and U28440 (N_28440,N_27382,N_27587);
xnor U28441 (N_28441,N_27093,N_27942);
and U28442 (N_28442,N_27334,N_27538);
xnor U28443 (N_28443,N_27857,N_27855);
or U28444 (N_28444,N_27312,N_27287);
and U28445 (N_28445,N_27737,N_27895);
nor U28446 (N_28446,N_27286,N_27815);
nand U28447 (N_28447,N_27706,N_27838);
nand U28448 (N_28448,N_27037,N_27260);
nand U28449 (N_28449,N_27028,N_27764);
and U28450 (N_28450,N_27171,N_27011);
xor U28451 (N_28451,N_27444,N_27948);
xnor U28452 (N_28452,N_27007,N_27723);
nor U28453 (N_28453,N_27157,N_27938);
nor U28454 (N_28454,N_27625,N_27831);
and U28455 (N_28455,N_27785,N_27090);
or U28456 (N_28456,N_27666,N_27248);
and U28457 (N_28457,N_27454,N_27450);
nor U28458 (N_28458,N_27134,N_27983);
nor U28459 (N_28459,N_27274,N_27207);
and U28460 (N_28460,N_27395,N_27040);
nor U28461 (N_28461,N_27554,N_27722);
or U28462 (N_28462,N_27550,N_27792);
xnor U28463 (N_28463,N_27430,N_27421);
and U28464 (N_28464,N_27278,N_27133);
and U28465 (N_28465,N_27012,N_27411);
and U28466 (N_28466,N_27796,N_27288);
nor U28467 (N_28467,N_27348,N_27511);
xor U28468 (N_28468,N_27629,N_27310);
and U28469 (N_28469,N_27875,N_27422);
and U28470 (N_28470,N_27910,N_27670);
xor U28471 (N_28471,N_27241,N_27899);
nand U28472 (N_28472,N_27655,N_27890);
and U28473 (N_28473,N_27918,N_27508);
nand U28474 (N_28474,N_27399,N_27681);
nor U28475 (N_28475,N_27413,N_27329);
and U28476 (N_28476,N_27077,N_27232);
or U28477 (N_28477,N_27958,N_27066);
nor U28478 (N_28478,N_27180,N_27097);
nand U28479 (N_28479,N_27390,N_27545);
nor U28480 (N_28480,N_27493,N_27213);
xor U28481 (N_28481,N_27615,N_27088);
or U28482 (N_28482,N_27864,N_27301);
or U28483 (N_28483,N_27752,N_27346);
nor U28484 (N_28484,N_27022,N_27523);
xnor U28485 (N_28485,N_27849,N_27257);
nor U28486 (N_28486,N_27821,N_27474);
or U28487 (N_28487,N_27593,N_27633);
or U28488 (N_28488,N_27541,N_27901);
xor U28489 (N_28489,N_27230,N_27300);
nand U28490 (N_28490,N_27483,N_27143);
nor U28491 (N_28491,N_27707,N_27169);
and U28492 (N_28492,N_27050,N_27386);
and U28493 (N_28493,N_27487,N_27185);
and U28494 (N_28494,N_27691,N_27081);
and U28495 (N_28495,N_27485,N_27973);
xnor U28496 (N_28496,N_27687,N_27643);
nand U28497 (N_28497,N_27816,N_27255);
nand U28498 (N_28498,N_27202,N_27405);
nand U28499 (N_28499,N_27912,N_27518);
and U28500 (N_28500,N_27788,N_27520);
and U28501 (N_28501,N_27525,N_27127);
and U28502 (N_28502,N_27681,N_27570);
nand U28503 (N_28503,N_27964,N_27147);
xor U28504 (N_28504,N_27739,N_27547);
nand U28505 (N_28505,N_27099,N_27953);
nand U28506 (N_28506,N_27951,N_27528);
or U28507 (N_28507,N_27263,N_27256);
nor U28508 (N_28508,N_27869,N_27366);
or U28509 (N_28509,N_27612,N_27555);
or U28510 (N_28510,N_27594,N_27510);
or U28511 (N_28511,N_27744,N_27785);
nand U28512 (N_28512,N_27829,N_27664);
nor U28513 (N_28513,N_27950,N_27214);
or U28514 (N_28514,N_27068,N_27020);
or U28515 (N_28515,N_27575,N_27288);
nand U28516 (N_28516,N_27398,N_27870);
nand U28517 (N_28517,N_27057,N_27290);
xnor U28518 (N_28518,N_27155,N_27544);
nand U28519 (N_28519,N_27015,N_27124);
nor U28520 (N_28520,N_27722,N_27131);
xnor U28521 (N_28521,N_27126,N_27501);
xnor U28522 (N_28522,N_27750,N_27139);
or U28523 (N_28523,N_27845,N_27627);
nor U28524 (N_28524,N_27955,N_27304);
and U28525 (N_28525,N_27093,N_27487);
or U28526 (N_28526,N_27712,N_27746);
and U28527 (N_28527,N_27018,N_27900);
nand U28528 (N_28528,N_27796,N_27978);
and U28529 (N_28529,N_27935,N_27566);
or U28530 (N_28530,N_27718,N_27507);
or U28531 (N_28531,N_27717,N_27524);
nor U28532 (N_28532,N_27251,N_27775);
nand U28533 (N_28533,N_27907,N_27559);
nor U28534 (N_28534,N_27358,N_27858);
or U28535 (N_28535,N_27054,N_27097);
xor U28536 (N_28536,N_27361,N_27919);
and U28537 (N_28537,N_27848,N_27836);
and U28538 (N_28538,N_27582,N_27617);
and U28539 (N_28539,N_27139,N_27086);
xnor U28540 (N_28540,N_27427,N_27490);
nand U28541 (N_28541,N_27087,N_27304);
xor U28542 (N_28542,N_27421,N_27903);
nand U28543 (N_28543,N_27921,N_27890);
and U28544 (N_28544,N_27892,N_27062);
nand U28545 (N_28545,N_27584,N_27892);
nand U28546 (N_28546,N_27815,N_27582);
nand U28547 (N_28547,N_27338,N_27815);
and U28548 (N_28548,N_27495,N_27425);
nand U28549 (N_28549,N_27702,N_27413);
nand U28550 (N_28550,N_27838,N_27261);
nor U28551 (N_28551,N_27166,N_27655);
and U28552 (N_28552,N_27606,N_27600);
xor U28553 (N_28553,N_27756,N_27373);
nor U28554 (N_28554,N_27601,N_27970);
nand U28555 (N_28555,N_27038,N_27272);
or U28556 (N_28556,N_27940,N_27188);
and U28557 (N_28557,N_27081,N_27398);
xor U28558 (N_28558,N_27401,N_27433);
nor U28559 (N_28559,N_27331,N_27268);
nand U28560 (N_28560,N_27534,N_27928);
or U28561 (N_28561,N_27780,N_27801);
and U28562 (N_28562,N_27893,N_27525);
nor U28563 (N_28563,N_27102,N_27018);
xor U28564 (N_28564,N_27817,N_27604);
xnor U28565 (N_28565,N_27850,N_27959);
and U28566 (N_28566,N_27791,N_27141);
nor U28567 (N_28567,N_27815,N_27528);
nor U28568 (N_28568,N_27023,N_27466);
xor U28569 (N_28569,N_27041,N_27012);
nor U28570 (N_28570,N_27769,N_27719);
and U28571 (N_28571,N_27591,N_27684);
nand U28572 (N_28572,N_27263,N_27493);
nor U28573 (N_28573,N_27709,N_27118);
and U28574 (N_28574,N_27535,N_27465);
or U28575 (N_28575,N_27734,N_27153);
nor U28576 (N_28576,N_27862,N_27222);
and U28577 (N_28577,N_27694,N_27340);
and U28578 (N_28578,N_27445,N_27010);
nand U28579 (N_28579,N_27639,N_27185);
xnor U28580 (N_28580,N_27406,N_27466);
nand U28581 (N_28581,N_27889,N_27335);
xnor U28582 (N_28582,N_27298,N_27544);
nor U28583 (N_28583,N_27939,N_27618);
nor U28584 (N_28584,N_27902,N_27009);
nand U28585 (N_28585,N_27607,N_27878);
or U28586 (N_28586,N_27807,N_27848);
and U28587 (N_28587,N_27615,N_27855);
nand U28588 (N_28588,N_27523,N_27909);
nand U28589 (N_28589,N_27438,N_27189);
and U28590 (N_28590,N_27653,N_27114);
xnor U28591 (N_28591,N_27291,N_27281);
or U28592 (N_28592,N_27853,N_27194);
nor U28593 (N_28593,N_27781,N_27121);
and U28594 (N_28594,N_27885,N_27812);
or U28595 (N_28595,N_27678,N_27084);
and U28596 (N_28596,N_27474,N_27927);
xnor U28597 (N_28597,N_27005,N_27190);
nand U28598 (N_28598,N_27832,N_27849);
and U28599 (N_28599,N_27479,N_27017);
and U28600 (N_28600,N_27899,N_27692);
xor U28601 (N_28601,N_27093,N_27637);
or U28602 (N_28602,N_27492,N_27009);
or U28603 (N_28603,N_27026,N_27578);
and U28604 (N_28604,N_27930,N_27719);
nand U28605 (N_28605,N_27101,N_27889);
or U28606 (N_28606,N_27388,N_27916);
or U28607 (N_28607,N_27827,N_27286);
or U28608 (N_28608,N_27966,N_27667);
and U28609 (N_28609,N_27538,N_27679);
or U28610 (N_28610,N_27712,N_27622);
xor U28611 (N_28611,N_27788,N_27040);
nand U28612 (N_28612,N_27280,N_27749);
and U28613 (N_28613,N_27044,N_27975);
and U28614 (N_28614,N_27533,N_27152);
and U28615 (N_28615,N_27274,N_27943);
or U28616 (N_28616,N_27421,N_27186);
and U28617 (N_28617,N_27545,N_27735);
nand U28618 (N_28618,N_27831,N_27766);
and U28619 (N_28619,N_27842,N_27616);
or U28620 (N_28620,N_27441,N_27831);
xor U28621 (N_28621,N_27587,N_27267);
nand U28622 (N_28622,N_27373,N_27737);
nand U28623 (N_28623,N_27519,N_27275);
and U28624 (N_28624,N_27747,N_27868);
or U28625 (N_28625,N_27120,N_27492);
nand U28626 (N_28626,N_27393,N_27843);
nor U28627 (N_28627,N_27151,N_27566);
or U28628 (N_28628,N_27065,N_27138);
and U28629 (N_28629,N_27628,N_27299);
and U28630 (N_28630,N_27263,N_27799);
or U28631 (N_28631,N_27150,N_27215);
xnor U28632 (N_28632,N_27680,N_27815);
nor U28633 (N_28633,N_27534,N_27324);
nand U28634 (N_28634,N_27916,N_27450);
nand U28635 (N_28635,N_27139,N_27688);
xnor U28636 (N_28636,N_27066,N_27427);
xor U28637 (N_28637,N_27458,N_27472);
and U28638 (N_28638,N_27886,N_27081);
or U28639 (N_28639,N_27212,N_27395);
nor U28640 (N_28640,N_27658,N_27604);
or U28641 (N_28641,N_27080,N_27485);
and U28642 (N_28642,N_27987,N_27048);
nand U28643 (N_28643,N_27514,N_27820);
or U28644 (N_28644,N_27777,N_27421);
nand U28645 (N_28645,N_27872,N_27521);
nor U28646 (N_28646,N_27437,N_27917);
or U28647 (N_28647,N_27359,N_27486);
nand U28648 (N_28648,N_27576,N_27727);
or U28649 (N_28649,N_27448,N_27765);
and U28650 (N_28650,N_27719,N_27362);
or U28651 (N_28651,N_27257,N_27782);
and U28652 (N_28652,N_27622,N_27432);
xnor U28653 (N_28653,N_27440,N_27079);
and U28654 (N_28654,N_27644,N_27385);
xnor U28655 (N_28655,N_27830,N_27025);
nor U28656 (N_28656,N_27840,N_27302);
nand U28657 (N_28657,N_27439,N_27837);
nor U28658 (N_28658,N_27562,N_27536);
xnor U28659 (N_28659,N_27398,N_27482);
nor U28660 (N_28660,N_27757,N_27713);
or U28661 (N_28661,N_27705,N_27402);
xnor U28662 (N_28662,N_27478,N_27438);
nand U28663 (N_28663,N_27333,N_27247);
and U28664 (N_28664,N_27471,N_27781);
nor U28665 (N_28665,N_27100,N_27732);
or U28666 (N_28666,N_27780,N_27730);
xor U28667 (N_28667,N_27762,N_27883);
or U28668 (N_28668,N_27179,N_27353);
nor U28669 (N_28669,N_27996,N_27434);
or U28670 (N_28670,N_27382,N_27118);
nand U28671 (N_28671,N_27233,N_27085);
and U28672 (N_28672,N_27803,N_27725);
xor U28673 (N_28673,N_27520,N_27065);
xnor U28674 (N_28674,N_27167,N_27657);
and U28675 (N_28675,N_27378,N_27253);
xor U28676 (N_28676,N_27635,N_27974);
or U28677 (N_28677,N_27687,N_27041);
or U28678 (N_28678,N_27414,N_27223);
xnor U28679 (N_28679,N_27974,N_27680);
xor U28680 (N_28680,N_27834,N_27385);
or U28681 (N_28681,N_27415,N_27510);
xor U28682 (N_28682,N_27252,N_27294);
xor U28683 (N_28683,N_27480,N_27056);
xnor U28684 (N_28684,N_27348,N_27061);
nor U28685 (N_28685,N_27647,N_27903);
or U28686 (N_28686,N_27945,N_27030);
and U28687 (N_28687,N_27531,N_27644);
xor U28688 (N_28688,N_27203,N_27136);
nand U28689 (N_28689,N_27202,N_27277);
nor U28690 (N_28690,N_27808,N_27722);
or U28691 (N_28691,N_27308,N_27210);
and U28692 (N_28692,N_27287,N_27838);
and U28693 (N_28693,N_27128,N_27433);
or U28694 (N_28694,N_27455,N_27632);
or U28695 (N_28695,N_27180,N_27448);
and U28696 (N_28696,N_27956,N_27057);
xnor U28697 (N_28697,N_27137,N_27995);
nor U28698 (N_28698,N_27334,N_27917);
and U28699 (N_28699,N_27171,N_27759);
and U28700 (N_28700,N_27406,N_27996);
nand U28701 (N_28701,N_27778,N_27022);
xnor U28702 (N_28702,N_27934,N_27114);
nor U28703 (N_28703,N_27680,N_27739);
xnor U28704 (N_28704,N_27835,N_27430);
and U28705 (N_28705,N_27022,N_27573);
or U28706 (N_28706,N_27802,N_27966);
and U28707 (N_28707,N_27619,N_27002);
and U28708 (N_28708,N_27737,N_27636);
and U28709 (N_28709,N_27649,N_27615);
nand U28710 (N_28710,N_27258,N_27848);
nor U28711 (N_28711,N_27442,N_27304);
nand U28712 (N_28712,N_27057,N_27945);
or U28713 (N_28713,N_27568,N_27786);
or U28714 (N_28714,N_27839,N_27458);
and U28715 (N_28715,N_27644,N_27186);
or U28716 (N_28716,N_27626,N_27230);
or U28717 (N_28717,N_27436,N_27702);
xnor U28718 (N_28718,N_27863,N_27107);
nor U28719 (N_28719,N_27353,N_27186);
or U28720 (N_28720,N_27191,N_27731);
and U28721 (N_28721,N_27147,N_27723);
or U28722 (N_28722,N_27685,N_27574);
or U28723 (N_28723,N_27383,N_27262);
and U28724 (N_28724,N_27978,N_27367);
xnor U28725 (N_28725,N_27213,N_27637);
or U28726 (N_28726,N_27541,N_27282);
nor U28727 (N_28727,N_27502,N_27583);
or U28728 (N_28728,N_27886,N_27757);
and U28729 (N_28729,N_27219,N_27448);
nand U28730 (N_28730,N_27664,N_27246);
nor U28731 (N_28731,N_27054,N_27186);
nor U28732 (N_28732,N_27288,N_27512);
nand U28733 (N_28733,N_27464,N_27895);
and U28734 (N_28734,N_27047,N_27360);
xnor U28735 (N_28735,N_27444,N_27764);
nor U28736 (N_28736,N_27900,N_27970);
nor U28737 (N_28737,N_27015,N_27307);
or U28738 (N_28738,N_27290,N_27732);
nand U28739 (N_28739,N_27226,N_27217);
xnor U28740 (N_28740,N_27546,N_27093);
or U28741 (N_28741,N_27535,N_27977);
nor U28742 (N_28742,N_27929,N_27549);
xor U28743 (N_28743,N_27919,N_27343);
nand U28744 (N_28744,N_27991,N_27186);
and U28745 (N_28745,N_27855,N_27786);
nand U28746 (N_28746,N_27250,N_27010);
or U28747 (N_28747,N_27961,N_27700);
and U28748 (N_28748,N_27341,N_27707);
xor U28749 (N_28749,N_27914,N_27158);
xnor U28750 (N_28750,N_27056,N_27844);
or U28751 (N_28751,N_27749,N_27628);
and U28752 (N_28752,N_27738,N_27838);
nand U28753 (N_28753,N_27714,N_27557);
nand U28754 (N_28754,N_27697,N_27644);
nand U28755 (N_28755,N_27307,N_27715);
xnor U28756 (N_28756,N_27550,N_27273);
xor U28757 (N_28757,N_27480,N_27436);
nand U28758 (N_28758,N_27444,N_27277);
and U28759 (N_28759,N_27878,N_27866);
nand U28760 (N_28760,N_27060,N_27355);
or U28761 (N_28761,N_27250,N_27923);
nor U28762 (N_28762,N_27930,N_27089);
and U28763 (N_28763,N_27777,N_27334);
and U28764 (N_28764,N_27967,N_27548);
nand U28765 (N_28765,N_27771,N_27504);
or U28766 (N_28766,N_27958,N_27514);
and U28767 (N_28767,N_27978,N_27771);
xnor U28768 (N_28768,N_27441,N_27613);
and U28769 (N_28769,N_27503,N_27725);
nand U28770 (N_28770,N_27617,N_27774);
or U28771 (N_28771,N_27592,N_27585);
and U28772 (N_28772,N_27873,N_27144);
and U28773 (N_28773,N_27030,N_27466);
nor U28774 (N_28774,N_27634,N_27990);
xnor U28775 (N_28775,N_27004,N_27773);
and U28776 (N_28776,N_27874,N_27849);
or U28777 (N_28777,N_27107,N_27144);
and U28778 (N_28778,N_27463,N_27251);
and U28779 (N_28779,N_27937,N_27348);
nor U28780 (N_28780,N_27119,N_27945);
nor U28781 (N_28781,N_27309,N_27454);
or U28782 (N_28782,N_27595,N_27893);
or U28783 (N_28783,N_27427,N_27017);
nand U28784 (N_28784,N_27088,N_27229);
and U28785 (N_28785,N_27872,N_27206);
or U28786 (N_28786,N_27455,N_27170);
and U28787 (N_28787,N_27520,N_27929);
nor U28788 (N_28788,N_27587,N_27153);
nand U28789 (N_28789,N_27100,N_27425);
xor U28790 (N_28790,N_27160,N_27334);
and U28791 (N_28791,N_27287,N_27773);
xor U28792 (N_28792,N_27469,N_27554);
nor U28793 (N_28793,N_27069,N_27530);
nand U28794 (N_28794,N_27604,N_27303);
nor U28795 (N_28795,N_27600,N_27475);
or U28796 (N_28796,N_27419,N_27094);
or U28797 (N_28797,N_27417,N_27191);
or U28798 (N_28798,N_27226,N_27247);
nor U28799 (N_28799,N_27609,N_27488);
nor U28800 (N_28800,N_27212,N_27454);
nor U28801 (N_28801,N_27990,N_27115);
or U28802 (N_28802,N_27271,N_27984);
or U28803 (N_28803,N_27473,N_27565);
nor U28804 (N_28804,N_27365,N_27167);
xnor U28805 (N_28805,N_27767,N_27647);
nor U28806 (N_28806,N_27435,N_27184);
and U28807 (N_28807,N_27545,N_27771);
xor U28808 (N_28808,N_27331,N_27006);
xor U28809 (N_28809,N_27745,N_27861);
xnor U28810 (N_28810,N_27251,N_27133);
or U28811 (N_28811,N_27143,N_27686);
xnor U28812 (N_28812,N_27508,N_27775);
nor U28813 (N_28813,N_27050,N_27466);
or U28814 (N_28814,N_27231,N_27248);
or U28815 (N_28815,N_27313,N_27498);
nand U28816 (N_28816,N_27590,N_27878);
nor U28817 (N_28817,N_27567,N_27171);
or U28818 (N_28818,N_27529,N_27203);
nand U28819 (N_28819,N_27875,N_27471);
xor U28820 (N_28820,N_27883,N_27323);
nor U28821 (N_28821,N_27944,N_27534);
nand U28822 (N_28822,N_27014,N_27788);
or U28823 (N_28823,N_27132,N_27602);
and U28824 (N_28824,N_27289,N_27740);
nand U28825 (N_28825,N_27565,N_27378);
nor U28826 (N_28826,N_27668,N_27665);
and U28827 (N_28827,N_27291,N_27190);
and U28828 (N_28828,N_27638,N_27061);
nor U28829 (N_28829,N_27255,N_27386);
nand U28830 (N_28830,N_27319,N_27412);
and U28831 (N_28831,N_27887,N_27685);
nor U28832 (N_28832,N_27649,N_27618);
nand U28833 (N_28833,N_27549,N_27308);
nand U28834 (N_28834,N_27933,N_27815);
and U28835 (N_28835,N_27289,N_27670);
and U28836 (N_28836,N_27060,N_27576);
nor U28837 (N_28837,N_27380,N_27348);
xnor U28838 (N_28838,N_27633,N_27194);
nor U28839 (N_28839,N_27186,N_27823);
and U28840 (N_28840,N_27351,N_27384);
or U28841 (N_28841,N_27276,N_27453);
or U28842 (N_28842,N_27624,N_27310);
or U28843 (N_28843,N_27511,N_27953);
and U28844 (N_28844,N_27371,N_27040);
nand U28845 (N_28845,N_27476,N_27010);
xnor U28846 (N_28846,N_27170,N_27964);
xnor U28847 (N_28847,N_27505,N_27586);
or U28848 (N_28848,N_27666,N_27926);
nand U28849 (N_28849,N_27550,N_27764);
xnor U28850 (N_28850,N_27967,N_27776);
xor U28851 (N_28851,N_27868,N_27385);
nor U28852 (N_28852,N_27221,N_27539);
nand U28853 (N_28853,N_27689,N_27546);
and U28854 (N_28854,N_27229,N_27827);
and U28855 (N_28855,N_27444,N_27382);
nor U28856 (N_28856,N_27386,N_27614);
or U28857 (N_28857,N_27321,N_27344);
xor U28858 (N_28858,N_27453,N_27389);
and U28859 (N_28859,N_27861,N_27322);
and U28860 (N_28860,N_27034,N_27080);
nor U28861 (N_28861,N_27328,N_27528);
nor U28862 (N_28862,N_27545,N_27309);
or U28863 (N_28863,N_27108,N_27931);
nor U28864 (N_28864,N_27869,N_27292);
xnor U28865 (N_28865,N_27182,N_27165);
xnor U28866 (N_28866,N_27132,N_27362);
or U28867 (N_28867,N_27740,N_27864);
xor U28868 (N_28868,N_27339,N_27741);
xor U28869 (N_28869,N_27766,N_27258);
xnor U28870 (N_28870,N_27697,N_27707);
or U28871 (N_28871,N_27309,N_27499);
xor U28872 (N_28872,N_27522,N_27214);
nand U28873 (N_28873,N_27219,N_27251);
xor U28874 (N_28874,N_27883,N_27387);
nand U28875 (N_28875,N_27005,N_27434);
or U28876 (N_28876,N_27160,N_27260);
nand U28877 (N_28877,N_27446,N_27696);
xor U28878 (N_28878,N_27304,N_27066);
nand U28879 (N_28879,N_27847,N_27321);
nor U28880 (N_28880,N_27662,N_27856);
nand U28881 (N_28881,N_27511,N_27699);
or U28882 (N_28882,N_27270,N_27600);
xor U28883 (N_28883,N_27600,N_27202);
or U28884 (N_28884,N_27250,N_27482);
xor U28885 (N_28885,N_27556,N_27510);
and U28886 (N_28886,N_27629,N_27624);
nor U28887 (N_28887,N_27772,N_27978);
nor U28888 (N_28888,N_27492,N_27797);
xnor U28889 (N_28889,N_27396,N_27567);
or U28890 (N_28890,N_27567,N_27647);
nor U28891 (N_28891,N_27942,N_27439);
nand U28892 (N_28892,N_27858,N_27559);
xor U28893 (N_28893,N_27924,N_27177);
nor U28894 (N_28894,N_27845,N_27010);
nor U28895 (N_28895,N_27636,N_27480);
xor U28896 (N_28896,N_27099,N_27915);
nor U28897 (N_28897,N_27655,N_27681);
nor U28898 (N_28898,N_27408,N_27392);
nand U28899 (N_28899,N_27198,N_27484);
nor U28900 (N_28900,N_27392,N_27875);
xor U28901 (N_28901,N_27128,N_27470);
or U28902 (N_28902,N_27936,N_27478);
and U28903 (N_28903,N_27620,N_27571);
nand U28904 (N_28904,N_27384,N_27527);
nand U28905 (N_28905,N_27332,N_27441);
or U28906 (N_28906,N_27926,N_27624);
or U28907 (N_28907,N_27178,N_27802);
xnor U28908 (N_28908,N_27698,N_27675);
nand U28909 (N_28909,N_27249,N_27053);
xor U28910 (N_28910,N_27576,N_27209);
or U28911 (N_28911,N_27260,N_27998);
xnor U28912 (N_28912,N_27860,N_27389);
or U28913 (N_28913,N_27079,N_27357);
xnor U28914 (N_28914,N_27833,N_27043);
nor U28915 (N_28915,N_27609,N_27588);
or U28916 (N_28916,N_27226,N_27118);
or U28917 (N_28917,N_27298,N_27543);
nand U28918 (N_28918,N_27205,N_27929);
and U28919 (N_28919,N_27111,N_27062);
or U28920 (N_28920,N_27567,N_27392);
or U28921 (N_28921,N_27651,N_27771);
nand U28922 (N_28922,N_27851,N_27829);
and U28923 (N_28923,N_27198,N_27820);
and U28924 (N_28924,N_27979,N_27178);
nand U28925 (N_28925,N_27908,N_27276);
xnor U28926 (N_28926,N_27925,N_27716);
nand U28927 (N_28927,N_27755,N_27822);
and U28928 (N_28928,N_27487,N_27603);
nor U28929 (N_28929,N_27167,N_27635);
nand U28930 (N_28930,N_27379,N_27221);
or U28931 (N_28931,N_27555,N_27426);
nor U28932 (N_28932,N_27423,N_27831);
xor U28933 (N_28933,N_27808,N_27434);
or U28934 (N_28934,N_27256,N_27942);
and U28935 (N_28935,N_27395,N_27525);
and U28936 (N_28936,N_27843,N_27230);
xnor U28937 (N_28937,N_27767,N_27853);
nand U28938 (N_28938,N_27878,N_27531);
or U28939 (N_28939,N_27016,N_27933);
nor U28940 (N_28940,N_27348,N_27831);
xnor U28941 (N_28941,N_27148,N_27427);
nand U28942 (N_28942,N_27791,N_27744);
nand U28943 (N_28943,N_27382,N_27860);
nand U28944 (N_28944,N_27975,N_27498);
or U28945 (N_28945,N_27773,N_27008);
xor U28946 (N_28946,N_27558,N_27410);
xor U28947 (N_28947,N_27431,N_27641);
nand U28948 (N_28948,N_27115,N_27823);
and U28949 (N_28949,N_27034,N_27375);
nor U28950 (N_28950,N_27935,N_27652);
nor U28951 (N_28951,N_27125,N_27804);
nor U28952 (N_28952,N_27000,N_27594);
nor U28953 (N_28953,N_27803,N_27756);
nor U28954 (N_28954,N_27372,N_27885);
nand U28955 (N_28955,N_27161,N_27844);
or U28956 (N_28956,N_27110,N_27551);
or U28957 (N_28957,N_27294,N_27906);
nor U28958 (N_28958,N_27081,N_27294);
xor U28959 (N_28959,N_27557,N_27303);
nor U28960 (N_28960,N_27713,N_27404);
nor U28961 (N_28961,N_27953,N_27571);
xor U28962 (N_28962,N_27152,N_27766);
nand U28963 (N_28963,N_27142,N_27874);
or U28964 (N_28964,N_27797,N_27413);
and U28965 (N_28965,N_27119,N_27684);
nand U28966 (N_28966,N_27374,N_27832);
nand U28967 (N_28967,N_27797,N_27479);
or U28968 (N_28968,N_27653,N_27746);
nor U28969 (N_28969,N_27294,N_27026);
nand U28970 (N_28970,N_27788,N_27277);
nor U28971 (N_28971,N_27878,N_27387);
nand U28972 (N_28972,N_27397,N_27131);
and U28973 (N_28973,N_27044,N_27180);
nor U28974 (N_28974,N_27018,N_27329);
xnor U28975 (N_28975,N_27428,N_27643);
nand U28976 (N_28976,N_27767,N_27352);
xnor U28977 (N_28977,N_27335,N_27325);
xnor U28978 (N_28978,N_27483,N_27360);
or U28979 (N_28979,N_27680,N_27066);
nor U28980 (N_28980,N_27716,N_27040);
or U28981 (N_28981,N_27128,N_27068);
nand U28982 (N_28982,N_27739,N_27029);
nor U28983 (N_28983,N_27660,N_27645);
nand U28984 (N_28984,N_27601,N_27673);
xor U28985 (N_28985,N_27318,N_27365);
or U28986 (N_28986,N_27787,N_27291);
nand U28987 (N_28987,N_27642,N_27609);
or U28988 (N_28988,N_27619,N_27167);
nor U28989 (N_28989,N_27592,N_27732);
nor U28990 (N_28990,N_27567,N_27600);
nor U28991 (N_28991,N_27960,N_27559);
nor U28992 (N_28992,N_27548,N_27970);
nor U28993 (N_28993,N_27541,N_27870);
xor U28994 (N_28994,N_27359,N_27295);
nor U28995 (N_28995,N_27388,N_27836);
nand U28996 (N_28996,N_27735,N_27482);
and U28997 (N_28997,N_27546,N_27675);
nand U28998 (N_28998,N_27357,N_27626);
or U28999 (N_28999,N_27023,N_27749);
and U29000 (N_29000,N_28701,N_28033);
nand U29001 (N_29001,N_28844,N_28586);
or U29002 (N_29002,N_28362,N_28029);
xor U29003 (N_29003,N_28183,N_28386);
nand U29004 (N_29004,N_28443,N_28768);
xor U29005 (N_29005,N_28621,N_28648);
nand U29006 (N_29006,N_28470,N_28451);
and U29007 (N_29007,N_28378,N_28323);
nor U29008 (N_29008,N_28619,N_28208);
nand U29009 (N_29009,N_28352,N_28391);
xnor U29010 (N_29010,N_28248,N_28992);
xor U29011 (N_29011,N_28583,N_28004);
and U29012 (N_29012,N_28698,N_28271);
nor U29013 (N_29013,N_28978,N_28186);
nand U29014 (N_29014,N_28348,N_28440);
or U29015 (N_29015,N_28150,N_28224);
or U29016 (N_29016,N_28901,N_28730);
xor U29017 (N_29017,N_28760,N_28260);
or U29018 (N_29018,N_28141,N_28840);
nor U29019 (N_29019,N_28708,N_28337);
nor U29020 (N_29020,N_28924,N_28031);
nand U29021 (N_29021,N_28842,N_28410);
or U29022 (N_29022,N_28125,N_28811);
nor U29023 (N_29023,N_28177,N_28776);
nand U29024 (N_29024,N_28148,N_28514);
nand U29025 (N_29025,N_28759,N_28839);
nand U29026 (N_29026,N_28302,N_28088);
xor U29027 (N_29027,N_28555,N_28489);
and U29028 (N_29028,N_28116,N_28762);
or U29029 (N_29029,N_28441,N_28749);
or U29030 (N_29030,N_28895,N_28641);
or U29031 (N_29031,N_28301,N_28794);
nand U29032 (N_29032,N_28676,N_28098);
nor U29033 (N_29033,N_28674,N_28020);
nand U29034 (N_29034,N_28897,N_28190);
and U29035 (N_29035,N_28015,N_28457);
or U29036 (N_29036,N_28905,N_28539);
nand U29037 (N_29037,N_28994,N_28615);
nand U29038 (N_29038,N_28587,N_28649);
xor U29039 (N_29039,N_28932,N_28739);
or U29040 (N_29040,N_28351,N_28767);
nor U29041 (N_29041,N_28949,N_28120);
nand U29042 (N_29042,N_28423,N_28666);
nand U29043 (N_29043,N_28947,N_28406);
nor U29044 (N_29044,N_28538,N_28564);
xnor U29045 (N_29045,N_28044,N_28558);
nor U29046 (N_29046,N_28919,N_28741);
nor U29047 (N_29047,N_28228,N_28569);
and U29048 (N_29048,N_28075,N_28926);
nor U29049 (N_29049,N_28213,N_28163);
xnor U29050 (N_29050,N_28403,N_28934);
xor U29051 (N_29051,N_28529,N_28182);
or U29052 (N_29052,N_28883,N_28609);
nor U29053 (N_29053,N_28942,N_28707);
xor U29054 (N_29054,N_28474,N_28589);
xnor U29055 (N_29055,N_28624,N_28900);
nor U29056 (N_29056,N_28812,N_28252);
and U29057 (N_29057,N_28039,N_28719);
and U29058 (N_29058,N_28726,N_28801);
or U29059 (N_29059,N_28548,N_28304);
nor U29060 (N_29060,N_28368,N_28953);
and U29061 (N_29061,N_28625,N_28736);
and U29062 (N_29062,N_28052,N_28399);
xor U29063 (N_29063,N_28518,N_28392);
nor U29064 (N_29064,N_28479,N_28508);
or U29065 (N_29065,N_28353,N_28076);
nor U29066 (N_29066,N_28772,N_28294);
nand U29067 (N_29067,N_28197,N_28357);
and U29068 (N_29068,N_28180,N_28439);
nor U29069 (N_29069,N_28500,N_28251);
nand U29070 (N_29070,N_28086,N_28981);
nand U29071 (N_29071,N_28792,N_28887);
xnor U29072 (N_29072,N_28258,N_28178);
nand U29073 (N_29073,N_28712,N_28280);
or U29074 (N_29074,N_28857,N_28774);
or U29075 (N_29075,N_28940,N_28402);
xor U29076 (N_29076,N_28255,N_28018);
nand U29077 (N_29077,N_28988,N_28911);
xor U29078 (N_29078,N_28702,N_28331);
or U29079 (N_29079,N_28377,N_28892);
or U29080 (N_29080,N_28700,N_28841);
or U29081 (N_29081,N_28893,N_28639);
and U29082 (N_29082,N_28101,N_28541);
or U29083 (N_29083,N_28425,N_28413);
and U29084 (N_29084,N_28724,N_28172);
xnor U29085 (N_29085,N_28584,N_28979);
nand U29086 (N_29086,N_28626,N_28788);
or U29087 (N_29087,N_28685,N_28671);
and U29088 (N_29088,N_28480,N_28446);
nand U29089 (N_29089,N_28318,N_28972);
xnor U29090 (N_29090,N_28153,N_28689);
or U29091 (N_29091,N_28176,N_28114);
nand U29092 (N_29092,N_28567,N_28537);
xnor U29093 (N_29093,N_28536,N_28313);
or U29094 (N_29094,N_28611,N_28886);
and U29095 (N_29095,N_28281,N_28613);
or U29096 (N_29096,N_28214,N_28206);
and U29097 (N_29097,N_28967,N_28960);
nand U29098 (N_29098,N_28291,N_28598);
nor U29099 (N_29099,N_28217,N_28123);
and U29100 (N_29100,N_28709,N_28264);
nor U29101 (N_29101,N_28814,N_28503);
and U29102 (N_29102,N_28372,N_28243);
or U29103 (N_29103,N_28417,N_28327);
and U29104 (N_29104,N_28822,N_28491);
or U29105 (N_29105,N_28629,N_28297);
xnor U29106 (N_29106,N_28232,N_28665);
nand U29107 (N_29107,N_28115,N_28209);
and U29108 (N_29108,N_28927,N_28531);
xor U29109 (N_29109,N_28225,N_28999);
xor U29110 (N_29110,N_28092,N_28546);
or U29111 (N_29111,N_28442,N_28469);
nor U29112 (N_29112,N_28129,N_28504);
and U29113 (N_29113,N_28156,N_28882);
xor U29114 (N_29114,N_28493,N_28340);
nor U29115 (N_29115,N_28652,N_28219);
xnor U29116 (N_29116,N_28144,N_28202);
nand U29117 (N_29117,N_28963,N_28663);
nand U29118 (N_29118,N_28694,N_28600);
xor U29119 (N_29119,N_28390,N_28863);
and U29120 (N_29120,N_28102,N_28152);
nor U29121 (N_29121,N_28053,N_28916);
xor U29122 (N_29122,N_28132,N_28850);
and U29123 (N_29123,N_28454,N_28941);
nand U29124 (N_29124,N_28317,N_28985);
and U29125 (N_29125,N_28644,N_28881);
or U29126 (N_29126,N_28358,N_28046);
and U29127 (N_29127,N_28211,N_28904);
nand U29128 (N_29128,N_28010,N_28827);
and U29129 (N_29129,N_28041,N_28025);
or U29130 (N_29130,N_28521,N_28055);
and U29131 (N_29131,N_28745,N_28743);
xor U29132 (N_29132,N_28912,N_28687);
nand U29133 (N_29133,N_28732,N_28858);
nor U29134 (N_29134,N_28710,N_28220);
or U29135 (N_29135,N_28865,N_28030);
xnor U29136 (N_29136,N_28133,N_28173);
nor U29137 (N_29137,N_28171,N_28524);
xor U29138 (N_29138,N_28825,N_28717);
or U29139 (N_29139,N_28049,N_28917);
nor U29140 (N_29140,N_28240,N_28166);
nor U29141 (N_29141,N_28433,N_28022);
or U29142 (N_29142,N_28308,N_28982);
or U29143 (N_29143,N_28013,N_28375);
xnor U29144 (N_29144,N_28311,N_28809);
or U29145 (N_29145,N_28421,N_28415);
xor U29146 (N_29146,N_28706,N_28691);
and U29147 (N_29147,N_28426,N_28488);
nor U29148 (N_29148,N_28727,N_28321);
nand U29149 (N_29149,N_28898,N_28203);
or U29150 (N_29150,N_28921,N_28870);
xor U29151 (N_29151,N_28593,N_28207);
or U29152 (N_29152,N_28515,N_28233);
nor U29153 (N_29153,N_28899,N_28349);
xnor U29154 (N_29154,N_28561,N_28779);
xnor U29155 (N_29155,N_28388,N_28411);
and U29156 (N_29156,N_28429,N_28944);
nor U29157 (N_29157,N_28109,N_28247);
xor U29158 (N_29158,N_28093,N_28974);
nand U29159 (N_29159,N_28250,N_28158);
nand U29160 (N_29160,N_28695,N_28930);
and U29161 (N_29161,N_28590,N_28062);
nand U29162 (N_29162,N_28786,N_28320);
xnor U29163 (N_29163,N_28275,N_28937);
and U29164 (N_29164,N_28167,N_28995);
or U29165 (N_29165,N_28789,N_28795);
nand U29166 (N_29166,N_28036,N_28189);
nor U29167 (N_29167,N_28819,N_28696);
nor U29168 (N_29168,N_28526,N_28490);
nor U29169 (N_29169,N_28501,N_28616);
xnor U29170 (N_29170,N_28533,N_28534);
and U29171 (N_29171,N_28545,N_28265);
nand U29172 (N_29172,N_28012,N_28079);
xnor U29173 (N_29173,N_28419,N_28766);
xor U29174 (N_29174,N_28699,N_28008);
nor U29175 (N_29175,N_28748,N_28506);
xnor U29176 (N_29176,N_28931,N_28945);
or U29177 (N_29177,N_28669,N_28601);
nand U29178 (N_29178,N_28959,N_28894);
xor U29179 (N_29179,N_28314,N_28026);
and U29180 (N_29180,N_28187,N_28690);
or U29181 (N_29181,N_28300,N_28520);
xnor U29182 (N_29182,N_28939,N_28492);
nor U29183 (N_29183,N_28752,N_28837);
nor U29184 (N_29184,N_28735,N_28085);
and U29185 (N_29185,N_28647,N_28113);
nand U29186 (N_29186,N_28513,N_28200);
and U29187 (N_29187,N_28913,N_28880);
or U29188 (N_29188,N_28268,N_28551);
nand U29189 (N_29189,N_28051,N_28175);
and U29190 (N_29190,N_28466,N_28742);
nand U29191 (N_29191,N_28071,N_28436);
nand U29192 (N_29192,N_28966,N_28229);
nand U29193 (N_29193,N_28293,N_28605);
and U29194 (N_29194,N_28188,N_28890);
or U29195 (N_29195,N_28778,N_28807);
xnor U29196 (N_29196,N_28284,N_28633);
nand U29197 (N_29197,N_28283,N_28461);
nor U29198 (N_29198,N_28336,N_28650);
nand U29199 (N_29199,N_28266,N_28753);
or U29200 (N_29200,N_28845,N_28090);
xor U29201 (N_29201,N_28456,N_28397);
and U29202 (N_29202,N_28968,N_28875);
nor U29203 (N_29203,N_28969,N_28903);
or U29204 (N_29204,N_28149,N_28874);
nor U29205 (N_29205,N_28427,N_28935);
xor U29206 (N_29206,N_28654,N_28747);
xor U29207 (N_29207,N_28846,N_28594);
and U29208 (N_29208,N_28612,N_28686);
nand U29209 (N_29209,N_28528,N_28094);
or U29210 (N_29210,N_28319,N_28553);
or U29211 (N_29211,N_28843,N_28169);
and U29212 (N_29212,N_28486,N_28798);
and U29213 (N_29213,N_28463,N_28962);
xor U29214 (N_29214,N_28783,N_28922);
or U29215 (N_29215,N_28389,N_28885);
nor U29216 (N_29216,N_28714,N_28073);
and U29217 (N_29217,N_28993,N_28196);
xnor U29218 (N_29218,N_28276,N_28261);
xor U29219 (N_29219,N_28914,N_28987);
nor U29220 (N_29220,N_28003,N_28918);
xnor U29221 (N_29221,N_28136,N_28366);
nand U29222 (N_29222,N_28552,N_28412);
nor U29223 (N_29223,N_28755,N_28159);
and U29224 (N_29224,N_28082,N_28731);
xnor U29225 (N_29225,N_28573,N_28864);
and U29226 (N_29226,N_28131,N_28285);
nor U29227 (N_29227,N_28928,N_28122);
xnor U29228 (N_29228,N_28634,N_28462);
nor U29229 (N_29229,N_28384,N_28958);
and U29230 (N_29230,N_28662,N_28856);
xnor U29231 (N_29231,N_28950,N_28562);
xnor U29232 (N_29232,N_28286,N_28836);
xor U29233 (N_29233,N_28103,N_28635);
nand U29234 (N_29234,N_28482,N_28269);
and U29235 (N_29235,N_28784,N_28230);
nand U29236 (N_29236,N_28356,N_28847);
nor U29237 (N_29237,N_28315,N_28316);
nand U29238 (N_29238,N_28438,N_28312);
xnor U29239 (N_29239,N_28394,N_28050);
nor U29240 (N_29240,N_28404,N_28105);
nor U29241 (N_29241,N_28374,N_28019);
or U29242 (N_29242,N_28016,N_28991);
or U29243 (N_29243,N_28869,N_28416);
nor U29244 (N_29244,N_28006,N_28771);
and U29245 (N_29245,N_28754,N_28568);
xnor U29246 (N_29246,N_28910,N_28236);
xnor U29247 (N_29247,N_28262,N_28127);
or U29248 (N_29248,N_28091,N_28174);
xor U29249 (N_29249,N_28065,N_28761);
or U29250 (N_29250,N_28263,N_28808);
nand U29251 (N_29251,N_28396,N_28606);
or U29252 (N_29252,N_28478,N_28201);
nor U29253 (N_29253,N_28867,N_28014);
or U29254 (N_29254,N_28305,N_28547);
nor U29255 (N_29255,N_28785,N_28081);
nor U29256 (N_29256,N_28298,N_28834);
and U29257 (N_29257,N_28603,N_28332);
nand U29258 (N_29258,N_28720,N_28673);
xor U29259 (N_29259,N_28151,N_28100);
or U29260 (N_29260,N_28288,N_28405);
and U29261 (N_29261,N_28853,N_28525);
nor U29262 (N_29262,N_28543,N_28891);
and U29263 (N_29263,N_28838,N_28078);
nor U29264 (N_29264,N_28817,N_28565);
xor U29265 (N_29265,N_28424,N_28385);
nand U29266 (N_29266,N_28848,N_28835);
or U29267 (N_29267,N_28072,N_28804);
nor U29268 (N_29268,N_28181,N_28162);
nor U29269 (N_29269,N_28990,N_28829);
nor U29270 (N_29270,N_28661,N_28566);
and U29271 (N_29271,N_28002,N_28401);
and U29272 (N_29272,N_28398,N_28477);
or U29273 (N_29273,N_28810,N_28303);
nand U29274 (N_29274,N_28715,N_28728);
nor U29275 (N_29275,N_28862,N_28638);
xor U29276 (N_29276,N_28483,N_28943);
and U29277 (N_29277,N_28367,N_28095);
and U29278 (N_29278,N_28195,N_28138);
and U29279 (N_29279,N_28588,N_28096);
nand U29280 (N_29280,N_28256,N_28341);
nor U29281 (N_29281,N_28110,N_28820);
nor U29282 (N_29282,N_28823,N_28227);
nor U29283 (N_29283,N_28338,N_28409);
or U29284 (N_29284,N_28360,N_28111);
nor U29285 (N_29285,N_28290,N_28976);
nand U29286 (N_29286,N_28664,N_28307);
nand U29287 (N_29287,N_28005,N_28637);
xor U29288 (N_29288,N_28145,N_28119);
nor U29289 (N_29289,N_28802,N_28764);
xor U29290 (N_29290,N_28769,N_28165);
nand U29291 (N_29291,N_28032,N_28408);
nand U29292 (N_29292,N_28879,N_28147);
xnor U29293 (N_29293,N_28067,N_28216);
or U29294 (N_29294,N_28936,N_28292);
nor U29295 (N_29295,N_28986,N_28502);
nor U29296 (N_29296,N_28007,N_28212);
nor U29297 (N_29297,N_28684,N_28756);
nor U29298 (N_29298,N_28581,N_28460);
or U29299 (N_29299,N_28400,N_28815);
or U29300 (N_29300,N_28485,N_28744);
and U29301 (N_29301,N_28713,N_28909);
and U29302 (N_29302,N_28956,N_28179);
xor U29303 (N_29303,N_28270,N_28575);
xor U29304 (N_29304,N_28254,N_28194);
xnor U29305 (N_29305,N_28117,N_28563);
or U29306 (N_29306,N_28437,N_28359);
or U29307 (N_29307,N_28984,N_28104);
or U29308 (N_29308,N_28192,N_28556);
and U29309 (N_29309,N_28902,N_28975);
and U29310 (N_29310,N_28831,N_28832);
xor U29311 (N_29311,N_28164,N_28738);
or U29312 (N_29312,N_28530,N_28198);
nor U29313 (N_29313,N_28459,N_28954);
or U29314 (N_29314,N_28585,N_28723);
and U29315 (N_29315,N_28045,N_28645);
or U29316 (N_29316,N_28080,N_28604);
nand U29317 (N_29317,N_28430,N_28607);
nor U29318 (N_29318,N_28274,N_28679);
nor U29319 (N_29319,N_28066,N_28907);
or U29320 (N_29320,N_28793,N_28204);
nor U29321 (N_29321,N_28328,N_28061);
nand U29322 (N_29322,N_28523,N_28657);
and U29323 (N_29323,N_28342,N_28383);
nand U29324 (N_29324,N_28023,N_28295);
nand U29325 (N_29325,N_28860,N_28231);
xor U29326 (N_29326,N_28035,N_28060);
and U29327 (N_29327,N_28519,N_28770);
xor U29328 (N_29328,N_28549,N_28757);
nor U29329 (N_29329,N_28722,N_28364);
or U29330 (N_29330,N_28697,N_28345);
nand U29331 (N_29331,N_28365,N_28868);
and U29332 (N_29332,N_28544,N_28309);
or U29333 (N_29333,N_28591,N_28758);
and U29334 (N_29334,N_28054,N_28849);
or U29335 (N_29335,N_28693,N_28047);
nand U29336 (N_29336,N_28199,N_28346);
nand U29337 (N_29337,N_28542,N_28729);
or U29338 (N_29338,N_28137,N_28112);
xnor U29339 (N_29339,N_28734,N_28777);
nand U29340 (N_29340,N_28787,N_28306);
and U29341 (N_29341,N_28226,N_28191);
and U29342 (N_29342,N_28161,N_28028);
nand U29343 (N_29343,N_28118,N_28021);
nor U29344 (N_29344,N_28861,N_28750);
nor U29345 (N_29345,N_28420,N_28130);
and U29346 (N_29346,N_28866,N_28097);
or U29347 (N_29347,N_28009,N_28571);
or U29348 (N_29348,N_28223,N_28718);
and U29349 (N_29349,N_28623,N_28938);
nand U29350 (N_29350,N_28933,N_28851);
nor U29351 (N_29351,N_28782,N_28929);
nand U29352 (N_29352,N_28678,N_28597);
nand U29353 (N_29353,N_28089,N_28622);
or U29354 (N_29354,N_28494,N_28681);
nor U29355 (N_29355,N_28373,N_28660);
xor U29356 (N_29356,N_28325,N_28040);
or U29357 (N_29357,N_28517,N_28688);
xor U29358 (N_29358,N_28682,N_28653);
nand U29359 (N_29359,N_28355,N_28393);
and U29360 (N_29360,N_28872,N_28107);
or U29361 (N_29361,N_28142,N_28422);
and U29362 (N_29362,N_28431,N_28554);
nor U29363 (N_29363,N_28608,N_28058);
xor U29364 (N_29364,N_28915,N_28560);
nand U29365 (N_29365,N_28627,N_28799);
nand U29366 (N_29366,N_28680,N_28821);
or U29367 (N_29367,N_28805,N_28121);
and U29368 (N_29368,N_28582,N_28733);
nand U29369 (N_29369,N_28580,N_28310);
nor U29370 (N_29370,N_28780,N_28279);
xor U29371 (N_29371,N_28803,N_28790);
nor U29372 (N_29372,N_28160,N_28579);
nor U29373 (N_29373,N_28063,N_28961);
and U29374 (N_29374,N_28692,N_28511);
nand U29375 (N_29375,N_28380,N_28134);
and U29376 (N_29376,N_28354,N_28299);
xnor U29377 (N_29377,N_28334,N_28326);
nor U29378 (N_29378,N_28464,N_28614);
nor U29379 (N_29379,N_28249,N_28599);
or U29380 (N_29380,N_28906,N_28527);
or U29381 (N_29381,N_28241,N_28826);
nor U29382 (N_29382,N_28576,N_28450);
xnor U29383 (N_29383,N_28570,N_28296);
or U29384 (N_29384,N_28472,N_28505);
and U29385 (N_29385,N_28476,N_28806);
xnor U29386 (N_29386,N_28484,N_28135);
and U29387 (N_29387,N_28740,N_28369);
nand U29388 (N_29388,N_28683,N_28452);
nand U29389 (N_29389,N_28185,N_28140);
nor U29390 (N_29390,N_28955,N_28572);
nor U29391 (N_29391,N_28077,N_28946);
nor U29392 (N_29392,N_28636,N_28499);
nand U29393 (N_29393,N_28667,N_28170);
and U29394 (N_29394,N_28871,N_28414);
xnor U29395 (N_29395,N_28467,N_28282);
xor U29396 (N_29396,N_28646,N_28106);
nor U29397 (N_29397,N_28828,N_28387);
nand U29398 (N_29398,N_28540,N_28672);
or U29399 (N_29399,N_28577,N_28221);
nor U29400 (N_29400,N_28746,N_28157);
or U29401 (N_29401,N_28287,N_28640);
xor U29402 (N_29402,N_28475,N_28655);
nor U29403 (N_29403,N_28343,N_28382);
nor U29404 (N_29404,N_28468,N_28083);
or U29405 (N_29405,N_28796,N_28830);
or U29406 (N_29406,N_28656,N_28516);
nor U29407 (N_29407,N_28108,N_28011);
nor U29408 (N_29408,N_28042,N_28833);
xor U29409 (N_29409,N_28458,N_28048);
xnor U29410 (N_29410,N_28428,N_28034);
and U29411 (N_29411,N_28878,N_28495);
and U29412 (N_29412,N_28658,N_28324);
or U29413 (N_29413,N_28363,N_28532);
xor U29414 (N_29414,N_28923,N_28084);
xor U29415 (N_29415,N_28595,N_28244);
or U29416 (N_29416,N_28329,N_28448);
nand U29417 (N_29417,N_28126,N_28957);
nand U29418 (N_29418,N_28964,N_28001);
nand U29419 (N_29419,N_28465,N_28610);
or U29420 (N_29420,N_28557,N_28574);
nand U29421 (N_29421,N_28813,N_28512);
nand U29422 (N_29422,N_28253,N_28068);
and U29423 (N_29423,N_28473,N_28259);
nor U29424 (N_29424,N_28215,N_28522);
xnor U29425 (N_29425,N_28535,N_28087);
nand U29426 (N_29426,N_28278,N_28361);
nand U29427 (N_29427,N_28238,N_28139);
nor U29428 (N_29428,N_28659,N_28407);
or U29429 (N_29429,N_28925,N_28453);
or U29430 (N_29430,N_28017,N_28617);
nand U29431 (N_29431,N_28797,N_28257);
xor U29432 (N_29432,N_28854,N_28000);
xor U29433 (N_29433,N_28432,N_28154);
xor U29434 (N_29434,N_28234,N_28059);
nor U29435 (N_29435,N_28876,N_28703);
or U29436 (N_29436,N_28481,N_28781);
nor U29437 (N_29437,N_28272,N_28246);
and U29438 (N_29438,N_28824,N_28330);
nand U29439 (N_29439,N_28381,N_28507);
or U29440 (N_29440,N_28642,N_28559);
nand U29441 (N_29441,N_28235,N_28592);
or U29442 (N_29442,N_28447,N_28496);
or U29443 (N_29443,N_28765,N_28996);
and U29444 (N_29444,N_28651,N_28435);
or U29445 (N_29445,N_28998,N_28970);
nand U29446 (N_29446,N_28498,N_28487);
nand U29447 (N_29447,N_28816,N_28376);
or U29448 (N_29448,N_28339,N_28889);
nor U29449 (N_29449,N_28668,N_28074);
or U29450 (N_29450,N_28952,N_28855);
nor U29451 (N_29451,N_28371,N_28859);
xnor U29452 (N_29452,N_28064,N_28510);
and U29453 (N_29453,N_28043,N_28509);
and U29454 (N_29454,N_28099,N_28070);
nor U29455 (N_29455,N_28948,N_28977);
xor U29456 (N_29456,N_28704,N_28818);
or U29457 (N_29457,N_28711,N_28980);
nand U29458 (N_29458,N_28983,N_28027);
xor U29459 (N_29459,N_28038,N_28193);
or U29460 (N_29460,N_28716,N_28370);
nor U29461 (N_29461,N_28971,N_28069);
and U29462 (N_29462,N_28350,N_28056);
nand U29463 (N_29463,N_28445,N_28210);
nor U29464 (N_29464,N_28578,N_28670);
nor U29465 (N_29465,N_28347,N_28973);
nand U29466 (N_29466,N_28155,N_28168);
xor U29467 (N_29467,N_28791,N_28497);
nor U29468 (N_29468,N_28965,N_28677);
nor U29469 (N_29469,N_28273,N_28037);
nor U29470 (N_29470,N_28379,N_28596);
or U29471 (N_29471,N_28024,N_28908);
xor U29472 (N_29472,N_28289,N_28705);
or U29473 (N_29473,N_28184,N_28344);
nor U29474 (N_29474,N_28920,N_28550);
nand U29475 (N_29475,N_28434,N_28800);
or U29476 (N_29476,N_28632,N_28143);
and U29477 (N_29477,N_28333,N_28471);
nor U29478 (N_29478,N_28444,N_28877);
and U29479 (N_29479,N_28335,N_28205);
and U29480 (N_29480,N_28128,N_28997);
nor U29481 (N_29481,N_28124,N_28628);
nand U29482 (N_29482,N_28618,N_28763);
and U29483 (N_29483,N_28455,N_28418);
nand U29484 (N_29484,N_28888,N_28725);
or U29485 (N_29485,N_28222,N_28873);
nor U29486 (N_29486,N_28395,N_28322);
xor U29487 (N_29487,N_28675,N_28218);
xnor U29488 (N_29488,N_28449,N_28751);
nand U29489 (N_29489,N_28245,N_28602);
or U29490 (N_29490,N_28239,N_28989);
xnor U29491 (N_29491,N_28630,N_28896);
nand U29492 (N_29492,N_28884,N_28775);
nand U29493 (N_29493,N_28643,N_28737);
or U29494 (N_29494,N_28852,N_28277);
nor U29495 (N_29495,N_28242,N_28237);
nor U29496 (N_29496,N_28951,N_28773);
nand U29497 (N_29497,N_28057,N_28631);
xnor U29498 (N_29498,N_28267,N_28620);
nand U29499 (N_29499,N_28146,N_28721);
nand U29500 (N_29500,N_28459,N_28200);
and U29501 (N_29501,N_28399,N_28907);
and U29502 (N_29502,N_28877,N_28629);
nand U29503 (N_29503,N_28815,N_28655);
nand U29504 (N_29504,N_28586,N_28532);
nor U29505 (N_29505,N_28267,N_28748);
nand U29506 (N_29506,N_28606,N_28289);
or U29507 (N_29507,N_28856,N_28603);
and U29508 (N_29508,N_28666,N_28627);
nand U29509 (N_29509,N_28307,N_28939);
xor U29510 (N_29510,N_28688,N_28806);
nand U29511 (N_29511,N_28699,N_28028);
xnor U29512 (N_29512,N_28460,N_28461);
nor U29513 (N_29513,N_28904,N_28075);
xnor U29514 (N_29514,N_28815,N_28018);
nor U29515 (N_29515,N_28409,N_28841);
or U29516 (N_29516,N_28873,N_28838);
nand U29517 (N_29517,N_28561,N_28629);
and U29518 (N_29518,N_28390,N_28918);
and U29519 (N_29519,N_28386,N_28309);
nand U29520 (N_29520,N_28615,N_28545);
nor U29521 (N_29521,N_28427,N_28001);
nand U29522 (N_29522,N_28414,N_28954);
or U29523 (N_29523,N_28757,N_28284);
nand U29524 (N_29524,N_28108,N_28035);
nand U29525 (N_29525,N_28255,N_28783);
nand U29526 (N_29526,N_28533,N_28047);
nor U29527 (N_29527,N_28878,N_28389);
nand U29528 (N_29528,N_28321,N_28689);
or U29529 (N_29529,N_28121,N_28459);
and U29530 (N_29530,N_28676,N_28207);
xor U29531 (N_29531,N_28232,N_28413);
or U29532 (N_29532,N_28518,N_28232);
xor U29533 (N_29533,N_28770,N_28398);
or U29534 (N_29534,N_28950,N_28564);
nor U29535 (N_29535,N_28381,N_28622);
or U29536 (N_29536,N_28011,N_28374);
nand U29537 (N_29537,N_28815,N_28747);
xor U29538 (N_29538,N_28210,N_28836);
nand U29539 (N_29539,N_28146,N_28434);
nand U29540 (N_29540,N_28613,N_28840);
and U29541 (N_29541,N_28284,N_28678);
nor U29542 (N_29542,N_28085,N_28249);
xor U29543 (N_29543,N_28652,N_28676);
xor U29544 (N_29544,N_28956,N_28772);
and U29545 (N_29545,N_28412,N_28545);
nor U29546 (N_29546,N_28683,N_28518);
nor U29547 (N_29547,N_28503,N_28676);
nand U29548 (N_29548,N_28536,N_28994);
xnor U29549 (N_29549,N_28706,N_28770);
or U29550 (N_29550,N_28284,N_28735);
nand U29551 (N_29551,N_28086,N_28076);
nor U29552 (N_29552,N_28973,N_28568);
xor U29553 (N_29553,N_28533,N_28760);
nor U29554 (N_29554,N_28893,N_28110);
or U29555 (N_29555,N_28011,N_28547);
xnor U29556 (N_29556,N_28278,N_28975);
or U29557 (N_29557,N_28575,N_28456);
xnor U29558 (N_29558,N_28726,N_28853);
nor U29559 (N_29559,N_28154,N_28471);
and U29560 (N_29560,N_28889,N_28394);
nor U29561 (N_29561,N_28406,N_28885);
xnor U29562 (N_29562,N_28505,N_28817);
nand U29563 (N_29563,N_28894,N_28965);
nand U29564 (N_29564,N_28593,N_28318);
nand U29565 (N_29565,N_28456,N_28809);
nand U29566 (N_29566,N_28989,N_28935);
or U29567 (N_29567,N_28072,N_28904);
nor U29568 (N_29568,N_28514,N_28607);
or U29569 (N_29569,N_28653,N_28671);
and U29570 (N_29570,N_28081,N_28799);
nand U29571 (N_29571,N_28407,N_28923);
nor U29572 (N_29572,N_28401,N_28570);
or U29573 (N_29573,N_28956,N_28600);
or U29574 (N_29574,N_28535,N_28427);
and U29575 (N_29575,N_28406,N_28039);
nand U29576 (N_29576,N_28260,N_28920);
nor U29577 (N_29577,N_28340,N_28460);
nand U29578 (N_29578,N_28494,N_28332);
and U29579 (N_29579,N_28103,N_28986);
nor U29580 (N_29580,N_28988,N_28922);
nor U29581 (N_29581,N_28520,N_28644);
and U29582 (N_29582,N_28081,N_28930);
and U29583 (N_29583,N_28192,N_28157);
nor U29584 (N_29584,N_28096,N_28744);
xor U29585 (N_29585,N_28587,N_28697);
and U29586 (N_29586,N_28239,N_28789);
nor U29587 (N_29587,N_28611,N_28156);
or U29588 (N_29588,N_28641,N_28283);
nand U29589 (N_29589,N_28002,N_28183);
or U29590 (N_29590,N_28299,N_28944);
nor U29591 (N_29591,N_28768,N_28335);
nand U29592 (N_29592,N_28876,N_28524);
or U29593 (N_29593,N_28506,N_28272);
xor U29594 (N_29594,N_28794,N_28243);
xnor U29595 (N_29595,N_28319,N_28692);
xor U29596 (N_29596,N_28951,N_28157);
nand U29597 (N_29597,N_28023,N_28340);
nand U29598 (N_29598,N_28150,N_28409);
or U29599 (N_29599,N_28123,N_28097);
or U29600 (N_29600,N_28636,N_28187);
xnor U29601 (N_29601,N_28099,N_28530);
or U29602 (N_29602,N_28079,N_28554);
and U29603 (N_29603,N_28247,N_28460);
and U29604 (N_29604,N_28229,N_28849);
and U29605 (N_29605,N_28246,N_28539);
nand U29606 (N_29606,N_28069,N_28890);
nand U29607 (N_29607,N_28116,N_28582);
nor U29608 (N_29608,N_28891,N_28695);
and U29609 (N_29609,N_28483,N_28870);
xor U29610 (N_29610,N_28142,N_28969);
nand U29611 (N_29611,N_28502,N_28878);
xor U29612 (N_29612,N_28973,N_28133);
and U29613 (N_29613,N_28517,N_28386);
nand U29614 (N_29614,N_28559,N_28977);
or U29615 (N_29615,N_28703,N_28925);
or U29616 (N_29616,N_28937,N_28599);
nand U29617 (N_29617,N_28213,N_28708);
nand U29618 (N_29618,N_28950,N_28373);
or U29619 (N_29619,N_28044,N_28383);
xnor U29620 (N_29620,N_28802,N_28877);
nor U29621 (N_29621,N_28180,N_28932);
or U29622 (N_29622,N_28642,N_28639);
xnor U29623 (N_29623,N_28273,N_28147);
or U29624 (N_29624,N_28778,N_28646);
nor U29625 (N_29625,N_28090,N_28665);
and U29626 (N_29626,N_28202,N_28097);
nor U29627 (N_29627,N_28226,N_28877);
nand U29628 (N_29628,N_28757,N_28099);
or U29629 (N_29629,N_28885,N_28306);
and U29630 (N_29630,N_28771,N_28895);
and U29631 (N_29631,N_28561,N_28042);
and U29632 (N_29632,N_28750,N_28560);
nor U29633 (N_29633,N_28981,N_28856);
nand U29634 (N_29634,N_28255,N_28011);
nand U29635 (N_29635,N_28728,N_28664);
nor U29636 (N_29636,N_28829,N_28735);
nand U29637 (N_29637,N_28802,N_28282);
nor U29638 (N_29638,N_28837,N_28125);
or U29639 (N_29639,N_28366,N_28958);
and U29640 (N_29640,N_28444,N_28246);
nor U29641 (N_29641,N_28831,N_28708);
xor U29642 (N_29642,N_28688,N_28057);
nor U29643 (N_29643,N_28906,N_28318);
xnor U29644 (N_29644,N_28952,N_28923);
and U29645 (N_29645,N_28570,N_28599);
or U29646 (N_29646,N_28150,N_28137);
nand U29647 (N_29647,N_28302,N_28551);
nand U29648 (N_29648,N_28258,N_28620);
nor U29649 (N_29649,N_28394,N_28166);
nor U29650 (N_29650,N_28439,N_28210);
nor U29651 (N_29651,N_28444,N_28532);
or U29652 (N_29652,N_28608,N_28475);
nand U29653 (N_29653,N_28320,N_28579);
nand U29654 (N_29654,N_28459,N_28654);
and U29655 (N_29655,N_28322,N_28971);
xor U29656 (N_29656,N_28681,N_28818);
nor U29657 (N_29657,N_28836,N_28797);
and U29658 (N_29658,N_28703,N_28961);
nor U29659 (N_29659,N_28635,N_28143);
xnor U29660 (N_29660,N_28626,N_28117);
xnor U29661 (N_29661,N_28644,N_28623);
xnor U29662 (N_29662,N_28519,N_28969);
nand U29663 (N_29663,N_28445,N_28171);
or U29664 (N_29664,N_28483,N_28635);
and U29665 (N_29665,N_28627,N_28049);
xnor U29666 (N_29666,N_28262,N_28418);
nor U29667 (N_29667,N_28293,N_28659);
nand U29668 (N_29668,N_28773,N_28517);
xnor U29669 (N_29669,N_28491,N_28974);
nor U29670 (N_29670,N_28163,N_28086);
xnor U29671 (N_29671,N_28129,N_28840);
nor U29672 (N_29672,N_28286,N_28079);
or U29673 (N_29673,N_28463,N_28488);
and U29674 (N_29674,N_28284,N_28596);
or U29675 (N_29675,N_28673,N_28366);
or U29676 (N_29676,N_28741,N_28066);
and U29677 (N_29677,N_28984,N_28066);
nand U29678 (N_29678,N_28625,N_28982);
nand U29679 (N_29679,N_28081,N_28551);
nand U29680 (N_29680,N_28820,N_28987);
or U29681 (N_29681,N_28686,N_28770);
nand U29682 (N_29682,N_28208,N_28530);
or U29683 (N_29683,N_28888,N_28290);
and U29684 (N_29684,N_28377,N_28076);
nand U29685 (N_29685,N_28518,N_28925);
or U29686 (N_29686,N_28086,N_28715);
or U29687 (N_29687,N_28554,N_28255);
or U29688 (N_29688,N_28225,N_28749);
nand U29689 (N_29689,N_28179,N_28732);
nand U29690 (N_29690,N_28505,N_28877);
xor U29691 (N_29691,N_28917,N_28707);
nor U29692 (N_29692,N_28281,N_28328);
and U29693 (N_29693,N_28850,N_28865);
nor U29694 (N_29694,N_28548,N_28915);
nand U29695 (N_29695,N_28560,N_28783);
nand U29696 (N_29696,N_28322,N_28481);
xnor U29697 (N_29697,N_28304,N_28188);
xnor U29698 (N_29698,N_28040,N_28290);
and U29699 (N_29699,N_28885,N_28382);
or U29700 (N_29700,N_28755,N_28414);
xnor U29701 (N_29701,N_28012,N_28607);
or U29702 (N_29702,N_28435,N_28403);
and U29703 (N_29703,N_28412,N_28299);
xor U29704 (N_29704,N_28210,N_28986);
nand U29705 (N_29705,N_28111,N_28839);
nand U29706 (N_29706,N_28134,N_28125);
or U29707 (N_29707,N_28875,N_28189);
nor U29708 (N_29708,N_28722,N_28363);
and U29709 (N_29709,N_28292,N_28832);
or U29710 (N_29710,N_28821,N_28428);
nor U29711 (N_29711,N_28650,N_28691);
nor U29712 (N_29712,N_28981,N_28937);
xnor U29713 (N_29713,N_28691,N_28719);
or U29714 (N_29714,N_28651,N_28184);
or U29715 (N_29715,N_28298,N_28645);
xor U29716 (N_29716,N_28030,N_28649);
nand U29717 (N_29717,N_28735,N_28513);
nor U29718 (N_29718,N_28415,N_28984);
nand U29719 (N_29719,N_28662,N_28104);
nand U29720 (N_29720,N_28249,N_28264);
and U29721 (N_29721,N_28022,N_28564);
nand U29722 (N_29722,N_28106,N_28617);
nor U29723 (N_29723,N_28022,N_28160);
and U29724 (N_29724,N_28451,N_28322);
nand U29725 (N_29725,N_28617,N_28820);
xnor U29726 (N_29726,N_28019,N_28045);
nand U29727 (N_29727,N_28190,N_28861);
and U29728 (N_29728,N_28014,N_28241);
xor U29729 (N_29729,N_28503,N_28073);
and U29730 (N_29730,N_28333,N_28303);
nor U29731 (N_29731,N_28566,N_28587);
xnor U29732 (N_29732,N_28857,N_28549);
and U29733 (N_29733,N_28696,N_28503);
or U29734 (N_29734,N_28481,N_28157);
and U29735 (N_29735,N_28035,N_28410);
and U29736 (N_29736,N_28236,N_28594);
and U29737 (N_29737,N_28047,N_28310);
and U29738 (N_29738,N_28694,N_28400);
or U29739 (N_29739,N_28364,N_28348);
and U29740 (N_29740,N_28750,N_28486);
xor U29741 (N_29741,N_28559,N_28357);
xnor U29742 (N_29742,N_28681,N_28840);
or U29743 (N_29743,N_28531,N_28765);
nand U29744 (N_29744,N_28503,N_28596);
or U29745 (N_29745,N_28115,N_28624);
nand U29746 (N_29746,N_28802,N_28872);
nand U29747 (N_29747,N_28881,N_28212);
nand U29748 (N_29748,N_28835,N_28516);
and U29749 (N_29749,N_28261,N_28981);
or U29750 (N_29750,N_28277,N_28737);
and U29751 (N_29751,N_28880,N_28174);
and U29752 (N_29752,N_28482,N_28273);
nor U29753 (N_29753,N_28773,N_28652);
xnor U29754 (N_29754,N_28140,N_28738);
xor U29755 (N_29755,N_28347,N_28584);
nor U29756 (N_29756,N_28894,N_28858);
nor U29757 (N_29757,N_28856,N_28826);
and U29758 (N_29758,N_28876,N_28411);
nand U29759 (N_29759,N_28608,N_28749);
nor U29760 (N_29760,N_28753,N_28116);
xor U29761 (N_29761,N_28492,N_28335);
or U29762 (N_29762,N_28526,N_28815);
xor U29763 (N_29763,N_28593,N_28083);
and U29764 (N_29764,N_28210,N_28850);
and U29765 (N_29765,N_28643,N_28881);
or U29766 (N_29766,N_28125,N_28688);
nor U29767 (N_29767,N_28662,N_28146);
xor U29768 (N_29768,N_28105,N_28382);
or U29769 (N_29769,N_28892,N_28430);
nor U29770 (N_29770,N_28620,N_28098);
xor U29771 (N_29771,N_28012,N_28943);
and U29772 (N_29772,N_28479,N_28251);
xor U29773 (N_29773,N_28013,N_28746);
and U29774 (N_29774,N_28534,N_28201);
and U29775 (N_29775,N_28566,N_28534);
and U29776 (N_29776,N_28098,N_28246);
and U29777 (N_29777,N_28915,N_28964);
and U29778 (N_29778,N_28878,N_28934);
nand U29779 (N_29779,N_28658,N_28951);
xor U29780 (N_29780,N_28634,N_28846);
xnor U29781 (N_29781,N_28693,N_28147);
or U29782 (N_29782,N_28729,N_28956);
or U29783 (N_29783,N_28185,N_28176);
nand U29784 (N_29784,N_28416,N_28801);
xnor U29785 (N_29785,N_28037,N_28489);
nor U29786 (N_29786,N_28701,N_28210);
nor U29787 (N_29787,N_28693,N_28842);
and U29788 (N_29788,N_28780,N_28562);
or U29789 (N_29789,N_28987,N_28143);
nand U29790 (N_29790,N_28609,N_28683);
xor U29791 (N_29791,N_28847,N_28072);
nor U29792 (N_29792,N_28053,N_28309);
nor U29793 (N_29793,N_28757,N_28573);
or U29794 (N_29794,N_28919,N_28641);
nor U29795 (N_29795,N_28070,N_28372);
nand U29796 (N_29796,N_28200,N_28700);
nand U29797 (N_29797,N_28081,N_28076);
nor U29798 (N_29798,N_28970,N_28250);
xor U29799 (N_29799,N_28778,N_28613);
and U29800 (N_29800,N_28732,N_28888);
xor U29801 (N_29801,N_28399,N_28877);
or U29802 (N_29802,N_28442,N_28764);
or U29803 (N_29803,N_28437,N_28108);
and U29804 (N_29804,N_28822,N_28739);
xnor U29805 (N_29805,N_28246,N_28736);
or U29806 (N_29806,N_28441,N_28170);
and U29807 (N_29807,N_28076,N_28986);
nand U29808 (N_29808,N_28687,N_28926);
nor U29809 (N_29809,N_28519,N_28546);
xor U29810 (N_29810,N_28939,N_28361);
and U29811 (N_29811,N_28011,N_28046);
or U29812 (N_29812,N_28805,N_28511);
xnor U29813 (N_29813,N_28734,N_28752);
xnor U29814 (N_29814,N_28894,N_28321);
nor U29815 (N_29815,N_28329,N_28659);
xnor U29816 (N_29816,N_28661,N_28943);
or U29817 (N_29817,N_28622,N_28554);
or U29818 (N_29818,N_28684,N_28700);
or U29819 (N_29819,N_28959,N_28700);
xor U29820 (N_29820,N_28515,N_28933);
nor U29821 (N_29821,N_28219,N_28321);
and U29822 (N_29822,N_28653,N_28039);
or U29823 (N_29823,N_28882,N_28188);
and U29824 (N_29824,N_28082,N_28093);
nor U29825 (N_29825,N_28170,N_28541);
xnor U29826 (N_29826,N_28168,N_28553);
and U29827 (N_29827,N_28117,N_28694);
and U29828 (N_29828,N_28687,N_28429);
or U29829 (N_29829,N_28880,N_28350);
xnor U29830 (N_29830,N_28499,N_28327);
and U29831 (N_29831,N_28652,N_28167);
and U29832 (N_29832,N_28637,N_28281);
or U29833 (N_29833,N_28180,N_28863);
and U29834 (N_29834,N_28486,N_28188);
or U29835 (N_29835,N_28004,N_28240);
or U29836 (N_29836,N_28669,N_28103);
and U29837 (N_29837,N_28584,N_28744);
and U29838 (N_29838,N_28528,N_28271);
and U29839 (N_29839,N_28482,N_28822);
xnor U29840 (N_29840,N_28041,N_28031);
nor U29841 (N_29841,N_28515,N_28084);
and U29842 (N_29842,N_28704,N_28713);
nor U29843 (N_29843,N_28662,N_28530);
xnor U29844 (N_29844,N_28691,N_28540);
nor U29845 (N_29845,N_28608,N_28751);
nand U29846 (N_29846,N_28243,N_28765);
nor U29847 (N_29847,N_28873,N_28952);
xnor U29848 (N_29848,N_28599,N_28419);
nand U29849 (N_29849,N_28450,N_28338);
or U29850 (N_29850,N_28859,N_28312);
nand U29851 (N_29851,N_28760,N_28045);
nor U29852 (N_29852,N_28180,N_28143);
and U29853 (N_29853,N_28010,N_28473);
or U29854 (N_29854,N_28795,N_28799);
or U29855 (N_29855,N_28867,N_28097);
xor U29856 (N_29856,N_28210,N_28662);
nor U29857 (N_29857,N_28415,N_28307);
nor U29858 (N_29858,N_28076,N_28333);
and U29859 (N_29859,N_28425,N_28344);
and U29860 (N_29860,N_28138,N_28374);
and U29861 (N_29861,N_28162,N_28396);
and U29862 (N_29862,N_28784,N_28352);
or U29863 (N_29863,N_28141,N_28901);
or U29864 (N_29864,N_28857,N_28657);
nand U29865 (N_29865,N_28494,N_28789);
nand U29866 (N_29866,N_28954,N_28641);
and U29867 (N_29867,N_28451,N_28248);
xor U29868 (N_29868,N_28491,N_28099);
xor U29869 (N_29869,N_28406,N_28646);
nor U29870 (N_29870,N_28459,N_28714);
nor U29871 (N_29871,N_28473,N_28516);
nor U29872 (N_29872,N_28269,N_28492);
and U29873 (N_29873,N_28972,N_28563);
nor U29874 (N_29874,N_28210,N_28373);
nand U29875 (N_29875,N_28188,N_28347);
xor U29876 (N_29876,N_28169,N_28752);
nand U29877 (N_29877,N_28411,N_28124);
nand U29878 (N_29878,N_28722,N_28960);
nand U29879 (N_29879,N_28604,N_28172);
xnor U29880 (N_29880,N_28773,N_28990);
or U29881 (N_29881,N_28845,N_28543);
nor U29882 (N_29882,N_28112,N_28466);
nand U29883 (N_29883,N_28408,N_28560);
nand U29884 (N_29884,N_28777,N_28251);
nor U29885 (N_29885,N_28793,N_28431);
and U29886 (N_29886,N_28016,N_28973);
and U29887 (N_29887,N_28206,N_28285);
nor U29888 (N_29888,N_28170,N_28785);
and U29889 (N_29889,N_28680,N_28924);
nand U29890 (N_29890,N_28984,N_28037);
nand U29891 (N_29891,N_28473,N_28896);
xnor U29892 (N_29892,N_28480,N_28278);
or U29893 (N_29893,N_28704,N_28361);
nor U29894 (N_29894,N_28554,N_28025);
nand U29895 (N_29895,N_28750,N_28141);
nand U29896 (N_29896,N_28911,N_28369);
xor U29897 (N_29897,N_28908,N_28129);
and U29898 (N_29898,N_28517,N_28361);
or U29899 (N_29899,N_28634,N_28834);
nor U29900 (N_29900,N_28860,N_28266);
xnor U29901 (N_29901,N_28101,N_28361);
nand U29902 (N_29902,N_28060,N_28992);
xnor U29903 (N_29903,N_28972,N_28930);
and U29904 (N_29904,N_28224,N_28658);
or U29905 (N_29905,N_28837,N_28657);
and U29906 (N_29906,N_28067,N_28436);
xnor U29907 (N_29907,N_28687,N_28230);
nor U29908 (N_29908,N_28112,N_28542);
xnor U29909 (N_29909,N_28749,N_28135);
and U29910 (N_29910,N_28466,N_28700);
and U29911 (N_29911,N_28314,N_28123);
nor U29912 (N_29912,N_28671,N_28004);
nor U29913 (N_29913,N_28119,N_28825);
and U29914 (N_29914,N_28568,N_28197);
nand U29915 (N_29915,N_28101,N_28979);
nor U29916 (N_29916,N_28633,N_28365);
and U29917 (N_29917,N_28842,N_28276);
nor U29918 (N_29918,N_28002,N_28403);
nand U29919 (N_29919,N_28833,N_28776);
nand U29920 (N_29920,N_28565,N_28666);
nand U29921 (N_29921,N_28109,N_28851);
nand U29922 (N_29922,N_28037,N_28256);
and U29923 (N_29923,N_28235,N_28300);
nand U29924 (N_29924,N_28415,N_28658);
nor U29925 (N_29925,N_28858,N_28856);
and U29926 (N_29926,N_28087,N_28328);
nor U29927 (N_29927,N_28337,N_28587);
nor U29928 (N_29928,N_28357,N_28927);
and U29929 (N_29929,N_28503,N_28938);
and U29930 (N_29930,N_28168,N_28918);
or U29931 (N_29931,N_28612,N_28808);
nor U29932 (N_29932,N_28862,N_28912);
xor U29933 (N_29933,N_28196,N_28931);
nor U29934 (N_29934,N_28929,N_28920);
nor U29935 (N_29935,N_28116,N_28474);
nand U29936 (N_29936,N_28571,N_28962);
xor U29937 (N_29937,N_28987,N_28190);
nor U29938 (N_29938,N_28926,N_28870);
xnor U29939 (N_29939,N_28799,N_28450);
nor U29940 (N_29940,N_28481,N_28873);
and U29941 (N_29941,N_28677,N_28382);
nand U29942 (N_29942,N_28866,N_28548);
and U29943 (N_29943,N_28907,N_28926);
or U29944 (N_29944,N_28132,N_28627);
xor U29945 (N_29945,N_28268,N_28120);
nand U29946 (N_29946,N_28138,N_28515);
xor U29947 (N_29947,N_28991,N_28114);
or U29948 (N_29948,N_28269,N_28951);
and U29949 (N_29949,N_28474,N_28689);
and U29950 (N_29950,N_28027,N_28647);
xor U29951 (N_29951,N_28986,N_28471);
or U29952 (N_29952,N_28705,N_28192);
xnor U29953 (N_29953,N_28194,N_28206);
nor U29954 (N_29954,N_28462,N_28793);
nor U29955 (N_29955,N_28900,N_28276);
xnor U29956 (N_29956,N_28983,N_28505);
nor U29957 (N_29957,N_28859,N_28081);
nand U29958 (N_29958,N_28950,N_28706);
nand U29959 (N_29959,N_28929,N_28719);
or U29960 (N_29960,N_28413,N_28751);
nand U29961 (N_29961,N_28323,N_28548);
and U29962 (N_29962,N_28187,N_28547);
and U29963 (N_29963,N_28400,N_28341);
or U29964 (N_29964,N_28630,N_28341);
xnor U29965 (N_29965,N_28751,N_28333);
nand U29966 (N_29966,N_28055,N_28750);
or U29967 (N_29967,N_28879,N_28217);
or U29968 (N_29968,N_28756,N_28690);
and U29969 (N_29969,N_28581,N_28570);
xor U29970 (N_29970,N_28871,N_28178);
or U29971 (N_29971,N_28151,N_28411);
nor U29972 (N_29972,N_28044,N_28741);
or U29973 (N_29973,N_28410,N_28202);
nor U29974 (N_29974,N_28480,N_28405);
and U29975 (N_29975,N_28169,N_28040);
nor U29976 (N_29976,N_28596,N_28919);
xor U29977 (N_29977,N_28209,N_28851);
and U29978 (N_29978,N_28907,N_28631);
or U29979 (N_29979,N_28267,N_28245);
and U29980 (N_29980,N_28390,N_28417);
and U29981 (N_29981,N_28872,N_28597);
nand U29982 (N_29982,N_28361,N_28926);
and U29983 (N_29983,N_28230,N_28535);
nand U29984 (N_29984,N_28950,N_28234);
or U29985 (N_29985,N_28544,N_28660);
or U29986 (N_29986,N_28463,N_28007);
nand U29987 (N_29987,N_28049,N_28610);
nor U29988 (N_29988,N_28214,N_28278);
or U29989 (N_29989,N_28925,N_28110);
or U29990 (N_29990,N_28856,N_28257);
nor U29991 (N_29991,N_28239,N_28682);
nor U29992 (N_29992,N_28342,N_28984);
or U29993 (N_29993,N_28059,N_28244);
nand U29994 (N_29994,N_28658,N_28675);
nor U29995 (N_29995,N_28436,N_28299);
and U29996 (N_29996,N_28185,N_28225);
nor U29997 (N_29997,N_28371,N_28306);
xnor U29998 (N_29998,N_28652,N_28647);
nand U29999 (N_29999,N_28765,N_28824);
nand U30000 (N_30000,N_29241,N_29206);
and U30001 (N_30001,N_29013,N_29530);
nand U30002 (N_30002,N_29141,N_29247);
or U30003 (N_30003,N_29531,N_29103);
nand U30004 (N_30004,N_29096,N_29200);
or U30005 (N_30005,N_29543,N_29738);
nor U30006 (N_30006,N_29763,N_29237);
and U30007 (N_30007,N_29725,N_29457);
nand U30008 (N_30008,N_29193,N_29204);
or U30009 (N_30009,N_29355,N_29707);
and U30010 (N_30010,N_29442,N_29106);
nand U30011 (N_30011,N_29694,N_29087);
and U30012 (N_30012,N_29742,N_29577);
and U30013 (N_30013,N_29722,N_29056);
xnor U30014 (N_30014,N_29240,N_29340);
xor U30015 (N_30015,N_29380,N_29149);
nand U30016 (N_30016,N_29085,N_29454);
and U30017 (N_30017,N_29469,N_29119);
nor U30018 (N_30018,N_29127,N_29867);
and U30019 (N_30019,N_29709,N_29811);
xnor U30020 (N_30020,N_29350,N_29639);
or U30021 (N_30021,N_29347,N_29177);
nor U30022 (N_30022,N_29134,N_29851);
nand U30023 (N_30023,N_29348,N_29325);
nor U30024 (N_30024,N_29769,N_29649);
xnor U30025 (N_30025,N_29928,N_29853);
and U30026 (N_30026,N_29429,N_29434);
nor U30027 (N_30027,N_29456,N_29636);
or U30028 (N_30028,N_29791,N_29637);
nand U30029 (N_30029,N_29597,N_29421);
xor U30030 (N_30030,N_29076,N_29662);
and U30031 (N_30031,N_29635,N_29813);
nor U30032 (N_30032,N_29745,N_29046);
nand U30033 (N_30033,N_29940,N_29887);
or U30034 (N_30034,N_29941,N_29006);
or U30035 (N_30035,N_29894,N_29688);
nor U30036 (N_30036,N_29107,N_29658);
or U30037 (N_30037,N_29497,N_29943);
nand U30038 (N_30038,N_29494,N_29807);
or U30039 (N_30039,N_29751,N_29196);
and U30040 (N_30040,N_29010,N_29672);
xnor U30041 (N_30041,N_29837,N_29564);
and U30042 (N_30042,N_29418,N_29059);
nand U30043 (N_30043,N_29323,N_29183);
and U30044 (N_30044,N_29728,N_29021);
or U30045 (N_30045,N_29897,N_29307);
or U30046 (N_30046,N_29631,N_29857);
nand U30047 (N_30047,N_29248,N_29341);
xor U30048 (N_30048,N_29091,N_29938);
and U30049 (N_30049,N_29023,N_29303);
and U30050 (N_30050,N_29559,N_29830);
nand U30051 (N_30051,N_29081,N_29990);
or U30052 (N_30052,N_29616,N_29819);
or U30053 (N_30053,N_29093,N_29845);
nor U30054 (N_30054,N_29891,N_29731);
nor U30055 (N_30055,N_29078,N_29432);
nor U30056 (N_30056,N_29279,N_29917);
and U30057 (N_30057,N_29986,N_29681);
and U30058 (N_30058,N_29332,N_29411);
nand U30059 (N_30059,N_29836,N_29806);
xor U30060 (N_30060,N_29854,N_29218);
xnor U30061 (N_30061,N_29174,N_29372);
and U30062 (N_30062,N_29109,N_29272);
and U30063 (N_30063,N_29646,N_29624);
and U30064 (N_30064,N_29039,N_29070);
nor U30065 (N_30065,N_29228,N_29000);
nand U30066 (N_30066,N_29808,N_29339);
or U30067 (N_30067,N_29191,N_29143);
nor U30068 (N_30068,N_29100,N_29608);
nor U30069 (N_30069,N_29654,N_29294);
or U30070 (N_30070,N_29858,N_29433);
or U30071 (N_30071,N_29114,N_29569);
nand U30072 (N_30072,N_29644,N_29926);
and U30073 (N_30073,N_29120,N_29280);
or U30074 (N_30074,N_29168,N_29505);
nor U30075 (N_30075,N_29310,N_29855);
nor U30076 (N_30076,N_29071,N_29762);
nor U30077 (N_30077,N_29596,N_29118);
nor U30078 (N_30078,N_29668,N_29800);
xor U30079 (N_30079,N_29550,N_29718);
nand U30080 (N_30080,N_29112,N_29485);
xnor U30081 (N_30081,N_29150,N_29225);
nand U30082 (N_30082,N_29483,N_29966);
or U30083 (N_30083,N_29529,N_29036);
or U30084 (N_30084,N_29501,N_29002);
nand U30085 (N_30085,N_29638,N_29264);
nand U30086 (N_30086,N_29804,N_29828);
and U30087 (N_30087,N_29030,N_29714);
nor U30088 (N_30088,N_29152,N_29378);
and U30089 (N_30089,N_29416,N_29669);
nand U30090 (N_30090,N_29359,N_29026);
nand U30091 (N_30091,N_29090,N_29523);
nand U30092 (N_30092,N_29562,N_29282);
and U30093 (N_30093,N_29367,N_29615);
nor U30094 (N_30094,N_29047,N_29233);
nand U30095 (N_30095,N_29661,N_29319);
xnor U30096 (N_30096,N_29872,N_29301);
nand U30097 (N_30097,N_29826,N_29765);
and U30098 (N_30098,N_29060,N_29989);
and U30099 (N_30099,N_29630,N_29787);
nand U30100 (N_30100,N_29749,N_29117);
and U30101 (N_30101,N_29219,N_29384);
nor U30102 (N_30102,N_29679,N_29674);
nor U30103 (N_30103,N_29601,N_29017);
xor U30104 (N_30104,N_29506,N_29981);
and U30105 (N_30105,N_29146,N_29353);
nand U30106 (N_30106,N_29609,N_29436);
xnor U30107 (N_30107,N_29817,N_29685);
nor U30108 (N_30108,N_29831,N_29580);
nand U30109 (N_30109,N_29708,N_29877);
or U30110 (N_30110,N_29859,N_29029);
xnor U30111 (N_30111,N_29073,N_29563);
nor U30112 (N_30112,N_29629,N_29781);
or U30113 (N_30113,N_29466,N_29249);
nand U30114 (N_30114,N_29678,N_29898);
or U30115 (N_30115,N_29227,N_29185);
xor U30116 (N_30116,N_29420,N_29074);
nor U30117 (N_30117,N_29581,N_29713);
nand U30118 (N_30118,N_29759,N_29541);
nor U30119 (N_30119,N_29527,N_29014);
nand U30120 (N_30120,N_29982,N_29903);
xor U30121 (N_30121,N_29479,N_29996);
nand U30122 (N_30122,N_29600,N_29299);
and U30123 (N_30123,N_29594,N_29613);
nand U30124 (N_30124,N_29290,N_29703);
or U30125 (N_30125,N_29198,N_29784);
nor U30126 (N_30126,N_29995,N_29803);
xnor U30127 (N_30127,N_29832,N_29660);
or U30128 (N_30128,N_29097,N_29452);
nand U30129 (N_30129,N_29827,N_29387);
nand U30130 (N_30130,N_29306,N_29463);
nor U30131 (N_30131,N_29049,N_29670);
or U30132 (N_30132,N_29656,N_29399);
and U30133 (N_30133,N_29650,N_29153);
or U30134 (N_30134,N_29179,N_29331);
or U30135 (N_30135,N_29480,N_29991);
nor U30136 (N_30136,N_29330,N_29627);
and U30137 (N_30137,N_29126,N_29522);
nand U30138 (N_30138,N_29889,N_29213);
nand U30139 (N_30139,N_29809,N_29269);
and U30140 (N_30140,N_29088,N_29519);
xor U30141 (N_30141,N_29890,N_29673);
nand U30142 (N_30142,N_29602,N_29614);
and U30143 (N_30143,N_29189,N_29318);
xnor U30144 (N_30144,N_29232,N_29050);
xnor U30145 (N_30145,N_29545,N_29470);
or U30146 (N_30146,N_29296,N_29801);
or U30147 (N_30147,N_29390,N_29625);
and U30148 (N_30148,N_29733,N_29508);
and U30149 (N_30149,N_29175,N_29415);
nand U30150 (N_30150,N_29715,N_29717);
nand U30151 (N_30151,N_29513,N_29360);
nor U30152 (N_30152,N_29203,N_29863);
and U30153 (N_30153,N_29285,N_29211);
or U30154 (N_30154,N_29992,N_29773);
or U30155 (N_30155,N_29839,N_29210);
and U30156 (N_30156,N_29895,N_29907);
and U30157 (N_30157,N_29351,N_29385);
nor U30158 (N_30158,N_29133,N_29166);
or U30159 (N_30159,N_29215,N_29675);
nand U30160 (N_30160,N_29553,N_29920);
and U30161 (N_30161,N_29697,N_29910);
or U30162 (N_30162,N_29362,N_29901);
nand U30163 (N_30163,N_29746,N_29862);
or U30164 (N_30164,N_29441,N_29524);
xnor U30165 (N_30165,N_29861,N_29162);
xnor U30166 (N_30166,N_29040,N_29651);
nand U30167 (N_30167,N_29590,N_29473);
nand U30168 (N_30168,N_29972,N_29790);
nor U30169 (N_30169,N_29968,N_29948);
xnor U30170 (N_30170,N_29267,N_29573);
nand U30171 (N_30171,N_29955,N_29435);
or U30172 (N_30172,N_29375,N_29274);
xor U30173 (N_30173,N_29221,N_29987);
nor U30174 (N_30174,N_29652,N_29263);
or U30175 (N_30175,N_29304,N_29558);
nor U30176 (N_30176,N_29666,N_29018);
and U30177 (N_30177,N_29067,N_29974);
nand U30178 (N_30178,N_29879,N_29882);
and U30179 (N_30179,N_29487,N_29758);
and U30180 (N_30180,N_29947,N_29755);
nor U30181 (N_30181,N_29683,N_29251);
or U30182 (N_30182,N_29727,N_29423);
xor U30183 (N_30183,N_29843,N_29967);
and U30184 (N_30184,N_29785,N_29507);
or U30185 (N_30185,N_29234,N_29253);
nand U30186 (N_30186,N_29407,N_29102);
nand U30187 (N_30187,N_29345,N_29422);
xnor U30188 (N_30188,N_29346,N_29985);
nand U30189 (N_30189,N_29481,N_29289);
nand U30190 (N_30190,N_29640,N_29159);
nor U30191 (N_30191,N_29767,N_29892);
or U30192 (N_30192,N_29025,N_29293);
nor U30193 (N_30193,N_29880,N_29057);
nor U30194 (N_30194,N_29593,N_29752);
nand U30195 (N_30195,N_29537,N_29104);
nand U30196 (N_30196,N_29748,N_29268);
nor U30197 (N_30197,N_29605,N_29729);
or U30198 (N_30198,N_29389,N_29934);
nand U30199 (N_30199,N_29089,N_29142);
xor U30200 (N_30200,N_29584,N_29007);
or U30201 (N_30201,N_29896,N_29334);
xnor U30202 (N_30202,N_29549,N_29316);
nand U30203 (N_30203,N_29489,N_29846);
xnor U30204 (N_30204,N_29116,N_29302);
or U30205 (N_30205,N_29413,N_29988);
xnor U30206 (N_30206,N_29032,N_29144);
or U30207 (N_30207,N_29566,N_29428);
xor U30208 (N_30208,N_29711,N_29044);
nand U30209 (N_30209,N_29064,N_29287);
nor U30210 (N_30210,N_29795,N_29327);
or U30211 (N_30211,N_29724,N_29165);
nor U30212 (N_30212,N_29386,N_29546);
nor U30213 (N_30213,N_29570,N_29214);
or U30214 (N_30214,N_29271,N_29771);
nor U30215 (N_30215,N_29490,N_29315);
nand U30216 (N_30216,N_29802,N_29099);
nor U30217 (N_30217,N_29052,N_29736);
xnor U30218 (N_30218,N_29217,N_29368);
nor U30219 (N_30219,N_29599,N_29446);
and U30220 (N_30220,N_29667,N_29042);
nand U30221 (N_30221,N_29510,N_29455);
nor U30222 (N_30222,N_29919,N_29937);
nor U30223 (N_30223,N_29259,N_29061);
nor U30224 (N_30224,N_29122,N_29354);
nand U30225 (N_30225,N_29381,N_29925);
nor U30226 (N_30226,N_29438,N_29701);
xor U30227 (N_30227,N_29170,N_29111);
and U30228 (N_30228,N_29439,N_29680);
and U30229 (N_30229,N_29884,N_29893);
nor U30230 (N_30230,N_29027,N_29978);
nor U30231 (N_30231,N_29376,N_29911);
and U30232 (N_30232,N_29835,N_29178);
and U30233 (N_30233,N_29222,N_29398);
nand U30234 (N_30234,N_29011,N_29147);
nand U30235 (N_30235,N_29720,N_29689);
or U30236 (N_30236,N_29041,N_29132);
xnor U30237 (N_30237,N_29923,N_29874);
and U30238 (N_30238,N_29001,N_29084);
xnor U30239 (N_30239,N_29883,N_29512);
xnor U30240 (N_30240,N_29798,N_29443);
nand U30241 (N_30241,N_29451,N_29462);
and U30242 (N_30242,N_29356,N_29419);
nor U30243 (N_30243,N_29676,N_29504);
nor U30244 (N_30244,N_29909,N_29246);
xor U30245 (N_30245,N_29944,N_29574);
xnor U30246 (N_30246,N_29514,N_29993);
or U30247 (N_30247,N_29012,N_29291);
and U30248 (N_30248,N_29365,N_29850);
and U30249 (N_30249,N_29431,N_29645);
xor U30250 (N_30250,N_29951,N_29735);
nor U30251 (N_30251,N_29699,N_29417);
and U30252 (N_30252,N_29467,N_29437);
xor U30253 (N_30253,N_29383,N_29870);
nand U30254 (N_30254,N_29493,N_29969);
nor U30255 (N_30255,N_29960,N_29677);
nand U30256 (N_30256,N_29912,N_29164);
or U30257 (N_30257,N_29959,N_29933);
xor U30258 (N_30258,N_29939,N_29607);
and U30259 (N_30259,N_29252,N_29539);
and U30260 (N_30260,N_29190,N_29337);
xnor U30261 (N_30261,N_29295,N_29403);
and U30262 (N_30262,N_29772,N_29961);
nand U30263 (N_30263,N_29066,N_29131);
or U30264 (N_30264,N_29886,N_29582);
or U30265 (N_30265,N_29068,N_29158);
or U30266 (N_30266,N_29156,N_29250);
nor U30267 (N_30267,N_29932,N_29592);
xnor U30268 (N_30268,N_29918,N_29517);
and U30269 (N_30269,N_29145,N_29598);
nand U30270 (N_30270,N_29611,N_29321);
xor U30271 (N_30271,N_29197,N_29623);
nor U30272 (N_30272,N_29548,N_29397);
and U30273 (N_30273,N_29230,N_29405);
xor U30274 (N_30274,N_29154,N_29700);
and U30275 (N_30275,N_29187,N_29072);
nor U30276 (N_30276,N_29976,N_29535);
xor U30277 (N_30277,N_29536,N_29364);
or U30278 (N_30278,N_29526,N_29245);
nor U30279 (N_30279,N_29994,N_29053);
nand U30280 (N_30280,N_29730,N_29571);
nand U30281 (N_30281,N_29764,N_29352);
and U30282 (N_30282,N_29556,N_29038);
nand U30283 (N_30283,N_29212,N_29136);
xnor U30284 (N_30284,N_29840,N_29184);
or U30285 (N_30285,N_29757,N_29015);
xnor U30286 (N_30286,N_29113,N_29157);
and U30287 (N_30287,N_29984,N_29873);
and U30288 (N_30288,N_29542,N_29461);
nor U30289 (N_30289,N_29964,N_29388);
and U30290 (N_30290,N_29004,N_29706);
nor U30291 (N_30291,N_29124,N_29612);
and U30292 (N_30292,N_29477,N_29780);
nor U30293 (N_30293,N_29821,N_29797);
xnor U30294 (N_30294,N_29016,N_29815);
and U30295 (N_30295,N_29603,N_29058);
and U30296 (N_30296,N_29336,N_29628);
or U30297 (N_30297,N_29833,N_29547);
or U30298 (N_30298,N_29472,N_29031);
or U30299 (N_30299,N_29243,N_29450);
or U30300 (N_30300,N_29176,N_29447);
nor U30301 (N_30301,N_29238,N_29488);
nor U30302 (N_30302,N_29400,N_29077);
nor U30303 (N_30303,N_29478,N_29254);
or U30304 (N_30304,N_29810,N_29999);
nand U30305 (N_30305,N_29482,N_29459);
nand U30306 (N_30306,N_29692,N_29888);
and U30307 (N_30307,N_29275,N_29043);
or U30308 (N_30308,N_29721,N_29820);
xor U30309 (N_30309,N_29180,N_29308);
nor U30310 (N_30310,N_29412,N_29292);
nand U30311 (N_30311,N_29648,N_29617);
or U30312 (N_30312,N_29474,N_29425);
and U30313 (N_30313,N_29902,N_29578);
nor U30314 (N_30314,N_29086,N_29444);
xor U30315 (N_30315,N_29151,N_29037);
nor U30316 (N_30316,N_29155,N_29363);
nand U30317 (N_30317,N_29684,N_29687);
and U30318 (N_30318,N_29869,N_29401);
nor U30319 (N_30319,N_29740,N_29783);
nor U30320 (N_30320,N_29782,N_29534);
or U30321 (N_30321,N_29975,N_29284);
nor U30322 (N_30322,N_29567,N_29286);
nor U30323 (N_30323,N_29621,N_29283);
or U30324 (N_30324,N_29796,N_29929);
or U30325 (N_30325,N_29194,N_29852);
nor U30326 (N_30326,N_29904,N_29406);
or U30327 (N_30327,N_29576,N_29949);
nor U30328 (N_30328,N_29110,N_29108);
nor U30329 (N_30329,N_29540,N_29051);
nor U30330 (N_30330,N_29135,N_29048);
nand U30331 (N_30331,N_29357,N_29220);
nand U30332 (N_30332,N_29300,N_29019);
or U30333 (N_30333,N_29201,N_29260);
nor U30334 (N_30334,N_29814,N_29956);
nand U30335 (N_30335,N_29818,N_29395);
and U30336 (N_30336,N_29983,N_29202);
nor U30337 (N_30337,N_29465,N_29468);
xor U30338 (N_30338,N_29970,N_29931);
nand U30339 (N_30339,N_29643,N_29445);
or U30340 (N_30340,N_29737,N_29619);
nand U30341 (N_30341,N_29426,N_29900);
xnor U30342 (N_30342,N_29003,N_29829);
nor U30343 (N_30343,N_29256,N_29080);
or U30344 (N_30344,N_29878,N_29544);
nor U30345 (N_30345,N_29063,N_29908);
xnor U30346 (N_30346,N_29020,N_29123);
nand U30347 (N_30347,N_29278,N_29172);
nand U30348 (N_30348,N_29865,N_29226);
nor U30349 (N_30349,N_29953,N_29954);
nor U30350 (N_30350,N_29361,N_29977);
or U30351 (N_30351,N_29079,N_29169);
and U30352 (N_30352,N_29794,N_29265);
nand U30353 (N_30353,N_29500,N_29326);
and U30354 (N_30354,N_29235,N_29864);
xor U30355 (N_30355,N_29297,N_29945);
nand U30356 (N_30356,N_29744,N_29822);
nor U30357 (N_30357,N_29034,N_29734);
xnor U30358 (N_30358,N_29320,N_29973);
nand U30359 (N_30359,N_29231,N_29690);
nand U30360 (N_30360,N_29776,N_29775);
nand U30361 (N_30361,N_29671,N_29834);
nor U30362 (N_30362,N_29653,N_29799);
xnor U30363 (N_30363,N_29393,N_29698);
xor U30364 (N_30364,N_29195,N_29528);
or U30365 (N_30365,N_29805,N_29324);
and U30366 (N_30366,N_29277,N_29216);
xor U30367 (N_30367,N_29761,N_29591);
nand U30368 (N_30368,N_29188,N_29333);
nor U30369 (N_30369,N_29595,N_29266);
xnor U30370 (N_30370,N_29704,N_29410);
or U30371 (N_30371,N_29496,N_29486);
nand U30372 (N_30372,N_29322,N_29062);
nor U30373 (N_30373,N_29695,N_29161);
or U30374 (N_30374,N_29009,N_29997);
and U30375 (N_30375,N_29464,N_29239);
nor U30376 (N_30376,N_29906,N_29101);
or U30377 (N_30377,N_29379,N_29665);
and U30378 (N_30378,N_29273,N_29786);
nor U30379 (N_30379,N_29816,N_29572);
nand U30380 (N_30380,N_29313,N_29881);
nand U30381 (N_30381,N_29575,N_29723);
and U30382 (N_30382,N_29921,N_29712);
nand U30383 (N_30383,N_29950,N_29957);
nand U30384 (N_30384,N_29634,N_29373);
xnor U30385 (N_30385,N_29663,N_29199);
and U30386 (N_30386,N_29223,N_29192);
or U30387 (N_30387,N_29588,N_29094);
and U30388 (N_30388,N_29682,N_29747);
and U30389 (N_30389,N_29024,N_29732);
nor U30390 (N_30390,N_29396,N_29208);
and U30391 (N_30391,N_29344,N_29792);
xor U30392 (N_30392,N_29942,N_29930);
xnor U30393 (N_30393,N_29209,N_29779);
and U30394 (N_30394,N_29622,N_29121);
or U30395 (N_30395,N_29716,N_29626);
nand U30396 (N_30396,N_29533,N_29655);
nor U30397 (N_30397,N_29309,N_29491);
nor U30398 (N_30398,N_29756,N_29860);
nand U30399 (N_30399,N_29404,N_29916);
xor U30400 (N_30400,N_29448,N_29008);
and U30401 (N_30401,N_29812,N_29965);
nor U30402 (N_30402,N_29255,N_29236);
xor U30403 (N_30403,N_29952,N_29370);
or U30404 (N_30404,N_29586,N_29579);
and U30405 (N_30405,N_29440,N_29998);
nand U30406 (N_30406,N_29092,N_29587);
xnor U30407 (N_30407,N_29604,N_29963);
or U30408 (N_30408,N_29750,N_29691);
nand U30409 (N_30409,N_29298,N_29139);
nor U30410 (N_30410,N_29657,N_29922);
xor U30411 (N_30411,N_29885,N_29585);
nand U30412 (N_30412,N_29664,N_29276);
or U30413 (N_30413,N_29028,N_29927);
or U30414 (N_30414,N_29620,N_29518);
and U30415 (N_30415,N_29719,N_29205);
nor U30416 (N_30416,N_29186,N_29207);
xor U30417 (N_30417,N_29659,N_29589);
nor U30418 (N_30418,N_29022,N_29128);
xnor U30419 (N_30419,N_29181,N_29686);
and U30420 (N_30420,N_29741,N_29696);
and U30421 (N_30421,N_29532,N_29824);
nor U30422 (N_30422,N_29160,N_29525);
xor U30423 (N_30423,N_29329,N_29743);
and U30424 (N_30424,N_29632,N_29754);
nand U30425 (N_30425,N_29130,N_29069);
nand U30426 (N_30426,N_29760,N_29229);
nand U30427 (N_30427,N_29382,N_29392);
nand U30428 (N_30428,N_29475,N_29856);
nand U30429 (N_30429,N_29045,N_29498);
nand U30430 (N_30430,N_29962,N_29391);
nand U30431 (N_30431,N_29560,N_29371);
xnor U30432 (N_30432,N_29035,N_29502);
xor U30433 (N_30433,N_29095,N_29914);
nand U30434 (N_30434,N_29270,N_29693);
or U30435 (N_30435,N_29115,N_29710);
nor U30436 (N_30436,N_29641,N_29182);
nand U30437 (N_30437,N_29328,N_29726);
and U30438 (N_30438,N_29129,N_29606);
nand U30439 (N_30439,N_29958,N_29516);
or U30440 (N_30440,N_29261,N_29557);
and U30441 (N_30441,N_29082,N_29847);
nor U30442 (N_30442,N_29366,N_29849);
xnor U30443 (N_30443,N_29935,N_29138);
nor U30444 (N_30444,N_29257,N_29148);
nand U30445 (N_30445,N_29905,N_29915);
xnor U30446 (N_30446,N_29377,N_29312);
xor U30447 (N_30447,N_29471,N_29633);
xor U30448 (N_30448,N_29841,N_29552);
nor U30449 (N_30449,N_29946,N_29642);
nand U30450 (N_30450,N_29460,N_29766);
or U30451 (N_30451,N_29848,N_29137);
and U30452 (N_30452,N_29647,N_29244);
nor U30453 (N_30453,N_29555,N_29789);
nand U30454 (N_30454,N_29503,N_29875);
nand U30455 (N_30455,N_29224,N_29342);
and U30456 (N_30456,N_29098,N_29777);
xnor U30457 (N_30457,N_29369,N_29866);
and U30458 (N_30458,N_29565,N_29054);
and U30459 (N_30459,N_29702,N_29338);
or U30460 (N_30460,N_29610,N_29305);
nor U30461 (N_30461,N_29476,N_29258);
nor U30462 (N_30462,N_29739,N_29033);
nand U30463 (N_30463,N_29825,N_29913);
nor U30464 (N_30464,N_29499,N_29453);
and U30465 (N_30465,N_29374,N_29458);
or U30466 (N_30466,N_29163,N_29055);
or U30467 (N_30467,N_29125,N_29561);
nand U30468 (N_30468,N_29408,N_29394);
nand U30469 (N_30469,N_29936,N_29083);
and U30470 (N_30470,N_29511,N_29430);
and U30471 (N_30471,N_29551,N_29924);
or U30472 (N_30472,N_29793,N_29075);
or U30473 (N_30473,N_29424,N_29971);
nor U30474 (N_30474,N_29844,N_29317);
and U30475 (N_30475,N_29774,N_29788);
nand U30476 (N_30476,N_29753,N_29242);
and U30477 (N_30477,N_29314,N_29838);
and U30478 (N_30478,N_29705,N_29065);
nor U30479 (N_30479,N_29876,N_29509);
and U30480 (N_30480,N_29538,N_29778);
nor U30481 (N_30481,N_29554,N_29358);
nor U30482 (N_30482,N_29770,N_29568);
nor U30483 (N_30483,N_29167,N_29495);
or U30484 (N_30484,N_29402,N_29515);
nand U30485 (N_30485,N_29311,N_29868);
nand U30486 (N_30486,N_29105,N_29171);
nor U30487 (N_30487,N_29414,N_29140);
nor U30488 (N_30488,N_29768,N_29281);
xor U30489 (N_30489,N_29871,N_29335);
or U30490 (N_30490,N_29980,N_29492);
nor U30491 (N_30491,N_29449,N_29005);
or U30492 (N_30492,N_29427,N_29262);
nor U30493 (N_30493,N_29173,N_29343);
nand U30494 (N_30494,N_29520,N_29618);
xor U30495 (N_30495,N_29409,N_29979);
and U30496 (N_30496,N_29842,N_29484);
and U30497 (N_30497,N_29899,N_29823);
or U30498 (N_30498,N_29583,N_29288);
and U30499 (N_30499,N_29521,N_29349);
or U30500 (N_30500,N_29671,N_29457);
or U30501 (N_30501,N_29244,N_29696);
xnor U30502 (N_30502,N_29547,N_29762);
xor U30503 (N_30503,N_29395,N_29552);
nand U30504 (N_30504,N_29410,N_29455);
nand U30505 (N_30505,N_29862,N_29132);
nand U30506 (N_30506,N_29940,N_29504);
and U30507 (N_30507,N_29535,N_29754);
nand U30508 (N_30508,N_29763,N_29220);
xor U30509 (N_30509,N_29162,N_29878);
nand U30510 (N_30510,N_29583,N_29775);
nor U30511 (N_30511,N_29524,N_29517);
xor U30512 (N_30512,N_29249,N_29912);
nand U30513 (N_30513,N_29342,N_29636);
xnor U30514 (N_30514,N_29858,N_29083);
xor U30515 (N_30515,N_29275,N_29521);
or U30516 (N_30516,N_29583,N_29069);
nor U30517 (N_30517,N_29706,N_29453);
xnor U30518 (N_30518,N_29212,N_29039);
nor U30519 (N_30519,N_29108,N_29850);
and U30520 (N_30520,N_29092,N_29229);
or U30521 (N_30521,N_29841,N_29256);
xor U30522 (N_30522,N_29222,N_29396);
xnor U30523 (N_30523,N_29880,N_29960);
xor U30524 (N_30524,N_29295,N_29028);
or U30525 (N_30525,N_29387,N_29113);
xor U30526 (N_30526,N_29472,N_29827);
nand U30527 (N_30527,N_29889,N_29866);
or U30528 (N_30528,N_29930,N_29221);
and U30529 (N_30529,N_29423,N_29442);
xor U30530 (N_30530,N_29733,N_29668);
xnor U30531 (N_30531,N_29970,N_29776);
xnor U30532 (N_30532,N_29024,N_29491);
or U30533 (N_30533,N_29837,N_29746);
nor U30534 (N_30534,N_29684,N_29373);
or U30535 (N_30535,N_29122,N_29027);
or U30536 (N_30536,N_29662,N_29044);
xor U30537 (N_30537,N_29868,N_29494);
xnor U30538 (N_30538,N_29089,N_29213);
nor U30539 (N_30539,N_29787,N_29746);
and U30540 (N_30540,N_29468,N_29119);
nand U30541 (N_30541,N_29997,N_29461);
xnor U30542 (N_30542,N_29338,N_29646);
nand U30543 (N_30543,N_29691,N_29818);
nor U30544 (N_30544,N_29349,N_29526);
nand U30545 (N_30545,N_29472,N_29324);
xor U30546 (N_30546,N_29107,N_29713);
xnor U30547 (N_30547,N_29162,N_29771);
or U30548 (N_30548,N_29743,N_29710);
nand U30549 (N_30549,N_29195,N_29597);
and U30550 (N_30550,N_29221,N_29809);
or U30551 (N_30551,N_29297,N_29484);
or U30552 (N_30552,N_29402,N_29526);
or U30553 (N_30553,N_29394,N_29216);
and U30554 (N_30554,N_29620,N_29733);
or U30555 (N_30555,N_29340,N_29972);
nand U30556 (N_30556,N_29227,N_29144);
xnor U30557 (N_30557,N_29698,N_29154);
nor U30558 (N_30558,N_29187,N_29890);
nor U30559 (N_30559,N_29994,N_29507);
or U30560 (N_30560,N_29338,N_29433);
nand U30561 (N_30561,N_29731,N_29050);
nor U30562 (N_30562,N_29292,N_29946);
or U30563 (N_30563,N_29015,N_29388);
and U30564 (N_30564,N_29548,N_29611);
or U30565 (N_30565,N_29714,N_29703);
xnor U30566 (N_30566,N_29973,N_29558);
nor U30567 (N_30567,N_29298,N_29537);
and U30568 (N_30568,N_29513,N_29415);
nor U30569 (N_30569,N_29976,N_29593);
or U30570 (N_30570,N_29317,N_29754);
nor U30571 (N_30571,N_29548,N_29990);
and U30572 (N_30572,N_29961,N_29726);
xnor U30573 (N_30573,N_29094,N_29036);
or U30574 (N_30574,N_29028,N_29229);
xnor U30575 (N_30575,N_29201,N_29310);
nand U30576 (N_30576,N_29959,N_29096);
xnor U30577 (N_30577,N_29268,N_29056);
or U30578 (N_30578,N_29477,N_29998);
nor U30579 (N_30579,N_29416,N_29122);
or U30580 (N_30580,N_29022,N_29659);
and U30581 (N_30581,N_29218,N_29116);
nand U30582 (N_30582,N_29946,N_29199);
nor U30583 (N_30583,N_29571,N_29492);
nand U30584 (N_30584,N_29169,N_29018);
or U30585 (N_30585,N_29858,N_29575);
or U30586 (N_30586,N_29491,N_29023);
nor U30587 (N_30587,N_29931,N_29633);
xnor U30588 (N_30588,N_29005,N_29475);
xnor U30589 (N_30589,N_29805,N_29034);
nand U30590 (N_30590,N_29165,N_29266);
or U30591 (N_30591,N_29895,N_29358);
xnor U30592 (N_30592,N_29150,N_29715);
nand U30593 (N_30593,N_29789,N_29715);
or U30594 (N_30594,N_29351,N_29712);
and U30595 (N_30595,N_29295,N_29647);
or U30596 (N_30596,N_29028,N_29317);
xnor U30597 (N_30597,N_29977,N_29281);
nand U30598 (N_30598,N_29465,N_29311);
xnor U30599 (N_30599,N_29688,N_29204);
nor U30600 (N_30600,N_29157,N_29947);
xor U30601 (N_30601,N_29014,N_29681);
nor U30602 (N_30602,N_29160,N_29818);
xnor U30603 (N_30603,N_29905,N_29737);
nor U30604 (N_30604,N_29745,N_29482);
nor U30605 (N_30605,N_29718,N_29894);
and U30606 (N_30606,N_29352,N_29704);
and U30607 (N_30607,N_29038,N_29097);
xnor U30608 (N_30608,N_29543,N_29458);
nand U30609 (N_30609,N_29184,N_29999);
xnor U30610 (N_30610,N_29947,N_29121);
nor U30611 (N_30611,N_29744,N_29570);
nand U30612 (N_30612,N_29322,N_29439);
and U30613 (N_30613,N_29411,N_29343);
nand U30614 (N_30614,N_29772,N_29343);
nor U30615 (N_30615,N_29108,N_29361);
nand U30616 (N_30616,N_29135,N_29822);
nor U30617 (N_30617,N_29262,N_29927);
or U30618 (N_30618,N_29733,N_29934);
nand U30619 (N_30619,N_29165,N_29483);
and U30620 (N_30620,N_29817,N_29896);
nor U30621 (N_30621,N_29999,N_29881);
nor U30622 (N_30622,N_29260,N_29880);
or U30623 (N_30623,N_29127,N_29853);
and U30624 (N_30624,N_29023,N_29490);
and U30625 (N_30625,N_29052,N_29808);
nand U30626 (N_30626,N_29826,N_29638);
nor U30627 (N_30627,N_29927,N_29217);
or U30628 (N_30628,N_29349,N_29731);
nor U30629 (N_30629,N_29485,N_29602);
nor U30630 (N_30630,N_29174,N_29675);
and U30631 (N_30631,N_29044,N_29581);
nand U30632 (N_30632,N_29905,N_29973);
and U30633 (N_30633,N_29820,N_29058);
or U30634 (N_30634,N_29487,N_29296);
xor U30635 (N_30635,N_29939,N_29444);
and U30636 (N_30636,N_29164,N_29443);
and U30637 (N_30637,N_29249,N_29443);
nand U30638 (N_30638,N_29242,N_29087);
nor U30639 (N_30639,N_29718,N_29082);
nor U30640 (N_30640,N_29970,N_29298);
or U30641 (N_30641,N_29492,N_29277);
xor U30642 (N_30642,N_29579,N_29289);
and U30643 (N_30643,N_29528,N_29031);
nand U30644 (N_30644,N_29980,N_29973);
or U30645 (N_30645,N_29028,N_29920);
xor U30646 (N_30646,N_29274,N_29484);
nor U30647 (N_30647,N_29257,N_29599);
or U30648 (N_30648,N_29725,N_29068);
nor U30649 (N_30649,N_29805,N_29982);
nor U30650 (N_30650,N_29274,N_29561);
xnor U30651 (N_30651,N_29798,N_29317);
nor U30652 (N_30652,N_29928,N_29898);
or U30653 (N_30653,N_29335,N_29263);
xnor U30654 (N_30654,N_29411,N_29226);
or U30655 (N_30655,N_29673,N_29141);
nor U30656 (N_30656,N_29316,N_29694);
and U30657 (N_30657,N_29881,N_29065);
nor U30658 (N_30658,N_29802,N_29223);
nand U30659 (N_30659,N_29351,N_29103);
nand U30660 (N_30660,N_29915,N_29682);
and U30661 (N_30661,N_29708,N_29919);
nor U30662 (N_30662,N_29449,N_29698);
xor U30663 (N_30663,N_29237,N_29080);
and U30664 (N_30664,N_29566,N_29243);
or U30665 (N_30665,N_29773,N_29395);
nand U30666 (N_30666,N_29211,N_29714);
or U30667 (N_30667,N_29529,N_29151);
nor U30668 (N_30668,N_29643,N_29350);
and U30669 (N_30669,N_29982,N_29441);
xor U30670 (N_30670,N_29229,N_29375);
and U30671 (N_30671,N_29987,N_29451);
xor U30672 (N_30672,N_29531,N_29204);
xor U30673 (N_30673,N_29001,N_29406);
or U30674 (N_30674,N_29714,N_29298);
or U30675 (N_30675,N_29783,N_29214);
nand U30676 (N_30676,N_29138,N_29595);
and U30677 (N_30677,N_29638,N_29694);
nor U30678 (N_30678,N_29819,N_29828);
or U30679 (N_30679,N_29788,N_29313);
xor U30680 (N_30680,N_29199,N_29219);
nor U30681 (N_30681,N_29489,N_29888);
nor U30682 (N_30682,N_29264,N_29415);
and U30683 (N_30683,N_29247,N_29828);
and U30684 (N_30684,N_29654,N_29960);
xnor U30685 (N_30685,N_29108,N_29932);
or U30686 (N_30686,N_29432,N_29108);
nor U30687 (N_30687,N_29381,N_29861);
nand U30688 (N_30688,N_29409,N_29903);
and U30689 (N_30689,N_29559,N_29770);
nor U30690 (N_30690,N_29097,N_29191);
nand U30691 (N_30691,N_29336,N_29833);
and U30692 (N_30692,N_29780,N_29486);
or U30693 (N_30693,N_29009,N_29646);
xor U30694 (N_30694,N_29811,N_29296);
xor U30695 (N_30695,N_29098,N_29571);
xnor U30696 (N_30696,N_29559,N_29623);
or U30697 (N_30697,N_29686,N_29488);
nor U30698 (N_30698,N_29773,N_29783);
nor U30699 (N_30699,N_29438,N_29317);
nor U30700 (N_30700,N_29893,N_29043);
xor U30701 (N_30701,N_29580,N_29464);
xnor U30702 (N_30702,N_29928,N_29098);
nor U30703 (N_30703,N_29302,N_29052);
nor U30704 (N_30704,N_29972,N_29229);
nand U30705 (N_30705,N_29323,N_29410);
or U30706 (N_30706,N_29970,N_29475);
nor U30707 (N_30707,N_29991,N_29236);
or U30708 (N_30708,N_29834,N_29625);
xnor U30709 (N_30709,N_29533,N_29774);
nor U30710 (N_30710,N_29691,N_29597);
nand U30711 (N_30711,N_29492,N_29466);
or U30712 (N_30712,N_29874,N_29035);
nand U30713 (N_30713,N_29377,N_29145);
and U30714 (N_30714,N_29697,N_29629);
or U30715 (N_30715,N_29173,N_29581);
nand U30716 (N_30716,N_29480,N_29855);
nor U30717 (N_30717,N_29899,N_29507);
xor U30718 (N_30718,N_29875,N_29223);
and U30719 (N_30719,N_29779,N_29542);
or U30720 (N_30720,N_29670,N_29089);
xnor U30721 (N_30721,N_29409,N_29729);
and U30722 (N_30722,N_29069,N_29245);
and U30723 (N_30723,N_29420,N_29429);
nor U30724 (N_30724,N_29189,N_29620);
and U30725 (N_30725,N_29017,N_29980);
or U30726 (N_30726,N_29106,N_29251);
or U30727 (N_30727,N_29588,N_29981);
xor U30728 (N_30728,N_29690,N_29792);
xnor U30729 (N_30729,N_29885,N_29322);
nand U30730 (N_30730,N_29265,N_29464);
or U30731 (N_30731,N_29953,N_29644);
xnor U30732 (N_30732,N_29455,N_29560);
xor U30733 (N_30733,N_29595,N_29055);
nor U30734 (N_30734,N_29100,N_29716);
xnor U30735 (N_30735,N_29348,N_29496);
or U30736 (N_30736,N_29489,N_29441);
nor U30737 (N_30737,N_29392,N_29126);
nand U30738 (N_30738,N_29284,N_29969);
and U30739 (N_30739,N_29787,N_29946);
nand U30740 (N_30740,N_29082,N_29110);
or U30741 (N_30741,N_29136,N_29551);
nand U30742 (N_30742,N_29002,N_29208);
nand U30743 (N_30743,N_29162,N_29538);
nor U30744 (N_30744,N_29093,N_29507);
nor U30745 (N_30745,N_29029,N_29521);
xnor U30746 (N_30746,N_29389,N_29822);
nor U30747 (N_30747,N_29239,N_29224);
nand U30748 (N_30748,N_29616,N_29506);
nor U30749 (N_30749,N_29369,N_29714);
nor U30750 (N_30750,N_29037,N_29859);
and U30751 (N_30751,N_29273,N_29296);
or U30752 (N_30752,N_29189,N_29478);
and U30753 (N_30753,N_29403,N_29189);
or U30754 (N_30754,N_29002,N_29930);
or U30755 (N_30755,N_29684,N_29668);
or U30756 (N_30756,N_29371,N_29607);
xnor U30757 (N_30757,N_29708,N_29852);
and U30758 (N_30758,N_29370,N_29268);
nor U30759 (N_30759,N_29582,N_29846);
nor U30760 (N_30760,N_29250,N_29399);
and U30761 (N_30761,N_29717,N_29490);
nand U30762 (N_30762,N_29310,N_29524);
and U30763 (N_30763,N_29631,N_29041);
nand U30764 (N_30764,N_29360,N_29860);
xor U30765 (N_30765,N_29926,N_29366);
nor U30766 (N_30766,N_29780,N_29082);
and U30767 (N_30767,N_29875,N_29906);
xnor U30768 (N_30768,N_29281,N_29615);
or U30769 (N_30769,N_29220,N_29998);
nand U30770 (N_30770,N_29925,N_29287);
nand U30771 (N_30771,N_29809,N_29451);
xor U30772 (N_30772,N_29184,N_29396);
and U30773 (N_30773,N_29883,N_29830);
nor U30774 (N_30774,N_29942,N_29357);
or U30775 (N_30775,N_29954,N_29515);
nand U30776 (N_30776,N_29438,N_29374);
or U30777 (N_30777,N_29069,N_29139);
nor U30778 (N_30778,N_29984,N_29426);
nand U30779 (N_30779,N_29409,N_29052);
and U30780 (N_30780,N_29765,N_29848);
and U30781 (N_30781,N_29818,N_29084);
and U30782 (N_30782,N_29784,N_29841);
xnor U30783 (N_30783,N_29297,N_29142);
nor U30784 (N_30784,N_29978,N_29544);
and U30785 (N_30785,N_29571,N_29943);
or U30786 (N_30786,N_29075,N_29422);
xor U30787 (N_30787,N_29785,N_29480);
or U30788 (N_30788,N_29108,N_29888);
xnor U30789 (N_30789,N_29023,N_29842);
or U30790 (N_30790,N_29307,N_29261);
nand U30791 (N_30791,N_29181,N_29890);
and U30792 (N_30792,N_29099,N_29507);
nand U30793 (N_30793,N_29433,N_29837);
nor U30794 (N_30794,N_29118,N_29527);
or U30795 (N_30795,N_29698,N_29696);
nand U30796 (N_30796,N_29035,N_29813);
or U30797 (N_30797,N_29064,N_29487);
nor U30798 (N_30798,N_29376,N_29339);
or U30799 (N_30799,N_29670,N_29825);
xnor U30800 (N_30800,N_29205,N_29609);
or U30801 (N_30801,N_29135,N_29973);
nand U30802 (N_30802,N_29509,N_29579);
xnor U30803 (N_30803,N_29652,N_29320);
or U30804 (N_30804,N_29190,N_29502);
xnor U30805 (N_30805,N_29291,N_29804);
nand U30806 (N_30806,N_29434,N_29787);
nor U30807 (N_30807,N_29435,N_29210);
or U30808 (N_30808,N_29523,N_29717);
and U30809 (N_30809,N_29154,N_29801);
xnor U30810 (N_30810,N_29331,N_29750);
xor U30811 (N_30811,N_29997,N_29673);
and U30812 (N_30812,N_29071,N_29307);
xnor U30813 (N_30813,N_29592,N_29286);
nor U30814 (N_30814,N_29707,N_29212);
and U30815 (N_30815,N_29028,N_29079);
xnor U30816 (N_30816,N_29351,N_29227);
nand U30817 (N_30817,N_29748,N_29556);
nor U30818 (N_30818,N_29889,N_29876);
xnor U30819 (N_30819,N_29495,N_29417);
nor U30820 (N_30820,N_29955,N_29378);
xnor U30821 (N_30821,N_29954,N_29006);
or U30822 (N_30822,N_29429,N_29135);
and U30823 (N_30823,N_29376,N_29787);
or U30824 (N_30824,N_29870,N_29118);
nand U30825 (N_30825,N_29823,N_29847);
or U30826 (N_30826,N_29008,N_29276);
xor U30827 (N_30827,N_29774,N_29623);
nor U30828 (N_30828,N_29836,N_29850);
nand U30829 (N_30829,N_29281,N_29690);
and U30830 (N_30830,N_29006,N_29503);
or U30831 (N_30831,N_29399,N_29361);
and U30832 (N_30832,N_29119,N_29514);
and U30833 (N_30833,N_29696,N_29187);
nor U30834 (N_30834,N_29704,N_29462);
nand U30835 (N_30835,N_29039,N_29169);
xor U30836 (N_30836,N_29669,N_29928);
and U30837 (N_30837,N_29941,N_29632);
xnor U30838 (N_30838,N_29380,N_29713);
nor U30839 (N_30839,N_29046,N_29214);
nand U30840 (N_30840,N_29490,N_29299);
xor U30841 (N_30841,N_29181,N_29616);
or U30842 (N_30842,N_29463,N_29747);
and U30843 (N_30843,N_29061,N_29358);
nand U30844 (N_30844,N_29677,N_29949);
xor U30845 (N_30845,N_29094,N_29722);
nand U30846 (N_30846,N_29156,N_29202);
or U30847 (N_30847,N_29725,N_29163);
xnor U30848 (N_30848,N_29911,N_29629);
nor U30849 (N_30849,N_29776,N_29766);
or U30850 (N_30850,N_29333,N_29125);
xnor U30851 (N_30851,N_29291,N_29915);
xor U30852 (N_30852,N_29343,N_29793);
nand U30853 (N_30853,N_29671,N_29123);
nand U30854 (N_30854,N_29070,N_29408);
or U30855 (N_30855,N_29678,N_29840);
or U30856 (N_30856,N_29543,N_29307);
xnor U30857 (N_30857,N_29413,N_29708);
nor U30858 (N_30858,N_29133,N_29013);
xor U30859 (N_30859,N_29592,N_29378);
or U30860 (N_30860,N_29395,N_29984);
nor U30861 (N_30861,N_29410,N_29909);
nand U30862 (N_30862,N_29886,N_29468);
nor U30863 (N_30863,N_29911,N_29990);
xor U30864 (N_30864,N_29643,N_29927);
nor U30865 (N_30865,N_29757,N_29498);
nand U30866 (N_30866,N_29853,N_29885);
nor U30867 (N_30867,N_29107,N_29811);
xor U30868 (N_30868,N_29706,N_29603);
nor U30869 (N_30869,N_29140,N_29241);
and U30870 (N_30870,N_29068,N_29364);
or U30871 (N_30871,N_29008,N_29247);
and U30872 (N_30872,N_29729,N_29799);
xor U30873 (N_30873,N_29803,N_29238);
nand U30874 (N_30874,N_29453,N_29502);
and U30875 (N_30875,N_29720,N_29977);
and U30876 (N_30876,N_29318,N_29873);
or U30877 (N_30877,N_29910,N_29181);
or U30878 (N_30878,N_29797,N_29822);
nor U30879 (N_30879,N_29080,N_29789);
xnor U30880 (N_30880,N_29690,N_29704);
or U30881 (N_30881,N_29447,N_29218);
nor U30882 (N_30882,N_29070,N_29587);
or U30883 (N_30883,N_29677,N_29137);
nor U30884 (N_30884,N_29757,N_29094);
xnor U30885 (N_30885,N_29936,N_29124);
and U30886 (N_30886,N_29193,N_29871);
and U30887 (N_30887,N_29283,N_29961);
nand U30888 (N_30888,N_29343,N_29155);
nor U30889 (N_30889,N_29189,N_29070);
and U30890 (N_30890,N_29575,N_29509);
or U30891 (N_30891,N_29885,N_29699);
and U30892 (N_30892,N_29228,N_29558);
nand U30893 (N_30893,N_29453,N_29567);
and U30894 (N_30894,N_29071,N_29888);
or U30895 (N_30895,N_29254,N_29613);
and U30896 (N_30896,N_29108,N_29546);
and U30897 (N_30897,N_29668,N_29538);
or U30898 (N_30898,N_29487,N_29718);
and U30899 (N_30899,N_29093,N_29363);
and U30900 (N_30900,N_29022,N_29821);
and U30901 (N_30901,N_29003,N_29865);
nor U30902 (N_30902,N_29910,N_29160);
and U30903 (N_30903,N_29526,N_29864);
and U30904 (N_30904,N_29083,N_29843);
nand U30905 (N_30905,N_29683,N_29049);
and U30906 (N_30906,N_29194,N_29100);
nand U30907 (N_30907,N_29533,N_29511);
and U30908 (N_30908,N_29790,N_29994);
xor U30909 (N_30909,N_29210,N_29034);
xnor U30910 (N_30910,N_29436,N_29171);
and U30911 (N_30911,N_29712,N_29212);
xor U30912 (N_30912,N_29576,N_29239);
or U30913 (N_30913,N_29592,N_29996);
nor U30914 (N_30914,N_29781,N_29750);
and U30915 (N_30915,N_29808,N_29608);
and U30916 (N_30916,N_29127,N_29845);
nor U30917 (N_30917,N_29948,N_29689);
nor U30918 (N_30918,N_29864,N_29629);
and U30919 (N_30919,N_29866,N_29661);
nand U30920 (N_30920,N_29588,N_29644);
nor U30921 (N_30921,N_29429,N_29382);
nor U30922 (N_30922,N_29053,N_29292);
xor U30923 (N_30923,N_29782,N_29744);
or U30924 (N_30924,N_29400,N_29861);
nor U30925 (N_30925,N_29017,N_29034);
nand U30926 (N_30926,N_29012,N_29366);
nand U30927 (N_30927,N_29545,N_29281);
xor U30928 (N_30928,N_29707,N_29266);
nor U30929 (N_30929,N_29164,N_29829);
nor U30930 (N_30930,N_29136,N_29926);
nand U30931 (N_30931,N_29138,N_29894);
nand U30932 (N_30932,N_29067,N_29533);
and U30933 (N_30933,N_29356,N_29012);
or U30934 (N_30934,N_29836,N_29233);
nor U30935 (N_30935,N_29467,N_29582);
and U30936 (N_30936,N_29168,N_29179);
xor U30937 (N_30937,N_29388,N_29059);
and U30938 (N_30938,N_29575,N_29128);
xnor U30939 (N_30939,N_29031,N_29965);
or U30940 (N_30940,N_29311,N_29361);
nor U30941 (N_30941,N_29673,N_29775);
nand U30942 (N_30942,N_29751,N_29052);
nor U30943 (N_30943,N_29179,N_29624);
and U30944 (N_30944,N_29591,N_29965);
or U30945 (N_30945,N_29001,N_29915);
and U30946 (N_30946,N_29117,N_29890);
nand U30947 (N_30947,N_29757,N_29130);
nand U30948 (N_30948,N_29192,N_29527);
or U30949 (N_30949,N_29549,N_29002);
and U30950 (N_30950,N_29207,N_29233);
nor U30951 (N_30951,N_29413,N_29433);
nor U30952 (N_30952,N_29545,N_29456);
or U30953 (N_30953,N_29260,N_29904);
or U30954 (N_30954,N_29641,N_29200);
or U30955 (N_30955,N_29189,N_29701);
nor U30956 (N_30956,N_29468,N_29812);
nor U30957 (N_30957,N_29336,N_29485);
and U30958 (N_30958,N_29917,N_29376);
nor U30959 (N_30959,N_29510,N_29061);
xor U30960 (N_30960,N_29840,N_29800);
nand U30961 (N_30961,N_29209,N_29998);
nand U30962 (N_30962,N_29010,N_29559);
or U30963 (N_30963,N_29708,N_29672);
or U30964 (N_30964,N_29637,N_29312);
or U30965 (N_30965,N_29558,N_29015);
xnor U30966 (N_30966,N_29206,N_29521);
nand U30967 (N_30967,N_29351,N_29800);
xor U30968 (N_30968,N_29018,N_29237);
xor U30969 (N_30969,N_29757,N_29150);
xnor U30970 (N_30970,N_29479,N_29264);
nand U30971 (N_30971,N_29902,N_29153);
and U30972 (N_30972,N_29775,N_29727);
or U30973 (N_30973,N_29245,N_29990);
nand U30974 (N_30974,N_29320,N_29252);
xnor U30975 (N_30975,N_29312,N_29721);
nand U30976 (N_30976,N_29572,N_29198);
and U30977 (N_30977,N_29297,N_29140);
nor U30978 (N_30978,N_29150,N_29396);
nor U30979 (N_30979,N_29120,N_29851);
nor U30980 (N_30980,N_29923,N_29541);
nor U30981 (N_30981,N_29025,N_29947);
nand U30982 (N_30982,N_29197,N_29605);
or U30983 (N_30983,N_29085,N_29300);
nor U30984 (N_30984,N_29085,N_29251);
nand U30985 (N_30985,N_29752,N_29761);
xor U30986 (N_30986,N_29424,N_29005);
or U30987 (N_30987,N_29443,N_29251);
nand U30988 (N_30988,N_29710,N_29454);
or U30989 (N_30989,N_29637,N_29590);
and U30990 (N_30990,N_29376,N_29647);
or U30991 (N_30991,N_29940,N_29789);
or U30992 (N_30992,N_29237,N_29169);
or U30993 (N_30993,N_29026,N_29370);
nand U30994 (N_30994,N_29893,N_29254);
or U30995 (N_30995,N_29465,N_29494);
and U30996 (N_30996,N_29056,N_29102);
xor U30997 (N_30997,N_29911,N_29311);
xor U30998 (N_30998,N_29266,N_29191);
xor U30999 (N_30999,N_29001,N_29705);
and U31000 (N_31000,N_30373,N_30046);
or U31001 (N_31001,N_30695,N_30062);
xnor U31002 (N_31002,N_30385,N_30261);
xnor U31003 (N_31003,N_30510,N_30964);
xnor U31004 (N_31004,N_30977,N_30195);
nand U31005 (N_31005,N_30281,N_30835);
or U31006 (N_31006,N_30871,N_30819);
nor U31007 (N_31007,N_30740,N_30343);
xor U31008 (N_31008,N_30122,N_30151);
nor U31009 (N_31009,N_30205,N_30033);
nor U31010 (N_31010,N_30217,N_30738);
nor U31011 (N_31011,N_30859,N_30282);
or U31012 (N_31012,N_30173,N_30066);
xor U31013 (N_31013,N_30279,N_30707);
nand U31014 (N_31014,N_30039,N_30488);
xnor U31015 (N_31015,N_30547,N_30833);
or U31016 (N_31016,N_30017,N_30928);
nand U31017 (N_31017,N_30537,N_30974);
and U31018 (N_31018,N_30721,N_30697);
nor U31019 (N_31019,N_30656,N_30240);
and U31020 (N_31020,N_30801,N_30274);
nand U31021 (N_31021,N_30834,N_30542);
and U31022 (N_31022,N_30919,N_30684);
nor U31023 (N_31023,N_30898,N_30090);
nor U31024 (N_31024,N_30321,N_30357);
nand U31025 (N_31025,N_30253,N_30007);
nand U31026 (N_31026,N_30647,N_30093);
and U31027 (N_31027,N_30899,N_30925);
or U31028 (N_31028,N_30138,N_30992);
and U31029 (N_31029,N_30862,N_30358);
xor U31030 (N_31030,N_30768,N_30519);
nor U31031 (N_31031,N_30569,N_30996);
xnor U31032 (N_31032,N_30784,N_30951);
nand U31033 (N_31033,N_30500,N_30592);
nor U31034 (N_31034,N_30089,N_30926);
xnor U31035 (N_31035,N_30502,N_30757);
or U31036 (N_31036,N_30437,N_30669);
or U31037 (N_31037,N_30418,N_30696);
or U31038 (N_31038,N_30599,N_30139);
nand U31039 (N_31039,N_30411,N_30248);
nor U31040 (N_31040,N_30233,N_30483);
nand U31041 (N_31041,N_30484,N_30178);
nand U31042 (N_31042,N_30566,N_30097);
or U31043 (N_31043,N_30280,N_30583);
nor U31044 (N_31044,N_30639,N_30296);
or U31045 (N_31045,N_30146,N_30242);
nand U31046 (N_31046,N_30962,N_30410);
nand U31047 (N_31047,N_30915,N_30297);
and U31048 (N_31048,N_30074,N_30155);
and U31049 (N_31049,N_30239,N_30931);
or U31050 (N_31050,N_30559,N_30092);
nand U31051 (N_31051,N_30235,N_30844);
nand U31052 (N_31052,N_30517,N_30783);
nand U31053 (N_31053,N_30210,N_30989);
or U31054 (N_31054,N_30060,N_30271);
nor U31055 (N_31055,N_30021,N_30107);
nor U31056 (N_31056,N_30312,N_30975);
nand U31057 (N_31057,N_30895,N_30886);
or U31058 (N_31058,N_30043,N_30446);
or U31059 (N_31059,N_30058,N_30885);
xor U31060 (N_31060,N_30169,N_30479);
and U31061 (N_31061,N_30106,N_30544);
nor U31062 (N_31062,N_30661,N_30606);
xor U31063 (N_31063,N_30643,N_30565);
xor U31064 (N_31064,N_30005,N_30352);
or U31065 (N_31065,N_30846,N_30777);
nor U31066 (N_31066,N_30476,N_30512);
xnor U31067 (N_31067,N_30737,N_30580);
nor U31068 (N_31068,N_30073,N_30831);
nand U31069 (N_31069,N_30393,N_30376);
or U31070 (N_31070,N_30191,N_30010);
and U31071 (N_31071,N_30515,N_30397);
or U31072 (N_31072,N_30957,N_30438);
xor U31073 (N_31073,N_30725,N_30382);
xnor U31074 (N_31074,N_30958,N_30826);
nor U31075 (N_31075,N_30897,N_30331);
nor U31076 (N_31076,N_30482,N_30621);
and U31077 (N_31077,N_30687,N_30563);
or U31078 (N_31078,N_30259,N_30460);
and U31079 (N_31079,N_30392,N_30270);
or U31080 (N_31080,N_30341,N_30099);
xnor U31081 (N_31081,N_30407,N_30377);
nand U31082 (N_31082,N_30558,N_30267);
xnor U31083 (N_31083,N_30396,N_30531);
nand U31084 (N_31084,N_30983,N_30703);
xnor U31085 (N_31085,N_30865,N_30199);
and U31086 (N_31086,N_30550,N_30944);
nand U31087 (N_31087,N_30568,N_30490);
and U31088 (N_31088,N_30809,N_30256);
and U31089 (N_31089,N_30234,N_30882);
or U31090 (N_31090,N_30820,N_30413);
and U31091 (N_31091,N_30444,N_30693);
or U31092 (N_31092,N_30328,N_30454);
and U31093 (N_31093,N_30469,N_30657);
nand U31094 (N_31094,N_30346,N_30405);
nor U31095 (N_31095,N_30749,N_30876);
xor U31096 (N_31096,N_30412,N_30244);
nor U31097 (N_31097,N_30228,N_30277);
xor U31098 (N_31098,N_30236,N_30634);
or U31099 (N_31099,N_30555,N_30604);
nor U31100 (N_31100,N_30430,N_30475);
or U31101 (N_31101,N_30748,N_30813);
and U31102 (N_31102,N_30466,N_30069);
or U31103 (N_31103,N_30193,N_30760);
and U31104 (N_31104,N_30736,N_30335);
or U31105 (N_31105,N_30627,N_30789);
xnor U31106 (N_31106,N_30215,N_30434);
nand U31107 (N_31107,N_30560,N_30160);
and U31108 (N_31108,N_30959,N_30858);
xor U31109 (N_31109,N_30116,N_30063);
nor U31110 (N_31110,N_30700,N_30708);
nor U31111 (N_31111,N_30121,N_30322);
nand U31112 (N_31112,N_30202,N_30573);
nor U31113 (N_31113,N_30528,N_30692);
or U31114 (N_31114,N_30241,N_30395);
or U31115 (N_31115,N_30579,N_30496);
xor U31116 (N_31116,N_30533,N_30286);
xnor U31117 (N_31117,N_30799,N_30201);
or U31118 (N_31118,N_30018,N_30132);
or U31119 (N_31119,N_30129,N_30214);
nand U31120 (N_31120,N_30796,N_30523);
xnor U31121 (N_31121,N_30632,N_30114);
and U31122 (N_31122,N_30812,N_30596);
nand U31123 (N_31123,N_30838,N_30663);
and U31124 (N_31124,N_30212,N_30671);
nand U31125 (N_31125,N_30781,N_30918);
xor U31126 (N_31126,N_30162,N_30753);
xnor U31127 (N_31127,N_30471,N_30028);
or U31128 (N_31128,N_30283,N_30176);
nor U31129 (N_31129,N_30751,N_30360);
nand U31130 (N_31130,N_30318,N_30874);
nand U31131 (N_31131,N_30586,N_30924);
and U31132 (N_31132,N_30896,N_30031);
or U31133 (N_31133,N_30183,N_30747);
or U31134 (N_31134,N_30589,N_30024);
or U31135 (N_31135,N_30694,N_30506);
xnor U31136 (N_31136,N_30238,N_30402);
or U31137 (N_31137,N_30965,N_30534);
nor U31138 (N_31138,N_30640,N_30367);
xor U31139 (N_31139,N_30997,N_30464);
nor U31140 (N_31140,N_30850,N_30029);
nor U31141 (N_31141,N_30674,N_30603);
nand U31142 (N_31142,N_30250,N_30733);
nor U31143 (N_31143,N_30546,N_30525);
nand U31144 (N_31144,N_30317,N_30845);
or U31145 (N_31145,N_30968,N_30648);
and U31146 (N_31146,N_30020,N_30439);
nor U31147 (N_31147,N_30272,N_30061);
xor U31148 (N_31148,N_30679,N_30999);
nand U31149 (N_31149,N_30219,N_30902);
and U31150 (N_31150,N_30495,N_30268);
and U31151 (N_31151,N_30980,N_30394);
and U31152 (N_31152,N_30750,N_30588);
nor U31153 (N_31153,N_30315,N_30243);
xor U31154 (N_31154,N_30463,N_30161);
or U31155 (N_31155,N_30800,N_30037);
nor U31156 (N_31156,N_30635,N_30729);
and U31157 (N_31157,N_30888,N_30120);
xor U31158 (N_31158,N_30856,N_30156);
nand U31159 (N_31159,N_30867,N_30730);
xnor U31160 (N_31160,N_30088,N_30404);
nand U31161 (N_31161,N_30969,N_30143);
or U31162 (N_31162,N_30184,N_30190);
or U31163 (N_31163,N_30347,N_30152);
nand U31164 (N_31164,N_30014,N_30879);
nand U31165 (N_31165,N_30816,N_30504);
xnor U31166 (N_31166,N_30213,N_30103);
and U31167 (N_31167,N_30487,N_30203);
nand U31168 (N_31168,N_30900,N_30262);
or U31169 (N_31169,N_30085,N_30079);
or U31170 (N_31170,N_30933,N_30456);
and U31171 (N_31171,N_30501,N_30094);
xor U31172 (N_31172,N_30970,N_30821);
or U31173 (N_31173,N_30231,N_30198);
or U31174 (N_31174,N_30769,N_30258);
or U31175 (N_31175,N_30609,N_30461);
nand U31176 (N_31176,N_30366,N_30709);
nor U31177 (N_31177,N_30817,N_30503);
or U31178 (N_31178,N_30319,N_30023);
or U31179 (N_31179,N_30247,N_30672);
nor U31180 (N_31180,N_30113,N_30414);
and U31181 (N_31181,N_30798,N_30167);
nand U31182 (N_31182,N_30788,N_30442);
nand U31183 (N_31183,N_30265,N_30077);
and U31184 (N_31184,N_30689,N_30935);
xnor U31185 (N_31185,N_30144,N_30520);
nor U31186 (N_31186,N_30422,N_30142);
and U31187 (N_31187,N_30150,N_30409);
xor U31188 (N_31188,N_30148,N_30207);
nand U31189 (N_31189,N_30130,N_30140);
nor U31190 (N_31190,N_30361,N_30389);
nand U31191 (N_31191,N_30954,N_30728);
or U31192 (N_31192,N_30543,N_30473);
xor U31193 (N_31193,N_30391,N_30901);
xnor U31194 (N_31194,N_30651,N_30163);
or U31195 (N_31195,N_30059,N_30292);
xnor U31196 (N_31196,N_30793,N_30978);
xor U31197 (N_31197,N_30995,N_30705);
and U31198 (N_31198,N_30403,N_30232);
or U31199 (N_31199,N_30314,N_30147);
or U31200 (N_31200,N_30932,N_30067);
xnor U31201 (N_31201,N_30904,N_30851);
and U31202 (N_31202,N_30134,N_30185);
nor U31203 (N_31203,N_30717,N_30050);
nand U31204 (N_31204,N_30513,N_30127);
or U31205 (N_31205,N_30522,N_30903);
xnor U31206 (N_31206,N_30329,N_30875);
nand U31207 (N_31207,N_30841,N_30189);
nor U31208 (N_31208,N_30594,N_30706);
nor U31209 (N_31209,N_30766,N_30741);
nor U31210 (N_31210,N_30115,N_30313);
and U31211 (N_31211,N_30006,N_30042);
nor U31212 (N_31212,N_30677,N_30457);
and U31213 (N_31213,N_30384,N_30309);
nand U31214 (N_31214,N_30655,N_30714);
nor U31215 (N_31215,N_30581,N_30363);
nor U31216 (N_31216,N_30963,N_30415);
xor U31217 (N_31217,N_30726,N_30387);
nor U31218 (N_31218,N_30790,N_30884);
nand U31219 (N_31219,N_30316,N_30474);
nand U31220 (N_31220,N_30839,N_30041);
or U31221 (N_31221,N_30036,N_30524);
and U31222 (N_31222,N_30260,N_30245);
and U31223 (N_31223,N_30535,N_30626);
and U31224 (N_31224,N_30837,N_30015);
or U31225 (N_31225,N_30814,N_30027);
nand U31226 (N_31226,N_30098,N_30157);
nor U31227 (N_31227,N_30356,N_30767);
xor U31228 (N_31228,N_30477,N_30938);
nand U31229 (N_31229,N_30096,N_30532);
and U31230 (N_31230,N_30470,N_30887);
xnor U31231 (N_31231,N_30302,N_30170);
or U31232 (N_31232,N_30001,N_30369);
xor U31233 (N_31233,N_30237,N_30664);
xor U31234 (N_31234,N_30907,N_30323);
and U31235 (N_31235,N_30072,N_30746);
and U31236 (N_31236,N_30371,N_30564);
or U31237 (N_31237,N_30774,N_30082);
or U31238 (N_31238,N_30340,N_30587);
and U31239 (N_31239,N_30861,N_30691);
and U31240 (N_31240,N_30802,N_30056);
nor U31241 (N_31241,N_30458,N_30852);
nor U31242 (N_31242,N_30792,N_30662);
xor U31243 (N_31243,N_30678,N_30022);
nor U31244 (N_31244,N_30670,N_30226);
nor U31245 (N_31245,N_30481,N_30688);
and U31246 (N_31246,N_30940,N_30857);
or U31247 (N_31247,N_30480,N_30934);
and U31248 (N_31248,N_30035,N_30683);
or U31249 (N_31249,N_30625,N_30338);
and U31250 (N_31250,N_30052,N_30723);
xor U31251 (N_31251,N_30493,N_30572);
and U31252 (N_31252,N_30222,N_30830);
nor U31253 (N_31253,N_30624,N_30443);
or U31254 (N_31254,N_30485,N_30827);
xnor U31255 (N_31255,N_30055,N_30386);
nand U31256 (N_31256,N_30803,N_30686);
nand U31257 (N_31257,N_30290,N_30776);
xor U31258 (N_31258,N_30453,N_30105);
nor U31259 (N_31259,N_30255,N_30514);
nand U31260 (N_31260,N_30922,N_30853);
or U31261 (N_31261,N_30891,N_30945);
nand U31262 (N_31262,N_30012,N_30780);
xor U31263 (N_31263,N_30497,N_30600);
nor U31264 (N_31264,N_30889,N_30771);
nand U31265 (N_31265,N_30131,N_30755);
or U31266 (N_31266,N_30921,N_30249);
nand U31267 (N_31267,N_30601,N_30204);
and U31268 (N_31268,N_30731,N_30472);
xnor U31269 (N_31269,N_30943,N_30383);
nor U31270 (N_31270,N_30787,N_30351);
or U31271 (N_31271,N_30349,N_30125);
nor U31272 (N_31272,N_30342,N_30435);
nor U31273 (N_31273,N_30071,N_30421);
nand U31274 (N_31274,N_30880,N_30892);
nor U31275 (N_31275,N_30177,N_30982);
and U31276 (N_31276,N_30641,N_30578);
nand U31277 (N_31277,N_30937,N_30216);
and U31278 (N_31278,N_30086,N_30873);
xor U31279 (N_31279,N_30136,N_30685);
xor U31280 (N_31280,N_30658,N_30665);
xor U31281 (N_31281,N_30773,N_30378);
xnor U31282 (N_31282,N_30562,N_30293);
nor U31283 (N_31283,N_30808,N_30870);
nor U31284 (N_31284,N_30981,N_30949);
or U31285 (N_31285,N_30192,N_30310);
xnor U31286 (N_31286,N_30300,N_30526);
nand U31287 (N_31287,N_30175,N_30530);
or U31288 (N_31288,N_30436,N_30571);
nor U31289 (N_31289,N_30305,N_30818);
or U31290 (N_31290,N_30124,N_30427);
xor U31291 (N_31291,N_30206,N_30976);
or U31292 (N_31292,N_30872,N_30570);
and U31293 (N_31293,N_30230,N_30673);
or U31294 (N_31294,N_30785,N_30284);
and U31295 (N_31295,N_30652,N_30223);
nand U31296 (N_31296,N_30986,N_30159);
or U31297 (N_31297,N_30307,N_30967);
and U31298 (N_31298,N_30631,N_30303);
xnor U31299 (N_31299,N_30053,N_30273);
and U31300 (N_31300,N_30539,N_30344);
xnor U31301 (N_31301,N_30843,N_30616);
or U31302 (N_31302,N_30939,N_30034);
xor U31303 (N_31303,N_30459,N_30637);
nand U31304 (N_31304,N_30339,N_30445);
xor U31305 (N_31305,N_30576,N_30388);
xnor U31306 (N_31306,N_30509,N_30102);
nor U31307 (N_31307,N_30905,N_30013);
xnor U31308 (N_31308,N_30511,N_30646);
and U31309 (N_31309,N_30083,N_30045);
or U31310 (N_31310,N_30716,N_30362);
xor U31311 (N_31311,N_30288,N_30521);
and U31312 (N_31312,N_30842,N_30979);
nor U31313 (N_31313,N_30772,N_30158);
xor U31314 (N_31314,N_30930,N_30087);
and U31315 (N_31315,N_30431,N_30440);
nand U31316 (N_31316,N_30807,N_30971);
nor U31317 (N_31317,N_30973,N_30629);
or U31318 (N_31318,N_30257,N_30735);
nand U31319 (N_31319,N_30929,N_30187);
nand U31320 (N_31320,N_30432,N_30585);
nand U31321 (N_31321,N_30540,N_30076);
nand U31322 (N_31322,N_30794,N_30135);
xor U31323 (N_31323,N_30119,N_30985);
nor U31324 (N_31324,N_30298,N_30486);
nand U31325 (N_31325,N_30091,N_30660);
nand U31326 (N_31326,N_30848,N_30910);
nor U31327 (N_31327,N_30133,N_30620);
or U31328 (N_31328,N_30615,N_30424);
and U31329 (N_31329,N_30659,N_30770);
nor U31330 (N_31330,N_30172,N_30109);
nand U31331 (N_31331,N_30375,N_30829);
or U31332 (N_31332,N_30081,N_30263);
and U31333 (N_31333,N_30220,N_30991);
nand U31334 (N_31334,N_30667,N_30353);
or U31335 (N_31335,N_30623,N_30491);
and U31336 (N_31336,N_30450,N_30551);
nand U31337 (N_31337,N_30854,N_30101);
nor U31338 (N_31338,N_30775,N_30864);
and U31339 (N_31339,N_30354,N_30153);
and U31340 (N_31340,N_30165,N_30334);
nor U31341 (N_31341,N_30617,N_30447);
nand U31342 (N_31342,N_30401,N_30478);
nor U31343 (N_31343,N_30294,N_30455);
nor U31344 (N_31344,N_30869,N_30619);
and U31345 (N_31345,N_30425,N_30953);
or U31346 (N_31346,N_30680,N_30426);
nor U31347 (N_31347,N_30682,N_30465);
and U31348 (N_31348,N_30266,N_30642);
xnor U31349 (N_31349,N_30374,N_30914);
nor U31350 (N_31350,N_30960,N_30269);
nand U31351 (N_31351,N_30308,N_30186);
nor U31352 (N_31352,N_30380,N_30002);
and U31353 (N_31353,N_30428,N_30112);
or U31354 (N_31354,N_30778,N_30883);
xor U31355 (N_31355,N_30348,N_30221);
nor U31356 (N_31356,N_30505,N_30840);
nor U31357 (N_31357,N_30350,N_30200);
or U31358 (N_31358,N_30337,N_30824);
nor U31359 (N_31359,N_30993,N_30498);
or U31360 (N_31360,N_30650,N_30049);
or U31361 (N_31361,N_30607,N_30998);
and U31362 (N_31362,N_30008,N_30164);
nand U31363 (N_31363,N_30032,N_30448);
and U31364 (N_31364,N_30499,N_30743);
and U31365 (N_31365,N_30645,N_30054);
and U31366 (N_31366,N_30764,N_30936);
nor U31367 (N_31367,N_30866,N_30420);
or U31368 (N_31368,N_30211,N_30275);
nand U31369 (N_31369,N_30759,N_30811);
and U31370 (N_31370,N_30111,N_30761);
xnor U31371 (N_31371,N_30994,N_30545);
nor U31372 (N_31372,N_30711,N_30591);
nor U31373 (N_31373,N_30196,N_30946);
nand U31374 (N_31374,N_30194,N_30003);
and U31375 (N_31375,N_30860,N_30855);
nor U31376 (N_31376,N_30719,N_30955);
and U31377 (N_31377,N_30877,N_30355);
nor U31378 (N_31378,N_30744,N_30359);
nand U31379 (N_31379,N_30868,N_30654);
and U31380 (N_31380,N_30141,N_30742);
and U31381 (N_31381,N_30666,N_30246);
nand U31382 (N_31382,N_30582,N_30561);
xnor U31383 (N_31383,N_30681,N_30698);
xnor U31384 (N_31384,N_30381,N_30878);
and U31385 (N_31385,N_30712,N_30557);
or U31386 (N_31386,N_30370,N_30597);
or U31387 (N_31387,N_30128,N_30462);
nand U31388 (N_31388,N_30429,N_30584);
nand U31389 (N_31389,N_30762,N_30786);
or U31390 (N_31390,N_30927,N_30038);
nor U31391 (N_31391,N_30218,N_30630);
nand U31392 (N_31392,N_30390,N_30618);
or U31393 (N_31393,N_30468,N_30966);
and U31394 (N_31394,N_30756,N_30507);
nor U31395 (N_31395,N_30011,N_30548);
nand U31396 (N_31396,N_30285,N_30416);
xor U31397 (N_31397,N_30400,N_30320);
and U31398 (N_31398,N_30251,N_30075);
nor U31399 (N_31399,N_30229,N_30311);
and U31400 (N_31400,N_30070,N_30026);
and U31401 (N_31401,N_30847,N_30299);
or U31402 (N_31402,N_30365,N_30145);
nand U31403 (N_31403,N_30084,N_30181);
xor U31404 (N_31404,N_30782,N_30598);
xor U31405 (N_31405,N_30208,N_30710);
nor U31406 (N_31406,N_30174,N_30863);
nor U31407 (N_31407,N_30467,N_30553);
or U31408 (N_31408,N_30330,N_30614);
or U31409 (N_31409,N_30988,N_30849);
or U31410 (N_31410,N_30752,N_30763);
nand U31411 (N_31411,N_30916,N_30990);
or U31412 (N_31412,N_30724,N_30123);
xor U31413 (N_31413,N_30702,N_30332);
or U31414 (N_31414,N_30291,N_30754);
and U31415 (N_31415,N_30913,N_30822);
xor U31416 (N_31416,N_30556,N_30306);
xor U31417 (N_31417,N_30690,N_30304);
nand U31418 (N_31418,N_30126,N_30948);
and U31419 (N_31419,N_30040,N_30209);
and U31420 (N_31420,N_30254,N_30984);
or U31421 (N_31421,N_30423,N_30000);
nand U31422 (N_31422,N_30554,N_30276);
and U31423 (N_31423,N_30739,N_30727);
nand U31424 (N_31424,N_30745,N_30612);
or U31425 (N_31425,N_30417,N_30704);
nand U31426 (N_31426,N_30715,N_30494);
and U31427 (N_31427,N_30188,N_30492);
nand U31428 (N_31428,N_30972,N_30909);
nand U31429 (N_31429,N_30489,N_30713);
nand U31430 (N_31430,N_30942,N_30823);
and U31431 (N_31431,N_30326,N_30920);
and U31432 (N_31432,N_30398,N_30516);
nor U31433 (N_31433,N_30518,N_30804);
nor U31434 (N_31434,N_30301,N_30336);
nor U31435 (N_31435,N_30137,N_30166);
and U31436 (N_31436,N_30825,N_30009);
xnor U31437 (N_31437,N_30225,N_30068);
nand U31438 (N_31438,N_30911,N_30168);
nor U31439 (N_31439,N_30718,N_30952);
and U31440 (N_31440,N_30590,N_30668);
and U31441 (N_31441,N_30224,N_30611);
nor U31442 (N_31442,N_30797,N_30765);
and U31443 (N_31443,N_30701,N_30441);
or U31444 (N_31444,N_30894,N_30508);
or U31445 (N_31445,N_30675,N_30016);
xor U31446 (N_31446,N_30264,N_30636);
and U31447 (N_31447,N_30104,N_30095);
xor U31448 (N_31448,N_30100,N_30118);
nor U31449 (N_31449,N_30004,N_30638);
nand U31450 (N_31450,N_30324,N_30433);
and U31451 (N_31451,N_30154,N_30252);
nand U31452 (N_31452,N_30368,N_30419);
xor U31453 (N_31453,N_30364,N_30549);
nor U31454 (N_31454,N_30567,N_30278);
or U31455 (N_31455,N_30828,N_30961);
and U31456 (N_31456,N_30064,N_30890);
xnor U31457 (N_31457,N_30628,N_30449);
nor U31458 (N_31458,N_30406,N_30644);
nor U31459 (N_31459,N_30180,N_30117);
nand U31460 (N_31460,N_30527,N_30197);
nand U31461 (N_31461,N_30602,N_30574);
and U31462 (N_31462,N_30917,N_30836);
nor U31463 (N_31463,N_30080,N_30595);
or U31464 (N_31464,N_30065,N_30613);
nor U31465 (N_31465,N_30171,N_30529);
nor U31466 (N_31466,N_30179,N_30805);
and U31467 (N_31467,N_30732,N_30912);
xnor U31468 (N_31468,N_30779,N_30893);
or U31469 (N_31469,N_30923,N_30722);
and U31470 (N_31470,N_30653,N_30025);
and U31471 (N_31471,N_30227,N_30956);
and U31472 (N_31472,N_30791,N_30408);
and U31473 (N_31473,N_30149,N_30110);
nand U31474 (N_31474,N_30795,N_30605);
xor U31475 (N_31475,N_30078,N_30947);
and U31476 (N_31476,N_30452,N_30622);
nor U31477 (N_31477,N_30720,N_30806);
nand U31478 (N_31478,N_30536,N_30950);
or U31479 (N_31479,N_30577,N_30399);
xor U31480 (N_31480,N_30019,N_30593);
or U31481 (N_31481,N_30289,N_30734);
xor U31482 (N_31482,N_30610,N_30333);
xnor U31483 (N_31483,N_30327,N_30044);
xnor U31484 (N_31484,N_30538,N_30047);
or U31485 (N_31485,N_30451,N_30699);
nor U31486 (N_31486,N_30832,N_30815);
nand U31487 (N_31487,N_30287,N_30325);
or U31488 (N_31488,N_30379,N_30541);
and U31489 (N_31489,N_30633,N_30182);
xnor U31490 (N_31490,N_30295,N_30881);
xnor U31491 (N_31491,N_30908,N_30552);
and U31492 (N_31492,N_30051,N_30108);
nor U31493 (N_31493,N_30030,N_30676);
or U31494 (N_31494,N_30372,N_30649);
or U31495 (N_31495,N_30608,N_30906);
or U31496 (N_31496,N_30057,N_30987);
nand U31497 (N_31497,N_30810,N_30048);
and U31498 (N_31498,N_30758,N_30345);
nor U31499 (N_31499,N_30941,N_30575);
and U31500 (N_31500,N_30760,N_30891);
xnor U31501 (N_31501,N_30305,N_30070);
and U31502 (N_31502,N_30458,N_30902);
nor U31503 (N_31503,N_30421,N_30699);
xor U31504 (N_31504,N_30713,N_30746);
nor U31505 (N_31505,N_30324,N_30732);
or U31506 (N_31506,N_30151,N_30421);
nand U31507 (N_31507,N_30552,N_30001);
xor U31508 (N_31508,N_30300,N_30593);
and U31509 (N_31509,N_30113,N_30657);
or U31510 (N_31510,N_30233,N_30771);
or U31511 (N_31511,N_30274,N_30554);
and U31512 (N_31512,N_30661,N_30153);
nor U31513 (N_31513,N_30984,N_30370);
or U31514 (N_31514,N_30330,N_30058);
and U31515 (N_31515,N_30747,N_30686);
and U31516 (N_31516,N_30678,N_30327);
nor U31517 (N_31517,N_30747,N_30390);
nor U31518 (N_31518,N_30495,N_30413);
xnor U31519 (N_31519,N_30815,N_30646);
and U31520 (N_31520,N_30869,N_30080);
xor U31521 (N_31521,N_30504,N_30786);
nor U31522 (N_31522,N_30583,N_30006);
and U31523 (N_31523,N_30736,N_30812);
xor U31524 (N_31524,N_30176,N_30804);
and U31525 (N_31525,N_30057,N_30288);
or U31526 (N_31526,N_30210,N_30774);
nand U31527 (N_31527,N_30955,N_30133);
or U31528 (N_31528,N_30515,N_30661);
or U31529 (N_31529,N_30642,N_30371);
nor U31530 (N_31530,N_30173,N_30381);
nor U31531 (N_31531,N_30556,N_30992);
nor U31532 (N_31532,N_30633,N_30118);
or U31533 (N_31533,N_30981,N_30174);
xnor U31534 (N_31534,N_30255,N_30287);
nand U31535 (N_31535,N_30585,N_30421);
or U31536 (N_31536,N_30881,N_30411);
nor U31537 (N_31537,N_30733,N_30561);
nor U31538 (N_31538,N_30281,N_30928);
and U31539 (N_31539,N_30507,N_30521);
nor U31540 (N_31540,N_30264,N_30368);
and U31541 (N_31541,N_30646,N_30678);
or U31542 (N_31542,N_30495,N_30896);
nor U31543 (N_31543,N_30128,N_30428);
or U31544 (N_31544,N_30031,N_30597);
and U31545 (N_31545,N_30113,N_30319);
nor U31546 (N_31546,N_30838,N_30555);
nand U31547 (N_31547,N_30385,N_30032);
xor U31548 (N_31548,N_30408,N_30192);
xnor U31549 (N_31549,N_30253,N_30625);
xnor U31550 (N_31550,N_30860,N_30390);
or U31551 (N_31551,N_30893,N_30074);
xor U31552 (N_31552,N_30735,N_30532);
nor U31553 (N_31553,N_30006,N_30388);
nand U31554 (N_31554,N_30120,N_30905);
and U31555 (N_31555,N_30812,N_30906);
nor U31556 (N_31556,N_30486,N_30805);
and U31557 (N_31557,N_30844,N_30144);
nor U31558 (N_31558,N_30560,N_30399);
or U31559 (N_31559,N_30932,N_30442);
xor U31560 (N_31560,N_30922,N_30980);
or U31561 (N_31561,N_30220,N_30877);
or U31562 (N_31562,N_30381,N_30376);
xnor U31563 (N_31563,N_30971,N_30006);
xor U31564 (N_31564,N_30671,N_30033);
nor U31565 (N_31565,N_30699,N_30121);
nand U31566 (N_31566,N_30383,N_30704);
xnor U31567 (N_31567,N_30530,N_30098);
or U31568 (N_31568,N_30040,N_30211);
or U31569 (N_31569,N_30626,N_30157);
nand U31570 (N_31570,N_30890,N_30528);
nor U31571 (N_31571,N_30972,N_30523);
nand U31572 (N_31572,N_30229,N_30934);
nand U31573 (N_31573,N_30027,N_30396);
xnor U31574 (N_31574,N_30645,N_30479);
or U31575 (N_31575,N_30849,N_30720);
or U31576 (N_31576,N_30686,N_30064);
nor U31577 (N_31577,N_30349,N_30957);
nand U31578 (N_31578,N_30223,N_30605);
and U31579 (N_31579,N_30298,N_30558);
or U31580 (N_31580,N_30647,N_30455);
or U31581 (N_31581,N_30198,N_30949);
nand U31582 (N_31582,N_30599,N_30106);
or U31583 (N_31583,N_30733,N_30677);
nand U31584 (N_31584,N_30936,N_30913);
nor U31585 (N_31585,N_30425,N_30305);
nand U31586 (N_31586,N_30139,N_30279);
or U31587 (N_31587,N_30602,N_30062);
nand U31588 (N_31588,N_30451,N_30752);
nand U31589 (N_31589,N_30455,N_30082);
and U31590 (N_31590,N_30914,N_30285);
nor U31591 (N_31591,N_30052,N_30147);
or U31592 (N_31592,N_30662,N_30699);
nand U31593 (N_31593,N_30385,N_30588);
nand U31594 (N_31594,N_30078,N_30517);
nor U31595 (N_31595,N_30615,N_30707);
and U31596 (N_31596,N_30739,N_30305);
nor U31597 (N_31597,N_30155,N_30028);
nand U31598 (N_31598,N_30525,N_30982);
and U31599 (N_31599,N_30129,N_30269);
or U31600 (N_31600,N_30772,N_30085);
nand U31601 (N_31601,N_30385,N_30708);
nor U31602 (N_31602,N_30082,N_30300);
nor U31603 (N_31603,N_30568,N_30945);
xnor U31604 (N_31604,N_30497,N_30599);
xnor U31605 (N_31605,N_30027,N_30398);
xnor U31606 (N_31606,N_30341,N_30838);
nor U31607 (N_31607,N_30782,N_30472);
nor U31608 (N_31608,N_30591,N_30737);
nand U31609 (N_31609,N_30333,N_30070);
and U31610 (N_31610,N_30074,N_30147);
or U31611 (N_31611,N_30035,N_30433);
and U31612 (N_31612,N_30367,N_30488);
nand U31613 (N_31613,N_30424,N_30774);
nand U31614 (N_31614,N_30918,N_30240);
nor U31615 (N_31615,N_30201,N_30851);
xnor U31616 (N_31616,N_30187,N_30636);
or U31617 (N_31617,N_30406,N_30898);
nand U31618 (N_31618,N_30458,N_30280);
or U31619 (N_31619,N_30370,N_30570);
nand U31620 (N_31620,N_30483,N_30482);
and U31621 (N_31621,N_30285,N_30874);
or U31622 (N_31622,N_30088,N_30253);
or U31623 (N_31623,N_30282,N_30157);
nor U31624 (N_31624,N_30676,N_30525);
or U31625 (N_31625,N_30040,N_30154);
xnor U31626 (N_31626,N_30746,N_30533);
and U31627 (N_31627,N_30753,N_30328);
nand U31628 (N_31628,N_30900,N_30267);
xor U31629 (N_31629,N_30098,N_30118);
nor U31630 (N_31630,N_30600,N_30912);
xnor U31631 (N_31631,N_30402,N_30330);
xnor U31632 (N_31632,N_30017,N_30194);
and U31633 (N_31633,N_30903,N_30478);
and U31634 (N_31634,N_30220,N_30082);
or U31635 (N_31635,N_30916,N_30695);
and U31636 (N_31636,N_30460,N_30832);
and U31637 (N_31637,N_30923,N_30735);
or U31638 (N_31638,N_30260,N_30684);
or U31639 (N_31639,N_30290,N_30345);
nand U31640 (N_31640,N_30304,N_30393);
and U31641 (N_31641,N_30666,N_30702);
and U31642 (N_31642,N_30627,N_30019);
nor U31643 (N_31643,N_30377,N_30353);
xnor U31644 (N_31644,N_30157,N_30782);
nor U31645 (N_31645,N_30731,N_30760);
xor U31646 (N_31646,N_30926,N_30180);
xnor U31647 (N_31647,N_30393,N_30271);
nor U31648 (N_31648,N_30384,N_30520);
and U31649 (N_31649,N_30492,N_30176);
nand U31650 (N_31650,N_30099,N_30491);
or U31651 (N_31651,N_30085,N_30914);
xnor U31652 (N_31652,N_30707,N_30476);
nand U31653 (N_31653,N_30959,N_30051);
nor U31654 (N_31654,N_30235,N_30212);
or U31655 (N_31655,N_30077,N_30083);
nor U31656 (N_31656,N_30973,N_30323);
and U31657 (N_31657,N_30483,N_30709);
nor U31658 (N_31658,N_30279,N_30036);
or U31659 (N_31659,N_30848,N_30049);
or U31660 (N_31660,N_30996,N_30330);
xnor U31661 (N_31661,N_30877,N_30461);
nand U31662 (N_31662,N_30375,N_30931);
xnor U31663 (N_31663,N_30568,N_30742);
nand U31664 (N_31664,N_30612,N_30210);
nor U31665 (N_31665,N_30200,N_30261);
and U31666 (N_31666,N_30009,N_30636);
nor U31667 (N_31667,N_30239,N_30879);
or U31668 (N_31668,N_30500,N_30757);
xnor U31669 (N_31669,N_30869,N_30097);
xnor U31670 (N_31670,N_30165,N_30635);
and U31671 (N_31671,N_30126,N_30529);
xnor U31672 (N_31672,N_30909,N_30268);
nor U31673 (N_31673,N_30476,N_30125);
nand U31674 (N_31674,N_30927,N_30052);
xnor U31675 (N_31675,N_30679,N_30682);
nand U31676 (N_31676,N_30279,N_30402);
xor U31677 (N_31677,N_30226,N_30393);
nand U31678 (N_31678,N_30404,N_30512);
nand U31679 (N_31679,N_30503,N_30461);
nor U31680 (N_31680,N_30394,N_30794);
nand U31681 (N_31681,N_30430,N_30946);
or U31682 (N_31682,N_30434,N_30558);
xor U31683 (N_31683,N_30054,N_30782);
nand U31684 (N_31684,N_30519,N_30456);
and U31685 (N_31685,N_30526,N_30431);
nand U31686 (N_31686,N_30396,N_30285);
and U31687 (N_31687,N_30555,N_30377);
xnor U31688 (N_31688,N_30205,N_30383);
or U31689 (N_31689,N_30020,N_30039);
or U31690 (N_31690,N_30272,N_30930);
nand U31691 (N_31691,N_30652,N_30763);
nor U31692 (N_31692,N_30853,N_30197);
or U31693 (N_31693,N_30787,N_30053);
xor U31694 (N_31694,N_30527,N_30876);
nor U31695 (N_31695,N_30622,N_30516);
xor U31696 (N_31696,N_30493,N_30517);
nor U31697 (N_31697,N_30307,N_30886);
nand U31698 (N_31698,N_30742,N_30262);
nor U31699 (N_31699,N_30735,N_30370);
xor U31700 (N_31700,N_30820,N_30000);
nor U31701 (N_31701,N_30357,N_30978);
and U31702 (N_31702,N_30942,N_30811);
or U31703 (N_31703,N_30343,N_30820);
xnor U31704 (N_31704,N_30501,N_30942);
nor U31705 (N_31705,N_30462,N_30794);
or U31706 (N_31706,N_30722,N_30174);
xor U31707 (N_31707,N_30607,N_30796);
nor U31708 (N_31708,N_30287,N_30327);
or U31709 (N_31709,N_30486,N_30465);
and U31710 (N_31710,N_30804,N_30540);
nor U31711 (N_31711,N_30945,N_30958);
xor U31712 (N_31712,N_30109,N_30992);
or U31713 (N_31713,N_30507,N_30788);
xor U31714 (N_31714,N_30321,N_30716);
xor U31715 (N_31715,N_30339,N_30517);
nor U31716 (N_31716,N_30827,N_30628);
nand U31717 (N_31717,N_30793,N_30745);
and U31718 (N_31718,N_30776,N_30011);
xnor U31719 (N_31719,N_30110,N_30432);
and U31720 (N_31720,N_30935,N_30787);
and U31721 (N_31721,N_30676,N_30755);
nand U31722 (N_31722,N_30737,N_30121);
and U31723 (N_31723,N_30440,N_30956);
nor U31724 (N_31724,N_30252,N_30083);
and U31725 (N_31725,N_30732,N_30539);
and U31726 (N_31726,N_30515,N_30440);
nor U31727 (N_31727,N_30039,N_30947);
nand U31728 (N_31728,N_30703,N_30103);
nor U31729 (N_31729,N_30371,N_30603);
and U31730 (N_31730,N_30375,N_30014);
nand U31731 (N_31731,N_30730,N_30654);
and U31732 (N_31732,N_30582,N_30815);
nand U31733 (N_31733,N_30662,N_30900);
and U31734 (N_31734,N_30330,N_30970);
and U31735 (N_31735,N_30364,N_30255);
or U31736 (N_31736,N_30916,N_30778);
and U31737 (N_31737,N_30460,N_30468);
nand U31738 (N_31738,N_30457,N_30534);
nand U31739 (N_31739,N_30638,N_30947);
and U31740 (N_31740,N_30178,N_30530);
or U31741 (N_31741,N_30548,N_30947);
xor U31742 (N_31742,N_30791,N_30402);
or U31743 (N_31743,N_30159,N_30690);
nor U31744 (N_31744,N_30006,N_30060);
nor U31745 (N_31745,N_30592,N_30310);
nor U31746 (N_31746,N_30176,N_30985);
and U31747 (N_31747,N_30875,N_30522);
and U31748 (N_31748,N_30909,N_30851);
and U31749 (N_31749,N_30522,N_30808);
xor U31750 (N_31750,N_30590,N_30145);
nand U31751 (N_31751,N_30225,N_30465);
or U31752 (N_31752,N_30152,N_30129);
and U31753 (N_31753,N_30621,N_30858);
and U31754 (N_31754,N_30698,N_30405);
xor U31755 (N_31755,N_30758,N_30733);
or U31756 (N_31756,N_30237,N_30788);
xnor U31757 (N_31757,N_30925,N_30150);
and U31758 (N_31758,N_30819,N_30852);
nor U31759 (N_31759,N_30761,N_30032);
nand U31760 (N_31760,N_30579,N_30096);
or U31761 (N_31761,N_30809,N_30701);
nor U31762 (N_31762,N_30799,N_30560);
or U31763 (N_31763,N_30762,N_30675);
xnor U31764 (N_31764,N_30089,N_30805);
xnor U31765 (N_31765,N_30890,N_30405);
or U31766 (N_31766,N_30682,N_30819);
nor U31767 (N_31767,N_30810,N_30589);
and U31768 (N_31768,N_30321,N_30126);
xnor U31769 (N_31769,N_30220,N_30729);
and U31770 (N_31770,N_30477,N_30529);
or U31771 (N_31771,N_30173,N_30793);
or U31772 (N_31772,N_30858,N_30191);
nor U31773 (N_31773,N_30641,N_30500);
nor U31774 (N_31774,N_30372,N_30714);
nor U31775 (N_31775,N_30982,N_30381);
xor U31776 (N_31776,N_30579,N_30392);
nor U31777 (N_31777,N_30553,N_30693);
and U31778 (N_31778,N_30740,N_30046);
and U31779 (N_31779,N_30150,N_30388);
nor U31780 (N_31780,N_30742,N_30819);
nand U31781 (N_31781,N_30277,N_30167);
or U31782 (N_31782,N_30933,N_30195);
xor U31783 (N_31783,N_30024,N_30355);
or U31784 (N_31784,N_30718,N_30682);
nor U31785 (N_31785,N_30016,N_30962);
nor U31786 (N_31786,N_30576,N_30991);
and U31787 (N_31787,N_30215,N_30591);
and U31788 (N_31788,N_30310,N_30308);
and U31789 (N_31789,N_30318,N_30160);
xor U31790 (N_31790,N_30932,N_30000);
xor U31791 (N_31791,N_30124,N_30020);
or U31792 (N_31792,N_30993,N_30411);
and U31793 (N_31793,N_30625,N_30024);
or U31794 (N_31794,N_30625,N_30049);
and U31795 (N_31795,N_30166,N_30804);
nor U31796 (N_31796,N_30357,N_30555);
xor U31797 (N_31797,N_30489,N_30977);
and U31798 (N_31798,N_30319,N_30833);
or U31799 (N_31799,N_30563,N_30665);
xnor U31800 (N_31800,N_30912,N_30513);
xnor U31801 (N_31801,N_30967,N_30248);
and U31802 (N_31802,N_30448,N_30606);
and U31803 (N_31803,N_30245,N_30250);
and U31804 (N_31804,N_30086,N_30809);
or U31805 (N_31805,N_30044,N_30439);
nor U31806 (N_31806,N_30610,N_30539);
and U31807 (N_31807,N_30361,N_30841);
xnor U31808 (N_31808,N_30402,N_30587);
xor U31809 (N_31809,N_30017,N_30687);
nor U31810 (N_31810,N_30554,N_30397);
nand U31811 (N_31811,N_30727,N_30864);
nor U31812 (N_31812,N_30170,N_30608);
nor U31813 (N_31813,N_30001,N_30338);
and U31814 (N_31814,N_30165,N_30361);
xnor U31815 (N_31815,N_30574,N_30914);
nand U31816 (N_31816,N_30075,N_30696);
or U31817 (N_31817,N_30424,N_30032);
nor U31818 (N_31818,N_30288,N_30867);
or U31819 (N_31819,N_30364,N_30534);
xor U31820 (N_31820,N_30858,N_30349);
nand U31821 (N_31821,N_30881,N_30739);
or U31822 (N_31822,N_30058,N_30690);
nand U31823 (N_31823,N_30250,N_30617);
xnor U31824 (N_31824,N_30692,N_30286);
nand U31825 (N_31825,N_30470,N_30226);
xnor U31826 (N_31826,N_30156,N_30104);
or U31827 (N_31827,N_30403,N_30934);
and U31828 (N_31828,N_30056,N_30083);
xnor U31829 (N_31829,N_30178,N_30734);
xor U31830 (N_31830,N_30905,N_30634);
nand U31831 (N_31831,N_30789,N_30873);
or U31832 (N_31832,N_30331,N_30297);
and U31833 (N_31833,N_30508,N_30486);
or U31834 (N_31834,N_30932,N_30340);
and U31835 (N_31835,N_30322,N_30049);
and U31836 (N_31836,N_30724,N_30814);
nand U31837 (N_31837,N_30839,N_30169);
xor U31838 (N_31838,N_30900,N_30905);
xnor U31839 (N_31839,N_30004,N_30444);
nor U31840 (N_31840,N_30865,N_30811);
or U31841 (N_31841,N_30831,N_30991);
xnor U31842 (N_31842,N_30504,N_30733);
xor U31843 (N_31843,N_30181,N_30629);
xnor U31844 (N_31844,N_30532,N_30132);
or U31845 (N_31845,N_30391,N_30323);
and U31846 (N_31846,N_30466,N_30536);
nor U31847 (N_31847,N_30847,N_30298);
and U31848 (N_31848,N_30882,N_30841);
or U31849 (N_31849,N_30125,N_30102);
nand U31850 (N_31850,N_30909,N_30926);
and U31851 (N_31851,N_30569,N_30824);
or U31852 (N_31852,N_30025,N_30941);
nand U31853 (N_31853,N_30567,N_30540);
nor U31854 (N_31854,N_30732,N_30249);
or U31855 (N_31855,N_30282,N_30172);
or U31856 (N_31856,N_30430,N_30344);
or U31857 (N_31857,N_30796,N_30593);
nor U31858 (N_31858,N_30625,N_30676);
xnor U31859 (N_31859,N_30646,N_30106);
and U31860 (N_31860,N_30435,N_30780);
nand U31861 (N_31861,N_30281,N_30353);
or U31862 (N_31862,N_30705,N_30680);
nand U31863 (N_31863,N_30293,N_30726);
nor U31864 (N_31864,N_30550,N_30746);
and U31865 (N_31865,N_30904,N_30074);
and U31866 (N_31866,N_30298,N_30195);
and U31867 (N_31867,N_30756,N_30589);
or U31868 (N_31868,N_30595,N_30020);
or U31869 (N_31869,N_30640,N_30305);
nor U31870 (N_31870,N_30804,N_30159);
and U31871 (N_31871,N_30540,N_30551);
xor U31872 (N_31872,N_30348,N_30423);
and U31873 (N_31873,N_30730,N_30181);
nand U31874 (N_31874,N_30438,N_30479);
xnor U31875 (N_31875,N_30282,N_30121);
nor U31876 (N_31876,N_30454,N_30009);
nand U31877 (N_31877,N_30898,N_30631);
xnor U31878 (N_31878,N_30944,N_30085);
nand U31879 (N_31879,N_30418,N_30641);
nand U31880 (N_31880,N_30120,N_30428);
and U31881 (N_31881,N_30894,N_30802);
or U31882 (N_31882,N_30909,N_30625);
or U31883 (N_31883,N_30352,N_30461);
nand U31884 (N_31884,N_30105,N_30509);
and U31885 (N_31885,N_30310,N_30762);
nand U31886 (N_31886,N_30439,N_30043);
xor U31887 (N_31887,N_30928,N_30328);
nand U31888 (N_31888,N_30596,N_30509);
or U31889 (N_31889,N_30461,N_30110);
nor U31890 (N_31890,N_30641,N_30232);
nand U31891 (N_31891,N_30001,N_30287);
xnor U31892 (N_31892,N_30649,N_30609);
nand U31893 (N_31893,N_30806,N_30243);
and U31894 (N_31894,N_30274,N_30241);
nor U31895 (N_31895,N_30631,N_30191);
xnor U31896 (N_31896,N_30371,N_30668);
or U31897 (N_31897,N_30980,N_30126);
or U31898 (N_31898,N_30419,N_30755);
xor U31899 (N_31899,N_30479,N_30047);
or U31900 (N_31900,N_30046,N_30094);
and U31901 (N_31901,N_30211,N_30442);
or U31902 (N_31902,N_30311,N_30716);
and U31903 (N_31903,N_30327,N_30047);
xnor U31904 (N_31904,N_30532,N_30318);
or U31905 (N_31905,N_30866,N_30328);
nand U31906 (N_31906,N_30625,N_30863);
nand U31907 (N_31907,N_30160,N_30968);
and U31908 (N_31908,N_30607,N_30591);
nand U31909 (N_31909,N_30360,N_30870);
nand U31910 (N_31910,N_30951,N_30147);
nor U31911 (N_31911,N_30344,N_30963);
and U31912 (N_31912,N_30267,N_30481);
and U31913 (N_31913,N_30787,N_30734);
or U31914 (N_31914,N_30803,N_30624);
and U31915 (N_31915,N_30123,N_30252);
nand U31916 (N_31916,N_30523,N_30030);
nand U31917 (N_31917,N_30167,N_30179);
and U31918 (N_31918,N_30043,N_30123);
and U31919 (N_31919,N_30680,N_30807);
nor U31920 (N_31920,N_30628,N_30485);
xor U31921 (N_31921,N_30583,N_30030);
xor U31922 (N_31922,N_30665,N_30670);
nand U31923 (N_31923,N_30130,N_30944);
xnor U31924 (N_31924,N_30861,N_30997);
xnor U31925 (N_31925,N_30110,N_30134);
and U31926 (N_31926,N_30116,N_30123);
and U31927 (N_31927,N_30203,N_30425);
nand U31928 (N_31928,N_30623,N_30463);
and U31929 (N_31929,N_30952,N_30866);
nand U31930 (N_31930,N_30634,N_30449);
nand U31931 (N_31931,N_30436,N_30414);
or U31932 (N_31932,N_30769,N_30953);
and U31933 (N_31933,N_30482,N_30110);
and U31934 (N_31934,N_30805,N_30728);
and U31935 (N_31935,N_30567,N_30565);
nor U31936 (N_31936,N_30381,N_30992);
nand U31937 (N_31937,N_30311,N_30068);
or U31938 (N_31938,N_30313,N_30482);
nand U31939 (N_31939,N_30003,N_30005);
nor U31940 (N_31940,N_30872,N_30877);
nand U31941 (N_31941,N_30192,N_30777);
xor U31942 (N_31942,N_30893,N_30081);
nand U31943 (N_31943,N_30601,N_30928);
nor U31944 (N_31944,N_30623,N_30214);
xor U31945 (N_31945,N_30107,N_30598);
nor U31946 (N_31946,N_30634,N_30909);
nor U31947 (N_31947,N_30929,N_30235);
xnor U31948 (N_31948,N_30163,N_30860);
or U31949 (N_31949,N_30317,N_30761);
nand U31950 (N_31950,N_30527,N_30914);
or U31951 (N_31951,N_30418,N_30971);
nor U31952 (N_31952,N_30394,N_30874);
nand U31953 (N_31953,N_30547,N_30140);
or U31954 (N_31954,N_30423,N_30205);
or U31955 (N_31955,N_30878,N_30998);
nand U31956 (N_31956,N_30318,N_30760);
or U31957 (N_31957,N_30384,N_30880);
and U31958 (N_31958,N_30021,N_30666);
nand U31959 (N_31959,N_30660,N_30445);
nand U31960 (N_31960,N_30011,N_30242);
nand U31961 (N_31961,N_30256,N_30992);
xor U31962 (N_31962,N_30360,N_30621);
and U31963 (N_31963,N_30533,N_30495);
or U31964 (N_31964,N_30089,N_30930);
and U31965 (N_31965,N_30263,N_30553);
xnor U31966 (N_31966,N_30811,N_30099);
nor U31967 (N_31967,N_30973,N_30158);
xnor U31968 (N_31968,N_30300,N_30722);
or U31969 (N_31969,N_30541,N_30445);
xnor U31970 (N_31970,N_30378,N_30114);
nand U31971 (N_31971,N_30259,N_30575);
nand U31972 (N_31972,N_30963,N_30138);
or U31973 (N_31973,N_30284,N_30600);
xor U31974 (N_31974,N_30168,N_30763);
and U31975 (N_31975,N_30993,N_30060);
nand U31976 (N_31976,N_30108,N_30040);
nor U31977 (N_31977,N_30079,N_30564);
xnor U31978 (N_31978,N_30679,N_30972);
and U31979 (N_31979,N_30067,N_30830);
nor U31980 (N_31980,N_30665,N_30793);
nor U31981 (N_31981,N_30084,N_30271);
nor U31982 (N_31982,N_30271,N_30432);
or U31983 (N_31983,N_30694,N_30402);
nand U31984 (N_31984,N_30150,N_30491);
xnor U31985 (N_31985,N_30580,N_30523);
nand U31986 (N_31986,N_30399,N_30206);
and U31987 (N_31987,N_30646,N_30528);
xor U31988 (N_31988,N_30248,N_30448);
nor U31989 (N_31989,N_30955,N_30957);
xor U31990 (N_31990,N_30057,N_30496);
nand U31991 (N_31991,N_30375,N_30021);
nand U31992 (N_31992,N_30479,N_30311);
nor U31993 (N_31993,N_30578,N_30598);
nand U31994 (N_31994,N_30403,N_30117);
or U31995 (N_31995,N_30057,N_30941);
nor U31996 (N_31996,N_30482,N_30591);
or U31997 (N_31997,N_30965,N_30583);
nand U31998 (N_31998,N_30300,N_30658);
and U31999 (N_31999,N_30254,N_30796);
nor U32000 (N_32000,N_31594,N_31558);
or U32001 (N_32001,N_31843,N_31503);
nand U32002 (N_32002,N_31160,N_31190);
and U32003 (N_32003,N_31880,N_31523);
nor U32004 (N_32004,N_31274,N_31159);
nand U32005 (N_32005,N_31429,N_31355);
nor U32006 (N_32006,N_31587,N_31833);
and U32007 (N_32007,N_31845,N_31075);
nand U32008 (N_32008,N_31773,N_31704);
nand U32009 (N_32009,N_31570,N_31488);
xor U32010 (N_32010,N_31179,N_31306);
nor U32011 (N_32011,N_31313,N_31433);
xnor U32012 (N_32012,N_31049,N_31392);
xnor U32013 (N_32013,N_31475,N_31099);
nor U32014 (N_32014,N_31838,N_31143);
nand U32015 (N_32015,N_31489,N_31320);
and U32016 (N_32016,N_31243,N_31809);
or U32017 (N_32017,N_31039,N_31056);
nor U32018 (N_32018,N_31032,N_31789);
nand U32019 (N_32019,N_31172,N_31742);
xnor U32020 (N_32020,N_31051,N_31768);
or U32021 (N_32021,N_31074,N_31364);
xnor U32022 (N_32022,N_31869,N_31389);
xnor U32023 (N_32023,N_31563,N_31571);
or U32024 (N_32024,N_31264,N_31628);
and U32025 (N_32025,N_31346,N_31211);
xor U32026 (N_32026,N_31971,N_31513);
xnor U32027 (N_32027,N_31886,N_31480);
and U32028 (N_32028,N_31082,N_31610);
and U32029 (N_32029,N_31341,N_31678);
nor U32030 (N_32030,N_31291,N_31194);
nand U32031 (N_32031,N_31506,N_31481);
nand U32032 (N_32032,N_31538,N_31415);
nor U32033 (N_32033,N_31474,N_31321);
nor U32034 (N_32034,N_31517,N_31634);
nor U32035 (N_32035,N_31713,N_31707);
nor U32036 (N_32036,N_31424,N_31081);
nand U32037 (N_32037,N_31453,N_31684);
xor U32038 (N_32038,N_31496,N_31230);
nor U32039 (N_32039,N_31013,N_31755);
and U32040 (N_32040,N_31554,N_31533);
xor U32041 (N_32041,N_31125,N_31458);
nand U32042 (N_32042,N_31246,N_31624);
nor U32043 (N_32043,N_31893,N_31991);
xnor U32044 (N_32044,N_31717,N_31912);
xnor U32045 (N_32045,N_31526,N_31823);
nand U32046 (N_32046,N_31793,N_31757);
and U32047 (N_32047,N_31418,N_31253);
xnor U32048 (N_32048,N_31780,N_31305);
and U32049 (N_32049,N_31941,N_31302);
nor U32050 (N_32050,N_31339,N_31808);
nand U32051 (N_32051,N_31701,N_31783);
or U32052 (N_32052,N_31703,N_31592);
and U32053 (N_32053,N_31981,N_31297);
and U32054 (N_32054,N_31955,N_31419);
and U32055 (N_32055,N_31390,N_31093);
xor U32056 (N_32056,N_31128,N_31402);
or U32057 (N_32057,N_31180,N_31799);
xnor U32058 (N_32058,N_31969,N_31575);
or U32059 (N_32059,N_31831,N_31500);
nor U32060 (N_32060,N_31650,N_31316);
nand U32061 (N_32061,N_31792,N_31658);
and U32062 (N_32062,N_31622,N_31399);
nand U32063 (N_32063,N_31599,N_31353);
xor U32064 (N_32064,N_31328,N_31784);
nand U32065 (N_32065,N_31655,N_31851);
nor U32066 (N_32066,N_31936,N_31370);
nor U32067 (N_32067,N_31478,N_31131);
xor U32068 (N_32068,N_31763,N_31537);
nor U32069 (N_32069,N_31816,N_31426);
and U32070 (N_32070,N_31470,N_31414);
xor U32071 (N_32071,N_31281,N_31300);
and U32072 (N_32072,N_31127,N_31031);
or U32073 (N_32073,N_31174,N_31868);
xnor U32074 (N_32074,N_31956,N_31293);
and U32075 (N_32075,N_31645,N_31195);
nor U32076 (N_32076,N_31050,N_31609);
nand U32077 (N_32077,N_31986,N_31895);
and U32078 (N_32078,N_31173,N_31689);
nor U32079 (N_32079,N_31114,N_31120);
nand U32080 (N_32080,N_31800,N_31657);
and U32081 (N_32081,N_31410,N_31830);
nand U32082 (N_32082,N_31731,N_31934);
nand U32083 (N_32083,N_31853,N_31349);
nand U32084 (N_32084,N_31303,N_31983);
or U32085 (N_32085,N_31358,N_31591);
xor U32086 (N_32086,N_31254,N_31191);
nor U32087 (N_32087,N_31965,N_31666);
nor U32088 (N_32088,N_31437,N_31862);
xor U32089 (N_32089,N_31069,N_31728);
or U32090 (N_32090,N_31690,N_31098);
nand U32091 (N_32091,N_31648,N_31425);
xor U32092 (N_32092,N_31372,N_31807);
nor U32093 (N_32093,N_31957,N_31361);
nand U32094 (N_32094,N_31858,N_31637);
nand U32095 (N_32095,N_31146,N_31597);
xor U32096 (N_32096,N_31483,N_31711);
or U32097 (N_32097,N_31931,N_31686);
nand U32098 (N_32098,N_31933,N_31497);
xnor U32099 (N_32099,N_31382,N_31391);
xor U32100 (N_32100,N_31046,N_31201);
and U32101 (N_32101,N_31982,N_31884);
nor U32102 (N_32102,N_31164,N_31631);
or U32103 (N_32103,N_31452,N_31920);
or U32104 (N_32104,N_31451,N_31815);
and U32105 (N_32105,N_31771,N_31133);
xnor U32106 (N_32106,N_31535,N_31136);
and U32107 (N_32107,N_31737,N_31457);
nand U32108 (N_32108,N_31882,N_31756);
xor U32109 (N_32109,N_31897,N_31092);
nand U32110 (N_32110,N_31566,N_31939);
xor U32111 (N_32111,N_31840,N_31747);
nand U32112 (N_32112,N_31058,N_31232);
nor U32113 (N_32113,N_31235,N_31922);
or U32114 (N_32114,N_31411,N_31450);
or U32115 (N_32115,N_31345,N_31687);
nand U32116 (N_32116,N_31902,N_31903);
nand U32117 (N_32117,N_31221,N_31002);
xor U32118 (N_32118,N_31205,N_31354);
nand U32119 (N_32119,N_31233,N_31826);
nand U32120 (N_32120,N_31852,N_31007);
nor U32121 (N_32121,N_31829,N_31071);
xor U32122 (N_32122,N_31342,N_31124);
or U32123 (N_32123,N_31461,N_31065);
and U32124 (N_32124,N_31151,N_31428);
and U32125 (N_32125,N_31109,N_31511);
nand U32126 (N_32126,N_31224,N_31856);
xor U32127 (N_32127,N_31870,N_31219);
nor U32128 (N_32128,N_31887,N_31844);
xor U32129 (N_32129,N_31619,N_31268);
nor U32130 (N_32130,N_31598,N_31629);
xor U32131 (N_32131,N_31968,N_31204);
nor U32132 (N_32132,N_31006,N_31021);
or U32133 (N_32133,N_31163,N_31691);
and U32134 (N_32134,N_31277,N_31604);
or U32135 (N_32135,N_31162,N_31288);
nor U32136 (N_32136,N_31603,N_31144);
nand U32137 (N_32137,N_31958,N_31175);
nor U32138 (N_32138,N_31168,N_31197);
and U32139 (N_32139,N_31256,N_31948);
nand U32140 (N_32140,N_31576,N_31189);
nand U32141 (N_32141,N_31859,N_31677);
and U32142 (N_32142,N_31652,N_31601);
xor U32143 (N_32143,N_31329,N_31123);
nand U32144 (N_32144,N_31664,N_31207);
nor U32145 (N_32145,N_31745,N_31000);
nor U32146 (N_32146,N_31181,N_31644);
nand U32147 (N_32147,N_31245,N_31748);
and U32148 (N_32148,N_31097,N_31605);
nand U32149 (N_32149,N_31375,N_31251);
nor U32150 (N_32150,N_31423,N_31085);
nand U32151 (N_32151,N_31149,N_31896);
nor U32152 (N_32152,N_31030,N_31953);
and U32153 (N_32153,N_31072,N_31834);
and U32154 (N_32154,N_31924,N_31805);
xor U32155 (N_32155,N_31660,N_31141);
and U32156 (N_32156,N_31596,N_31722);
or U32157 (N_32157,N_31616,N_31386);
nand U32158 (N_32158,N_31269,N_31620);
xnor U32159 (N_32159,N_31908,N_31248);
nor U32160 (N_32160,N_31581,N_31753);
or U32161 (N_32161,N_31209,N_31979);
and U32162 (N_32162,N_31290,N_31493);
xor U32163 (N_32163,N_31440,N_31029);
or U32164 (N_32164,N_31095,N_31665);
nand U32165 (N_32165,N_31841,N_31590);
xor U32166 (N_32166,N_31762,N_31777);
or U32167 (N_32167,N_31153,N_31989);
or U32168 (N_32168,N_31324,N_31932);
or U32169 (N_32169,N_31132,N_31573);
or U32170 (N_32170,N_31491,N_31155);
xnor U32171 (N_32171,N_31409,N_31460);
nor U32172 (N_32172,N_31724,N_31241);
and U32173 (N_32173,N_31695,N_31121);
or U32174 (N_32174,N_31282,N_31294);
and U32175 (N_32175,N_31089,N_31994);
and U32176 (N_32176,N_31166,N_31387);
and U32177 (N_32177,N_31801,N_31275);
and U32178 (N_32178,N_31279,N_31111);
or U32179 (N_32179,N_31649,N_31720);
and U32180 (N_32180,N_31977,N_31651);
nor U32181 (N_32181,N_31812,N_31502);
and U32182 (N_32182,N_31292,N_31338);
xnor U32183 (N_32183,N_31646,N_31915);
nor U32184 (N_32184,N_31514,N_31161);
xor U32185 (N_32185,N_31066,N_31505);
nand U32186 (N_32186,N_31413,N_31921);
or U32187 (N_32187,N_31662,N_31875);
nand U32188 (N_32188,N_31044,N_31565);
nor U32189 (N_32189,N_31556,N_31381);
nor U32190 (N_32190,N_31879,N_31216);
or U32191 (N_32191,N_31518,N_31984);
or U32192 (N_32192,N_31220,N_31890);
xnor U32193 (N_32193,N_31947,N_31733);
and U32194 (N_32194,N_31184,N_31422);
nand U32195 (N_32195,N_31997,N_31954);
nand U32196 (N_32196,N_31560,N_31530);
or U32197 (N_32197,N_31479,N_31696);
nor U32198 (N_32198,N_31842,N_31527);
nand U32199 (N_32199,N_31817,N_31116);
and U32200 (N_32200,N_31020,N_31850);
and U32201 (N_32201,N_31770,N_31196);
or U32202 (N_32202,N_31775,N_31210);
xnor U32203 (N_32203,N_31814,N_31679);
and U32204 (N_32204,N_31962,N_31945);
and U32205 (N_32205,N_31906,N_31688);
xnor U32206 (N_32206,N_31307,N_31016);
xor U32207 (N_32207,N_31001,N_31010);
nor U32208 (N_32208,N_31023,N_31215);
xor U32209 (N_32209,N_31676,N_31091);
and U32210 (N_32210,N_31944,N_31519);
xnor U32211 (N_32211,N_31996,N_31498);
nand U32212 (N_32212,N_31228,N_31167);
nor U32213 (N_32213,N_31607,N_31572);
or U32214 (N_32214,N_31445,N_31298);
nor U32215 (N_32215,N_31557,N_31905);
nand U32216 (N_32216,N_31786,N_31463);
nor U32217 (N_32217,N_31212,N_31871);
nand U32218 (N_32218,N_31632,N_31014);
xnor U32219 (N_32219,N_31206,N_31904);
nand U32220 (N_32220,N_31559,N_31606);
and U32221 (N_32221,N_31378,N_31289);
nand U32222 (N_32222,N_31308,N_31767);
and U32223 (N_32223,N_31471,N_31692);
nor U32224 (N_32224,N_31395,N_31992);
and U32225 (N_32225,N_31521,N_31112);
nor U32226 (N_32226,N_31589,N_31318);
nand U32227 (N_32227,N_31052,N_31003);
nor U32228 (N_32228,N_31761,N_31796);
nand U32229 (N_32229,N_31960,N_31693);
and U32230 (N_32230,N_31614,N_31656);
nor U32231 (N_32231,N_31626,N_31034);
and U32232 (N_32232,N_31863,N_31446);
nor U32233 (N_32233,N_31267,N_31694);
xnor U32234 (N_32234,N_31988,N_31147);
nor U32235 (N_32235,N_31015,N_31340);
and U32236 (N_32236,N_31919,N_31385);
nand U32237 (N_32237,N_31961,N_31012);
or U32238 (N_32238,N_31079,N_31396);
nor U32239 (N_32239,N_31080,N_31710);
or U32240 (N_32240,N_31405,N_31176);
and U32241 (N_32241,N_31585,N_31331);
nor U32242 (N_32242,N_31482,N_31213);
or U32243 (N_32243,N_31705,N_31447);
or U32244 (N_32244,N_31200,N_31730);
nor U32245 (N_32245,N_31795,N_31490);
or U32246 (N_32246,N_31974,N_31810);
or U32247 (N_32247,N_31117,N_31836);
or U32248 (N_32248,N_31907,N_31492);
xor U32249 (N_32249,N_31273,N_31827);
or U32250 (N_32250,N_31416,N_31152);
nand U32251 (N_32251,N_31284,N_31462);
or U32252 (N_32252,N_31673,N_31244);
or U32253 (N_32253,N_31726,N_31739);
xor U32254 (N_32254,N_31716,N_31102);
and U32255 (N_32255,N_31477,N_31772);
and U32256 (N_32256,N_31749,N_31107);
xor U32257 (N_32257,N_31438,N_31516);
or U32258 (N_32258,N_31547,N_31053);
xnor U32259 (N_32259,N_31846,N_31885);
xor U32260 (N_32260,N_31295,N_31380);
nor U32261 (N_32261,N_31073,N_31042);
or U32262 (N_32262,N_31319,N_31406);
nand U32263 (N_32263,N_31579,N_31055);
and U32264 (N_32264,N_31327,N_31776);
nand U32265 (N_32265,N_31140,N_31824);
xnor U32266 (N_32266,N_31837,N_31129);
xor U32267 (N_32267,N_31252,N_31854);
xnor U32268 (N_32268,N_31317,N_31171);
or U32269 (N_32269,N_31980,N_31323);
nor U32270 (N_32270,N_31718,N_31315);
or U32271 (N_32271,N_31229,N_31529);
and U32272 (N_32272,N_31369,N_31441);
nand U32273 (N_32273,N_31876,N_31881);
or U32274 (N_32274,N_31790,N_31584);
and U32275 (N_32275,N_31134,N_31636);
xnor U32276 (N_32276,N_31043,N_31891);
and U32277 (N_32277,N_31577,N_31068);
or U32278 (N_32278,N_31976,N_31262);
or U32279 (N_32279,N_31334,N_31304);
xnor U32280 (N_32280,N_31754,N_31487);
nor U32281 (N_32281,N_31464,N_31779);
or U32282 (N_32282,N_31286,N_31825);
nor U32283 (N_32283,N_31914,N_31363);
nand U32284 (N_32284,N_31735,N_31113);
xnor U32285 (N_32285,N_31063,N_31916);
and U32286 (N_32286,N_31999,N_31087);
nand U32287 (N_32287,N_31588,N_31857);
or U32288 (N_32288,N_31698,N_31105);
nand U32289 (N_32289,N_31613,N_31371);
or U32290 (N_32290,N_31028,N_31524);
nor U32291 (N_32291,N_31811,N_31541);
xor U32292 (N_32292,N_31938,N_31674);
nand U32293 (N_32293,N_31642,N_31612);
nor U32294 (N_32294,N_31118,N_31401);
nand U32295 (N_32295,N_31449,N_31439);
and U32296 (N_32296,N_31347,N_31721);
or U32297 (N_32297,N_31059,N_31928);
xor U32298 (N_32298,N_31064,N_31333);
and U32299 (N_32299,N_31356,N_31417);
nand U32300 (N_32300,N_31336,N_31913);
or U32301 (N_32301,N_31680,N_31765);
nand U32302 (N_32302,N_31344,N_31335);
nor U32303 (N_32303,N_31746,N_31054);
nand U32304 (N_32304,N_31683,N_31158);
and U32305 (N_32305,N_31266,N_31199);
and U32306 (N_32306,N_31729,N_31431);
xnor U32307 (N_32307,N_31548,N_31217);
nand U32308 (N_32308,N_31484,N_31045);
nor U32309 (N_32309,N_31608,N_31026);
or U32310 (N_32310,N_31549,N_31978);
and U32311 (N_32311,N_31122,N_31100);
xnor U32312 (N_32312,N_31250,N_31485);
and U32313 (N_32313,N_31510,N_31719);
xor U32314 (N_32314,N_31672,N_31027);
nand U32315 (N_32315,N_31964,N_31018);
nand U32316 (N_32316,N_31515,N_31630);
or U32317 (N_32317,N_31156,N_31236);
nand U32318 (N_32318,N_31917,N_31787);
nor U32319 (N_32319,N_31086,N_31476);
nand U32320 (N_32320,N_31106,N_31643);
nor U32321 (N_32321,N_31828,N_31060);
nand U32322 (N_32322,N_31009,N_31670);
nand U32323 (N_32323,N_31101,N_31377);
or U32324 (N_32324,N_31734,N_31806);
xor U32325 (N_32325,N_31580,N_31231);
xor U32326 (N_32326,N_31367,N_31888);
xor U32327 (N_32327,N_31911,N_31866);
or U32328 (N_32328,N_31935,N_31725);
nor U32329 (N_32329,N_31077,N_31070);
nor U32330 (N_32330,N_31108,N_31899);
xor U32331 (N_32331,N_31486,N_31110);
and U32332 (N_32332,N_31552,N_31697);
and U32333 (N_32333,N_31368,N_31750);
nor U32334 (N_32334,N_31708,N_31017);
nand U32335 (N_32335,N_31785,N_31169);
or U32336 (N_32336,N_31094,N_31821);
nor U32337 (N_32337,N_31640,N_31848);
or U32338 (N_32338,N_31272,N_31067);
nand U32339 (N_32339,N_31436,N_31802);
and U32340 (N_32340,N_31813,N_31430);
and U32341 (N_32341,N_31661,N_31647);
or U32342 (N_32342,N_31532,N_31578);
xnor U32343 (N_32343,N_31376,N_31467);
nand U32344 (N_32344,N_31918,N_31443);
xor U32345 (N_32345,N_31038,N_31384);
nand U32346 (N_32346,N_31967,N_31008);
or U32347 (N_32347,N_31138,N_31987);
nor U32348 (N_32348,N_31551,N_31078);
nand U32349 (N_32349,N_31973,N_31247);
nor U32350 (N_32350,N_31040,N_31995);
xnor U32351 (N_32351,N_31421,N_31312);
xor U32352 (N_32352,N_31309,N_31872);
xor U32353 (N_32353,N_31280,N_31641);
and U32354 (N_32354,N_31627,N_31226);
or U32355 (N_32355,N_31203,N_31104);
or U32356 (N_32356,N_31702,N_31170);
nor U32357 (N_32357,N_31835,N_31208);
or U32358 (N_32358,N_31459,N_31407);
nand U32359 (N_32359,N_31740,N_31263);
nand U32360 (N_32360,N_31178,N_31659);
and U32361 (N_32361,N_31883,N_31555);
xor U32362 (N_32362,N_31225,N_31260);
and U32363 (N_32363,N_31706,N_31760);
or U32364 (N_32364,N_31283,N_31154);
or U32365 (N_32365,N_31314,N_31847);
nor U32366 (N_32366,N_31867,N_31198);
nor U32367 (N_32367,N_31663,N_31258);
nand U32368 (N_32368,N_31096,N_31671);
and U32369 (N_32369,N_31736,N_31709);
xnor U32370 (N_32370,N_31330,N_31432);
nand U32371 (N_32371,N_31393,N_31359);
xnor U32372 (N_32372,N_31145,N_31357);
nand U32373 (N_32373,N_31011,N_31926);
nor U32374 (N_32374,N_31574,N_31240);
xnor U32375 (N_32375,N_31427,N_31383);
nand U32376 (N_32376,N_31041,N_31033);
and U32377 (N_32377,N_31797,N_31600);
xor U32378 (N_32378,N_31139,N_31985);
xnor U32379 (N_32379,N_31257,N_31473);
nand U32380 (N_32380,N_31398,N_31832);
or U32381 (N_32381,N_31712,N_31420);
or U32382 (N_32382,N_31700,N_31865);
nor U32383 (N_32383,N_31522,N_31504);
or U32384 (N_32384,N_31512,N_31562);
and U32385 (N_32385,N_31188,N_31894);
nand U32386 (N_32386,N_31047,N_31923);
xor U32387 (N_32387,N_31781,N_31455);
or U32388 (N_32388,N_31299,N_31638);
nor U32389 (N_32389,N_31301,N_31593);
nor U32390 (N_32390,N_31855,N_31752);
nand U32391 (N_32391,N_31925,N_31654);
xnor U32392 (N_32392,N_31860,N_31946);
or U32393 (N_32393,N_31326,N_31185);
and U32394 (N_32394,N_31550,N_31466);
nor U32395 (N_32395,N_31397,N_31076);
and U32396 (N_32396,N_31183,N_31403);
and U32397 (N_32397,N_31501,N_31766);
or U32398 (N_32398,N_31019,N_31536);
xor U32399 (N_32399,N_31611,N_31468);
and U32400 (N_32400,N_31499,N_31877);
or U32401 (N_32401,N_31822,N_31177);
xnor U32402 (N_32402,N_31525,N_31150);
nor U32403 (N_32403,N_31667,N_31022);
xnor U32404 (N_32404,N_31618,N_31937);
nor U32405 (N_32405,N_31699,N_31115);
or U32406 (N_32406,N_31534,N_31803);
and U32407 (N_32407,N_31311,N_31543);
nor U32408 (N_32408,N_31544,N_31322);
or U32409 (N_32409,N_31864,N_31348);
xor U32410 (N_32410,N_31929,N_31782);
and U32411 (N_32411,N_31930,N_31744);
nor U32412 (N_32412,N_31553,N_31255);
nand U32413 (N_32413,N_31061,N_31623);
nor U32414 (N_32414,N_31727,N_31909);
xor U32415 (N_32415,N_31222,N_31900);
nand U32416 (N_32416,N_31901,N_31249);
and U32417 (N_32417,N_31448,N_31508);
or U32418 (N_32418,N_31394,N_31972);
nand U32419 (N_32419,N_31963,N_31561);
nor U32420 (N_32420,N_31849,N_31352);
nor U32421 (N_32421,N_31949,N_31759);
xor U32422 (N_32422,N_31239,N_31715);
nor U32423 (N_32423,N_31025,N_31373);
nand U32424 (N_32424,N_31165,N_31595);
or U32425 (N_32425,N_31769,N_31296);
and U32426 (N_32426,N_31435,N_31337);
nand U32427 (N_32427,N_31669,N_31975);
nand U32428 (N_32428,N_31531,N_31940);
and U32429 (N_32429,N_31998,N_31743);
and U32430 (N_32430,N_31540,N_31265);
xnor U32431 (N_32431,N_31951,N_31653);
nor U32432 (N_32432,N_31362,N_31412);
nand U32433 (N_32433,N_31625,N_31270);
and U32434 (N_32434,N_31528,N_31682);
xnor U32435 (N_32435,N_31366,N_31732);
and U32436 (N_32436,N_31048,N_31259);
and U32437 (N_32437,N_31993,N_31223);
or U32438 (N_32438,N_31285,N_31186);
xnor U32439 (N_32439,N_31583,N_31142);
or U32440 (N_32440,N_31005,N_31090);
or U32441 (N_32441,N_31218,N_31738);
xor U32442 (N_32442,N_31582,N_31950);
nand U32443 (N_32443,N_31035,N_31820);
nor U32444 (N_32444,N_31057,N_31454);
nor U32445 (N_32445,N_31861,N_31126);
nor U32446 (N_32446,N_31024,N_31764);
or U32447 (N_32447,N_31088,N_31714);
and U32448 (N_32448,N_31633,N_31343);
nor U32449 (N_32449,N_31271,N_31192);
xor U32450 (N_32450,N_31520,N_31379);
nor U32451 (N_32451,N_31408,N_31791);
xnor U32452 (N_32452,N_31788,N_31892);
nor U32453 (N_32453,N_31037,N_31276);
and U32454 (N_32454,N_31325,N_31365);
xnor U32455 (N_32455,N_31214,N_31839);
or U32456 (N_32456,N_31202,N_31617);
or U32457 (N_32457,N_31182,N_31287);
nor U32458 (N_32458,N_31568,N_31130);
or U32459 (N_32459,N_31942,N_31187);
or U32460 (N_32460,N_31675,N_31569);
nor U32461 (N_32461,N_31360,N_31148);
nor U32462 (N_32462,N_31602,N_31751);
and U32463 (N_32463,N_31494,N_31062);
nor U32464 (N_32464,N_31388,N_31469);
nor U32465 (N_32465,N_31400,N_31723);
xor U32466 (N_32466,N_31970,N_31350);
nand U32467 (N_32467,N_31434,N_31507);
nand U32468 (N_32468,N_31878,N_31456);
and U32469 (N_32469,N_31567,N_31278);
xnor U32470 (N_32470,N_31310,N_31586);
xor U32471 (N_32471,N_31818,N_31119);
nor U32472 (N_32472,N_31444,N_31794);
xnor U32473 (N_32473,N_31261,N_31545);
and U32474 (N_32474,N_31990,N_31135);
xnor U32475 (N_32475,N_31804,N_31910);
and U32476 (N_32476,N_31332,N_31758);
or U32477 (N_32477,N_31778,N_31952);
nand U32478 (N_32478,N_31615,N_31242);
nand U32479 (N_32479,N_31542,N_31084);
nor U32480 (N_32480,N_31546,N_31741);
nor U32481 (N_32481,N_31898,N_31774);
nor U32482 (N_32482,N_31966,N_31351);
nand U32483 (N_32483,N_31472,N_31635);
or U32484 (N_32484,N_31668,N_31234);
nand U32485 (N_32485,N_31959,N_31681);
nor U32486 (N_32486,N_31621,N_31495);
xor U32487 (N_32487,N_31442,N_31819);
or U32488 (N_32488,N_31227,N_31874);
xor U32489 (N_32489,N_31943,N_31404);
or U32490 (N_32490,N_31137,N_31083);
xnor U32491 (N_32491,N_31103,N_31238);
xnor U32492 (N_32492,N_31685,N_31465);
and U32493 (N_32493,N_31889,N_31509);
nand U32494 (N_32494,N_31237,N_31004);
nor U32495 (N_32495,N_31927,N_31539);
and U32496 (N_32496,N_31564,N_31036);
and U32497 (N_32497,N_31193,N_31157);
nor U32498 (N_32498,N_31798,N_31873);
xnor U32499 (N_32499,N_31639,N_31374);
nand U32500 (N_32500,N_31738,N_31938);
nand U32501 (N_32501,N_31277,N_31274);
or U32502 (N_32502,N_31191,N_31587);
and U32503 (N_32503,N_31893,N_31714);
or U32504 (N_32504,N_31631,N_31177);
and U32505 (N_32505,N_31575,N_31625);
or U32506 (N_32506,N_31140,N_31745);
and U32507 (N_32507,N_31234,N_31333);
and U32508 (N_32508,N_31619,N_31464);
xor U32509 (N_32509,N_31921,N_31915);
and U32510 (N_32510,N_31767,N_31470);
nand U32511 (N_32511,N_31694,N_31340);
xor U32512 (N_32512,N_31993,N_31091);
xnor U32513 (N_32513,N_31163,N_31737);
and U32514 (N_32514,N_31955,N_31212);
or U32515 (N_32515,N_31048,N_31555);
xnor U32516 (N_32516,N_31380,N_31837);
xnor U32517 (N_32517,N_31125,N_31183);
nor U32518 (N_32518,N_31908,N_31389);
xnor U32519 (N_32519,N_31714,N_31668);
nand U32520 (N_32520,N_31347,N_31370);
xor U32521 (N_32521,N_31076,N_31562);
nand U32522 (N_32522,N_31732,N_31836);
xor U32523 (N_32523,N_31146,N_31003);
or U32524 (N_32524,N_31939,N_31418);
and U32525 (N_32525,N_31941,N_31713);
nand U32526 (N_32526,N_31606,N_31399);
nand U32527 (N_32527,N_31563,N_31608);
xor U32528 (N_32528,N_31538,N_31084);
nand U32529 (N_32529,N_31280,N_31980);
nand U32530 (N_32530,N_31254,N_31920);
xnor U32531 (N_32531,N_31852,N_31417);
and U32532 (N_32532,N_31934,N_31770);
or U32533 (N_32533,N_31743,N_31828);
xor U32534 (N_32534,N_31859,N_31111);
nor U32535 (N_32535,N_31702,N_31612);
and U32536 (N_32536,N_31876,N_31510);
nand U32537 (N_32537,N_31644,N_31795);
nand U32538 (N_32538,N_31302,N_31065);
nor U32539 (N_32539,N_31086,N_31340);
or U32540 (N_32540,N_31541,N_31285);
and U32541 (N_32541,N_31535,N_31754);
and U32542 (N_32542,N_31787,N_31949);
nand U32543 (N_32543,N_31075,N_31081);
nand U32544 (N_32544,N_31985,N_31308);
nand U32545 (N_32545,N_31681,N_31246);
nor U32546 (N_32546,N_31411,N_31063);
nand U32547 (N_32547,N_31963,N_31686);
or U32548 (N_32548,N_31817,N_31514);
or U32549 (N_32549,N_31016,N_31328);
and U32550 (N_32550,N_31015,N_31431);
nand U32551 (N_32551,N_31666,N_31262);
xor U32552 (N_32552,N_31273,N_31385);
or U32553 (N_32553,N_31765,N_31072);
or U32554 (N_32554,N_31146,N_31619);
nor U32555 (N_32555,N_31399,N_31488);
and U32556 (N_32556,N_31822,N_31529);
xor U32557 (N_32557,N_31625,N_31698);
nor U32558 (N_32558,N_31254,N_31573);
and U32559 (N_32559,N_31756,N_31236);
nand U32560 (N_32560,N_31477,N_31085);
or U32561 (N_32561,N_31580,N_31936);
or U32562 (N_32562,N_31784,N_31729);
nor U32563 (N_32563,N_31689,N_31604);
nor U32564 (N_32564,N_31820,N_31180);
xor U32565 (N_32565,N_31217,N_31645);
and U32566 (N_32566,N_31298,N_31215);
xor U32567 (N_32567,N_31572,N_31571);
nor U32568 (N_32568,N_31344,N_31652);
nor U32569 (N_32569,N_31715,N_31140);
xor U32570 (N_32570,N_31224,N_31063);
and U32571 (N_32571,N_31696,N_31016);
nor U32572 (N_32572,N_31453,N_31288);
nand U32573 (N_32573,N_31108,N_31517);
xnor U32574 (N_32574,N_31947,N_31688);
and U32575 (N_32575,N_31835,N_31809);
xor U32576 (N_32576,N_31800,N_31527);
nand U32577 (N_32577,N_31483,N_31974);
and U32578 (N_32578,N_31684,N_31081);
xnor U32579 (N_32579,N_31167,N_31401);
and U32580 (N_32580,N_31800,N_31395);
and U32581 (N_32581,N_31874,N_31658);
xnor U32582 (N_32582,N_31694,N_31020);
xor U32583 (N_32583,N_31800,N_31549);
and U32584 (N_32584,N_31850,N_31974);
nand U32585 (N_32585,N_31678,N_31672);
and U32586 (N_32586,N_31503,N_31037);
nor U32587 (N_32587,N_31828,N_31613);
nand U32588 (N_32588,N_31691,N_31386);
or U32589 (N_32589,N_31123,N_31718);
or U32590 (N_32590,N_31023,N_31689);
or U32591 (N_32591,N_31524,N_31801);
nand U32592 (N_32592,N_31015,N_31345);
and U32593 (N_32593,N_31975,N_31833);
and U32594 (N_32594,N_31415,N_31165);
or U32595 (N_32595,N_31615,N_31866);
nor U32596 (N_32596,N_31246,N_31513);
nand U32597 (N_32597,N_31713,N_31330);
or U32598 (N_32598,N_31731,N_31378);
xnor U32599 (N_32599,N_31342,N_31768);
and U32600 (N_32600,N_31887,N_31039);
nor U32601 (N_32601,N_31559,N_31368);
nor U32602 (N_32602,N_31021,N_31134);
nand U32603 (N_32603,N_31859,N_31309);
and U32604 (N_32604,N_31988,N_31776);
xnor U32605 (N_32605,N_31479,N_31875);
nor U32606 (N_32606,N_31366,N_31051);
xor U32607 (N_32607,N_31491,N_31659);
nand U32608 (N_32608,N_31662,N_31407);
or U32609 (N_32609,N_31638,N_31632);
nor U32610 (N_32610,N_31920,N_31890);
nor U32611 (N_32611,N_31576,N_31293);
nand U32612 (N_32612,N_31309,N_31650);
nand U32613 (N_32613,N_31893,N_31538);
nand U32614 (N_32614,N_31537,N_31737);
xnor U32615 (N_32615,N_31753,N_31548);
or U32616 (N_32616,N_31573,N_31629);
and U32617 (N_32617,N_31893,N_31380);
xor U32618 (N_32618,N_31800,N_31141);
nand U32619 (N_32619,N_31558,N_31796);
nand U32620 (N_32620,N_31652,N_31161);
nand U32621 (N_32621,N_31125,N_31561);
xnor U32622 (N_32622,N_31607,N_31325);
xnor U32623 (N_32623,N_31524,N_31332);
or U32624 (N_32624,N_31112,N_31111);
and U32625 (N_32625,N_31341,N_31849);
nand U32626 (N_32626,N_31762,N_31616);
nor U32627 (N_32627,N_31330,N_31528);
nand U32628 (N_32628,N_31124,N_31094);
or U32629 (N_32629,N_31206,N_31770);
and U32630 (N_32630,N_31577,N_31522);
or U32631 (N_32631,N_31373,N_31069);
nor U32632 (N_32632,N_31344,N_31108);
nor U32633 (N_32633,N_31092,N_31952);
xor U32634 (N_32634,N_31653,N_31985);
or U32635 (N_32635,N_31095,N_31817);
nor U32636 (N_32636,N_31626,N_31483);
xnor U32637 (N_32637,N_31463,N_31040);
nor U32638 (N_32638,N_31836,N_31083);
xor U32639 (N_32639,N_31774,N_31260);
or U32640 (N_32640,N_31343,N_31817);
nand U32641 (N_32641,N_31558,N_31023);
and U32642 (N_32642,N_31549,N_31271);
nand U32643 (N_32643,N_31143,N_31139);
and U32644 (N_32644,N_31161,N_31385);
or U32645 (N_32645,N_31358,N_31908);
nor U32646 (N_32646,N_31406,N_31258);
xor U32647 (N_32647,N_31340,N_31885);
or U32648 (N_32648,N_31208,N_31555);
or U32649 (N_32649,N_31902,N_31400);
nor U32650 (N_32650,N_31932,N_31615);
xor U32651 (N_32651,N_31504,N_31434);
xor U32652 (N_32652,N_31721,N_31846);
nand U32653 (N_32653,N_31197,N_31749);
xnor U32654 (N_32654,N_31348,N_31379);
nor U32655 (N_32655,N_31085,N_31306);
nor U32656 (N_32656,N_31611,N_31808);
nand U32657 (N_32657,N_31415,N_31562);
nor U32658 (N_32658,N_31043,N_31783);
and U32659 (N_32659,N_31318,N_31887);
nor U32660 (N_32660,N_31627,N_31362);
nor U32661 (N_32661,N_31884,N_31608);
nand U32662 (N_32662,N_31540,N_31193);
nor U32663 (N_32663,N_31309,N_31456);
or U32664 (N_32664,N_31537,N_31170);
nand U32665 (N_32665,N_31319,N_31129);
and U32666 (N_32666,N_31431,N_31126);
and U32667 (N_32667,N_31969,N_31956);
xor U32668 (N_32668,N_31354,N_31806);
nand U32669 (N_32669,N_31757,N_31329);
nand U32670 (N_32670,N_31091,N_31576);
xnor U32671 (N_32671,N_31617,N_31475);
and U32672 (N_32672,N_31255,N_31695);
and U32673 (N_32673,N_31250,N_31940);
nand U32674 (N_32674,N_31548,N_31747);
nand U32675 (N_32675,N_31170,N_31491);
nand U32676 (N_32676,N_31817,N_31691);
or U32677 (N_32677,N_31436,N_31900);
nor U32678 (N_32678,N_31764,N_31310);
and U32679 (N_32679,N_31979,N_31060);
and U32680 (N_32680,N_31047,N_31115);
xor U32681 (N_32681,N_31519,N_31432);
nor U32682 (N_32682,N_31079,N_31121);
xor U32683 (N_32683,N_31307,N_31887);
xnor U32684 (N_32684,N_31424,N_31734);
nor U32685 (N_32685,N_31834,N_31518);
xnor U32686 (N_32686,N_31109,N_31436);
nand U32687 (N_32687,N_31486,N_31374);
nand U32688 (N_32688,N_31143,N_31818);
xor U32689 (N_32689,N_31980,N_31138);
nor U32690 (N_32690,N_31145,N_31431);
and U32691 (N_32691,N_31972,N_31362);
nand U32692 (N_32692,N_31521,N_31868);
nor U32693 (N_32693,N_31364,N_31305);
and U32694 (N_32694,N_31868,N_31897);
or U32695 (N_32695,N_31611,N_31695);
nor U32696 (N_32696,N_31738,N_31844);
and U32697 (N_32697,N_31783,N_31681);
nand U32698 (N_32698,N_31249,N_31894);
xnor U32699 (N_32699,N_31176,N_31222);
xnor U32700 (N_32700,N_31386,N_31450);
nand U32701 (N_32701,N_31338,N_31176);
and U32702 (N_32702,N_31631,N_31627);
and U32703 (N_32703,N_31251,N_31554);
xor U32704 (N_32704,N_31519,N_31199);
xor U32705 (N_32705,N_31383,N_31052);
nand U32706 (N_32706,N_31022,N_31029);
nand U32707 (N_32707,N_31889,N_31103);
and U32708 (N_32708,N_31634,N_31248);
nand U32709 (N_32709,N_31137,N_31543);
and U32710 (N_32710,N_31134,N_31661);
or U32711 (N_32711,N_31846,N_31686);
nand U32712 (N_32712,N_31441,N_31951);
and U32713 (N_32713,N_31857,N_31697);
xnor U32714 (N_32714,N_31946,N_31648);
nand U32715 (N_32715,N_31948,N_31967);
xor U32716 (N_32716,N_31403,N_31478);
xor U32717 (N_32717,N_31827,N_31235);
or U32718 (N_32718,N_31370,N_31937);
xnor U32719 (N_32719,N_31521,N_31890);
nand U32720 (N_32720,N_31156,N_31430);
nor U32721 (N_32721,N_31370,N_31846);
nand U32722 (N_32722,N_31968,N_31359);
nand U32723 (N_32723,N_31636,N_31435);
nand U32724 (N_32724,N_31744,N_31497);
and U32725 (N_32725,N_31298,N_31323);
nor U32726 (N_32726,N_31081,N_31753);
nor U32727 (N_32727,N_31848,N_31675);
or U32728 (N_32728,N_31877,N_31268);
nand U32729 (N_32729,N_31909,N_31176);
xnor U32730 (N_32730,N_31643,N_31262);
and U32731 (N_32731,N_31136,N_31683);
or U32732 (N_32732,N_31743,N_31479);
and U32733 (N_32733,N_31547,N_31737);
nor U32734 (N_32734,N_31078,N_31759);
or U32735 (N_32735,N_31613,N_31549);
nand U32736 (N_32736,N_31410,N_31283);
nor U32737 (N_32737,N_31703,N_31794);
and U32738 (N_32738,N_31662,N_31588);
and U32739 (N_32739,N_31263,N_31659);
nand U32740 (N_32740,N_31513,N_31062);
nand U32741 (N_32741,N_31932,N_31115);
nor U32742 (N_32742,N_31927,N_31712);
or U32743 (N_32743,N_31135,N_31522);
or U32744 (N_32744,N_31615,N_31540);
and U32745 (N_32745,N_31655,N_31813);
xor U32746 (N_32746,N_31289,N_31421);
and U32747 (N_32747,N_31617,N_31488);
nand U32748 (N_32748,N_31980,N_31764);
nor U32749 (N_32749,N_31916,N_31811);
nand U32750 (N_32750,N_31965,N_31532);
nor U32751 (N_32751,N_31939,N_31232);
xor U32752 (N_32752,N_31000,N_31874);
xnor U32753 (N_32753,N_31920,N_31220);
nor U32754 (N_32754,N_31331,N_31102);
and U32755 (N_32755,N_31889,N_31197);
nand U32756 (N_32756,N_31473,N_31191);
and U32757 (N_32757,N_31949,N_31784);
or U32758 (N_32758,N_31508,N_31679);
nand U32759 (N_32759,N_31638,N_31754);
or U32760 (N_32760,N_31024,N_31458);
and U32761 (N_32761,N_31670,N_31808);
nand U32762 (N_32762,N_31559,N_31713);
or U32763 (N_32763,N_31194,N_31565);
xor U32764 (N_32764,N_31640,N_31533);
nand U32765 (N_32765,N_31340,N_31599);
xnor U32766 (N_32766,N_31753,N_31475);
or U32767 (N_32767,N_31133,N_31107);
and U32768 (N_32768,N_31441,N_31132);
nor U32769 (N_32769,N_31416,N_31835);
nand U32770 (N_32770,N_31641,N_31658);
or U32771 (N_32771,N_31276,N_31688);
or U32772 (N_32772,N_31062,N_31889);
or U32773 (N_32773,N_31235,N_31015);
or U32774 (N_32774,N_31277,N_31033);
xnor U32775 (N_32775,N_31655,N_31582);
and U32776 (N_32776,N_31449,N_31725);
nor U32777 (N_32777,N_31493,N_31313);
or U32778 (N_32778,N_31199,N_31935);
nor U32779 (N_32779,N_31959,N_31265);
or U32780 (N_32780,N_31807,N_31104);
xnor U32781 (N_32781,N_31376,N_31104);
nand U32782 (N_32782,N_31013,N_31621);
or U32783 (N_32783,N_31826,N_31745);
xnor U32784 (N_32784,N_31607,N_31068);
nand U32785 (N_32785,N_31686,N_31669);
and U32786 (N_32786,N_31197,N_31973);
or U32787 (N_32787,N_31059,N_31943);
xor U32788 (N_32788,N_31007,N_31608);
nand U32789 (N_32789,N_31009,N_31880);
xnor U32790 (N_32790,N_31282,N_31736);
or U32791 (N_32791,N_31231,N_31471);
or U32792 (N_32792,N_31465,N_31213);
and U32793 (N_32793,N_31611,N_31956);
nand U32794 (N_32794,N_31306,N_31474);
xnor U32795 (N_32795,N_31969,N_31801);
xor U32796 (N_32796,N_31626,N_31243);
nand U32797 (N_32797,N_31453,N_31904);
nor U32798 (N_32798,N_31267,N_31558);
nor U32799 (N_32799,N_31954,N_31379);
xnor U32800 (N_32800,N_31593,N_31801);
nand U32801 (N_32801,N_31976,N_31859);
xnor U32802 (N_32802,N_31036,N_31671);
xnor U32803 (N_32803,N_31780,N_31815);
or U32804 (N_32804,N_31773,N_31491);
nand U32805 (N_32805,N_31542,N_31623);
and U32806 (N_32806,N_31837,N_31646);
xnor U32807 (N_32807,N_31907,N_31444);
and U32808 (N_32808,N_31463,N_31860);
nand U32809 (N_32809,N_31456,N_31280);
nor U32810 (N_32810,N_31130,N_31429);
nand U32811 (N_32811,N_31426,N_31720);
or U32812 (N_32812,N_31894,N_31507);
nand U32813 (N_32813,N_31238,N_31569);
nand U32814 (N_32814,N_31606,N_31489);
or U32815 (N_32815,N_31856,N_31395);
nor U32816 (N_32816,N_31151,N_31807);
nand U32817 (N_32817,N_31080,N_31411);
xor U32818 (N_32818,N_31749,N_31134);
or U32819 (N_32819,N_31645,N_31980);
nor U32820 (N_32820,N_31516,N_31490);
xor U32821 (N_32821,N_31914,N_31067);
xor U32822 (N_32822,N_31809,N_31115);
xnor U32823 (N_32823,N_31111,N_31402);
or U32824 (N_32824,N_31018,N_31072);
xor U32825 (N_32825,N_31447,N_31829);
and U32826 (N_32826,N_31757,N_31371);
xor U32827 (N_32827,N_31530,N_31213);
or U32828 (N_32828,N_31125,N_31397);
nor U32829 (N_32829,N_31908,N_31995);
or U32830 (N_32830,N_31597,N_31598);
or U32831 (N_32831,N_31862,N_31602);
or U32832 (N_32832,N_31568,N_31613);
or U32833 (N_32833,N_31681,N_31121);
xnor U32834 (N_32834,N_31200,N_31278);
nor U32835 (N_32835,N_31556,N_31830);
and U32836 (N_32836,N_31712,N_31323);
nor U32837 (N_32837,N_31747,N_31816);
nand U32838 (N_32838,N_31195,N_31565);
nand U32839 (N_32839,N_31704,N_31519);
or U32840 (N_32840,N_31969,N_31108);
xnor U32841 (N_32841,N_31122,N_31816);
or U32842 (N_32842,N_31886,N_31232);
xnor U32843 (N_32843,N_31826,N_31799);
nand U32844 (N_32844,N_31094,N_31268);
nand U32845 (N_32845,N_31817,N_31015);
nand U32846 (N_32846,N_31507,N_31356);
nand U32847 (N_32847,N_31388,N_31373);
or U32848 (N_32848,N_31925,N_31772);
or U32849 (N_32849,N_31756,N_31430);
or U32850 (N_32850,N_31525,N_31569);
nor U32851 (N_32851,N_31665,N_31569);
or U32852 (N_32852,N_31232,N_31843);
and U32853 (N_32853,N_31808,N_31247);
nor U32854 (N_32854,N_31942,N_31337);
xor U32855 (N_32855,N_31748,N_31438);
xor U32856 (N_32856,N_31681,N_31451);
nand U32857 (N_32857,N_31738,N_31819);
nor U32858 (N_32858,N_31974,N_31053);
xnor U32859 (N_32859,N_31677,N_31464);
and U32860 (N_32860,N_31178,N_31261);
nand U32861 (N_32861,N_31558,N_31086);
nand U32862 (N_32862,N_31923,N_31019);
or U32863 (N_32863,N_31460,N_31311);
or U32864 (N_32864,N_31251,N_31169);
nor U32865 (N_32865,N_31477,N_31434);
nand U32866 (N_32866,N_31587,N_31096);
nor U32867 (N_32867,N_31063,N_31196);
nor U32868 (N_32868,N_31974,N_31014);
nand U32869 (N_32869,N_31315,N_31082);
or U32870 (N_32870,N_31487,N_31859);
nor U32871 (N_32871,N_31879,N_31457);
xnor U32872 (N_32872,N_31415,N_31262);
xnor U32873 (N_32873,N_31381,N_31132);
xnor U32874 (N_32874,N_31851,N_31719);
and U32875 (N_32875,N_31365,N_31990);
nor U32876 (N_32876,N_31085,N_31148);
xnor U32877 (N_32877,N_31257,N_31759);
xor U32878 (N_32878,N_31890,N_31700);
or U32879 (N_32879,N_31731,N_31994);
nand U32880 (N_32880,N_31982,N_31153);
nor U32881 (N_32881,N_31932,N_31255);
or U32882 (N_32882,N_31279,N_31856);
nand U32883 (N_32883,N_31126,N_31897);
xor U32884 (N_32884,N_31882,N_31279);
and U32885 (N_32885,N_31832,N_31566);
or U32886 (N_32886,N_31943,N_31808);
or U32887 (N_32887,N_31830,N_31114);
or U32888 (N_32888,N_31308,N_31651);
nand U32889 (N_32889,N_31029,N_31574);
xnor U32890 (N_32890,N_31566,N_31308);
and U32891 (N_32891,N_31374,N_31846);
nand U32892 (N_32892,N_31935,N_31657);
or U32893 (N_32893,N_31620,N_31089);
xor U32894 (N_32894,N_31727,N_31471);
xor U32895 (N_32895,N_31937,N_31604);
nor U32896 (N_32896,N_31275,N_31016);
xnor U32897 (N_32897,N_31591,N_31704);
xor U32898 (N_32898,N_31454,N_31947);
or U32899 (N_32899,N_31526,N_31562);
xnor U32900 (N_32900,N_31076,N_31868);
xor U32901 (N_32901,N_31619,N_31486);
nand U32902 (N_32902,N_31903,N_31853);
nor U32903 (N_32903,N_31803,N_31889);
or U32904 (N_32904,N_31170,N_31504);
nor U32905 (N_32905,N_31724,N_31352);
and U32906 (N_32906,N_31534,N_31994);
nor U32907 (N_32907,N_31087,N_31354);
or U32908 (N_32908,N_31330,N_31162);
and U32909 (N_32909,N_31140,N_31699);
or U32910 (N_32910,N_31690,N_31777);
nor U32911 (N_32911,N_31967,N_31864);
or U32912 (N_32912,N_31385,N_31145);
nand U32913 (N_32913,N_31411,N_31651);
nor U32914 (N_32914,N_31241,N_31398);
xor U32915 (N_32915,N_31675,N_31382);
xnor U32916 (N_32916,N_31226,N_31324);
xor U32917 (N_32917,N_31172,N_31789);
nor U32918 (N_32918,N_31274,N_31733);
xnor U32919 (N_32919,N_31493,N_31404);
xnor U32920 (N_32920,N_31342,N_31901);
xor U32921 (N_32921,N_31146,N_31541);
nand U32922 (N_32922,N_31924,N_31835);
nor U32923 (N_32923,N_31940,N_31644);
or U32924 (N_32924,N_31305,N_31559);
or U32925 (N_32925,N_31533,N_31814);
xor U32926 (N_32926,N_31418,N_31853);
or U32927 (N_32927,N_31691,N_31993);
nand U32928 (N_32928,N_31311,N_31991);
xnor U32929 (N_32929,N_31439,N_31699);
xor U32930 (N_32930,N_31675,N_31097);
nor U32931 (N_32931,N_31688,N_31824);
and U32932 (N_32932,N_31967,N_31795);
nor U32933 (N_32933,N_31566,N_31386);
nand U32934 (N_32934,N_31043,N_31787);
xnor U32935 (N_32935,N_31627,N_31415);
and U32936 (N_32936,N_31465,N_31603);
nand U32937 (N_32937,N_31112,N_31296);
nor U32938 (N_32938,N_31321,N_31250);
nand U32939 (N_32939,N_31564,N_31627);
and U32940 (N_32940,N_31221,N_31043);
nand U32941 (N_32941,N_31514,N_31419);
xor U32942 (N_32942,N_31452,N_31817);
or U32943 (N_32943,N_31520,N_31230);
or U32944 (N_32944,N_31694,N_31337);
and U32945 (N_32945,N_31431,N_31480);
and U32946 (N_32946,N_31491,N_31380);
nand U32947 (N_32947,N_31534,N_31282);
xor U32948 (N_32948,N_31641,N_31647);
xnor U32949 (N_32949,N_31363,N_31244);
or U32950 (N_32950,N_31792,N_31935);
or U32951 (N_32951,N_31342,N_31201);
nand U32952 (N_32952,N_31336,N_31618);
xor U32953 (N_32953,N_31000,N_31423);
or U32954 (N_32954,N_31986,N_31855);
nor U32955 (N_32955,N_31361,N_31711);
or U32956 (N_32956,N_31442,N_31354);
xor U32957 (N_32957,N_31532,N_31357);
nor U32958 (N_32958,N_31838,N_31129);
nor U32959 (N_32959,N_31361,N_31731);
xnor U32960 (N_32960,N_31826,N_31809);
and U32961 (N_32961,N_31611,N_31333);
nand U32962 (N_32962,N_31817,N_31773);
or U32963 (N_32963,N_31807,N_31210);
nor U32964 (N_32964,N_31004,N_31081);
nand U32965 (N_32965,N_31734,N_31649);
nor U32966 (N_32966,N_31451,N_31341);
nor U32967 (N_32967,N_31807,N_31680);
nand U32968 (N_32968,N_31998,N_31808);
nand U32969 (N_32969,N_31821,N_31506);
xnor U32970 (N_32970,N_31878,N_31655);
nand U32971 (N_32971,N_31520,N_31243);
or U32972 (N_32972,N_31624,N_31613);
nand U32973 (N_32973,N_31426,N_31185);
and U32974 (N_32974,N_31820,N_31306);
nand U32975 (N_32975,N_31014,N_31888);
and U32976 (N_32976,N_31816,N_31929);
or U32977 (N_32977,N_31722,N_31875);
nor U32978 (N_32978,N_31476,N_31972);
xnor U32979 (N_32979,N_31397,N_31310);
nand U32980 (N_32980,N_31875,N_31239);
or U32981 (N_32981,N_31357,N_31573);
nor U32982 (N_32982,N_31707,N_31705);
xor U32983 (N_32983,N_31678,N_31992);
or U32984 (N_32984,N_31208,N_31024);
nand U32985 (N_32985,N_31684,N_31762);
or U32986 (N_32986,N_31983,N_31132);
and U32987 (N_32987,N_31899,N_31042);
xnor U32988 (N_32988,N_31140,N_31495);
or U32989 (N_32989,N_31625,N_31027);
or U32990 (N_32990,N_31863,N_31882);
or U32991 (N_32991,N_31806,N_31708);
and U32992 (N_32992,N_31167,N_31264);
xnor U32993 (N_32993,N_31709,N_31328);
nor U32994 (N_32994,N_31816,N_31982);
xor U32995 (N_32995,N_31373,N_31111);
or U32996 (N_32996,N_31486,N_31926);
nor U32997 (N_32997,N_31409,N_31744);
and U32998 (N_32998,N_31228,N_31638);
and U32999 (N_32999,N_31889,N_31331);
xor U33000 (N_33000,N_32315,N_32346);
nand U33001 (N_33001,N_32010,N_32092);
or U33002 (N_33002,N_32850,N_32424);
nor U33003 (N_33003,N_32517,N_32061);
nor U33004 (N_33004,N_32725,N_32633);
nand U33005 (N_33005,N_32772,N_32863);
or U33006 (N_33006,N_32866,N_32071);
xor U33007 (N_33007,N_32780,N_32649);
xnor U33008 (N_33008,N_32371,N_32964);
and U33009 (N_33009,N_32020,N_32472);
nor U33010 (N_33010,N_32502,N_32597);
nand U33011 (N_33011,N_32841,N_32901);
nor U33012 (N_33012,N_32756,N_32192);
nor U33013 (N_33013,N_32821,N_32105);
xnor U33014 (N_33014,N_32180,N_32706);
or U33015 (N_33015,N_32859,N_32318);
nand U33016 (N_33016,N_32551,N_32735);
and U33017 (N_33017,N_32126,N_32323);
nor U33018 (N_33018,N_32816,N_32164);
xor U33019 (N_33019,N_32610,N_32256);
nand U33020 (N_33020,N_32055,N_32119);
or U33021 (N_33021,N_32096,N_32792);
nand U33022 (N_33022,N_32081,N_32334);
nor U33023 (N_33023,N_32052,N_32337);
and U33024 (N_33024,N_32263,N_32991);
or U33025 (N_33025,N_32047,N_32496);
xor U33026 (N_33026,N_32468,N_32769);
nand U33027 (N_33027,N_32778,N_32703);
and U33028 (N_33028,N_32264,N_32483);
and U33029 (N_33029,N_32045,N_32057);
and U33030 (N_33030,N_32719,N_32667);
nand U33031 (N_33031,N_32993,N_32062);
nor U33032 (N_33032,N_32390,N_32786);
xnor U33033 (N_33033,N_32986,N_32043);
and U33034 (N_33034,N_32473,N_32632);
xnor U33035 (N_33035,N_32783,N_32414);
nor U33036 (N_33036,N_32282,N_32983);
or U33037 (N_33037,N_32287,N_32560);
and U33038 (N_33038,N_32295,N_32275);
nand U33039 (N_33039,N_32104,N_32569);
and U33040 (N_33040,N_32467,N_32357);
xnor U33041 (N_33041,N_32117,N_32135);
xnor U33042 (N_33042,N_32504,N_32031);
nor U33043 (N_33043,N_32625,N_32647);
nand U33044 (N_33044,N_32013,N_32130);
nor U33045 (N_33045,N_32358,N_32524);
nand U33046 (N_33046,N_32186,N_32338);
nor U33047 (N_33047,N_32366,N_32181);
xnor U33048 (N_33048,N_32133,N_32507);
nand U33049 (N_33049,N_32865,N_32406);
or U33050 (N_33050,N_32505,N_32776);
and U33051 (N_33051,N_32845,N_32405);
xor U33052 (N_33052,N_32768,N_32539);
and U33053 (N_33053,N_32286,N_32876);
nand U33054 (N_33054,N_32101,N_32965);
and U33055 (N_33055,N_32210,N_32039);
and U33056 (N_33056,N_32306,N_32021);
nor U33057 (N_33057,N_32954,N_32987);
nand U33058 (N_33058,N_32736,N_32946);
nor U33059 (N_33059,N_32397,N_32121);
or U33060 (N_33060,N_32277,N_32134);
or U33061 (N_33061,N_32852,N_32149);
or U33062 (N_33062,N_32826,N_32738);
nor U33063 (N_33063,N_32076,N_32402);
xnor U33064 (N_33064,N_32737,N_32503);
xnor U33065 (N_33065,N_32990,N_32142);
nor U33066 (N_33066,N_32747,N_32856);
nand U33067 (N_33067,N_32743,N_32682);
or U33068 (N_33068,N_32162,N_32928);
nand U33069 (N_33069,N_32545,N_32877);
xor U33070 (N_33070,N_32403,N_32373);
nand U33071 (N_33071,N_32675,N_32871);
nor U33072 (N_33072,N_32757,N_32910);
xnor U33073 (N_33073,N_32217,N_32543);
xnor U33074 (N_33074,N_32511,N_32691);
xnor U33075 (N_33075,N_32289,N_32345);
and U33076 (N_33076,N_32308,N_32956);
and U33077 (N_33077,N_32343,N_32069);
and U33078 (N_33078,N_32512,N_32083);
nand U33079 (N_33079,N_32435,N_32755);
nor U33080 (N_33080,N_32457,N_32578);
xor U33081 (N_33081,N_32670,N_32618);
nor U33082 (N_33082,N_32479,N_32762);
xor U33083 (N_33083,N_32836,N_32589);
nor U33084 (N_33084,N_32898,N_32733);
and U33085 (N_33085,N_32448,N_32564);
and U33086 (N_33086,N_32353,N_32899);
and U33087 (N_33087,N_32949,N_32860);
or U33088 (N_33088,N_32236,N_32594);
and U33089 (N_33089,N_32331,N_32407);
and U33090 (N_33090,N_32616,N_32066);
xnor U33091 (N_33091,N_32771,N_32570);
nand U33092 (N_33092,N_32113,N_32966);
xor U33093 (N_33093,N_32720,N_32015);
and U33094 (N_33094,N_32163,N_32182);
and U33095 (N_33095,N_32660,N_32563);
nor U33096 (N_33096,N_32328,N_32196);
and U33097 (N_33097,N_32557,N_32423);
nand U33098 (N_33098,N_32639,N_32927);
and U33099 (N_33099,N_32394,N_32879);
or U33100 (N_33100,N_32829,N_32332);
nand U33101 (N_33101,N_32279,N_32515);
nor U33102 (N_33102,N_32100,N_32432);
xor U33103 (N_33103,N_32311,N_32476);
nand U33104 (N_33104,N_32443,N_32112);
nand U33105 (N_33105,N_32996,N_32360);
xor U33106 (N_33106,N_32108,N_32685);
xor U33107 (N_33107,N_32385,N_32544);
xnor U33108 (N_33108,N_32292,N_32453);
and U33109 (N_33109,N_32739,N_32035);
and U33110 (N_33110,N_32437,N_32042);
or U33111 (N_33111,N_32090,N_32693);
xnor U33112 (N_33112,N_32382,N_32365);
xor U33113 (N_33113,N_32349,N_32046);
and U33114 (N_33114,N_32599,N_32098);
nand U33115 (N_33115,N_32583,N_32540);
xor U33116 (N_33116,N_32077,N_32086);
nor U33117 (N_33117,N_32754,N_32802);
nand U33118 (N_33118,N_32652,N_32980);
or U33119 (N_33119,N_32729,N_32781);
nor U33120 (N_33120,N_32225,N_32984);
xor U33121 (N_33121,N_32731,N_32644);
nor U33122 (N_33122,N_32344,N_32678);
nand U33123 (N_33123,N_32692,N_32333);
xnor U33124 (N_33124,N_32622,N_32867);
nand U33125 (N_33125,N_32410,N_32974);
xnor U33126 (N_33126,N_32489,N_32601);
nand U33127 (N_33127,N_32482,N_32005);
and U33128 (N_33128,N_32316,N_32145);
nor U33129 (N_33129,N_32619,N_32269);
nor U33130 (N_33130,N_32326,N_32232);
or U33131 (N_33131,N_32520,N_32658);
or U33132 (N_33132,N_32070,N_32324);
xor U33133 (N_33133,N_32129,N_32226);
and U33134 (N_33134,N_32266,N_32408);
nor U33135 (N_33135,N_32469,N_32183);
xor U33136 (N_33136,N_32235,N_32559);
nor U33137 (N_33137,N_32151,N_32789);
and U33138 (N_33138,N_32033,N_32078);
xnor U33139 (N_33139,N_32029,N_32642);
and U33140 (N_33140,N_32761,N_32419);
nor U33141 (N_33141,N_32440,N_32607);
or U33142 (N_33142,N_32227,N_32645);
and U33143 (N_33143,N_32700,N_32218);
or U33144 (N_33144,N_32770,N_32716);
xnor U33145 (N_33145,N_32925,N_32817);
and U33146 (N_33146,N_32612,N_32808);
or U33147 (N_33147,N_32962,N_32679);
xor U33148 (N_33148,N_32726,N_32935);
xnor U33149 (N_33149,N_32748,N_32937);
nand U33150 (N_33150,N_32857,N_32024);
nor U33151 (N_33151,N_32442,N_32629);
nand U33152 (N_33152,N_32456,N_32596);
or U33153 (N_33153,N_32466,N_32364);
xnor U33154 (N_33154,N_32111,N_32915);
xor U33155 (N_33155,N_32027,N_32454);
nand U33156 (N_33156,N_32339,N_32734);
nand U33157 (N_33157,N_32474,N_32751);
and U33158 (N_33158,N_32006,N_32438);
xor U33159 (N_33159,N_32088,N_32140);
or U33160 (N_33160,N_32291,N_32294);
nor U33161 (N_33161,N_32582,N_32961);
xnor U33162 (N_33162,N_32745,N_32830);
or U33163 (N_33163,N_32942,N_32815);
or U33164 (N_33164,N_32458,N_32461);
nand U33165 (N_33165,N_32952,N_32073);
nor U33166 (N_33166,N_32978,N_32257);
nor U33167 (N_33167,N_32951,N_32272);
nand U33168 (N_33168,N_32004,N_32686);
xor U33169 (N_33169,N_32621,N_32262);
nor U33170 (N_33170,N_32905,N_32753);
nor U33171 (N_33171,N_32605,N_32941);
nand U33172 (N_33172,N_32203,N_32902);
and U33173 (N_33173,N_32797,N_32016);
and U33174 (N_33174,N_32565,N_32944);
xnor U33175 (N_33175,N_32573,N_32132);
or U33176 (N_33176,N_32285,N_32506);
and U33177 (N_33177,N_32766,N_32298);
nor U33178 (N_33178,N_32653,N_32034);
and U33179 (N_33179,N_32842,N_32820);
nor U33180 (N_33180,N_32425,N_32303);
nor U33181 (N_33181,N_32814,N_32635);
nor U33182 (N_33182,N_32518,N_32477);
nand U33183 (N_33183,N_32431,N_32854);
or U33184 (N_33184,N_32415,N_32873);
nor U33185 (N_33185,N_32525,N_32819);
xnor U33186 (N_33186,N_32422,N_32411);
xnor U33187 (N_33187,N_32413,N_32148);
xor U33188 (N_33188,N_32418,N_32932);
nand U33189 (N_33189,N_32259,N_32439);
and U33190 (N_33190,N_32463,N_32680);
xnor U33191 (N_33191,N_32288,N_32153);
nand U33192 (N_33192,N_32392,N_32002);
xnor U33193 (N_33193,N_32886,N_32586);
and U33194 (N_33194,N_32498,N_32810);
nand U33195 (N_33195,N_32038,N_32891);
or U33196 (N_33196,N_32401,N_32136);
or U33197 (N_33197,N_32009,N_32556);
and U33198 (N_33198,N_32904,N_32106);
nand U33199 (N_33199,N_32643,N_32727);
xnor U33200 (N_33200,N_32094,N_32212);
nand U33201 (N_33201,N_32903,N_32330);
xnor U33202 (N_33202,N_32892,N_32150);
nor U33203 (N_33203,N_32141,N_32156);
xnor U33204 (N_33204,N_32249,N_32386);
or U33205 (N_33205,N_32319,N_32896);
nor U33206 (N_33206,N_32278,N_32837);
xnor U33207 (N_33207,N_32208,N_32933);
xnor U33208 (N_33208,N_32805,N_32659);
nor U33209 (N_33209,N_32958,N_32585);
nand U33210 (N_33210,N_32994,N_32875);
xnor U33211 (N_33211,N_32803,N_32624);
nand U33212 (N_33212,N_32206,N_32939);
nor U33213 (N_33213,N_32157,N_32229);
and U33214 (N_33214,N_32451,N_32801);
xnor U33215 (N_33215,N_32603,N_32509);
and U33216 (N_33216,N_32889,N_32674);
or U33217 (N_33217,N_32920,N_32809);
or U33218 (N_33218,N_32341,N_32237);
and U33219 (N_33219,N_32926,N_32017);
nand U33220 (N_33220,N_32452,N_32895);
nand U33221 (N_33221,N_32243,N_32960);
or U33222 (N_33222,N_32715,N_32963);
or U33223 (N_33223,N_32239,N_32982);
and U33224 (N_33224,N_32554,N_32989);
nand U33225 (N_33225,N_32530,N_32590);
or U33226 (N_33226,N_32097,N_32600);
nor U33227 (N_33227,N_32059,N_32305);
or U33228 (N_33228,N_32433,N_32051);
nand U33229 (N_33229,N_32434,N_32048);
xor U33230 (N_33230,N_32626,N_32205);
and U33231 (N_33231,N_32553,N_32999);
or U33232 (N_33232,N_32872,N_32628);
nor U33233 (N_33233,N_32416,N_32722);
and U33234 (N_33234,N_32103,N_32193);
and U33235 (N_33235,N_32350,N_32465);
xnor U33236 (N_33236,N_32934,N_32484);
nand U33237 (N_33237,N_32270,N_32317);
nand U33238 (N_33238,N_32807,N_32724);
xnor U33239 (N_33239,N_32267,N_32445);
xnor U33240 (N_33240,N_32798,N_32231);
or U33241 (N_33241,N_32765,N_32152);
or U33242 (N_33242,N_32250,N_32172);
and U33243 (N_33243,N_32742,N_32701);
xnor U33244 (N_33244,N_32255,N_32537);
and U33245 (N_33245,N_32710,N_32704);
and U33246 (N_33246,N_32032,N_32767);
nor U33247 (N_33247,N_32302,N_32475);
or U33248 (N_33248,N_32219,N_32110);
and U33249 (N_33249,N_32421,N_32462);
or U33250 (N_33250,N_32646,N_32900);
or U33251 (N_33251,N_32116,N_32713);
nor U33252 (N_33252,N_32201,N_32884);
xnor U33253 (N_33253,N_32124,N_32361);
or U33254 (N_33254,N_32216,N_32493);
nor U33255 (N_33255,N_32500,N_32080);
nor U33256 (N_33256,N_32222,N_32948);
nand U33257 (N_33257,N_32579,N_32791);
or U33258 (N_33258,N_32587,N_32001);
nor U33259 (N_33259,N_32398,N_32519);
xor U33260 (N_33260,N_32492,N_32995);
or U33261 (N_33261,N_32521,N_32914);
or U33262 (N_33262,N_32146,N_32623);
nand U33263 (N_33263,N_32668,N_32179);
or U33264 (N_33264,N_32168,N_32120);
nor U33265 (N_33265,N_32940,N_32712);
or U33266 (N_33266,N_32717,N_32936);
and U33267 (N_33267,N_32014,N_32155);
nand U33268 (N_33268,N_32296,N_32887);
nor U33269 (N_33269,N_32567,N_32060);
xnor U33270 (N_33270,N_32568,N_32207);
or U33271 (N_33271,N_32728,N_32271);
nor U33272 (N_33272,N_32662,N_32855);
nor U33273 (N_33273,N_32075,N_32387);
nand U33274 (N_33274,N_32947,N_32347);
xor U33275 (N_33275,N_32118,N_32878);
xor U33276 (N_33276,N_32671,N_32019);
or U33277 (N_33277,N_32165,N_32516);
xor U33278 (N_33278,N_32127,N_32026);
xor U33279 (N_33279,N_32718,N_32188);
nand U33280 (N_33280,N_32037,N_32615);
xor U33281 (N_33281,N_32955,N_32064);
nor U33282 (N_33282,N_32528,N_32917);
nor U33283 (N_33283,N_32109,N_32195);
or U33284 (N_33284,N_32436,N_32806);
xnor U33285 (N_33285,N_32592,N_32732);
nand U33286 (N_33286,N_32684,N_32664);
xor U33287 (N_33287,N_32312,N_32834);
xnor U33288 (N_33288,N_32846,N_32730);
xnor U33289 (N_33289,N_32550,N_32694);
xor U33290 (N_33290,N_32079,N_32897);
and U33291 (N_33291,N_32487,N_32787);
nand U33292 (N_33292,N_32923,N_32758);
or U33293 (N_33293,N_32908,N_32087);
xor U33294 (N_33294,N_32028,N_32495);
xnor U33295 (N_33295,N_32510,N_32139);
and U33296 (N_33296,N_32058,N_32273);
nand U33297 (N_33297,N_32023,N_32552);
or U33298 (N_33298,N_32352,N_32374);
nand U33299 (N_33299,N_32907,N_32336);
nor U33300 (N_33300,N_32672,N_32838);
or U33301 (N_33301,N_32340,N_32547);
nand U33302 (N_33302,N_32888,N_32818);
or U33303 (N_33303,N_32348,N_32699);
or U33304 (N_33304,N_32655,N_32242);
nand U33305 (N_33305,N_32380,N_32584);
or U33306 (N_33306,N_32189,N_32301);
nor U33307 (N_33307,N_32300,N_32396);
and U33308 (N_33308,N_32174,N_32158);
nand U33309 (N_33309,N_32535,N_32566);
nand U33310 (N_33310,N_32696,N_32840);
xor U33311 (N_33311,N_32575,N_32541);
nand U33312 (N_33312,N_32906,N_32741);
or U33313 (N_33313,N_32084,N_32823);
or U33314 (N_33314,N_32882,N_32973);
nand U33315 (N_33315,N_32214,N_32630);
nand U33316 (N_33316,N_32847,N_32501);
or U33317 (N_33317,N_32919,N_32945);
or U33318 (N_33318,N_32874,N_32839);
xor U33319 (N_33319,N_32998,N_32131);
or U33320 (N_33320,N_32844,N_32428);
xnor U33321 (N_33321,N_32523,N_32608);
nand U33322 (N_33322,N_32447,N_32215);
and U33323 (N_33323,N_32170,N_32025);
nor U33324 (N_33324,N_32246,N_32714);
nand U33325 (N_33325,N_32471,N_32253);
nand U33326 (N_33326,N_32393,N_32977);
and U33327 (N_33327,N_32202,N_32053);
xor U33328 (N_33328,N_32399,N_32943);
or U33329 (N_33329,N_32363,N_32602);
nor U33330 (N_33330,N_32063,N_32641);
nor U33331 (N_33331,N_32320,N_32782);
and U33332 (N_33332,N_32233,N_32008);
xnor U33333 (N_33333,N_32763,N_32325);
or U33334 (N_33334,N_32067,N_32938);
xnor U33335 (N_33335,N_32224,N_32161);
and U33336 (N_33336,N_32388,N_32527);
nor U33337 (N_33337,N_32369,N_32293);
and U33338 (N_33338,N_32593,N_32309);
and U33339 (N_33339,N_32784,N_32281);
and U33340 (N_33340,N_32444,N_32409);
or U33341 (N_33341,N_32211,N_32811);
and U33342 (N_33342,N_32307,N_32687);
and U33343 (N_33343,N_32238,N_32957);
nand U33344 (N_33344,N_32634,N_32377);
or U33345 (N_33345,N_32683,N_32221);
xnor U33346 (N_33346,N_32513,N_32744);
nand U33347 (N_33347,N_32843,N_32265);
nor U33348 (N_33348,N_32427,N_32122);
and U33349 (N_33349,N_32752,N_32209);
or U33350 (N_33350,N_32853,N_32804);
nand U33351 (N_33351,N_32909,N_32831);
xor U33352 (N_33352,N_32160,N_32572);
nor U33353 (N_33353,N_32372,N_32676);
and U33354 (N_33354,N_32997,N_32656);
xnor U33355 (N_33355,N_32178,N_32950);
nand U33356 (N_33356,N_32381,N_32972);
or U33357 (N_33357,N_32379,N_32795);
nor U33358 (N_33358,N_32190,N_32197);
nand U33359 (N_33359,N_32412,N_32979);
nand U33360 (N_33360,N_32611,N_32204);
xnor U33361 (N_33361,N_32709,N_32669);
xnor U33362 (N_33362,N_32123,N_32184);
nor U33363 (N_33363,N_32627,N_32894);
or U33364 (N_33364,N_32470,N_32522);
xor U33365 (N_33365,N_32562,N_32681);
nor U33366 (N_33366,N_32598,N_32749);
xor U33367 (N_33367,N_32574,N_32147);
xor U33368 (N_33368,N_32533,N_32144);
nand U33369 (N_33369,N_32446,N_32708);
xor U33370 (N_33370,N_32449,N_32661);
or U33371 (N_33371,N_32370,N_32992);
or U33372 (N_33372,N_32880,N_32918);
nand U33373 (N_33373,N_32138,N_32159);
nand U33374 (N_33374,N_32812,N_32125);
or U33375 (N_33375,N_32491,N_32790);
nand U33376 (N_33376,N_32698,N_32665);
xnor U33377 (N_33377,N_32775,N_32234);
or U33378 (N_33378,N_32800,N_32930);
nand U33379 (N_33379,N_32760,N_32280);
or U33380 (N_33380,N_32555,N_32970);
or U33381 (N_33381,N_32050,N_32114);
or U33382 (N_33382,N_32796,N_32012);
or U33383 (N_33383,N_32480,N_32198);
or U33384 (N_33384,N_32604,N_32975);
and U33385 (N_33385,N_32581,N_32774);
nor U33386 (N_33386,N_32391,N_32988);
or U33387 (N_33387,N_32187,N_32514);
nor U33388 (N_33388,N_32534,N_32143);
and U33389 (N_33389,N_32441,N_32430);
nand U33390 (N_33390,N_32030,N_32091);
nor U33391 (N_33391,N_32223,N_32931);
or U33392 (N_33392,N_32723,N_32200);
nand U33393 (N_33393,N_32885,N_32044);
nor U33394 (N_33394,N_32356,N_32404);
nand U33395 (N_33395,N_32881,N_32526);
or U33396 (N_33396,N_32228,N_32959);
xor U33397 (N_33397,N_32327,N_32759);
or U33398 (N_33398,N_32137,N_32711);
and U33399 (N_33399,N_32191,N_32536);
and U33400 (N_33400,N_32690,N_32799);
nor U33401 (N_33401,N_32702,N_32697);
xnor U33402 (N_33402,N_32813,N_32663);
or U33403 (N_33403,N_32673,N_32304);
xnor U33404 (N_33404,N_32869,N_32777);
nand U33405 (N_33405,N_32929,N_32689);
nand U33406 (N_33406,N_32283,N_32529);
xor U33407 (N_33407,N_32638,N_32011);
nand U33408 (N_33408,N_32240,N_32072);
or U33409 (N_33409,N_32464,N_32588);
nand U33410 (N_33410,N_32089,N_32383);
and U33411 (N_33411,N_32746,N_32354);
and U33412 (N_33412,N_32082,N_32499);
xnor U33413 (N_33413,N_32538,N_32613);
or U33414 (N_33414,N_32252,N_32362);
nor U33415 (N_33415,N_32128,N_32054);
xor U33416 (N_33416,N_32740,N_32115);
nor U33417 (N_33417,N_32321,N_32166);
nor U33418 (N_33418,N_32849,N_32705);
nand U33419 (N_33419,N_32185,N_32245);
xor U33420 (N_33420,N_32494,N_32022);
xnor U33421 (N_33421,N_32169,N_32640);
xor U33422 (N_33422,N_32244,N_32968);
xor U33423 (N_33423,N_32868,N_32953);
nand U33424 (N_33424,N_32794,N_32862);
xor U33425 (N_33425,N_32003,N_32355);
or U33426 (N_33426,N_32041,N_32870);
and U33427 (N_33427,N_32376,N_32851);
nor U33428 (N_33428,N_32450,N_32532);
nand U33429 (N_33429,N_32912,N_32102);
and U33430 (N_33430,N_32367,N_32558);
xnor U33431 (N_33431,N_32864,N_32368);
or U33432 (N_33432,N_32893,N_32213);
nor U33433 (N_33433,N_32651,N_32486);
nand U33434 (N_33434,N_32173,N_32107);
xnor U33435 (N_33435,N_32788,N_32695);
nor U33436 (N_33436,N_32508,N_32637);
or U33437 (N_33437,N_32176,N_32395);
nor U33438 (N_33438,N_32258,N_32576);
and U33439 (N_33439,N_32577,N_32251);
and U33440 (N_33440,N_32389,N_32636);
nand U33441 (N_33441,N_32921,N_32542);
xnor U33442 (N_33442,N_32199,N_32459);
and U33443 (N_33443,N_32548,N_32260);
xnor U33444 (N_33444,N_32848,N_32721);
or U33445 (N_33445,N_32351,N_32617);
nor U33446 (N_33446,N_32000,N_32314);
and U33447 (N_33447,N_32220,N_32420);
and U33448 (N_33448,N_32976,N_32688);
xor U33449 (N_33449,N_32764,N_32861);
nor U33450 (N_33450,N_32322,N_32247);
or U33451 (N_33451,N_32378,N_32261);
or U33452 (N_33452,N_32171,N_32631);
nor U33453 (N_33453,N_32065,N_32154);
nor U33454 (N_33454,N_32359,N_32175);
xor U33455 (N_33455,N_32549,N_32384);
and U33456 (N_33456,N_32890,N_32481);
nand U33457 (N_33457,N_32194,N_32248);
nand U33458 (N_33458,N_32614,N_32313);
or U33459 (N_33459,N_32429,N_32707);
and U33460 (N_33460,N_32981,N_32230);
or U33461 (N_33461,N_32167,N_32824);
nor U33462 (N_33462,N_32924,N_32099);
xnor U33463 (N_33463,N_32241,N_32335);
xnor U33464 (N_33464,N_32254,N_32985);
and U33465 (N_33465,N_32400,N_32056);
xor U33466 (N_33466,N_32832,N_32375);
xnor U33467 (N_33467,N_32268,N_32785);
or U33468 (N_33468,N_32883,N_32654);
xnor U33469 (N_33469,N_32561,N_32049);
and U33470 (N_33470,N_32591,N_32822);
xnor U33471 (N_33471,N_32490,N_32828);
xor U33472 (N_33472,N_32342,N_32036);
nand U33473 (N_33473,N_32297,N_32580);
nor U33474 (N_33474,N_32967,N_32773);
and U33475 (N_33475,N_32488,N_32093);
nor U33476 (N_33476,N_32284,N_32455);
xnor U33477 (N_33477,N_32276,N_32074);
nor U33478 (N_33478,N_32040,N_32007);
nand U33479 (N_33479,N_32299,N_32916);
xnor U33480 (N_33480,N_32648,N_32018);
and U33481 (N_33481,N_32095,N_32531);
nor U33482 (N_33482,N_32571,N_32650);
nand U33483 (N_33483,N_32595,N_32497);
or U33484 (N_33484,N_32620,N_32911);
nand U33485 (N_33485,N_32290,N_32825);
nand U33486 (N_33486,N_32858,N_32666);
and U33487 (N_33487,N_32478,N_32922);
and U33488 (N_33488,N_32426,N_32971);
nor U33489 (N_33489,N_32177,N_32677);
and U33490 (N_33490,N_32779,N_32606);
or U33491 (N_33491,N_32827,N_32460);
nor U33492 (N_33492,N_32068,N_32833);
or U33493 (N_33493,N_32485,N_32546);
xor U33494 (N_33494,N_32310,N_32657);
and U33495 (N_33495,N_32609,N_32274);
and U33496 (N_33496,N_32417,N_32750);
xnor U33497 (N_33497,N_32793,N_32085);
nor U33498 (N_33498,N_32835,N_32969);
nand U33499 (N_33499,N_32913,N_32329);
nand U33500 (N_33500,N_32362,N_32530);
or U33501 (N_33501,N_32981,N_32311);
and U33502 (N_33502,N_32241,N_32257);
xor U33503 (N_33503,N_32325,N_32848);
nand U33504 (N_33504,N_32605,N_32565);
and U33505 (N_33505,N_32032,N_32755);
nor U33506 (N_33506,N_32137,N_32953);
nor U33507 (N_33507,N_32556,N_32888);
and U33508 (N_33508,N_32227,N_32917);
and U33509 (N_33509,N_32995,N_32554);
nor U33510 (N_33510,N_32149,N_32605);
or U33511 (N_33511,N_32051,N_32791);
and U33512 (N_33512,N_32988,N_32132);
or U33513 (N_33513,N_32099,N_32017);
nand U33514 (N_33514,N_32873,N_32322);
or U33515 (N_33515,N_32514,N_32956);
and U33516 (N_33516,N_32430,N_32120);
and U33517 (N_33517,N_32132,N_32218);
nand U33518 (N_33518,N_32539,N_32348);
xnor U33519 (N_33519,N_32272,N_32962);
nor U33520 (N_33520,N_32348,N_32041);
nand U33521 (N_33521,N_32960,N_32755);
and U33522 (N_33522,N_32287,N_32672);
nor U33523 (N_33523,N_32758,N_32204);
or U33524 (N_33524,N_32437,N_32822);
or U33525 (N_33525,N_32632,N_32707);
and U33526 (N_33526,N_32059,N_32606);
and U33527 (N_33527,N_32738,N_32301);
or U33528 (N_33528,N_32308,N_32688);
nand U33529 (N_33529,N_32261,N_32376);
and U33530 (N_33530,N_32193,N_32537);
nand U33531 (N_33531,N_32423,N_32021);
or U33532 (N_33532,N_32436,N_32137);
nor U33533 (N_33533,N_32263,N_32291);
nand U33534 (N_33534,N_32372,N_32601);
nor U33535 (N_33535,N_32674,N_32119);
nor U33536 (N_33536,N_32701,N_32681);
or U33537 (N_33537,N_32494,N_32606);
nor U33538 (N_33538,N_32152,N_32755);
nor U33539 (N_33539,N_32133,N_32463);
and U33540 (N_33540,N_32440,N_32938);
or U33541 (N_33541,N_32296,N_32700);
and U33542 (N_33542,N_32411,N_32804);
xnor U33543 (N_33543,N_32695,N_32054);
and U33544 (N_33544,N_32480,N_32545);
nand U33545 (N_33545,N_32672,N_32191);
nand U33546 (N_33546,N_32569,N_32106);
or U33547 (N_33547,N_32683,N_32265);
and U33548 (N_33548,N_32141,N_32557);
xor U33549 (N_33549,N_32399,N_32468);
nor U33550 (N_33550,N_32691,N_32836);
xor U33551 (N_33551,N_32117,N_32440);
nor U33552 (N_33552,N_32506,N_32780);
xor U33553 (N_33553,N_32761,N_32075);
and U33554 (N_33554,N_32128,N_32885);
xor U33555 (N_33555,N_32657,N_32718);
nor U33556 (N_33556,N_32750,N_32429);
and U33557 (N_33557,N_32161,N_32394);
nor U33558 (N_33558,N_32959,N_32606);
xor U33559 (N_33559,N_32034,N_32859);
nand U33560 (N_33560,N_32824,N_32477);
xnor U33561 (N_33561,N_32135,N_32778);
xor U33562 (N_33562,N_32198,N_32942);
nand U33563 (N_33563,N_32227,N_32129);
or U33564 (N_33564,N_32606,N_32373);
nand U33565 (N_33565,N_32359,N_32031);
nand U33566 (N_33566,N_32515,N_32786);
nor U33567 (N_33567,N_32557,N_32355);
or U33568 (N_33568,N_32765,N_32463);
nor U33569 (N_33569,N_32217,N_32608);
nand U33570 (N_33570,N_32460,N_32003);
xnor U33571 (N_33571,N_32542,N_32243);
nor U33572 (N_33572,N_32148,N_32285);
nand U33573 (N_33573,N_32018,N_32843);
xnor U33574 (N_33574,N_32751,N_32974);
nand U33575 (N_33575,N_32447,N_32403);
and U33576 (N_33576,N_32601,N_32102);
nor U33577 (N_33577,N_32636,N_32588);
and U33578 (N_33578,N_32662,N_32490);
xnor U33579 (N_33579,N_32803,N_32246);
nor U33580 (N_33580,N_32905,N_32932);
and U33581 (N_33581,N_32437,N_32981);
nor U33582 (N_33582,N_32909,N_32695);
xnor U33583 (N_33583,N_32394,N_32535);
nand U33584 (N_33584,N_32165,N_32940);
and U33585 (N_33585,N_32418,N_32882);
xor U33586 (N_33586,N_32399,N_32071);
nand U33587 (N_33587,N_32608,N_32852);
nor U33588 (N_33588,N_32434,N_32252);
xor U33589 (N_33589,N_32577,N_32797);
and U33590 (N_33590,N_32722,N_32899);
or U33591 (N_33591,N_32338,N_32443);
nand U33592 (N_33592,N_32331,N_32552);
nor U33593 (N_33593,N_32838,N_32129);
or U33594 (N_33594,N_32916,N_32509);
xor U33595 (N_33595,N_32304,N_32460);
or U33596 (N_33596,N_32906,N_32666);
nand U33597 (N_33597,N_32592,N_32022);
xor U33598 (N_33598,N_32804,N_32625);
or U33599 (N_33599,N_32140,N_32783);
nor U33600 (N_33600,N_32542,N_32804);
nor U33601 (N_33601,N_32428,N_32927);
xnor U33602 (N_33602,N_32574,N_32510);
nor U33603 (N_33603,N_32234,N_32256);
or U33604 (N_33604,N_32669,N_32342);
or U33605 (N_33605,N_32795,N_32832);
nand U33606 (N_33606,N_32134,N_32326);
and U33607 (N_33607,N_32424,N_32976);
xnor U33608 (N_33608,N_32023,N_32472);
and U33609 (N_33609,N_32933,N_32221);
xor U33610 (N_33610,N_32695,N_32685);
xor U33611 (N_33611,N_32591,N_32848);
nand U33612 (N_33612,N_32507,N_32790);
xnor U33613 (N_33613,N_32859,N_32914);
nor U33614 (N_33614,N_32607,N_32599);
and U33615 (N_33615,N_32796,N_32025);
nand U33616 (N_33616,N_32309,N_32583);
xnor U33617 (N_33617,N_32500,N_32887);
and U33618 (N_33618,N_32166,N_32934);
or U33619 (N_33619,N_32910,N_32392);
nor U33620 (N_33620,N_32314,N_32579);
and U33621 (N_33621,N_32921,N_32858);
xor U33622 (N_33622,N_32616,N_32698);
or U33623 (N_33623,N_32182,N_32020);
xor U33624 (N_33624,N_32666,N_32020);
or U33625 (N_33625,N_32178,N_32349);
xor U33626 (N_33626,N_32080,N_32197);
xor U33627 (N_33627,N_32660,N_32908);
or U33628 (N_33628,N_32224,N_32164);
or U33629 (N_33629,N_32891,N_32864);
nor U33630 (N_33630,N_32280,N_32717);
xor U33631 (N_33631,N_32998,N_32707);
nor U33632 (N_33632,N_32814,N_32731);
or U33633 (N_33633,N_32604,N_32866);
or U33634 (N_33634,N_32995,N_32714);
nor U33635 (N_33635,N_32676,N_32689);
nand U33636 (N_33636,N_32702,N_32226);
nor U33637 (N_33637,N_32777,N_32178);
or U33638 (N_33638,N_32511,N_32164);
nor U33639 (N_33639,N_32070,N_32267);
nand U33640 (N_33640,N_32263,N_32404);
nand U33641 (N_33641,N_32651,N_32021);
xnor U33642 (N_33642,N_32208,N_32919);
xnor U33643 (N_33643,N_32749,N_32288);
or U33644 (N_33644,N_32420,N_32603);
nor U33645 (N_33645,N_32765,N_32950);
or U33646 (N_33646,N_32390,N_32449);
xnor U33647 (N_33647,N_32393,N_32178);
and U33648 (N_33648,N_32726,N_32234);
nor U33649 (N_33649,N_32130,N_32848);
or U33650 (N_33650,N_32073,N_32318);
nand U33651 (N_33651,N_32206,N_32038);
or U33652 (N_33652,N_32020,N_32538);
or U33653 (N_33653,N_32450,N_32232);
nand U33654 (N_33654,N_32962,N_32913);
nand U33655 (N_33655,N_32885,N_32521);
nor U33656 (N_33656,N_32594,N_32720);
or U33657 (N_33657,N_32217,N_32962);
nand U33658 (N_33658,N_32705,N_32145);
nand U33659 (N_33659,N_32312,N_32195);
and U33660 (N_33660,N_32848,N_32438);
and U33661 (N_33661,N_32793,N_32439);
nand U33662 (N_33662,N_32218,N_32576);
nor U33663 (N_33663,N_32369,N_32635);
or U33664 (N_33664,N_32816,N_32127);
nand U33665 (N_33665,N_32109,N_32651);
or U33666 (N_33666,N_32703,N_32008);
xnor U33667 (N_33667,N_32074,N_32304);
or U33668 (N_33668,N_32273,N_32700);
or U33669 (N_33669,N_32674,N_32585);
nor U33670 (N_33670,N_32346,N_32569);
nor U33671 (N_33671,N_32534,N_32606);
nor U33672 (N_33672,N_32148,N_32367);
nand U33673 (N_33673,N_32207,N_32735);
or U33674 (N_33674,N_32943,N_32976);
and U33675 (N_33675,N_32734,N_32420);
nor U33676 (N_33676,N_32492,N_32845);
nand U33677 (N_33677,N_32921,N_32401);
and U33678 (N_33678,N_32473,N_32627);
nor U33679 (N_33679,N_32529,N_32794);
xor U33680 (N_33680,N_32250,N_32940);
or U33681 (N_33681,N_32690,N_32058);
nand U33682 (N_33682,N_32791,N_32933);
nor U33683 (N_33683,N_32459,N_32210);
nand U33684 (N_33684,N_32956,N_32735);
and U33685 (N_33685,N_32218,N_32535);
xnor U33686 (N_33686,N_32457,N_32716);
xnor U33687 (N_33687,N_32434,N_32011);
and U33688 (N_33688,N_32516,N_32361);
nand U33689 (N_33689,N_32330,N_32331);
nand U33690 (N_33690,N_32106,N_32574);
and U33691 (N_33691,N_32317,N_32452);
or U33692 (N_33692,N_32375,N_32486);
nor U33693 (N_33693,N_32561,N_32805);
xnor U33694 (N_33694,N_32338,N_32453);
xor U33695 (N_33695,N_32010,N_32813);
and U33696 (N_33696,N_32976,N_32237);
xor U33697 (N_33697,N_32854,N_32299);
and U33698 (N_33698,N_32269,N_32967);
nand U33699 (N_33699,N_32521,N_32745);
nor U33700 (N_33700,N_32699,N_32106);
xor U33701 (N_33701,N_32873,N_32069);
or U33702 (N_33702,N_32752,N_32787);
and U33703 (N_33703,N_32354,N_32337);
xor U33704 (N_33704,N_32310,N_32130);
and U33705 (N_33705,N_32416,N_32205);
and U33706 (N_33706,N_32050,N_32102);
xnor U33707 (N_33707,N_32619,N_32286);
nand U33708 (N_33708,N_32835,N_32213);
or U33709 (N_33709,N_32327,N_32100);
or U33710 (N_33710,N_32688,N_32603);
or U33711 (N_33711,N_32366,N_32531);
nor U33712 (N_33712,N_32497,N_32502);
nor U33713 (N_33713,N_32916,N_32482);
or U33714 (N_33714,N_32797,N_32834);
nor U33715 (N_33715,N_32639,N_32759);
and U33716 (N_33716,N_32862,N_32470);
xor U33717 (N_33717,N_32668,N_32446);
nor U33718 (N_33718,N_32335,N_32636);
xnor U33719 (N_33719,N_32463,N_32864);
and U33720 (N_33720,N_32951,N_32841);
or U33721 (N_33721,N_32575,N_32846);
nand U33722 (N_33722,N_32594,N_32716);
xor U33723 (N_33723,N_32415,N_32225);
or U33724 (N_33724,N_32159,N_32638);
or U33725 (N_33725,N_32276,N_32585);
and U33726 (N_33726,N_32715,N_32400);
xor U33727 (N_33727,N_32998,N_32447);
nor U33728 (N_33728,N_32475,N_32385);
nand U33729 (N_33729,N_32798,N_32715);
or U33730 (N_33730,N_32626,N_32848);
or U33731 (N_33731,N_32732,N_32359);
and U33732 (N_33732,N_32757,N_32153);
or U33733 (N_33733,N_32532,N_32847);
or U33734 (N_33734,N_32460,N_32070);
nor U33735 (N_33735,N_32093,N_32803);
or U33736 (N_33736,N_32709,N_32172);
or U33737 (N_33737,N_32210,N_32717);
nand U33738 (N_33738,N_32991,N_32357);
or U33739 (N_33739,N_32414,N_32773);
or U33740 (N_33740,N_32887,N_32793);
nor U33741 (N_33741,N_32321,N_32907);
and U33742 (N_33742,N_32919,N_32361);
nor U33743 (N_33743,N_32572,N_32079);
and U33744 (N_33744,N_32485,N_32583);
nor U33745 (N_33745,N_32035,N_32852);
nand U33746 (N_33746,N_32832,N_32967);
and U33747 (N_33747,N_32111,N_32785);
nor U33748 (N_33748,N_32316,N_32433);
and U33749 (N_33749,N_32599,N_32537);
nand U33750 (N_33750,N_32061,N_32289);
nor U33751 (N_33751,N_32839,N_32493);
and U33752 (N_33752,N_32210,N_32999);
nor U33753 (N_33753,N_32203,N_32168);
nand U33754 (N_33754,N_32723,N_32482);
nor U33755 (N_33755,N_32144,N_32903);
nor U33756 (N_33756,N_32111,N_32751);
nor U33757 (N_33757,N_32778,N_32686);
and U33758 (N_33758,N_32604,N_32582);
xnor U33759 (N_33759,N_32212,N_32497);
nor U33760 (N_33760,N_32753,N_32701);
or U33761 (N_33761,N_32777,N_32012);
nand U33762 (N_33762,N_32462,N_32008);
and U33763 (N_33763,N_32957,N_32834);
xnor U33764 (N_33764,N_32919,N_32868);
xor U33765 (N_33765,N_32189,N_32203);
and U33766 (N_33766,N_32854,N_32626);
xnor U33767 (N_33767,N_32272,N_32075);
nor U33768 (N_33768,N_32706,N_32208);
xor U33769 (N_33769,N_32733,N_32585);
xor U33770 (N_33770,N_32123,N_32883);
or U33771 (N_33771,N_32245,N_32890);
nand U33772 (N_33772,N_32429,N_32499);
xor U33773 (N_33773,N_32657,N_32968);
nor U33774 (N_33774,N_32991,N_32778);
and U33775 (N_33775,N_32812,N_32153);
or U33776 (N_33776,N_32496,N_32842);
xnor U33777 (N_33777,N_32378,N_32686);
nor U33778 (N_33778,N_32858,N_32174);
and U33779 (N_33779,N_32163,N_32381);
xnor U33780 (N_33780,N_32302,N_32201);
nand U33781 (N_33781,N_32178,N_32958);
nor U33782 (N_33782,N_32745,N_32033);
nand U33783 (N_33783,N_32400,N_32059);
xor U33784 (N_33784,N_32935,N_32285);
xnor U33785 (N_33785,N_32042,N_32448);
nor U33786 (N_33786,N_32783,N_32610);
xor U33787 (N_33787,N_32156,N_32472);
and U33788 (N_33788,N_32550,N_32490);
and U33789 (N_33789,N_32316,N_32389);
nor U33790 (N_33790,N_32825,N_32103);
xor U33791 (N_33791,N_32967,N_32996);
xor U33792 (N_33792,N_32539,N_32406);
nand U33793 (N_33793,N_32771,N_32728);
nand U33794 (N_33794,N_32278,N_32336);
nor U33795 (N_33795,N_32973,N_32904);
nand U33796 (N_33796,N_32641,N_32080);
nand U33797 (N_33797,N_32470,N_32176);
nand U33798 (N_33798,N_32570,N_32341);
or U33799 (N_33799,N_32453,N_32417);
and U33800 (N_33800,N_32837,N_32856);
xnor U33801 (N_33801,N_32303,N_32122);
or U33802 (N_33802,N_32678,N_32345);
or U33803 (N_33803,N_32651,N_32139);
xnor U33804 (N_33804,N_32979,N_32638);
nand U33805 (N_33805,N_32217,N_32303);
xnor U33806 (N_33806,N_32865,N_32093);
nor U33807 (N_33807,N_32832,N_32452);
or U33808 (N_33808,N_32043,N_32231);
xnor U33809 (N_33809,N_32472,N_32439);
xnor U33810 (N_33810,N_32353,N_32846);
and U33811 (N_33811,N_32202,N_32905);
nand U33812 (N_33812,N_32487,N_32533);
and U33813 (N_33813,N_32598,N_32186);
xnor U33814 (N_33814,N_32788,N_32346);
or U33815 (N_33815,N_32134,N_32708);
or U33816 (N_33816,N_32213,N_32030);
and U33817 (N_33817,N_32054,N_32469);
and U33818 (N_33818,N_32318,N_32826);
and U33819 (N_33819,N_32659,N_32145);
and U33820 (N_33820,N_32903,N_32244);
xnor U33821 (N_33821,N_32837,N_32279);
or U33822 (N_33822,N_32891,N_32670);
and U33823 (N_33823,N_32882,N_32900);
and U33824 (N_33824,N_32463,N_32697);
nor U33825 (N_33825,N_32419,N_32238);
or U33826 (N_33826,N_32534,N_32985);
nand U33827 (N_33827,N_32694,N_32659);
xnor U33828 (N_33828,N_32919,N_32305);
nor U33829 (N_33829,N_32314,N_32021);
and U33830 (N_33830,N_32374,N_32210);
nand U33831 (N_33831,N_32644,N_32025);
nor U33832 (N_33832,N_32187,N_32131);
nor U33833 (N_33833,N_32242,N_32083);
or U33834 (N_33834,N_32841,N_32969);
xor U33835 (N_33835,N_32230,N_32636);
nand U33836 (N_33836,N_32967,N_32629);
nor U33837 (N_33837,N_32339,N_32138);
nor U33838 (N_33838,N_32340,N_32917);
xor U33839 (N_33839,N_32206,N_32836);
nor U33840 (N_33840,N_32964,N_32370);
or U33841 (N_33841,N_32391,N_32557);
and U33842 (N_33842,N_32278,N_32707);
nand U33843 (N_33843,N_32852,N_32701);
xnor U33844 (N_33844,N_32289,N_32943);
xnor U33845 (N_33845,N_32733,N_32852);
xor U33846 (N_33846,N_32638,N_32498);
nand U33847 (N_33847,N_32852,N_32097);
and U33848 (N_33848,N_32281,N_32265);
and U33849 (N_33849,N_32581,N_32248);
xor U33850 (N_33850,N_32131,N_32722);
and U33851 (N_33851,N_32585,N_32176);
and U33852 (N_33852,N_32526,N_32623);
or U33853 (N_33853,N_32774,N_32174);
nor U33854 (N_33854,N_32198,N_32363);
nand U33855 (N_33855,N_32318,N_32674);
nand U33856 (N_33856,N_32923,N_32392);
or U33857 (N_33857,N_32255,N_32942);
nand U33858 (N_33858,N_32675,N_32813);
or U33859 (N_33859,N_32766,N_32357);
and U33860 (N_33860,N_32615,N_32461);
or U33861 (N_33861,N_32405,N_32071);
nand U33862 (N_33862,N_32129,N_32802);
or U33863 (N_33863,N_32942,N_32761);
or U33864 (N_33864,N_32842,N_32430);
xnor U33865 (N_33865,N_32925,N_32684);
or U33866 (N_33866,N_32996,N_32457);
xnor U33867 (N_33867,N_32449,N_32438);
nand U33868 (N_33868,N_32761,N_32226);
or U33869 (N_33869,N_32073,N_32304);
nand U33870 (N_33870,N_32984,N_32672);
nand U33871 (N_33871,N_32117,N_32176);
xnor U33872 (N_33872,N_32197,N_32748);
nor U33873 (N_33873,N_32505,N_32946);
xnor U33874 (N_33874,N_32170,N_32265);
nor U33875 (N_33875,N_32194,N_32481);
xor U33876 (N_33876,N_32746,N_32515);
or U33877 (N_33877,N_32388,N_32220);
xor U33878 (N_33878,N_32520,N_32549);
xnor U33879 (N_33879,N_32312,N_32229);
xor U33880 (N_33880,N_32570,N_32904);
or U33881 (N_33881,N_32096,N_32440);
nor U33882 (N_33882,N_32816,N_32852);
nor U33883 (N_33883,N_32981,N_32710);
nand U33884 (N_33884,N_32074,N_32640);
and U33885 (N_33885,N_32390,N_32454);
nand U33886 (N_33886,N_32256,N_32213);
xor U33887 (N_33887,N_32416,N_32371);
or U33888 (N_33888,N_32690,N_32930);
xor U33889 (N_33889,N_32498,N_32249);
nor U33890 (N_33890,N_32481,N_32416);
nor U33891 (N_33891,N_32244,N_32485);
nand U33892 (N_33892,N_32087,N_32246);
nor U33893 (N_33893,N_32232,N_32349);
nand U33894 (N_33894,N_32999,N_32026);
and U33895 (N_33895,N_32946,N_32973);
nor U33896 (N_33896,N_32941,N_32507);
or U33897 (N_33897,N_32195,N_32325);
nor U33898 (N_33898,N_32537,N_32928);
or U33899 (N_33899,N_32409,N_32965);
or U33900 (N_33900,N_32135,N_32457);
nor U33901 (N_33901,N_32234,N_32891);
xnor U33902 (N_33902,N_32162,N_32479);
nand U33903 (N_33903,N_32581,N_32116);
and U33904 (N_33904,N_32148,N_32156);
nand U33905 (N_33905,N_32920,N_32394);
xor U33906 (N_33906,N_32842,N_32473);
or U33907 (N_33907,N_32935,N_32808);
nand U33908 (N_33908,N_32477,N_32621);
or U33909 (N_33909,N_32953,N_32500);
or U33910 (N_33910,N_32543,N_32552);
xnor U33911 (N_33911,N_32826,N_32301);
nor U33912 (N_33912,N_32058,N_32972);
and U33913 (N_33913,N_32639,N_32853);
nand U33914 (N_33914,N_32797,N_32516);
and U33915 (N_33915,N_32117,N_32202);
xnor U33916 (N_33916,N_32176,N_32033);
or U33917 (N_33917,N_32962,N_32330);
nor U33918 (N_33918,N_32123,N_32619);
or U33919 (N_33919,N_32159,N_32292);
xnor U33920 (N_33920,N_32695,N_32233);
or U33921 (N_33921,N_32677,N_32393);
or U33922 (N_33922,N_32495,N_32938);
nand U33923 (N_33923,N_32823,N_32411);
xnor U33924 (N_33924,N_32804,N_32814);
nor U33925 (N_33925,N_32912,N_32297);
or U33926 (N_33926,N_32436,N_32102);
or U33927 (N_33927,N_32187,N_32991);
xnor U33928 (N_33928,N_32190,N_32357);
nor U33929 (N_33929,N_32876,N_32884);
nor U33930 (N_33930,N_32386,N_32470);
and U33931 (N_33931,N_32045,N_32698);
nand U33932 (N_33932,N_32927,N_32730);
or U33933 (N_33933,N_32285,N_32916);
and U33934 (N_33934,N_32802,N_32584);
xor U33935 (N_33935,N_32157,N_32172);
and U33936 (N_33936,N_32731,N_32022);
and U33937 (N_33937,N_32386,N_32975);
or U33938 (N_33938,N_32449,N_32931);
xnor U33939 (N_33939,N_32937,N_32814);
or U33940 (N_33940,N_32924,N_32373);
or U33941 (N_33941,N_32106,N_32008);
or U33942 (N_33942,N_32241,N_32317);
nand U33943 (N_33943,N_32408,N_32644);
nand U33944 (N_33944,N_32685,N_32868);
and U33945 (N_33945,N_32788,N_32565);
xor U33946 (N_33946,N_32422,N_32587);
xnor U33947 (N_33947,N_32301,N_32455);
and U33948 (N_33948,N_32428,N_32024);
or U33949 (N_33949,N_32776,N_32947);
xnor U33950 (N_33950,N_32262,N_32280);
nor U33951 (N_33951,N_32302,N_32289);
and U33952 (N_33952,N_32127,N_32699);
and U33953 (N_33953,N_32549,N_32426);
xnor U33954 (N_33954,N_32754,N_32913);
nor U33955 (N_33955,N_32827,N_32337);
nand U33956 (N_33956,N_32056,N_32706);
nand U33957 (N_33957,N_32418,N_32058);
or U33958 (N_33958,N_32072,N_32818);
and U33959 (N_33959,N_32378,N_32964);
or U33960 (N_33960,N_32405,N_32358);
and U33961 (N_33961,N_32555,N_32873);
and U33962 (N_33962,N_32743,N_32191);
nand U33963 (N_33963,N_32567,N_32646);
or U33964 (N_33964,N_32898,N_32862);
and U33965 (N_33965,N_32486,N_32230);
nand U33966 (N_33966,N_32894,N_32373);
nand U33967 (N_33967,N_32908,N_32581);
and U33968 (N_33968,N_32469,N_32976);
or U33969 (N_33969,N_32283,N_32949);
xnor U33970 (N_33970,N_32899,N_32630);
and U33971 (N_33971,N_32048,N_32060);
or U33972 (N_33972,N_32634,N_32730);
or U33973 (N_33973,N_32034,N_32644);
and U33974 (N_33974,N_32062,N_32906);
or U33975 (N_33975,N_32886,N_32307);
and U33976 (N_33976,N_32206,N_32938);
xnor U33977 (N_33977,N_32508,N_32316);
nor U33978 (N_33978,N_32397,N_32114);
nor U33979 (N_33979,N_32550,N_32296);
nand U33980 (N_33980,N_32818,N_32222);
or U33981 (N_33981,N_32385,N_32897);
xor U33982 (N_33982,N_32117,N_32236);
xnor U33983 (N_33983,N_32034,N_32546);
nor U33984 (N_33984,N_32228,N_32435);
and U33985 (N_33985,N_32074,N_32720);
or U33986 (N_33986,N_32293,N_32288);
xor U33987 (N_33987,N_32838,N_32828);
nand U33988 (N_33988,N_32213,N_32443);
or U33989 (N_33989,N_32616,N_32301);
or U33990 (N_33990,N_32745,N_32105);
nor U33991 (N_33991,N_32343,N_32831);
nand U33992 (N_33992,N_32644,N_32807);
nand U33993 (N_33993,N_32932,N_32252);
or U33994 (N_33994,N_32972,N_32733);
nor U33995 (N_33995,N_32892,N_32043);
xnor U33996 (N_33996,N_32140,N_32808);
and U33997 (N_33997,N_32350,N_32292);
nand U33998 (N_33998,N_32338,N_32226);
xnor U33999 (N_33999,N_32940,N_32845);
nor U34000 (N_34000,N_33606,N_33753);
nor U34001 (N_34001,N_33302,N_33337);
xor U34002 (N_34002,N_33038,N_33636);
xor U34003 (N_34003,N_33679,N_33761);
xnor U34004 (N_34004,N_33994,N_33573);
and U34005 (N_34005,N_33059,N_33001);
and U34006 (N_34006,N_33156,N_33673);
and U34007 (N_34007,N_33411,N_33977);
and U34008 (N_34008,N_33103,N_33381);
nor U34009 (N_34009,N_33541,N_33987);
or U34010 (N_34010,N_33019,N_33435);
nor U34011 (N_34011,N_33667,N_33420);
or U34012 (N_34012,N_33908,N_33115);
nand U34013 (N_34013,N_33783,N_33543);
and U34014 (N_34014,N_33562,N_33384);
nor U34015 (N_34015,N_33932,N_33132);
nand U34016 (N_34016,N_33522,N_33821);
or U34017 (N_34017,N_33093,N_33315);
or U34018 (N_34018,N_33317,N_33427);
and U34019 (N_34019,N_33054,N_33854);
xnor U34020 (N_34020,N_33814,N_33474);
and U34021 (N_34021,N_33726,N_33790);
nor U34022 (N_34022,N_33355,N_33188);
and U34023 (N_34023,N_33508,N_33599);
nor U34024 (N_34024,N_33570,N_33086);
and U34025 (N_34025,N_33918,N_33473);
nand U34026 (N_34026,N_33819,N_33741);
or U34027 (N_34027,N_33476,N_33099);
and U34028 (N_34028,N_33223,N_33561);
nor U34029 (N_34029,N_33364,N_33763);
nor U34030 (N_34030,N_33641,N_33836);
nand U34031 (N_34031,N_33300,N_33074);
or U34032 (N_34032,N_33715,N_33713);
nand U34033 (N_34033,N_33815,N_33375);
or U34034 (N_34034,N_33149,N_33898);
xnor U34035 (N_34035,N_33775,N_33702);
nand U34036 (N_34036,N_33332,N_33963);
nor U34037 (N_34037,N_33523,N_33557);
or U34038 (N_34038,N_33346,N_33799);
nor U34039 (N_34039,N_33654,N_33047);
or U34040 (N_34040,N_33944,N_33878);
xnor U34041 (N_34041,N_33619,N_33926);
nor U34042 (N_34042,N_33436,N_33005);
or U34043 (N_34043,N_33170,N_33382);
nand U34044 (N_34044,N_33579,N_33181);
xnor U34045 (N_34045,N_33246,N_33540);
nand U34046 (N_34046,N_33488,N_33356);
nand U34047 (N_34047,N_33928,N_33394);
xor U34048 (N_34048,N_33198,N_33786);
nand U34049 (N_34049,N_33416,N_33716);
xnor U34050 (N_34050,N_33004,N_33970);
nor U34051 (N_34051,N_33512,N_33992);
or U34052 (N_34052,N_33247,N_33527);
or U34053 (N_34053,N_33470,N_33958);
and U34054 (N_34054,N_33409,N_33901);
nor U34055 (N_34055,N_33389,N_33145);
and U34056 (N_34056,N_33362,N_33954);
nor U34057 (N_34057,N_33805,N_33640);
nor U34058 (N_34058,N_33091,N_33428);
nand U34059 (N_34059,N_33688,N_33581);
and U34060 (N_34060,N_33913,N_33144);
xnor U34061 (N_34061,N_33957,N_33672);
and U34062 (N_34062,N_33870,N_33165);
and U34063 (N_34063,N_33754,N_33485);
nand U34064 (N_34064,N_33275,N_33361);
nor U34065 (N_34065,N_33161,N_33873);
and U34066 (N_34066,N_33069,N_33909);
nor U34067 (N_34067,N_33976,N_33883);
nand U34068 (N_34068,N_33240,N_33016);
nand U34069 (N_34069,N_33772,N_33452);
or U34070 (N_34070,N_33044,N_33244);
nor U34071 (N_34071,N_33169,N_33596);
xnor U34072 (N_34072,N_33830,N_33006);
nor U34073 (N_34073,N_33861,N_33796);
and U34074 (N_34074,N_33351,N_33979);
xor U34075 (N_34075,N_33564,N_33851);
nor U34076 (N_34076,N_33724,N_33229);
or U34077 (N_34077,N_33566,N_33014);
xor U34078 (N_34078,N_33285,N_33127);
nand U34079 (N_34079,N_33270,N_33891);
nor U34080 (N_34080,N_33410,N_33365);
or U34081 (N_34081,N_33077,N_33446);
xnor U34082 (N_34082,N_33262,N_33822);
nand U34083 (N_34083,N_33043,N_33100);
xor U34084 (N_34084,N_33844,N_33113);
nand U34085 (N_34085,N_33139,N_33066);
or U34086 (N_34086,N_33274,N_33785);
nor U34087 (N_34087,N_33721,N_33207);
and U34088 (N_34088,N_33533,N_33261);
nor U34089 (N_34089,N_33937,N_33680);
or U34090 (N_34090,N_33128,N_33493);
nand U34091 (N_34091,N_33153,N_33303);
nor U34092 (N_34092,N_33714,N_33924);
xnor U34093 (N_34093,N_33792,N_33813);
nand U34094 (N_34094,N_33208,N_33960);
and U34095 (N_34095,N_33894,N_33466);
nor U34096 (N_34096,N_33458,N_33867);
xor U34097 (N_34097,N_33310,N_33340);
and U34098 (N_34098,N_33272,N_33020);
or U34099 (N_34099,N_33444,N_33063);
nand U34100 (N_34100,N_33569,N_33395);
and U34101 (N_34101,N_33098,N_33542);
xor U34102 (N_34102,N_33820,N_33407);
nor U34103 (N_34103,N_33853,N_33610);
nor U34104 (N_34104,N_33347,N_33184);
nor U34105 (N_34105,N_33968,N_33053);
and U34106 (N_34106,N_33119,N_33871);
and U34107 (N_34107,N_33973,N_33385);
xnor U34108 (N_34108,N_33808,N_33131);
and U34109 (N_34109,N_33439,N_33108);
nor U34110 (N_34110,N_33765,N_33150);
nand U34111 (N_34111,N_33556,N_33779);
and U34112 (N_34112,N_33035,N_33010);
nor U34113 (N_34113,N_33400,N_33287);
nor U34114 (N_34114,N_33825,N_33391);
xor U34115 (N_34115,N_33612,N_33017);
and U34116 (N_34116,N_33288,N_33218);
nand U34117 (N_34117,N_33080,N_33665);
nand U34118 (N_34118,N_33744,N_33650);
xnor U34119 (N_34119,N_33609,N_33831);
or U34120 (N_34120,N_33434,N_33371);
and U34121 (N_34121,N_33081,N_33794);
nand U34122 (N_34122,N_33206,N_33535);
nor U34123 (N_34123,N_33567,N_33104);
xnor U34124 (N_34124,N_33030,N_33055);
nor U34125 (N_34125,N_33027,N_33191);
nand U34126 (N_34126,N_33848,N_33530);
nand U34127 (N_34127,N_33491,N_33768);
xor U34128 (N_34128,N_33195,N_33734);
nand U34129 (N_34129,N_33157,N_33256);
or U34130 (N_34130,N_33232,N_33866);
and U34131 (N_34131,N_33626,N_33424);
and U34132 (N_34132,N_33746,N_33585);
and U34133 (N_34133,N_33480,N_33777);
and U34134 (N_34134,N_33787,N_33524);
xnor U34135 (N_34135,N_33965,N_33438);
nor U34136 (N_34136,N_33258,N_33986);
xor U34137 (N_34137,N_33216,N_33374);
xor U34138 (N_34138,N_33980,N_33843);
or U34139 (N_34139,N_33916,N_33703);
xor U34140 (N_34140,N_33598,N_33372);
nor U34141 (N_34141,N_33594,N_33348);
or U34142 (N_34142,N_33946,N_33758);
and U34143 (N_34143,N_33600,N_33345);
and U34144 (N_34144,N_33057,N_33141);
xor U34145 (N_34145,N_33631,N_33056);
xnor U34146 (N_34146,N_33759,N_33551);
nand U34147 (N_34147,N_33478,N_33296);
xnor U34148 (N_34148,N_33990,N_33278);
xnor U34149 (N_34149,N_33516,N_33875);
xnor U34150 (N_34150,N_33942,N_33943);
and U34151 (N_34151,N_33972,N_33215);
xor U34152 (N_34152,N_33988,N_33211);
nand U34153 (N_34153,N_33041,N_33290);
nor U34154 (N_34154,N_33621,N_33282);
or U34155 (N_34155,N_33513,N_33496);
nand U34156 (N_34156,N_33902,N_33064);
or U34157 (N_34157,N_33021,N_33964);
xnor U34158 (N_34158,N_33192,N_33605);
nor U34159 (N_34159,N_33417,N_33344);
nor U34160 (N_34160,N_33917,N_33587);
xor U34161 (N_34161,N_33323,N_33118);
xnor U34162 (N_34162,N_33185,N_33291);
or U34163 (N_34163,N_33083,N_33483);
nor U34164 (N_34164,N_33387,N_33430);
and U34165 (N_34165,N_33967,N_33202);
and U34166 (N_34166,N_33433,N_33595);
nor U34167 (N_34167,N_33314,N_33694);
and U34168 (N_34168,N_33525,N_33900);
and U34169 (N_34169,N_33257,N_33903);
and U34170 (N_34170,N_33051,N_33350);
nand U34171 (N_34171,N_33793,N_33255);
nor U34172 (N_34172,N_33766,N_33437);
xnor U34173 (N_34173,N_33975,N_33892);
xor U34174 (N_34174,N_33735,N_33601);
nor U34175 (N_34175,N_33239,N_33137);
nand U34176 (N_34176,N_33869,N_33896);
or U34177 (N_34177,N_33733,N_33868);
nand U34178 (N_34178,N_33187,N_33238);
and U34179 (N_34179,N_33107,N_33668);
xor U34180 (N_34180,N_33426,N_33940);
and U34181 (N_34181,N_33071,N_33265);
or U34182 (N_34182,N_33450,N_33520);
or U34183 (N_34183,N_33408,N_33818);
and U34184 (N_34184,N_33951,N_33681);
xor U34185 (N_34185,N_33653,N_33840);
nand U34186 (N_34186,N_33865,N_33547);
or U34187 (N_34187,N_33085,N_33658);
xnor U34188 (N_34188,N_33927,N_33369);
nor U34189 (N_34189,N_33635,N_33582);
or U34190 (N_34190,N_33817,N_33058);
and U34191 (N_34191,N_33178,N_33518);
nor U34192 (N_34192,N_33778,N_33443);
nor U34193 (N_34193,N_33402,N_33835);
xor U34194 (N_34194,N_33173,N_33620);
and U34195 (N_34195,N_33874,N_33034);
nor U34196 (N_34196,N_33969,N_33625);
nand U34197 (N_34197,N_33396,N_33719);
nor U34198 (N_34198,N_33477,N_33008);
nand U34199 (N_34199,N_33956,N_33329);
nor U34200 (N_34200,N_33463,N_33076);
nor U34201 (N_34201,N_33552,N_33319);
nor U34202 (N_34202,N_33536,N_33320);
or U34203 (N_34203,N_33695,N_33007);
and U34204 (N_34204,N_33683,N_33592);
nand U34205 (N_34205,N_33228,N_33070);
nand U34206 (N_34206,N_33286,N_33684);
and U34207 (N_34207,N_33690,N_33950);
and U34208 (N_34208,N_33897,N_33328);
nor U34209 (N_34209,N_33386,N_33190);
nor U34210 (N_34210,N_33614,N_33697);
xnor U34211 (N_34211,N_33534,N_33560);
nand U34212 (N_34212,N_33378,N_33849);
and U34213 (N_34213,N_33632,N_33171);
and U34214 (N_34214,N_33045,N_33390);
xor U34215 (N_34215,N_33029,N_33294);
nand U34216 (N_34216,N_33441,N_33914);
xnor U34217 (N_34217,N_33116,N_33889);
and U34218 (N_34218,N_33788,N_33728);
xnor U34219 (N_34219,N_33693,N_33698);
nand U34220 (N_34220,N_33800,N_33484);
and U34221 (N_34221,N_33002,N_33780);
or U34222 (N_34222,N_33549,N_33349);
or U34223 (N_34223,N_33062,N_33360);
nand U34224 (N_34224,N_33353,N_33225);
or U34225 (N_34225,N_33826,N_33468);
nand U34226 (N_34226,N_33406,N_33487);
nor U34227 (N_34227,N_33829,N_33065);
nand U34228 (N_34228,N_33706,N_33106);
xnor U34229 (N_34229,N_33893,N_33249);
xnor U34230 (N_34230,N_33529,N_33254);
xor U34231 (N_34231,N_33532,N_33613);
nor U34232 (N_34232,N_33922,N_33597);
nor U34233 (N_34233,N_33399,N_33481);
and U34234 (N_34234,N_33164,N_33642);
nand U34235 (N_34235,N_33061,N_33911);
nand U34236 (N_34236,N_33842,N_33838);
xor U34237 (N_34237,N_33462,N_33284);
and U34238 (N_34238,N_33180,N_33864);
xnor U34239 (N_34239,N_33459,N_33174);
or U34240 (N_34240,N_33649,N_33637);
xnor U34241 (N_34241,N_33243,N_33366);
nand U34242 (N_34242,N_33504,N_33471);
or U34243 (N_34243,N_33558,N_33519);
xor U34244 (N_34244,N_33414,N_33638);
xor U34245 (N_34245,N_33806,N_33890);
nor U34246 (N_34246,N_33862,N_33152);
nand U34247 (N_34247,N_33072,N_33791);
xnor U34248 (N_34248,N_33887,N_33046);
and U34249 (N_34249,N_33906,N_33148);
or U34250 (N_34250,N_33961,N_33507);
xor U34251 (N_34251,N_33280,N_33750);
xnor U34252 (N_34252,N_33380,N_33671);
nor U34253 (N_34253,N_33872,N_33773);
and U34254 (N_34254,N_33945,N_33803);
or U34255 (N_34255,N_33602,N_33431);
nor U34256 (N_34256,N_33675,N_33298);
nor U34257 (N_34257,N_33226,N_33647);
nand U34258 (N_34258,N_33336,N_33096);
nand U34259 (N_34259,N_33774,N_33135);
or U34260 (N_34260,N_33879,N_33196);
nor U34261 (N_34261,N_33939,N_33949);
or U34262 (N_34262,N_33832,N_33451);
nand U34263 (N_34263,N_33616,N_33309);
xor U34264 (N_34264,N_33816,N_33105);
or U34265 (N_34265,N_33357,N_33933);
nor U34266 (N_34266,N_33024,N_33037);
xnor U34267 (N_34267,N_33266,N_33938);
nor U34268 (N_34268,N_33634,N_33651);
nor U34269 (N_34269,N_33147,N_33877);
nor U34270 (N_34270,N_33925,N_33531);
and U34271 (N_34271,N_33730,N_33500);
nand U34272 (N_34272,N_33498,N_33717);
nor U34273 (N_34273,N_33823,N_33517);
nand U34274 (N_34274,N_33656,N_33971);
or U34275 (N_34275,N_33859,N_33112);
nand U34276 (N_34276,N_33807,N_33018);
nand U34277 (N_34277,N_33789,N_33678);
and U34278 (N_34278,N_33326,N_33962);
nor U34279 (N_34279,N_33367,N_33448);
nor U34280 (N_34280,N_33456,N_33904);
and U34281 (N_34281,N_33453,N_33705);
nor U34282 (N_34282,N_33769,N_33253);
and U34283 (N_34283,N_33151,N_33510);
nor U34284 (N_34284,N_33028,N_33335);
nand U34285 (N_34285,N_33669,N_33686);
nor U34286 (N_34286,N_33248,N_33049);
xnor U34287 (N_34287,N_33292,N_33251);
xnor U34288 (N_34288,N_33186,N_33584);
xnor U34289 (N_34289,N_33760,N_33022);
xnor U34290 (N_34290,N_33930,N_33359);
nor U34291 (N_34291,N_33460,N_33267);
nand U34292 (N_34292,N_33664,N_33075);
nor U34293 (N_34293,N_33486,N_33515);
or U34294 (N_34294,N_33179,N_33422);
xnor U34295 (N_34295,N_33217,N_33306);
and U34296 (N_34296,N_33503,N_33289);
nand U34297 (N_34297,N_33997,N_33465);
xnor U34298 (N_34298,N_33200,N_33670);
nor U34299 (N_34299,N_33068,N_33092);
nor U34300 (N_34300,N_33729,N_33123);
and U34301 (N_34301,N_33129,N_33245);
nor U34302 (N_34302,N_33464,N_33089);
nor U34303 (N_34303,N_33067,N_33553);
and U34304 (N_34304,N_33559,N_33078);
nor U34305 (N_34305,N_33824,N_33160);
and U34306 (N_34306,N_33241,N_33327);
and U34307 (N_34307,N_33052,N_33798);
xnor U34308 (N_34308,N_33528,N_33745);
nor U34309 (N_34309,N_33845,N_33795);
and U34310 (N_34310,N_33991,N_33710);
xnor U34311 (N_34311,N_33899,N_33699);
xor U34312 (N_34312,N_33301,N_33757);
nor U34313 (N_34313,N_33628,N_33674);
xnor U34314 (N_34314,N_33687,N_33405);
nand U34315 (N_34315,N_33415,N_33120);
nor U34316 (N_34316,N_33324,N_33172);
xnor U34317 (N_34317,N_33250,N_33401);
xor U34318 (N_34318,N_33989,N_33885);
and U34319 (N_34319,N_33026,N_33648);
and U34320 (N_34320,N_33555,N_33544);
and U34321 (N_34321,N_33727,N_33124);
nand U34322 (N_34322,N_33948,N_33154);
or U34323 (N_34323,N_33352,N_33331);
nor U34324 (N_34324,N_33492,N_33138);
nor U34325 (N_34325,N_33393,N_33125);
and U34326 (N_34326,N_33659,N_33227);
xnor U34327 (N_34327,N_33087,N_33603);
xnor U34328 (N_34328,N_33403,N_33756);
xor U34329 (N_34329,N_33213,N_33645);
xor U34330 (N_34330,N_33677,N_33264);
nand U34331 (N_34331,N_33497,N_33905);
nor U34332 (N_34332,N_33776,N_33935);
and U34333 (N_34333,N_33388,N_33271);
or U34334 (N_34334,N_33999,N_33281);
or U34335 (N_34335,N_33313,N_33880);
and U34336 (N_34336,N_33219,N_33580);
and U34337 (N_34337,N_33804,N_33921);
and U34338 (N_34338,N_33321,N_33467);
or U34339 (N_34339,N_33322,N_33283);
xor U34340 (N_34340,N_33882,N_33575);
and U34341 (N_34341,N_33033,N_33277);
nand U34342 (N_34342,N_33571,N_33847);
and U34343 (N_34343,N_33511,N_33998);
or U34344 (N_34344,N_33852,N_33888);
nor U34345 (N_34345,N_33712,N_33489);
nor U34346 (N_34346,N_33501,N_33031);
and U34347 (N_34347,N_33009,N_33545);
xnor U34348 (N_34348,N_33354,N_33423);
and U34349 (N_34349,N_33259,N_33143);
or U34350 (N_34350,N_33748,N_33182);
or U34351 (N_34351,N_33343,N_33404);
nor U34352 (N_34352,N_33652,N_33781);
xor U34353 (N_34353,N_33981,N_33711);
or U34354 (N_34354,N_33947,N_33455);
xnor U34355 (N_34355,N_33134,N_33234);
xnor U34356 (N_34356,N_33363,N_33368);
nor U34357 (N_34357,N_33342,N_33203);
and U34358 (N_34358,N_33738,N_33725);
and U34359 (N_34359,N_33023,N_33392);
nor U34360 (N_34360,N_33624,N_33231);
and U34361 (N_34361,N_33718,N_33235);
and U34362 (N_34362,N_33025,N_33036);
nor U34363 (N_34363,N_33886,N_33655);
and U34364 (N_34364,N_33111,N_33472);
and U34365 (N_34365,N_33856,N_33447);
nand U34366 (N_34366,N_33577,N_33011);
nand U34367 (N_34367,N_33696,N_33809);
nand U34368 (N_34368,N_33993,N_33136);
nand U34369 (N_34369,N_33088,N_33090);
or U34370 (N_34370,N_33782,N_33884);
and U34371 (N_34371,N_33646,N_33521);
nor U34372 (N_34372,N_33242,N_33784);
or U34373 (N_34373,N_33858,N_33966);
nand U34374 (N_34374,N_33308,N_33316);
nand U34375 (N_34375,N_33469,N_33015);
or U34376 (N_34376,N_33163,N_33742);
nand U34377 (N_34377,N_33048,N_33514);
nor U34378 (N_34378,N_33252,N_33623);
nor U34379 (N_34379,N_33707,N_33537);
nand U34380 (N_34380,N_33212,N_33923);
xnor U34381 (N_34381,N_33617,N_33482);
and U34382 (N_34382,N_33846,N_33221);
and U34383 (N_34383,N_33660,N_33810);
nand U34384 (N_34384,N_33214,N_33565);
and U34385 (N_34385,N_33554,N_33109);
nand U34386 (N_34386,N_33996,N_33931);
and U34387 (N_34387,N_33383,N_33418);
nor U34388 (N_34388,N_33175,N_33593);
and U34389 (N_34389,N_33588,N_33548);
nor U34390 (N_34390,N_33629,N_33692);
nand U34391 (N_34391,N_33627,N_33689);
nor U34392 (N_34392,N_33370,N_33142);
and U34393 (N_34393,N_33012,N_33751);
nor U34394 (N_34394,N_33802,N_33121);
or U34395 (N_34395,N_33722,N_33295);
nor U34396 (N_34396,N_33586,N_33210);
or U34397 (N_34397,N_33102,N_33604);
or U34398 (N_34398,N_33333,N_33495);
and U34399 (N_34399,N_33590,N_33122);
xnor U34400 (N_34400,N_33622,N_33413);
nor U34401 (N_34401,N_33158,N_33506);
xor U34402 (N_34402,N_33701,N_33000);
nor U34403 (N_34403,N_33376,N_33839);
or U34404 (N_34404,N_33720,N_33747);
nor U34405 (N_34405,N_33318,N_33662);
xnor U34406 (N_34406,N_33633,N_33442);
and U34407 (N_34407,N_33984,N_33419);
or U34408 (N_34408,N_33307,N_33084);
nor U34409 (N_34409,N_33140,N_33700);
nor U34410 (N_34410,N_33685,N_33338);
nor U34411 (N_34411,N_33334,N_33490);
nand U34412 (N_34412,N_33762,N_33097);
and U34413 (N_34413,N_33639,N_33339);
nand U34414 (N_34414,N_33572,N_33168);
nor U34415 (N_34415,N_33740,N_33801);
nor U34416 (N_34416,N_33607,N_33855);
or U34417 (N_34417,N_33833,N_33177);
and U34418 (N_34418,N_33297,N_33412);
nor U34419 (N_34419,N_33857,N_33193);
or U34420 (N_34420,N_33941,N_33920);
or U34421 (N_34421,N_33032,N_33094);
xnor U34422 (N_34422,N_33755,N_33978);
xnor U34423 (N_34423,N_33907,N_33189);
and U34424 (N_34424,N_33079,N_33736);
and U34425 (N_34425,N_33919,N_33040);
or U34426 (N_34426,N_33358,N_33276);
or U34427 (N_34427,N_33162,N_33194);
nor U34428 (N_34428,N_33591,N_33657);
xor U34429 (N_34429,N_33666,N_33834);
or U34430 (N_34430,N_33881,N_33305);
nor U34431 (N_34431,N_33130,N_33183);
and U34432 (N_34432,N_33312,N_33959);
or U34433 (N_34433,N_33550,N_33583);
or U34434 (N_34434,N_33159,N_33739);
nor U34435 (N_34435,N_33425,N_33743);
and U34436 (N_34436,N_33475,N_33039);
nor U34437 (N_34437,N_33505,N_33325);
xor U34438 (N_34438,N_33876,N_33379);
nor U34439 (N_34439,N_33863,N_33953);
nand U34440 (N_34440,N_33201,N_33709);
nand U34441 (N_34441,N_33233,N_33767);
and U34442 (N_34442,N_33457,N_33563);
xnor U34443 (N_34443,N_33895,N_33663);
xnor U34444 (N_34444,N_33101,N_33260);
nand U34445 (N_34445,N_33454,N_33828);
nor U34446 (N_34446,N_33220,N_33176);
or U34447 (N_34447,N_33146,N_33731);
and U34448 (N_34448,N_33691,N_33060);
nand U34449 (N_34449,N_33373,N_33910);
nand U34450 (N_34450,N_33797,N_33539);
and U34451 (N_34451,N_33204,N_33311);
or U34452 (N_34452,N_33827,N_33155);
nand U34453 (N_34453,N_33095,N_33749);
and U34454 (N_34454,N_33985,N_33167);
and U34455 (N_34455,N_33509,N_33546);
nand U34456 (N_34456,N_33126,N_33268);
or U34457 (N_34457,N_33421,N_33197);
and U34458 (N_34458,N_33936,N_33279);
and U34459 (N_34459,N_33708,N_33611);
and U34460 (N_34460,N_33723,N_33912);
nand U34461 (N_34461,N_33643,N_33661);
nor U34462 (N_34462,N_33732,N_33538);
and U34463 (N_34463,N_33110,N_33114);
nor U34464 (N_34464,N_33479,N_33752);
and U34465 (N_34465,N_33263,N_33224);
or U34466 (N_34466,N_33502,N_33526);
xor U34467 (N_34467,N_33209,N_33397);
nand U34468 (N_34468,N_33199,N_33704);
nand U34469 (N_34469,N_33952,N_33568);
or U34470 (N_34470,N_33615,N_33133);
and U34471 (N_34471,N_33440,N_33682);
or U34472 (N_34472,N_33737,N_33073);
or U34473 (N_34473,N_33771,N_33013);
nand U34474 (N_34474,N_33578,N_33995);
nor U34475 (N_34475,N_33236,N_33082);
nand U34476 (N_34476,N_33398,N_33983);
nand U34477 (N_34477,N_33330,N_33432);
nor U34478 (N_34478,N_33589,N_33955);
xor U34479 (N_34479,N_33915,N_33166);
or U34480 (N_34480,N_33237,N_33273);
nor U34481 (N_34481,N_33461,N_33841);
nand U34482 (N_34482,N_33449,N_33812);
nand U34483 (N_34483,N_33770,N_33003);
and U34484 (N_34484,N_33304,N_33850);
or U34485 (N_34485,N_33837,N_33630);
and U34486 (N_34486,N_33445,N_33429);
nor U34487 (N_34487,N_33574,N_33042);
nand U34488 (N_34488,N_33974,N_33618);
nor U34489 (N_34489,N_33764,N_33269);
xnor U34490 (N_34490,N_33293,N_33499);
nor U34491 (N_34491,N_33050,N_33934);
nor U34492 (N_34492,N_33576,N_33676);
nand U34493 (N_34493,N_33860,N_33377);
nor U34494 (N_34494,N_33608,N_33230);
and U34495 (N_34495,N_33117,N_33982);
and U34496 (N_34496,N_33811,N_33205);
or U34497 (N_34497,N_33494,N_33299);
nor U34498 (N_34498,N_33929,N_33644);
nand U34499 (N_34499,N_33222,N_33341);
xor U34500 (N_34500,N_33054,N_33734);
or U34501 (N_34501,N_33237,N_33754);
xor U34502 (N_34502,N_33538,N_33428);
nand U34503 (N_34503,N_33724,N_33577);
or U34504 (N_34504,N_33018,N_33219);
and U34505 (N_34505,N_33529,N_33869);
nor U34506 (N_34506,N_33799,N_33595);
or U34507 (N_34507,N_33175,N_33490);
xnor U34508 (N_34508,N_33030,N_33972);
nand U34509 (N_34509,N_33436,N_33302);
nand U34510 (N_34510,N_33568,N_33836);
nor U34511 (N_34511,N_33476,N_33054);
or U34512 (N_34512,N_33849,N_33312);
nand U34513 (N_34513,N_33500,N_33198);
and U34514 (N_34514,N_33810,N_33424);
nor U34515 (N_34515,N_33276,N_33692);
nand U34516 (N_34516,N_33671,N_33284);
and U34517 (N_34517,N_33657,N_33380);
nor U34518 (N_34518,N_33977,N_33175);
nand U34519 (N_34519,N_33287,N_33984);
or U34520 (N_34520,N_33192,N_33607);
or U34521 (N_34521,N_33052,N_33381);
or U34522 (N_34522,N_33195,N_33613);
xor U34523 (N_34523,N_33427,N_33862);
nand U34524 (N_34524,N_33725,N_33719);
and U34525 (N_34525,N_33136,N_33601);
xor U34526 (N_34526,N_33795,N_33416);
xnor U34527 (N_34527,N_33905,N_33738);
xnor U34528 (N_34528,N_33609,N_33296);
or U34529 (N_34529,N_33594,N_33740);
nand U34530 (N_34530,N_33895,N_33227);
and U34531 (N_34531,N_33626,N_33242);
nor U34532 (N_34532,N_33647,N_33578);
xor U34533 (N_34533,N_33547,N_33479);
xnor U34534 (N_34534,N_33213,N_33001);
xnor U34535 (N_34535,N_33301,N_33673);
nand U34536 (N_34536,N_33573,N_33745);
xor U34537 (N_34537,N_33580,N_33054);
nand U34538 (N_34538,N_33433,N_33270);
and U34539 (N_34539,N_33412,N_33520);
nor U34540 (N_34540,N_33479,N_33827);
or U34541 (N_34541,N_33191,N_33703);
nor U34542 (N_34542,N_33116,N_33392);
nand U34543 (N_34543,N_33236,N_33696);
nand U34544 (N_34544,N_33308,N_33093);
or U34545 (N_34545,N_33939,N_33512);
xor U34546 (N_34546,N_33992,N_33484);
and U34547 (N_34547,N_33184,N_33270);
xnor U34548 (N_34548,N_33510,N_33845);
and U34549 (N_34549,N_33981,N_33225);
nand U34550 (N_34550,N_33993,N_33946);
nor U34551 (N_34551,N_33212,N_33314);
xnor U34552 (N_34552,N_33083,N_33599);
or U34553 (N_34553,N_33134,N_33431);
or U34554 (N_34554,N_33361,N_33293);
nor U34555 (N_34555,N_33548,N_33665);
nand U34556 (N_34556,N_33119,N_33916);
nand U34557 (N_34557,N_33015,N_33933);
nand U34558 (N_34558,N_33880,N_33995);
nor U34559 (N_34559,N_33865,N_33739);
nand U34560 (N_34560,N_33612,N_33341);
xor U34561 (N_34561,N_33831,N_33647);
and U34562 (N_34562,N_33359,N_33602);
nor U34563 (N_34563,N_33597,N_33311);
or U34564 (N_34564,N_33338,N_33545);
or U34565 (N_34565,N_33414,N_33062);
xnor U34566 (N_34566,N_33867,N_33052);
or U34567 (N_34567,N_33700,N_33068);
nor U34568 (N_34568,N_33021,N_33135);
and U34569 (N_34569,N_33881,N_33787);
nor U34570 (N_34570,N_33319,N_33784);
nor U34571 (N_34571,N_33723,N_33119);
and U34572 (N_34572,N_33246,N_33316);
xnor U34573 (N_34573,N_33682,N_33423);
nor U34574 (N_34574,N_33073,N_33877);
nor U34575 (N_34575,N_33060,N_33114);
xnor U34576 (N_34576,N_33530,N_33808);
or U34577 (N_34577,N_33970,N_33643);
xor U34578 (N_34578,N_33294,N_33099);
or U34579 (N_34579,N_33196,N_33854);
or U34580 (N_34580,N_33129,N_33877);
nand U34581 (N_34581,N_33680,N_33819);
xnor U34582 (N_34582,N_33132,N_33741);
nor U34583 (N_34583,N_33438,N_33057);
or U34584 (N_34584,N_33511,N_33778);
or U34585 (N_34585,N_33649,N_33319);
nand U34586 (N_34586,N_33264,N_33551);
xor U34587 (N_34587,N_33787,N_33208);
and U34588 (N_34588,N_33085,N_33296);
nand U34589 (N_34589,N_33342,N_33668);
or U34590 (N_34590,N_33137,N_33743);
or U34591 (N_34591,N_33502,N_33977);
and U34592 (N_34592,N_33729,N_33072);
nand U34593 (N_34593,N_33953,N_33877);
and U34594 (N_34594,N_33445,N_33996);
nand U34595 (N_34595,N_33824,N_33090);
or U34596 (N_34596,N_33941,N_33132);
nor U34597 (N_34597,N_33291,N_33540);
and U34598 (N_34598,N_33422,N_33926);
or U34599 (N_34599,N_33394,N_33417);
or U34600 (N_34600,N_33979,N_33617);
nor U34601 (N_34601,N_33634,N_33423);
and U34602 (N_34602,N_33490,N_33455);
or U34603 (N_34603,N_33598,N_33479);
and U34604 (N_34604,N_33541,N_33983);
nor U34605 (N_34605,N_33730,N_33405);
xnor U34606 (N_34606,N_33407,N_33595);
or U34607 (N_34607,N_33391,N_33517);
and U34608 (N_34608,N_33549,N_33511);
xor U34609 (N_34609,N_33210,N_33473);
nand U34610 (N_34610,N_33455,N_33447);
and U34611 (N_34611,N_33328,N_33112);
and U34612 (N_34612,N_33170,N_33277);
xnor U34613 (N_34613,N_33829,N_33316);
xnor U34614 (N_34614,N_33531,N_33950);
or U34615 (N_34615,N_33141,N_33259);
and U34616 (N_34616,N_33808,N_33248);
nand U34617 (N_34617,N_33165,N_33779);
nand U34618 (N_34618,N_33686,N_33323);
or U34619 (N_34619,N_33101,N_33298);
nor U34620 (N_34620,N_33656,N_33283);
nor U34621 (N_34621,N_33052,N_33672);
and U34622 (N_34622,N_33684,N_33710);
and U34623 (N_34623,N_33371,N_33648);
nand U34624 (N_34624,N_33352,N_33414);
nand U34625 (N_34625,N_33413,N_33753);
or U34626 (N_34626,N_33745,N_33100);
nor U34627 (N_34627,N_33916,N_33120);
nor U34628 (N_34628,N_33073,N_33758);
and U34629 (N_34629,N_33786,N_33278);
nor U34630 (N_34630,N_33728,N_33105);
or U34631 (N_34631,N_33389,N_33273);
and U34632 (N_34632,N_33545,N_33574);
or U34633 (N_34633,N_33268,N_33638);
nor U34634 (N_34634,N_33055,N_33740);
and U34635 (N_34635,N_33939,N_33384);
nand U34636 (N_34636,N_33540,N_33810);
nand U34637 (N_34637,N_33912,N_33638);
xnor U34638 (N_34638,N_33471,N_33631);
xor U34639 (N_34639,N_33333,N_33126);
xor U34640 (N_34640,N_33797,N_33873);
or U34641 (N_34641,N_33696,N_33110);
or U34642 (N_34642,N_33188,N_33832);
and U34643 (N_34643,N_33261,N_33739);
and U34644 (N_34644,N_33677,N_33905);
xor U34645 (N_34645,N_33079,N_33419);
nand U34646 (N_34646,N_33435,N_33398);
and U34647 (N_34647,N_33515,N_33301);
nor U34648 (N_34648,N_33313,N_33164);
nand U34649 (N_34649,N_33544,N_33517);
or U34650 (N_34650,N_33386,N_33788);
and U34651 (N_34651,N_33488,N_33089);
xnor U34652 (N_34652,N_33493,N_33322);
nand U34653 (N_34653,N_33181,N_33269);
and U34654 (N_34654,N_33890,N_33759);
and U34655 (N_34655,N_33691,N_33226);
nor U34656 (N_34656,N_33705,N_33416);
or U34657 (N_34657,N_33634,N_33835);
nor U34658 (N_34658,N_33537,N_33541);
nor U34659 (N_34659,N_33126,N_33754);
and U34660 (N_34660,N_33650,N_33001);
and U34661 (N_34661,N_33907,N_33311);
xor U34662 (N_34662,N_33062,N_33995);
and U34663 (N_34663,N_33354,N_33550);
xor U34664 (N_34664,N_33232,N_33762);
nand U34665 (N_34665,N_33352,N_33165);
nand U34666 (N_34666,N_33764,N_33361);
and U34667 (N_34667,N_33671,N_33974);
nor U34668 (N_34668,N_33604,N_33764);
and U34669 (N_34669,N_33542,N_33260);
and U34670 (N_34670,N_33419,N_33267);
and U34671 (N_34671,N_33369,N_33169);
nand U34672 (N_34672,N_33967,N_33154);
and U34673 (N_34673,N_33006,N_33368);
and U34674 (N_34674,N_33496,N_33137);
xnor U34675 (N_34675,N_33444,N_33941);
or U34676 (N_34676,N_33091,N_33634);
and U34677 (N_34677,N_33811,N_33338);
and U34678 (N_34678,N_33278,N_33125);
and U34679 (N_34679,N_33984,N_33505);
nor U34680 (N_34680,N_33412,N_33234);
and U34681 (N_34681,N_33546,N_33777);
nor U34682 (N_34682,N_33289,N_33234);
nand U34683 (N_34683,N_33743,N_33305);
nand U34684 (N_34684,N_33635,N_33637);
nor U34685 (N_34685,N_33965,N_33090);
nand U34686 (N_34686,N_33917,N_33742);
nand U34687 (N_34687,N_33290,N_33156);
or U34688 (N_34688,N_33296,N_33650);
and U34689 (N_34689,N_33014,N_33586);
and U34690 (N_34690,N_33979,N_33265);
or U34691 (N_34691,N_33400,N_33896);
nand U34692 (N_34692,N_33414,N_33135);
and U34693 (N_34693,N_33368,N_33095);
nor U34694 (N_34694,N_33037,N_33515);
nor U34695 (N_34695,N_33991,N_33429);
xor U34696 (N_34696,N_33931,N_33829);
nand U34697 (N_34697,N_33180,N_33741);
xnor U34698 (N_34698,N_33045,N_33488);
nor U34699 (N_34699,N_33426,N_33929);
or U34700 (N_34700,N_33908,N_33085);
or U34701 (N_34701,N_33595,N_33468);
or U34702 (N_34702,N_33238,N_33257);
xor U34703 (N_34703,N_33826,N_33405);
nand U34704 (N_34704,N_33067,N_33760);
nand U34705 (N_34705,N_33661,N_33445);
and U34706 (N_34706,N_33080,N_33434);
nand U34707 (N_34707,N_33347,N_33197);
nand U34708 (N_34708,N_33319,N_33943);
and U34709 (N_34709,N_33434,N_33381);
nand U34710 (N_34710,N_33487,N_33218);
xor U34711 (N_34711,N_33621,N_33105);
nor U34712 (N_34712,N_33294,N_33011);
nand U34713 (N_34713,N_33585,N_33782);
or U34714 (N_34714,N_33808,N_33848);
nand U34715 (N_34715,N_33008,N_33763);
nor U34716 (N_34716,N_33976,N_33326);
xnor U34717 (N_34717,N_33951,N_33465);
nand U34718 (N_34718,N_33742,N_33714);
nand U34719 (N_34719,N_33427,N_33712);
xnor U34720 (N_34720,N_33474,N_33336);
nand U34721 (N_34721,N_33911,N_33127);
or U34722 (N_34722,N_33980,N_33631);
or U34723 (N_34723,N_33422,N_33771);
or U34724 (N_34724,N_33530,N_33035);
nand U34725 (N_34725,N_33158,N_33222);
nor U34726 (N_34726,N_33957,N_33119);
nor U34727 (N_34727,N_33631,N_33077);
and U34728 (N_34728,N_33316,N_33517);
or U34729 (N_34729,N_33150,N_33369);
or U34730 (N_34730,N_33507,N_33139);
nand U34731 (N_34731,N_33695,N_33566);
nand U34732 (N_34732,N_33628,N_33602);
nand U34733 (N_34733,N_33271,N_33658);
and U34734 (N_34734,N_33251,N_33226);
nor U34735 (N_34735,N_33273,N_33966);
or U34736 (N_34736,N_33382,N_33899);
nor U34737 (N_34737,N_33800,N_33095);
or U34738 (N_34738,N_33631,N_33661);
or U34739 (N_34739,N_33372,N_33494);
nor U34740 (N_34740,N_33989,N_33895);
xnor U34741 (N_34741,N_33632,N_33817);
nor U34742 (N_34742,N_33750,N_33213);
nor U34743 (N_34743,N_33687,N_33642);
or U34744 (N_34744,N_33912,N_33820);
nor U34745 (N_34745,N_33938,N_33392);
nand U34746 (N_34746,N_33134,N_33283);
nor U34747 (N_34747,N_33655,N_33748);
nor U34748 (N_34748,N_33721,N_33024);
xor U34749 (N_34749,N_33254,N_33684);
xnor U34750 (N_34750,N_33028,N_33759);
nand U34751 (N_34751,N_33703,N_33643);
xor U34752 (N_34752,N_33284,N_33841);
xor U34753 (N_34753,N_33885,N_33622);
and U34754 (N_34754,N_33807,N_33712);
nand U34755 (N_34755,N_33898,N_33790);
and U34756 (N_34756,N_33290,N_33670);
nor U34757 (N_34757,N_33216,N_33152);
nand U34758 (N_34758,N_33092,N_33757);
nor U34759 (N_34759,N_33470,N_33095);
or U34760 (N_34760,N_33907,N_33709);
and U34761 (N_34761,N_33987,N_33095);
or U34762 (N_34762,N_33573,N_33496);
nor U34763 (N_34763,N_33718,N_33825);
xnor U34764 (N_34764,N_33287,N_33006);
nand U34765 (N_34765,N_33603,N_33140);
and U34766 (N_34766,N_33245,N_33356);
xor U34767 (N_34767,N_33173,N_33879);
xor U34768 (N_34768,N_33119,N_33309);
or U34769 (N_34769,N_33591,N_33491);
nand U34770 (N_34770,N_33817,N_33779);
nor U34771 (N_34771,N_33906,N_33133);
nor U34772 (N_34772,N_33987,N_33788);
nand U34773 (N_34773,N_33989,N_33941);
nand U34774 (N_34774,N_33071,N_33094);
nor U34775 (N_34775,N_33687,N_33081);
or U34776 (N_34776,N_33603,N_33039);
or U34777 (N_34777,N_33377,N_33337);
or U34778 (N_34778,N_33644,N_33806);
and U34779 (N_34779,N_33298,N_33175);
nand U34780 (N_34780,N_33580,N_33330);
nand U34781 (N_34781,N_33884,N_33200);
and U34782 (N_34782,N_33042,N_33258);
or U34783 (N_34783,N_33843,N_33446);
and U34784 (N_34784,N_33956,N_33562);
or U34785 (N_34785,N_33766,N_33323);
or U34786 (N_34786,N_33255,N_33773);
or U34787 (N_34787,N_33387,N_33213);
or U34788 (N_34788,N_33875,N_33696);
and U34789 (N_34789,N_33629,N_33882);
or U34790 (N_34790,N_33342,N_33657);
nand U34791 (N_34791,N_33723,N_33903);
nand U34792 (N_34792,N_33121,N_33663);
nor U34793 (N_34793,N_33344,N_33761);
xnor U34794 (N_34794,N_33376,N_33923);
nand U34795 (N_34795,N_33347,N_33487);
or U34796 (N_34796,N_33114,N_33443);
or U34797 (N_34797,N_33489,N_33909);
nor U34798 (N_34798,N_33030,N_33304);
nand U34799 (N_34799,N_33377,N_33629);
nand U34800 (N_34800,N_33116,N_33668);
or U34801 (N_34801,N_33970,N_33506);
nor U34802 (N_34802,N_33185,N_33678);
and U34803 (N_34803,N_33693,N_33431);
nand U34804 (N_34804,N_33656,N_33096);
nand U34805 (N_34805,N_33832,N_33397);
nand U34806 (N_34806,N_33897,N_33626);
nand U34807 (N_34807,N_33950,N_33434);
or U34808 (N_34808,N_33048,N_33076);
nor U34809 (N_34809,N_33142,N_33242);
or U34810 (N_34810,N_33861,N_33262);
nor U34811 (N_34811,N_33926,N_33578);
nor U34812 (N_34812,N_33672,N_33336);
nand U34813 (N_34813,N_33533,N_33684);
or U34814 (N_34814,N_33991,N_33507);
nor U34815 (N_34815,N_33267,N_33691);
nor U34816 (N_34816,N_33044,N_33169);
nor U34817 (N_34817,N_33628,N_33953);
nand U34818 (N_34818,N_33732,N_33946);
nor U34819 (N_34819,N_33868,N_33983);
xor U34820 (N_34820,N_33952,N_33432);
and U34821 (N_34821,N_33500,N_33598);
nand U34822 (N_34822,N_33621,N_33245);
nor U34823 (N_34823,N_33372,N_33684);
nand U34824 (N_34824,N_33350,N_33783);
nand U34825 (N_34825,N_33018,N_33178);
nor U34826 (N_34826,N_33635,N_33279);
nand U34827 (N_34827,N_33564,N_33731);
nand U34828 (N_34828,N_33359,N_33164);
nor U34829 (N_34829,N_33129,N_33043);
and U34830 (N_34830,N_33095,N_33762);
and U34831 (N_34831,N_33806,N_33620);
nor U34832 (N_34832,N_33378,N_33837);
xor U34833 (N_34833,N_33189,N_33331);
xnor U34834 (N_34834,N_33842,N_33050);
and U34835 (N_34835,N_33905,N_33048);
or U34836 (N_34836,N_33918,N_33176);
nand U34837 (N_34837,N_33737,N_33226);
or U34838 (N_34838,N_33896,N_33273);
nor U34839 (N_34839,N_33361,N_33224);
nand U34840 (N_34840,N_33444,N_33187);
xnor U34841 (N_34841,N_33823,N_33726);
nand U34842 (N_34842,N_33869,N_33032);
or U34843 (N_34843,N_33426,N_33552);
and U34844 (N_34844,N_33836,N_33994);
nor U34845 (N_34845,N_33511,N_33925);
xnor U34846 (N_34846,N_33955,N_33692);
nand U34847 (N_34847,N_33757,N_33277);
and U34848 (N_34848,N_33430,N_33840);
or U34849 (N_34849,N_33175,N_33351);
xnor U34850 (N_34850,N_33806,N_33427);
and U34851 (N_34851,N_33382,N_33291);
xor U34852 (N_34852,N_33388,N_33525);
nor U34853 (N_34853,N_33159,N_33788);
xnor U34854 (N_34854,N_33872,N_33479);
xor U34855 (N_34855,N_33197,N_33390);
and U34856 (N_34856,N_33373,N_33132);
or U34857 (N_34857,N_33345,N_33074);
and U34858 (N_34858,N_33311,N_33030);
nand U34859 (N_34859,N_33908,N_33987);
nor U34860 (N_34860,N_33683,N_33694);
and U34861 (N_34861,N_33785,N_33618);
and U34862 (N_34862,N_33074,N_33491);
and U34863 (N_34863,N_33135,N_33430);
nand U34864 (N_34864,N_33853,N_33674);
or U34865 (N_34865,N_33389,N_33793);
and U34866 (N_34866,N_33622,N_33331);
or U34867 (N_34867,N_33541,N_33258);
and U34868 (N_34868,N_33416,N_33809);
nor U34869 (N_34869,N_33887,N_33242);
nor U34870 (N_34870,N_33033,N_33479);
nor U34871 (N_34871,N_33073,N_33393);
nor U34872 (N_34872,N_33942,N_33173);
and U34873 (N_34873,N_33824,N_33374);
nor U34874 (N_34874,N_33991,N_33224);
and U34875 (N_34875,N_33451,N_33093);
and U34876 (N_34876,N_33435,N_33463);
xor U34877 (N_34877,N_33975,N_33903);
xor U34878 (N_34878,N_33307,N_33384);
xnor U34879 (N_34879,N_33643,N_33173);
xnor U34880 (N_34880,N_33809,N_33209);
or U34881 (N_34881,N_33599,N_33648);
and U34882 (N_34882,N_33318,N_33360);
nand U34883 (N_34883,N_33320,N_33251);
or U34884 (N_34884,N_33005,N_33455);
or U34885 (N_34885,N_33837,N_33062);
nand U34886 (N_34886,N_33671,N_33983);
and U34887 (N_34887,N_33231,N_33651);
nand U34888 (N_34888,N_33644,N_33378);
nand U34889 (N_34889,N_33506,N_33665);
xor U34890 (N_34890,N_33447,N_33982);
or U34891 (N_34891,N_33085,N_33854);
xnor U34892 (N_34892,N_33014,N_33758);
xnor U34893 (N_34893,N_33519,N_33643);
or U34894 (N_34894,N_33945,N_33323);
and U34895 (N_34895,N_33766,N_33177);
nor U34896 (N_34896,N_33681,N_33825);
nor U34897 (N_34897,N_33835,N_33749);
nand U34898 (N_34898,N_33153,N_33380);
nor U34899 (N_34899,N_33705,N_33618);
xnor U34900 (N_34900,N_33092,N_33418);
and U34901 (N_34901,N_33958,N_33568);
xnor U34902 (N_34902,N_33696,N_33779);
nand U34903 (N_34903,N_33124,N_33955);
nor U34904 (N_34904,N_33841,N_33830);
and U34905 (N_34905,N_33714,N_33731);
or U34906 (N_34906,N_33702,N_33360);
nand U34907 (N_34907,N_33500,N_33873);
nand U34908 (N_34908,N_33187,N_33734);
nand U34909 (N_34909,N_33192,N_33183);
nand U34910 (N_34910,N_33545,N_33167);
or U34911 (N_34911,N_33985,N_33168);
nor U34912 (N_34912,N_33189,N_33696);
nor U34913 (N_34913,N_33127,N_33966);
and U34914 (N_34914,N_33528,N_33501);
nand U34915 (N_34915,N_33979,N_33071);
nand U34916 (N_34916,N_33797,N_33299);
nand U34917 (N_34917,N_33367,N_33606);
nor U34918 (N_34918,N_33804,N_33146);
nor U34919 (N_34919,N_33864,N_33962);
nand U34920 (N_34920,N_33944,N_33415);
nand U34921 (N_34921,N_33557,N_33071);
and U34922 (N_34922,N_33865,N_33156);
xor U34923 (N_34923,N_33356,N_33007);
and U34924 (N_34924,N_33712,N_33162);
xnor U34925 (N_34925,N_33455,N_33887);
or U34926 (N_34926,N_33527,N_33822);
xnor U34927 (N_34927,N_33959,N_33189);
nand U34928 (N_34928,N_33049,N_33428);
or U34929 (N_34929,N_33870,N_33238);
xnor U34930 (N_34930,N_33271,N_33775);
and U34931 (N_34931,N_33899,N_33565);
and U34932 (N_34932,N_33263,N_33992);
nand U34933 (N_34933,N_33662,N_33600);
nand U34934 (N_34934,N_33072,N_33455);
nor U34935 (N_34935,N_33150,N_33890);
nor U34936 (N_34936,N_33105,N_33216);
xnor U34937 (N_34937,N_33918,N_33150);
nand U34938 (N_34938,N_33883,N_33997);
nor U34939 (N_34939,N_33894,N_33751);
nor U34940 (N_34940,N_33884,N_33181);
nand U34941 (N_34941,N_33593,N_33634);
or U34942 (N_34942,N_33527,N_33535);
and U34943 (N_34943,N_33987,N_33108);
xor U34944 (N_34944,N_33186,N_33361);
xnor U34945 (N_34945,N_33959,N_33251);
or U34946 (N_34946,N_33044,N_33035);
and U34947 (N_34947,N_33837,N_33195);
and U34948 (N_34948,N_33625,N_33428);
and U34949 (N_34949,N_33848,N_33356);
and U34950 (N_34950,N_33349,N_33777);
nand U34951 (N_34951,N_33691,N_33802);
xnor U34952 (N_34952,N_33497,N_33123);
nand U34953 (N_34953,N_33568,N_33519);
nor U34954 (N_34954,N_33446,N_33113);
nor U34955 (N_34955,N_33344,N_33716);
and U34956 (N_34956,N_33912,N_33243);
or U34957 (N_34957,N_33345,N_33863);
and U34958 (N_34958,N_33669,N_33743);
nor U34959 (N_34959,N_33255,N_33283);
nor U34960 (N_34960,N_33619,N_33291);
nor U34961 (N_34961,N_33151,N_33673);
xnor U34962 (N_34962,N_33678,N_33686);
and U34963 (N_34963,N_33114,N_33441);
xnor U34964 (N_34964,N_33887,N_33520);
xnor U34965 (N_34965,N_33381,N_33481);
or U34966 (N_34966,N_33618,N_33827);
nor U34967 (N_34967,N_33019,N_33605);
xor U34968 (N_34968,N_33379,N_33975);
and U34969 (N_34969,N_33002,N_33474);
and U34970 (N_34970,N_33445,N_33531);
nor U34971 (N_34971,N_33862,N_33595);
nand U34972 (N_34972,N_33802,N_33771);
nor U34973 (N_34973,N_33470,N_33884);
nor U34974 (N_34974,N_33484,N_33784);
nor U34975 (N_34975,N_33711,N_33585);
nor U34976 (N_34976,N_33672,N_33407);
or U34977 (N_34977,N_33926,N_33345);
and U34978 (N_34978,N_33056,N_33574);
nor U34979 (N_34979,N_33204,N_33256);
or U34980 (N_34980,N_33195,N_33046);
and U34981 (N_34981,N_33065,N_33123);
and U34982 (N_34982,N_33939,N_33277);
nand U34983 (N_34983,N_33608,N_33494);
or U34984 (N_34984,N_33154,N_33684);
nand U34985 (N_34985,N_33728,N_33045);
nand U34986 (N_34986,N_33543,N_33296);
nor U34987 (N_34987,N_33174,N_33382);
nor U34988 (N_34988,N_33247,N_33038);
and U34989 (N_34989,N_33841,N_33723);
nand U34990 (N_34990,N_33960,N_33127);
and U34991 (N_34991,N_33129,N_33158);
and U34992 (N_34992,N_33100,N_33242);
and U34993 (N_34993,N_33245,N_33054);
or U34994 (N_34994,N_33356,N_33492);
or U34995 (N_34995,N_33907,N_33691);
xor U34996 (N_34996,N_33047,N_33961);
xnor U34997 (N_34997,N_33725,N_33514);
nor U34998 (N_34998,N_33954,N_33411);
and U34999 (N_34999,N_33958,N_33791);
or U35000 (N_35000,N_34269,N_34637);
nand U35001 (N_35001,N_34194,N_34654);
nor U35002 (N_35002,N_34569,N_34847);
nand U35003 (N_35003,N_34386,N_34243);
nand U35004 (N_35004,N_34490,N_34000);
and U35005 (N_35005,N_34079,N_34875);
xor U35006 (N_35006,N_34617,N_34122);
nand U35007 (N_35007,N_34533,N_34994);
nor U35008 (N_35008,N_34987,N_34305);
nor U35009 (N_35009,N_34620,N_34754);
xnor U35010 (N_35010,N_34717,N_34737);
nor U35011 (N_35011,N_34170,N_34995);
and U35012 (N_35012,N_34306,N_34325);
nand U35013 (N_35013,N_34117,N_34380);
nand U35014 (N_35014,N_34034,N_34059);
xor U35015 (N_35015,N_34822,N_34403);
nor U35016 (N_35016,N_34963,N_34732);
or U35017 (N_35017,N_34169,N_34765);
nor U35018 (N_35018,N_34558,N_34268);
or U35019 (N_35019,N_34592,N_34369);
xor U35020 (N_35020,N_34708,N_34265);
nand U35021 (N_35021,N_34772,N_34488);
nand U35022 (N_35022,N_34580,N_34352);
nor U35023 (N_35023,N_34090,N_34223);
nand U35024 (N_35024,N_34158,N_34573);
or U35025 (N_35025,N_34334,N_34843);
or U35026 (N_35026,N_34798,N_34048);
nand U35027 (N_35027,N_34162,N_34249);
nor U35028 (N_35028,N_34586,N_34433);
and U35029 (N_35029,N_34092,N_34939);
nand U35030 (N_35030,N_34787,N_34021);
nor U35031 (N_35031,N_34493,N_34944);
xnor U35032 (N_35032,N_34201,N_34685);
nand U35033 (N_35033,N_34814,N_34665);
or U35034 (N_35034,N_34166,N_34662);
or U35035 (N_35035,N_34590,N_34983);
or U35036 (N_35036,N_34095,N_34979);
xor U35037 (N_35037,N_34553,N_34360);
xnor U35038 (N_35038,N_34474,N_34686);
nand U35039 (N_35039,N_34317,N_34485);
nand U35040 (N_35040,N_34093,N_34812);
or U35041 (N_35041,N_34005,N_34509);
xor U35042 (N_35042,N_34709,N_34807);
nand U35043 (N_35043,N_34964,N_34755);
nand U35044 (N_35044,N_34228,N_34257);
nor U35045 (N_35045,N_34751,N_34954);
and U35046 (N_35046,N_34328,N_34153);
xor U35047 (N_35047,N_34279,N_34706);
nand U35048 (N_35048,N_34358,N_34029);
nor U35049 (N_35049,N_34237,N_34703);
nor U35050 (N_35050,N_34978,N_34546);
nand U35051 (N_35051,N_34027,N_34714);
xnor U35052 (N_35052,N_34813,N_34971);
or U35053 (N_35053,N_34037,N_34862);
nand U35054 (N_35054,N_34625,N_34072);
nor U35055 (N_35055,N_34436,N_34652);
or U35056 (N_35056,N_34486,N_34332);
nor U35057 (N_35057,N_34702,N_34348);
nor U35058 (N_35058,N_34596,N_34389);
and U35059 (N_35059,N_34776,N_34628);
nor U35060 (N_35060,N_34977,N_34413);
or U35061 (N_35061,N_34478,N_34871);
and U35062 (N_35062,N_34529,N_34456);
and U35063 (N_35063,N_34922,N_34442);
xor U35064 (N_35064,N_34152,N_34541);
nand U35065 (N_35065,N_34868,N_34672);
nand U35066 (N_35066,N_34653,N_34361);
xnor U35067 (N_35067,N_34700,N_34479);
xnor U35068 (N_35068,N_34163,N_34668);
and U35069 (N_35069,N_34552,N_34419);
xnor U35070 (N_35070,N_34125,N_34324);
nor U35071 (N_35071,N_34658,N_34312);
nand U35072 (N_35072,N_34659,N_34086);
nor U35073 (N_35073,N_34316,N_34976);
xor U35074 (N_35074,N_34118,N_34213);
and U35075 (N_35075,N_34376,N_34182);
or U35076 (N_35076,N_34252,N_34982);
and U35077 (N_35077,N_34323,N_34344);
nor U35078 (N_35078,N_34864,N_34736);
and U35079 (N_35079,N_34715,N_34180);
and U35080 (N_35080,N_34865,N_34101);
nor U35081 (N_35081,N_34384,N_34804);
or U35082 (N_35082,N_34970,N_34632);
nand U35083 (N_35083,N_34296,N_34743);
nor U35084 (N_35084,N_34444,N_34147);
nor U35085 (N_35085,N_34164,N_34599);
nor U35086 (N_35086,N_34365,N_34933);
xor U35087 (N_35087,N_34796,N_34450);
nand U35088 (N_35088,N_34507,N_34004);
and U35089 (N_35089,N_34378,N_34565);
xnor U35090 (N_35090,N_34886,N_34629);
or U35091 (N_35091,N_34713,N_34974);
nand U35092 (N_35092,N_34575,N_34879);
and U35093 (N_35093,N_34260,N_34908);
nor U35094 (N_35094,N_34689,N_34400);
or U35095 (N_35095,N_34791,N_34402);
or U35096 (N_35096,N_34461,N_34351);
and U35097 (N_35097,N_34115,N_34530);
nand U35098 (N_35098,N_34189,N_34275);
xor U35099 (N_35099,N_34437,N_34267);
nor U35100 (N_35100,N_34966,N_34300);
or U35101 (N_35101,N_34844,N_34506);
nand U35102 (N_35102,N_34564,N_34199);
nor U35103 (N_35103,N_34934,N_34354);
nand U35104 (N_35104,N_34539,N_34462);
nand U35105 (N_35105,N_34256,N_34457);
xor U35106 (N_35106,N_34128,N_34587);
and U35107 (N_35107,N_34941,N_34283);
and U35108 (N_35108,N_34497,N_34947);
nor U35109 (N_35109,N_34626,N_34366);
or U35110 (N_35110,N_34320,N_34621);
nand U35111 (N_35111,N_34061,N_34399);
xnor U35112 (N_35112,N_34661,N_34721);
nand U35113 (N_35113,N_34171,N_34640);
and U35114 (N_35114,N_34234,N_34028);
xnor U35115 (N_35115,N_34921,N_34423);
nor U35116 (N_35116,N_34192,N_34741);
and U35117 (N_35117,N_34014,N_34438);
xnor U35118 (N_35118,N_34742,N_34286);
nor U35119 (N_35119,N_34955,N_34285);
nand U35120 (N_35120,N_34032,N_34420);
and U35121 (N_35121,N_34321,N_34889);
xor U35122 (N_35122,N_34753,N_34815);
or U35123 (N_35123,N_34288,N_34677);
nand U35124 (N_35124,N_34657,N_34730);
or U35125 (N_35125,N_34915,N_34408);
nor U35126 (N_35126,N_34129,N_34867);
nand U35127 (N_35127,N_34045,N_34549);
nand U35128 (N_35128,N_34912,N_34893);
nand U35129 (N_35129,N_34501,N_34074);
and U35130 (N_35130,N_34774,N_34885);
nand U35131 (N_35131,N_34405,N_34528);
or U35132 (N_35132,N_34345,N_34310);
xnor U35133 (N_35133,N_34655,N_34836);
xnor U35134 (N_35134,N_34451,N_34264);
and U35135 (N_35135,N_34341,N_34425);
nand U35136 (N_35136,N_34165,N_34584);
and U35137 (N_35137,N_34135,N_34303);
nor U35138 (N_35138,N_34510,N_34538);
nor U35139 (N_35139,N_34126,N_34077);
xnor U35140 (N_35140,N_34576,N_34195);
and U35141 (N_35141,N_34293,N_34877);
xnor U35142 (N_35142,N_34673,N_34968);
nand U35143 (N_35143,N_34797,N_34988);
xnor U35144 (N_35144,N_34203,N_34374);
xnor U35145 (N_35145,N_34113,N_34534);
and U35146 (N_35146,N_34740,N_34562);
and U35147 (N_35147,N_34775,N_34866);
nor U35148 (N_35148,N_34896,N_34500);
and U35149 (N_35149,N_34899,N_34806);
and U35150 (N_35150,N_34981,N_34980);
or U35151 (N_35151,N_34383,N_34733);
nand U35152 (N_35152,N_34087,N_34174);
nand U35153 (N_35153,N_34650,N_34874);
xor U35154 (N_35154,N_34311,N_34817);
nand U35155 (N_35155,N_34010,N_34484);
nand U35156 (N_35156,N_34103,N_34055);
xor U35157 (N_35157,N_34287,N_34091);
nor U35158 (N_35158,N_34834,N_34544);
or U35159 (N_35159,N_34177,N_34353);
or U35160 (N_35160,N_34390,N_34082);
or U35161 (N_35161,N_34594,N_34643);
nor U35162 (N_35162,N_34215,N_34618);
or U35163 (N_35163,N_34747,N_34134);
nor U35164 (N_35164,N_34100,N_34773);
and U35165 (N_35165,N_34585,N_34639);
and U35166 (N_35166,N_34319,N_34638);
or U35167 (N_35167,N_34377,N_34527);
nor U35168 (N_35168,N_34953,N_34602);
nand U35169 (N_35169,N_34127,N_34855);
and U35170 (N_35170,N_34582,N_34503);
nor U35171 (N_35171,N_34239,N_34508);
and U35172 (N_35172,N_34161,N_34133);
nand U35173 (N_35173,N_34487,N_34779);
and U35174 (N_35174,N_34363,N_34697);
or U35175 (N_35175,N_34958,N_34805);
or U35176 (N_35176,N_34492,N_34802);
xor U35177 (N_35177,N_34062,N_34758);
and U35178 (N_35178,N_34928,N_34013);
nand U35179 (N_35179,N_34785,N_34902);
or U35180 (N_35180,N_34827,N_34230);
and U35181 (N_35181,N_34943,N_34609);
or U35182 (N_35182,N_34710,N_34060);
and U35183 (N_35183,N_34176,N_34211);
or U35184 (N_35184,N_34309,N_34494);
xor U35185 (N_35185,N_34900,N_34612);
xnor U35186 (N_35186,N_34036,N_34856);
and U35187 (N_35187,N_34929,N_34704);
nand U35188 (N_35188,N_34477,N_34421);
nor U35189 (N_35189,N_34997,N_34107);
nor U35190 (N_35190,N_34903,N_34924);
and U35191 (N_35191,N_34999,N_34156);
nand U35192 (N_35192,N_34726,N_34897);
nor U35193 (N_35193,N_34986,N_34973);
xor U35194 (N_35194,N_34894,N_34063);
nand U35195 (N_35195,N_34241,N_34543);
or U35196 (N_35196,N_34920,N_34996);
and U35197 (N_35197,N_34409,N_34106);
and U35198 (N_35198,N_34627,N_34949);
nand U35199 (N_35199,N_34009,N_34031);
xnor U35200 (N_35200,N_34671,N_34210);
xnor U35201 (N_35201,N_34570,N_34387);
and U35202 (N_35202,N_34800,N_34168);
nor U35203 (N_35203,N_34942,N_34187);
nor U35204 (N_35204,N_34362,N_34250);
xnor U35205 (N_35205,N_34863,N_34646);
nor U35206 (N_35206,N_34453,N_34424);
nor U35207 (N_35207,N_34071,N_34216);
nor U35208 (N_35208,N_34829,N_34711);
nor U35209 (N_35209,N_34607,N_34962);
nor U35210 (N_35210,N_34839,N_34936);
or U35211 (N_35211,N_34025,N_34615);
nor U35212 (N_35212,N_34276,N_34222);
nand U35213 (N_35213,N_34085,N_34120);
and U35214 (N_35214,N_34645,N_34830);
nand U35215 (N_35215,N_34990,N_34696);
and U35216 (N_35216,N_34322,N_34038);
nor U35217 (N_35217,N_34058,N_34614);
xnor U35218 (N_35218,N_34604,N_34729);
xor U35219 (N_35219,N_34155,N_34340);
and U35220 (N_35220,N_34396,N_34097);
xor U35221 (N_35221,N_34233,N_34610);
xor U35222 (N_35222,N_34019,N_34852);
or U35223 (N_35223,N_34757,N_34298);
or U35224 (N_35224,N_34066,N_34660);
nor U35225 (N_35225,N_34551,N_34819);
and U35226 (N_35226,N_34600,N_34845);
nand U35227 (N_35227,N_34853,N_34667);
and U35228 (N_35228,N_34183,N_34820);
nand U35229 (N_35229,N_34145,N_34967);
or U35230 (N_35230,N_34748,N_34373);
and U35231 (N_35231,N_34395,N_34972);
and U35232 (N_35232,N_34190,N_34434);
or U35233 (N_35233,N_34854,N_34872);
nand U35234 (N_35234,N_34301,N_34540);
xnor U35235 (N_35235,N_34725,N_34302);
and U35236 (N_35236,N_34364,N_34532);
nand U35237 (N_35237,N_34745,N_34560);
xnor U35238 (N_35238,N_34039,N_34116);
nand U35239 (N_35239,N_34795,N_34932);
or U35240 (N_35240,N_34465,N_34559);
or U35241 (N_35241,N_34382,N_34948);
or U35242 (N_35242,N_34959,N_34531);
or U35243 (N_35243,N_34297,N_34720);
nor U35244 (N_35244,N_34124,N_34350);
nor U35245 (N_35245,N_34925,N_34482);
xnor U35246 (N_35246,N_34235,N_34960);
xnor U35247 (N_35247,N_34537,N_34567);
and U35248 (N_35248,N_34043,N_34469);
xnor U35249 (N_35249,N_34781,N_34270);
or U35250 (N_35250,N_34992,N_34206);
or U35251 (N_35251,N_34246,N_34040);
and U35252 (N_35252,N_34790,N_34664);
nand U35253 (N_35253,N_34712,N_34068);
or U35254 (N_35254,N_34033,N_34335);
and U35255 (N_35255,N_34148,N_34574);
and U35256 (N_35256,N_34067,N_34227);
or U35257 (N_35257,N_34881,N_34911);
xnor U35258 (N_35258,N_34229,N_34426);
or U35259 (N_35259,N_34761,N_34273);
nand U35260 (N_35260,N_34763,N_34857);
or U35261 (N_35261,N_34220,N_34890);
nor U35262 (N_35262,N_34111,N_34056);
nand U35263 (N_35263,N_34398,N_34518);
or U35264 (N_35264,N_34130,N_34024);
or U35265 (N_35265,N_34262,N_34792);
and U35266 (N_35266,N_34723,N_34054);
nor U35267 (N_35267,N_34381,N_34630);
or U35268 (N_35268,N_34007,N_34691);
nor U35269 (N_35269,N_34613,N_34483);
nand U35270 (N_35270,N_34261,N_34002);
or U35271 (N_35271,N_34780,N_34226);
nor U35272 (N_35272,N_34718,N_34916);
xor U35273 (N_35273,N_34053,N_34255);
or U35274 (N_35274,N_34695,N_34680);
and U35275 (N_35275,N_34075,N_34247);
or U35276 (N_35276,N_34096,N_34221);
and U35277 (N_35277,N_34523,N_34244);
xor U35278 (N_35278,N_34331,N_34349);
xor U35279 (N_35279,N_34304,N_34011);
nand U35280 (N_35280,N_34811,N_34887);
xnor U35281 (N_35281,N_34181,N_34020);
xnor U35282 (N_35282,N_34906,N_34006);
xnor U35283 (N_35283,N_34326,N_34536);
and U35284 (N_35284,N_34232,N_34835);
xor U35285 (N_35285,N_34589,N_34513);
xnor U35286 (N_35286,N_34674,N_34577);
and U35287 (N_35287,N_34571,N_34563);
nor U35288 (N_35288,N_34330,N_34368);
or U35289 (N_35289,N_34608,N_34277);
xnor U35290 (N_35290,N_34078,N_34017);
and U35291 (N_35291,N_34200,N_34821);
nand U35292 (N_35292,N_34050,N_34459);
xor U35293 (N_35293,N_34901,N_34282);
xor U35294 (N_35294,N_34289,N_34678);
xnor U35295 (N_35295,N_34568,N_34511);
and U35296 (N_35296,N_34514,N_34644);
nor U35297 (N_35297,N_34749,N_34825);
xor U35298 (N_35298,N_34504,N_34198);
xor U35299 (N_35299,N_34003,N_34080);
nor U35300 (N_35300,N_34769,N_34150);
and U35301 (N_35301,N_34572,N_34149);
nand U35302 (N_35302,N_34338,N_34648);
nor U35303 (N_35303,N_34370,N_34705);
and U35304 (N_35304,N_34692,N_34404);
nand U35305 (N_35305,N_34417,N_34946);
nor U35306 (N_35306,N_34883,N_34460);
xnor U35307 (N_35307,N_34375,N_34651);
nand U35308 (N_35308,N_34193,N_34832);
xnor U35309 (N_35309,N_34052,N_34888);
or U35310 (N_35310,N_34957,N_34858);
and U35311 (N_35311,N_34550,N_34379);
or U35312 (N_35312,N_34965,N_34892);
nand U35313 (N_35313,N_34119,N_34641);
and U35314 (N_35314,N_34212,N_34473);
xor U35315 (N_35315,N_34468,N_34698);
xnor U35316 (N_35316,N_34635,N_34598);
nor U35317 (N_35317,N_34784,N_34524);
xor U35318 (N_35318,N_34123,N_34624);
or U35319 (N_35319,N_34505,N_34401);
and U35320 (N_35320,N_34556,N_34407);
nand U35321 (N_35321,N_34329,N_34098);
xnor U35322 (N_35322,N_34141,N_34209);
nor U35323 (N_35323,N_34860,N_34512);
nor U35324 (N_35324,N_34517,N_34428);
nor U35325 (N_35325,N_34076,N_34826);
and U35326 (N_35326,N_34343,N_34634);
and U35327 (N_35327,N_34266,N_34831);
nor U35328 (N_35328,N_34385,N_34931);
and U35329 (N_35329,N_34356,N_34258);
nand U35330 (N_35330,N_34333,N_34727);
nor U35331 (N_35331,N_34993,N_34913);
and U35332 (N_35332,N_34891,N_34272);
nor U35333 (N_35333,N_34926,N_34579);
and U35334 (N_35334,N_34471,N_34292);
nand U35335 (N_35335,N_34372,N_34138);
xnor U35336 (N_35336,N_34956,N_34647);
xnor U35337 (N_35337,N_34496,N_34047);
or U35338 (N_35338,N_34869,N_34547);
and U35339 (N_35339,N_34525,N_34416);
nor U35340 (N_35340,N_34016,N_34770);
or U35341 (N_35341,N_34809,N_34476);
xor U35342 (N_35342,N_34688,N_34065);
nor U35343 (N_35343,N_34756,N_34793);
nand U35344 (N_35344,N_34597,N_34789);
xor U35345 (N_35345,N_34905,N_34391);
nor U35346 (N_35346,N_34173,N_34406);
nand U35347 (N_35347,N_34073,N_34035);
or U35348 (N_35348,N_34281,N_34768);
nand U35349 (N_35349,N_34882,N_34104);
xor U35350 (N_35350,N_34904,N_34204);
nand U35351 (N_35351,N_34945,N_34088);
nand U35352 (N_35352,N_34859,N_34681);
or U35353 (N_35353,N_34669,N_34838);
or U35354 (N_35354,N_34015,N_34475);
nand U35355 (N_35355,N_34327,N_34084);
and U35356 (N_35356,N_34984,N_34861);
and U35357 (N_35357,N_34760,N_34397);
nor U35358 (N_35358,N_34526,N_34466);
xor U35359 (N_35359,N_34411,N_34810);
or U35360 (N_35360,N_34099,N_34693);
nor U35361 (N_35361,N_34030,N_34415);
and U35362 (N_35362,N_34927,N_34690);
xnor U35363 (N_35363,N_34998,N_34786);
nor U35364 (N_35364,N_34185,N_34018);
xor U35365 (N_35365,N_34782,N_34225);
nor U35366 (N_35366,N_34291,N_34263);
nor U35367 (N_35367,N_34884,N_34394);
and U35368 (N_35368,N_34516,N_34422);
nand U35369 (N_35369,N_34601,N_34519);
nand U35370 (N_35370,N_34259,N_34961);
and U35371 (N_35371,N_34694,N_34245);
nor U35372 (N_35372,N_34184,N_34799);
nand U35373 (N_35373,N_34824,N_34178);
nand U35374 (N_35374,N_34441,N_34224);
or U35375 (N_35375,N_34159,N_34935);
nor U35376 (N_35376,N_34342,N_34636);
xnor U35377 (N_35377,N_34026,N_34849);
nand U35378 (N_35378,N_34499,N_34764);
nor U35379 (N_35379,N_34307,N_34347);
nand U35380 (N_35380,N_34548,N_34808);
and U35381 (N_35381,N_34914,N_34427);
nor U35382 (N_35382,N_34290,N_34253);
nand U35383 (N_35383,N_34367,N_34132);
and U35384 (N_35384,N_34445,N_34139);
and U35385 (N_35385,N_34828,N_34294);
and U35386 (N_35386,N_34777,N_34606);
nand U35387 (N_35387,N_34846,N_34136);
nor U35388 (N_35388,N_34143,N_34359);
xor U35389 (N_35389,N_34412,N_34895);
nor U35390 (N_35390,N_34898,N_34137);
xor U35391 (N_35391,N_34495,N_34752);
nor U35392 (N_35392,N_34778,N_34205);
nor U35393 (N_35393,N_34841,N_34489);
nor U35394 (N_35394,N_34430,N_34472);
nor U35395 (N_35395,N_34675,N_34670);
and U35396 (N_35396,N_34917,N_34446);
nor U35397 (N_35397,N_34022,N_34154);
or U35398 (N_35398,N_34001,N_34070);
xor U35399 (N_35399,N_34151,N_34656);
nor U35400 (N_35400,N_34684,N_34208);
xnor U35401 (N_35401,N_34642,N_34801);
nand U35402 (N_35402,N_34012,N_34850);
or U35403 (N_35403,N_34236,N_34595);
nand U35404 (N_35404,N_34788,N_34299);
nand U35405 (N_35405,N_34274,N_34794);
and U35406 (N_35406,N_34663,N_34930);
nor U35407 (N_35407,N_34448,N_34619);
and U35408 (N_35408,N_34464,N_34454);
or U35409 (N_35409,N_34179,N_34443);
and U35410 (N_35410,N_34623,N_34701);
xor U35411 (N_35411,N_34676,N_34231);
nand U35412 (N_35412,N_34046,N_34566);
or U35413 (N_35413,N_34728,N_34452);
nor U35414 (N_35414,N_34593,N_34611);
nor U35415 (N_35415,N_34969,N_34975);
and U35416 (N_35416,N_34146,N_34545);
xnor U35417 (N_35417,N_34746,N_34919);
or U35418 (N_35418,N_34783,N_34042);
or U35419 (N_35419,N_34160,N_34023);
xnor U35420 (N_35420,N_34217,N_34388);
xor U35421 (N_35421,N_34991,N_34502);
nand U35422 (N_35422,N_34498,N_34435);
nand U35423 (N_35423,N_34481,N_34214);
nand U35424 (N_35424,N_34295,N_34766);
nand U35425 (N_35425,N_34196,N_34759);
and U35426 (N_35426,N_34561,N_34081);
xor U35427 (N_35427,N_34251,N_34631);
nor U35428 (N_35428,N_34816,N_34355);
nor U35429 (N_35429,N_34699,N_34167);
and U35430 (N_35430,N_34431,N_34089);
and U35431 (N_35431,N_34142,N_34480);
and U35432 (N_35432,N_34719,N_34909);
xnor U35433 (N_35433,N_34197,N_34207);
or U35434 (N_35434,N_34284,N_34734);
and U35435 (N_35435,N_34083,N_34837);
nor U35436 (N_35436,N_34716,N_34952);
xnor U35437 (N_35437,N_34581,N_34622);
nor U35438 (N_35438,N_34554,N_34940);
nor U35439 (N_35439,N_34108,N_34833);
nor U35440 (N_35440,N_34414,N_34041);
and U35441 (N_35441,N_34731,N_34851);
and U35442 (N_35442,N_34682,N_34842);
nor U35443 (N_35443,N_34649,N_34951);
and U35444 (N_35444,N_34542,N_34271);
and U35445 (N_35445,N_34449,N_34873);
xor U35446 (N_35446,N_34771,N_34131);
or U35447 (N_35447,N_34094,N_34616);
xnor U35448 (N_35448,N_34938,N_34458);
and U35449 (N_35449,N_34557,N_34238);
nor U35450 (N_35450,N_34110,N_34429);
and U35451 (N_35451,N_34102,N_34280);
or U35452 (N_35452,N_34175,N_34186);
or U35453 (N_35453,N_34840,N_34687);
and U35454 (N_35454,N_34989,N_34470);
or U35455 (N_35455,N_34064,N_34069);
and U35456 (N_35456,N_34467,N_34393);
nor U35457 (N_35457,N_34218,N_34985);
nand U35458 (N_35458,N_34707,N_34144);
nand U35459 (N_35459,N_34633,N_34418);
nand U35460 (N_35460,N_34313,N_34337);
nand U35461 (N_35461,N_34907,N_34202);
nand U35462 (N_35462,N_34308,N_34491);
and U35463 (N_35463,N_34278,N_34439);
nand U35464 (N_35464,N_34172,N_34722);
or U35465 (N_35465,N_34191,N_34910);
nor U35466 (N_35466,N_34583,N_34463);
and U35467 (N_35467,N_34219,N_34044);
nor U35468 (N_35468,N_34520,N_34392);
xnor U35469 (N_35469,N_34410,N_34318);
nand U35470 (N_35470,N_34923,N_34605);
nor U35471 (N_35471,N_34818,N_34346);
nand U35472 (N_35472,N_34937,N_34870);
or U35473 (N_35473,N_34515,N_34432);
nand U35474 (N_35474,N_34735,N_34157);
nor U35475 (N_35475,N_34591,N_34522);
and U35476 (N_35476,N_34188,N_34588);
nor U35477 (N_35477,N_34140,N_34049);
nor U35478 (N_35478,N_34314,N_34848);
nand U35479 (N_35479,N_34109,N_34823);
or U35480 (N_35480,N_34357,N_34535);
nor U35481 (N_35481,N_34455,N_34339);
nor U35482 (N_35482,N_34112,N_34918);
nand U35483 (N_35483,N_34447,N_34105);
nor U35484 (N_35484,N_34114,N_34521);
nor U35485 (N_35485,N_34744,N_34121);
and U35486 (N_35486,N_34762,N_34240);
nand U35487 (N_35487,N_34371,N_34666);
or U35488 (N_35488,N_34242,N_34876);
or U35489 (N_35489,N_34578,N_34555);
and U35490 (N_35490,N_34315,N_34440);
nand U35491 (N_35491,N_34950,N_34254);
nand U35492 (N_35492,N_34679,N_34767);
and U35493 (N_35493,N_34738,N_34878);
nand U35494 (N_35494,N_34248,N_34336);
or U35495 (N_35495,N_34683,N_34739);
nor U35496 (N_35496,N_34057,N_34880);
nor U35497 (N_35497,N_34750,N_34603);
xnor U35498 (N_35498,N_34724,N_34008);
xnor U35499 (N_35499,N_34051,N_34803);
nand U35500 (N_35500,N_34840,N_34926);
or U35501 (N_35501,N_34340,N_34707);
and U35502 (N_35502,N_34154,N_34643);
and U35503 (N_35503,N_34020,N_34725);
xor U35504 (N_35504,N_34334,N_34947);
xnor U35505 (N_35505,N_34398,N_34065);
and U35506 (N_35506,N_34124,N_34899);
xor U35507 (N_35507,N_34809,N_34274);
or U35508 (N_35508,N_34891,N_34409);
and U35509 (N_35509,N_34212,N_34302);
and U35510 (N_35510,N_34585,N_34097);
or U35511 (N_35511,N_34795,N_34231);
nor U35512 (N_35512,N_34214,N_34397);
and U35513 (N_35513,N_34280,N_34967);
and U35514 (N_35514,N_34901,N_34245);
or U35515 (N_35515,N_34715,N_34494);
nand U35516 (N_35516,N_34982,N_34890);
xor U35517 (N_35517,N_34031,N_34318);
nor U35518 (N_35518,N_34300,N_34668);
nor U35519 (N_35519,N_34524,N_34739);
or U35520 (N_35520,N_34036,N_34677);
nand U35521 (N_35521,N_34749,N_34802);
xor U35522 (N_35522,N_34927,N_34194);
and U35523 (N_35523,N_34740,N_34210);
and U35524 (N_35524,N_34994,N_34250);
or U35525 (N_35525,N_34359,N_34182);
and U35526 (N_35526,N_34513,N_34816);
and U35527 (N_35527,N_34456,N_34561);
or U35528 (N_35528,N_34467,N_34531);
xnor U35529 (N_35529,N_34424,N_34397);
nor U35530 (N_35530,N_34384,N_34672);
nor U35531 (N_35531,N_34854,N_34408);
xor U35532 (N_35532,N_34555,N_34548);
nand U35533 (N_35533,N_34928,N_34343);
and U35534 (N_35534,N_34246,N_34458);
xnor U35535 (N_35535,N_34363,N_34325);
and U35536 (N_35536,N_34520,N_34397);
or U35537 (N_35537,N_34333,N_34777);
nor U35538 (N_35538,N_34857,N_34491);
nor U35539 (N_35539,N_34364,N_34536);
nand U35540 (N_35540,N_34238,N_34943);
or U35541 (N_35541,N_34263,N_34236);
xor U35542 (N_35542,N_34164,N_34975);
nor U35543 (N_35543,N_34491,N_34871);
and U35544 (N_35544,N_34625,N_34462);
or U35545 (N_35545,N_34750,N_34930);
nand U35546 (N_35546,N_34154,N_34607);
nand U35547 (N_35547,N_34505,N_34301);
xnor U35548 (N_35548,N_34840,N_34370);
xor U35549 (N_35549,N_34974,N_34811);
or U35550 (N_35550,N_34520,N_34752);
or U35551 (N_35551,N_34429,N_34104);
nand U35552 (N_35552,N_34075,N_34618);
or U35553 (N_35553,N_34963,N_34105);
or U35554 (N_35554,N_34359,N_34620);
or U35555 (N_35555,N_34373,N_34755);
nor U35556 (N_35556,N_34140,N_34597);
xor U35557 (N_35557,N_34455,N_34228);
nor U35558 (N_35558,N_34902,N_34024);
and U35559 (N_35559,N_34815,N_34085);
or U35560 (N_35560,N_34244,N_34664);
xnor U35561 (N_35561,N_34487,N_34213);
and U35562 (N_35562,N_34359,N_34193);
nand U35563 (N_35563,N_34932,N_34397);
xnor U35564 (N_35564,N_34336,N_34193);
nor U35565 (N_35565,N_34467,N_34562);
xor U35566 (N_35566,N_34020,N_34272);
nor U35567 (N_35567,N_34064,N_34346);
and U35568 (N_35568,N_34899,N_34639);
nor U35569 (N_35569,N_34419,N_34067);
nand U35570 (N_35570,N_34369,N_34865);
xnor U35571 (N_35571,N_34468,N_34253);
and U35572 (N_35572,N_34545,N_34687);
or U35573 (N_35573,N_34260,N_34387);
xor U35574 (N_35574,N_34681,N_34385);
nor U35575 (N_35575,N_34204,N_34793);
or U35576 (N_35576,N_34186,N_34634);
nor U35577 (N_35577,N_34020,N_34976);
xnor U35578 (N_35578,N_34210,N_34715);
nand U35579 (N_35579,N_34216,N_34170);
nand U35580 (N_35580,N_34096,N_34142);
or U35581 (N_35581,N_34739,N_34161);
nand U35582 (N_35582,N_34906,N_34783);
nor U35583 (N_35583,N_34940,N_34262);
and U35584 (N_35584,N_34188,N_34145);
nor U35585 (N_35585,N_34618,N_34360);
and U35586 (N_35586,N_34281,N_34806);
nand U35587 (N_35587,N_34532,N_34061);
and U35588 (N_35588,N_34332,N_34884);
nand U35589 (N_35589,N_34904,N_34378);
nor U35590 (N_35590,N_34511,N_34554);
xnor U35591 (N_35591,N_34789,N_34115);
nand U35592 (N_35592,N_34747,N_34997);
nand U35593 (N_35593,N_34302,N_34317);
or U35594 (N_35594,N_34351,N_34336);
xnor U35595 (N_35595,N_34456,N_34391);
nand U35596 (N_35596,N_34020,N_34756);
nor U35597 (N_35597,N_34147,N_34468);
nand U35598 (N_35598,N_34718,N_34229);
or U35599 (N_35599,N_34536,N_34565);
nand U35600 (N_35600,N_34196,N_34474);
xnor U35601 (N_35601,N_34013,N_34456);
and U35602 (N_35602,N_34686,N_34854);
nand U35603 (N_35603,N_34687,N_34571);
nor U35604 (N_35604,N_34054,N_34539);
xor U35605 (N_35605,N_34261,N_34742);
nor U35606 (N_35606,N_34150,N_34313);
and U35607 (N_35607,N_34976,N_34533);
xnor U35608 (N_35608,N_34237,N_34486);
nor U35609 (N_35609,N_34698,N_34133);
nor U35610 (N_35610,N_34308,N_34772);
xor U35611 (N_35611,N_34594,N_34765);
nor U35612 (N_35612,N_34542,N_34349);
xor U35613 (N_35613,N_34757,N_34964);
or U35614 (N_35614,N_34025,N_34495);
and U35615 (N_35615,N_34859,N_34235);
nand U35616 (N_35616,N_34378,N_34555);
and U35617 (N_35617,N_34677,N_34398);
nand U35618 (N_35618,N_34477,N_34218);
xor U35619 (N_35619,N_34093,N_34380);
xnor U35620 (N_35620,N_34517,N_34765);
nand U35621 (N_35621,N_34793,N_34028);
or U35622 (N_35622,N_34999,N_34896);
nor U35623 (N_35623,N_34618,N_34946);
or U35624 (N_35624,N_34871,N_34456);
nor U35625 (N_35625,N_34354,N_34912);
xnor U35626 (N_35626,N_34703,N_34762);
xor U35627 (N_35627,N_34796,N_34496);
xnor U35628 (N_35628,N_34588,N_34515);
and U35629 (N_35629,N_34778,N_34615);
xnor U35630 (N_35630,N_34268,N_34609);
xor U35631 (N_35631,N_34516,N_34550);
or U35632 (N_35632,N_34036,N_34506);
and U35633 (N_35633,N_34583,N_34447);
nand U35634 (N_35634,N_34639,N_34375);
nand U35635 (N_35635,N_34930,N_34060);
nand U35636 (N_35636,N_34578,N_34199);
nand U35637 (N_35637,N_34094,N_34016);
or U35638 (N_35638,N_34591,N_34726);
or U35639 (N_35639,N_34590,N_34224);
nand U35640 (N_35640,N_34216,N_34020);
nand U35641 (N_35641,N_34598,N_34676);
nand U35642 (N_35642,N_34674,N_34475);
xor U35643 (N_35643,N_34200,N_34651);
or U35644 (N_35644,N_34382,N_34349);
or U35645 (N_35645,N_34250,N_34324);
and U35646 (N_35646,N_34595,N_34903);
and U35647 (N_35647,N_34670,N_34492);
xnor U35648 (N_35648,N_34518,N_34151);
xnor U35649 (N_35649,N_34305,N_34014);
nand U35650 (N_35650,N_34718,N_34944);
nand U35651 (N_35651,N_34385,N_34271);
and U35652 (N_35652,N_34161,N_34253);
nor U35653 (N_35653,N_34755,N_34008);
nor U35654 (N_35654,N_34675,N_34055);
nor U35655 (N_35655,N_34881,N_34571);
and U35656 (N_35656,N_34683,N_34060);
and U35657 (N_35657,N_34463,N_34116);
and U35658 (N_35658,N_34228,N_34803);
nand U35659 (N_35659,N_34458,N_34696);
nor U35660 (N_35660,N_34524,N_34513);
and U35661 (N_35661,N_34289,N_34009);
or U35662 (N_35662,N_34311,N_34081);
or U35663 (N_35663,N_34471,N_34558);
and U35664 (N_35664,N_34426,N_34785);
nor U35665 (N_35665,N_34563,N_34884);
and U35666 (N_35666,N_34926,N_34501);
and U35667 (N_35667,N_34725,N_34756);
or U35668 (N_35668,N_34070,N_34390);
nor U35669 (N_35669,N_34675,N_34500);
nor U35670 (N_35670,N_34863,N_34054);
nor U35671 (N_35671,N_34649,N_34947);
and U35672 (N_35672,N_34125,N_34691);
nor U35673 (N_35673,N_34960,N_34664);
and U35674 (N_35674,N_34973,N_34712);
and U35675 (N_35675,N_34386,N_34528);
or U35676 (N_35676,N_34701,N_34866);
or U35677 (N_35677,N_34950,N_34412);
and U35678 (N_35678,N_34496,N_34452);
xnor U35679 (N_35679,N_34465,N_34852);
xnor U35680 (N_35680,N_34711,N_34388);
nor U35681 (N_35681,N_34266,N_34543);
or U35682 (N_35682,N_34973,N_34519);
xor U35683 (N_35683,N_34892,N_34692);
and U35684 (N_35684,N_34874,N_34581);
nand U35685 (N_35685,N_34477,N_34027);
and U35686 (N_35686,N_34608,N_34611);
nor U35687 (N_35687,N_34914,N_34129);
or U35688 (N_35688,N_34768,N_34689);
or U35689 (N_35689,N_34130,N_34309);
xnor U35690 (N_35690,N_34684,N_34204);
xor U35691 (N_35691,N_34213,N_34416);
nand U35692 (N_35692,N_34149,N_34084);
xor U35693 (N_35693,N_34465,N_34706);
nor U35694 (N_35694,N_34197,N_34537);
nor U35695 (N_35695,N_34357,N_34402);
and U35696 (N_35696,N_34375,N_34927);
xnor U35697 (N_35697,N_34214,N_34511);
xnor U35698 (N_35698,N_34512,N_34010);
or U35699 (N_35699,N_34800,N_34437);
and U35700 (N_35700,N_34942,N_34721);
and U35701 (N_35701,N_34096,N_34800);
or U35702 (N_35702,N_34286,N_34729);
nor U35703 (N_35703,N_34456,N_34769);
and U35704 (N_35704,N_34908,N_34530);
xnor U35705 (N_35705,N_34429,N_34068);
nor U35706 (N_35706,N_34459,N_34700);
and U35707 (N_35707,N_34135,N_34326);
or U35708 (N_35708,N_34324,N_34699);
and U35709 (N_35709,N_34253,N_34457);
nand U35710 (N_35710,N_34826,N_34238);
and U35711 (N_35711,N_34351,N_34452);
xor U35712 (N_35712,N_34538,N_34478);
and U35713 (N_35713,N_34403,N_34110);
xnor U35714 (N_35714,N_34276,N_34107);
xor U35715 (N_35715,N_34848,N_34056);
xor U35716 (N_35716,N_34486,N_34927);
nor U35717 (N_35717,N_34806,N_34880);
xor U35718 (N_35718,N_34195,N_34133);
xor U35719 (N_35719,N_34843,N_34976);
and U35720 (N_35720,N_34058,N_34379);
nor U35721 (N_35721,N_34885,N_34248);
nor U35722 (N_35722,N_34895,N_34592);
or U35723 (N_35723,N_34393,N_34966);
nor U35724 (N_35724,N_34200,N_34246);
or U35725 (N_35725,N_34481,N_34867);
nor U35726 (N_35726,N_34760,N_34641);
xor U35727 (N_35727,N_34203,N_34837);
or U35728 (N_35728,N_34584,N_34548);
or U35729 (N_35729,N_34852,N_34420);
nand U35730 (N_35730,N_34752,N_34128);
nor U35731 (N_35731,N_34066,N_34897);
nand U35732 (N_35732,N_34857,N_34721);
or U35733 (N_35733,N_34417,N_34233);
or U35734 (N_35734,N_34086,N_34799);
or U35735 (N_35735,N_34204,N_34063);
or U35736 (N_35736,N_34645,N_34868);
and U35737 (N_35737,N_34907,N_34680);
nand U35738 (N_35738,N_34178,N_34987);
and U35739 (N_35739,N_34813,N_34682);
xor U35740 (N_35740,N_34701,N_34004);
nand U35741 (N_35741,N_34939,N_34325);
xnor U35742 (N_35742,N_34129,N_34563);
nand U35743 (N_35743,N_34794,N_34272);
or U35744 (N_35744,N_34306,N_34262);
nand U35745 (N_35745,N_34500,N_34991);
nor U35746 (N_35746,N_34827,N_34321);
and U35747 (N_35747,N_34479,N_34080);
nand U35748 (N_35748,N_34857,N_34945);
xnor U35749 (N_35749,N_34475,N_34210);
nor U35750 (N_35750,N_34982,N_34007);
or U35751 (N_35751,N_34306,N_34132);
or U35752 (N_35752,N_34348,N_34061);
or U35753 (N_35753,N_34330,N_34925);
and U35754 (N_35754,N_34453,N_34730);
nor U35755 (N_35755,N_34850,N_34515);
or U35756 (N_35756,N_34316,N_34280);
nor U35757 (N_35757,N_34801,N_34117);
and U35758 (N_35758,N_34799,N_34521);
nor U35759 (N_35759,N_34164,N_34006);
and U35760 (N_35760,N_34998,N_34147);
nor U35761 (N_35761,N_34604,N_34503);
xnor U35762 (N_35762,N_34106,N_34342);
xor U35763 (N_35763,N_34917,N_34038);
xnor U35764 (N_35764,N_34806,N_34975);
xnor U35765 (N_35765,N_34836,N_34498);
xor U35766 (N_35766,N_34361,N_34966);
and U35767 (N_35767,N_34764,N_34046);
nor U35768 (N_35768,N_34420,N_34464);
and U35769 (N_35769,N_34451,N_34958);
and U35770 (N_35770,N_34832,N_34144);
or U35771 (N_35771,N_34271,N_34746);
nand U35772 (N_35772,N_34354,N_34531);
and U35773 (N_35773,N_34580,N_34358);
xor U35774 (N_35774,N_34610,N_34429);
and U35775 (N_35775,N_34536,N_34928);
nand U35776 (N_35776,N_34136,N_34084);
nor U35777 (N_35777,N_34771,N_34510);
or U35778 (N_35778,N_34749,N_34741);
and U35779 (N_35779,N_34030,N_34688);
and U35780 (N_35780,N_34429,N_34836);
xor U35781 (N_35781,N_34091,N_34615);
and U35782 (N_35782,N_34088,N_34046);
xnor U35783 (N_35783,N_34979,N_34425);
nand U35784 (N_35784,N_34027,N_34776);
nor U35785 (N_35785,N_34657,N_34680);
or U35786 (N_35786,N_34263,N_34025);
nor U35787 (N_35787,N_34043,N_34607);
xor U35788 (N_35788,N_34685,N_34460);
nor U35789 (N_35789,N_34122,N_34303);
or U35790 (N_35790,N_34243,N_34780);
nor U35791 (N_35791,N_34905,N_34375);
and U35792 (N_35792,N_34395,N_34635);
xor U35793 (N_35793,N_34465,N_34177);
nor U35794 (N_35794,N_34245,N_34073);
xor U35795 (N_35795,N_34727,N_34480);
nor U35796 (N_35796,N_34984,N_34765);
and U35797 (N_35797,N_34892,N_34390);
nand U35798 (N_35798,N_34367,N_34745);
xor U35799 (N_35799,N_34921,N_34051);
and U35800 (N_35800,N_34785,N_34068);
and U35801 (N_35801,N_34079,N_34220);
nor U35802 (N_35802,N_34781,N_34231);
and U35803 (N_35803,N_34723,N_34394);
nor U35804 (N_35804,N_34854,N_34066);
or U35805 (N_35805,N_34461,N_34934);
nand U35806 (N_35806,N_34214,N_34058);
and U35807 (N_35807,N_34105,N_34031);
or U35808 (N_35808,N_34121,N_34272);
and U35809 (N_35809,N_34489,N_34963);
and U35810 (N_35810,N_34414,N_34030);
or U35811 (N_35811,N_34232,N_34849);
nor U35812 (N_35812,N_34573,N_34661);
and U35813 (N_35813,N_34636,N_34929);
or U35814 (N_35814,N_34610,N_34384);
nand U35815 (N_35815,N_34417,N_34296);
and U35816 (N_35816,N_34062,N_34934);
and U35817 (N_35817,N_34564,N_34902);
or U35818 (N_35818,N_34083,N_34902);
or U35819 (N_35819,N_34103,N_34174);
xor U35820 (N_35820,N_34927,N_34730);
and U35821 (N_35821,N_34132,N_34438);
and U35822 (N_35822,N_34657,N_34796);
or U35823 (N_35823,N_34605,N_34631);
nor U35824 (N_35824,N_34414,N_34140);
nand U35825 (N_35825,N_34534,N_34439);
xor U35826 (N_35826,N_34331,N_34266);
and U35827 (N_35827,N_34262,N_34983);
nand U35828 (N_35828,N_34697,N_34980);
nor U35829 (N_35829,N_34257,N_34860);
xor U35830 (N_35830,N_34614,N_34350);
nor U35831 (N_35831,N_34277,N_34713);
and U35832 (N_35832,N_34202,N_34379);
nand U35833 (N_35833,N_34430,N_34848);
xor U35834 (N_35834,N_34331,N_34626);
or U35835 (N_35835,N_34167,N_34673);
xor U35836 (N_35836,N_34928,N_34820);
and U35837 (N_35837,N_34152,N_34334);
or U35838 (N_35838,N_34829,N_34592);
nand U35839 (N_35839,N_34894,N_34034);
xor U35840 (N_35840,N_34239,N_34443);
nor U35841 (N_35841,N_34756,N_34923);
and U35842 (N_35842,N_34815,N_34196);
and U35843 (N_35843,N_34648,N_34250);
and U35844 (N_35844,N_34053,N_34828);
and U35845 (N_35845,N_34412,N_34990);
and U35846 (N_35846,N_34659,N_34462);
or U35847 (N_35847,N_34514,N_34109);
and U35848 (N_35848,N_34548,N_34754);
or U35849 (N_35849,N_34397,N_34555);
xnor U35850 (N_35850,N_34038,N_34339);
nand U35851 (N_35851,N_34645,N_34120);
nand U35852 (N_35852,N_34889,N_34085);
xor U35853 (N_35853,N_34509,N_34674);
nor U35854 (N_35854,N_34409,N_34849);
xor U35855 (N_35855,N_34996,N_34156);
and U35856 (N_35856,N_34950,N_34803);
nor U35857 (N_35857,N_34428,N_34138);
xor U35858 (N_35858,N_34408,N_34538);
or U35859 (N_35859,N_34584,N_34115);
or U35860 (N_35860,N_34076,N_34283);
xnor U35861 (N_35861,N_34511,N_34004);
nand U35862 (N_35862,N_34744,N_34671);
nor U35863 (N_35863,N_34829,N_34150);
nor U35864 (N_35864,N_34705,N_34192);
xnor U35865 (N_35865,N_34099,N_34445);
and U35866 (N_35866,N_34813,N_34528);
xnor U35867 (N_35867,N_34410,N_34380);
or U35868 (N_35868,N_34299,N_34551);
xor U35869 (N_35869,N_34920,N_34070);
nand U35870 (N_35870,N_34752,N_34809);
nor U35871 (N_35871,N_34760,N_34616);
nor U35872 (N_35872,N_34690,N_34319);
nand U35873 (N_35873,N_34235,N_34182);
or U35874 (N_35874,N_34862,N_34423);
xor U35875 (N_35875,N_34955,N_34353);
and U35876 (N_35876,N_34323,N_34430);
xnor U35877 (N_35877,N_34030,N_34881);
and U35878 (N_35878,N_34263,N_34113);
or U35879 (N_35879,N_34714,N_34238);
or U35880 (N_35880,N_34181,N_34311);
nand U35881 (N_35881,N_34128,N_34486);
xnor U35882 (N_35882,N_34696,N_34944);
nor U35883 (N_35883,N_34633,N_34209);
and U35884 (N_35884,N_34455,N_34366);
nand U35885 (N_35885,N_34823,N_34224);
or U35886 (N_35886,N_34563,N_34449);
nor U35887 (N_35887,N_34784,N_34641);
and U35888 (N_35888,N_34697,N_34389);
nor U35889 (N_35889,N_34949,N_34372);
and U35890 (N_35890,N_34476,N_34301);
nor U35891 (N_35891,N_34320,N_34024);
or U35892 (N_35892,N_34153,N_34407);
nand U35893 (N_35893,N_34250,N_34002);
or U35894 (N_35894,N_34595,N_34533);
nand U35895 (N_35895,N_34866,N_34710);
nand U35896 (N_35896,N_34232,N_34006);
xor U35897 (N_35897,N_34157,N_34915);
nor U35898 (N_35898,N_34119,N_34829);
nor U35899 (N_35899,N_34154,N_34951);
and U35900 (N_35900,N_34362,N_34970);
and U35901 (N_35901,N_34343,N_34757);
nand U35902 (N_35902,N_34702,N_34710);
nor U35903 (N_35903,N_34141,N_34683);
nand U35904 (N_35904,N_34309,N_34387);
xnor U35905 (N_35905,N_34890,N_34762);
and U35906 (N_35906,N_34382,N_34175);
xor U35907 (N_35907,N_34840,N_34115);
or U35908 (N_35908,N_34388,N_34628);
nor U35909 (N_35909,N_34900,N_34058);
nand U35910 (N_35910,N_34209,N_34533);
nand U35911 (N_35911,N_34277,N_34629);
and U35912 (N_35912,N_34890,N_34172);
nand U35913 (N_35913,N_34071,N_34768);
or U35914 (N_35914,N_34838,N_34104);
nand U35915 (N_35915,N_34843,N_34772);
or U35916 (N_35916,N_34659,N_34658);
nand U35917 (N_35917,N_34037,N_34951);
nor U35918 (N_35918,N_34776,N_34377);
and U35919 (N_35919,N_34673,N_34488);
and U35920 (N_35920,N_34240,N_34772);
xnor U35921 (N_35921,N_34116,N_34314);
nand U35922 (N_35922,N_34208,N_34056);
or U35923 (N_35923,N_34221,N_34483);
and U35924 (N_35924,N_34275,N_34033);
or U35925 (N_35925,N_34243,N_34441);
or U35926 (N_35926,N_34808,N_34344);
and U35927 (N_35927,N_34099,N_34214);
or U35928 (N_35928,N_34216,N_34731);
and U35929 (N_35929,N_34639,N_34999);
and U35930 (N_35930,N_34927,N_34228);
or U35931 (N_35931,N_34823,N_34397);
and U35932 (N_35932,N_34107,N_34747);
and U35933 (N_35933,N_34455,N_34723);
nor U35934 (N_35934,N_34662,N_34862);
nand U35935 (N_35935,N_34875,N_34370);
nand U35936 (N_35936,N_34529,N_34285);
and U35937 (N_35937,N_34591,N_34018);
xor U35938 (N_35938,N_34808,N_34676);
nor U35939 (N_35939,N_34931,N_34340);
nand U35940 (N_35940,N_34356,N_34362);
and U35941 (N_35941,N_34547,N_34535);
nand U35942 (N_35942,N_34569,N_34134);
or U35943 (N_35943,N_34985,N_34340);
and U35944 (N_35944,N_34587,N_34332);
nor U35945 (N_35945,N_34790,N_34010);
or U35946 (N_35946,N_34805,N_34751);
nor U35947 (N_35947,N_34437,N_34835);
nand U35948 (N_35948,N_34133,N_34845);
xnor U35949 (N_35949,N_34131,N_34115);
or U35950 (N_35950,N_34400,N_34729);
nor U35951 (N_35951,N_34958,N_34653);
nor U35952 (N_35952,N_34692,N_34900);
or U35953 (N_35953,N_34917,N_34083);
xnor U35954 (N_35954,N_34118,N_34210);
nor U35955 (N_35955,N_34010,N_34553);
xnor U35956 (N_35956,N_34937,N_34072);
xor U35957 (N_35957,N_34664,N_34898);
nor U35958 (N_35958,N_34547,N_34266);
nor U35959 (N_35959,N_34961,N_34734);
xnor U35960 (N_35960,N_34041,N_34008);
and U35961 (N_35961,N_34113,N_34549);
and U35962 (N_35962,N_34447,N_34065);
nor U35963 (N_35963,N_34329,N_34725);
nor U35964 (N_35964,N_34802,N_34845);
nand U35965 (N_35965,N_34211,N_34015);
and U35966 (N_35966,N_34655,N_34670);
nand U35967 (N_35967,N_34611,N_34551);
nand U35968 (N_35968,N_34947,N_34506);
or U35969 (N_35969,N_34181,N_34540);
nand U35970 (N_35970,N_34148,N_34916);
nor U35971 (N_35971,N_34122,N_34253);
nand U35972 (N_35972,N_34824,N_34240);
nor U35973 (N_35973,N_34031,N_34195);
and U35974 (N_35974,N_34935,N_34340);
nor U35975 (N_35975,N_34345,N_34637);
xor U35976 (N_35976,N_34182,N_34422);
or U35977 (N_35977,N_34655,N_34889);
nand U35978 (N_35978,N_34136,N_34400);
nor U35979 (N_35979,N_34217,N_34247);
nand U35980 (N_35980,N_34147,N_34774);
xor U35981 (N_35981,N_34074,N_34963);
or U35982 (N_35982,N_34114,N_34940);
nor U35983 (N_35983,N_34769,N_34785);
nand U35984 (N_35984,N_34082,N_34991);
or U35985 (N_35985,N_34130,N_34909);
nand U35986 (N_35986,N_34444,N_34653);
xnor U35987 (N_35987,N_34073,N_34272);
or U35988 (N_35988,N_34834,N_34348);
and U35989 (N_35989,N_34577,N_34960);
xor U35990 (N_35990,N_34514,N_34264);
or U35991 (N_35991,N_34327,N_34318);
and U35992 (N_35992,N_34049,N_34096);
nor U35993 (N_35993,N_34557,N_34008);
nor U35994 (N_35994,N_34994,N_34701);
nor U35995 (N_35995,N_34726,N_34465);
xor U35996 (N_35996,N_34412,N_34479);
nor U35997 (N_35997,N_34116,N_34087);
or U35998 (N_35998,N_34423,N_34100);
xnor U35999 (N_35999,N_34670,N_34733);
xnor U36000 (N_36000,N_35744,N_35150);
xor U36001 (N_36001,N_35510,N_35090);
nor U36002 (N_36002,N_35783,N_35854);
xor U36003 (N_36003,N_35392,N_35784);
nand U36004 (N_36004,N_35277,N_35944);
or U36005 (N_36005,N_35565,N_35776);
nand U36006 (N_36006,N_35694,N_35999);
nand U36007 (N_36007,N_35559,N_35575);
nand U36008 (N_36008,N_35096,N_35019);
xor U36009 (N_36009,N_35189,N_35493);
nand U36010 (N_36010,N_35582,N_35601);
xor U36011 (N_36011,N_35847,N_35233);
and U36012 (N_36012,N_35059,N_35679);
nor U36013 (N_36013,N_35683,N_35162);
xor U36014 (N_36014,N_35614,N_35142);
xnor U36015 (N_36015,N_35182,N_35304);
and U36016 (N_36016,N_35197,N_35455);
xnor U36017 (N_36017,N_35836,N_35775);
nor U36018 (N_36018,N_35320,N_35237);
and U36019 (N_36019,N_35037,N_35617);
or U36020 (N_36020,N_35957,N_35312);
xnor U36021 (N_36021,N_35170,N_35193);
nor U36022 (N_36022,N_35066,N_35507);
nor U36023 (N_36023,N_35456,N_35763);
xor U36024 (N_36024,N_35378,N_35923);
xor U36025 (N_36025,N_35281,N_35438);
xor U36026 (N_36026,N_35805,N_35143);
and U36027 (N_36027,N_35140,N_35508);
and U36028 (N_36028,N_35433,N_35983);
nand U36029 (N_36029,N_35905,N_35893);
nor U36030 (N_36030,N_35722,N_35223);
nor U36031 (N_36031,N_35502,N_35819);
and U36032 (N_36032,N_35914,N_35731);
xnor U36033 (N_36033,N_35425,N_35877);
nor U36034 (N_36034,N_35930,N_35029);
nor U36035 (N_36035,N_35327,N_35603);
and U36036 (N_36036,N_35286,N_35138);
nand U36037 (N_36037,N_35837,N_35301);
or U36038 (N_36038,N_35106,N_35955);
nand U36039 (N_36039,N_35466,N_35405);
or U36040 (N_36040,N_35191,N_35872);
and U36041 (N_36041,N_35423,N_35751);
and U36042 (N_36042,N_35366,N_35483);
or U36043 (N_36043,N_35319,N_35082);
or U36044 (N_36044,N_35710,N_35398);
nor U36045 (N_36045,N_35463,N_35219);
or U36046 (N_36046,N_35401,N_35504);
and U36047 (N_36047,N_35210,N_35501);
or U36048 (N_36048,N_35512,N_35895);
and U36049 (N_36049,N_35478,N_35678);
xnor U36050 (N_36050,N_35546,N_35645);
nor U36051 (N_36051,N_35748,N_35639);
and U36052 (N_36052,N_35095,N_35781);
nand U36053 (N_36053,N_35214,N_35061);
and U36054 (N_36054,N_35618,N_35026);
nor U36055 (N_36055,N_35631,N_35410);
or U36056 (N_36056,N_35995,N_35093);
nor U36057 (N_36057,N_35755,N_35929);
or U36058 (N_36058,N_35782,N_35712);
and U36059 (N_36059,N_35531,N_35229);
nand U36060 (N_36060,N_35012,N_35899);
xnor U36061 (N_36061,N_35988,N_35462);
nor U36062 (N_36062,N_35823,N_35180);
or U36063 (N_36063,N_35584,N_35457);
and U36064 (N_36064,N_35109,N_35033);
and U36065 (N_36065,N_35567,N_35244);
nor U36066 (N_36066,N_35856,N_35717);
xor U36067 (N_36067,N_35358,N_35183);
and U36068 (N_36068,N_35939,N_35052);
and U36069 (N_36069,N_35652,N_35777);
nor U36070 (N_36070,N_35144,N_35393);
and U36071 (N_36071,N_35676,N_35533);
or U36072 (N_36072,N_35857,N_35175);
nand U36073 (N_36073,N_35650,N_35928);
nand U36074 (N_36074,N_35972,N_35389);
xor U36075 (N_36075,N_35373,N_35453);
or U36076 (N_36076,N_35450,N_35900);
and U36077 (N_36077,N_35660,N_35025);
or U36078 (N_36078,N_35412,N_35843);
or U36079 (N_36079,N_35612,N_35677);
or U36080 (N_36080,N_35635,N_35297);
or U36081 (N_36081,N_35815,N_35613);
nand U36082 (N_36082,N_35806,N_35201);
nand U36083 (N_36083,N_35813,N_35176);
or U36084 (N_36084,N_35675,N_35111);
and U36085 (N_36085,N_35699,N_35786);
nand U36086 (N_36086,N_35043,N_35121);
nand U36087 (N_36087,N_35313,N_35913);
or U36088 (N_36088,N_35049,N_35765);
nand U36089 (N_36089,N_35147,N_35658);
and U36090 (N_36090,N_35761,N_35842);
and U36091 (N_36091,N_35442,N_35368);
nand U36092 (N_36092,N_35374,N_35728);
nor U36093 (N_36093,N_35561,N_35271);
nor U36094 (N_36094,N_35866,N_35719);
xnor U36095 (N_36095,N_35758,N_35942);
nor U36096 (N_36096,N_35355,N_35384);
or U36097 (N_36097,N_35894,N_35338);
nand U36098 (N_36098,N_35283,N_35752);
and U36099 (N_36099,N_35377,N_35104);
nand U36100 (N_36100,N_35464,N_35657);
and U36101 (N_36101,N_35080,N_35245);
nor U36102 (N_36102,N_35888,N_35114);
nor U36103 (N_36103,N_35647,N_35395);
and U36104 (N_36104,N_35476,N_35760);
or U36105 (N_36105,N_35159,N_35194);
and U36106 (N_36106,N_35001,N_35703);
or U36107 (N_36107,N_35726,N_35360);
xnor U36108 (N_36108,N_35949,N_35526);
or U36109 (N_36109,N_35042,N_35585);
and U36110 (N_36110,N_35808,N_35127);
nand U36111 (N_36111,N_35824,N_35352);
nand U36112 (N_36112,N_35571,N_35495);
xor U36113 (N_36113,N_35284,N_35084);
nand U36114 (N_36114,N_35048,N_35349);
nor U36115 (N_36115,N_35821,N_35853);
or U36116 (N_36116,N_35308,N_35077);
nor U36117 (N_36117,N_35800,N_35723);
nor U36118 (N_36118,N_35616,N_35344);
and U36119 (N_36119,N_35480,N_35240);
and U36120 (N_36120,N_35000,N_35732);
nand U36121 (N_36121,N_35296,N_35890);
xnor U36122 (N_36122,N_35740,N_35727);
or U36123 (N_36123,N_35709,N_35474);
nand U36124 (N_36124,N_35513,N_35257);
xor U36125 (N_36125,N_35950,N_35880);
nand U36126 (N_36126,N_35573,N_35139);
xnor U36127 (N_36127,N_35145,N_35058);
nor U36128 (N_36128,N_35619,N_35970);
nor U36129 (N_36129,N_35185,N_35943);
nand U36130 (N_36130,N_35045,N_35413);
xnor U36131 (N_36131,N_35769,N_35499);
or U36132 (N_36132,N_35644,N_35115);
and U36133 (N_36133,N_35586,N_35009);
nand U36134 (N_36134,N_35372,N_35060);
or U36135 (N_36135,N_35874,N_35956);
or U36136 (N_36136,N_35278,N_35216);
and U36137 (N_36137,N_35295,N_35449);
or U36138 (N_36138,N_35576,N_35506);
nand U36139 (N_36139,N_35226,N_35404);
xor U36140 (N_36140,N_35103,N_35259);
nand U36141 (N_36141,N_35430,N_35535);
and U36142 (N_36142,N_35509,N_35399);
or U36143 (N_36143,N_35231,N_35912);
nor U36144 (N_36144,N_35055,N_35908);
and U36145 (N_36145,N_35460,N_35884);
nand U36146 (N_36146,N_35873,N_35337);
nand U36147 (N_36147,N_35332,N_35641);
xnor U36148 (N_36148,N_35864,N_35518);
or U36149 (N_36149,N_35239,N_35486);
xor U36150 (N_36150,N_35705,N_35555);
nand U36151 (N_36151,N_35896,N_35918);
xnor U36152 (N_36152,N_35081,N_35353);
nor U36153 (N_36153,N_35437,N_35065);
or U36154 (N_36154,N_35982,N_35276);
nor U36155 (N_36155,N_35217,N_35467);
nor U36156 (N_36156,N_35347,N_35521);
or U36157 (N_36157,N_35580,N_35110);
nand U36158 (N_36158,N_35620,N_35346);
nor U36159 (N_36159,N_35729,N_35316);
or U36160 (N_36160,N_35633,N_35632);
and U36161 (N_36161,N_35906,N_35323);
or U36162 (N_36162,N_35876,N_35051);
or U36163 (N_36163,N_35730,N_35623);
nand U36164 (N_36164,N_35196,N_35306);
or U36165 (N_36165,N_35882,N_35814);
and U36166 (N_36166,N_35247,N_35889);
nand U36167 (N_36167,N_35964,N_35701);
nor U36168 (N_36168,N_35519,N_35577);
nor U36169 (N_36169,N_35054,N_35883);
nor U36170 (N_36170,N_35131,N_35285);
nand U36171 (N_36171,N_35097,N_35596);
nor U36172 (N_36172,N_35962,N_35282);
nand U36173 (N_36173,N_35440,N_35544);
nand U36174 (N_36174,N_35046,N_35788);
and U36175 (N_36175,N_35700,N_35479);
nor U36176 (N_36176,N_35790,N_35976);
nor U36177 (N_36177,N_35269,N_35870);
and U36178 (N_36178,N_35021,N_35141);
nand U36179 (N_36179,N_35868,N_35986);
nand U36180 (N_36180,N_35572,N_35164);
nor U36181 (N_36181,N_35047,N_35005);
nand U36182 (N_36182,N_35382,N_35706);
nand U36183 (N_36183,N_35648,N_35032);
xor U36184 (N_36184,N_35628,N_35322);
xnor U36185 (N_36185,N_35498,N_35738);
and U36186 (N_36186,N_35465,N_35985);
or U36187 (N_36187,N_35579,N_35746);
nand U36188 (N_36188,N_35148,N_35318);
and U36189 (N_36189,N_35951,N_35023);
nor U36190 (N_36190,N_35340,N_35898);
or U36191 (N_36191,N_35330,N_35625);
or U36192 (N_36192,N_35414,N_35887);
xnor U36193 (N_36193,N_35200,N_35852);
or U36194 (N_36194,N_35671,N_35960);
xnor U36195 (N_36195,N_35325,N_35522);
and U36196 (N_36196,N_35451,N_35803);
nor U36197 (N_36197,N_35538,N_35188);
or U36198 (N_36198,N_35356,N_35865);
nand U36199 (N_36199,N_35469,N_35850);
and U36200 (N_36200,N_35024,N_35946);
nand U36201 (N_36201,N_35711,N_35454);
or U36202 (N_36202,N_35428,N_35006);
xor U36203 (N_36203,N_35926,N_35030);
nand U36204 (N_36204,N_35303,N_35569);
nor U36205 (N_36205,N_35932,N_35720);
xnor U36206 (N_36206,N_35416,N_35621);
nand U36207 (N_36207,N_35181,N_35400);
nand U36208 (N_36208,N_35708,N_35801);
and U36209 (N_36209,N_35593,N_35941);
and U36210 (N_36210,N_35468,N_35246);
and U36211 (N_36211,N_35750,N_35497);
nand U36212 (N_36212,N_35792,N_35691);
and U36213 (N_36213,N_35947,N_35473);
nor U36214 (N_36214,N_35937,N_35481);
nand U36215 (N_36215,N_35073,N_35636);
or U36216 (N_36216,N_35491,N_35132);
nor U36217 (N_36217,N_35161,N_35662);
nor U36218 (N_36218,N_35967,N_35979);
nand U36219 (N_36219,N_35044,N_35153);
nand U36220 (N_36220,N_35489,N_35445);
nor U36221 (N_36221,N_35721,N_35387);
nand U36222 (N_36222,N_35698,N_35064);
nand U36223 (N_36223,N_35258,N_35380);
nand U36224 (N_36224,N_35687,N_35275);
or U36225 (N_36225,N_35654,N_35213);
xor U36226 (N_36226,N_35600,N_35343);
nand U36227 (N_36227,N_35554,N_35050);
and U36228 (N_36228,N_35403,N_35235);
nand U36229 (N_36229,N_35597,N_35371);
xor U36230 (N_36230,N_35649,N_35326);
nor U36231 (N_36231,N_35102,N_35133);
and U36232 (N_36232,N_35520,N_35830);
nand U36233 (N_36233,N_35968,N_35293);
or U36234 (N_36234,N_35839,N_35379);
xnor U36235 (N_36235,N_35749,N_35838);
or U36236 (N_36236,N_35485,N_35190);
or U36237 (N_36237,N_35958,N_35350);
or U36238 (N_36238,N_35171,N_35622);
and U36239 (N_36239,N_35891,N_35859);
xor U36240 (N_36240,N_35039,N_35415);
nor U36241 (N_36241,N_35434,N_35411);
nand U36242 (N_36242,N_35664,N_35990);
xnor U36243 (N_36243,N_35359,N_35804);
xor U36244 (N_36244,N_35195,N_35424);
nor U36245 (N_36245,N_35910,N_35909);
and U36246 (N_36246,N_35270,N_35779);
and U36247 (N_36247,N_35028,N_35989);
and U36248 (N_36248,N_35288,N_35100);
and U36249 (N_36249,N_35653,N_35503);
nor U36250 (N_36250,N_35690,N_35655);
nor U36251 (N_36251,N_35470,N_35177);
xor U36252 (N_36252,N_35695,N_35108);
or U36253 (N_36253,N_35643,N_35391);
xor U36254 (N_36254,N_35232,N_35530);
or U36255 (N_36255,N_35552,N_35785);
nor U36256 (N_36256,N_35178,N_35529);
and U36257 (N_36257,N_35444,N_35797);
xnor U36258 (N_36258,N_35205,N_35290);
and U36259 (N_36259,N_35915,N_35543);
nand U36260 (N_36260,N_35668,N_35250);
nor U36261 (N_36261,N_35608,N_35835);
xnor U36262 (N_36262,N_35329,N_35809);
nor U36263 (N_36263,N_35274,N_35828);
nor U36264 (N_36264,N_35459,N_35624);
nand U36265 (N_36265,N_35163,N_35432);
xor U36266 (N_36266,N_35266,N_35822);
nand U36267 (N_36267,N_35085,N_35407);
or U36268 (N_36268,N_35532,N_35560);
and U36269 (N_36269,N_35638,N_35419);
nand U36270 (N_36270,N_35673,N_35260);
xnor U36271 (N_36271,N_35994,N_35186);
nor U36272 (N_36272,N_35766,N_35092);
nand U36273 (N_36273,N_35362,N_35429);
xor U36274 (N_36274,N_35844,N_35475);
nand U36275 (N_36275,N_35057,N_35581);
or U36276 (N_36276,N_35772,N_35072);
nor U36277 (N_36277,N_35435,N_35919);
xor U36278 (N_36278,N_35827,N_35574);
and U36279 (N_36279,N_35524,N_35137);
xnor U36280 (N_36280,N_35665,N_35667);
or U36281 (N_36281,N_35484,N_35680);
nand U36282 (N_36282,N_35354,N_35611);
nor U36283 (N_36283,N_35056,N_35551);
xnor U36284 (N_36284,N_35192,N_35659);
nand U36285 (N_36285,N_35487,N_35692);
and U36286 (N_36286,N_35774,N_35166);
nand U36287 (N_36287,N_35089,N_35417);
nor U36288 (N_36288,N_35242,N_35490);
or U36289 (N_36289,N_35129,N_35158);
nand U36290 (N_36290,N_35291,N_35672);
xor U36291 (N_36291,N_35074,N_35079);
nor U36292 (N_36292,N_35627,N_35549);
and U36293 (N_36293,N_35292,N_35402);
or U36294 (N_36294,N_35020,N_35253);
nand U36295 (N_36295,N_35793,N_35591);
nor U36296 (N_36296,N_35878,N_35458);
and U36297 (N_36297,N_35369,N_35826);
nand U36298 (N_36298,N_35441,N_35336);
and U36299 (N_36299,N_35851,N_35390);
nand U36300 (N_36300,N_35034,N_35307);
nor U36301 (N_36301,N_35254,N_35916);
and U36302 (N_36302,N_35965,N_35992);
or U36303 (N_36303,N_35791,N_35626);
xor U36304 (N_36304,N_35169,N_35642);
xor U36305 (N_36305,N_35564,N_35743);
and U36306 (N_36306,N_35394,N_35220);
or U36307 (N_36307,N_35681,N_35126);
nor U36308 (N_36308,N_35385,N_35871);
and U36309 (N_36309,N_35505,N_35426);
or U36310 (N_36310,N_35963,N_35041);
nor U36311 (N_36311,N_35810,N_35798);
nor U36312 (N_36312,N_35255,N_35452);
and U36313 (N_36313,N_35768,N_35155);
xor U36314 (N_36314,N_35829,N_35607);
and U36315 (N_36315,N_35834,N_35527);
and U36316 (N_36316,N_35536,N_35725);
nor U36317 (N_36317,N_35845,N_35818);
and U36318 (N_36318,N_35091,N_35172);
or U36319 (N_36319,N_35892,N_35855);
nor U36320 (N_36320,N_35609,N_35764);
and U36321 (N_36321,N_35015,N_35563);
nor U36322 (N_36322,N_35817,N_35339);
nand U36323 (N_36323,N_35718,N_35787);
xnor U36324 (N_36324,N_35209,N_35971);
xnor U36325 (N_36325,N_35832,N_35173);
nand U36326 (N_36326,N_35361,N_35228);
nand U36327 (N_36327,N_35767,N_35849);
or U36328 (N_36328,N_35541,N_35098);
xnor U36329 (N_36329,N_35737,N_35969);
nor U36330 (N_36330,N_35966,N_35702);
or U36331 (N_36331,N_35334,N_35348);
nor U36332 (N_36332,N_35934,N_35206);
nand U36333 (N_36333,N_35436,N_35500);
and U36334 (N_36334,N_35027,N_35472);
nor U36335 (N_36335,N_35003,N_35997);
or U36336 (N_36336,N_35342,N_35207);
and U36337 (N_36337,N_35867,N_35187);
nor U36338 (N_36338,N_35588,N_35224);
nand U36339 (N_36339,N_35101,N_35911);
nand U36340 (N_36340,N_35300,N_35525);
xnor U36341 (N_36341,N_35940,N_35007);
or U36342 (N_36342,N_35446,N_35494);
nand U36343 (N_36343,N_35540,N_35184);
or U36344 (N_36344,N_35086,N_35036);
nand U36345 (N_36345,N_35553,N_35149);
nor U36346 (N_36346,N_35230,N_35595);
xor U36347 (N_36347,N_35396,N_35674);
nor U36348 (N_36348,N_35302,N_35053);
nand U36349 (N_36349,N_35714,N_35202);
or U36350 (N_36350,N_35321,N_35125);
nor U36351 (N_36351,N_35087,N_35901);
nand U36352 (N_36352,N_35907,N_35038);
nor U36353 (N_36353,N_35461,N_35208);
or U36354 (N_36354,N_35167,N_35328);
xnor U36355 (N_36355,N_35747,N_35663);
or U36356 (N_36356,N_35534,N_35248);
xnor U36357 (N_36357,N_35981,N_35067);
nor U36358 (N_36358,N_35482,N_35795);
xor U36359 (N_36359,N_35756,N_35954);
and U36360 (N_36360,N_35629,N_35587);
and U36361 (N_36361,N_35933,N_35789);
and U36362 (N_36362,N_35980,N_35757);
nand U36363 (N_36363,N_35682,N_35365);
or U36364 (N_36364,N_35861,N_35204);
nand U36365 (N_36365,N_35739,N_35151);
xor U36366 (N_36366,N_35222,N_35686);
nand U36367 (N_36367,N_35715,N_35961);
or U36368 (N_36368,N_35754,N_35707);
nor U36369 (N_36369,N_35589,N_35936);
or U36370 (N_36370,N_35528,N_35548);
xnor U36371 (N_36371,N_35018,N_35031);
xor U36372 (N_36372,N_35345,N_35071);
xnor U36373 (N_36373,N_35279,N_35218);
or U36374 (N_36374,N_35203,N_35816);
and U36375 (N_36375,N_35397,N_35566);
nand U36376 (N_36376,N_35212,N_35116);
nand U36377 (N_36377,N_35124,N_35938);
xor U36378 (N_36378,N_35558,N_35174);
and U36379 (N_36379,N_35858,N_35802);
or U36380 (N_36380,N_35696,N_35753);
xnor U36381 (N_36381,N_35762,N_35078);
and U36382 (N_36382,N_35615,N_35386);
or U36383 (N_36383,N_35408,N_35122);
and U36384 (N_36384,N_35119,N_35160);
xor U36385 (N_36385,N_35118,N_35381);
nand U36386 (N_36386,N_35807,N_35123);
xnor U36387 (N_36387,N_35651,N_35902);
xnor U36388 (N_36388,N_35846,N_35735);
or U36389 (N_36389,N_35341,N_35697);
or U36390 (N_36390,N_35040,N_35448);
xor U36391 (N_36391,N_35152,N_35825);
xor U36392 (N_36392,N_35070,N_35076);
and U36393 (N_36393,N_35917,N_35897);
nand U36394 (N_36394,N_35011,N_35570);
and U36395 (N_36395,N_35146,N_35831);
and U36396 (N_36396,N_35948,N_35606);
or U36397 (N_36397,N_35733,N_35557);
or U36398 (N_36398,N_35578,N_35771);
xnor U36399 (N_36399,N_35590,N_35920);
nor U36400 (N_36400,N_35075,N_35684);
and U36401 (N_36401,N_35602,N_35511);
or U36402 (N_36402,N_35812,N_35646);
xor U36403 (N_36403,N_35305,N_35351);
xnor U36404 (N_36404,N_35977,N_35427);
or U36405 (N_36405,N_35973,N_35267);
xor U36406 (N_36406,N_35922,N_35273);
and U36407 (N_36407,N_35311,N_35656);
nor U36408 (N_36408,N_35666,N_35252);
nor U36409 (N_36409,N_35156,N_35885);
nand U36410 (N_36410,N_35243,N_35736);
or U36411 (N_36411,N_35693,N_35068);
nand U36412 (N_36412,N_35241,N_35251);
and U36413 (N_36413,N_35539,N_35376);
or U36414 (N_36414,N_35991,N_35324);
or U36415 (N_36415,N_35496,N_35516);
nand U36416 (N_36416,N_35357,N_35780);
nand U36417 (N_36417,N_35713,N_35099);
nor U36418 (N_36418,N_35105,N_35848);
nor U36419 (N_36419,N_35136,N_35741);
and U36420 (N_36420,N_35724,N_35331);
nor U36421 (N_36421,N_35333,N_35262);
or U36422 (N_36422,N_35375,N_35863);
nand U36423 (N_36423,N_35904,N_35925);
or U36424 (N_36424,N_35309,N_35370);
or U36425 (N_36425,N_35869,N_35592);
xnor U36426 (N_36426,N_35154,N_35335);
or U36427 (N_36427,N_35661,N_35094);
nand U36428 (N_36428,N_35537,N_35112);
nor U36429 (N_36429,N_35975,N_35583);
or U36430 (N_36430,N_35996,N_35117);
nor U36431 (N_36431,N_35562,N_35249);
nand U36432 (N_36432,N_35069,N_35299);
or U36433 (N_36433,N_35264,N_35841);
nand U36434 (N_36434,N_35179,N_35310);
nand U36435 (N_36435,N_35594,N_35272);
xnor U36436 (N_36436,N_35685,N_35022);
xor U36437 (N_36437,N_35545,N_35833);
or U36438 (N_36438,N_35261,N_35704);
nand U36439 (N_36439,N_35669,N_35688);
or U36440 (N_36440,N_35935,N_35013);
nand U36441 (N_36441,N_35931,N_35927);
and U36442 (N_36442,N_35168,N_35383);
nand U36443 (N_36443,N_35514,N_35016);
or U36444 (N_36444,N_35517,N_35014);
xnor U36445 (N_36445,N_35130,N_35924);
nand U36446 (N_36446,N_35364,N_35263);
xor U36447 (N_36447,N_35234,N_35875);
nand U36448 (N_36448,N_35820,N_35998);
nand U36449 (N_36449,N_35550,N_35879);
nand U36450 (N_36450,N_35598,N_35280);
or U36451 (N_36451,N_35811,N_35083);
and U36452 (N_36452,N_35640,N_35881);
nor U36453 (N_36453,N_35120,N_35984);
or U36454 (N_36454,N_35689,N_35294);
and U36455 (N_36455,N_35388,N_35987);
nor U36456 (N_36456,N_35317,N_35409);
and U36457 (N_36457,N_35716,N_35225);
nor U36458 (N_36458,N_35135,N_35974);
nor U36459 (N_36459,N_35978,N_35447);
and U36460 (N_36460,N_35599,N_35422);
nand U36461 (N_36461,N_35017,N_35742);
or U36462 (N_36462,N_35157,N_35421);
or U36463 (N_36463,N_35605,N_35418);
and U36464 (N_36464,N_35420,N_35406);
nor U36465 (N_36465,N_35315,N_35314);
xnor U36466 (N_36466,N_35556,N_35637);
or U36467 (N_36467,N_35604,N_35945);
and U36468 (N_36468,N_35063,N_35128);
xor U36469 (N_36469,N_35265,N_35903);
nand U36470 (N_36470,N_35745,N_35367);
and U36471 (N_36471,N_35993,N_35547);
and U36472 (N_36472,N_35778,N_35008);
nand U36473 (N_36473,N_35298,N_35840);
nor U36474 (N_36474,N_35238,N_35471);
nor U36475 (N_36475,N_35134,N_35035);
and U36476 (N_36476,N_35488,N_35799);
or U36477 (N_36477,N_35492,N_35953);
or U36478 (N_36478,N_35268,N_35515);
nor U36479 (N_36479,N_35431,N_35004);
nor U36480 (N_36480,N_35634,N_35796);
or U36481 (N_36481,N_35165,N_35568);
nand U36482 (N_36482,N_35062,N_35088);
or U36483 (N_36483,N_35477,N_35256);
and U36484 (N_36484,N_35921,N_35002);
and U36485 (N_36485,N_35670,N_35443);
xor U36486 (N_36486,N_35959,N_35952);
xnor U36487 (N_36487,N_35113,N_35107);
nand U36488 (N_36488,N_35221,N_35363);
xor U36489 (N_36489,N_35630,N_35734);
nand U36490 (N_36490,N_35770,N_35862);
nand U36491 (N_36491,N_35199,N_35227);
or U36492 (N_36492,N_35794,N_35198);
and U36493 (N_36493,N_35287,N_35236);
nand U36494 (N_36494,N_35215,N_35289);
xnor U36495 (N_36495,N_35773,N_35610);
nand U36496 (N_36496,N_35542,N_35211);
xor U36497 (N_36497,N_35523,N_35759);
xor U36498 (N_36498,N_35886,N_35860);
nand U36499 (N_36499,N_35010,N_35439);
nor U36500 (N_36500,N_35301,N_35503);
or U36501 (N_36501,N_35106,N_35763);
nand U36502 (N_36502,N_35352,N_35019);
xnor U36503 (N_36503,N_35264,N_35792);
nand U36504 (N_36504,N_35689,N_35698);
xor U36505 (N_36505,N_35284,N_35267);
nand U36506 (N_36506,N_35113,N_35701);
and U36507 (N_36507,N_35911,N_35176);
and U36508 (N_36508,N_35904,N_35943);
xnor U36509 (N_36509,N_35039,N_35345);
nor U36510 (N_36510,N_35613,N_35135);
nor U36511 (N_36511,N_35974,N_35258);
xor U36512 (N_36512,N_35865,N_35315);
xnor U36513 (N_36513,N_35168,N_35069);
xnor U36514 (N_36514,N_35964,N_35500);
and U36515 (N_36515,N_35372,N_35898);
xor U36516 (N_36516,N_35414,N_35663);
xor U36517 (N_36517,N_35683,N_35937);
nand U36518 (N_36518,N_35250,N_35134);
xor U36519 (N_36519,N_35036,N_35831);
and U36520 (N_36520,N_35684,N_35507);
nor U36521 (N_36521,N_35045,N_35766);
nand U36522 (N_36522,N_35180,N_35791);
nor U36523 (N_36523,N_35759,N_35289);
or U36524 (N_36524,N_35332,N_35268);
or U36525 (N_36525,N_35651,N_35494);
and U36526 (N_36526,N_35963,N_35337);
xnor U36527 (N_36527,N_35562,N_35883);
or U36528 (N_36528,N_35830,N_35392);
xor U36529 (N_36529,N_35439,N_35166);
nor U36530 (N_36530,N_35451,N_35047);
xor U36531 (N_36531,N_35213,N_35470);
nor U36532 (N_36532,N_35540,N_35197);
nor U36533 (N_36533,N_35887,N_35059);
nand U36534 (N_36534,N_35138,N_35812);
nor U36535 (N_36535,N_35839,N_35996);
or U36536 (N_36536,N_35479,N_35812);
nor U36537 (N_36537,N_35177,N_35361);
xor U36538 (N_36538,N_35544,N_35703);
nor U36539 (N_36539,N_35675,N_35244);
and U36540 (N_36540,N_35346,N_35324);
xor U36541 (N_36541,N_35958,N_35888);
xor U36542 (N_36542,N_35771,N_35057);
and U36543 (N_36543,N_35337,N_35226);
nand U36544 (N_36544,N_35131,N_35871);
nor U36545 (N_36545,N_35959,N_35262);
nand U36546 (N_36546,N_35881,N_35551);
xor U36547 (N_36547,N_35899,N_35622);
nor U36548 (N_36548,N_35608,N_35990);
nand U36549 (N_36549,N_35999,N_35913);
nor U36550 (N_36550,N_35854,N_35550);
nand U36551 (N_36551,N_35727,N_35195);
nor U36552 (N_36552,N_35998,N_35425);
nand U36553 (N_36553,N_35375,N_35585);
and U36554 (N_36554,N_35564,N_35687);
and U36555 (N_36555,N_35037,N_35461);
xor U36556 (N_36556,N_35203,N_35350);
xnor U36557 (N_36557,N_35493,N_35685);
or U36558 (N_36558,N_35998,N_35057);
nor U36559 (N_36559,N_35101,N_35750);
or U36560 (N_36560,N_35578,N_35965);
nand U36561 (N_36561,N_35816,N_35519);
nand U36562 (N_36562,N_35057,N_35016);
nor U36563 (N_36563,N_35028,N_35086);
or U36564 (N_36564,N_35707,N_35670);
or U36565 (N_36565,N_35722,N_35431);
nand U36566 (N_36566,N_35808,N_35796);
nor U36567 (N_36567,N_35810,N_35550);
and U36568 (N_36568,N_35601,N_35741);
and U36569 (N_36569,N_35978,N_35364);
or U36570 (N_36570,N_35104,N_35014);
and U36571 (N_36571,N_35804,N_35757);
nor U36572 (N_36572,N_35207,N_35940);
or U36573 (N_36573,N_35311,N_35173);
and U36574 (N_36574,N_35694,N_35267);
and U36575 (N_36575,N_35074,N_35483);
and U36576 (N_36576,N_35083,N_35419);
nor U36577 (N_36577,N_35257,N_35701);
and U36578 (N_36578,N_35699,N_35332);
xor U36579 (N_36579,N_35846,N_35368);
and U36580 (N_36580,N_35684,N_35486);
nor U36581 (N_36581,N_35279,N_35819);
nor U36582 (N_36582,N_35401,N_35563);
xor U36583 (N_36583,N_35769,N_35827);
xnor U36584 (N_36584,N_35122,N_35018);
xnor U36585 (N_36585,N_35372,N_35316);
and U36586 (N_36586,N_35133,N_35474);
xnor U36587 (N_36587,N_35974,N_35129);
nor U36588 (N_36588,N_35662,N_35464);
nand U36589 (N_36589,N_35270,N_35864);
or U36590 (N_36590,N_35321,N_35562);
xor U36591 (N_36591,N_35794,N_35126);
nand U36592 (N_36592,N_35925,N_35815);
or U36593 (N_36593,N_35302,N_35469);
nand U36594 (N_36594,N_35922,N_35854);
or U36595 (N_36595,N_35189,N_35753);
xnor U36596 (N_36596,N_35737,N_35896);
nand U36597 (N_36597,N_35783,N_35320);
nor U36598 (N_36598,N_35531,N_35629);
nand U36599 (N_36599,N_35294,N_35653);
and U36600 (N_36600,N_35620,N_35660);
nand U36601 (N_36601,N_35064,N_35281);
xnor U36602 (N_36602,N_35034,N_35437);
nor U36603 (N_36603,N_35522,N_35786);
nand U36604 (N_36604,N_35719,N_35985);
nor U36605 (N_36605,N_35951,N_35857);
or U36606 (N_36606,N_35442,N_35264);
nor U36607 (N_36607,N_35205,N_35431);
or U36608 (N_36608,N_35137,N_35878);
or U36609 (N_36609,N_35849,N_35856);
and U36610 (N_36610,N_35473,N_35811);
or U36611 (N_36611,N_35742,N_35974);
nand U36612 (N_36612,N_35427,N_35707);
and U36613 (N_36613,N_35006,N_35217);
nand U36614 (N_36614,N_35967,N_35044);
or U36615 (N_36615,N_35431,N_35621);
nor U36616 (N_36616,N_35508,N_35088);
and U36617 (N_36617,N_35150,N_35184);
or U36618 (N_36618,N_35289,N_35221);
or U36619 (N_36619,N_35275,N_35671);
nand U36620 (N_36620,N_35999,N_35235);
xor U36621 (N_36621,N_35759,N_35232);
nor U36622 (N_36622,N_35557,N_35087);
nand U36623 (N_36623,N_35556,N_35268);
xor U36624 (N_36624,N_35782,N_35662);
and U36625 (N_36625,N_35207,N_35195);
or U36626 (N_36626,N_35103,N_35744);
or U36627 (N_36627,N_35992,N_35346);
xnor U36628 (N_36628,N_35407,N_35322);
nand U36629 (N_36629,N_35251,N_35830);
nor U36630 (N_36630,N_35216,N_35968);
nor U36631 (N_36631,N_35617,N_35437);
nand U36632 (N_36632,N_35474,N_35044);
nor U36633 (N_36633,N_35966,N_35652);
nand U36634 (N_36634,N_35468,N_35471);
xnor U36635 (N_36635,N_35427,N_35023);
nand U36636 (N_36636,N_35062,N_35665);
or U36637 (N_36637,N_35059,N_35675);
and U36638 (N_36638,N_35627,N_35629);
nand U36639 (N_36639,N_35560,N_35824);
and U36640 (N_36640,N_35713,N_35055);
nand U36641 (N_36641,N_35199,N_35402);
nor U36642 (N_36642,N_35948,N_35101);
or U36643 (N_36643,N_35622,N_35102);
nor U36644 (N_36644,N_35041,N_35241);
or U36645 (N_36645,N_35586,N_35708);
or U36646 (N_36646,N_35236,N_35105);
and U36647 (N_36647,N_35370,N_35627);
nor U36648 (N_36648,N_35630,N_35227);
nor U36649 (N_36649,N_35477,N_35764);
and U36650 (N_36650,N_35205,N_35625);
or U36651 (N_36651,N_35894,N_35230);
xnor U36652 (N_36652,N_35329,N_35109);
nand U36653 (N_36653,N_35366,N_35230);
or U36654 (N_36654,N_35916,N_35988);
xor U36655 (N_36655,N_35204,N_35917);
nor U36656 (N_36656,N_35095,N_35660);
xor U36657 (N_36657,N_35282,N_35452);
nor U36658 (N_36658,N_35860,N_35387);
nand U36659 (N_36659,N_35746,N_35363);
nor U36660 (N_36660,N_35167,N_35922);
or U36661 (N_36661,N_35469,N_35186);
nand U36662 (N_36662,N_35349,N_35408);
and U36663 (N_36663,N_35263,N_35766);
nor U36664 (N_36664,N_35548,N_35723);
nor U36665 (N_36665,N_35680,N_35199);
and U36666 (N_36666,N_35168,N_35326);
nor U36667 (N_36667,N_35067,N_35999);
or U36668 (N_36668,N_35343,N_35981);
nor U36669 (N_36669,N_35355,N_35820);
nor U36670 (N_36670,N_35823,N_35481);
xnor U36671 (N_36671,N_35909,N_35072);
and U36672 (N_36672,N_35075,N_35871);
and U36673 (N_36673,N_35030,N_35228);
nor U36674 (N_36674,N_35311,N_35843);
and U36675 (N_36675,N_35117,N_35337);
xor U36676 (N_36676,N_35534,N_35037);
or U36677 (N_36677,N_35958,N_35440);
xor U36678 (N_36678,N_35019,N_35920);
xnor U36679 (N_36679,N_35413,N_35753);
xor U36680 (N_36680,N_35355,N_35163);
xor U36681 (N_36681,N_35850,N_35631);
and U36682 (N_36682,N_35967,N_35584);
nand U36683 (N_36683,N_35750,N_35166);
nor U36684 (N_36684,N_35191,N_35645);
nor U36685 (N_36685,N_35816,N_35663);
nor U36686 (N_36686,N_35816,N_35446);
and U36687 (N_36687,N_35864,N_35266);
and U36688 (N_36688,N_35439,N_35046);
nand U36689 (N_36689,N_35921,N_35314);
nand U36690 (N_36690,N_35722,N_35330);
nand U36691 (N_36691,N_35904,N_35435);
nand U36692 (N_36692,N_35759,N_35578);
xor U36693 (N_36693,N_35736,N_35850);
or U36694 (N_36694,N_35722,N_35309);
and U36695 (N_36695,N_35631,N_35982);
and U36696 (N_36696,N_35574,N_35074);
nand U36697 (N_36697,N_35112,N_35557);
and U36698 (N_36698,N_35469,N_35432);
nor U36699 (N_36699,N_35412,N_35921);
nor U36700 (N_36700,N_35816,N_35698);
and U36701 (N_36701,N_35559,N_35199);
nor U36702 (N_36702,N_35545,N_35804);
xnor U36703 (N_36703,N_35655,N_35735);
or U36704 (N_36704,N_35018,N_35220);
xor U36705 (N_36705,N_35202,N_35507);
xor U36706 (N_36706,N_35053,N_35369);
nor U36707 (N_36707,N_35258,N_35573);
or U36708 (N_36708,N_35376,N_35441);
xnor U36709 (N_36709,N_35542,N_35139);
or U36710 (N_36710,N_35622,N_35515);
nand U36711 (N_36711,N_35210,N_35830);
nor U36712 (N_36712,N_35953,N_35449);
xor U36713 (N_36713,N_35400,N_35388);
or U36714 (N_36714,N_35746,N_35555);
nor U36715 (N_36715,N_35584,N_35075);
xor U36716 (N_36716,N_35565,N_35733);
nand U36717 (N_36717,N_35763,N_35917);
and U36718 (N_36718,N_35826,N_35637);
or U36719 (N_36719,N_35967,N_35802);
or U36720 (N_36720,N_35117,N_35017);
or U36721 (N_36721,N_35862,N_35711);
nor U36722 (N_36722,N_35011,N_35504);
nand U36723 (N_36723,N_35159,N_35783);
nor U36724 (N_36724,N_35764,N_35184);
nor U36725 (N_36725,N_35557,N_35848);
nor U36726 (N_36726,N_35867,N_35296);
and U36727 (N_36727,N_35004,N_35592);
xor U36728 (N_36728,N_35819,N_35291);
nor U36729 (N_36729,N_35159,N_35677);
nand U36730 (N_36730,N_35696,N_35122);
or U36731 (N_36731,N_35382,N_35606);
or U36732 (N_36732,N_35024,N_35351);
and U36733 (N_36733,N_35271,N_35920);
nand U36734 (N_36734,N_35682,N_35134);
and U36735 (N_36735,N_35456,N_35366);
nand U36736 (N_36736,N_35736,N_35253);
and U36737 (N_36737,N_35936,N_35393);
and U36738 (N_36738,N_35880,N_35892);
nand U36739 (N_36739,N_35701,N_35879);
or U36740 (N_36740,N_35493,N_35014);
or U36741 (N_36741,N_35305,N_35287);
xor U36742 (N_36742,N_35425,N_35959);
xnor U36743 (N_36743,N_35113,N_35431);
nor U36744 (N_36744,N_35054,N_35311);
nand U36745 (N_36745,N_35874,N_35992);
or U36746 (N_36746,N_35144,N_35244);
or U36747 (N_36747,N_35899,N_35767);
or U36748 (N_36748,N_35398,N_35094);
nor U36749 (N_36749,N_35833,N_35920);
xor U36750 (N_36750,N_35295,N_35866);
nor U36751 (N_36751,N_35323,N_35193);
nand U36752 (N_36752,N_35832,N_35709);
xnor U36753 (N_36753,N_35809,N_35122);
and U36754 (N_36754,N_35689,N_35598);
and U36755 (N_36755,N_35577,N_35120);
nand U36756 (N_36756,N_35372,N_35616);
and U36757 (N_36757,N_35192,N_35723);
xor U36758 (N_36758,N_35330,N_35968);
or U36759 (N_36759,N_35325,N_35608);
and U36760 (N_36760,N_35736,N_35260);
xnor U36761 (N_36761,N_35552,N_35005);
xnor U36762 (N_36762,N_35843,N_35273);
or U36763 (N_36763,N_35808,N_35004);
and U36764 (N_36764,N_35858,N_35416);
nand U36765 (N_36765,N_35209,N_35370);
nand U36766 (N_36766,N_35402,N_35953);
xnor U36767 (N_36767,N_35390,N_35504);
and U36768 (N_36768,N_35472,N_35361);
nor U36769 (N_36769,N_35754,N_35842);
nand U36770 (N_36770,N_35081,N_35113);
xor U36771 (N_36771,N_35813,N_35862);
xor U36772 (N_36772,N_35505,N_35647);
xor U36773 (N_36773,N_35173,N_35424);
nor U36774 (N_36774,N_35759,N_35105);
nor U36775 (N_36775,N_35889,N_35982);
xnor U36776 (N_36776,N_35072,N_35402);
and U36777 (N_36777,N_35863,N_35796);
nor U36778 (N_36778,N_35575,N_35701);
nand U36779 (N_36779,N_35525,N_35821);
xnor U36780 (N_36780,N_35207,N_35514);
and U36781 (N_36781,N_35922,N_35825);
nor U36782 (N_36782,N_35100,N_35064);
nor U36783 (N_36783,N_35995,N_35260);
nand U36784 (N_36784,N_35549,N_35673);
and U36785 (N_36785,N_35683,N_35087);
and U36786 (N_36786,N_35484,N_35152);
xnor U36787 (N_36787,N_35095,N_35320);
nor U36788 (N_36788,N_35441,N_35505);
xor U36789 (N_36789,N_35147,N_35054);
xnor U36790 (N_36790,N_35027,N_35034);
or U36791 (N_36791,N_35859,N_35155);
and U36792 (N_36792,N_35750,N_35533);
nand U36793 (N_36793,N_35675,N_35983);
xor U36794 (N_36794,N_35032,N_35244);
or U36795 (N_36795,N_35916,N_35086);
nor U36796 (N_36796,N_35166,N_35180);
and U36797 (N_36797,N_35153,N_35684);
and U36798 (N_36798,N_35314,N_35158);
and U36799 (N_36799,N_35545,N_35174);
xor U36800 (N_36800,N_35738,N_35730);
xnor U36801 (N_36801,N_35466,N_35968);
nor U36802 (N_36802,N_35726,N_35137);
nand U36803 (N_36803,N_35207,N_35881);
nor U36804 (N_36804,N_35495,N_35178);
xor U36805 (N_36805,N_35310,N_35701);
and U36806 (N_36806,N_35288,N_35962);
nand U36807 (N_36807,N_35211,N_35482);
and U36808 (N_36808,N_35116,N_35106);
nor U36809 (N_36809,N_35645,N_35409);
or U36810 (N_36810,N_35552,N_35259);
nand U36811 (N_36811,N_35075,N_35865);
or U36812 (N_36812,N_35893,N_35948);
or U36813 (N_36813,N_35181,N_35758);
nor U36814 (N_36814,N_35408,N_35295);
or U36815 (N_36815,N_35033,N_35331);
nand U36816 (N_36816,N_35751,N_35770);
xnor U36817 (N_36817,N_35884,N_35493);
or U36818 (N_36818,N_35991,N_35854);
or U36819 (N_36819,N_35674,N_35890);
and U36820 (N_36820,N_35880,N_35088);
or U36821 (N_36821,N_35189,N_35988);
nor U36822 (N_36822,N_35862,N_35525);
and U36823 (N_36823,N_35450,N_35689);
nand U36824 (N_36824,N_35622,N_35701);
nor U36825 (N_36825,N_35939,N_35190);
nor U36826 (N_36826,N_35877,N_35674);
and U36827 (N_36827,N_35043,N_35966);
xor U36828 (N_36828,N_35353,N_35407);
or U36829 (N_36829,N_35572,N_35037);
nor U36830 (N_36830,N_35734,N_35364);
xnor U36831 (N_36831,N_35129,N_35556);
nor U36832 (N_36832,N_35714,N_35590);
nand U36833 (N_36833,N_35581,N_35286);
xnor U36834 (N_36834,N_35028,N_35357);
and U36835 (N_36835,N_35987,N_35234);
nor U36836 (N_36836,N_35660,N_35956);
nand U36837 (N_36837,N_35332,N_35057);
and U36838 (N_36838,N_35808,N_35811);
xor U36839 (N_36839,N_35659,N_35807);
nor U36840 (N_36840,N_35925,N_35950);
nor U36841 (N_36841,N_35165,N_35390);
nand U36842 (N_36842,N_35763,N_35473);
nand U36843 (N_36843,N_35001,N_35651);
xor U36844 (N_36844,N_35547,N_35700);
nor U36845 (N_36845,N_35712,N_35936);
xor U36846 (N_36846,N_35573,N_35805);
xnor U36847 (N_36847,N_35166,N_35208);
nor U36848 (N_36848,N_35294,N_35491);
nor U36849 (N_36849,N_35450,N_35298);
or U36850 (N_36850,N_35274,N_35420);
and U36851 (N_36851,N_35262,N_35330);
nand U36852 (N_36852,N_35129,N_35449);
xnor U36853 (N_36853,N_35344,N_35953);
xnor U36854 (N_36854,N_35119,N_35161);
xnor U36855 (N_36855,N_35642,N_35161);
and U36856 (N_36856,N_35523,N_35037);
nand U36857 (N_36857,N_35491,N_35673);
or U36858 (N_36858,N_35016,N_35797);
and U36859 (N_36859,N_35062,N_35524);
nor U36860 (N_36860,N_35116,N_35023);
and U36861 (N_36861,N_35206,N_35923);
and U36862 (N_36862,N_35208,N_35653);
nor U36863 (N_36863,N_35267,N_35870);
nor U36864 (N_36864,N_35261,N_35453);
xnor U36865 (N_36865,N_35046,N_35049);
or U36866 (N_36866,N_35055,N_35919);
nor U36867 (N_36867,N_35700,N_35092);
nand U36868 (N_36868,N_35329,N_35013);
nor U36869 (N_36869,N_35319,N_35540);
and U36870 (N_36870,N_35545,N_35055);
or U36871 (N_36871,N_35738,N_35314);
xnor U36872 (N_36872,N_35187,N_35550);
and U36873 (N_36873,N_35581,N_35329);
nand U36874 (N_36874,N_35572,N_35399);
nor U36875 (N_36875,N_35709,N_35717);
and U36876 (N_36876,N_35207,N_35156);
nor U36877 (N_36877,N_35256,N_35522);
nor U36878 (N_36878,N_35540,N_35094);
xor U36879 (N_36879,N_35519,N_35896);
and U36880 (N_36880,N_35691,N_35725);
nor U36881 (N_36881,N_35322,N_35654);
or U36882 (N_36882,N_35305,N_35610);
or U36883 (N_36883,N_35339,N_35719);
and U36884 (N_36884,N_35147,N_35613);
nand U36885 (N_36885,N_35758,N_35375);
or U36886 (N_36886,N_35515,N_35657);
nand U36887 (N_36887,N_35837,N_35283);
and U36888 (N_36888,N_35945,N_35740);
or U36889 (N_36889,N_35878,N_35478);
xnor U36890 (N_36890,N_35302,N_35054);
or U36891 (N_36891,N_35182,N_35617);
nand U36892 (N_36892,N_35889,N_35282);
and U36893 (N_36893,N_35470,N_35953);
and U36894 (N_36894,N_35149,N_35543);
or U36895 (N_36895,N_35046,N_35058);
and U36896 (N_36896,N_35892,N_35216);
or U36897 (N_36897,N_35792,N_35348);
xor U36898 (N_36898,N_35968,N_35151);
xnor U36899 (N_36899,N_35876,N_35264);
nand U36900 (N_36900,N_35469,N_35221);
or U36901 (N_36901,N_35825,N_35696);
and U36902 (N_36902,N_35530,N_35098);
xnor U36903 (N_36903,N_35064,N_35172);
or U36904 (N_36904,N_35533,N_35394);
or U36905 (N_36905,N_35727,N_35788);
or U36906 (N_36906,N_35185,N_35420);
xnor U36907 (N_36907,N_35954,N_35105);
xor U36908 (N_36908,N_35371,N_35162);
xnor U36909 (N_36909,N_35122,N_35078);
and U36910 (N_36910,N_35626,N_35453);
and U36911 (N_36911,N_35983,N_35553);
nand U36912 (N_36912,N_35854,N_35903);
nor U36913 (N_36913,N_35325,N_35392);
and U36914 (N_36914,N_35185,N_35902);
and U36915 (N_36915,N_35586,N_35782);
or U36916 (N_36916,N_35228,N_35679);
nor U36917 (N_36917,N_35816,N_35691);
or U36918 (N_36918,N_35080,N_35050);
nand U36919 (N_36919,N_35343,N_35936);
nor U36920 (N_36920,N_35209,N_35748);
nor U36921 (N_36921,N_35513,N_35091);
xnor U36922 (N_36922,N_35186,N_35663);
or U36923 (N_36923,N_35522,N_35216);
xor U36924 (N_36924,N_35818,N_35604);
nor U36925 (N_36925,N_35413,N_35317);
and U36926 (N_36926,N_35073,N_35869);
nor U36927 (N_36927,N_35328,N_35771);
nor U36928 (N_36928,N_35494,N_35460);
or U36929 (N_36929,N_35567,N_35390);
nand U36930 (N_36930,N_35994,N_35260);
xnor U36931 (N_36931,N_35262,N_35005);
nor U36932 (N_36932,N_35118,N_35714);
nor U36933 (N_36933,N_35794,N_35877);
and U36934 (N_36934,N_35312,N_35041);
or U36935 (N_36935,N_35072,N_35707);
or U36936 (N_36936,N_35649,N_35833);
xor U36937 (N_36937,N_35107,N_35754);
nor U36938 (N_36938,N_35120,N_35762);
nor U36939 (N_36939,N_35312,N_35086);
or U36940 (N_36940,N_35800,N_35805);
nor U36941 (N_36941,N_35122,N_35510);
xnor U36942 (N_36942,N_35063,N_35210);
or U36943 (N_36943,N_35182,N_35200);
nand U36944 (N_36944,N_35419,N_35278);
nand U36945 (N_36945,N_35899,N_35410);
xor U36946 (N_36946,N_35103,N_35472);
nor U36947 (N_36947,N_35714,N_35391);
or U36948 (N_36948,N_35051,N_35503);
and U36949 (N_36949,N_35558,N_35892);
nand U36950 (N_36950,N_35020,N_35170);
xnor U36951 (N_36951,N_35410,N_35950);
and U36952 (N_36952,N_35522,N_35061);
nor U36953 (N_36953,N_35692,N_35976);
nor U36954 (N_36954,N_35466,N_35303);
xnor U36955 (N_36955,N_35932,N_35507);
and U36956 (N_36956,N_35769,N_35796);
nand U36957 (N_36957,N_35928,N_35757);
and U36958 (N_36958,N_35374,N_35391);
xor U36959 (N_36959,N_35249,N_35140);
xor U36960 (N_36960,N_35413,N_35178);
xnor U36961 (N_36961,N_35606,N_35025);
nand U36962 (N_36962,N_35877,N_35708);
xnor U36963 (N_36963,N_35572,N_35279);
nor U36964 (N_36964,N_35789,N_35027);
xor U36965 (N_36965,N_35332,N_35888);
nand U36966 (N_36966,N_35975,N_35505);
nor U36967 (N_36967,N_35666,N_35394);
or U36968 (N_36968,N_35519,N_35797);
or U36969 (N_36969,N_35748,N_35278);
or U36970 (N_36970,N_35361,N_35705);
nand U36971 (N_36971,N_35075,N_35759);
nand U36972 (N_36972,N_35680,N_35628);
or U36973 (N_36973,N_35598,N_35501);
nand U36974 (N_36974,N_35043,N_35059);
nand U36975 (N_36975,N_35701,N_35423);
and U36976 (N_36976,N_35444,N_35626);
nand U36977 (N_36977,N_35586,N_35234);
nor U36978 (N_36978,N_35458,N_35740);
xor U36979 (N_36979,N_35361,N_35442);
nor U36980 (N_36980,N_35998,N_35239);
nor U36981 (N_36981,N_35080,N_35568);
nor U36982 (N_36982,N_35877,N_35105);
and U36983 (N_36983,N_35540,N_35060);
nand U36984 (N_36984,N_35259,N_35273);
or U36985 (N_36985,N_35780,N_35717);
xor U36986 (N_36986,N_35198,N_35926);
nor U36987 (N_36987,N_35959,N_35155);
nor U36988 (N_36988,N_35582,N_35117);
and U36989 (N_36989,N_35540,N_35144);
nor U36990 (N_36990,N_35705,N_35128);
or U36991 (N_36991,N_35136,N_35857);
and U36992 (N_36992,N_35895,N_35532);
nand U36993 (N_36993,N_35229,N_35626);
or U36994 (N_36994,N_35159,N_35705);
nand U36995 (N_36995,N_35398,N_35944);
or U36996 (N_36996,N_35009,N_35659);
nor U36997 (N_36997,N_35169,N_35771);
xnor U36998 (N_36998,N_35220,N_35445);
xor U36999 (N_36999,N_35169,N_35069);
and U37000 (N_37000,N_36617,N_36534);
nand U37001 (N_37001,N_36983,N_36893);
and U37002 (N_37002,N_36355,N_36524);
nor U37003 (N_37003,N_36265,N_36705);
nor U37004 (N_37004,N_36327,N_36414);
and U37005 (N_37005,N_36647,N_36215);
xnor U37006 (N_37006,N_36956,N_36973);
and U37007 (N_37007,N_36292,N_36251);
nor U37008 (N_37008,N_36106,N_36779);
and U37009 (N_37009,N_36066,N_36429);
or U37010 (N_37010,N_36827,N_36198);
nor U37011 (N_37011,N_36366,N_36299);
xnor U37012 (N_37012,N_36216,N_36924);
nand U37013 (N_37013,N_36758,N_36621);
and U37014 (N_37014,N_36386,N_36682);
and U37015 (N_37015,N_36103,N_36137);
xor U37016 (N_37016,N_36741,N_36563);
nor U37017 (N_37017,N_36116,N_36456);
nor U37018 (N_37018,N_36584,N_36683);
or U37019 (N_37019,N_36290,N_36120);
nand U37020 (N_37020,N_36599,N_36517);
nand U37021 (N_37021,N_36556,N_36908);
and U37022 (N_37022,N_36028,N_36166);
and U37023 (N_37023,N_36281,N_36496);
nand U37024 (N_37024,N_36262,N_36536);
nand U37025 (N_37025,N_36441,N_36587);
nand U37026 (N_37026,N_36760,N_36903);
xor U37027 (N_37027,N_36448,N_36443);
or U37028 (N_37028,N_36296,N_36541);
and U37029 (N_37029,N_36709,N_36364);
xor U37030 (N_37030,N_36527,N_36822);
nor U37031 (N_37031,N_36037,N_36272);
nand U37032 (N_37032,N_36479,N_36119);
nor U37033 (N_37033,N_36884,N_36655);
nand U37034 (N_37034,N_36865,N_36904);
or U37035 (N_37035,N_36189,N_36150);
or U37036 (N_37036,N_36784,N_36252);
nor U37037 (N_37037,N_36177,N_36726);
nor U37038 (N_37038,N_36229,N_36075);
nand U37039 (N_37039,N_36543,N_36487);
xnor U37040 (N_37040,N_36305,N_36521);
nand U37041 (N_37041,N_36812,N_36522);
and U37042 (N_37042,N_36007,N_36986);
nand U37043 (N_37043,N_36424,N_36469);
nand U37044 (N_37044,N_36490,N_36854);
nor U37045 (N_37045,N_36227,N_36768);
nand U37046 (N_37046,N_36248,N_36692);
or U37047 (N_37047,N_36668,N_36352);
and U37048 (N_37048,N_36157,N_36084);
and U37049 (N_37049,N_36025,N_36987);
nand U37050 (N_37050,N_36284,N_36153);
nand U37051 (N_37051,N_36307,N_36205);
nand U37052 (N_37052,N_36373,N_36003);
nor U37053 (N_37053,N_36401,N_36319);
nand U37054 (N_37054,N_36914,N_36143);
xor U37055 (N_37055,N_36944,N_36439);
nand U37056 (N_37056,N_36808,N_36869);
nor U37057 (N_37057,N_36957,N_36354);
or U37058 (N_37058,N_36099,N_36494);
nand U37059 (N_37059,N_36141,N_36491);
and U37060 (N_37060,N_36510,N_36035);
nor U37061 (N_37061,N_36585,N_36308);
xnor U37062 (N_37062,N_36291,N_36253);
or U37063 (N_37063,N_36937,N_36547);
xnor U37064 (N_37064,N_36195,N_36090);
and U37065 (N_37065,N_36169,N_36529);
nor U37066 (N_37066,N_36159,N_36213);
and U37067 (N_37067,N_36241,N_36371);
nand U37068 (N_37068,N_36526,N_36823);
and U37069 (N_37069,N_36151,N_36950);
nand U37070 (N_37070,N_36943,N_36730);
and U37071 (N_37071,N_36382,N_36897);
nand U37072 (N_37072,N_36656,N_36721);
nand U37073 (N_37073,N_36470,N_36498);
and U37074 (N_37074,N_36097,N_36278);
and U37075 (N_37075,N_36481,N_36452);
nand U37076 (N_37076,N_36044,N_36693);
and U37077 (N_37077,N_36385,N_36661);
xnor U37078 (N_37078,N_36791,N_36652);
and U37079 (N_37079,N_36672,N_36107);
or U37080 (N_37080,N_36129,N_36212);
nor U37081 (N_37081,N_36380,N_36597);
and U37082 (N_37082,N_36442,N_36091);
and U37083 (N_37083,N_36562,N_36052);
nor U37084 (N_37084,N_36112,N_36829);
and U37085 (N_37085,N_36646,N_36776);
nor U37086 (N_37086,N_36499,N_36444);
nand U37087 (N_37087,N_36863,N_36847);
and U37088 (N_37088,N_36036,N_36068);
or U37089 (N_37089,N_36088,N_36886);
xnor U37090 (N_37090,N_36340,N_36042);
nand U37091 (N_37091,N_36144,N_36316);
and U37092 (N_37092,N_36894,N_36817);
and U37093 (N_37093,N_36796,N_36834);
or U37094 (N_37094,N_36845,N_36819);
xor U37095 (N_37095,N_36326,N_36882);
and U37096 (N_37096,N_36321,N_36639);
nor U37097 (N_37097,N_36422,N_36853);
nand U37098 (N_37098,N_36773,N_36858);
xor U37099 (N_37099,N_36832,N_36867);
or U37100 (N_37100,N_36875,N_36034);
nor U37101 (N_37101,N_36349,N_36467);
or U37102 (N_37102,N_36336,N_36109);
nand U37103 (N_37103,N_36057,N_36230);
or U37104 (N_37104,N_36322,N_36335);
or U37105 (N_37105,N_36744,N_36079);
xnor U37106 (N_37106,N_36539,N_36952);
nand U37107 (N_37107,N_36070,N_36892);
nand U37108 (N_37108,N_36558,N_36073);
nor U37109 (N_37109,N_36483,N_36977);
or U37110 (N_37110,N_36581,N_36907);
or U37111 (N_37111,N_36619,N_36282);
nand U37112 (N_37112,N_36734,N_36690);
or U37113 (N_37113,N_36675,N_36649);
xor U37114 (N_37114,N_36165,N_36446);
and U37115 (N_37115,N_36023,N_36978);
xor U37116 (N_37116,N_36979,N_36178);
and U37117 (N_37117,N_36715,N_36256);
xnor U37118 (N_37118,N_36011,N_36047);
nor U37119 (N_37119,N_36641,N_36155);
or U37120 (N_37120,N_36206,N_36182);
nor U37121 (N_37121,N_36679,N_36163);
nand U37122 (N_37122,N_36085,N_36849);
xnor U37123 (N_37123,N_36942,N_36799);
xnor U37124 (N_37124,N_36232,N_36502);
or U37125 (N_37125,N_36833,N_36830);
and U37126 (N_37126,N_36664,N_36797);
and U37127 (N_37127,N_36226,N_36633);
nand U37128 (N_37128,N_36008,N_36820);
or U37129 (N_37129,N_36005,N_36301);
or U37130 (N_37130,N_36194,N_36312);
xor U37131 (N_37131,N_36293,N_36379);
or U37132 (N_37132,N_36064,N_36427);
nor U37133 (N_37133,N_36781,N_36273);
and U37134 (N_37134,N_36631,N_36131);
nor U37135 (N_37135,N_36389,N_36866);
xor U37136 (N_37136,N_36501,N_36644);
xor U37137 (N_37137,N_36793,N_36482);
xnor U37138 (N_37138,N_36976,N_36828);
nand U37139 (N_37139,N_36570,N_36686);
xnor U37140 (N_37140,N_36890,N_36304);
or U37141 (N_37141,N_36609,N_36700);
and U37142 (N_37142,N_36771,N_36592);
or U37143 (N_37143,N_36345,N_36513);
nor U37144 (N_37144,N_36925,N_36728);
and U37145 (N_37145,N_36887,N_36255);
xnor U37146 (N_37146,N_36809,N_36782);
and U37147 (N_37147,N_36125,N_36917);
and U37148 (N_37148,N_36571,N_36259);
or U37149 (N_37149,N_36569,N_36939);
or U37150 (N_37150,N_36287,N_36717);
or U37151 (N_37151,N_36329,N_36086);
nand U37152 (N_37152,N_36601,N_36236);
and U37153 (N_37153,N_36121,N_36302);
nor U37154 (N_37154,N_36045,N_36628);
or U37155 (N_37155,N_36818,N_36020);
or U37156 (N_37156,N_36990,N_36916);
xor U37157 (N_37157,N_36605,N_36725);
or U37158 (N_37158,N_36474,N_36146);
nor U37159 (N_37159,N_36362,N_36593);
nand U37160 (N_37160,N_36638,N_36477);
nor U37161 (N_37161,N_36505,N_36409);
or U37162 (N_37162,N_36525,N_36982);
nand U37163 (N_37163,N_36787,N_36283);
or U37164 (N_37164,N_36836,N_36674);
or U37165 (N_37165,N_36673,N_36275);
nand U37166 (N_37166,N_36266,N_36356);
or U37167 (N_37167,N_36685,N_36303);
and U37168 (N_37168,N_36767,N_36486);
nor U37169 (N_37169,N_36136,N_36040);
and U37170 (N_37170,N_36357,N_36101);
or U37171 (N_37171,N_36495,N_36017);
nor U37172 (N_37172,N_36093,N_36413);
xor U37173 (N_37173,N_36848,N_36528);
or U37174 (N_37174,N_36559,N_36161);
nand U37175 (N_37175,N_36430,N_36620);
nor U37176 (N_37176,N_36270,N_36405);
nand U37177 (N_37177,N_36816,N_36004);
and U37178 (N_37178,N_36221,N_36384);
xnor U37179 (N_37179,N_36873,N_36348);
and U37180 (N_37180,N_36122,N_36678);
and U37181 (N_37181,N_36936,N_36995);
nor U37182 (N_37182,N_36190,N_36410);
or U37183 (N_37183,N_36923,N_36915);
nor U37184 (N_37184,N_36723,N_36244);
or U37185 (N_37185,N_36504,N_36999);
nor U37186 (N_37186,N_36343,N_36394);
or U37187 (N_37187,N_36688,N_36934);
nor U37188 (N_37188,N_36269,N_36072);
and U37189 (N_37189,N_36964,N_36802);
and U37190 (N_37190,N_36684,N_36332);
and U37191 (N_37191,N_36350,N_36440);
nor U37192 (N_37192,N_36960,N_36049);
or U37193 (N_37193,N_36399,N_36523);
and U37194 (N_37194,N_36564,N_36026);
nand U37195 (N_37195,N_36984,N_36931);
nand U37196 (N_37196,N_36933,N_36835);
or U37197 (N_37197,N_36650,N_36716);
nand U37198 (N_37198,N_36860,N_36134);
or U37199 (N_37199,N_36298,N_36014);
nor U37200 (N_37200,N_36761,N_36218);
xnor U37201 (N_37201,N_36168,N_36824);
or U37202 (N_37202,N_36503,N_36805);
nor U37203 (N_37203,N_36223,N_36862);
or U37204 (N_37204,N_36344,N_36390);
nand U37205 (N_37205,N_36663,N_36043);
or U37206 (N_37206,N_36268,N_36476);
nor U37207 (N_37207,N_36100,N_36598);
and U37208 (N_37208,N_36162,N_36009);
nand U37209 (N_37209,N_36798,N_36347);
nand U37210 (N_37210,N_36185,N_36825);
and U37211 (N_37211,N_36135,N_36078);
nor U37212 (N_37212,N_36110,N_36772);
nand U37213 (N_37213,N_36718,N_36472);
xor U37214 (N_37214,N_36276,N_36637);
nand U37215 (N_37215,N_36289,N_36220);
and U37216 (N_37216,N_36993,N_36060);
nor U37217 (N_37217,N_36337,N_36128);
nor U37218 (N_37218,N_36083,N_36142);
and U37219 (N_37219,N_36861,N_36224);
xor U37220 (N_37220,N_36967,N_36374);
or U37221 (N_37221,N_36596,N_36065);
and U37222 (N_37222,N_36209,N_36048);
or U37223 (N_37223,N_36665,N_36560);
nor U37224 (N_37224,N_36545,N_36613);
and U37225 (N_37225,N_36234,N_36018);
xnor U37226 (N_37226,N_36520,N_36900);
xnor U37227 (N_37227,N_36397,N_36777);
xnor U37228 (N_37228,N_36500,N_36087);
xor U37229 (N_37229,N_36994,N_36955);
and U37230 (N_37230,N_36192,N_36426);
nor U37231 (N_37231,N_36911,N_36363);
and U37232 (N_37232,N_36445,N_36737);
and U37233 (N_37233,N_36077,N_36659);
xor U37234 (N_37234,N_36738,N_36971);
and U37235 (N_37235,N_36032,N_36434);
nor U37236 (N_37236,N_36877,N_36435);
or U37237 (N_37237,N_36056,N_36774);
nand U37238 (N_37238,N_36970,N_36062);
xnor U37239 (N_37239,N_36881,N_36704);
nor U37240 (N_37240,N_36412,N_36214);
or U37241 (N_37241,N_36670,N_36901);
nor U37242 (N_37242,N_36888,N_36896);
or U37243 (N_37243,N_36616,N_36323);
nor U37244 (N_37244,N_36311,N_36375);
and U37245 (N_37245,N_36769,N_36455);
xnor U37246 (N_37246,N_36515,N_36530);
nand U37247 (N_37247,N_36170,N_36544);
xnor U37248 (N_37248,N_36764,N_36810);
and U37249 (N_37249,N_36436,N_36358);
nand U37250 (N_37250,N_36489,N_36876);
and U37251 (N_37251,N_36181,N_36567);
and U37252 (N_37252,N_36997,N_36369);
and U37253 (N_37253,N_36548,N_36694);
and U37254 (N_37254,N_36801,N_36067);
xor U37255 (N_37255,N_36864,N_36871);
nand U37256 (N_37256,N_36148,N_36315);
or U37257 (N_37257,N_36257,N_36247);
and U37258 (N_37258,N_36200,N_36578);
or U37259 (N_37259,N_36130,N_36203);
or U37260 (N_37260,N_36731,N_36745);
xor U37261 (N_37261,N_36803,N_36565);
or U37262 (N_37262,N_36765,N_36219);
or U37263 (N_37263,N_36603,N_36856);
xor U37264 (N_37264,N_36951,N_36660);
nand U37265 (N_37265,N_36063,N_36635);
nand U37266 (N_37266,N_36857,N_36353);
nand U37267 (N_37267,N_36383,N_36550);
or U37268 (N_37268,N_36297,N_36158);
nand U37269 (N_37269,N_36574,N_36191);
xor U37270 (N_37270,N_36419,N_36411);
nand U37271 (N_37271,N_36147,N_36462);
or U37272 (N_37272,N_36531,N_36838);
and U37273 (N_37273,N_36623,N_36002);
nor U37274 (N_37274,N_36642,N_36627);
and U37275 (N_37275,N_36814,N_36677);
nor U37276 (N_37276,N_36611,N_36594);
nor U37277 (N_37277,N_36339,N_36509);
xnor U37278 (N_37278,N_36583,N_36277);
or U37279 (N_37279,N_36920,N_36186);
or U37280 (N_37280,N_36590,N_36294);
nor U37281 (N_37281,N_36098,N_36154);
xnor U37282 (N_37282,N_36546,N_36418);
or U37283 (N_37283,N_36905,N_36309);
nor U37284 (N_37284,N_36300,N_36961);
xnor U37285 (N_37285,N_36965,N_36279);
or U37286 (N_37286,N_36946,N_36172);
or U37287 (N_37287,N_36645,N_36954);
or U37288 (N_37288,N_36789,N_36497);
or U37289 (N_37289,N_36855,N_36105);
and U37290 (N_37290,N_36577,N_36449);
nor U37291 (N_37291,N_36250,N_36962);
or U37292 (N_37292,N_36880,N_36183);
or U37293 (N_37293,N_36111,N_36217);
nand U37294 (N_37294,N_36000,N_36325);
nor U37295 (N_37295,N_36792,N_36636);
or U37296 (N_37296,N_36512,N_36766);
xor U37297 (N_37297,N_36464,N_36164);
nand U37298 (N_37298,N_36376,N_36138);
and U37299 (N_37299,N_36460,N_36826);
and U37300 (N_37300,N_36514,N_36945);
xor U37301 (N_37301,N_36237,N_36669);
nand U37302 (N_37302,N_36899,N_36420);
nor U37303 (N_37303,N_36210,N_36551);
nor U37304 (N_37304,N_36199,N_36972);
nor U37305 (N_37305,N_36204,N_36696);
and U37306 (N_37306,N_36421,N_36566);
nor U37307 (N_37307,N_36699,N_36859);
and U37308 (N_37308,N_36837,N_36184);
nand U37309 (N_37309,N_36975,N_36310);
nor U37310 (N_37310,N_36969,N_36102);
and U37311 (N_37311,N_36807,N_36451);
nand U37312 (N_37312,N_36607,N_36941);
and U37313 (N_37313,N_36478,N_36701);
or U37314 (N_37314,N_36437,N_36263);
nand U37315 (N_37315,N_36459,N_36114);
nand U37316 (N_37316,N_36852,N_36330);
nand U37317 (N_37317,N_36267,N_36815);
nand U37318 (N_37318,N_36910,N_36841);
xnor U37319 (N_37319,N_36367,N_36532);
or U37320 (N_37320,N_36233,N_36680);
and U37321 (N_37321,N_36051,N_36974);
and U37322 (N_37322,N_36197,N_36788);
xnor U37323 (N_37323,N_36465,N_36179);
xnor U37324 (N_37324,N_36622,N_36295);
and U37325 (N_37325,N_36949,N_36274);
nand U37326 (N_37326,N_36608,N_36821);
nor U37327 (N_37327,N_36913,N_36708);
xor U37328 (N_37328,N_36634,N_36604);
and U37329 (N_37329,N_36804,N_36115);
or U37330 (N_37330,N_36403,N_36338);
xnor U37331 (N_37331,N_36466,N_36795);
and U37332 (N_37332,N_36407,N_36519);
or U37333 (N_37333,N_36264,N_36341);
or U37334 (N_37334,N_36707,N_36733);
nand U37335 (N_37335,N_36388,N_36288);
xor U37336 (N_37336,N_36408,N_36484);
or U37337 (N_37337,N_36368,N_36076);
xor U37338 (N_37338,N_36387,N_36985);
nand U37339 (N_37339,N_36334,N_36992);
nand U37340 (N_37340,N_36968,N_36433);
and U37341 (N_37341,N_36038,N_36400);
or U37342 (N_37342,N_36447,N_36013);
nand U37343 (N_37343,N_36019,N_36959);
xnor U37344 (N_37344,N_36850,N_36480);
nand U37345 (N_37345,N_36930,N_36912);
nand U37346 (N_37346,N_36549,N_36780);
and U37347 (N_37347,N_36729,N_36082);
xnor U37348 (N_37348,N_36724,N_36196);
nor U37349 (N_37349,N_36658,N_36488);
and U37350 (N_37350,N_36800,N_36595);
nor U37351 (N_37351,N_36331,N_36508);
and U37352 (N_37352,N_36071,N_36242);
xor U37353 (N_37353,N_36966,N_36171);
xor U37354 (N_37354,N_36235,N_36671);
nor U37355 (N_37355,N_36461,N_36706);
nor U37356 (N_37356,N_36417,N_36012);
nand U37357 (N_37357,N_36024,N_36676);
and U37358 (N_37358,N_36395,N_36260);
xnor U37359 (N_37359,N_36759,N_36538);
xnor U37360 (N_37360,N_36285,N_36602);
xor U37361 (N_37361,N_36180,N_36695);
or U37362 (N_37362,N_36313,N_36402);
nor U37363 (N_37363,N_36653,N_36722);
nor U37364 (N_37364,N_36328,N_36015);
and U37365 (N_37365,N_36778,N_36228);
and U37366 (N_37366,N_36697,N_36240);
xor U37367 (N_37367,N_36874,N_36535);
and U37368 (N_37368,N_36540,N_36714);
nand U37369 (N_37369,N_36842,N_36902);
and U37370 (N_37370,N_36041,N_36492);
or U37371 (N_37371,N_36280,N_36552);
xor U37372 (N_37372,N_36475,N_36981);
nand U37373 (N_37373,N_36485,N_36909);
nand U37374 (N_37374,N_36160,N_36124);
nor U37375 (N_37375,N_36365,N_36868);
xor U37376 (N_37376,N_36872,N_36187);
nor U37377 (N_37377,N_36739,N_36458);
xnor U37378 (N_37378,N_36748,N_36457);
or U37379 (N_37379,N_36625,N_36736);
and U37380 (N_37380,N_36927,N_36554);
nand U37381 (N_37381,N_36149,N_36589);
nand U37382 (N_37382,N_36030,N_36557);
and U37383 (N_37383,N_36691,N_36225);
nor U37384 (N_37384,N_36001,N_36719);
nor U37385 (N_37385,N_36940,N_36081);
and U37386 (N_37386,N_36839,N_36468);
or U37387 (N_37387,N_36561,N_36404);
and U37388 (N_37388,N_36702,N_36346);
nor U37389 (N_37389,N_36046,N_36753);
or U37390 (N_37390,N_36537,N_36996);
or U37391 (N_37391,N_36710,N_36428);
and U37392 (N_37392,N_36883,N_36630);
nand U37393 (N_37393,N_36027,N_36919);
and U37394 (N_37394,N_36786,N_36568);
xnor U37395 (N_37395,N_36506,N_36021);
xnor U37396 (N_37396,N_36342,N_36453);
xnor U37397 (N_37397,N_36406,N_36432);
and U37398 (N_37398,N_36948,N_36775);
nor U37399 (N_37399,N_36022,N_36193);
nor U37400 (N_37400,N_36615,N_36053);
xor U37401 (N_37401,N_36988,N_36359);
xor U37402 (N_37402,N_36840,N_36846);
nor U37403 (N_37403,N_36133,N_36749);
xnor U37404 (N_37404,N_36132,N_36963);
or U37405 (N_37405,N_36317,N_36306);
nand U37406 (N_37406,N_36320,N_36126);
nor U37407 (N_37407,N_36055,N_36742);
xnor U37408 (N_37408,N_36156,N_36104);
nand U37409 (N_37409,N_36770,N_36878);
nand U37410 (N_37410,N_36127,N_36763);
nand U37411 (N_37411,N_36953,N_36794);
and U37412 (N_37412,N_36991,N_36703);
or U37413 (N_37413,N_36643,N_36416);
and U37414 (N_37414,N_36732,N_36687);
nor U37415 (N_37415,N_36438,N_36811);
and U37416 (N_37416,N_36752,N_36454);
nor U37417 (N_37417,N_36870,N_36626);
nor U37418 (N_37418,N_36713,N_36576);
nor U37419 (N_37419,N_36118,N_36879);
xor U37420 (N_37420,N_36921,N_36392);
or U37421 (N_37421,N_36174,N_36096);
nor U37422 (N_37422,N_36727,N_36579);
xor U37423 (N_37423,N_36516,N_36333);
or U37424 (N_37424,N_36039,N_36207);
nand U37425 (N_37425,N_36667,N_36932);
nand U37426 (N_37426,N_36555,N_36712);
nand U37427 (N_37427,N_36391,N_36935);
xor U37428 (N_37428,N_36239,N_36922);
nor U37429 (N_37429,N_36471,N_36069);
nor U37430 (N_37430,N_36600,N_36271);
or U37431 (N_37431,N_36238,N_36947);
xnor U37432 (N_37432,N_36998,N_36648);
and U37433 (N_37433,N_36425,N_36372);
nor U37434 (N_37434,N_36286,N_36381);
or U37435 (N_37435,N_36572,N_36926);
and U37436 (N_37436,N_36370,N_36553);
or U37437 (N_37437,N_36089,N_36906);
xor U37438 (N_37438,N_36612,N_36231);
nand U37439 (N_37439,N_36754,N_36361);
and U37440 (N_37440,N_36586,N_36891);
nand U37441 (N_37441,N_36746,N_36059);
xor U37442 (N_37442,N_36351,N_36895);
nand U37443 (N_37443,N_36246,N_36751);
and U37444 (N_37444,N_36606,N_36757);
xor U37445 (N_37445,N_36094,N_36324);
nor U37446 (N_37446,N_36640,N_36314);
nand U37447 (N_37447,N_36618,N_36844);
or U37448 (N_37448,N_36050,N_36033);
nor U37449 (N_37449,N_36423,N_36629);
nand U37450 (N_37450,N_36398,N_36785);
nand U37451 (N_37451,N_36167,N_36591);
or U37452 (N_37452,N_36542,N_36145);
and U37453 (N_37453,N_36254,N_36681);
or U37454 (N_37454,N_36898,N_36666);
and U37455 (N_37455,N_36507,N_36031);
nor U37456 (N_37456,N_36518,N_36074);
nand U37457 (N_37457,N_36006,N_36783);
or U37458 (N_37458,N_36918,N_36061);
and U37459 (N_37459,N_36010,N_36582);
or U37460 (N_37460,N_36588,N_36511);
nand U37461 (N_37461,N_36140,N_36396);
xnor U37462 (N_37462,N_36533,N_36806);
and U37463 (N_37463,N_36463,N_36208);
nand U37464 (N_37464,N_36202,N_36755);
nand U37465 (N_37465,N_36657,N_36735);
or U37466 (N_37466,N_36211,N_36493);
nor U37467 (N_37467,N_36258,N_36176);
nor U37468 (N_37468,N_36473,N_36095);
nand U37469 (N_37469,N_36851,N_36058);
xnor U37470 (N_37470,N_36928,N_36831);
nor U37471 (N_37471,N_36393,N_36415);
or U37472 (N_37472,N_36632,N_36450);
and U37473 (N_37473,N_36889,N_36813);
xor U37474 (N_37474,N_36624,N_36790);
or U37475 (N_37475,N_36117,N_36711);
and U37476 (N_37476,N_36188,N_36980);
xor U37477 (N_37477,N_36113,N_36989);
or U37478 (N_37478,N_36614,N_36175);
or U37479 (N_37479,N_36123,N_36747);
nor U37480 (N_37480,N_36651,N_36938);
and U37481 (N_37481,N_36378,N_36318);
nand U37482 (N_37482,N_36698,N_36885);
or U37483 (N_37483,N_36573,N_36929);
and U37484 (N_37484,N_36245,N_36750);
xnor U37485 (N_37485,N_36740,N_36720);
or U37486 (N_37486,N_36243,N_36360);
nor U37487 (N_37487,N_36575,N_36762);
xor U37488 (N_37488,N_36843,N_36080);
xor U37489 (N_37489,N_36054,N_36152);
or U37490 (N_37490,N_36222,N_36108);
or U37491 (N_37491,N_36756,N_36431);
or U37492 (N_37492,N_36173,N_36610);
and U37493 (N_37493,N_36029,N_36662);
or U37494 (N_37494,N_36580,N_36249);
xor U37495 (N_37495,N_36689,N_36654);
nor U37496 (N_37496,N_36261,N_36201);
or U37497 (N_37497,N_36958,N_36377);
xnor U37498 (N_37498,N_36092,N_36743);
nor U37499 (N_37499,N_36139,N_36016);
or U37500 (N_37500,N_36716,N_36804);
nor U37501 (N_37501,N_36316,N_36060);
nand U37502 (N_37502,N_36205,N_36450);
nor U37503 (N_37503,N_36389,N_36247);
and U37504 (N_37504,N_36316,N_36351);
or U37505 (N_37505,N_36671,N_36340);
nor U37506 (N_37506,N_36124,N_36199);
and U37507 (N_37507,N_36990,N_36628);
and U37508 (N_37508,N_36268,N_36049);
nor U37509 (N_37509,N_36539,N_36357);
or U37510 (N_37510,N_36110,N_36360);
nand U37511 (N_37511,N_36803,N_36901);
nor U37512 (N_37512,N_36293,N_36383);
xor U37513 (N_37513,N_36841,N_36653);
nor U37514 (N_37514,N_36391,N_36064);
or U37515 (N_37515,N_36054,N_36139);
and U37516 (N_37516,N_36712,N_36393);
nor U37517 (N_37517,N_36877,N_36175);
or U37518 (N_37518,N_36708,N_36891);
nor U37519 (N_37519,N_36826,N_36289);
and U37520 (N_37520,N_36309,N_36852);
and U37521 (N_37521,N_36310,N_36117);
nor U37522 (N_37522,N_36903,N_36204);
nand U37523 (N_37523,N_36481,N_36762);
or U37524 (N_37524,N_36225,N_36492);
nor U37525 (N_37525,N_36652,N_36164);
nand U37526 (N_37526,N_36638,N_36313);
xnor U37527 (N_37527,N_36698,N_36233);
xnor U37528 (N_37528,N_36445,N_36177);
xnor U37529 (N_37529,N_36621,N_36405);
nand U37530 (N_37530,N_36260,N_36910);
and U37531 (N_37531,N_36395,N_36985);
or U37532 (N_37532,N_36845,N_36736);
or U37533 (N_37533,N_36365,N_36907);
xnor U37534 (N_37534,N_36940,N_36041);
nor U37535 (N_37535,N_36673,N_36060);
or U37536 (N_37536,N_36666,N_36538);
xnor U37537 (N_37537,N_36266,N_36037);
xnor U37538 (N_37538,N_36040,N_36117);
and U37539 (N_37539,N_36164,N_36928);
and U37540 (N_37540,N_36804,N_36183);
and U37541 (N_37541,N_36802,N_36772);
xnor U37542 (N_37542,N_36955,N_36710);
and U37543 (N_37543,N_36920,N_36101);
nand U37544 (N_37544,N_36014,N_36508);
xnor U37545 (N_37545,N_36212,N_36753);
nand U37546 (N_37546,N_36678,N_36576);
xnor U37547 (N_37547,N_36442,N_36565);
and U37548 (N_37548,N_36883,N_36879);
or U37549 (N_37549,N_36462,N_36918);
nand U37550 (N_37550,N_36710,N_36268);
and U37551 (N_37551,N_36474,N_36633);
or U37552 (N_37552,N_36910,N_36576);
nor U37553 (N_37553,N_36457,N_36361);
nor U37554 (N_37554,N_36287,N_36049);
and U37555 (N_37555,N_36170,N_36491);
or U37556 (N_37556,N_36968,N_36888);
or U37557 (N_37557,N_36601,N_36357);
nor U37558 (N_37558,N_36751,N_36332);
nand U37559 (N_37559,N_36544,N_36251);
nand U37560 (N_37560,N_36866,N_36033);
xnor U37561 (N_37561,N_36219,N_36490);
xor U37562 (N_37562,N_36766,N_36013);
nand U37563 (N_37563,N_36091,N_36997);
and U37564 (N_37564,N_36142,N_36742);
nand U37565 (N_37565,N_36409,N_36732);
nor U37566 (N_37566,N_36104,N_36972);
or U37567 (N_37567,N_36545,N_36855);
and U37568 (N_37568,N_36731,N_36490);
nand U37569 (N_37569,N_36855,N_36322);
nand U37570 (N_37570,N_36634,N_36966);
and U37571 (N_37571,N_36841,N_36695);
or U37572 (N_37572,N_36552,N_36329);
nand U37573 (N_37573,N_36663,N_36053);
nor U37574 (N_37574,N_36812,N_36646);
nand U37575 (N_37575,N_36581,N_36415);
xor U37576 (N_37576,N_36476,N_36924);
nand U37577 (N_37577,N_36225,N_36136);
or U37578 (N_37578,N_36785,N_36086);
nand U37579 (N_37579,N_36397,N_36940);
xor U37580 (N_37580,N_36510,N_36953);
xnor U37581 (N_37581,N_36184,N_36149);
nor U37582 (N_37582,N_36741,N_36094);
and U37583 (N_37583,N_36290,N_36324);
xnor U37584 (N_37584,N_36178,N_36951);
or U37585 (N_37585,N_36865,N_36075);
nor U37586 (N_37586,N_36455,N_36579);
or U37587 (N_37587,N_36669,N_36811);
nand U37588 (N_37588,N_36099,N_36001);
or U37589 (N_37589,N_36456,N_36740);
nor U37590 (N_37590,N_36315,N_36371);
nand U37591 (N_37591,N_36085,N_36475);
nor U37592 (N_37592,N_36277,N_36336);
and U37593 (N_37593,N_36688,N_36534);
nand U37594 (N_37594,N_36866,N_36465);
and U37595 (N_37595,N_36543,N_36374);
and U37596 (N_37596,N_36569,N_36332);
nor U37597 (N_37597,N_36656,N_36867);
xor U37598 (N_37598,N_36646,N_36713);
xor U37599 (N_37599,N_36090,N_36449);
xnor U37600 (N_37600,N_36391,N_36536);
nor U37601 (N_37601,N_36979,N_36440);
or U37602 (N_37602,N_36518,N_36728);
and U37603 (N_37603,N_36738,N_36636);
xnor U37604 (N_37604,N_36521,N_36810);
or U37605 (N_37605,N_36267,N_36717);
or U37606 (N_37606,N_36818,N_36382);
xor U37607 (N_37607,N_36328,N_36290);
xor U37608 (N_37608,N_36272,N_36241);
nand U37609 (N_37609,N_36969,N_36133);
nand U37610 (N_37610,N_36081,N_36571);
and U37611 (N_37611,N_36479,N_36358);
xor U37612 (N_37612,N_36134,N_36115);
xnor U37613 (N_37613,N_36992,N_36776);
nand U37614 (N_37614,N_36395,N_36425);
and U37615 (N_37615,N_36590,N_36472);
and U37616 (N_37616,N_36912,N_36024);
and U37617 (N_37617,N_36503,N_36578);
xnor U37618 (N_37618,N_36374,N_36220);
or U37619 (N_37619,N_36147,N_36970);
nor U37620 (N_37620,N_36694,N_36538);
nor U37621 (N_37621,N_36342,N_36885);
or U37622 (N_37622,N_36660,N_36511);
and U37623 (N_37623,N_36837,N_36428);
or U37624 (N_37624,N_36547,N_36055);
nand U37625 (N_37625,N_36416,N_36484);
and U37626 (N_37626,N_36125,N_36877);
nand U37627 (N_37627,N_36433,N_36497);
nor U37628 (N_37628,N_36934,N_36657);
nor U37629 (N_37629,N_36264,N_36343);
or U37630 (N_37630,N_36156,N_36632);
nand U37631 (N_37631,N_36736,N_36628);
nand U37632 (N_37632,N_36661,N_36908);
and U37633 (N_37633,N_36797,N_36937);
xor U37634 (N_37634,N_36812,N_36295);
xor U37635 (N_37635,N_36819,N_36994);
nand U37636 (N_37636,N_36142,N_36091);
or U37637 (N_37637,N_36077,N_36488);
nand U37638 (N_37638,N_36189,N_36198);
nor U37639 (N_37639,N_36782,N_36522);
nor U37640 (N_37640,N_36414,N_36535);
nand U37641 (N_37641,N_36414,N_36155);
and U37642 (N_37642,N_36816,N_36617);
xnor U37643 (N_37643,N_36646,N_36373);
or U37644 (N_37644,N_36478,N_36120);
nor U37645 (N_37645,N_36453,N_36569);
nand U37646 (N_37646,N_36023,N_36127);
and U37647 (N_37647,N_36033,N_36689);
and U37648 (N_37648,N_36904,N_36956);
or U37649 (N_37649,N_36768,N_36659);
nand U37650 (N_37650,N_36412,N_36785);
nand U37651 (N_37651,N_36584,N_36472);
nand U37652 (N_37652,N_36485,N_36271);
nand U37653 (N_37653,N_36159,N_36545);
or U37654 (N_37654,N_36362,N_36725);
xnor U37655 (N_37655,N_36954,N_36417);
and U37656 (N_37656,N_36916,N_36691);
nand U37657 (N_37657,N_36747,N_36873);
xor U37658 (N_37658,N_36914,N_36602);
nor U37659 (N_37659,N_36874,N_36573);
nand U37660 (N_37660,N_36121,N_36400);
or U37661 (N_37661,N_36029,N_36371);
and U37662 (N_37662,N_36449,N_36648);
nor U37663 (N_37663,N_36013,N_36272);
or U37664 (N_37664,N_36168,N_36833);
xnor U37665 (N_37665,N_36350,N_36482);
or U37666 (N_37666,N_36441,N_36367);
or U37667 (N_37667,N_36013,N_36893);
nor U37668 (N_37668,N_36691,N_36704);
xnor U37669 (N_37669,N_36721,N_36159);
or U37670 (N_37670,N_36127,N_36312);
and U37671 (N_37671,N_36671,N_36833);
xor U37672 (N_37672,N_36844,N_36099);
or U37673 (N_37673,N_36652,N_36429);
and U37674 (N_37674,N_36044,N_36993);
nor U37675 (N_37675,N_36225,N_36658);
or U37676 (N_37676,N_36187,N_36959);
or U37677 (N_37677,N_36345,N_36928);
and U37678 (N_37678,N_36774,N_36650);
nor U37679 (N_37679,N_36003,N_36123);
nor U37680 (N_37680,N_36141,N_36302);
xor U37681 (N_37681,N_36092,N_36864);
nor U37682 (N_37682,N_36053,N_36135);
xnor U37683 (N_37683,N_36037,N_36617);
nand U37684 (N_37684,N_36570,N_36055);
and U37685 (N_37685,N_36047,N_36653);
xnor U37686 (N_37686,N_36720,N_36738);
nor U37687 (N_37687,N_36201,N_36906);
nand U37688 (N_37688,N_36394,N_36112);
and U37689 (N_37689,N_36501,N_36840);
nand U37690 (N_37690,N_36035,N_36553);
xor U37691 (N_37691,N_36179,N_36803);
nand U37692 (N_37692,N_36654,N_36294);
nor U37693 (N_37693,N_36205,N_36822);
nor U37694 (N_37694,N_36231,N_36239);
nand U37695 (N_37695,N_36376,N_36073);
or U37696 (N_37696,N_36994,N_36721);
or U37697 (N_37697,N_36331,N_36330);
xor U37698 (N_37698,N_36061,N_36916);
nor U37699 (N_37699,N_36868,N_36001);
xnor U37700 (N_37700,N_36403,N_36846);
nor U37701 (N_37701,N_36786,N_36231);
and U37702 (N_37702,N_36554,N_36545);
xnor U37703 (N_37703,N_36001,N_36807);
or U37704 (N_37704,N_36349,N_36000);
and U37705 (N_37705,N_36468,N_36380);
or U37706 (N_37706,N_36870,N_36824);
or U37707 (N_37707,N_36218,N_36132);
and U37708 (N_37708,N_36602,N_36981);
or U37709 (N_37709,N_36537,N_36640);
or U37710 (N_37710,N_36385,N_36104);
and U37711 (N_37711,N_36062,N_36628);
xnor U37712 (N_37712,N_36169,N_36764);
and U37713 (N_37713,N_36348,N_36565);
nor U37714 (N_37714,N_36336,N_36422);
or U37715 (N_37715,N_36417,N_36549);
nand U37716 (N_37716,N_36997,N_36057);
or U37717 (N_37717,N_36034,N_36389);
or U37718 (N_37718,N_36962,N_36109);
or U37719 (N_37719,N_36927,N_36769);
xnor U37720 (N_37720,N_36220,N_36502);
and U37721 (N_37721,N_36073,N_36118);
and U37722 (N_37722,N_36855,N_36430);
nor U37723 (N_37723,N_36002,N_36669);
xor U37724 (N_37724,N_36606,N_36163);
nor U37725 (N_37725,N_36112,N_36345);
nor U37726 (N_37726,N_36651,N_36957);
and U37727 (N_37727,N_36404,N_36787);
and U37728 (N_37728,N_36090,N_36491);
xor U37729 (N_37729,N_36707,N_36167);
and U37730 (N_37730,N_36362,N_36747);
and U37731 (N_37731,N_36801,N_36536);
nand U37732 (N_37732,N_36266,N_36554);
xnor U37733 (N_37733,N_36147,N_36277);
nand U37734 (N_37734,N_36841,N_36949);
nor U37735 (N_37735,N_36973,N_36635);
xnor U37736 (N_37736,N_36307,N_36448);
and U37737 (N_37737,N_36447,N_36640);
or U37738 (N_37738,N_36222,N_36355);
and U37739 (N_37739,N_36934,N_36875);
nor U37740 (N_37740,N_36339,N_36766);
xor U37741 (N_37741,N_36587,N_36100);
and U37742 (N_37742,N_36395,N_36797);
and U37743 (N_37743,N_36656,N_36081);
nand U37744 (N_37744,N_36107,N_36944);
nand U37745 (N_37745,N_36133,N_36653);
xor U37746 (N_37746,N_36083,N_36295);
or U37747 (N_37747,N_36967,N_36296);
xor U37748 (N_37748,N_36763,N_36207);
or U37749 (N_37749,N_36206,N_36759);
and U37750 (N_37750,N_36687,N_36908);
or U37751 (N_37751,N_36845,N_36599);
xor U37752 (N_37752,N_36405,N_36947);
nor U37753 (N_37753,N_36634,N_36435);
and U37754 (N_37754,N_36530,N_36156);
nor U37755 (N_37755,N_36919,N_36036);
or U37756 (N_37756,N_36031,N_36063);
nor U37757 (N_37757,N_36187,N_36312);
or U37758 (N_37758,N_36463,N_36042);
or U37759 (N_37759,N_36813,N_36700);
nand U37760 (N_37760,N_36314,N_36892);
or U37761 (N_37761,N_36215,N_36760);
and U37762 (N_37762,N_36104,N_36061);
xor U37763 (N_37763,N_36361,N_36764);
nor U37764 (N_37764,N_36276,N_36167);
nor U37765 (N_37765,N_36931,N_36271);
and U37766 (N_37766,N_36260,N_36960);
or U37767 (N_37767,N_36827,N_36807);
nand U37768 (N_37768,N_36355,N_36104);
nor U37769 (N_37769,N_36228,N_36907);
and U37770 (N_37770,N_36709,N_36631);
nand U37771 (N_37771,N_36497,N_36348);
nor U37772 (N_37772,N_36335,N_36406);
nand U37773 (N_37773,N_36577,N_36953);
or U37774 (N_37774,N_36198,N_36300);
and U37775 (N_37775,N_36352,N_36620);
nand U37776 (N_37776,N_36137,N_36221);
xor U37777 (N_37777,N_36773,N_36044);
xor U37778 (N_37778,N_36408,N_36304);
and U37779 (N_37779,N_36839,N_36695);
or U37780 (N_37780,N_36533,N_36090);
xor U37781 (N_37781,N_36861,N_36295);
nand U37782 (N_37782,N_36039,N_36795);
nor U37783 (N_37783,N_36196,N_36564);
xor U37784 (N_37784,N_36918,N_36076);
or U37785 (N_37785,N_36344,N_36785);
or U37786 (N_37786,N_36898,N_36510);
nand U37787 (N_37787,N_36000,N_36743);
xor U37788 (N_37788,N_36217,N_36941);
nand U37789 (N_37789,N_36484,N_36653);
nand U37790 (N_37790,N_36253,N_36271);
or U37791 (N_37791,N_36957,N_36395);
or U37792 (N_37792,N_36218,N_36139);
and U37793 (N_37793,N_36038,N_36390);
nand U37794 (N_37794,N_36649,N_36738);
nand U37795 (N_37795,N_36457,N_36772);
xnor U37796 (N_37796,N_36289,N_36120);
nand U37797 (N_37797,N_36461,N_36530);
xnor U37798 (N_37798,N_36628,N_36624);
or U37799 (N_37799,N_36821,N_36887);
and U37800 (N_37800,N_36441,N_36089);
and U37801 (N_37801,N_36111,N_36348);
and U37802 (N_37802,N_36255,N_36838);
nor U37803 (N_37803,N_36468,N_36404);
and U37804 (N_37804,N_36773,N_36903);
nand U37805 (N_37805,N_36740,N_36641);
xnor U37806 (N_37806,N_36698,N_36214);
nand U37807 (N_37807,N_36514,N_36258);
xor U37808 (N_37808,N_36647,N_36683);
nor U37809 (N_37809,N_36787,N_36854);
xnor U37810 (N_37810,N_36068,N_36281);
or U37811 (N_37811,N_36924,N_36073);
xor U37812 (N_37812,N_36521,N_36654);
and U37813 (N_37813,N_36745,N_36497);
nor U37814 (N_37814,N_36007,N_36361);
nor U37815 (N_37815,N_36810,N_36036);
xor U37816 (N_37816,N_36873,N_36193);
and U37817 (N_37817,N_36044,N_36772);
nand U37818 (N_37818,N_36371,N_36349);
and U37819 (N_37819,N_36527,N_36045);
xor U37820 (N_37820,N_36521,N_36258);
xor U37821 (N_37821,N_36001,N_36206);
nand U37822 (N_37822,N_36157,N_36194);
nand U37823 (N_37823,N_36069,N_36506);
xor U37824 (N_37824,N_36702,N_36942);
nand U37825 (N_37825,N_36395,N_36579);
xnor U37826 (N_37826,N_36892,N_36012);
and U37827 (N_37827,N_36174,N_36549);
nor U37828 (N_37828,N_36593,N_36950);
xnor U37829 (N_37829,N_36611,N_36675);
xnor U37830 (N_37830,N_36849,N_36838);
or U37831 (N_37831,N_36734,N_36170);
and U37832 (N_37832,N_36637,N_36716);
and U37833 (N_37833,N_36018,N_36461);
or U37834 (N_37834,N_36887,N_36702);
or U37835 (N_37835,N_36649,N_36088);
and U37836 (N_37836,N_36205,N_36180);
nand U37837 (N_37837,N_36078,N_36948);
nor U37838 (N_37838,N_36145,N_36010);
nor U37839 (N_37839,N_36512,N_36698);
nand U37840 (N_37840,N_36595,N_36226);
nand U37841 (N_37841,N_36043,N_36995);
nor U37842 (N_37842,N_36892,N_36482);
nand U37843 (N_37843,N_36796,N_36842);
or U37844 (N_37844,N_36558,N_36263);
nor U37845 (N_37845,N_36718,N_36121);
nand U37846 (N_37846,N_36466,N_36596);
and U37847 (N_37847,N_36037,N_36114);
and U37848 (N_37848,N_36801,N_36469);
or U37849 (N_37849,N_36571,N_36274);
xnor U37850 (N_37850,N_36524,N_36044);
or U37851 (N_37851,N_36765,N_36393);
or U37852 (N_37852,N_36363,N_36999);
xnor U37853 (N_37853,N_36957,N_36875);
nor U37854 (N_37854,N_36735,N_36559);
nand U37855 (N_37855,N_36773,N_36373);
or U37856 (N_37856,N_36761,N_36741);
and U37857 (N_37857,N_36565,N_36748);
nand U37858 (N_37858,N_36184,N_36312);
nand U37859 (N_37859,N_36329,N_36462);
and U37860 (N_37860,N_36726,N_36899);
nand U37861 (N_37861,N_36815,N_36773);
xor U37862 (N_37862,N_36303,N_36423);
and U37863 (N_37863,N_36450,N_36144);
nand U37864 (N_37864,N_36567,N_36019);
nand U37865 (N_37865,N_36684,N_36696);
nor U37866 (N_37866,N_36269,N_36349);
nor U37867 (N_37867,N_36361,N_36423);
or U37868 (N_37868,N_36077,N_36506);
nand U37869 (N_37869,N_36269,N_36403);
and U37870 (N_37870,N_36018,N_36623);
nand U37871 (N_37871,N_36227,N_36266);
or U37872 (N_37872,N_36283,N_36043);
and U37873 (N_37873,N_36409,N_36302);
xor U37874 (N_37874,N_36107,N_36252);
or U37875 (N_37875,N_36165,N_36433);
and U37876 (N_37876,N_36481,N_36968);
nand U37877 (N_37877,N_36127,N_36809);
xnor U37878 (N_37878,N_36707,N_36385);
nor U37879 (N_37879,N_36722,N_36944);
and U37880 (N_37880,N_36398,N_36410);
or U37881 (N_37881,N_36872,N_36272);
or U37882 (N_37882,N_36846,N_36746);
xor U37883 (N_37883,N_36650,N_36152);
nand U37884 (N_37884,N_36582,N_36387);
or U37885 (N_37885,N_36073,N_36359);
or U37886 (N_37886,N_36326,N_36713);
and U37887 (N_37887,N_36483,N_36695);
xnor U37888 (N_37888,N_36726,N_36178);
and U37889 (N_37889,N_36544,N_36223);
xnor U37890 (N_37890,N_36774,N_36133);
and U37891 (N_37891,N_36985,N_36753);
nand U37892 (N_37892,N_36320,N_36452);
or U37893 (N_37893,N_36401,N_36806);
nor U37894 (N_37894,N_36504,N_36482);
nor U37895 (N_37895,N_36532,N_36473);
nor U37896 (N_37896,N_36616,N_36046);
xnor U37897 (N_37897,N_36951,N_36174);
and U37898 (N_37898,N_36760,N_36183);
and U37899 (N_37899,N_36133,N_36915);
xor U37900 (N_37900,N_36205,N_36547);
and U37901 (N_37901,N_36925,N_36764);
nand U37902 (N_37902,N_36118,N_36275);
and U37903 (N_37903,N_36129,N_36011);
nand U37904 (N_37904,N_36757,N_36334);
nand U37905 (N_37905,N_36083,N_36812);
or U37906 (N_37906,N_36080,N_36086);
nor U37907 (N_37907,N_36655,N_36162);
xnor U37908 (N_37908,N_36609,N_36940);
xnor U37909 (N_37909,N_36208,N_36821);
and U37910 (N_37910,N_36706,N_36532);
or U37911 (N_37911,N_36482,N_36050);
xnor U37912 (N_37912,N_36937,N_36777);
and U37913 (N_37913,N_36570,N_36670);
nand U37914 (N_37914,N_36328,N_36299);
and U37915 (N_37915,N_36341,N_36014);
or U37916 (N_37916,N_36506,N_36414);
xnor U37917 (N_37917,N_36521,N_36550);
nand U37918 (N_37918,N_36332,N_36888);
nor U37919 (N_37919,N_36744,N_36529);
or U37920 (N_37920,N_36464,N_36380);
xnor U37921 (N_37921,N_36641,N_36613);
and U37922 (N_37922,N_36021,N_36545);
xor U37923 (N_37923,N_36698,N_36309);
and U37924 (N_37924,N_36024,N_36643);
xnor U37925 (N_37925,N_36713,N_36278);
and U37926 (N_37926,N_36536,N_36338);
and U37927 (N_37927,N_36090,N_36653);
nand U37928 (N_37928,N_36290,N_36869);
nor U37929 (N_37929,N_36259,N_36017);
nand U37930 (N_37930,N_36948,N_36706);
or U37931 (N_37931,N_36752,N_36920);
or U37932 (N_37932,N_36425,N_36276);
or U37933 (N_37933,N_36386,N_36875);
xnor U37934 (N_37934,N_36023,N_36148);
nand U37935 (N_37935,N_36146,N_36440);
and U37936 (N_37936,N_36714,N_36864);
nand U37937 (N_37937,N_36435,N_36055);
or U37938 (N_37938,N_36103,N_36321);
nand U37939 (N_37939,N_36427,N_36638);
xnor U37940 (N_37940,N_36402,N_36252);
and U37941 (N_37941,N_36121,N_36916);
xnor U37942 (N_37942,N_36154,N_36424);
or U37943 (N_37943,N_36474,N_36433);
xor U37944 (N_37944,N_36713,N_36786);
nor U37945 (N_37945,N_36035,N_36292);
xnor U37946 (N_37946,N_36531,N_36652);
nand U37947 (N_37947,N_36708,N_36093);
and U37948 (N_37948,N_36820,N_36496);
xor U37949 (N_37949,N_36480,N_36595);
or U37950 (N_37950,N_36247,N_36476);
nand U37951 (N_37951,N_36054,N_36385);
nor U37952 (N_37952,N_36265,N_36305);
nand U37953 (N_37953,N_36626,N_36812);
or U37954 (N_37954,N_36182,N_36779);
nand U37955 (N_37955,N_36217,N_36819);
nand U37956 (N_37956,N_36506,N_36350);
nor U37957 (N_37957,N_36700,N_36594);
nand U37958 (N_37958,N_36389,N_36662);
xor U37959 (N_37959,N_36960,N_36771);
nor U37960 (N_37960,N_36086,N_36355);
nand U37961 (N_37961,N_36955,N_36401);
and U37962 (N_37962,N_36435,N_36772);
nor U37963 (N_37963,N_36620,N_36622);
and U37964 (N_37964,N_36494,N_36872);
and U37965 (N_37965,N_36985,N_36038);
nand U37966 (N_37966,N_36082,N_36001);
xor U37967 (N_37967,N_36448,N_36571);
xor U37968 (N_37968,N_36534,N_36332);
xor U37969 (N_37969,N_36375,N_36345);
xor U37970 (N_37970,N_36348,N_36224);
or U37971 (N_37971,N_36207,N_36812);
or U37972 (N_37972,N_36749,N_36379);
nand U37973 (N_37973,N_36898,N_36632);
or U37974 (N_37974,N_36687,N_36747);
nor U37975 (N_37975,N_36056,N_36706);
nor U37976 (N_37976,N_36439,N_36090);
nor U37977 (N_37977,N_36756,N_36175);
nor U37978 (N_37978,N_36700,N_36893);
nor U37979 (N_37979,N_36179,N_36842);
or U37980 (N_37980,N_36254,N_36857);
xor U37981 (N_37981,N_36625,N_36154);
or U37982 (N_37982,N_36602,N_36833);
nand U37983 (N_37983,N_36095,N_36216);
nor U37984 (N_37984,N_36861,N_36254);
nor U37985 (N_37985,N_36498,N_36602);
xor U37986 (N_37986,N_36234,N_36599);
nand U37987 (N_37987,N_36310,N_36716);
or U37988 (N_37988,N_36610,N_36648);
nand U37989 (N_37989,N_36843,N_36202);
xnor U37990 (N_37990,N_36981,N_36689);
nor U37991 (N_37991,N_36035,N_36872);
nand U37992 (N_37992,N_36845,N_36079);
xor U37993 (N_37993,N_36292,N_36606);
xor U37994 (N_37994,N_36772,N_36997);
and U37995 (N_37995,N_36145,N_36266);
xor U37996 (N_37996,N_36012,N_36254);
and U37997 (N_37997,N_36130,N_36806);
and U37998 (N_37998,N_36054,N_36680);
nor U37999 (N_37999,N_36837,N_36533);
xor U38000 (N_38000,N_37127,N_37817);
and U38001 (N_38001,N_37257,N_37727);
and U38002 (N_38002,N_37442,N_37347);
or U38003 (N_38003,N_37646,N_37688);
or U38004 (N_38004,N_37224,N_37937);
nand U38005 (N_38005,N_37046,N_37306);
and U38006 (N_38006,N_37865,N_37896);
xnor U38007 (N_38007,N_37636,N_37664);
nor U38008 (N_38008,N_37287,N_37707);
or U38009 (N_38009,N_37831,N_37209);
nor U38010 (N_38010,N_37634,N_37648);
xor U38011 (N_38011,N_37551,N_37457);
nor U38012 (N_38012,N_37732,N_37972);
nor U38013 (N_38013,N_37004,N_37180);
or U38014 (N_38014,N_37050,N_37542);
or U38015 (N_38015,N_37844,N_37168);
nor U38016 (N_38016,N_37757,N_37230);
nand U38017 (N_38017,N_37850,N_37008);
xor U38018 (N_38018,N_37875,N_37156);
xor U38019 (N_38019,N_37995,N_37369);
xor U38020 (N_38020,N_37419,N_37091);
nand U38021 (N_38021,N_37205,N_37760);
nand U38022 (N_38022,N_37506,N_37137);
xnor U38023 (N_38023,N_37181,N_37093);
or U38024 (N_38024,N_37649,N_37497);
and U38025 (N_38025,N_37984,N_37809);
nand U38026 (N_38026,N_37019,N_37170);
and U38027 (N_38027,N_37924,N_37283);
or U38028 (N_38028,N_37228,N_37679);
and U38029 (N_38029,N_37612,N_37053);
and U38030 (N_38030,N_37808,N_37343);
xor U38031 (N_38031,N_37864,N_37070);
xnor U38032 (N_38032,N_37201,N_37239);
nand U38033 (N_38033,N_37951,N_37481);
nand U38034 (N_38034,N_37938,N_37988);
nor U38035 (N_38035,N_37321,N_37929);
nor U38036 (N_38036,N_37952,N_37790);
or U38037 (N_38037,N_37453,N_37219);
and U38038 (N_38038,N_37811,N_37604);
and U38039 (N_38039,N_37367,N_37271);
and U38040 (N_38040,N_37121,N_37072);
nand U38041 (N_38041,N_37490,N_37444);
nand U38042 (N_38042,N_37241,N_37307);
and U38043 (N_38043,N_37392,N_37515);
xnor U38044 (N_38044,N_37778,N_37350);
or U38045 (N_38045,N_37179,N_37883);
nor U38046 (N_38046,N_37456,N_37439);
nand U38047 (N_38047,N_37701,N_37379);
or U38048 (N_38048,N_37917,N_37068);
xor U38049 (N_38049,N_37521,N_37683);
nand U38050 (N_38050,N_37142,N_37944);
or U38051 (N_38051,N_37880,N_37484);
nand U38052 (N_38052,N_37366,N_37829);
and U38053 (N_38053,N_37178,N_37527);
xor U38054 (N_38054,N_37189,N_37532);
or U38055 (N_38055,N_37736,N_37992);
and U38056 (N_38056,N_37788,N_37591);
nor U38057 (N_38057,N_37657,N_37799);
nor U38058 (N_38058,N_37730,N_37362);
nor U38059 (N_38059,N_37780,N_37772);
or U38060 (N_38060,N_37318,N_37285);
xnor U38061 (N_38061,N_37833,N_37948);
nand U38062 (N_38062,N_37061,N_37204);
or U38063 (N_38063,N_37842,N_37411);
or U38064 (N_38064,N_37196,N_37786);
nor U38065 (N_38065,N_37940,N_37403);
and U38066 (N_38066,N_37956,N_37274);
nand U38067 (N_38067,N_37432,N_37460);
nand U38068 (N_38068,N_37601,N_37489);
nand U38069 (N_38069,N_37709,N_37559);
xor U38070 (N_38070,N_37576,N_37928);
nor U38071 (N_38071,N_37609,N_37335);
nand U38072 (N_38072,N_37278,N_37867);
or U38073 (N_38073,N_37923,N_37964);
nand U38074 (N_38074,N_37085,N_37038);
xor U38075 (N_38075,N_37611,N_37578);
nor U38076 (N_38076,N_37090,N_37000);
xnor U38077 (N_38077,N_37596,N_37968);
or U38078 (N_38078,N_37024,N_37650);
nand U38079 (N_38079,N_37961,N_37686);
or U38080 (N_38080,N_37986,N_37889);
nor U38081 (N_38081,N_37037,N_37512);
and U38082 (N_38082,N_37293,N_37377);
and U38083 (N_38083,N_37710,N_37910);
and U38084 (N_38084,N_37191,N_37435);
or U38085 (N_38085,N_37821,N_37492);
xor U38086 (N_38086,N_37389,N_37603);
xnor U38087 (N_38087,N_37966,N_37304);
or U38088 (N_38088,N_37704,N_37983);
and U38089 (N_38089,N_37577,N_37644);
nand U38090 (N_38090,N_37280,N_37065);
and U38091 (N_38091,N_37147,N_37312);
or U38092 (N_38092,N_37922,N_37822);
nor U38093 (N_38093,N_37394,N_37176);
nor U38094 (N_38094,N_37141,N_37627);
nor U38095 (N_38095,N_37613,N_37438);
nand U38096 (N_38096,N_37398,N_37353);
and U38097 (N_38097,N_37508,N_37502);
nand U38098 (N_38098,N_37535,N_37186);
nand U38099 (N_38099,N_37782,N_37893);
nand U38100 (N_38100,N_37826,N_37313);
xnor U38101 (N_38101,N_37381,N_37915);
xor U38102 (N_38102,N_37395,N_37740);
xor U38103 (N_38103,N_37486,N_37214);
nand U38104 (N_38104,N_37900,N_37721);
or U38105 (N_38105,N_37668,N_37877);
or U38106 (N_38106,N_37197,N_37661);
xor U38107 (N_38107,N_37621,N_37473);
and U38108 (N_38108,N_37815,N_37400);
xor U38109 (N_38109,N_37422,N_37582);
and U38110 (N_38110,N_37546,N_37773);
nor U38111 (N_38111,N_37825,N_37076);
xnor U38112 (N_38112,N_37282,N_37054);
nand U38113 (N_38113,N_37526,N_37469);
or U38114 (N_38114,N_37265,N_37311);
nand U38115 (N_38115,N_37338,N_37588);
nand U38116 (N_38116,N_37795,N_37638);
xor U38117 (N_38117,N_37244,N_37245);
xor U38118 (N_38118,N_37056,N_37474);
nor U38119 (N_38119,N_37433,N_37305);
or U38120 (N_38120,N_37839,N_37458);
nand U38121 (N_38121,N_37441,N_37912);
nor U38122 (N_38122,N_37860,N_37423);
nor U38123 (N_38123,N_37327,N_37216);
nor U38124 (N_38124,N_37510,N_37911);
nand U38125 (N_38125,N_37530,N_37361);
nand U38126 (N_38126,N_37059,N_37269);
xnor U38127 (N_38127,N_37292,N_37409);
xor U38128 (N_38128,N_37518,N_37151);
or U38129 (N_38129,N_37349,N_37479);
nand U38130 (N_38130,N_37820,N_37404);
xnor U38131 (N_38131,N_37697,N_37619);
nand U38132 (N_38132,N_37408,N_37982);
xnor U38133 (N_38133,N_37372,N_37894);
or U38134 (N_38134,N_37027,N_37999);
nand U38135 (N_38135,N_37284,N_37602);
and U38136 (N_38136,N_37348,N_37459);
or U38137 (N_38137,N_37847,N_37035);
nor U38138 (N_38138,N_37098,N_37385);
or U38139 (N_38139,N_37776,N_37500);
xor U38140 (N_38140,N_37745,N_37317);
or U38141 (N_38141,N_37505,N_37116);
nand U38142 (N_38142,N_37913,N_37213);
and U38143 (N_38143,N_37364,N_37017);
and U38144 (N_38144,N_37887,N_37629);
or U38145 (N_38145,N_37112,N_37870);
nor U38146 (N_38146,N_37901,N_37060);
or U38147 (N_38147,N_37352,N_37837);
xor U38148 (N_38148,N_37888,N_37846);
and U38149 (N_38149,N_37451,N_37848);
and U38150 (N_38150,N_37359,N_37045);
and U38151 (N_38151,N_37762,N_37718);
and U38152 (N_38152,N_37957,N_37803);
xnor U38153 (N_38153,N_37885,N_37371);
or U38154 (N_38154,N_37002,N_37029);
xnor U38155 (N_38155,N_37009,N_37715);
xnor U38156 (N_38156,N_37726,N_37162);
nor U38157 (N_38157,N_37339,N_37712);
nor U38158 (N_38158,N_37699,N_37491);
nand U38159 (N_38159,N_37775,N_37391);
or U38160 (N_38160,N_37332,N_37614);
or U38161 (N_38161,N_37063,N_37696);
and U38162 (N_38162,N_37291,N_37493);
nor U38163 (N_38163,N_37028,N_37084);
or U38164 (N_38164,N_37096,N_37495);
xor U38165 (N_38165,N_37014,N_37674);
and U38166 (N_38166,N_37855,N_37628);
xor U38167 (N_38167,N_37568,N_37416);
nand U38168 (N_38168,N_37044,N_37080);
nor U38169 (N_38169,N_37520,N_37851);
nand U38170 (N_38170,N_37597,N_37804);
and U38171 (N_38171,N_37909,N_37461);
and U38172 (N_38172,N_37570,N_37583);
nand U38173 (N_38173,N_37079,N_37333);
nor U38174 (N_38174,N_37529,N_37058);
nor U38175 (N_38175,N_37471,N_37711);
nor U38176 (N_38176,N_37823,N_37088);
or U38177 (N_38177,N_37286,N_37368);
and U38178 (N_38178,N_37933,N_37669);
nor U38179 (N_38179,N_37810,N_37415);
nand U38180 (N_38180,N_37902,N_37914);
nand U38181 (N_38181,N_37086,N_37798);
nand U38182 (N_38182,N_37319,N_37190);
and U38183 (N_38183,N_37246,N_37516);
and U38184 (N_38184,N_37766,N_37676);
and U38185 (N_38185,N_37288,N_37905);
or U38186 (N_38186,N_37382,N_37700);
nor U38187 (N_38187,N_37608,N_37466);
nand U38188 (N_38188,N_37488,N_37159);
nor U38189 (N_38189,N_37005,N_37206);
and U38190 (N_38190,N_37040,N_37262);
nor U38191 (N_38191,N_37256,N_37344);
xnor U38192 (N_38192,N_37525,N_37212);
or U38193 (N_38193,N_37586,N_37172);
nand U38194 (N_38194,N_37862,N_37606);
xor U38195 (N_38195,N_37025,N_37610);
xor U38196 (N_38196,N_37099,N_37852);
xnor U38197 (N_38197,N_37077,N_37100);
xnor U38198 (N_38198,N_37323,N_37953);
nand U38199 (N_38199,N_37198,N_37266);
and U38200 (N_38200,N_37118,N_37547);
nand U38201 (N_38201,N_37954,N_37504);
and U38202 (N_38202,N_37430,N_37464);
xnor U38203 (N_38203,N_37331,N_37316);
nor U38204 (N_38204,N_37531,N_37450);
nand U38205 (N_38205,N_37215,N_37690);
nor U38206 (N_38206,N_37449,N_37918);
nand U38207 (N_38207,N_37921,N_37134);
or U38208 (N_38208,N_37543,N_37247);
nor U38209 (N_38209,N_37554,N_37341);
nand U38210 (N_38210,N_37974,N_37259);
xor U38211 (N_38211,N_37012,N_37320);
or U38212 (N_38212,N_37660,N_37477);
nand U38213 (N_38213,N_37754,N_37232);
nor U38214 (N_38214,N_37425,N_37145);
nand U38215 (N_38215,N_37571,N_37496);
xnor U38216 (N_38216,N_37315,N_37555);
and U38217 (N_38217,N_37748,N_37468);
or U38218 (N_38218,N_37545,N_37994);
nand U38219 (N_38219,N_37448,N_37673);
nor U38220 (N_38220,N_37838,N_37272);
nand U38221 (N_38221,N_37926,N_37946);
xnor U38222 (N_38222,N_37979,N_37976);
and U38223 (N_38223,N_37802,N_37281);
nand U38224 (N_38224,N_37796,N_37689);
xor U38225 (N_38225,N_37463,N_37238);
and U38226 (N_38226,N_37598,N_37665);
nor U38227 (N_38227,N_37478,N_37074);
or U38228 (N_38228,N_37599,N_37685);
or U38229 (N_38229,N_37069,N_37600);
xor U38230 (N_38230,N_37763,N_37779);
xor U38231 (N_38231,N_37594,N_37396);
xor U38232 (N_38232,N_37932,N_37062);
nor U38233 (N_38233,N_37724,N_37617);
nor U38234 (N_38234,N_37858,N_37537);
xnor U38235 (N_38235,N_37373,N_37095);
xnor U38236 (N_38236,N_37943,N_37123);
nor U38237 (N_38237,N_37250,N_37472);
and U38238 (N_38238,N_37182,N_37637);
nand U38239 (N_38239,N_37174,N_37106);
nor U38240 (N_38240,N_37378,N_37861);
xnor U38241 (N_38241,N_37414,N_37947);
nand U38242 (N_38242,N_37753,N_37436);
nor U38243 (N_38243,N_37955,N_37625);
or U38244 (N_38244,N_37445,N_37022);
xor U38245 (N_38245,N_37797,N_37393);
xnor U38246 (N_38246,N_37565,N_37148);
nand U38247 (N_38247,N_37903,N_37544);
and U38248 (N_38248,N_37624,N_37226);
nand U38249 (N_38249,N_37248,N_37334);
and U38250 (N_38250,N_37931,N_37067);
or U38251 (N_38251,N_37593,N_37030);
nor U38252 (N_38252,N_37052,N_37356);
nand U38253 (N_38253,N_37655,N_37302);
and U38254 (N_38254,N_37310,N_37539);
and U38255 (N_38255,N_37082,N_37483);
or U38256 (N_38256,N_37540,N_37714);
nand U38257 (N_38257,N_37651,N_37705);
nor U38258 (N_38258,N_37819,N_37171);
or U38259 (N_38259,N_37767,N_37263);
xnor U38260 (N_38260,N_37702,N_37217);
xor U38261 (N_38261,N_37183,N_37242);
or U38262 (N_38262,N_37131,N_37203);
or U38263 (N_38263,N_37267,N_37039);
nand U38264 (N_38264,N_37958,N_37399);
or U38265 (N_38265,N_37210,N_37001);
or U38266 (N_38266,N_37703,N_37290);
nand U38267 (N_38267,N_37401,N_37807);
and U38268 (N_38268,N_37750,N_37985);
or U38269 (N_38269,N_37443,N_37384);
nand U38270 (N_38270,N_37370,N_37687);
and U38271 (N_38271,N_37980,N_37073);
xor U38272 (N_38272,N_37942,N_37834);
and U38273 (N_38273,N_37941,N_37978);
xor U38274 (N_38274,N_37410,N_37254);
xnor U38275 (N_38275,N_37556,N_37326);
and U38276 (N_38276,N_37160,N_37616);
and U38277 (N_38277,N_37358,N_37078);
nand U38278 (N_38278,N_37869,N_37879);
or U38279 (N_38279,N_37351,N_37365);
nor U38280 (N_38280,N_37211,N_37965);
and U38281 (N_38281,N_37330,N_37828);
and U38282 (N_38282,N_37698,N_37276);
nand U38283 (N_38283,N_37927,N_37042);
and U38284 (N_38284,N_37866,N_37114);
nor U38285 (N_38285,N_37470,N_37827);
and U38286 (N_38286,N_37742,N_37755);
nand U38287 (N_38287,N_37173,N_37751);
and U38288 (N_38288,N_37626,N_37694);
nor U38289 (N_38289,N_37429,N_37882);
or U38290 (N_38290,N_37681,N_37166);
nor U38291 (N_38291,N_37218,N_37092);
and U38292 (N_38292,N_37632,N_37087);
or U38293 (N_38293,N_37939,N_37871);
nor U38294 (N_38294,N_37360,N_37240);
nand U38295 (N_38295,N_37769,N_37514);
xor U38296 (N_38296,N_37405,N_37107);
and U38297 (N_38297,N_37440,N_37615);
xnor U38298 (N_38298,N_37764,N_37397);
nor U38299 (N_38299,N_37034,N_37417);
nand U38300 (N_38300,N_37607,N_37249);
or U38301 (N_38301,N_37595,N_37195);
or U38302 (N_38302,N_37642,N_37236);
xor U38303 (N_38303,N_37043,N_37164);
xor U38304 (N_38304,N_37185,N_37252);
nor U38305 (N_38305,N_37667,N_37904);
nor U38306 (N_38306,N_37298,N_37564);
or U38307 (N_38307,N_37428,N_37890);
nor U38308 (N_38308,N_37777,N_37789);
nand U38309 (N_38309,N_37412,N_37691);
nor U38310 (N_38310,N_37066,N_37048);
and U38311 (N_38311,N_37845,N_37297);
and U38312 (N_38312,N_37452,N_37522);
and U38313 (N_38313,N_37906,N_37227);
and U38314 (N_38314,N_37421,N_37562);
xor U38315 (N_38315,N_37723,N_37258);
and U38316 (N_38316,N_37950,N_37678);
xor U38317 (N_38317,N_37041,N_37569);
nor U38318 (N_38318,N_37108,N_37011);
nand U38319 (N_38319,N_37550,N_37390);
or U38320 (N_38320,N_37971,N_37010);
and U38321 (N_38321,N_37152,N_37692);
and U38322 (N_38322,N_37639,N_37585);
nor U38323 (N_38323,N_37032,N_37975);
and U38324 (N_38324,N_37243,N_37580);
and U38325 (N_38325,N_37150,N_37336);
or U38326 (N_38326,N_37325,N_37733);
nand U38327 (N_38327,N_37824,N_37169);
nor U38328 (N_38328,N_37670,N_37140);
or U38329 (N_38329,N_37235,N_37970);
and U38330 (N_38330,N_37158,N_37731);
or U38331 (N_38331,N_37758,N_37841);
or U38332 (N_38332,N_37886,N_37047);
and U38333 (N_38333,N_37574,N_37402);
and U38334 (N_38334,N_37907,N_37346);
nand U38335 (N_38335,N_37936,N_37354);
or U38336 (N_38336,N_37155,N_37794);
and U38337 (N_38337,N_37973,N_37407);
nand U38338 (N_38338,N_37653,N_37801);
or U38339 (N_38339,N_37725,N_37006);
or U38340 (N_38340,N_37538,N_37584);
or U38341 (N_38341,N_37800,N_37342);
nor U38342 (N_38342,N_37981,N_37097);
and U38343 (N_38343,N_37739,N_37813);
or U38344 (N_38344,N_37963,N_37418);
and U38345 (N_38345,N_37622,N_37089);
and U38346 (N_38346,N_37892,N_37749);
or U38347 (N_38347,N_37765,N_37130);
nor U38348 (N_38348,N_37620,N_37920);
or U38349 (N_38349,N_37363,N_37192);
and U38350 (N_38350,N_37094,N_37768);
xor U38351 (N_38351,N_37735,N_37519);
nor U38352 (N_38352,N_37572,N_37260);
nor U38353 (N_38353,N_37783,N_37806);
and U38354 (N_38354,N_37706,N_37781);
xnor U38355 (N_38355,N_37722,N_37388);
nand U38356 (N_38356,N_37876,N_37908);
and U38357 (N_38357,N_37314,N_37561);
and U38358 (N_38358,N_37534,N_37117);
and U38359 (N_38359,N_37083,N_37934);
nand U38360 (N_38360,N_37233,N_37881);
xor U38361 (N_38361,N_37863,N_37849);
or U38362 (N_38362,N_37447,N_37355);
nor U38363 (N_38363,N_37303,N_37671);
nor U38364 (N_38364,N_37296,N_37264);
nand U38365 (N_38365,N_37139,N_37566);
or U38366 (N_38366,N_37567,N_37253);
nor U38367 (N_38367,N_37427,N_37208);
nor U38368 (N_38368,N_37462,N_37013);
and U38369 (N_38369,N_37279,N_37840);
or U38370 (N_38370,N_37793,N_37835);
and U38371 (N_38371,N_37308,N_37785);
xnor U38372 (N_38372,N_37935,N_37136);
or U38373 (N_38373,N_37075,N_37329);
xnor U38374 (N_38374,N_37144,N_37376);
xor U38375 (N_38375,N_37261,N_37575);
and U38376 (N_38376,N_37275,N_37787);
nand U38377 (N_38377,N_37187,N_37916);
and U38378 (N_38378,N_37055,N_37071);
and U38379 (N_38379,N_37872,N_37507);
and U38380 (N_38380,N_37579,N_37684);
or U38381 (N_38381,N_37374,N_37814);
nand U38382 (N_38382,N_37498,N_37656);
nor U38383 (N_38383,N_37163,N_37509);
nand U38384 (N_38384,N_37207,N_37729);
xnor U38385 (N_38385,N_37843,N_37791);
or U38386 (N_38386,N_37124,N_37143);
nor U38387 (N_38387,N_37563,N_37895);
nor U38388 (N_38388,N_37064,N_37122);
or U38389 (N_38389,N_37884,N_37289);
nor U38390 (N_38390,N_37663,N_37475);
nor U38391 (N_38391,N_37434,N_37549);
nor U38392 (N_38392,N_37517,N_37300);
and U38393 (N_38393,N_37949,N_37033);
nor U38394 (N_38394,N_37830,N_37719);
or U38395 (N_38395,N_37188,N_37728);
xnor U38396 (N_38396,N_37200,N_37523);
and U38397 (N_38397,N_37454,N_37194);
or U38398 (N_38398,N_37128,N_37680);
xor U38399 (N_38399,N_37126,N_37658);
or U38400 (N_38400,N_37590,N_37560);
nand U38401 (N_38401,N_37102,N_37345);
or U38402 (N_38402,N_37337,N_37026);
nor U38403 (N_38403,N_37552,N_37499);
nand U38404 (N_38404,N_37268,N_37734);
and U38405 (N_38405,N_37874,N_37003);
nor U38406 (N_38406,N_37640,N_37270);
and U38407 (N_38407,N_37741,N_37592);
or U38408 (N_38408,N_37511,N_37135);
nor U38409 (N_38409,N_37357,N_37770);
nor U38410 (N_38410,N_37424,N_37771);
nor U38411 (N_38411,N_37643,N_37476);
nand U38412 (N_38412,N_37105,N_37647);
or U38413 (N_38413,N_37744,N_37202);
or U38414 (N_38414,N_37487,N_37111);
nor U38415 (N_38415,N_37482,N_37573);
nand U38416 (N_38416,N_37277,N_37220);
xnor U38417 (N_38417,N_37049,N_37878);
nand U38418 (N_38418,N_37184,N_37533);
or U38419 (N_38419,N_37132,N_37672);
or U38420 (N_38420,N_37129,N_37836);
nor U38421 (N_38421,N_37618,N_37752);
or U38422 (N_38422,N_37120,N_37161);
nand U38423 (N_38423,N_37633,N_37666);
nor U38424 (N_38424,N_37746,N_37386);
and U38425 (N_38425,N_37993,N_37177);
or U38426 (N_38426,N_37383,N_37426);
and U38427 (N_38427,N_37654,N_37125);
or U38428 (N_38428,N_37501,N_37406);
nor U38429 (N_38429,N_37541,N_37007);
or U38430 (N_38430,N_37221,N_37962);
nor U38431 (N_38431,N_37146,N_37859);
nand U38432 (N_38432,N_37309,N_37536);
nand U38433 (N_38433,N_37747,N_37455);
and U38434 (N_38434,N_37255,N_37021);
nor U38435 (N_38435,N_37222,N_37322);
and U38436 (N_38436,N_37513,N_37897);
or U38437 (N_38437,N_37018,N_37605);
nor U38438 (N_38438,N_37020,N_37057);
nand U38439 (N_38439,N_37989,N_37991);
nor U38440 (N_38440,N_37645,N_37324);
and U38441 (N_38441,N_37717,N_37662);
xnor U38442 (N_38442,N_37716,N_37969);
and U38443 (N_38443,N_37524,N_37115);
and U38444 (N_38444,N_37437,N_37199);
xnor U38445 (N_38445,N_37558,N_37868);
nand U38446 (N_38446,N_37138,N_37465);
nand U38447 (N_38447,N_37682,N_37967);
or U38448 (N_38448,N_37237,N_37635);
nand U38449 (N_38449,N_37652,N_37856);
xor U38450 (N_38450,N_37494,N_37375);
xor U38451 (N_38451,N_37154,N_37225);
nor U38452 (N_38452,N_37631,N_37340);
nor U38453 (N_38453,N_37110,N_37630);
nand U38454 (N_38454,N_37157,N_37119);
nand U38455 (N_38455,N_37693,N_37175);
xor U38456 (N_38456,N_37023,N_37623);
and U38457 (N_38457,N_37485,N_37818);
and U38458 (N_38458,N_37251,N_37977);
xor U38459 (N_38459,N_37413,N_37223);
xnor U38460 (N_38460,N_37133,N_37193);
and U38461 (N_38461,N_37857,N_37959);
and U38462 (N_38462,N_37675,N_37853);
or U38463 (N_38463,N_37743,N_37812);
or U38464 (N_38464,N_37553,N_37036);
and U38465 (N_38465,N_37016,N_37101);
and U38466 (N_38466,N_37945,N_37548);
nor U38467 (N_38467,N_37930,N_37104);
xnor U38468 (N_38468,N_37738,N_37713);
or U38469 (N_38469,N_37774,N_37708);
nor U38470 (N_38470,N_37557,N_37051);
nand U38471 (N_38471,N_37149,N_37299);
and U38472 (N_38472,N_37659,N_37113);
nand U38473 (N_38473,N_37832,N_37756);
nor U38474 (N_38474,N_37759,N_37737);
or U38475 (N_38475,N_37328,N_37103);
and U38476 (N_38476,N_37720,N_37420);
and U38477 (N_38477,N_37229,N_37792);
or U38478 (N_38478,N_37873,N_37167);
nand U38479 (N_38479,N_37919,N_37015);
or U38480 (N_38480,N_37998,N_37925);
or U38481 (N_38481,N_37677,N_37480);
nor U38482 (N_38482,N_37589,N_37805);
nor U38483 (N_38483,N_37891,N_37031);
xnor U38484 (N_38484,N_37695,N_37587);
xor U38485 (N_38485,N_37784,N_37996);
nand U38486 (N_38486,N_37503,N_37153);
nand U38487 (N_38487,N_37387,N_37960);
nand U38488 (N_38488,N_37431,N_37294);
and U38489 (N_38489,N_37231,N_37446);
and U38490 (N_38490,N_37109,N_37467);
nand U38491 (N_38491,N_37273,N_37295);
nand U38492 (N_38492,N_37898,N_37528);
and U38493 (N_38493,N_37380,N_37165);
xor U38494 (N_38494,N_37761,N_37990);
xor U38495 (N_38495,N_37641,N_37997);
and U38496 (N_38496,N_37816,N_37081);
nor U38497 (N_38497,N_37301,N_37581);
and U38498 (N_38498,N_37899,N_37234);
or U38499 (N_38499,N_37987,N_37854);
xnor U38500 (N_38500,N_37706,N_37074);
nand U38501 (N_38501,N_37210,N_37878);
nand U38502 (N_38502,N_37148,N_37142);
or U38503 (N_38503,N_37945,N_37035);
nor U38504 (N_38504,N_37607,N_37401);
xor U38505 (N_38505,N_37300,N_37898);
and U38506 (N_38506,N_37953,N_37128);
nand U38507 (N_38507,N_37954,N_37919);
or U38508 (N_38508,N_37438,N_37759);
nand U38509 (N_38509,N_37479,N_37405);
xor U38510 (N_38510,N_37510,N_37194);
nor U38511 (N_38511,N_37188,N_37797);
nor U38512 (N_38512,N_37881,N_37137);
nand U38513 (N_38513,N_37654,N_37353);
nand U38514 (N_38514,N_37053,N_37755);
or U38515 (N_38515,N_37781,N_37597);
xor U38516 (N_38516,N_37404,N_37368);
and U38517 (N_38517,N_37569,N_37795);
or U38518 (N_38518,N_37287,N_37957);
xor U38519 (N_38519,N_37388,N_37641);
or U38520 (N_38520,N_37377,N_37774);
nor U38521 (N_38521,N_37546,N_37510);
xor U38522 (N_38522,N_37329,N_37146);
nand U38523 (N_38523,N_37381,N_37266);
nand U38524 (N_38524,N_37693,N_37302);
xnor U38525 (N_38525,N_37934,N_37889);
and U38526 (N_38526,N_37324,N_37635);
nor U38527 (N_38527,N_37904,N_37997);
nand U38528 (N_38528,N_37345,N_37569);
nor U38529 (N_38529,N_37194,N_37434);
nand U38530 (N_38530,N_37790,N_37999);
xnor U38531 (N_38531,N_37160,N_37785);
nand U38532 (N_38532,N_37920,N_37185);
and U38533 (N_38533,N_37350,N_37258);
and U38534 (N_38534,N_37268,N_37026);
nand U38535 (N_38535,N_37881,N_37749);
or U38536 (N_38536,N_37221,N_37010);
and U38537 (N_38537,N_37976,N_37301);
or U38538 (N_38538,N_37580,N_37107);
nand U38539 (N_38539,N_37697,N_37652);
or U38540 (N_38540,N_37004,N_37688);
or U38541 (N_38541,N_37261,N_37849);
nand U38542 (N_38542,N_37737,N_37467);
or U38543 (N_38543,N_37123,N_37207);
or U38544 (N_38544,N_37405,N_37789);
nand U38545 (N_38545,N_37090,N_37568);
xnor U38546 (N_38546,N_37444,N_37094);
and U38547 (N_38547,N_37680,N_37817);
nand U38548 (N_38548,N_37907,N_37371);
and U38549 (N_38549,N_37144,N_37256);
xnor U38550 (N_38550,N_37799,N_37349);
and U38551 (N_38551,N_37542,N_37897);
and U38552 (N_38552,N_37016,N_37139);
and U38553 (N_38553,N_37586,N_37502);
nand U38554 (N_38554,N_37118,N_37688);
or U38555 (N_38555,N_37010,N_37257);
nor U38556 (N_38556,N_37103,N_37016);
or U38557 (N_38557,N_37893,N_37292);
xor U38558 (N_38558,N_37907,N_37506);
xnor U38559 (N_38559,N_37677,N_37508);
or U38560 (N_38560,N_37828,N_37225);
nand U38561 (N_38561,N_37513,N_37765);
xor U38562 (N_38562,N_37863,N_37967);
and U38563 (N_38563,N_37030,N_37148);
nand U38564 (N_38564,N_37060,N_37789);
nor U38565 (N_38565,N_37105,N_37914);
nand U38566 (N_38566,N_37072,N_37344);
nand U38567 (N_38567,N_37236,N_37159);
or U38568 (N_38568,N_37209,N_37119);
xor U38569 (N_38569,N_37431,N_37382);
and U38570 (N_38570,N_37255,N_37169);
nand U38571 (N_38571,N_37576,N_37364);
nand U38572 (N_38572,N_37863,N_37327);
nand U38573 (N_38573,N_37692,N_37552);
nor U38574 (N_38574,N_37985,N_37209);
xor U38575 (N_38575,N_37636,N_37110);
nor U38576 (N_38576,N_37075,N_37502);
and U38577 (N_38577,N_37063,N_37598);
and U38578 (N_38578,N_37272,N_37476);
nand U38579 (N_38579,N_37915,N_37791);
nand U38580 (N_38580,N_37805,N_37330);
nor U38581 (N_38581,N_37935,N_37024);
nor U38582 (N_38582,N_37246,N_37554);
nor U38583 (N_38583,N_37462,N_37988);
nor U38584 (N_38584,N_37760,N_37592);
nand U38585 (N_38585,N_37495,N_37009);
and U38586 (N_38586,N_37543,N_37430);
or U38587 (N_38587,N_37377,N_37783);
xnor U38588 (N_38588,N_37738,N_37628);
xnor U38589 (N_38589,N_37238,N_37219);
nor U38590 (N_38590,N_37380,N_37800);
nand U38591 (N_38591,N_37990,N_37656);
or U38592 (N_38592,N_37022,N_37060);
nor U38593 (N_38593,N_37028,N_37707);
nand U38594 (N_38594,N_37664,N_37765);
and U38595 (N_38595,N_37726,N_37962);
nand U38596 (N_38596,N_37236,N_37639);
nand U38597 (N_38597,N_37605,N_37484);
nand U38598 (N_38598,N_37893,N_37302);
and U38599 (N_38599,N_37364,N_37098);
xnor U38600 (N_38600,N_37962,N_37887);
and U38601 (N_38601,N_37826,N_37656);
or U38602 (N_38602,N_37736,N_37356);
and U38603 (N_38603,N_37446,N_37547);
nor U38604 (N_38604,N_37327,N_37105);
nor U38605 (N_38605,N_37594,N_37853);
and U38606 (N_38606,N_37584,N_37670);
nand U38607 (N_38607,N_37071,N_37529);
nor U38608 (N_38608,N_37236,N_37919);
nand U38609 (N_38609,N_37751,N_37197);
xnor U38610 (N_38610,N_37085,N_37182);
nand U38611 (N_38611,N_37830,N_37098);
xor U38612 (N_38612,N_37025,N_37399);
and U38613 (N_38613,N_37610,N_37498);
nand U38614 (N_38614,N_37459,N_37791);
xor U38615 (N_38615,N_37322,N_37538);
nor U38616 (N_38616,N_37865,N_37249);
nor U38617 (N_38617,N_37066,N_37063);
xnor U38618 (N_38618,N_37503,N_37710);
nor U38619 (N_38619,N_37448,N_37714);
nor U38620 (N_38620,N_37361,N_37190);
nand U38621 (N_38621,N_37865,N_37220);
nand U38622 (N_38622,N_37332,N_37641);
nor U38623 (N_38623,N_37901,N_37595);
or U38624 (N_38624,N_37447,N_37677);
or U38625 (N_38625,N_37512,N_37496);
xor U38626 (N_38626,N_37539,N_37427);
and U38627 (N_38627,N_37828,N_37069);
xnor U38628 (N_38628,N_37070,N_37162);
or U38629 (N_38629,N_37994,N_37686);
nor U38630 (N_38630,N_37442,N_37188);
or U38631 (N_38631,N_37842,N_37928);
and U38632 (N_38632,N_37290,N_37908);
or U38633 (N_38633,N_37380,N_37683);
or U38634 (N_38634,N_37651,N_37997);
nor U38635 (N_38635,N_37906,N_37549);
or U38636 (N_38636,N_37807,N_37682);
or U38637 (N_38637,N_37889,N_37108);
and U38638 (N_38638,N_37752,N_37542);
xnor U38639 (N_38639,N_37448,N_37813);
or U38640 (N_38640,N_37236,N_37990);
or U38641 (N_38641,N_37502,N_37836);
nor U38642 (N_38642,N_37532,N_37184);
xnor U38643 (N_38643,N_37212,N_37921);
nor U38644 (N_38644,N_37026,N_37136);
xor U38645 (N_38645,N_37299,N_37296);
nand U38646 (N_38646,N_37538,N_37806);
nor U38647 (N_38647,N_37193,N_37739);
and U38648 (N_38648,N_37858,N_37058);
and U38649 (N_38649,N_37862,N_37214);
or U38650 (N_38650,N_37793,N_37932);
xnor U38651 (N_38651,N_37476,N_37894);
xnor U38652 (N_38652,N_37138,N_37359);
nand U38653 (N_38653,N_37793,N_37032);
and U38654 (N_38654,N_37242,N_37626);
and U38655 (N_38655,N_37604,N_37148);
and U38656 (N_38656,N_37369,N_37810);
and U38657 (N_38657,N_37529,N_37930);
or U38658 (N_38658,N_37889,N_37426);
xnor U38659 (N_38659,N_37727,N_37476);
nor U38660 (N_38660,N_37074,N_37841);
nand U38661 (N_38661,N_37127,N_37392);
or U38662 (N_38662,N_37105,N_37790);
nand U38663 (N_38663,N_37110,N_37694);
nor U38664 (N_38664,N_37040,N_37320);
nand U38665 (N_38665,N_37300,N_37294);
nor U38666 (N_38666,N_37818,N_37177);
xor U38667 (N_38667,N_37504,N_37669);
xor U38668 (N_38668,N_37330,N_37274);
nor U38669 (N_38669,N_37321,N_37080);
nor U38670 (N_38670,N_37834,N_37746);
nand U38671 (N_38671,N_37484,N_37458);
nand U38672 (N_38672,N_37786,N_37615);
nor U38673 (N_38673,N_37341,N_37932);
nand U38674 (N_38674,N_37279,N_37734);
and U38675 (N_38675,N_37841,N_37256);
nand U38676 (N_38676,N_37040,N_37275);
or U38677 (N_38677,N_37879,N_37953);
and U38678 (N_38678,N_37236,N_37111);
xnor U38679 (N_38679,N_37918,N_37309);
and U38680 (N_38680,N_37947,N_37967);
or U38681 (N_38681,N_37742,N_37230);
and U38682 (N_38682,N_37095,N_37072);
nor U38683 (N_38683,N_37379,N_37602);
or U38684 (N_38684,N_37161,N_37925);
or U38685 (N_38685,N_37489,N_37048);
or U38686 (N_38686,N_37925,N_37221);
xor U38687 (N_38687,N_37771,N_37625);
and U38688 (N_38688,N_37903,N_37401);
and U38689 (N_38689,N_37479,N_37549);
nor U38690 (N_38690,N_37564,N_37667);
or U38691 (N_38691,N_37706,N_37496);
and U38692 (N_38692,N_37052,N_37677);
nor U38693 (N_38693,N_37867,N_37173);
and U38694 (N_38694,N_37174,N_37314);
nand U38695 (N_38695,N_37467,N_37497);
nand U38696 (N_38696,N_37034,N_37057);
nor U38697 (N_38697,N_37872,N_37647);
xor U38698 (N_38698,N_37659,N_37292);
nand U38699 (N_38699,N_37089,N_37674);
or U38700 (N_38700,N_37929,N_37500);
and U38701 (N_38701,N_37996,N_37646);
xnor U38702 (N_38702,N_37920,N_37881);
xnor U38703 (N_38703,N_37654,N_37227);
and U38704 (N_38704,N_37995,N_37016);
nand U38705 (N_38705,N_37019,N_37473);
and U38706 (N_38706,N_37604,N_37249);
xor U38707 (N_38707,N_37837,N_37831);
nand U38708 (N_38708,N_37991,N_37774);
and U38709 (N_38709,N_37536,N_37690);
nand U38710 (N_38710,N_37544,N_37177);
and U38711 (N_38711,N_37052,N_37644);
or U38712 (N_38712,N_37223,N_37593);
or U38713 (N_38713,N_37800,N_37866);
or U38714 (N_38714,N_37589,N_37712);
or U38715 (N_38715,N_37717,N_37851);
nand U38716 (N_38716,N_37955,N_37602);
nand U38717 (N_38717,N_37361,N_37736);
xnor U38718 (N_38718,N_37033,N_37689);
nand U38719 (N_38719,N_37410,N_37073);
nor U38720 (N_38720,N_37787,N_37585);
nand U38721 (N_38721,N_37203,N_37885);
nor U38722 (N_38722,N_37059,N_37912);
xor U38723 (N_38723,N_37892,N_37504);
nand U38724 (N_38724,N_37787,N_37587);
or U38725 (N_38725,N_37094,N_37704);
and U38726 (N_38726,N_37112,N_37930);
nor U38727 (N_38727,N_37814,N_37318);
xnor U38728 (N_38728,N_37750,N_37565);
xnor U38729 (N_38729,N_37597,N_37679);
xnor U38730 (N_38730,N_37433,N_37858);
xnor U38731 (N_38731,N_37941,N_37803);
nand U38732 (N_38732,N_37671,N_37237);
or U38733 (N_38733,N_37947,N_37127);
nand U38734 (N_38734,N_37292,N_37008);
nand U38735 (N_38735,N_37526,N_37381);
xor U38736 (N_38736,N_37988,N_37067);
xor U38737 (N_38737,N_37670,N_37883);
or U38738 (N_38738,N_37225,N_37772);
or U38739 (N_38739,N_37421,N_37271);
xor U38740 (N_38740,N_37931,N_37952);
or U38741 (N_38741,N_37301,N_37184);
nor U38742 (N_38742,N_37424,N_37950);
nor U38743 (N_38743,N_37808,N_37777);
xnor U38744 (N_38744,N_37445,N_37141);
nand U38745 (N_38745,N_37508,N_37305);
or U38746 (N_38746,N_37200,N_37896);
nor U38747 (N_38747,N_37665,N_37650);
nor U38748 (N_38748,N_37396,N_37452);
and U38749 (N_38749,N_37820,N_37927);
and U38750 (N_38750,N_37717,N_37867);
nor U38751 (N_38751,N_37898,N_37131);
or U38752 (N_38752,N_37129,N_37343);
or U38753 (N_38753,N_37524,N_37739);
nor U38754 (N_38754,N_37106,N_37108);
nand U38755 (N_38755,N_37278,N_37047);
nand U38756 (N_38756,N_37674,N_37728);
xnor U38757 (N_38757,N_37963,N_37360);
nor U38758 (N_38758,N_37198,N_37850);
or U38759 (N_38759,N_37686,N_37821);
nor U38760 (N_38760,N_37117,N_37829);
nand U38761 (N_38761,N_37253,N_37708);
and U38762 (N_38762,N_37376,N_37288);
and U38763 (N_38763,N_37701,N_37467);
nand U38764 (N_38764,N_37893,N_37045);
or U38765 (N_38765,N_37838,N_37429);
or U38766 (N_38766,N_37338,N_37170);
xor U38767 (N_38767,N_37663,N_37960);
nor U38768 (N_38768,N_37992,N_37335);
or U38769 (N_38769,N_37426,N_37202);
and U38770 (N_38770,N_37413,N_37023);
and U38771 (N_38771,N_37370,N_37856);
xor U38772 (N_38772,N_37466,N_37246);
nand U38773 (N_38773,N_37154,N_37893);
nand U38774 (N_38774,N_37429,N_37534);
or U38775 (N_38775,N_37395,N_37877);
nand U38776 (N_38776,N_37801,N_37641);
or U38777 (N_38777,N_37721,N_37616);
nor U38778 (N_38778,N_37364,N_37077);
nand U38779 (N_38779,N_37999,N_37586);
or U38780 (N_38780,N_37114,N_37298);
nor U38781 (N_38781,N_37123,N_37600);
or U38782 (N_38782,N_37560,N_37337);
nand U38783 (N_38783,N_37537,N_37514);
and U38784 (N_38784,N_37672,N_37946);
nand U38785 (N_38785,N_37894,N_37157);
xor U38786 (N_38786,N_37251,N_37381);
and U38787 (N_38787,N_37853,N_37802);
xor U38788 (N_38788,N_37867,N_37533);
nor U38789 (N_38789,N_37610,N_37018);
nand U38790 (N_38790,N_37788,N_37914);
and U38791 (N_38791,N_37849,N_37985);
or U38792 (N_38792,N_37266,N_37150);
and U38793 (N_38793,N_37274,N_37471);
nor U38794 (N_38794,N_37405,N_37603);
nand U38795 (N_38795,N_37399,N_37349);
nand U38796 (N_38796,N_37003,N_37154);
nor U38797 (N_38797,N_37551,N_37752);
or U38798 (N_38798,N_37876,N_37194);
and U38799 (N_38799,N_37614,N_37582);
xor U38800 (N_38800,N_37304,N_37280);
and U38801 (N_38801,N_37842,N_37758);
nand U38802 (N_38802,N_37180,N_37917);
nand U38803 (N_38803,N_37481,N_37630);
or U38804 (N_38804,N_37121,N_37833);
nand U38805 (N_38805,N_37275,N_37305);
and U38806 (N_38806,N_37695,N_37035);
and U38807 (N_38807,N_37047,N_37810);
nor U38808 (N_38808,N_37733,N_37708);
xnor U38809 (N_38809,N_37233,N_37392);
and U38810 (N_38810,N_37973,N_37639);
or U38811 (N_38811,N_37664,N_37187);
nand U38812 (N_38812,N_37634,N_37352);
or U38813 (N_38813,N_37680,N_37470);
and U38814 (N_38814,N_37684,N_37692);
xor U38815 (N_38815,N_37347,N_37764);
and U38816 (N_38816,N_37761,N_37508);
nor U38817 (N_38817,N_37669,N_37045);
or U38818 (N_38818,N_37518,N_37574);
or U38819 (N_38819,N_37399,N_37553);
nand U38820 (N_38820,N_37818,N_37010);
nand U38821 (N_38821,N_37384,N_37456);
and U38822 (N_38822,N_37142,N_37812);
nor U38823 (N_38823,N_37079,N_37270);
xnor U38824 (N_38824,N_37879,N_37313);
nor U38825 (N_38825,N_37888,N_37270);
xnor U38826 (N_38826,N_37591,N_37790);
and U38827 (N_38827,N_37028,N_37131);
nor U38828 (N_38828,N_37027,N_37412);
nand U38829 (N_38829,N_37566,N_37900);
nor U38830 (N_38830,N_37823,N_37026);
nand U38831 (N_38831,N_37884,N_37798);
nor U38832 (N_38832,N_37320,N_37275);
or U38833 (N_38833,N_37446,N_37329);
or U38834 (N_38834,N_37301,N_37846);
or U38835 (N_38835,N_37012,N_37928);
nor U38836 (N_38836,N_37138,N_37846);
and U38837 (N_38837,N_37713,N_37044);
nand U38838 (N_38838,N_37017,N_37020);
nand U38839 (N_38839,N_37172,N_37785);
nor U38840 (N_38840,N_37626,N_37552);
or U38841 (N_38841,N_37053,N_37603);
nor U38842 (N_38842,N_37496,N_37379);
nor U38843 (N_38843,N_37280,N_37153);
and U38844 (N_38844,N_37784,N_37579);
nor U38845 (N_38845,N_37773,N_37315);
nor U38846 (N_38846,N_37437,N_37763);
or U38847 (N_38847,N_37747,N_37893);
nand U38848 (N_38848,N_37161,N_37223);
and U38849 (N_38849,N_37766,N_37506);
nor U38850 (N_38850,N_37069,N_37354);
and U38851 (N_38851,N_37601,N_37023);
nor U38852 (N_38852,N_37066,N_37455);
or U38853 (N_38853,N_37259,N_37629);
or U38854 (N_38854,N_37761,N_37449);
or U38855 (N_38855,N_37923,N_37875);
xnor U38856 (N_38856,N_37051,N_37063);
and U38857 (N_38857,N_37851,N_37544);
or U38858 (N_38858,N_37387,N_37274);
nand U38859 (N_38859,N_37050,N_37661);
xnor U38860 (N_38860,N_37564,N_37387);
and U38861 (N_38861,N_37768,N_37873);
nand U38862 (N_38862,N_37758,N_37190);
nor U38863 (N_38863,N_37378,N_37503);
and U38864 (N_38864,N_37982,N_37967);
xnor U38865 (N_38865,N_37537,N_37558);
or U38866 (N_38866,N_37771,N_37195);
nand U38867 (N_38867,N_37165,N_37966);
nor U38868 (N_38868,N_37944,N_37238);
or U38869 (N_38869,N_37467,N_37566);
nor U38870 (N_38870,N_37459,N_37958);
and U38871 (N_38871,N_37587,N_37247);
nand U38872 (N_38872,N_37691,N_37817);
nor U38873 (N_38873,N_37090,N_37614);
xnor U38874 (N_38874,N_37312,N_37907);
and U38875 (N_38875,N_37619,N_37342);
nand U38876 (N_38876,N_37377,N_37678);
or U38877 (N_38877,N_37604,N_37941);
nor U38878 (N_38878,N_37256,N_37738);
and U38879 (N_38879,N_37885,N_37445);
or U38880 (N_38880,N_37702,N_37252);
and U38881 (N_38881,N_37482,N_37470);
or U38882 (N_38882,N_37898,N_37262);
nand U38883 (N_38883,N_37816,N_37566);
nor U38884 (N_38884,N_37961,N_37337);
and U38885 (N_38885,N_37164,N_37195);
nand U38886 (N_38886,N_37007,N_37199);
or U38887 (N_38887,N_37759,N_37726);
and U38888 (N_38888,N_37029,N_37482);
and U38889 (N_38889,N_37421,N_37307);
xor U38890 (N_38890,N_37585,N_37592);
nand U38891 (N_38891,N_37926,N_37347);
xnor U38892 (N_38892,N_37728,N_37649);
and U38893 (N_38893,N_37270,N_37016);
xor U38894 (N_38894,N_37093,N_37057);
and U38895 (N_38895,N_37062,N_37789);
xnor U38896 (N_38896,N_37289,N_37965);
xnor U38897 (N_38897,N_37021,N_37065);
or U38898 (N_38898,N_37512,N_37527);
and U38899 (N_38899,N_37160,N_37905);
and U38900 (N_38900,N_37539,N_37749);
or U38901 (N_38901,N_37826,N_37850);
nor U38902 (N_38902,N_37919,N_37397);
or U38903 (N_38903,N_37833,N_37736);
or U38904 (N_38904,N_37441,N_37368);
xnor U38905 (N_38905,N_37855,N_37364);
nand U38906 (N_38906,N_37430,N_37141);
nor U38907 (N_38907,N_37021,N_37151);
xnor U38908 (N_38908,N_37493,N_37309);
xor U38909 (N_38909,N_37716,N_37107);
xor U38910 (N_38910,N_37684,N_37765);
and U38911 (N_38911,N_37946,N_37001);
and U38912 (N_38912,N_37082,N_37663);
nand U38913 (N_38913,N_37523,N_37226);
nand U38914 (N_38914,N_37627,N_37784);
and U38915 (N_38915,N_37498,N_37995);
xor U38916 (N_38916,N_37603,N_37682);
or U38917 (N_38917,N_37123,N_37786);
or U38918 (N_38918,N_37206,N_37014);
nand U38919 (N_38919,N_37734,N_37560);
nor U38920 (N_38920,N_37764,N_37374);
and U38921 (N_38921,N_37945,N_37747);
xnor U38922 (N_38922,N_37636,N_37020);
nand U38923 (N_38923,N_37355,N_37661);
xor U38924 (N_38924,N_37666,N_37220);
nor U38925 (N_38925,N_37560,N_37767);
nand U38926 (N_38926,N_37152,N_37918);
xnor U38927 (N_38927,N_37534,N_37712);
nor U38928 (N_38928,N_37058,N_37264);
xnor U38929 (N_38929,N_37207,N_37182);
or U38930 (N_38930,N_37278,N_37005);
nand U38931 (N_38931,N_37201,N_37969);
and U38932 (N_38932,N_37012,N_37821);
nor U38933 (N_38933,N_37595,N_37729);
nor U38934 (N_38934,N_37553,N_37529);
or U38935 (N_38935,N_37430,N_37537);
or U38936 (N_38936,N_37206,N_37149);
or U38937 (N_38937,N_37648,N_37587);
nand U38938 (N_38938,N_37306,N_37004);
nor U38939 (N_38939,N_37751,N_37404);
xor U38940 (N_38940,N_37179,N_37540);
nor U38941 (N_38941,N_37564,N_37078);
xnor U38942 (N_38942,N_37947,N_37736);
and U38943 (N_38943,N_37975,N_37064);
and U38944 (N_38944,N_37073,N_37493);
xor U38945 (N_38945,N_37724,N_37277);
xor U38946 (N_38946,N_37576,N_37660);
nor U38947 (N_38947,N_37817,N_37953);
xor U38948 (N_38948,N_37847,N_37004);
or U38949 (N_38949,N_37386,N_37404);
xor U38950 (N_38950,N_37686,N_37125);
and U38951 (N_38951,N_37905,N_37814);
nor U38952 (N_38952,N_37742,N_37241);
or U38953 (N_38953,N_37681,N_37646);
nand U38954 (N_38954,N_37612,N_37365);
nand U38955 (N_38955,N_37300,N_37664);
nand U38956 (N_38956,N_37269,N_37864);
nand U38957 (N_38957,N_37326,N_37378);
xnor U38958 (N_38958,N_37695,N_37398);
xnor U38959 (N_38959,N_37190,N_37173);
or U38960 (N_38960,N_37209,N_37022);
nor U38961 (N_38961,N_37134,N_37090);
and U38962 (N_38962,N_37435,N_37269);
xor U38963 (N_38963,N_37416,N_37811);
or U38964 (N_38964,N_37075,N_37316);
or U38965 (N_38965,N_37071,N_37347);
xor U38966 (N_38966,N_37885,N_37812);
nor U38967 (N_38967,N_37934,N_37243);
and U38968 (N_38968,N_37246,N_37567);
nand U38969 (N_38969,N_37598,N_37465);
nand U38970 (N_38970,N_37232,N_37477);
nor U38971 (N_38971,N_37382,N_37587);
xnor U38972 (N_38972,N_37127,N_37940);
nand U38973 (N_38973,N_37947,N_37175);
or U38974 (N_38974,N_37283,N_37079);
xor U38975 (N_38975,N_37370,N_37931);
nand U38976 (N_38976,N_37420,N_37257);
nand U38977 (N_38977,N_37948,N_37495);
and U38978 (N_38978,N_37657,N_37637);
nand U38979 (N_38979,N_37436,N_37083);
nand U38980 (N_38980,N_37728,N_37181);
nor U38981 (N_38981,N_37319,N_37485);
and U38982 (N_38982,N_37754,N_37484);
or U38983 (N_38983,N_37596,N_37833);
and U38984 (N_38984,N_37964,N_37845);
and U38985 (N_38985,N_37940,N_37945);
or U38986 (N_38986,N_37392,N_37419);
and U38987 (N_38987,N_37247,N_37257);
xnor U38988 (N_38988,N_37547,N_37470);
nor U38989 (N_38989,N_37394,N_37558);
and U38990 (N_38990,N_37047,N_37150);
nand U38991 (N_38991,N_37916,N_37256);
nand U38992 (N_38992,N_37878,N_37477);
xor U38993 (N_38993,N_37670,N_37607);
xor U38994 (N_38994,N_37199,N_37027);
and U38995 (N_38995,N_37516,N_37778);
xor U38996 (N_38996,N_37567,N_37664);
or U38997 (N_38997,N_37905,N_37356);
and U38998 (N_38998,N_37423,N_37086);
or U38999 (N_38999,N_37021,N_37236);
nor U39000 (N_39000,N_38407,N_38309);
xnor U39001 (N_39001,N_38960,N_38063);
nor U39002 (N_39002,N_38489,N_38593);
xnor U39003 (N_39003,N_38260,N_38040);
xnor U39004 (N_39004,N_38302,N_38797);
and U39005 (N_39005,N_38706,N_38197);
or U39006 (N_39006,N_38947,N_38699);
xnor U39007 (N_39007,N_38564,N_38130);
nand U39008 (N_39008,N_38323,N_38060);
or U39009 (N_39009,N_38740,N_38567);
nand U39010 (N_39010,N_38349,N_38565);
or U39011 (N_39011,N_38529,N_38111);
and U39012 (N_39012,N_38480,N_38575);
and U39013 (N_39013,N_38850,N_38647);
nand U39014 (N_39014,N_38073,N_38666);
xnor U39015 (N_39015,N_38044,N_38064);
xnor U39016 (N_39016,N_38746,N_38041);
nor U39017 (N_39017,N_38872,N_38570);
and U39018 (N_39018,N_38681,N_38750);
and U39019 (N_39019,N_38475,N_38227);
or U39020 (N_39020,N_38134,N_38618);
xor U39021 (N_39021,N_38853,N_38720);
nand U39022 (N_39022,N_38043,N_38312);
and U39023 (N_39023,N_38836,N_38365);
or U39024 (N_39024,N_38255,N_38616);
nor U39025 (N_39025,N_38627,N_38758);
and U39026 (N_39026,N_38362,N_38074);
xor U39027 (N_39027,N_38672,N_38865);
xor U39028 (N_39028,N_38327,N_38526);
and U39029 (N_39029,N_38752,N_38334);
xnor U39030 (N_39030,N_38430,N_38726);
and U39031 (N_39031,N_38711,N_38289);
nand U39032 (N_39032,N_38221,N_38014);
and U39033 (N_39033,N_38154,N_38093);
and U39034 (N_39034,N_38488,N_38590);
and U39035 (N_39035,N_38251,N_38902);
xnor U39036 (N_39036,N_38248,N_38188);
xnor U39037 (N_39037,N_38846,N_38701);
nor U39038 (N_39038,N_38719,N_38025);
nor U39039 (N_39039,N_38199,N_38031);
nor U39040 (N_39040,N_38801,N_38363);
or U39041 (N_39041,N_38462,N_38767);
xor U39042 (N_39042,N_38001,N_38374);
and U39043 (N_39043,N_38625,N_38694);
or U39044 (N_39044,N_38211,N_38149);
or U39045 (N_39045,N_38538,N_38057);
or U39046 (N_39046,N_38795,N_38447);
nor U39047 (N_39047,N_38626,N_38971);
nor U39048 (N_39048,N_38079,N_38989);
nand U39049 (N_39049,N_38721,N_38898);
and U39050 (N_39050,N_38875,N_38770);
nand U39051 (N_39051,N_38459,N_38937);
nor U39052 (N_39052,N_38174,N_38743);
xnor U39053 (N_39053,N_38406,N_38279);
and U39054 (N_39054,N_38152,N_38737);
and U39055 (N_39055,N_38926,N_38912);
or U39056 (N_39056,N_38804,N_38696);
and U39057 (N_39057,N_38753,N_38051);
or U39058 (N_39058,N_38654,N_38559);
nor U39059 (N_39059,N_38536,N_38092);
nor U39060 (N_39060,N_38889,N_38669);
nor U39061 (N_39061,N_38950,N_38324);
or U39062 (N_39062,N_38004,N_38532);
or U39063 (N_39063,N_38765,N_38725);
xnor U39064 (N_39064,N_38470,N_38858);
nand U39065 (N_39065,N_38042,N_38441);
or U39066 (N_39066,N_38288,N_38422);
and U39067 (N_39067,N_38683,N_38942);
nand U39068 (N_39068,N_38397,N_38688);
and U39069 (N_39069,N_38281,N_38698);
and U39070 (N_39070,N_38817,N_38034);
xor U39071 (N_39071,N_38990,N_38945);
nand U39072 (N_39072,N_38477,N_38261);
xnor U39073 (N_39073,N_38471,N_38563);
or U39074 (N_39074,N_38774,N_38476);
and U39075 (N_39075,N_38209,N_38777);
and U39076 (N_39076,N_38649,N_38491);
or U39077 (N_39077,N_38574,N_38921);
or U39078 (N_39078,N_38998,N_38062);
or U39079 (N_39079,N_38651,N_38375);
xor U39080 (N_39080,N_38038,N_38298);
nand U39081 (N_39081,N_38794,N_38586);
nand U39082 (N_39082,N_38333,N_38613);
nand U39083 (N_39083,N_38037,N_38581);
and U39084 (N_39084,N_38700,N_38854);
and U39085 (N_39085,N_38604,N_38112);
or U39086 (N_39086,N_38506,N_38523);
nand U39087 (N_39087,N_38445,N_38030);
and U39088 (N_39088,N_38633,N_38249);
and U39089 (N_39089,N_38120,N_38515);
nand U39090 (N_39090,N_38301,N_38754);
nor U39091 (N_39091,N_38216,N_38479);
and U39092 (N_39092,N_38167,N_38424);
xnor U39093 (N_39093,N_38553,N_38493);
or U39094 (N_39094,N_38531,N_38356);
or U39095 (N_39095,N_38002,N_38252);
and U39096 (N_39096,N_38687,N_38439);
xor U39097 (N_39097,N_38233,N_38451);
nand U39098 (N_39098,N_38572,N_38440);
nand U39099 (N_39099,N_38602,N_38929);
and U39100 (N_39100,N_38418,N_38376);
xor U39101 (N_39101,N_38524,N_38876);
or U39102 (N_39102,N_38219,N_38163);
and U39103 (N_39103,N_38139,N_38552);
nor U39104 (N_39104,N_38083,N_38528);
nand U39105 (N_39105,N_38562,N_38592);
nand U39106 (N_39106,N_38748,N_38463);
or U39107 (N_39107,N_38355,N_38114);
or U39108 (N_39108,N_38343,N_38319);
nand U39109 (N_39109,N_38186,N_38224);
nand U39110 (N_39110,N_38100,N_38996);
and U39111 (N_39111,N_38107,N_38049);
or U39112 (N_39112,N_38534,N_38554);
or U39113 (N_39113,N_38772,N_38709);
or U39114 (N_39114,N_38591,N_38845);
or U39115 (N_39115,N_38123,N_38839);
and U39116 (N_39116,N_38697,N_38816);
or U39117 (N_39117,N_38793,N_38657);
xnor U39118 (N_39118,N_38980,N_38663);
nand U39119 (N_39119,N_38915,N_38566);
nor U39120 (N_39120,N_38861,N_38165);
xor U39121 (N_39121,N_38315,N_38690);
xor U39122 (N_39122,N_38196,N_38595);
or U39123 (N_39123,N_38612,N_38603);
nand U39124 (N_39124,N_38432,N_38253);
or U39125 (N_39125,N_38851,N_38168);
and U39126 (N_39126,N_38667,N_38398);
nand U39127 (N_39127,N_38478,N_38230);
nand U39128 (N_39128,N_38502,N_38803);
nor U39129 (N_39129,N_38766,N_38949);
or U39130 (N_39130,N_38503,N_38704);
nand U39131 (N_39131,N_38620,N_38443);
nand U39132 (N_39132,N_38905,N_38871);
xnor U39133 (N_39133,N_38778,N_38548);
or U39134 (N_39134,N_38358,N_38710);
xnor U39135 (N_39135,N_38967,N_38756);
xnor U39136 (N_39136,N_38294,N_38383);
and U39137 (N_39137,N_38232,N_38886);
xor U39138 (N_39138,N_38660,N_38017);
and U39139 (N_39139,N_38306,N_38968);
xnor U39140 (N_39140,N_38285,N_38438);
xnor U39141 (N_39141,N_38320,N_38741);
nand U39142 (N_39142,N_38582,N_38150);
nand U39143 (N_39143,N_38576,N_38692);
or U39144 (N_39144,N_38205,N_38070);
nand U39145 (N_39145,N_38594,N_38065);
or U39146 (N_39146,N_38055,N_38304);
nand U39147 (N_39147,N_38852,N_38664);
nor U39148 (N_39148,N_38371,N_38512);
or U39149 (N_39149,N_38317,N_38678);
xor U39150 (N_39150,N_38173,N_38519);
xor U39151 (N_39151,N_38452,N_38608);
xor U39152 (N_39152,N_38705,N_38913);
or U39153 (N_39153,N_38089,N_38550);
xnor U39154 (N_39154,N_38991,N_38466);
nor U39155 (N_39155,N_38088,N_38372);
nand U39156 (N_39156,N_38113,N_38557);
and U39157 (N_39157,N_38464,N_38105);
xnor U39158 (N_39158,N_38855,N_38033);
and U39159 (N_39159,N_38344,N_38067);
or U39160 (N_39160,N_38533,N_38670);
nor U39161 (N_39161,N_38568,N_38832);
nor U39162 (N_39162,N_38357,N_38952);
xnor U39163 (N_39163,N_38988,N_38609);
nor U39164 (N_39164,N_38190,N_38715);
nand U39165 (N_39165,N_38164,N_38596);
or U39166 (N_39166,N_38779,N_38822);
nor U39167 (N_39167,N_38976,N_38290);
and U39168 (N_39168,N_38614,N_38521);
and U39169 (N_39169,N_38146,N_38059);
or U39170 (N_39170,N_38717,N_38340);
and U39171 (N_39171,N_38322,N_38425);
or U39172 (N_39172,N_38456,N_38053);
or U39173 (N_39173,N_38192,N_38155);
or U39174 (N_39174,N_38361,N_38964);
and U39175 (N_39175,N_38360,N_38218);
xor U39176 (N_39176,N_38234,N_38203);
nand U39177 (N_39177,N_38399,N_38645);
xnor U39178 (N_39178,N_38090,N_38800);
nor U39179 (N_39179,N_38142,N_38035);
nand U39180 (N_39180,N_38181,N_38008);
or U39181 (N_39181,N_38169,N_38556);
nand U39182 (N_39182,N_38069,N_38702);
xor U39183 (N_39183,N_38023,N_38983);
or U39184 (N_39184,N_38525,N_38946);
and U39185 (N_39185,N_38729,N_38416);
nor U39186 (N_39186,N_38426,N_38421);
nor U39187 (N_39187,N_38879,N_38351);
or U39188 (N_39188,N_38668,N_38036);
and U39189 (N_39189,N_38339,N_38337);
and U39190 (N_39190,N_38148,N_38578);
and U39191 (N_39191,N_38631,N_38623);
nand U39192 (N_39192,N_38204,N_38785);
and U39193 (N_39193,N_38435,N_38436);
xor U39194 (N_39194,N_38895,N_38265);
xnor U39195 (N_39195,N_38768,N_38147);
or U39196 (N_39196,N_38540,N_38085);
and U39197 (N_39197,N_38500,N_38264);
and U39198 (N_39198,N_38182,N_38643);
nand U39199 (N_39199,N_38104,N_38597);
or U39200 (N_39200,N_38605,N_38560);
nor U39201 (N_39201,N_38128,N_38347);
nor U39202 (N_39202,N_38119,N_38217);
nand U39203 (N_39203,N_38823,N_38691);
or U39204 (N_39204,N_38350,N_38894);
or U39205 (N_39205,N_38775,N_38712);
or U39206 (N_39206,N_38162,N_38757);
and U39207 (N_39207,N_38959,N_38262);
xor U39208 (N_39208,N_38966,N_38684);
nor U39209 (N_39209,N_38487,N_38573);
or U39210 (N_39210,N_38254,N_38086);
nand U39211 (N_39211,N_38263,N_38117);
nor U39212 (N_39212,N_38394,N_38732);
and U39213 (N_39213,N_38207,N_38071);
or U39214 (N_39214,N_38364,N_38241);
xnor U39215 (N_39215,N_38882,N_38972);
or U39216 (N_39216,N_38222,N_38316);
nand U39217 (N_39217,N_38933,N_38180);
and U39218 (N_39218,N_38226,N_38297);
and U39219 (N_39219,N_38813,N_38970);
nand U39220 (N_39220,N_38948,N_38050);
nor U39221 (N_39221,N_38267,N_38583);
xnor U39222 (N_39222,N_38610,N_38501);
nor U39223 (N_39223,N_38009,N_38856);
xnor U39224 (N_39224,N_38830,N_38716);
and U39225 (N_39225,N_38136,N_38229);
nand U39226 (N_39226,N_38733,N_38314);
or U39227 (N_39227,N_38077,N_38587);
and U39228 (N_39228,N_38273,N_38965);
nor U39229 (N_39229,N_38282,N_38919);
nand U39230 (N_39230,N_38909,N_38140);
nand U39231 (N_39231,N_38513,N_38903);
nand U39232 (N_39232,N_38601,N_38098);
and U39233 (N_39233,N_38096,N_38893);
xor U39234 (N_39234,N_38481,N_38392);
nor U39235 (N_39235,N_38724,N_38133);
nor U39236 (N_39236,N_38621,N_38434);
or U39237 (N_39237,N_38240,N_38786);
xnor U39238 (N_39238,N_38212,N_38930);
or U39239 (N_39239,N_38877,N_38420);
or U39240 (N_39240,N_38170,N_38874);
or U39241 (N_39241,N_38448,N_38808);
xnor U39242 (N_39242,N_38006,N_38276);
and U39243 (N_39243,N_38455,N_38429);
nor U39244 (N_39244,N_38973,N_38607);
xor U39245 (N_39245,N_38331,N_38409);
and U39246 (N_39246,N_38838,N_38728);
nor U39247 (N_39247,N_38175,N_38600);
xnor U39248 (N_39248,N_38236,N_38266);
nor U39249 (N_39249,N_38849,N_38047);
or U39250 (N_39250,N_38588,N_38326);
xor U39251 (N_39251,N_38495,N_38280);
nand U39252 (N_39252,N_38271,N_38888);
nand U39253 (N_39253,N_38644,N_38395);
xor U39254 (N_39254,N_38121,N_38245);
nor U39255 (N_39255,N_38641,N_38239);
xor U39256 (N_39256,N_38256,N_38918);
and U39257 (N_39257,N_38228,N_38431);
and U39258 (N_39258,N_38453,N_38954);
and U39259 (N_39259,N_38798,N_38992);
nand U39260 (N_39260,N_38143,N_38934);
nor U39261 (N_39261,N_38126,N_38805);
nand U39262 (N_39262,N_38235,N_38387);
or U39263 (N_39263,N_38806,N_38561);
or U39264 (N_39264,N_38780,N_38999);
and U39265 (N_39265,N_38827,N_38187);
xnor U39266 (N_39266,N_38868,N_38735);
xor U39267 (N_39267,N_38076,N_38308);
xor U39268 (N_39268,N_38714,N_38007);
xor U39269 (N_39269,N_38734,N_38642);
nor U39270 (N_39270,N_38080,N_38648);
nor U39271 (N_39271,N_38313,N_38811);
nor U39272 (N_39272,N_38807,N_38242);
nor U39273 (N_39273,N_38348,N_38482);
nand U39274 (N_39274,N_38046,N_38437);
xor U39275 (N_39275,N_38799,N_38833);
xnor U39276 (N_39276,N_38744,N_38962);
xor U39277 (N_39277,N_38408,N_38961);
and U39278 (N_39278,N_38160,N_38137);
xor U39279 (N_39279,N_38403,N_38019);
nand U39280 (N_39280,N_38878,N_38102);
xnor U39281 (N_39281,N_38659,N_38474);
nand U39282 (N_39282,N_38951,N_38859);
nand U39283 (N_39283,N_38873,N_38981);
xnor U39284 (N_39284,N_38755,N_38490);
or U39285 (N_39285,N_38527,N_38099);
or U39286 (N_39286,N_38115,N_38907);
nand U39287 (N_39287,N_38810,N_38393);
xnor U39288 (N_39288,N_38458,N_38072);
nor U39289 (N_39289,N_38247,N_38880);
nor U39290 (N_39290,N_38243,N_38045);
or U39291 (N_39291,N_38274,N_38826);
or U39292 (N_39292,N_38884,N_38747);
or U39293 (N_39293,N_38027,N_38995);
nor U39294 (N_39294,N_38159,N_38213);
nor U39295 (N_39295,N_38354,N_38419);
nand U39296 (N_39296,N_38116,N_38442);
and U39297 (N_39297,N_38891,N_38924);
nand U39298 (N_39298,N_38555,N_38377);
nand U39299 (N_39299,N_38200,N_38367);
or U39300 (N_39300,N_38124,N_38378);
or U39301 (N_39301,N_38020,N_38821);
xnor U39302 (N_39302,N_38015,N_38738);
xnor U39303 (N_39303,N_38412,N_38646);
and U39304 (N_39304,N_38819,N_38457);
and U39305 (N_39305,N_38788,N_38269);
nor U39306 (N_39306,N_38246,N_38917);
nand U39307 (N_39307,N_38283,N_38828);
or U39308 (N_39308,N_38718,N_38400);
or U39309 (N_39309,N_38078,N_38796);
nor U39310 (N_39310,N_38492,N_38792);
and U39311 (N_39311,N_38940,N_38195);
and U39312 (N_39312,N_38032,N_38286);
xnor U39313 (N_39313,N_38369,N_38454);
nor U39314 (N_39314,N_38505,N_38382);
and U39315 (N_39315,N_38141,N_38825);
or U39316 (N_39316,N_38277,N_38783);
xnor U39317 (N_39317,N_38151,N_38287);
or U39318 (N_39318,N_38997,N_38809);
or U39319 (N_39319,N_38335,N_38016);
nor U39320 (N_39320,N_38250,N_38837);
and U39321 (N_39321,N_38225,N_38656);
xor U39322 (N_39322,N_38087,N_38391);
nor U39323 (N_39323,N_38673,N_38359);
nor U39324 (N_39324,N_38584,N_38179);
nor U39325 (N_39325,N_38682,N_38026);
xnor U39326 (N_39326,N_38762,N_38622);
and U39327 (N_39327,N_38010,N_38908);
and U39328 (N_39328,N_38184,N_38841);
nand U39329 (N_39329,N_38193,N_38975);
or U39330 (N_39330,N_38336,N_38415);
and U39331 (N_39331,N_38346,N_38955);
xor U39332 (N_39332,N_38498,N_38864);
or U39333 (N_39333,N_38223,N_38925);
and U39334 (N_39334,N_38402,N_38900);
nand U39335 (N_39335,N_38847,N_38685);
nand U39336 (N_39336,N_38091,N_38024);
or U39337 (N_39337,N_38106,N_38520);
and U39338 (N_39338,N_38916,N_38829);
nand U39339 (N_39339,N_38923,N_38606);
nor U39340 (N_39340,N_38514,N_38977);
nand U39341 (N_39341,N_38310,N_38144);
or U39342 (N_39342,N_38761,N_38763);
xor U39343 (N_39343,N_38084,N_38958);
and U39344 (N_39344,N_38386,N_38000);
and U39345 (N_39345,N_38380,N_38048);
nand U39346 (N_39346,N_38284,N_38097);
nand U39347 (N_39347,N_38467,N_38011);
or U39348 (N_39348,N_38161,N_38636);
and U39349 (N_39349,N_38496,N_38650);
nand U39350 (N_39350,N_38820,N_38068);
nand U39351 (N_39351,N_38537,N_38214);
and U39352 (N_39352,N_38544,N_38866);
or U39353 (N_39353,N_38835,N_38066);
nand U39354 (N_39354,N_38194,N_38259);
or U39355 (N_39355,N_38637,N_38885);
xor U39356 (N_39356,N_38703,N_38423);
xnor U39357 (N_39357,N_38473,N_38275);
nor U39358 (N_39358,N_38787,N_38624);
xor U39359 (N_39359,N_38617,N_38485);
nand U39360 (N_39360,N_38338,N_38630);
xnor U39361 (N_39361,N_38634,N_38887);
nor U39362 (N_39362,N_38330,N_38366);
or U39363 (N_39363,N_38215,N_38052);
nand U39364 (N_39364,N_38742,N_38713);
xor U39365 (N_39365,N_38411,N_38901);
xor U39366 (N_39366,N_38611,N_38985);
and U39367 (N_39367,N_38892,N_38307);
xor U39368 (N_39368,N_38508,N_38103);
nor U39369 (N_39369,N_38848,N_38486);
and U39370 (N_39370,N_38176,N_38890);
nand U39371 (N_39371,N_38577,N_38417);
nand U39372 (N_39372,N_38270,N_38831);
and U39373 (N_39373,N_38910,N_38029);
or U39374 (N_39374,N_38599,N_38639);
xor U39375 (N_39375,N_38405,N_38723);
nand U39376 (N_39376,N_38790,N_38095);
or U39377 (N_39377,N_38295,N_38278);
nand U39378 (N_39378,N_38177,N_38469);
nor U39379 (N_39379,N_38815,N_38081);
nand U39380 (N_39380,N_38652,N_38427);
or U39381 (N_39381,N_38928,N_38094);
and U39382 (N_39382,N_38546,N_38296);
xor U39383 (N_39383,N_38863,N_38516);
xnor U39384 (N_39384,N_38157,N_38629);
or U39385 (N_39385,N_38510,N_38818);
and U39386 (N_39386,N_38210,N_38299);
nor U39387 (N_39387,N_38658,N_38677);
and U39388 (N_39388,N_38944,N_38941);
and U39389 (N_39389,N_38003,N_38268);
or U39390 (N_39390,N_38695,N_38237);
or U39391 (N_39391,N_38158,N_38543);
nor U39392 (N_39392,N_38201,N_38497);
or U39393 (N_39393,N_38771,N_38722);
nor U39394 (N_39394,N_38039,N_38483);
and U39395 (N_39395,N_38013,N_38058);
and U39396 (N_39396,N_38370,N_38745);
nor U39397 (N_39397,N_38504,N_38812);
or U39398 (N_39398,N_38342,N_38185);
nor U39399 (N_39399,N_38824,N_38675);
nor U39400 (N_39400,N_38547,N_38679);
or U39401 (N_39401,N_38206,N_38539);
nand U39402 (N_39402,N_38166,N_38870);
nor U39403 (N_39403,N_38589,N_38075);
or U39404 (N_39404,N_38661,N_38936);
and U39405 (N_39405,N_38110,N_38325);
and U39406 (N_39406,N_38332,N_38028);
nor U39407 (N_39407,N_38231,N_38404);
or U39408 (N_39408,N_38773,N_38468);
and U39409 (N_39409,N_38125,N_38686);
or U39410 (N_39410,N_38956,N_38410);
xnor U39411 (N_39411,N_38178,N_38638);
xnor U39412 (N_39412,N_38938,N_38984);
and U39413 (N_39413,N_38802,N_38054);
nor U39414 (N_39414,N_38781,N_38986);
or U39415 (N_39415,N_38769,N_38653);
or U39416 (N_39416,N_38300,N_38082);
and U39417 (N_39417,N_38842,N_38444);
or U39418 (N_39418,N_38982,N_38676);
nand U39419 (N_39419,N_38736,N_38145);
and U39420 (N_39420,N_38198,N_38328);
xor U39421 (N_39421,N_38381,N_38665);
nor U39422 (N_39422,N_38922,N_38522);
and U39423 (N_39423,N_38021,N_38293);
and U39424 (N_39424,N_38433,N_38385);
nor U39425 (N_39425,N_38862,N_38238);
xnor U39426 (N_39426,N_38896,N_38396);
xor U39427 (N_39427,N_38542,N_38953);
or U39428 (N_39428,N_38927,N_38834);
nor U39429 (N_39429,N_38414,N_38022);
nor U39430 (N_39430,N_38739,N_38545);
or U39431 (N_39431,N_38311,N_38153);
nor U39432 (N_39432,N_38680,N_38131);
and U39433 (N_39433,N_38957,N_38018);
nor U39434 (N_39434,N_38291,N_38484);
nand U39435 (N_39435,N_38707,N_38987);
or U39436 (N_39436,N_38693,N_38138);
or U39437 (N_39437,N_38585,N_38580);
nor U39438 (N_39438,N_38005,N_38558);
xnor U39439 (N_39439,N_38571,N_38844);
xnor U39440 (N_39440,N_38122,N_38867);
and U39441 (N_39441,N_38183,N_38551);
and U39442 (N_39442,N_38446,N_38881);
xor U39443 (N_39443,N_38318,N_38305);
and U39444 (N_39444,N_38635,N_38974);
xor U39445 (N_39445,N_38598,N_38857);
or U39446 (N_39446,N_38272,N_38628);
and U39447 (N_39447,N_38897,N_38135);
or U39448 (N_39448,N_38499,N_38784);
or U39449 (N_39449,N_38329,N_38511);
nor U39450 (N_39450,N_38883,N_38899);
or U39451 (N_39451,N_38632,N_38202);
and U39452 (N_39452,N_38764,N_38208);
nand U39453 (N_39453,N_38353,N_38840);
or U39454 (N_39454,N_38662,N_38932);
and U39455 (N_39455,N_38994,N_38731);
xnor U39456 (N_39456,N_38911,N_38906);
and U39457 (N_39457,N_38869,N_38759);
nand U39458 (N_39458,N_38931,N_38978);
xor U39459 (N_39459,N_38920,N_38012);
and U39460 (N_39460,N_38056,N_38109);
or U39461 (N_39461,N_38530,N_38101);
or U39462 (N_39462,N_38671,N_38814);
nor U39463 (N_39463,N_38517,N_38535);
nor U39464 (N_39464,N_38730,N_38341);
and U39465 (N_39465,N_38388,N_38172);
nor U39466 (N_39466,N_38368,N_38156);
or U39467 (N_39467,N_38345,N_38751);
nand U39468 (N_39468,N_38303,N_38655);
nor U39469 (N_39469,N_38220,N_38549);
xor U39470 (N_39470,N_38460,N_38789);
nand U39471 (N_39471,N_38674,N_38450);
or U39472 (N_39472,N_38171,N_38569);
xnor U39473 (N_39473,N_38579,N_38129);
and U39474 (N_39474,N_38061,N_38352);
xor U39475 (N_39475,N_38993,N_38321);
xor U39476 (N_39476,N_38390,N_38132);
and U39477 (N_39477,N_38401,N_38472);
nand U39478 (N_39478,N_38979,N_38244);
nand U39479 (N_39479,N_38615,N_38127);
nor U39480 (N_39480,N_38413,N_38689);
nor U39481 (N_39481,N_38379,N_38969);
nand U39482 (N_39482,N_38518,N_38939);
xnor U39483 (N_39483,N_38108,N_38914);
nand U39484 (N_39484,N_38389,N_38760);
and U39485 (N_39485,N_38189,N_38494);
nand U39486 (N_39486,N_38507,N_38373);
nor U39487 (N_39487,N_38776,N_38465);
or U39488 (N_39488,N_38118,N_38782);
or U39489 (N_39489,N_38640,N_38258);
and U39490 (N_39490,N_38619,N_38509);
and U39491 (N_39491,N_38791,N_38904);
nor U39492 (N_39492,N_38191,N_38963);
or U39493 (N_39493,N_38292,N_38843);
or U39494 (N_39494,N_38384,N_38860);
nand U39495 (N_39495,N_38749,N_38257);
xor U39496 (N_39496,N_38708,N_38461);
nor U39497 (N_39497,N_38541,N_38935);
nor U39498 (N_39498,N_38428,N_38449);
or U39499 (N_39499,N_38727,N_38943);
xnor U39500 (N_39500,N_38381,N_38492);
nand U39501 (N_39501,N_38955,N_38044);
nor U39502 (N_39502,N_38000,N_38400);
nand U39503 (N_39503,N_38556,N_38439);
nand U39504 (N_39504,N_38485,N_38953);
xor U39505 (N_39505,N_38615,N_38967);
or U39506 (N_39506,N_38094,N_38219);
nor U39507 (N_39507,N_38321,N_38769);
and U39508 (N_39508,N_38976,N_38696);
or U39509 (N_39509,N_38824,N_38538);
nor U39510 (N_39510,N_38282,N_38107);
nand U39511 (N_39511,N_38073,N_38209);
xor U39512 (N_39512,N_38827,N_38621);
xor U39513 (N_39513,N_38551,N_38372);
nor U39514 (N_39514,N_38719,N_38519);
nand U39515 (N_39515,N_38688,N_38883);
or U39516 (N_39516,N_38911,N_38879);
or U39517 (N_39517,N_38176,N_38596);
or U39518 (N_39518,N_38909,N_38728);
or U39519 (N_39519,N_38434,N_38706);
xor U39520 (N_39520,N_38309,N_38146);
or U39521 (N_39521,N_38517,N_38556);
or U39522 (N_39522,N_38804,N_38870);
nor U39523 (N_39523,N_38307,N_38328);
xor U39524 (N_39524,N_38220,N_38096);
and U39525 (N_39525,N_38679,N_38496);
or U39526 (N_39526,N_38471,N_38221);
or U39527 (N_39527,N_38454,N_38455);
or U39528 (N_39528,N_38869,N_38784);
nor U39529 (N_39529,N_38487,N_38751);
xnor U39530 (N_39530,N_38604,N_38714);
or U39531 (N_39531,N_38629,N_38217);
and U39532 (N_39532,N_38656,N_38122);
and U39533 (N_39533,N_38895,N_38814);
xnor U39534 (N_39534,N_38948,N_38085);
and U39535 (N_39535,N_38867,N_38978);
nand U39536 (N_39536,N_38051,N_38968);
nand U39537 (N_39537,N_38187,N_38732);
nand U39538 (N_39538,N_38742,N_38006);
and U39539 (N_39539,N_38925,N_38313);
nand U39540 (N_39540,N_38396,N_38613);
and U39541 (N_39541,N_38480,N_38373);
or U39542 (N_39542,N_38261,N_38013);
nand U39543 (N_39543,N_38172,N_38499);
nand U39544 (N_39544,N_38107,N_38505);
xnor U39545 (N_39545,N_38767,N_38937);
xor U39546 (N_39546,N_38944,N_38551);
and U39547 (N_39547,N_38172,N_38474);
nor U39548 (N_39548,N_38063,N_38239);
and U39549 (N_39549,N_38052,N_38228);
xor U39550 (N_39550,N_38755,N_38259);
nand U39551 (N_39551,N_38407,N_38244);
and U39552 (N_39552,N_38090,N_38223);
nor U39553 (N_39553,N_38478,N_38995);
nor U39554 (N_39554,N_38389,N_38839);
nor U39555 (N_39555,N_38101,N_38056);
nor U39556 (N_39556,N_38733,N_38083);
xor U39557 (N_39557,N_38255,N_38032);
xnor U39558 (N_39558,N_38014,N_38549);
nand U39559 (N_39559,N_38374,N_38425);
xor U39560 (N_39560,N_38644,N_38048);
nand U39561 (N_39561,N_38983,N_38881);
or U39562 (N_39562,N_38671,N_38470);
nand U39563 (N_39563,N_38569,N_38643);
or U39564 (N_39564,N_38367,N_38660);
nand U39565 (N_39565,N_38496,N_38897);
and U39566 (N_39566,N_38992,N_38620);
nor U39567 (N_39567,N_38808,N_38278);
nor U39568 (N_39568,N_38214,N_38503);
and U39569 (N_39569,N_38726,N_38481);
xnor U39570 (N_39570,N_38655,N_38962);
nor U39571 (N_39571,N_38044,N_38528);
nor U39572 (N_39572,N_38871,N_38846);
nor U39573 (N_39573,N_38208,N_38123);
xnor U39574 (N_39574,N_38636,N_38808);
nand U39575 (N_39575,N_38488,N_38170);
and U39576 (N_39576,N_38256,N_38933);
or U39577 (N_39577,N_38288,N_38612);
xor U39578 (N_39578,N_38749,N_38174);
or U39579 (N_39579,N_38005,N_38653);
nor U39580 (N_39580,N_38028,N_38916);
nor U39581 (N_39581,N_38428,N_38303);
nor U39582 (N_39582,N_38026,N_38360);
nor U39583 (N_39583,N_38002,N_38815);
nand U39584 (N_39584,N_38418,N_38256);
xor U39585 (N_39585,N_38627,N_38129);
xor U39586 (N_39586,N_38316,N_38620);
nor U39587 (N_39587,N_38786,N_38844);
nor U39588 (N_39588,N_38625,N_38204);
and U39589 (N_39589,N_38580,N_38713);
nor U39590 (N_39590,N_38792,N_38295);
nor U39591 (N_39591,N_38806,N_38786);
and U39592 (N_39592,N_38524,N_38359);
and U39593 (N_39593,N_38119,N_38658);
xnor U39594 (N_39594,N_38609,N_38068);
xnor U39595 (N_39595,N_38499,N_38040);
or U39596 (N_39596,N_38911,N_38319);
nor U39597 (N_39597,N_38550,N_38512);
nor U39598 (N_39598,N_38111,N_38094);
nor U39599 (N_39599,N_38001,N_38933);
or U39600 (N_39600,N_38548,N_38438);
nor U39601 (N_39601,N_38209,N_38947);
or U39602 (N_39602,N_38680,N_38991);
nand U39603 (N_39603,N_38752,N_38565);
nand U39604 (N_39604,N_38012,N_38873);
or U39605 (N_39605,N_38998,N_38409);
nor U39606 (N_39606,N_38191,N_38212);
nor U39607 (N_39607,N_38130,N_38330);
and U39608 (N_39608,N_38883,N_38317);
or U39609 (N_39609,N_38126,N_38067);
or U39610 (N_39610,N_38740,N_38688);
or U39611 (N_39611,N_38305,N_38168);
or U39612 (N_39612,N_38820,N_38593);
xor U39613 (N_39613,N_38571,N_38286);
nand U39614 (N_39614,N_38732,N_38196);
and U39615 (N_39615,N_38982,N_38581);
nand U39616 (N_39616,N_38504,N_38193);
nor U39617 (N_39617,N_38748,N_38861);
xor U39618 (N_39618,N_38188,N_38989);
nand U39619 (N_39619,N_38403,N_38713);
nor U39620 (N_39620,N_38127,N_38383);
nor U39621 (N_39621,N_38777,N_38989);
xor U39622 (N_39622,N_38934,N_38446);
xor U39623 (N_39623,N_38747,N_38707);
nor U39624 (N_39624,N_38864,N_38734);
nand U39625 (N_39625,N_38395,N_38393);
or U39626 (N_39626,N_38255,N_38131);
xor U39627 (N_39627,N_38386,N_38146);
or U39628 (N_39628,N_38053,N_38905);
nor U39629 (N_39629,N_38417,N_38932);
nand U39630 (N_39630,N_38630,N_38520);
nand U39631 (N_39631,N_38650,N_38787);
and U39632 (N_39632,N_38234,N_38910);
xnor U39633 (N_39633,N_38433,N_38493);
xor U39634 (N_39634,N_38353,N_38997);
or U39635 (N_39635,N_38117,N_38236);
and U39636 (N_39636,N_38267,N_38143);
nand U39637 (N_39637,N_38304,N_38224);
or U39638 (N_39638,N_38747,N_38489);
nand U39639 (N_39639,N_38484,N_38856);
or U39640 (N_39640,N_38677,N_38023);
nor U39641 (N_39641,N_38132,N_38512);
or U39642 (N_39642,N_38388,N_38769);
xor U39643 (N_39643,N_38388,N_38801);
nor U39644 (N_39644,N_38476,N_38468);
xor U39645 (N_39645,N_38500,N_38357);
and U39646 (N_39646,N_38558,N_38057);
nor U39647 (N_39647,N_38588,N_38877);
or U39648 (N_39648,N_38463,N_38124);
or U39649 (N_39649,N_38655,N_38531);
xor U39650 (N_39650,N_38770,N_38122);
or U39651 (N_39651,N_38189,N_38996);
or U39652 (N_39652,N_38453,N_38741);
nor U39653 (N_39653,N_38843,N_38167);
nor U39654 (N_39654,N_38823,N_38725);
and U39655 (N_39655,N_38779,N_38520);
and U39656 (N_39656,N_38951,N_38601);
nor U39657 (N_39657,N_38087,N_38474);
xnor U39658 (N_39658,N_38746,N_38768);
xnor U39659 (N_39659,N_38767,N_38971);
nand U39660 (N_39660,N_38618,N_38181);
or U39661 (N_39661,N_38980,N_38396);
and U39662 (N_39662,N_38828,N_38167);
xnor U39663 (N_39663,N_38000,N_38367);
nand U39664 (N_39664,N_38666,N_38398);
xnor U39665 (N_39665,N_38337,N_38627);
nor U39666 (N_39666,N_38045,N_38506);
and U39667 (N_39667,N_38015,N_38254);
and U39668 (N_39668,N_38338,N_38518);
or U39669 (N_39669,N_38938,N_38023);
nand U39670 (N_39670,N_38054,N_38585);
nor U39671 (N_39671,N_38306,N_38678);
and U39672 (N_39672,N_38693,N_38728);
and U39673 (N_39673,N_38310,N_38941);
or U39674 (N_39674,N_38344,N_38288);
nor U39675 (N_39675,N_38642,N_38540);
xnor U39676 (N_39676,N_38180,N_38958);
nor U39677 (N_39677,N_38732,N_38956);
or U39678 (N_39678,N_38264,N_38050);
xnor U39679 (N_39679,N_38797,N_38847);
nor U39680 (N_39680,N_38173,N_38410);
nand U39681 (N_39681,N_38516,N_38683);
nor U39682 (N_39682,N_38936,N_38942);
nor U39683 (N_39683,N_38412,N_38250);
nor U39684 (N_39684,N_38861,N_38066);
nor U39685 (N_39685,N_38861,N_38245);
xnor U39686 (N_39686,N_38053,N_38227);
xor U39687 (N_39687,N_38509,N_38924);
nand U39688 (N_39688,N_38328,N_38973);
and U39689 (N_39689,N_38001,N_38416);
and U39690 (N_39690,N_38728,N_38163);
nor U39691 (N_39691,N_38999,N_38459);
nand U39692 (N_39692,N_38243,N_38273);
and U39693 (N_39693,N_38777,N_38113);
xnor U39694 (N_39694,N_38109,N_38371);
nand U39695 (N_39695,N_38132,N_38021);
nand U39696 (N_39696,N_38945,N_38442);
nand U39697 (N_39697,N_38477,N_38070);
and U39698 (N_39698,N_38873,N_38480);
nor U39699 (N_39699,N_38943,N_38809);
or U39700 (N_39700,N_38071,N_38556);
nand U39701 (N_39701,N_38678,N_38997);
and U39702 (N_39702,N_38149,N_38631);
and U39703 (N_39703,N_38787,N_38918);
nand U39704 (N_39704,N_38231,N_38672);
nor U39705 (N_39705,N_38880,N_38808);
nor U39706 (N_39706,N_38519,N_38540);
xor U39707 (N_39707,N_38846,N_38743);
xor U39708 (N_39708,N_38064,N_38218);
nor U39709 (N_39709,N_38586,N_38657);
nand U39710 (N_39710,N_38053,N_38776);
xor U39711 (N_39711,N_38629,N_38158);
or U39712 (N_39712,N_38733,N_38384);
and U39713 (N_39713,N_38341,N_38661);
xnor U39714 (N_39714,N_38506,N_38808);
xor U39715 (N_39715,N_38154,N_38363);
or U39716 (N_39716,N_38656,N_38319);
xor U39717 (N_39717,N_38404,N_38900);
or U39718 (N_39718,N_38469,N_38517);
or U39719 (N_39719,N_38813,N_38368);
and U39720 (N_39720,N_38613,N_38518);
xor U39721 (N_39721,N_38631,N_38188);
xnor U39722 (N_39722,N_38627,N_38947);
and U39723 (N_39723,N_38068,N_38122);
xor U39724 (N_39724,N_38071,N_38991);
nor U39725 (N_39725,N_38151,N_38730);
nand U39726 (N_39726,N_38155,N_38144);
xnor U39727 (N_39727,N_38422,N_38567);
xor U39728 (N_39728,N_38735,N_38751);
or U39729 (N_39729,N_38990,N_38004);
xor U39730 (N_39730,N_38017,N_38728);
xnor U39731 (N_39731,N_38055,N_38394);
xor U39732 (N_39732,N_38115,N_38570);
xnor U39733 (N_39733,N_38215,N_38695);
nand U39734 (N_39734,N_38855,N_38306);
nand U39735 (N_39735,N_38353,N_38306);
or U39736 (N_39736,N_38300,N_38193);
nor U39737 (N_39737,N_38668,N_38150);
or U39738 (N_39738,N_38384,N_38965);
or U39739 (N_39739,N_38977,N_38903);
or U39740 (N_39740,N_38133,N_38983);
nor U39741 (N_39741,N_38017,N_38026);
nand U39742 (N_39742,N_38293,N_38500);
or U39743 (N_39743,N_38554,N_38768);
nor U39744 (N_39744,N_38696,N_38233);
nor U39745 (N_39745,N_38251,N_38995);
or U39746 (N_39746,N_38316,N_38436);
xor U39747 (N_39747,N_38052,N_38830);
xor U39748 (N_39748,N_38569,N_38126);
nand U39749 (N_39749,N_38906,N_38063);
nand U39750 (N_39750,N_38039,N_38116);
nand U39751 (N_39751,N_38388,N_38254);
nor U39752 (N_39752,N_38999,N_38164);
xor U39753 (N_39753,N_38046,N_38462);
nor U39754 (N_39754,N_38802,N_38462);
or U39755 (N_39755,N_38419,N_38871);
or U39756 (N_39756,N_38641,N_38091);
nor U39757 (N_39757,N_38714,N_38719);
or U39758 (N_39758,N_38109,N_38529);
xor U39759 (N_39759,N_38767,N_38615);
or U39760 (N_39760,N_38479,N_38283);
and U39761 (N_39761,N_38247,N_38565);
xnor U39762 (N_39762,N_38933,N_38906);
xor U39763 (N_39763,N_38465,N_38831);
or U39764 (N_39764,N_38422,N_38569);
or U39765 (N_39765,N_38355,N_38662);
or U39766 (N_39766,N_38412,N_38301);
nor U39767 (N_39767,N_38201,N_38416);
or U39768 (N_39768,N_38224,N_38975);
xnor U39769 (N_39769,N_38528,N_38279);
nand U39770 (N_39770,N_38334,N_38255);
nor U39771 (N_39771,N_38030,N_38565);
and U39772 (N_39772,N_38218,N_38477);
or U39773 (N_39773,N_38748,N_38202);
nor U39774 (N_39774,N_38040,N_38398);
nand U39775 (N_39775,N_38444,N_38323);
and U39776 (N_39776,N_38751,N_38059);
or U39777 (N_39777,N_38945,N_38009);
and U39778 (N_39778,N_38793,N_38105);
and U39779 (N_39779,N_38350,N_38041);
or U39780 (N_39780,N_38901,N_38567);
nor U39781 (N_39781,N_38846,N_38117);
and U39782 (N_39782,N_38877,N_38172);
or U39783 (N_39783,N_38859,N_38350);
and U39784 (N_39784,N_38005,N_38969);
nand U39785 (N_39785,N_38735,N_38296);
nand U39786 (N_39786,N_38236,N_38432);
xnor U39787 (N_39787,N_38436,N_38202);
xnor U39788 (N_39788,N_38228,N_38748);
and U39789 (N_39789,N_38685,N_38301);
xnor U39790 (N_39790,N_38019,N_38428);
and U39791 (N_39791,N_38137,N_38855);
nand U39792 (N_39792,N_38842,N_38131);
nand U39793 (N_39793,N_38909,N_38399);
and U39794 (N_39794,N_38655,N_38375);
nand U39795 (N_39795,N_38176,N_38983);
nor U39796 (N_39796,N_38813,N_38227);
nor U39797 (N_39797,N_38795,N_38394);
and U39798 (N_39798,N_38682,N_38971);
and U39799 (N_39799,N_38618,N_38004);
xor U39800 (N_39800,N_38312,N_38790);
xor U39801 (N_39801,N_38116,N_38219);
nand U39802 (N_39802,N_38179,N_38684);
or U39803 (N_39803,N_38726,N_38362);
nor U39804 (N_39804,N_38777,N_38237);
or U39805 (N_39805,N_38866,N_38233);
xnor U39806 (N_39806,N_38130,N_38180);
or U39807 (N_39807,N_38613,N_38263);
and U39808 (N_39808,N_38231,N_38994);
nand U39809 (N_39809,N_38940,N_38154);
xnor U39810 (N_39810,N_38153,N_38600);
nand U39811 (N_39811,N_38052,N_38884);
xnor U39812 (N_39812,N_38632,N_38901);
nor U39813 (N_39813,N_38110,N_38335);
nand U39814 (N_39814,N_38681,N_38702);
nor U39815 (N_39815,N_38698,N_38524);
xor U39816 (N_39816,N_38574,N_38401);
nor U39817 (N_39817,N_38798,N_38775);
nor U39818 (N_39818,N_38405,N_38318);
or U39819 (N_39819,N_38906,N_38464);
nor U39820 (N_39820,N_38773,N_38925);
xnor U39821 (N_39821,N_38231,N_38241);
or U39822 (N_39822,N_38940,N_38427);
xnor U39823 (N_39823,N_38345,N_38857);
or U39824 (N_39824,N_38601,N_38208);
and U39825 (N_39825,N_38400,N_38041);
xor U39826 (N_39826,N_38695,N_38279);
nor U39827 (N_39827,N_38717,N_38731);
or U39828 (N_39828,N_38404,N_38518);
and U39829 (N_39829,N_38690,N_38004);
nor U39830 (N_39830,N_38047,N_38115);
xor U39831 (N_39831,N_38381,N_38716);
nor U39832 (N_39832,N_38633,N_38582);
nor U39833 (N_39833,N_38194,N_38364);
xnor U39834 (N_39834,N_38741,N_38953);
xnor U39835 (N_39835,N_38126,N_38486);
xor U39836 (N_39836,N_38072,N_38008);
nand U39837 (N_39837,N_38365,N_38410);
nand U39838 (N_39838,N_38434,N_38630);
and U39839 (N_39839,N_38892,N_38402);
nor U39840 (N_39840,N_38541,N_38694);
xor U39841 (N_39841,N_38886,N_38210);
or U39842 (N_39842,N_38544,N_38305);
or U39843 (N_39843,N_38720,N_38478);
xor U39844 (N_39844,N_38283,N_38093);
xnor U39845 (N_39845,N_38579,N_38291);
xnor U39846 (N_39846,N_38538,N_38905);
nand U39847 (N_39847,N_38726,N_38970);
or U39848 (N_39848,N_38242,N_38209);
and U39849 (N_39849,N_38095,N_38744);
nor U39850 (N_39850,N_38665,N_38786);
nand U39851 (N_39851,N_38378,N_38706);
and U39852 (N_39852,N_38100,N_38818);
xnor U39853 (N_39853,N_38152,N_38630);
or U39854 (N_39854,N_38361,N_38505);
and U39855 (N_39855,N_38343,N_38103);
nand U39856 (N_39856,N_38432,N_38167);
nand U39857 (N_39857,N_38816,N_38388);
nor U39858 (N_39858,N_38105,N_38495);
nor U39859 (N_39859,N_38926,N_38513);
nand U39860 (N_39860,N_38147,N_38843);
nand U39861 (N_39861,N_38326,N_38812);
nor U39862 (N_39862,N_38815,N_38177);
nand U39863 (N_39863,N_38967,N_38376);
nand U39864 (N_39864,N_38931,N_38210);
or U39865 (N_39865,N_38434,N_38802);
or U39866 (N_39866,N_38587,N_38417);
and U39867 (N_39867,N_38485,N_38044);
and U39868 (N_39868,N_38115,N_38335);
nor U39869 (N_39869,N_38808,N_38167);
xnor U39870 (N_39870,N_38233,N_38736);
xor U39871 (N_39871,N_38238,N_38058);
or U39872 (N_39872,N_38653,N_38907);
nor U39873 (N_39873,N_38269,N_38461);
and U39874 (N_39874,N_38473,N_38503);
nor U39875 (N_39875,N_38319,N_38510);
nor U39876 (N_39876,N_38708,N_38215);
and U39877 (N_39877,N_38578,N_38919);
nor U39878 (N_39878,N_38177,N_38186);
or U39879 (N_39879,N_38293,N_38254);
or U39880 (N_39880,N_38403,N_38140);
nand U39881 (N_39881,N_38690,N_38993);
nor U39882 (N_39882,N_38097,N_38838);
and U39883 (N_39883,N_38428,N_38580);
and U39884 (N_39884,N_38986,N_38121);
and U39885 (N_39885,N_38838,N_38659);
or U39886 (N_39886,N_38081,N_38168);
xnor U39887 (N_39887,N_38250,N_38156);
nand U39888 (N_39888,N_38442,N_38683);
and U39889 (N_39889,N_38725,N_38784);
or U39890 (N_39890,N_38627,N_38846);
nand U39891 (N_39891,N_38680,N_38443);
nor U39892 (N_39892,N_38683,N_38572);
or U39893 (N_39893,N_38252,N_38243);
nor U39894 (N_39894,N_38595,N_38324);
and U39895 (N_39895,N_38084,N_38378);
xor U39896 (N_39896,N_38344,N_38768);
nand U39897 (N_39897,N_38344,N_38888);
nor U39898 (N_39898,N_38532,N_38462);
nand U39899 (N_39899,N_38067,N_38621);
nand U39900 (N_39900,N_38488,N_38123);
nand U39901 (N_39901,N_38611,N_38517);
or U39902 (N_39902,N_38773,N_38884);
nor U39903 (N_39903,N_38298,N_38989);
nand U39904 (N_39904,N_38090,N_38859);
nor U39905 (N_39905,N_38660,N_38515);
nor U39906 (N_39906,N_38112,N_38131);
xor U39907 (N_39907,N_38984,N_38319);
xor U39908 (N_39908,N_38577,N_38553);
or U39909 (N_39909,N_38613,N_38849);
xor U39910 (N_39910,N_38212,N_38130);
xnor U39911 (N_39911,N_38153,N_38090);
nand U39912 (N_39912,N_38450,N_38018);
nand U39913 (N_39913,N_38764,N_38783);
and U39914 (N_39914,N_38059,N_38836);
or U39915 (N_39915,N_38925,N_38996);
xnor U39916 (N_39916,N_38497,N_38506);
or U39917 (N_39917,N_38808,N_38211);
nand U39918 (N_39918,N_38043,N_38966);
xor U39919 (N_39919,N_38488,N_38229);
xor U39920 (N_39920,N_38443,N_38539);
nor U39921 (N_39921,N_38810,N_38661);
xor U39922 (N_39922,N_38800,N_38779);
xnor U39923 (N_39923,N_38179,N_38343);
nand U39924 (N_39924,N_38118,N_38241);
nor U39925 (N_39925,N_38749,N_38586);
nor U39926 (N_39926,N_38209,N_38961);
or U39927 (N_39927,N_38161,N_38015);
and U39928 (N_39928,N_38661,N_38214);
nor U39929 (N_39929,N_38686,N_38289);
or U39930 (N_39930,N_38983,N_38249);
or U39931 (N_39931,N_38632,N_38446);
or U39932 (N_39932,N_38545,N_38255);
nand U39933 (N_39933,N_38127,N_38473);
nand U39934 (N_39934,N_38206,N_38729);
xor U39935 (N_39935,N_38171,N_38053);
and U39936 (N_39936,N_38185,N_38268);
and U39937 (N_39937,N_38809,N_38637);
and U39938 (N_39938,N_38340,N_38422);
nand U39939 (N_39939,N_38947,N_38813);
and U39940 (N_39940,N_38077,N_38701);
nand U39941 (N_39941,N_38105,N_38977);
nor U39942 (N_39942,N_38828,N_38548);
and U39943 (N_39943,N_38062,N_38245);
nor U39944 (N_39944,N_38524,N_38387);
nor U39945 (N_39945,N_38045,N_38700);
nand U39946 (N_39946,N_38176,N_38390);
xnor U39947 (N_39947,N_38703,N_38478);
nand U39948 (N_39948,N_38590,N_38388);
nand U39949 (N_39949,N_38966,N_38440);
nand U39950 (N_39950,N_38107,N_38758);
xnor U39951 (N_39951,N_38750,N_38749);
xnor U39952 (N_39952,N_38528,N_38297);
or U39953 (N_39953,N_38594,N_38021);
xor U39954 (N_39954,N_38699,N_38349);
and U39955 (N_39955,N_38572,N_38331);
nand U39956 (N_39956,N_38898,N_38694);
and U39957 (N_39957,N_38768,N_38565);
nor U39958 (N_39958,N_38591,N_38848);
nor U39959 (N_39959,N_38372,N_38356);
or U39960 (N_39960,N_38312,N_38543);
and U39961 (N_39961,N_38822,N_38572);
nor U39962 (N_39962,N_38059,N_38742);
or U39963 (N_39963,N_38185,N_38474);
or U39964 (N_39964,N_38847,N_38361);
xor U39965 (N_39965,N_38714,N_38542);
nor U39966 (N_39966,N_38513,N_38389);
nor U39967 (N_39967,N_38865,N_38033);
xnor U39968 (N_39968,N_38504,N_38634);
nor U39969 (N_39969,N_38280,N_38219);
and U39970 (N_39970,N_38937,N_38201);
or U39971 (N_39971,N_38220,N_38635);
xnor U39972 (N_39972,N_38477,N_38344);
nor U39973 (N_39973,N_38242,N_38222);
nand U39974 (N_39974,N_38516,N_38084);
xnor U39975 (N_39975,N_38859,N_38412);
nand U39976 (N_39976,N_38989,N_38060);
nor U39977 (N_39977,N_38255,N_38677);
or U39978 (N_39978,N_38188,N_38801);
nor U39979 (N_39979,N_38183,N_38027);
and U39980 (N_39980,N_38224,N_38872);
nor U39981 (N_39981,N_38912,N_38286);
nand U39982 (N_39982,N_38595,N_38840);
and U39983 (N_39983,N_38403,N_38689);
xnor U39984 (N_39984,N_38288,N_38905);
or U39985 (N_39985,N_38901,N_38805);
nor U39986 (N_39986,N_38039,N_38388);
or U39987 (N_39987,N_38081,N_38290);
nor U39988 (N_39988,N_38307,N_38103);
nand U39989 (N_39989,N_38927,N_38700);
nand U39990 (N_39990,N_38926,N_38109);
xnor U39991 (N_39991,N_38909,N_38908);
xnor U39992 (N_39992,N_38638,N_38205);
and U39993 (N_39993,N_38274,N_38257);
nor U39994 (N_39994,N_38476,N_38220);
nand U39995 (N_39995,N_38327,N_38502);
nand U39996 (N_39996,N_38153,N_38847);
xnor U39997 (N_39997,N_38911,N_38259);
or U39998 (N_39998,N_38418,N_38914);
or U39999 (N_39999,N_38649,N_38444);
or U40000 (N_40000,N_39337,N_39405);
nand U40001 (N_40001,N_39835,N_39294);
xor U40002 (N_40002,N_39624,N_39872);
or U40003 (N_40003,N_39332,N_39052);
nand U40004 (N_40004,N_39787,N_39164);
xnor U40005 (N_40005,N_39860,N_39087);
nand U40006 (N_40006,N_39029,N_39976);
nor U40007 (N_40007,N_39113,N_39211);
or U40008 (N_40008,N_39418,N_39383);
and U40009 (N_40009,N_39119,N_39913);
nand U40010 (N_40010,N_39465,N_39990);
or U40011 (N_40011,N_39472,N_39669);
or U40012 (N_40012,N_39583,N_39060);
or U40013 (N_40013,N_39174,N_39981);
nor U40014 (N_40014,N_39566,N_39628);
xnor U40015 (N_40015,N_39637,N_39414);
xor U40016 (N_40016,N_39996,N_39995);
nor U40017 (N_40017,N_39058,N_39593);
or U40018 (N_40018,N_39623,N_39235);
or U40019 (N_40019,N_39469,N_39030);
and U40020 (N_40020,N_39042,N_39272);
or U40021 (N_40021,N_39543,N_39240);
or U40022 (N_40022,N_39947,N_39803);
and U40023 (N_40023,N_39175,N_39117);
nor U40024 (N_40024,N_39424,N_39810);
nand U40025 (N_40025,N_39054,N_39553);
or U40026 (N_40026,N_39367,N_39843);
nor U40027 (N_40027,N_39766,N_39892);
xnor U40028 (N_40028,N_39186,N_39894);
xor U40029 (N_40029,N_39541,N_39570);
and U40030 (N_40030,N_39417,N_39299);
nand U40031 (N_40031,N_39846,N_39551);
or U40032 (N_40032,N_39490,N_39396);
xnor U40033 (N_40033,N_39244,N_39330);
nand U40034 (N_40034,N_39497,N_39676);
nor U40035 (N_40035,N_39454,N_39525);
nor U40036 (N_40036,N_39813,N_39256);
nor U40037 (N_40037,N_39094,N_39865);
nor U40038 (N_40038,N_39612,N_39136);
nand U40039 (N_40039,N_39851,N_39768);
or U40040 (N_40040,N_39677,N_39730);
or U40041 (N_40041,N_39779,N_39538);
nor U40042 (N_40042,N_39507,N_39021);
nand U40043 (N_40043,N_39190,N_39982);
xnor U40044 (N_40044,N_39125,N_39671);
nor U40045 (N_40045,N_39301,N_39882);
xor U40046 (N_40046,N_39084,N_39934);
xor U40047 (N_40047,N_39361,N_39009);
xor U40048 (N_40048,N_39091,N_39733);
and U40049 (N_40049,N_39399,N_39078);
nor U40050 (N_40050,N_39505,N_39287);
or U40051 (N_40051,N_39620,N_39528);
xor U40052 (N_40052,N_39834,N_39395);
and U40053 (N_40053,N_39280,N_39877);
xnor U40054 (N_40054,N_39617,N_39740);
xor U40055 (N_40055,N_39736,N_39679);
nor U40056 (N_40056,N_39110,N_39043);
xnor U40057 (N_40057,N_39828,N_39868);
or U40058 (N_40058,N_39710,N_39071);
nor U40059 (N_40059,N_39121,N_39576);
nand U40060 (N_40060,N_39216,N_39440);
and U40061 (N_40061,N_39019,N_39005);
and U40062 (N_40062,N_39602,N_39459);
xor U40063 (N_40063,N_39638,N_39461);
nor U40064 (N_40064,N_39821,N_39520);
or U40065 (N_40065,N_39426,N_39375);
and U40066 (N_40066,N_39652,N_39758);
nand U40067 (N_40067,N_39006,N_39312);
nor U40068 (N_40068,N_39184,N_39519);
xnor U40069 (N_40069,N_39518,N_39967);
or U40070 (N_40070,N_39802,N_39928);
or U40071 (N_40071,N_39784,N_39951);
xor U40072 (N_40072,N_39082,N_39309);
and U40073 (N_40073,N_39295,N_39757);
or U40074 (N_40074,N_39448,N_39980);
nand U40075 (N_40075,N_39717,N_39713);
or U40076 (N_40076,N_39942,N_39975);
nor U40077 (N_40077,N_39999,N_39728);
nand U40078 (N_40078,N_39269,N_39419);
nand U40079 (N_40079,N_39754,N_39065);
and U40080 (N_40080,N_39645,N_39989);
and U40081 (N_40081,N_39031,N_39798);
nor U40082 (N_40082,N_39574,N_39756);
nand U40083 (N_40083,N_39722,N_39083);
or U40084 (N_40084,N_39516,N_39561);
nor U40085 (N_40085,N_39857,N_39388);
nand U40086 (N_40086,N_39304,N_39435);
nor U40087 (N_40087,N_39836,N_39242);
or U40088 (N_40088,N_39711,N_39342);
and U40089 (N_40089,N_39935,N_39438);
or U40090 (N_40090,N_39883,N_39946);
nand U40091 (N_40091,N_39000,N_39780);
or U40092 (N_40092,N_39849,N_39051);
nor U40093 (N_40093,N_39111,N_39323);
and U40094 (N_40094,N_39526,N_39255);
nor U40095 (N_40095,N_39221,N_39471);
and U40096 (N_40096,N_39511,N_39558);
nand U40097 (N_40097,N_39866,N_39959);
nor U40098 (N_40098,N_39326,N_39983);
nor U40099 (N_40099,N_39365,N_39613);
nand U40100 (N_40100,N_39694,N_39243);
and U40101 (N_40101,N_39675,N_39660);
xor U40102 (N_40102,N_39099,N_39270);
xor U40103 (N_40103,N_39131,N_39151);
and U40104 (N_40104,N_39993,N_39837);
or U40105 (N_40105,N_39986,N_39708);
or U40106 (N_40106,N_39037,N_39143);
and U40107 (N_40107,N_39283,N_39259);
xor U40108 (N_40108,N_39004,N_39806);
nor U40109 (N_40109,N_39841,N_39463);
nor U40110 (N_40110,N_39819,N_39066);
or U40111 (N_40111,N_39443,N_39619);
nor U40112 (N_40112,N_39689,N_39929);
and U40113 (N_40113,N_39489,N_39402);
and U40114 (N_40114,N_39902,N_39478);
xor U40115 (N_40115,N_39401,N_39978);
nand U40116 (N_40116,N_39362,N_39218);
xnor U40117 (N_40117,N_39715,N_39812);
xor U40118 (N_40118,N_39321,N_39686);
nor U40119 (N_40119,N_39556,N_39804);
or U40120 (N_40120,N_39941,N_39276);
nor U40121 (N_40121,N_39925,N_39464);
and U40122 (N_40122,N_39124,N_39963);
nand U40123 (N_40123,N_39739,N_39920);
nor U40124 (N_40124,N_39200,N_39373);
nor U40125 (N_40125,N_39562,N_39759);
and U40126 (N_40126,N_39250,N_39842);
nand U40127 (N_40127,N_39010,N_39354);
nor U40128 (N_40128,N_39477,N_39227);
and U40129 (N_40129,N_39041,N_39668);
nor U40130 (N_40130,N_39302,N_39639);
and U40131 (N_40131,N_39927,N_39161);
and U40132 (N_40132,N_39232,N_39888);
xnor U40133 (N_40133,N_39411,N_39932);
nor U40134 (N_40134,N_39564,N_39410);
or U40135 (N_40135,N_39264,N_39634);
nor U40136 (N_40136,N_39884,N_39277);
nand U40137 (N_40137,N_39069,N_39421);
and U40138 (N_40138,N_39171,N_39392);
nand U40139 (N_40139,N_39653,N_39745);
or U40140 (N_40140,N_39817,N_39486);
xor U40141 (N_40141,N_39288,N_39147);
xor U40142 (N_40142,N_39627,N_39056);
nor U40143 (N_40143,N_39987,N_39297);
xor U40144 (N_40144,N_39921,N_39788);
nor U40145 (N_40145,N_39618,N_39797);
nor U40146 (N_40146,N_39933,N_39429);
nor U40147 (N_40147,N_39595,N_39891);
nand U40148 (N_40148,N_39662,N_39633);
and U40149 (N_40149,N_39859,N_39948);
nor U40150 (N_40150,N_39425,N_39251);
xnor U40151 (N_40151,N_39818,N_39449);
nand U40152 (N_40152,N_39610,N_39239);
nor U40153 (N_40153,N_39345,N_39917);
nor U40154 (N_40154,N_39257,N_39880);
nand U40155 (N_40155,N_39651,N_39353);
and U40156 (N_40156,N_39844,N_39038);
nand U40157 (N_40157,N_39546,N_39318);
and U40158 (N_40158,N_39278,N_39643);
and U40159 (N_40159,N_39580,N_39830);
nand U40160 (N_40160,N_39195,N_39632);
nand U40161 (N_40161,N_39355,N_39444);
xnor U40162 (N_40162,N_39327,N_39437);
and U40163 (N_40163,N_39391,N_39020);
nor U40164 (N_40164,N_39678,N_39086);
and U40165 (N_40165,N_39075,N_39485);
or U40166 (N_40166,N_39688,N_39807);
nor U40167 (N_40167,N_39303,N_39744);
or U40168 (N_40168,N_39696,N_39977);
and U40169 (N_40169,N_39336,N_39625);
nand U40170 (N_40170,N_39879,N_39560);
nand U40171 (N_40171,N_39389,N_39045);
nand U40172 (N_40172,N_39994,N_39382);
nor U40173 (N_40173,N_39053,N_39313);
or U40174 (N_40174,N_39349,N_39281);
or U40175 (N_40175,N_39607,N_39260);
xor U40176 (N_40176,N_39245,N_39498);
xor U40177 (N_40177,N_39363,N_39441);
nor U40178 (N_40178,N_39827,N_39666);
and U40179 (N_40179,N_39796,N_39286);
xnor U40180 (N_40180,N_39199,N_39371);
xnor U40181 (N_40181,N_39964,N_39621);
and U40182 (N_40182,N_39014,N_39016);
and U40183 (N_40183,N_39919,N_39222);
nand U40184 (N_40184,N_39296,N_39291);
nand U40185 (N_40185,N_39614,N_39504);
nand U40186 (N_40186,N_39700,N_39755);
nor U40187 (N_40187,N_39611,N_39413);
or U40188 (N_40188,N_39962,N_39537);
nor U40189 (N_40189,N_39816,N_39753);
and U40190 (N_40190,N_39196,N_39059);
or U40191 (N_40191,N_39875,N_39547);
or U40192 (N_40192,N_39070,N_39629);
and U40193 (N_40193,N_39462,N_39018);
nor U40194 (N_40194,N_39185,N_39166);
nor U40195 (N_40195,N_39521,N_39542);
xor U40196 (N_40196,N_39726,N_39731);
nand U40197 (N_40197,N_39737,N_39776);
xnor U40198 (N_40198,N_39039,N_39640);
nand U40199 (N_40199,N_39017,N_39115);
and U40200 (N_40200,N_39529,N_39198);
and U40201 (N_40201,N_39792,N_39565);
nand U40202 (N_40202,N_39957,N_39644);
nor U40203 (N_40203,N_39535,N_39635);
nor U40204 (N_40204,N_39552,N_39144);
or U40205 (N_40205,N_39606,N_39252);
nand U40206 (N_40206,N_39032,N_39394);
xor U40207 (N_40207,N_39012,N_39109);
nand U40208 (N_40208,N_39145,N_39630);
and U40209 (N_40209,N_39126,N_39589);
nand U40210 (N_40210,N_39522,N_39135);
and U40211 (N_40211,N_39956,N_39467);
or U40212 (N_40212,N_39366,N_39578);
or U40213 (N_40213,N_39046,N_39530);
or U40214 (N_40214,N_39025,N_39335);
xor U40215 (N_40215,N_39263,N_39899);
nor U40216 (N_40216,N_39442,N_39539);
or U40217 (N_40217,N_39400,N_39081);
or U40218 (N_40218,N_39887,N_39709);
nand U40219 (N_40219,N_39746,N_39149);
nand U40220 (N_40220,N_39773,N_39393);
or U40221 (N_40221,N_39725,N_39153);
nand U40222 (N_40222,N_39955,N_39930);
or U40223 (N_40223,N_39064,N_39491);
nor U40224 (N_40224,N_39650,N_39738);
nor U40225 (N_40225,N_39923,N_39910);
and U40226 (N_40226,N_39483,N_39191);
xor U40227 (N_40227,N_39150,N_39063);
and U40228 (N_40228,N_39512,N_39501);
or U40229 (N_40229,N_39428,N_39750);
xor U40230 (N_40230,N_39238,N_39447);
nor U40231 (N_40231,N_39517,N_39712);
xnor U40232 (N_40232,N_39789,N_39549);
xnor U40233 (N_40233,N_39210,N_39101);
nand U40234 (N_40234,N_39889,N_39890);
and U40235 (N_40235,N_39307,N_39436);
nand U40236 (N_40236,N_39116,N_39322);
nor U40237 (N_40237,N_39456,N_39748);
nand U40238 (N_40238,N_39961,N_39601);
and U40239 (N_40239,N_39687,N_39495);
nor U40240 (N_40240,N_39333,N_39331);
and U40241 (N_40241,N_39655,N_39735);
nand U40242 (N_40242,N_39432,N_39201);
or U40243 (N_40243,N_39673,N_39188);
or U40244 (N_40244,N_39905,N_39108);
and U40245 (N_40245,N_39824,N_39893);
nor U40246 (N_40246,N_39112,N_39514);
and U40247 (N_40247,N_39189,N_39914);
or U40248 (N_40248,N_39699,N_39691);
nand U40249 (N_40249,N_39104,N_39197);
xor U40250 (N_40250,N_39204,N_39954);
and U40251 (N_40251,N_39953,N_39540);
or U40252 (N_40252,N_39702,N_39672);
nor U40253 (N_40253,N_39845,N_39767);
and U40254 (N_40254,N_39506,N_39073);
xnor U40255 (N_40255,N_39647,N_39002);
and U40256 (N_40256,N_39008,N_39596);
and U40257 (N_40257,N_39412,N_39509);
or U40258 (N_40258,N_39918,N_39581);
and U40259 (N_40259,N_39575,N_39369);
nand U40260 (N_40260,N_39106,N_39968);
nor U40261 (N_40261,N_39300,N_39832);
nand U40262 (N_40262,N_39714,N_39001);
nand U40263 (N_40263,N_39984,N_39028);
xor U40264 (N_40264,N_39765,N_39912);
nand U40265 (N_40265,N_39707,N_39727);
nor U40266 (N_40266,N_39723,N_39455);
nor U40267 (N_40267,N_39206,N_39568);
or U40268 (N_40268,N_39949,N_39873);
nor U40269 (N_40269,N_39503,N_39183);
xnor U40270 (N_40270,N_39027,N_39194);
xor U40271 (N_40271,N_39178,N_39203);
nor U40272 (N_40272,N_39446,N_39998);
or U40273 (N_40273,N_39579,N_39434);
nor U40274 (N_40274,N_39907,N_39062);
or U40275 (N_40275,N_39352,N_39681);
and U40276 (N_40276,N_39034,N_39850);
nor U40277 (N_40277,N_39572,N_39657);
and U40278 (N_40278,N_39217,N_39351);
xor U40279 (N_40279,N_39690,N_39513);
and U40280 (N_40280,N_39732,N_39093);
nand U40281 (N_40281,N_39372,N_39403);
nand U40282 (N_40282,N_39481,N_39114);
or U40283 (N_40283,N_39105,N_39786);
or U40284 (N_40284,N_39800,N_39328);
or U40285 (N_40285,N_39406,N_39636);
and U40286 (N_40286,N_39534,N_39665);
and U40287 (N_40287,N_39305,N_39407);
or U40288 (N_40288,N_39176,N_39600);
and U40289 (N_40289,N_39790,N_39015);
nand U40290 (N_40290,N_39049,N_39329);
nor U40291 (N_40291,N_39654,N_39840);
nand U40292 (N_40292,N_39897,N_39292);
and U40293 (N_40293,N_39128,N_39182);
or U40294 (N_40294,N_39230,N_39480);
or U40295 (N_40295,N_39316,N_39903);
and U40296 (N_40296,N_39778,N_39152);
nor U40297 (N_40297,N_39848,N_39508);
xnor U40298 (N_40298,N_39346,N_39311);
and U40299 (N_40299,N_39777,N_39663);
or U40300 (N_40300,N_39626,N_39347);
xor U40301 (N_40301,N_39500,N_39704);
nor U40302 (N_40302,N_39939,N_39805);
or U40303 (N_40303,N_39420,N_39076);
and U40304 (N_40304,N_39165,N_39167);
nand U40305 (N_40305,N_39341,N_39588);
or U40306 (N_40306,N_39271,N_39548);
and U40307 (N_40307,N_39047,N_39493);
or U40308 (N_40308,N_39384,N_39077);
nor U40309 (N_40309,N_39555,N_39095);
nand U40310 (N_40310,N_39473,N_39705);
nor U40311 (N_40311,N_39979,N_39847);
or U40312 (N_40312,N_39692,N_39385);
nand U40313 (N_40313,N_39192,N_39901);
and U40314 (N_40314,N_39213,N_39864);
nor U40315 (N_40315,N_39215,N_39088);
nand U40316 (N_40316,N_39867,N_39282);
xnor U40317 (N_40317,N_39599,N_39033);
and U40318 (N_40318,N_39229,N_39772);
or U40319 (N_40319,N_39915,N_39139);
xnor U40320 (N_40320,N_39181,N_39854);
xor U40321 (N_40321,N_39693,N_39874);
nor U40322 (N_40322,N_39180,N_39761);
nor U40323 (N_40323,N_39762,N_39487);
or U40324 (N_40324,N_39582,N_39340);
xor U40325 (N_40325,N_39187,N_39376);
nand U40326 (N_40326,N_39499,N_39074);
nor U40327 (N_40327,N_39571,N_39157);
nand U40328 (N_40328,N_39496,N_39785);
xnor U40329 (N_40329,N_39764,N_39958);
nor U40330 (N_40330,N_39390,N_39701);
nor U40331 (N_40331,N_39439,N_39616);
or U40332 (N_40332,N_39682,N_39168);
and U40333 (N_40333,N_39950,N_39224);
nor U40334 (N_40334,N_39118,N_39922);
nand U40335 (N_40335,N_39140,N_39752);
nor U40336 (N_40336,N_39985,N_39855);
xor U40337 (N_40337,N_39973,N_39479);
xor U40338 (N_40338,N_39743,N_39348);
nand U40339 (N_40339,N_39044,N_39484);
nand U40340 (N_40340,N_39885,N_39386);
nand U40341 (N_40341,N_39554,N_39703);
xnor U40342 (N_40342,N_39916,N_39408);
nor U40343 (N_40343,N_39760,N_39475);
nand U40344 (N_40344,N_39254,N_39524);
nor U40345 (N_40345,N_39067,N_39670);
nand U40346 (N_40346,N_39097,N_39308);
xnor U40347 (N_40347,N_39404,N_39246);
nand U40348 (N_40348,N_39965,N_39011);
or U40349 (N_40349,N_39133,N_39173);
or U40350 (N_40350,N_39148,N_39527);
xor U40351 (N_40351,N_39862,N_39234);
nand U40352 (N_40352,N_39544,N_39380);
nor U40353 (N_40353,N_39236,N_39586);
nand U40354 (N_40354,N_39172,N_39969);
xor U40355 (N_40355,N_39368,N_39557);
nand U40356 (N_40356,N_39100,N_39207);
xnor U40357 (N_40357,N_39974,N_39577);
and U40358 (N_40358,N_39466,N_39594);
or U40359 (N_40359,N_39022,N_39631);
nor U40360 (N_40360,N_39971,N_39724);
nor U40361 (N_40361,N_39991,N_39770);
nand U40362 (N_40362,N_39488,N_39266);
nor U40363 (N_40363,N_39035,N_39988);
nor U40364 (N_40364,N_39036,N_39261);
xnor U40365 (N_40365,N_39815,N_39603);
and U40366 (N_40366,N_39158,N_39944);
or U40367 (N_40367,N_39068,N_39926);
xor U40368 (N_40368,N_39820,N_39646);
or U40369 (N_40369,N_39584,N_39782);
and U40370 (N_40370,N_39334,N_39608);
or U40371 (N_40371,N_39852,N_39876);
nor U40372 (N_40372,N_39451,N_39642);
xnor U40373 (N_40373,N_39729,N_39262);
nand U40374 (N_40374,N_39683,N_39559);
or U40375 (N_40375,N_39536,N_39226);
nand U40376 (N_40376,N_39641,N_39409);
xnor U40377 (N_40377,N_39205,N_39248);
nand U40378 (N_40378,N_39751,N_39344);
xnor U40379 (N_40379,N_39055,N_39123);
and U40380 (N_40380,N_39381,N_39374);
nand U40381 (N_40381,N_39057,N_39871);
or U40382 (N_40382,N_39658,N_39900);
or U40383 (N_40383,N_39127,N_39040);
and U40384 (N_40384,N_39587,N_39179);
xnor U40385 (N_40385,N_39208,N_39268);
or U40386 (N_40386,N_39431,N_39911);
nand U40387 (N_40387,N_39833,N_39853);
nor U40388 (N_40388,N_39997,N_39156);
nor U40389 (N_40389,N_39622,N_39881);
or U40390 (N_40390,N_39719,N_39482);
nand U40391 (N_40391,N_39339,N_39120);
nor U40392 (N_40392,N_39423,N_39427);
xnor U40393 (N_40393,N_39285,N_39648);
and U40394 (N_40394,N_39769,N_39096);
and U40395 (N_40395,N_39952,N_39476);
or U40396 (N_40396,N_39741,N_39159);
xor U40397 (N_40397,N_39155,N_39775);
nor U40398 (N_40398,N_39253,N_39398);
or U40399 (N_40399,N_39122,N_39839);
and U40400 (N_40400,N_39154,N_39350);
or U40401 (N_40401,N_39450,N_39293);
or U40402 (N_40402,N_39415,N_39233);
nand U40403 (N_40403,N_39898,N_39823);
or U40404 (N_40404,N_39664,N_39290);
or U40405 (N_40405,N_39799,N_39494);
nor U40406 (N_40406,N_39960,N_39904);
and U40407 (N_40407,N_39430,N_39649);
nand U40408 (N_40408,N_39924,N_39468);
and U40409 (N_40409,N_39275,N_39258);
nand U40410 (N_40410,N_39397,N_39667);
nor U40411 (N_40411,N_39138,N_39416);
and U40412 (N_40412,N_39680,N_39085);
or U40413 (N_40413,N_39433,N_39089);
nor U40414 (N_40414,N_39223,N_39202);
xor U40415 (N_40415,N_39134,N_39163);
nor U40416 (N_40416,N_39567,N_39858);
and U40417 (N_40417,N_39209,N_39357);
and U40418 (N_40418,N_39314,N_39747);
or U40419 (N_40419,N_39231,N_39869);
nand U40420 (N_40420,N_39510,N_39310);
or U40421 (N_40421,N_39825,N_39050);
nor U40422 (N_40422,N_39377,N_39720);
nor U40423 (N_40423,N_39938,N_39007);
and U40424 (N_40424,N_39169,N_39598);
and U40425 (N_40425,N_39228,N_39225);
and U40426 (N_40426,N_39791,N_39170);
nand U40427 (N_40427,N_39458,N_39177);
nand U40428 (N_40428,N_39793,N_39515);
nor U40429 (N_40429,N_39605,N_39364);
or U40430 (N_40430,N_39160,N_39861);
xor U40431 (N_40431,N_39742,N_39289);
and U40432 (N_40432,N_39453,N_39107);
or U40433 (N_40433,N_39298,N_39763);
nand U40434 (N_40434,N_39319,N_39721);
or U40435 (N_40435,N_39695,N_39531);
or U40436 (N_40436,N_39597,N_39870);
nand U40437 (N_40437,N_39931,N_39343);
xnor U40438 (N_40438,N_39906,N_39360);
xor U40439 (N_40439,N_39214,N_39102);
or U40440 (N_40440,N_39718,N_39706);
nor U40441 (N_40441,N_39220,N_39822);
and U40442 (N_40442,N_39716,N_39265);
nand U40443 (N_40443,N_39137,N_39684);
and U40444 (N_40444,N_39972,N_39129);
nor U40445 (N_40445,N_39826,N_39532);
nor U40446 (N_40446,N_39545,N_39162);
xnor U40447 (N_40447,N_39359,N_39609);
nand U40448 (N_40448,N_39685,N_39966);
xor U40449 (N_40449,N_39338,N_39940);
or U40450 (N_40450,N_39098,N_39387);
nor U40451 (N_40451,N_39771,N_39146);
nand U40452 (N_40452,N_39838,N_39697);
nand U40453 (N_40453,N_39615,N_39219);
or U40454 (N_40454,N_39563,N_39674);
nor U40455 (N_40455,N_39460,N_39237);
and U40456 (N_40456,N_39774,N_39550);
xor U40457 (N_40457,N_39783,N_39422);
nand U40458 (N_40458,N_39523,N_39474);
nand U40459 (N_40459,N_39279,N_39781);
and U40460 (N_40460,N_39943,N_39795);
and U40461 (N_40461,N_39734,N_39132);
nor U40462 (N_40462,N_39061,N_39585);
xor U40463 (N_40463,N_39325,N_39856);
nand U40464 (N_40464,N_39315,N_39809);
nor U40465 (N_40465,N_39698,N_39013);
nand U40466 (N_40466,N_39130,N_39533);
nand U40467 (N_40467,N_39592,N_39080);
nand U40468 (N_40468,N_39378,N_39142);
nand U40469 (N_40469,N_39604,N_39445);
xor U40470 (N_40470,N_39814,N_39896);
xnor U40471 (N_40471,N_39886,N_39659);
and U40472 (N_40472,N_39267,N_39141);
nor U40473 (N_40473,N_39452,N_39811);
or U40474 (N_40474,N_39249,N_39024);
xnor U40475 (N_40475,N_39241,N_39808);
nor U40476 (N_40476,N_39026,N_39457);
and U40477 (N_40477,N_39358,N_39831);
and U40478 (N_40478,N_39306,N_39284);
nand U40479 (N_40479,N_39212,N_39023);
nand U40480 (N_40480,N_39656,N_39749);
xnor U40481 (N_40481,N_39569,N_39320);
or U40482 (N_40482,N_39379,N_39324);
nor U40483 (N_40483,N_39794,N_39048);
xnor U40484 (N_40484,N_39492,N_39247);
xor U40485 (N_40485,N_39003,N_39661);
or U40486 (N_40486,N_39072,N_39092);
nor U40487 (N_40487,N_39829,N_39193);
and U40488 (N_40488,N_39937,N_39273);
or U40489 (N_40489,N_39936,N_39863);
and U40490 (N_40490,N_39590,N_39370);
nand U40491 (N_40491,N_39090,N_39274);
and U40492 (N_40492,N_39591,N_39908);
nor U40493 (N_40493,N_39317,N_39970);
xor U40494 (N_40494,N_39356,N_39502);
and U40495 (N_40495,N_39895,N_39470);
or U40496 (N_40496,N_39992,N_39573);
and U40497 (N_40497,N_39079,N_39945);
or U40498 (N_40498,N_39909,N_39801);
xor U40499 (N_40499,N_39878,N_39103);
or U40500 (N_40500,N_39865,N_39982);
or U40501 (N_40501,N_39309,N_39319);
xnor U40502 (N_40502,N_39663,N_39791);
xor U40503 (N_40503,N_39635,N_39912);
xor U40504 (N_40504,N_39555,N_39843);
and U40505 (N_40505,N_39190,N_39424);
or U40506 (N_40506,N_39034,N_39674);
nand U40507 (N_40507,N_39704,N_39154);
nor U40508 (N_40508,N_39131,N_39159);
xor U40509 (N_40509,N_39813,N_39176);
nand U40510 (N_40510,N_39964,N_39278);
nand U40511 (N_40511,N_39369,N_39780);
and U40512 (N_40512,N_39690,N_39250);
nand U40513 (N_40513,N_39433,N_39323);
nand U40514 (N_40514,N_39111,N_39754);
nor U40515 (N_40515,N_39656,N_39489);
nor U40516 (N_40516,N_39078,N_39943);
nand U40517 (N_40517,N_39362,N_39987);
nor U40518 (N_40518,N_39359,N_39349);
or U40519 (N_40519,N_39046,N_39402);
nand U40520 (N_40520,N_39104,N_39224);
nor U40521 (N_40521,N_39294,N_39593);
or U40522 (N_40522,N_39972,N_39099);
nand U40523 (N_40523,N_39480,N_39952);
xnor U40524 (N_40524,N_39735,N_39616);
xnor U40525 (N_40525,N_39739,N_39156);
xnor U40526 (N_40526,N_39435,N_39099);
xnor U40527 (N_40527,N_39951,N_39603);
nor U40528 (N_40528,N_39066,N_39621);
nor U40529 (N_40529,N_39191,N_39911);
nor U40530 (N_40530,N_39276,N_39477);
nand U40531 (N_40531,N_39338,N_39791);
xnor U40532 (N_40532,N_39683,N_39089);
nor U40533 (N_40533,N_39250,N_39955);
nor U40534 (N_40534,N_39193,N_39445);
nand U40535 (N_40535,N_39815,N_39707);
xnor U40536 (N_40536,N_39766,N_39731);
or U40537 (N_40537,N_39685,N_39372);
nor U40538 (N_40538,N_39868,N_39535);
nor U40539 (N_40539,N_39977,N_39737);
xnor U40540 (N_40540,N_39562,N_39617);
xnor U40541 (N_40541,N_39699,N_39766);
nand U40542 (N_40542,N_39052,N_39924);
nand U40543 (N_40543,N_39439,N_39803);
and U40544 (N_40544,N_39999,N_39278);
or U40545 (N_40545,N_39475,N_39168);
or U40546 (N_40546,N_39785,N_39476);
xnor U40547 (N_40547,N_39104,N_39222);
nand U40548 (N_40548,N_39969,N_39229);
and U40549 (N_40549,N_39068,N_39425);
and U40550 (N_40550,N_39088,N_39039);
and U40551 (N_40551,N_39867,N_39893);
and U40552 (N_40552,N_39663,N_39051);
nand U40553 (N_40553,N_39078,N_39568);
nor U40554 (N_40554,N_39858,N_39968);
or U40555 (N_40555,N_39614,N_39959);
nor U40556 (N_40556,N_39444,N_39585);
nand U40557 (N_40557,N_39279,N_39697);
and U40558 (N_40558,N_39697,N_39046);
and U40559 (N_40559,N_39574,N_39541);
xnor U40560 (N_40560,N_39079,N_39159);
or U40561 (N_40561,N_39503,N_39228);
nor U40562 (N_40562,N_39315,N_39084);
nor U40563 (N_40563,N_39844,N_39967);
xnor U40564 (N_40564,N_39406,N_39348);
nor U40565 (N_40565,N_39449,N_39234);
nand U40566 (N_40566,N_39583,N_39972);
and U40567 (N_40567,N_39553,N_39410);
and U40568 (N_40568,N_39784,N_39856);
and U40569 (N_40569,N_39091,N_39601);
nor U40570 (N_40570,N_39550,N_39547);
xor U40571 (N_40571,N_39186,N_39418);
or U40572 (N_40572,N_39063,N_39825);
nor U40573 (N_40573,N_39127,N_39774);
or U40574 (N_40574,N_39823,N_39427);
or U40575 (N_40575,N_39246,N_39244);
or U40576 (N_40576,N_39839,N_39913);
nor U40577 (N_40577,N_39983,N_39717);
or U40578 (N_40578,N_39283,N_39569);
nor U40579 (N_40579,N_39013,N_39304);
or U40580 (N_40580,N_39037,N_39011);
and U40581 (N_40581,N_39814,N_39505);
or U40582 (N_40582,N_39966,N_39803);
nor U40583 (N_40583,N_39377,N_39678);
nand U40584 (N_40584,N_39538,N_39505);
nand U40585 (N_40585,N_39228,N_39686);
nand U40586 (N_40586,N_39989,N_39780);
nand U40587 (N_40587,N_39593,N_39387);
nand U40588 (N_40588,N_39315,N_39757);
xnor U40589 (N_40589,N_39069,N_39959);
and U40590 (N_40590,N_39631,N_39008);
nand U40591 (N_40591,N_39757,N_39393);
nand U40592 (N_40592,N_39775,N_39729);
nor U40593 (N_40593,N_39450,N_39980);
or U40594 (N_40594,N_39226,N_39673);
or U40595 (N_40595,N_39364,N_39616);
or U40596 (N_40596,N_39039,N_39236);
xor U40597 (N_40597,N_39324,N_39188);
or U40598 (N_40598,N_39492,N_39442);
or U40599 (N_40599,N_39270,N_39150);
or U40600 (N_40600,N_39571,N_39002);
xnor U40601 (N_40601,N_39712,N_39259);
xor U40602 (N_40602,N_39124,N_39467);
xnor U40603 (N_40603,N_39639,N_39893);
and U40604 (N_40604,N_39692,N_39099);
nor U40605 (N_40605,N_39318,N_39283);
nand U40606 (N_40606,N_39773,N_39427);
xnor U40607 (N_40607,N_39251,N_39311);
xnor U40608 (N_40608,N_39189,N_39423);
xnor U40609 (N_40609,N_39792,N_39335);
nand U40610 (N_40610,N_39398,N_39286);
nand U40611 (N_40611,N_39832,N_39773);
and U40612 (N_40612,N_39361,N_39558);
or U40613 (N_40613,N_39170,N_39027);
and U40614 (N_40614,N_39425,N_39441);
and U40615 (N_40615,N_39893,N_39825);
or U40616 (N_40616,N_39433,N_39031);
or U40617 (N_40617,N_39038,N_39753);
or U40618 (N_40618,N_39072,N_39149);
or U40619 (N_40619,N_39181,N_39903);
and U40620 (N_40620,N_39834,N_39903);
xnor U40621 (N_40621,N_39787,N_39186);
nand U40622 (N_40622,N_39696,N_39660);
nand U40623 (N_40623,N_39992,N_39936);
nor U40624 (N_40624,N_39150,N_39537);
and U40625 (N_40625,N_39309,N_39097);
and U40626 (N_40626,N_39967,N_39786);
xnor U40627 (N_40627,N_39624,N_39114);
nand U40628 (N_40628,N_39503,N_39268);
nand U40629 (N_40629,N_39435,N_39483);
and U40630 (N_40630,N_39986,N_39677);
or U40631 (N_40631,N_39679,N_39499);
or U40632 (N_40632,N_39986,N_39813);
or U40633 (N_40633,N_39613,N_39778);
or U40634 (N_40634,N_39289,N_39873);
nor U40635 (N_40635,N_39349,N_39020);
and U40636 (N_40636,N_39784,N_39459);
nor U40637 (N_40637,N_39099,N_39608);
nand U40638 (N_40638,N_39307,N_39606);
nor U40639 (N_40639,N_39605,N_39651);
nor U40640 (N_40640,N_39587,N_39815);
and U40641 (N_40641,N_39307,N_39074);
and U40642 (N_40642,N_39436,N_39684);
or U40643 (N_40643,N_39659,N_39887);
nor U40644 (N_40644,N_39221,N_39163);
or U40645 (N_40645,N_39603,N_39519);
or U40646 (N_40646,N_39785,N_39823);
nor U40647 (N_40647,N_39744,N_39814);
nand U40648 (N_40648,N_39448,N_39536);
and U40649 (N_40649,N_39528,N_39574);
nand U40650 (N_40650,N_39851,N_39621);
and U40651 (N_40651,N_39519,N_39023);
or U40652 (N_40652,N_39780,N_39912);
and U40653 (N_40653,N_39428,N_39440);
nand U40654 (N_40654,N_39795,N_39979);
xor U40655 (N_40655,N_39034,N_39391);
or U40656 (N_40656,N_39919,N_39981);
or U40657 (N_40657,N_39740,N_39483);
nor U40658 (N_40658,N_39720,N_39508);
and U40659 (N_40659,N_39504,N_39017);
and U40660 (N_40660,N_39129,N_39872);
nand U40661 (N_40661,N_39235,N_39514);
xor U40662 (N_40662,N_39130,N_39642);
nand U40663 (N_40663,N_39655,N_39027);
or U40664 (N_40664,N_39217,N_39160);
nor U40665 (N_40665,N_39504,N_39183);
nand U40666 (N_40666,N_39812,N_39819);
nor U40667 (N_40667,N_39122,N_39097);
xor U40668 (N_40668,N_39105,N_39263);
or U40669 (N_40669,N_39370,N_39022);
xnor U40670 (N_40670,N_39273,N_39951);
and U40671 (N_40671,N_39350,N_39550);
nor U40672 (N_40672,N_39232,N_39319);
and U40673 (N_40673,N_39461,N_39559);
or U40674 (N_40674,N_39215,N_39327);
nand U40675 (N_40675,N_39069,N_39435);
and U40676 (N_40676,N_39719,N_39324);
or U40677 (N_40677,N_39846,N_39315);
or U40678 (N_40678,N_39945,N_39738);
xor U40679 (N_40679,N_39919,N_39285);
nand U40680 (N_40680,N_39537,N_39867);
and U40681 (N_40681,N_39575,N_39601);
or U40682 (N_40682,N_39807,N_39470);
nand U40683 (N_40683,N_39512,N_39385);
nand U40684 (N_40684,N_39782,N_39144);
nand U40685 (N_40685,N_39433,N_39706);
xnor U40686 (N_40686,N_39410,N_39785);
or U40687 (N_40687,N_39562,N_39499);
xor U40688 (N_40688,N_39527,N_39338);
and U40689 (N_40689,N_39125,N_39978);
or U40690 (N_40690,N_39675,N_39016);
and U40691 (N_40691,N_39031,N_39158);
nand U40692 (N_40692,N_39726,N_39919);
and U40693 (N_40693,N_39811,N_39199);
nand U40694 (N_40694,N_39643,N_39667);
nor U40695 (N_40695,N_39734,N_39255);
xor U40696 (N_40696,N_39789,N_39056);
xor U40697 (N_40697,N_39360,N_39236);
xnor U40698 (N_40698,N_39748,N_39978);
nand U40699 (N_40699,N_39619,N_39532);
or U40700 (N_40700,N_39995,N_39634);
or U40701 (N_40701,N_39770,N_39727);
or U40702 (N_40702,N_39380,N_39034);
or U40703 (N_40703,N_39846,N_39429);
xnor U40704 (N_40704,N_39251,N_39176);
nand U40705 (N_40705,N_39531,N_39667);
and U40706 (N_40706,N_39862,N_39656);
and U40707 (N_40707,N_39939,N_39196);
nand U40708 (N_40708,N_39758,N_39967);
nor U40709 (N_40709,N_39370,N_39946);
nand U40710 (N_40710,N_39316,N_39654);
or U40711 (N_40711,N_39822,N_39175);
or U40712 (N_40712,N_39792,N_39646);
nand U40713 (N_40713,N_39024,N_39371);
or U40714 (N_40714,N_39164,N_39232);
nand U40715 (N_40715,N_39869,N_39204);
or U40716 (N_40716,N_39929,N_39090);
or U40717 (N_40717,N_39908,N_39257);
nand U40718 (N_40718,N_39860,N_39112);
nor U40719 (N_40719,N_39506,N_39158);
nor U40720 (N_40720,N_39004,N_39951);
or U40721 (N_40721,N_39453,N_39235);
or U40722 (N_40722,N_39930,N_39306);
xnor U40723 (N_40723,N_39360,N_39910);
xor U40724 (N_40724,N_39617,N_39055);
and U40725 (N_40725,N_39716,N_39173);
nand U40726 (N_40726,N_39020,N_39944);
nor U40727 (N_40727,N_39912,N_39462);
nor U40728 (N_40728,N_39547,N_39255);
and U40729 (N_40729,N_39122,N_39576);
and U40730 (N_40730,N_39981,N_39762);
nor U40731 (N_40731,N_39723,N_39886);
nor U40732 (N_40732,N_39879,N_39957);
or U40733 (N_40733,N_39510,N_39742);
nor U40734 (N_40734,N_39063,N_39191);
and U40735 (N_40735,N_39788,N_39837);
nand U40736 (N_40736,N_39793,N_39459);
xnor U40737 (N_40737,N_39711,N_39233);
nand U40738 (N_40738,N_39875,N_39485);
nand U40739 (N_40739,N_39876,N_39291);
nand U40740 (N_40740,N_39799,N_39741);
and U40741 (N_40741,N_39923,N_39127);
nor U40742 (N_40742,N_39764,N_39950);
nor U40743 (N_40743,N_39938,N_39595);
and U40744 (N_40744,N_39845,N_39322);
or U40745 (N_40745,N_39616,N_39435);
xor U40746 (N_40746,N_39713,N_39535);
nor U40747 (N_40747,N_39554,N_39127);
nor U40748 (N_40748,N_39351,N_39368);
xnor U40749 (N_40749,N_39217,N_39775);
xnor U40750 (N_40750,N_39633,N_39271);
nor U40751 (N_40751,N_39192,N_39336);
nor U40752 (N_40752,N_39270,N_39367);
xor U40753 (N_40753,N_39050,N_39578);
nand U40754 (N_40754,N_39188,N_39410);
and U40755 (N_40755,N_39688,N_39753);
xnor U40756 (N_40756,N_39510,N_39136);
xor U40757 (N_40757,N_39267,N_39378);
nand U40758 (N_40758,N_39900,N_39768);
and U40759 (N_40759,N_39613,N_39342);
and U40760 (N_40760,N_39968,N_39674);
nand U40761 (N_40761,N_39256,N_39967);
and U40762 (N_40762,N_39919,N_39667);
xnor U40763 (N_40763,N_39448,N_39172);
nor U40764 (N_40764,N_39332,N_39172);
xor U40765 (N_40765,N_39647,N_39755);
nand U40766 (N_40766,N_39048,N_39163);
nand U40767 (N_40767,N_39398,N_39675);
nand U40768 (N_40768,N_39798,N_39588);
and U40769 (N_40769,N_39278,N_39127);
nor U40770 (N_40770,N_39443,N_39060);
xnor U40771 (N_40771,N_39200,N_39998);
nand U40772 (N_40772,N_39346,N_39563);
nor U40773 (N_40773,N_39536,N_39565);
or U40774 (N_40774,N_39925,N_39222);
xor U40775 (N_40775,N_39257,N_39813);
nand U40776 (N_40776,N_39235,N_39162);
nand U40777 (N_40777,N_39485,N_39364);
nand U40778 (N_40778,N_39918,N_39675);
or U40779 (N_40779,N_39703,N_39856);
or U40780 (N_40780,N_39306,N_39245);
nor U40781 (N_40781,N_39500,N_39473);
nor U40782 (N_40782,N_39169,N_39655);
nand U40783 (N_40783,N_39611,N_39959);
and U40784 (N_40784,N_39391,N_39963);
xnor U40785 (N_40785,N_39331,N_39490);
and U40786 (N_40786,N_39621,N_39002);
xnor U40787 (N_40787,N_39134,N_39672);
nor U40788 (N_40788,N_39763,N_39755);
or U40789 (N_40789,N_39635,N_39676);
or U40790 (N_40790,N_39087,N_39566);
or U40791 (N_40791,N_39393,N_39288);
nor U40792 (N_40792,N_39274,N_39751);
xor U40793 (N_40793,N_39037,N_39604);
xor U40794 (N_40794,N_39482,N_39481);
or U40795 (N_40795,N_39403,N_39661);
nand U40796 (N_40796,N_39109,N_39396);
nor U40797 (N_40797,N_39078,N_39650);
and U40798 (N_40798,N_39564,N_39922);
nand U40799 (N_40799,N_39327,N_39242);
and U40800 (N_40800,N_39073,N_39915);
xnor U40801 (N_40801,N_39512,N_39972);
nand U40802 (N_40802,N_39124,N_39877);
and U40803 (N_40803,N_39726,N_39693);
or U40804 (N_40804,N_39472,N_39000);
nand U40805 (N_40805,N_39092,N_39891);
xnor U40806 (N_40806,N_39459,N_39539);
and U40807 (N_40807,N_39529,N_39488);
xnor U40808 (N_40808,N_39171,N_39476);
xor U40809 (N_40809,N_39509,N_39980);
nand U40810 (N_40810,N_39032,N_39726);
nand U40811 (N_40811,N_39319,N_39191);
nand U40812 (N_40812,N_39694,N_39619);
nor U40813 (N_40813,N_39934,N_39894);
xor U40814 (N_40814,N_39775,N_39099);
xnor U40815 (N_40815,N_39814,N_39056);
nor U40816 (N_40816,N_39461,N_39733);
nand U40817 (N_40817,N_39923,N_39216);
nor U40818 (N_40818,N_39476,N_39707);
and U40819 (N_40819,N_39878,N_39699);
and U40820 (N_40820,N_39091,N_39398);
nor U40821 (N_40821,N_39799,N_39041);
nor U40822 (N_40822,N_39349,N_39464);
nand U40823 (N_40823,N_39275,N_39777);
and U40824 (N_40824,N_39992,N_39596);
nor U40825 (N_40825,N_39121,N_39867);
xor U40826 (N_40826,N_39277,N_39293);
or U40827 (N_40827,N_39744,N_39815);
nand U40828 (N_40828,N_39735,N_39474);
nor U40829 (N_40829,N_39134,N_39115);
xor U40830 (N_40830,N_39355,N_39555);
nor U40831 (N_40831,N_39632,N_39925);
nand U40832 (N_40832,N_39826,N_39933);
and U40833 (N_40833,N_39734,N_39726);
nor U40834 (N_40834,N_39814,N_39103);
xor U40835 (N_40835,N_39039,N_39304);
and U40836 (N_40836,N_39901,N_39363);
or U40837 (N_40837,N_39445,N_39168);
or U40838 (N_40838,N_39080,N_39477);
or U40839 (N_40839,N_39881,N_39925);
nor U40840 (N_40840,N_39650,N_39202);
xnor U40841 (N_40841,N_39411,N_39883);
nor U40842 (N_40842,N_39767,N_39244);
or U40843 (N_40843,N_39678,N_39512);
and U40844 (N_40844,N_39202,N_39234);
nor U40845 (N_40845,N_39218,N_39496);
or U40846 (N_40846,N_39482,N_39730);
nand U40847 (N_40847,N_39162,N_39330);
or U40848 (N_40848,N_39740,N_39844);
and U40849 (N_40849,N_39481,N_39828);
nand U40850 (N_40850,N_39344,N_39628);
and U40851 (N_40851,N_39062,N_39763);
xnor U40852 (N_40852,N_39786,N_39207);
xnor U40853 (N_40853,N_39056,N_39201);
xnor U40854 (N_40854,N_39318,N_39296);
nor U40855 (N_40855,N_39878,N_39419);
xnor U40856 (N_40856,N_39314,N_39186);
xnor U40857 (N_40857,N_39546,N_39355);
and U40858 (N_40858,N_39350,N_39242);
xor U40859 (N_40859,N_39665,N_39118);
xnor U40860 (N_40860,N_39425,N_39906);
or U40861 (N_40861,N_39667,N_39634);
nand U40862 (N_40862,N_39233,N_39167);
nand U40863 (N_40863,N_39759,N_39305);
and U40864 (N_40864,N_39406,N_39474);
or U40865 (N_40865,N_39144,N_39340);
nor U40866 (N_40866,N_39320,N_39383);
xnor U40867 (N_40867,N_39052,N_39948);
xnor U40868 (N_40868,N_39565,N_39490);
or U40869 (N_40869,N_39261,N_39053);
or U40870 (N_40870,N_39687,N_39998);
xor U40871 (N_40871,N_39971,N_39152);
nor U40872 (N_40872,N_39201,N_39217);
or U40873 (N_40873,N_39991,N_39813);
and U40874 (N_40874,N_39335,N_39759);
nor U40875 (N_40875,N_39643,N_39007);
and U40876 (N_40876,N_39014,N_39728);
nor U40877 (N_40877,N_39327,N_39216);
and U40878 (N_40878,N_39304,N_39913);
nor U40879 (N_40879,N_39564,N_39635);
and U40880 (N_40880,N_39758,N_39817);
xor U40881 (N_40881,N_39667,N_39094);
xor U40882 (N_40882,N_39516,N_39002);
xnor U40883 (N_40883,N_39176,N_39719);
xor U40884 (N_40884,N_39817,N_39421);
nand U40885 (N_40885,N_39351,N_39778);
or U40886 (N_40886,N_39983,N_39578);
and U40887 (N_40887,N_39504,N_39724);
xor U40888 (N_40888,N_39517,N_39213);
and U40889 (N_40889,N_39503,N_39303);
or U40890 (N_40890,N_39114,N_39653);
or U40891 (N_40891,N_39002,N_39694);
or U40892 (N_40892,N_39499,N_39608);
and U40893 (N_40893,N_39180,N_39539);
nand U40894 (N_40894,N_39156,N_39688);
nor U40895 (N_40895,N_39812,N_39598);
xor U40896 (N_40896,N_39168,N_39925);
nand U40897 (N_40897,N_39943,N_39299);
nor U40898 (N_40898,N_39848,N_39991);
or U40899 (N_40899,N_39768,N_39336);
and U40900 (N_40900,N_39861,N_39506);
nor U40901 (N_40901,N_39107,N_39934);
and U40902 (N_40902,N_39040,N_39902);
xor U40903 (N_40903,N_39782,N_39902);
and U40904 (N_40904,N_39020,N_39035);
or U40905 (N_40905,N_39044,N_39431);
nor U40906 (N_40906,N_39958,N_39624);
xnor U40907 (N_40907,N_39468,N_39176);
nand U40908 (N_40908,N_39454,N_39489);
or U40909 (N_40909,N_39411,N_39348);
nor U40910 (N_40910,N_39365,N_39583);
and U40911 (N_40911,N_39217,N_39648);
nand U40912 (N_40912,N_39070,N_39688);
xor U40913 (N_40913,N_39644,N_39082);
and U40914 (N_40914,N_39963,N_39947);
nand U40915 (N_40915,N_39992,N_39115);
or U40916 (N_40916,N_39319,N_39070);
and U40917 (N_40917,N_39602,N_39929);
and U40918 (N_40918,N_39003,N_39325);
xnor U40919 (N_40919,N_39217,N_39066);
and U40920 (N_40920,N_39129,N_39380);
nor U40921 (N_40921,N_39824,N_39485);
nand U40922 (N_40922,N_39051,N_39325);
nor U40923 (N_40923,N_39101,N_39447);
and U40924 (N_40924,N_39675,N_39593);
nor U40925 (N_40925,N_39534,N_39493);
nand U40926 (N_40926,N_39590,N_39875);
and U40927 (N_40927,N_39295,N_39805);
nor U40928 (N_40928,N_39413,N_39013);
or U40929 (N_40929,N_39400,N_39243);
xor U40930 (N_40930,N_39070,N_39266);
xor U40931 (N_40931,N_39473,N_39652);
nand U40932 (N_40932,N_39147,N_39001);
nor U40933 (N_40933,N_39368,N_39370);
and U40934 (N_40934,N_39430,N_39655);
and U40935 (N_40935,N_39612,N_39336);
and U40936 (N_40936,N_39179,N_39706);
xor U40937 (N_40937,N_39487,N_39067);
nand U40938 (N_40938,N_39231,N_39462);
nor U40939 (N_40939,N_39943,N_39318);
nand U40940 (N_40940,N_39394,N_39431);
or U40941 (N_40941,N_39101,N_39732);
nor U40942 (N_40942,N_39523,N_39864);
or U40943 (N_40943,N_39990,N_39462);
xnor U40944 (N_40944,N_39223,N_39493);
xor U40945 (N_40945,N_39234,N_39892);
or U40946 (N_40946,N_39227,N_39621);
xnor U40947 (N_40947,N_39695,N_39254);
and U40948 (N_40948,N_39053,N_39907);
nand U40949 (N_40949,N_39583,N_39641);
xor U40950 (N_40950,N_39546,N_39207);
or U40951 (N_40951,N_39699,N_39323);
nand U40952 (N_40952,N_39295,N_39321);
and U40953 (N_40953,N_39985,N_39271);
and U40954 (N_40954,N_39386,N_39371);
and U40955 (N_40955,N_39789,N_39073);
xnor U40956 (N_40956,N_39571,N_39707);
xor U40957 (N_40957,N_39140,N_39528);
nor U40958 (N_40958,N_39336,N_39993);
or U40959 (N_40959,N_39063,N_39391);
xor U40960 (N_40960,N_39974,N_39726);
xor U40961 (N_40961,N_39081,N_39487);
xor U40962 (N_40962,N_39638,N_39657);
or U40963 (N_40963,N_39112,N_39140);
nand U40964 (N_40964,N_39122,N_39608);
and U40965 (N_40965,N_39295,N_39588);
nand U40966 (N_40966,N_39075,N_39319);
nor U40967 (N_40967,N_39190,N_39167);
or U40968 (N_40968,N_39514,N_39218);
and U40969 (N_40969,N_39547,N_39493);
nor U40970 (N_40970,N_39908,N_39806);
and U40971 (N_40971,N_39142,N_39569);
nand U40972 (N_40972,N_39176,N_39605);
xnor U40973 (N_40973,N_39004,N_39805);
or U40974 (N_40974,N_39906,N_39500);
xnor U40975 (N_40975,N_39039,N_39776);
or U40976 (N_40976,N_39097,N_39438);
nor U40977 (N_40977,N_39835,N_39362);
or U40978 (N_40978,N_39398,N_39698);
or U40979 (N_40979,N_39996,N_39206);
nor U40980 (N_40980,N_39360,N_39998);
nor U40981 (N_40981,N_39746,N_39009);
or U40982 (N_40982,N_39066,N_39482);
nand U40983 (N_40983,N_39413,N_39410);
or U40984 (N_40984,N_39620,N_39226);
nand U40985 (N_40985,N_39335,N_39502);
xnor U40986 (N_40986,N_39684,N_39654);
and U40987 (N_40987,N_39946,N_39419);
and U40988 (N_40988,N_39743,N_39263);
and U40989 (N_40989,N_39184,N_39818);
xnor U40990 (N_40990,N_39157,N_39545);
nor U40991 (N_40991,N_39532,N_39382);
and U40992 (N_40992,N_39635,N_39190);
nor U40993 (N_40993,N_39633,N_39274);
nor U40994 (N_40994,N_39029,N_39569);
nand U40995 (N_40995,N_39518,N_39905);
nor U40996 (N_40996,N_39170,N_39745);
or U40997 (N_40997,N_39944,N_39683);
xnor U40998 (N_40998,N_39806,N_39168);
xnor U40999 (N_40999,N_39927,N_39048);
nor U41000 (N_41000,N_40467,N_40508);
nand U41001 (N_41001,N_40484,N_40059);
nor U41002 (N_41002,N_40157,N_40928);
and U41003 (N_41003,N_40586,N_40333);
nand U41004 (N_41004,N_40271,N_40347);
xnor U41005 (N_41005,N_40133,N_40732);
xor U41006 (N_41006,N_40552,N_40772);
nor U41007 (N_41007,N_40022,N_40023);
and U41008 (N_41008,N_40219,N_40120);
xor U41009 (N_41009,N_40436,N_40388);
nor U41010 (N_41010,N_40101,N_40797);
nor U41011 (N_41011,N_40870,N_40202);
nand U41012 (N_41012,N_40128,N_40233);
or U41013 (N_41013,N_40414,N_40683);
nor U41014 (N_41014,N_40661,N_40764);
xor U41015 (N_41015,N_40415,N_40925);
or U41016 (N_41016,N_40030,N_40911);
xnor U41017 (N_41017,N_40882,N_40153);
xnor U41018 (N_41018,N_40151,N_40813);
and U41019 (N_41019,N_40042,N_40439);
nor U41020 (N_41020,N_40770,N_40221);
or U41021 (N_41021,N_40284,N_40631);
nor U41022 (N_41022,N_40741,N_40418);
nand U41023 (N_41023,N_40431,N_40684);
nor U41024 (N_41024,N_40368,N_40419);
xor U41025 (N_41025,N_40601,N_40465);
nor U41026 (N_41026,N_40659,N_40315);
or U41027 (N_41027,N_40780,N_40759);
nor U41028 (N_41028,N_40097,N_40213);
nand U41029 (N_41029,N_40862,N_40432);
or U41030 (N_41030,N_40913,N_40855);
or U41031 (N_41031,N_40671,N_40196);
nor U41032 (N_41032,N_40406,N_40424);
nand U41033 (N_41033,N_40905,N_40959);
xnor U41034 (N_41034,N_40075,N_40280);
nand U41035 (N_41035,N_40978,N_40255);
and U41036 (N_41036,N_40635,N_40955);
nand U41037 (N_41037,N_40539,N_40585);
and U41038 (N_41038,N_40794,N_40125);
xor U41039 (N_41039,N_40223,N_40081);
or U41040 (N_41040,N_40938,N_40037);
nand U41041 (N_41041,N_40853,N_40496);
and U41042 (N_41042,N_40940,N_40718);
and U41043 (N_41043,N_40294,N_40766);
xor U41044 (N_41044,N_40869,N_40685);
and U41045 (N_41045,N_40815,N_40933);
nand U41046 (N_41046,N_40458,N_40632);
or U41047 (N_41047,N_40274,N_40131);
nor U41048 (N_41048,N_40584,N_40437);
xor U41049 (N_41049,N_40946,N_40111);
or U41050 (N_41050,N_40245,N_40006);
and U41051 (N_41051,N_40642,N_40653);
nand U41052 (N_41052,N_40500,N_40445);
nor U41053 (N_41053,N_40316,N_40681);
or U41054 (N_41054,N_40690,N_40839);
or U41055 (N_41055,N_40654,N_40040);
and U41056 (N_41056,N_40660,N_40567);
nor U41057 (N_41057,N_40198,N_40719);
xor U41058 (N_41058,N_40450,N_40178);
and U41059 (N_41059,N_40738,N_40616);
nor U41060 (N_41060,N_40045,N_40725);
nor U41061 (N_41061,N_40537,N_40995);
nand U41062 (N_41062,N_40655,N_40737);
nor U41063 (N_41063,N_40008,N_40234);
xnor U41064 (N_41064,N_40474,N_40723);
xor U41065 (N_41065,N_40173,N_40997);
xor U41066 (N_41066,N_40808,N_40645);
or U41067 (N_41067,N_40957,N_40872);
and U41068 (N_41068,N_40582,N_40866);
and U41069 (N_41069,N_40481,N_40201);
nor U41070 (N_41070,N_40954,N_40695);
nor U41071 (N_41071,N_40972,N_40887);
xnor U41072 (N_41072,N_40319,N_40354);
or U41073 (N_41073,N_40346,N_40307);
nand U41074 (N_41074,N_40158,N_40374);
and U41075 (N_41075,N_40921,N_40848);
nor U41076 (N_41076,N_40636,N_40868);
and U41077 (N_41077,N_40998,N_40569);
nand U41078 (N_41078,N_40247,N_40657);
nor U41079 (N_41079,N_40630,N_40523);
nor U41080 (N_41080,N_40041,N_40625);
and U41081 (N_41081,N_40289,N_40126);
or U41082 (N_41082,N_40005,N_40892);
xor U41083 (N_41083,N_40429,N_40485);
or U41084 (N_41084,N_40580,N_40417);
nand U41085 (N_41085,N_40146,N_40413);
and U41086 (N_41086,N_40825,N_40947);
or U41087 (N_41087,N_40299,N_40345);
and U41088 (N_41088,N_40204,N_40934);
xnor U41089 (N_41089,N_40114,N_40190);
nor U41090 (N_41090,N_40034,N_40177);
nor U41091 (N_41091,N_40894,N_40889);
or U41092 (N_41092,N_40533,N_40590);
xor U41093 (N_41093,N_40740,N_40364);
and U41094 (N_41094,N_40142,N_40138);
or U41095 (N_41095,N_40704,N_40506);
nor U41096 (N_41096,N_40207,N_40819);
xor U41097 (N_41097,N_40407,N_40149);
nor U41098 (N_41098,N_40952,N_40669);
nor U41099 (N_41099,N_40052,N_40646);
nor U41100 (N_41100,N_40795,N_40408);
or U41101 (N_41101,N_40127,N_40501);
and U41102 (N_41102,N_40534,N_40489);
nor U41103 (N_41103,N_40517,N_40471);
xnor U41104 (N_41104,N_40265,N_40001);
and U41105 (N_41105,N_40675,N_40656);
nand U41106 (N_41106,N_40773,N_40224);
xor U41107 (N_41107,N_40516,N_40726);
nor U41108 (N_41108,N_40067,N_40141);
and U41109 (N_41109,N_40077,N_40867);
or U41110 (N_41110,N_40055,N_40000);
xor U41111 (N_41111,N_40864,N_40236);
nand U41112 (N_41112,N_40438,N_40139);
nand U41113 (N_41113,N_40960,N_40464);
or U41114 (N_41114,N_40554,N_40261);
xnor U41115 (N_41115,N_40162,N_40382);
nand U41116 (N_41116,N_40781,N_40387);
nand U41117 (N_41117,N_40812,N_40348);
nand U41118 (N_41118,N_40383,N_40011);
nand U41119 (N_41119,N_40589,N_40020);
nor U41120 (N_41120,N_40604,N_40666);
xnor U41121 (N_41121,N_40943,N_40673);
xnor U41122 (N_41122,N_40254,N_40576);
or U41123 (N_41123,N_40999,N_40462);
and U41124 (N_41124,N_40287,N_40412);
nor U41125 (N_41125,N_40950,N_40817);
nand U41126 (N_41126,N_40252,N_40748);
and U41127 (N_41127,N_40229,N_40927);
nand U41128 (N_41128,N_40956,N_40248);
xor U41129 (N_41129,N_40594,N_40273);
nand U41130 (N_41130,N_40851,N_40235);
nor U41131 (N_41131,N_40013,N_40066);
nand U41132 (N_41132,N_40355,N_40935);
or U41133 (N_41133,N_40608,N_40974);
xnor U41134 (N_41134,N_40434,N_40473);
xnor U41135 (N_41135,N_40860,N_40854);
and U41136 (N_41136,N_40401,N_40623);
nor U41137 (N_41137,N_40391,N_40033);
xnor U41138 (N_41138,N_40511,N_40026);
nand U41139 (N_41139,N_40472,N_40237);
nor U41140 (N_41140,N_40342,N_40155);
xnor U41141 (N_41141,N_40370,N_40038);
nand U41142 (N_41142,N_40863,N_40277);
nor U41143 (N_41143,N_40615,N_40563);
nor U41144 (N_41144,N_40735,N_40832);
nor U41145 (N_41145,N_40961,N_40626);
xor U41146 (N_41146,N_40593,N_40612);
or U41147 (N_41147,N_40542,N_40605);
or U41148 (N_41148,N_40416,N_40880);
and U41149 (N_41149,N_40015,N_40981);
nor U41150 (N_41150,N_40587,N_40885);
xnor U41151 (N_41151,N_40099,N_40330);
or U41152 (N_41152,N_40478,N_40686);
xor U41153 (N_41153,N_40620,N_40044);
nor U41154 (N_41154,N_40375,N_40682);
xor U41155 (N_41155,N_40268,N_40639);
nand U41156 (N_41156,N_40694,N_40072);
nor U41157 (N_41157,N_40744,N_40509);
or U41158 (N_41158,N_40352,N_40025);
or U41159 (N_41159,N_40640,N_40137);
nand U41160 (N_41160,N_40842,N_40877);
nand U41161 (N_41161,N_40336,N_40806);
nand U41162 (N_41162,N_40761,N_40123);
or U41163 (N_41163,N_40278,N_40185);
nand U41164 (N_41164,N_40166,N_40087);
nor U41165 (N_41165,N_40226,N_40937);
and U41166 (N_41166,N_40134,N_40633);
xnor U41167 (N_41167,N_40621,N_40822);
nor U41168 (N_41168,N_40180,N_40917);
nand U41169 (N_41169,N_40003,N_40012);
or U41170 (N_41170,N_40065,N_40930);
nand U41171 (N_41171,N_40189,N_40688);
nor U41172 (N_41172,N_40801,N_40831);
or U41173 (N_41173,N_40859,N_40024);
nor U41174 (N_41174,N_40269,N_40969);
or U41175 (N_41175,N_40308,N_40420);
and U41176 (N_41176,N_40811,N_40263);
and U41177 (N_41177,N_40386,N_40175);
nand U41178 (N_41178,N_40170,N_40774);
nand U41179 (N_41179,N_40596,N_40792);
or U41180 (N_41180,N_40964,N_40507);
xnor U41181 (N_41181,N_40919,N_40241);
xnor U41182 (N_41182,N_40266,N_40729);
and U41183 (N_41183,N_40222,N_40035);
or U41184 (N_41184,N_40080,N_40893);
xor U41185 (N_41185,N_40897,N_40966);
xor U41186 (N_41186,N_40152,N_40427);
nand U41187 (N_41187,N_40062,N_40169);
or U41188 (N_41188,N_40830,N_40376);
nor U41189 (N_41189,N_40514,N_40791);
nand U41190 (N_41190,N_40109,N_40494);
or U41191 (N_41191,N_40670,N_40147);
xnor U41192 (N_41192,N_40083,N_40130);
nand U41193 (N_41193,N_40503,N_40550);
or U41194 (N_41194,N_40122,N_40548);
nand U41195 (N_41195,N_40292,N_40852);
and U41196 (N_41196,N_40692,N_40334);
xnor U41197 (N_41197,N_40426,N_40807);
xnor U41198 (N_41198,N_40054,N_40578);
nor U41199 (N_41199,N_40398,N_40297);
or U41200 (N_41200,N_40982,N_40619);
and U41201 (N_41201,N_40228,N_40209);
nand U41202 (N_41202,N_40039,N_40384);
and U41203 (N_41203,N_40144,N_40086);
nand U41204 (N_41204,N_40161,N_40136);
nor U41205 (N_41205,N_40350,N_40168);
nor U41206 (N_41206,N_40486,N_40225);
xnor U41207 (N_41207,N_40665,N_40283);
and U41208 (N_41208,N_40971,N_40325);
nand U41209 (N_41209,N_40423,N_40805);
or U41210 (N_41210,N_40409,N_40676);
nand U41211 (N_41211,N_40159,N_40218);
nand U41212 (N_41212,N_40984,N_40778);
nand U41213 (N_41213,N_40487,N_40073);
or U41214 (N_41214,N_40727,N_40390);
nor U41215 (N_41215,N_40480,N_40891);
xor U41216 (N_41216,N_40979,N_40344);
or U41217 (N_41217,N_40541,N_40743);
nor U41218 (N_41218,N_40896,N_40793);
and U41219 (N_41219,N_40712,N_40321);
or U41220 (N_41220,N_40389,N_40574);
xnor U41221 (N_41221,N_40611,N_40078);
or U41222 (N_41222,N_40910,N_40318);
xnor U41223 (N_41223,N_40016,N_40754);
nor U41224 (N_41224,N_40353,N_40181);
nand U41225 (N_41225,N_40703,N_40405);
and U41226 (N_41226,N_40524,N_40296);
nor U41227 (N_41227,N_40205,N_40543);
nor U41228 (N_41228,N_40483,N_40179);
xor U41229 (N_41229,N_40105,N_40710);
xor U41230 (N_41230,N_40525,N_40371);
xor U41231 (N_41231,N_40488,N_40309);
nand U41232 (N_41232,N_40396,N_40460);
xnor U41233 (N_41233,N_40555,N_40798);
and U41234 (N_41234,N_40809,N_40706);
and U41235 (N_41235,N_40053,N_40929);
xor U41236 (N_41236,N_40156,N_40785);
and U41237 (N_41237,N_40206,N_40886);
and U41238 (N_41238,N_40124,N_40977);
xor U41239 (N_41239,N_40617,N_40068);
nand U41240 (N_41240,N_40728,N_40988);
nor U41241 (N_41241,N_40923,N_40824);
and U41242 (N_41242,N_40753,N_40449);
or U41243 (N_41243,N_40777,N_40239);
xnor U41244 (N_41244,N_40702,N_40377);
or U41245 (N_41245,N_40084,N_40932);
xnor U41246 (N_41246,N_40027,N_40820);
xor U41247 (N_41247,N_40678,N_40441);
nand U41248 (N_41248,N_40823,N_40519);
or U41249 (N_41249,N_40644,N_40597);
xnor U41250 (N_41250,N_40323,N_40463);
and U41251 (N_41251,N_40402,N_40936);
xnor U41252 (N_41252,N_40606,N_40610);
and U41253 (N_41253,N_40570,N_40212);
and U41254 (N_41254,N_40902,N_40322);
nand U41255 (N_41255,N_40556,N_40057);
nor U41256 (N_41256,N_40453,N_40652);
nand U41257 (N_41257,N_40253,N_40028);
or U41258 (N_41258,N_40010,N_40337);
and U41259 (N_41259,N_40428,N_40691);
or U41260 (N_41260,N_40967,N_40672);
nor U41261 (N_41261,N_40711,N_40260);
nor U41262 (N_41262,N_40571,N_40931);
nor U41263 (N_41263,N_40833,N_40843);
nor U41264 (N_41264,N_40121,N_40581);
xor U41265 (N_41265,N_40118,N_40722);
and U41266 (N_41266,N_40214,N_40461);
xnor U41267 (N_41267,N_40454,N_40746);
nor U41268 (N_41268,N_40435,N_40536);
xor U41269 (N_41269,N_40721,N_40535);
or U41270 (N_41270,N_40312,N_40951);
or U41271 (N_41271,N_40107,N_40561);
or U41272 (N_41272,N_40883,N_40160);
nand U41273 (N_41273,N_40965,N_40775);
or U41274 (N_41274,N_40021,N_40298);
and U41275 (N_41275,N_40527,N_40477);
and U41276 (N_41276,N_40340,N_40165);
nand U41277 (N_41277,N_40240,N_40306);
nand U41278 (N_41278,N_40091,N_40980);
nor U41279 (N_41279,N_40926,N_40858);
nand U41280 (N_41280,N_40779,N_40904);
or U41281 (N_41281,N_40100,N_40243);
and U41282 (N_41282,N_40267,N_40258);
nand U41283 (N_41283,N_40143,N_40575);
xor U41284 (N_41284,N_40140,N_40835);
and U41285 (N_41285,N_40787,N_40939);
or U41286 (N_41286,N_40985,N_40069);
xor U41287 (N_41287,N_40357,N_40343);
xor U41288 (N_41288,N_40032,N_40171);
xor U41289 (N_41289,N_40989,N_40865);
nor U41290 (N_41290,N_40900,N_40079);
or U41291 (N_41291,N_40758,N_40518);
or U41292 (N_41292,N_40530,N_40092);
and U41293 (N_41293,N_40440,N_40095);
nor U41294 (N_41294,N_40650,N_40279);
and U41295 (N_41295,N_40522,N_40515);
nor U41296 (N_41296,N_40285,N_40215);
or U41297 (N_41297,N_40840,N_40186);
nand U41298 (N_41298,N_40498,N_40958);
nor U41299 (N_41299,N_40948,N_40814);
nand U41300 (N_41300,N_40276,N_40845);
nand U41301 (N_41301,N_40579,N_40510);
or U41302 (N_41302,N_40211,N_40804);
nor U41303 (N_41303,N_40901,N_40145);
or U41304 (N_41304,N_40399,N_40526);
and U41305 (N_41305,N_40549,N_40050);
nand U41306 (N_41306,N_40802,N_40007);
xnor U41307 (N_41307,N_40755,N_40031);
and U41308 (N_41308,N_40907,N_40693);
nor U41309 (N_41309,N_40898,N_40104);
nand U41310 (N_41310,N_40113,N_40873);
nor U41311 (N_41311,N_40455,N_40987);
or U41312 (N_41312,N_40098,N_40970);
nand U41313 (N_41313,N_40349,N_40739);
and U41314 (N_41314,N_40459,N_40912);
or U41315 (N_41315,N_40332,N_40089);
xnor U41316 (N_41316,N_40183,N_40899);
nor U41317 (N_41317,N_40529,N_40360);
and U41318 (N_41318,N_40895,N_40208);
or U41319 (N_41319,N_40668,N_40259);
xnor U41320 (N_41320,N_40816,N_40217);
nand U41321 (N_41321,N_40492,N_40720);
nand U41322 (N_41322,N_40918,N_40700);
nand U41323 (N_41323,N_40456,N_40944);
xor U41324 (N_41324,N_40358,N_40150);
xor U41325 (N_41325,N_40915,N_40641);
xnor U41326 (N_41326,N_40609,N_40962);
and U41327 (N_41327,N_40504,N_40112);
xor U41328 (N_41328,N_40857,N_40093);
nand U41329 (N_41329,N_40874,N_40745);
nor U41330 (N_41330,N_40953,N_40532);
nor U41331 (N_41331,N_40992,N_40275);
xor U41332 (N_41332,N_40789,N_40366);
nor U41333 (N_41333,N_40362,N_40622);
xor U41334 (N_41334,N_40071,N_40572);
or U41335 (N_41335,N_40547,N_40110);
and U41336 (N_41336,N_40838,N_40699);
nor U41337 (N_41337,N_40762,N_40829);
and U41338 (N_41338,N_40782,N_40602);
or U41339 (N_41339,N_40291,N_40600);
nand U41340 (N_41340,N_40116,N_40017);
xnor U41341 (N_41341,N_40861,N_40757);
nand U41342 (N_41342,N_40760,N_40447);
and U41343 (N_41343,N_40577,N_40187);
or U41344 (N_41344,N_40736,N_40174);
nor U41345 (N_41345,N_40771,N_40647);
nand U41346 (N_41346,N_40164,N_40074);
nor U41347 (N_41347,N_40210,N_40430);
and U41348 (N_41348,N_40314,N_40986);
xor U41349 (N_41349,N_40476,N_40879);
and U41350 (N_41350,N_40520,N_40421);
nor U41351 (N_41351,N_40320,N_40090);
nand U41352 (N_41352,N_40176,N_40697);
xnor U41353 (N_41353,N_40397,N_40272);
and U41354 (N_41354,N_40172,N_40624);
nand U41355 (N_41355,N_40191,N_40890);
nor U41356 (N_41356,N_40061,N_40493);
xor U41357 (N_41357,N_40331,N_40784);
and U41358 (N_41358,N_40167,N_40553);
nor U41359 (N_41359,N_40378,N_40076);
nand U41360 (N_41360,N_40649,N_40628);
xor U41361 (N_41361,N_40531,N_40834);
and U41362 (N_41362,N_40803,N_40199);
nand U41363 (N_41363,N_40513,N_40663);
nor U41364 (N_41364,N_40058,N_40991);
nor U41365 (N_41365,N_40192,N_40546);
xnor U41366 (N_41366,N_40871,N_40920);
nor U41367 (N_41367,N_40195,N_40103);
nand U41368 (N_41368,N_40922,N_40651);
nand U41369 (N_41369,N_40115,N_40776);
nand U41370 (N_41370,N_40048,N_40043);
xnor U41371 (N_41371,N_40752,N_40715);
xnor U41372 (N_41372,N_40148,N_40994);
nand U41373 (N_41373,N_40497,N_40102);
nand U41374 (N_41374,N_40790,N_40106);
or U41375 (N_41375,N_40566,N_40341);
or U41376 (N_41376,N_40317,N_40495);
and U41377 (N_41377,N_40004,N_40818);
nand U41378 (N_41378,N_40286,N_40713);
nor U41379 (N_41379,N_40878,N_40182);
or U41380 (N_41380,N_40282,N_40359);
or U41381 (N_41381,N_40230,N_40701);
or U41382 (N_41382,N_40502,N_40750);
or U41383 (N_41383,N_40385,N_40749);
or U41384 (N_41384,N_40696,N_40443);
or U41385 (N_41385,N_40365,N_40714);
nand U41386 (N_41386,N_40788,N_40521);
nor U41387 (N_41387,N_40643,N_40444);
nand U41388 (N_41388,N_40849,N_40457);
and U41389 (N_41389,N_40231,N_40875);
nand U41390 (N_41390,N_40303,N_40876);
or U41391 (N_41391,N_40193,N_40648);
and U41392 (N_41392,N_40490,N_40257);
nand U41393 (N_41393,N_40302,N_40242);
or U41394 (N_41394,N_40422,N_40968);
or U41395 (N_41395,N_40996,N_40361);
and U41396 (N_41396,N_40560,N_40810);
xnor U41397 (N_41397,N_40884,N_40117);
xor U41398 (N_41398,N_40949,N_40724);
xor U41399 (N_41399,N_40403,N_40448);
xor U41400 (N_41400,N_40446,N_40888);
nor U41401 (N_41401,N_40301,N_40433);
and U41402 (N_41402,N_40990,N_40742);
nand U41403 (N_41403,N_40270,N_40599);
nand U41404 (N_41404,N_40705,N_40468);
nand U41405 (N_41405,N_40796,N_40051);
or U41406 (N_41406,N_40154,N_40827);
and U41407 (N_41407,N_40404,N_40380);
nand U41408 (N_41408,N_40310,N_40551);
nor U41409 (N_41409,N_40592,N_40512);
nand U41410 (N_41410,N_40466,N_40942);
or U41411 (N_41411,N_40338,N_40559);
and U41412 (N_41412,N_40800,N_40680);
or U41413 (N_41413,N_40324,N_40295);
or U41414 (N_41414,N_40914,N_40847);
and U41415 (N_41415,N_40367,N_40328);
or U41416 (N_41416,N_40410,N_40329);
nand U41417 (N_41417,N_40941,N_40634);
nor U41418 (N_41418,N_40305,N_40841);
nor U41419 (N_41419,N_40135,N_40046);
and U41420 (N_41420,N_40395,N_40769);
or U41421 (N_41421,N_40019,N_40730);
xor U41422 (N_41422,N_40588,N_40227);
nand U41423 (N_41423,N_40288,N_40372);
nand U41424 (N_41424,N_40197,N_40002);
xnor U41425 (N_41425,N_40558,N_40351);
nor U41426 (N_41426,N_40326,N_40482);
nand U41427 (N_41427,N_40163,N_40846);
xnor U41428 (N_41428,N_40251,N_40184);
or U41429 (N_41429,N_40733,N_40194);
and U41430 (N_41430,N_40369,N_40658);
or U41431 (N_41431,N_40629,N_40356);
xnor U41432 (N_41432,N_40627,N_40573);
xor U41433 (N_41433,N_40264,N_40614);
nor U41434 (N_41434,N_40844,N_40763);
nand U41435 (N_41435,N_40618,N_40014);
nand U41436 (N_41436,N_40828,N_40060);
nor U41437 (N_41437,N_40363,N_40470);
nand U41438 (N_41438,N_40392,N_40491);
and U41439 (N_41439,N_40903,N_40018);
or U41440 (N_41440,N_40064,N_40400);
nand U41441 (N_41441,N_40036,N_40096);
nor U41442 (N_41442,N_40250,N_40707);
xnor U41443 (N_41443,N_40747,N_40505);
or U41444 (N_41444,N_40708,N_40607);
or U41445 (N_41445,N_40544,N_40603);
and U41446 (N_41446,N_40765,N_40881);
nand U41447 (N_41447,N_40916,N_40783);
and U41448 (N_41448,N_40565,N_40232);
xnor U41449 (N_41449,N_40246,N_40598);
nand U41450 (N_41450,N_40411,N_40469);
and U41451 (N_41451,N_40442,N_40698);
nor U41452 (N_41452,N_40734,N_40339);
xor U41453 (N_41453,N_40756,N_40499);
nor U41454 (N_41454,N_40056,N_40088);
nor U41455 (N_41455,N_40394,N_40637);
and U41456 (N_41456,N_40837,N_40029);
nor U41457 (N_41457,N_40595,N_40709);
or U41458 (N_41458,N_40799,N_40821);
and U41459 (N_41459,N_40049,N_40300);
xnor U41460 (N_41460,N_40850,N_40129);
nand U41461 (N_41461,N_40751,N_40613);
nor U41462 (N_41462,N_40188,N_40768);
nand U41463 (N_41463,N_40203,N_40856);
nand U41464 (N_41464,N_40381,N_40674);
xnor U41465 (N_41465,N_40538,N_40216);
and U41466 (N_41466,N_40667,N_40311);
nor U41467 (N_41467,N_40479,N_40557);
and U41468 (N_41468,N_40290,N_40583);
or U41469 (N_41469,N_40976,N_40047);
nor U41470 (N_41470,N_40108,N_40906);
and U41471 (N_41471,N_40716,N_40327);
xor U41472 (N_41472,N_40379,N_40475);
and U41473 (N_41473,N_40085,N_40540);
xnor U41474 (N_41474,N_40528,N_40220);
nand U41475 (N_41475,N_40909,N_40945);
nand U41476 (N_41476,N_40452,N_40983);
nor U41477 (N_41477,N_40238,N_40767);
xnor U41478 (N_41478,N_40664,N_40731);
nand U41479 (N_41479,N_40082,N_40826);
nor U41480 (N_41480,N_40249,N_40119);
or U41481 (N_41481,N_40836,N_40993);
nor U41482 (N_41482,N_40244,N_40963);
xor U41483 (N_41483,N_40313,N_40679);
nor U41484 (N_41484,N_40393,N_40281);
and U41485 (N_41485,N_40335,N_40304);
or U41486 (N_41486,N_40373,N_40568);
nor U41487 (N_41487,N_40070,N_40293);
nor U41488 (N_41488,N_40262,N_40689);
nor U41489 (N_41489,N_40677,N_40662);
nor U41490 (N_41490,N_40451,N_40132);
nand U41491 (N_41491,N_40786,N_40973);
and U41492 (N_41492,N_40564,N_40924);
xnor U41493 (N_41493,N_40562,N_40638);
or U41494 (N_41494,N_40975,N_40425);
nor U41495 (N_41495,N_40908,N_40009);
or U41496 (N_41496,N_40094,N_40256);
and U41497 (N_41497,N_40687,N_40545);
xor U41498 (N_41498,N_40591,N_40717);
and U41499 (N_41499,N_40200,N_40063);
xnor U41500 (N_41500,N_40347,N_40514);
and U41501 (N_41501,N_40618,N_40442);
xor U41502 (N_41502,N_40525,N_40291);
nand U41503 (N_41503,N_40125,N_40243);
or U41504 (N_41504,N_40616,N_40213);
nor U41505 (N_41505,N_40679,N_40723);
nor U41506 (N_41506,N_40625,N_40290);
or U41507 (N_41507,N_40800,N_40047);
or U41508 (N_41508,N_40692,N_40021);
or U41509 (N_41509,N_40227,N_40918);
xnor U41510 (N_41510,N_40028,N_40816);
nand U41511 (N_41511,N_40356,N_40290);
and U41512 (N_41512,N_40972,N_40847);
and U41513 (N_41513,N_40553,N_40746);
nor U41514 (N_41514,N_40289,N_40102);
nand U41515 (N_41515,N_40980,N_40872);
xnor U41516 (N_41516,N_40699,N_40678);
or U41517 (N_41517,N_40928,N_40775);
nand U41518 (N_41518,N_40729,N_40725);
nor U41519 (N_41519,N_40496,N_40867);
and U41520 (N_41520,N_40511,N_40908);
nor U41521 (N_41521,N_40896,N_40716);
nand U41522 (N_41522,N_40088,N_40701);
nor U41523 (N_41523,N_40230,N_40955);
or U41524 (N_41524,N_40628,N_40986);
nand U41525 (N_41525,N_40020,N_40205);
xor U41526 (N_41526,N_40702,N_40441);
xnor U41527 (N_41527,N_40807,N_40915);
nand U41528 (N_41528,N_40566,N_40103);
or U41529 (N_41529,N_40837,N_40603);
nor U41530 (N_41530,N_40230,N_40144);
nand U41531 (N_41531,N_40825,N_40296);
xnor U41532 (N_41532,N_40659,N_40536);
and U41533 (N_41533,N_40156,N_40641);
and U41534 (N_41534,N_40610,N_40484);
xor U41535 (N_41535,N_40890,N_40541);
xnor U41536 (N_41536,N_40335,N_40574);
xnor U41537 (N_41537,N_40139,N_40881);
nand U41538 (N_41538,N_40051,N_40515);
and U41539 (N_41539,N_40305,N_40794);
xnor U41540 (N_41540,N_40541,N_40768);
xnor U41541 (N_41541,N_40048,N_40608);
xor U41542 (N_41542,N_40085,N_40811);
and U41543 (N_41543,N_40528,N_40316);
or U41544 (N_41544,N_40177,N_40092);
or U41545 (N_41545,N_40516,N_40443);
and U41546 (N_41546,N_40926,N_40514);
or U41547 (N_41547,N_40494,N_40728);
nand U41548 (N_41548,N_40659,N_40541);
nor U41549 (N_41549,N_40040,N_40324);
xor U41550 (N_41550,N_40209,N_40677);
nor U41551 (N_41551,N_40480,N_40973);
or U41552 (N_41552,N_40112,N_40134);
xor U41553 (N_41553,N_40687,N_40744);
xor U41554 (N_41554,N_40407,N_40493);
nand U41555 (N_41555,N_40894,N_40217);
xnor U41556 (N_41556,N_40076,N_40413);
xor U41557 (N_41557,N_40999,N_40780);
nor U41558 (N_41558,N_40287,N_40537);
nor U41559 (N_41559,N_40031,N_40217);
nor U41560 (N_41560,N_40970,N_40879);
nand U41561 (N_41561,N_40717,N_40636);
nor U41562 (N_41562,N_40075,N_40206);
and U41563 (N_41563,N_40631,N_40331);
nand U41564 (N_41564,N_40293,N_40549);
and U41565 (N_41565,N_40252,N_40967);
and U41566 (N_41566,N_40155,N_40467);
nand U41567 (N_41567,N_40930,N_40887);
xnor U41568 (N_41568,N_40546,N_40368);
nor U41569 (N_41569,N_40091,N_40481);
and U41570 (N_41570,N_40021,N_40198);
nand U41571 (N_41571,N_40799,N_40556);
and U41572 (N_41572,N_40604,N_40807);
nand U41573 (N_41573,N_40294,N_40794);
or U41574 (N_41574,N_40051,N_40869);
or U41575 (N_41575,N_40912,N_40217);
and U41576 (N_41576,N_40053,N_40385);
and U41577 (N_41577,N_40721,N_40822);
and U41578 (N_41578,N_40415,N_40268);
and U41579 (N_41579,N_40318,N_40958);
nor U41580 (N_41580,N_40605,N_40176);
and U41581 (N_41581,N_40349,N_40861);
nand U41582 (N_41582,N_40403,N_40854);
xor U41583 (N_41583,N_40727,N_40879);
or U41584 (N_41584,N_40822,N_40340);
or U41585 (N_41585,N_40607,N_40913);
xnor U41586 (N_41586,N_40676,N_40408);
nor U41587 (N_41587,N_40961,N_40529);
and U41588 (N_41588,N_40778,N_40485);
nand U41589 (N_41589,N_40918,N_40027);
or U41590 (N_41590,N_40645,N_40375);
and U41591 (N_41591,N_40887,N_40483);
nor U41592 (N_41592,N_40192,N_40455);
or U41593 (N_41593,N_40215,N_40423);
xor U41594 (N_41594,N_40722,N_40425);
nor U41595 (N_41595,N_40377,N_40853);
nor U41596 (N_41596,N_40718,N_40986);
nand U41597 (N_41597,N_40096,N_40535);
nor U41598 (N_41598,N_40903,N_40839);
nor U41599 (N_41599,N_40942,N_40314);
xor U41600 (N_41600,N_40854,N_40598);
nand U41601 (N_41601,N_40901,N_40685);
nand U41602 (N_41602,N_40416,N_40614);
xor U41603 (N_41603,N_40249,N_40955);
or U41604 (N_41604,N_40947,N_40405);
nor U41605 (N_41605,N_40495,N_40203);
or U41606 (N_41606,N_40319,N_40306);
nor U41607 (N_41607,N_40716,N_40699);
and U41608 (N_41608,N_40399,N_40617);
or U41609 (N_41609,N_40088,N_40612);
xor U41610 (N_41610,N_40831,N_40988);
and U41611 (N_41611,N_40689,N_40848);
or U41612 (N_41612,N_40035,N_40937);
xnor U41613 (N_41613,N_40036,N_40412);
nand U41614 (N_41614,N_40611,N_40966);
or U41615 (N_41615,N_40547,N_40273);
xor U41616 (N_41616,N_40293,N_40885);
and U41617 (N_41617,N_40474,N_40596);
and U41618 (N_41618,N_40265,N_40495);
nand U41619 (N_41619,N_40989,N_40281);
nor U41620 (N_41620,N_40956,N_40972);
nor U41621 (N_41621,N_40292,N_40205);
or U41622 (N_41622,N_40867,N_40895);
nor U41623 (N_41623,N_40387,N_40232);
and U41624 (N_41624,N_40999,N_40504);
and U41625 (N_41625,N_40371,N_40054);
nand U41626 (N_41626,N_40988,N_40507);
and U41627 (N_41627,N_40492,N_40589);
xnor U41628 (N_41628,N_40677,N_40752);
nor U41629 (N_41629,N_40354,N_40888);
nor U41630 (N_41630,N_40416,N_40575);
and U41631 (N_41631,N_40908,N_40206);
xor U41632 (N_41632,N_40476,N_40832);
nor U41633 (N_41633,N_40847,N_40383);
or U41634 (N_41634,N_40334,N_40917);
xor U41635 (N_41635,N_40607,N_40329);
nor U41636 (N_41636,N_40198,N_40253);
and U41637 (N_41637,N_40640,N_40435);
nor U41638 (N_41638,N_40214,N_40106);
or U41639 (N_41639,N_40637,N_40935);
and U41640 (N_41640,N_40214,N_40383);
or U41641 (N_41641,N_40584,N_40775);
xor U41642 (N_41642,N_40955,N_40877);
xor U41643 (N_41643,N_40569,N_40292);
and U41644 (N_41644,N_40745,N_40396);
xor U41645 (N_41645,N_40076,N_40863);
nand U41646 (N_41646,N_40297,N_40228);
xnor U41647 (N_41647,N_40228,N_40199);
xnor U41648 (N_41648,N_40995,N_40246);
nand U41649 (N_41649,N_40942,N_40712);
and U41650 (N_41650,N_40635,N_40407);
xnor U41651 (N_41651,N_40332,N_40923);
xor U41652 (N_41652,N_40550,N_40111);
or U41653 (N_41653,N_40970,N_40972);
nand U41654 (N_41654,N_40656,N_40526);
xnor U41655 (N_41655,N_40778,N_40213);
nor U41656 (N_41656,N_40150,N_40763);
nor U41657 (N_41657,N_40734,N_40335);
or U41658 (N_41658,N_40789,N_40560);
or U41659 (N_41659,N_40190,N_40004);
or U41660 (N_41660,N_40413,N_40850);
xor U41661 (N_41661,N_40098,N_40880);
or U41662 (N_41662,N_40634,N_40188);
or U41663 (N_41663,N_40508,N_40993);
nor U41664 (N_41664,N_40438,N_40883);
and U41665 (N_41665,N_40102,N_40264);
nor U41666 (N_41666,N_40646,N_40909);
nor U41667 (N_41667,N_40240,N_40640);
and U41668 (N_41668,N_40472,N_40710);
and U41669 (N_41669,N_40018,N_40533);
xor U41670 (N_41670,N_40799,N_40105);
and U41671 (N_41671,N_40735,N_40840);
or U41672 (N_41672,N_40635,N_40372);
and U41673 (N_41673,N_40595,N_40353);
or U41674 (N_41674,N_40211,N_40346);
nand U41675 (N_41675,N_40166,N_40918);
nor U41676 (N_41676,N_40051,N_40645);
or U41677 (N_41677,N_40803,N_40409);
and U41678 (N_41678,N_40960,N_40047);
or U41679 (N_41679,N_40341,N_40942);
xor U41680 (N_41680,N_40897,N_40202);
nor U41681 (N_41681,N_40890,N_40727);
or U41682 (N_41682,N_40094,N_40178);
or U41683 (N_41683,N_40822,N_40579);
and U41684 (N_41684,N_40134,N_40760);
nor U41685 (N_41685,N_40136,N_40856);
nor U41686 (N_41686,N_40242,N_40324);
and U41687 (N_41687,N_40621,N_40548);
or U41688 (N_41688,N_40027,N_40028);
nand U41689 (N_41689,N_40598,N_40207);
and U41690 (N_41690,N_40131,N_40084);
and U41691 (N_41691,N_40448,N_40494);
xor U41692 (N_41692,N_40813,N_40819);
nand U41693 (N_41693,N_40086,N_40769);
or U41694 (N_41694,N_40233,N_40053);
or U41695 (N_41695,N_40014,N_40579);
nand U41696 (N_41696,N_40928,N_40893);
nor U41697 (N_41697,N_40409,N_40705);
and U41698 (N_41698,N_40832,N_40780);
and U41699 (N_41699,N_40354,N_40246);
or U41700 (N_41700,N_40815,N_40444);
nor U41701 (N_41701,N_40356,N_40245);
or U41702 (N_41702,N_40207,N_40193);
nand U41703 (N_41703,N_40399,N_40469);
and U41704 (N_41704,N_40525,N_40406);
and U41705 (N_41705,N_40380,N_40401);
nand U41706 (N_41706,N_40646,N_40065);
or U41707 (N_41707,N_40379,N_40484);
or U41708 (N_41708,N_40757,N_40453);
and U41709 (N_41709,N_40134,N_40532);
or U41710 (N_41710,N_40352,N_40999);
nand U41711 (N_41711,N_40438,N_40260);
or U41712 (N_41712,N_40289,N_40835);
xor U41713 (N_41713,N_40823,N_40622);
nand U41714 (N_41714,N_40596,N_40091);
or U41715 (N_41715,N_40429,N_40141);
and U41716 (N_41716,N_40260,N_40429);
or U41717 (N_41717,N_40115,N_40440);
nand U41718 (N_41718,N_40144,N_40147);
xnor U41719 (N_41719,N_40199,N_40515);
or U41720 (N_41720,N_40224,N_40067);
nor U41721 (N_41721,N_40147,N_40213);
xor U41722 (N_41722,N_40489,N_40224);
nand U41723 (N_41723,N_40588,N_40158);
xnor U41724 (N_41724,N_40585,N_40933);
nand U41725 (N_41725,N_40907,N_40832);
nor U41726 (N_41726,N_40412,N_40501);
and U41727 (N_41727,N_40205,N_40557);
nor U41728 (N_41728,N_40952,N_40609);
xor U41729 (N_41729,N_40315,N_40294);
or U41730 (N_41730,N_40894,N_40178);
nand U41731 (N_41731,N_40268,N_40798);
xor U41732 (N_41732,N_40732,N_40422);
nand U41733 (N_41733,N_40563,N_40789);
xnor U41734 (N_41734,N_40237,N_40242);
nor U41735 (N_41735,N_40601,N_40287);
nand U41736 (N_41736,N_40917,N_40753);
and U41737 (N_41737,N_40534,N_40790);
or U41738 (N_41738,N_40622,N_40504);
or U41739 (N_41739,N_40164,N_40319);
nor U41740 (N_41740,N_40223,N_40939);
nand U41741 (N_41741,N_40738,N_40241);
or U41742 (N_41742,N_40571,N_40278);
nor U41743 (N_41743,N_40144,N_40662);
xnor U41744 (N_41744,N_40135,N_40866);
nor U41745 (N_41745,N_40249,N_40150);
xnor U41746 (N_41746,N_40857,N_40617);
and U41747 (N_41747,N_40055,N_40343);
xnor U41748 (N_41748,N_40508,N_40261);
nand U41749 (N_41749,N_40615,N_40095);
xnor U41750 (N_41750,N_40076,N_40362);
nand U41751 (N_41751,N_40500,N_40735);
or U41752 (N_41752,N_40202,N_40873);
or U41753 (N_41753,N_40198,N_40283);
xor U41754 (N_41754,N_40569,N_40100);
or U41755 (N_41755,N_40383,N_40402);
and U41756 (N_41756,N_40140,N_40759);
nand U41757 (N_41757,N_40034,N_40172);
nand U41758 (N_41758,N_40046,N_40755);
nand U41759 (N_41759,N_40530,N_40271);
xor U41760 (N_41760,N_40216,N_40726);
xor U41761 (N_41761,N_40795,N_40705);
nor U41762 (N_41762,N_40696,N_40738);
nand U41763 (N_41763,N_40878,N_40102);
xnor U41764 (N_41764,N_40355,N_40820);
nand U41765 (N_41765,N_40462,N_40079);
and U41766 (N_41766,N_40005,N_40600);
nor U41767 (N_41767,N_40049,N_40362);
and U41768 (N_41768,N_40207,N_40397);
nand U41769 (N_41769,N_40556,N_40834);
nor U41770 (N_41770,N_40859,N_40875);
nand U41771 (N_41771,N_40731,N_40897);
nand U41772 (N_41772,N_40553,N_40079);
xor U41773 (N_41773,N_40472,N_40390);
and U41774 (N_41774,N_40337,N_40177);
nor U41775 (N_41775,N_40363,N_40713);
nor U41776 (N_41776,N_40820,N_40100);
or U41777 (N_41777,N_40060,N_40302);
nand U41778 (N_41778,N_40376,N_40912);
xnor U41779 (N_41779,N_40504,N_40781);
nand U41780 (N_41780,N_40922,N_40650);
xor U41781 (N_41781,N_40014,N_40710);
and U41782 (N_41782,N_40032,N_40338);
and U41783 (N_41783,N_40481,N_40516);
nand U41784 (N_41784,N_40181,N_40042);
xor U41785 (N_41785,N_40585,N_40830);
or U41786 (N_41786,N_40923,N_40213);
nor U41787 (N_41787,N_40949,N_40883);
nand U41788 (N_41788,N_40257,N_40440);
xor U41789 (N_41789,N_40058,N_40386);
and U41790 (N_41790,N_40399,N_40885);
xnor U41791 (N_41791,N_40263,N_40271);
or U41792 (N_41792,N_40191,N_40107);
nor U41793 (N_41793,N_40833,N_40737);
xnor U41794 (N_41794,N_40184,N_40104);
nand U41795 (N_41795,N_40734,N_40178);
or U41796 (N_41796,N_40268,N_40047);
nand U41797 (N_41797,N_40860,N_40953);
nand U41798 (N_41798,N_40144,N_40219);
xor U41799 (N_41799,N_40175,N_40695);
and U41800 (N_41800,N_40443,N_40168);
xor U41801 (N_41801,N_40051,N_40962);
and U41802 (N_41802,N_40536,N_40458);
and U41803 (N_41803,N_40356,N_40052);
nor U41804 (N_41804,N_40846,N_40629);
or U41805 (N_41805,N_40449,N_40180);
or U41806 (N_41806,N_40536,N_40187);
nor U41807 (N_41807,N_40722,N_40857);
nor U41808 (N_41808,N_40810,N_40185);
nor U41809 (N_41809,N_40803,N_40450);
and U41810 (N_41810,N_40608,N_40875);
nor U41811 (N_41811,N_40272,N_40056);
or U41812 (N_41812,N_40439,N_40848);
nor U41813 (N_41813,N_40831,N_40592);
xnor U41814 (N_41814,N_40604,N_40490);
or U41815 (N_41815,N_40770,N_40001);
nand U41816 (N_41816,N_40986,N_40029);
nor U41817 (N_41817,N_40892,N_40182);
xor U41818 (N_41818,N_40449,N_40270);
or U41819 (N_41819,N_40068,N_40608);
and U41820 (N_41820,N_40274,N_40704);
and U41821 (N_41821,N_40612,N_40892);
or U41822 (N_41822,N_40488,N_40027);
or U41823 (N_41823,N_40168,N_40752);
nand U41824 (N_41824,N_40616,N_40994);
nand U41825 (N_41825,N_40548,N_40317);
nor U41826 (N_41826,N_40527,N_40234);
xnor U41827 (N_41827,N_40757,N_40233);
xnor U41828 (N_41828,N_40990,N_40431);
nand U41829 (N_41829,N_40478,N_40302);
nand U41830 (N_41830,N_40411,N_40658);
xnor U41831 (N_41831,N_40671,N_40140);
and U41832 (N_41832,N_40807,N_40226);
or U41833 (N_41833,N_40797,N_40617);
or U41834 (N_41834,N_40328,N_40487);
xnor U41835 (N_41835,N_40052,N_40060);
and U41836 (N_41836,N_40392,N_40141);
and U41837 (N_41837,N_40890,N_40869);
xor U41838 (N_41838,N_40977,N_40271);
nor U41839 (N_41839,N_40037,N_40622);
or U41840 (N_41840,N_40267,N_40008);
nand U41841 (N_41841,N_40263,N_40462);
or U41842 (N_41842,N_40080,N_40692);
or U41843 (N_41843,N_40826,N_40344);
or U41844 (N_41844,N_40586,N_40999);
or U41845 (N_41845,N_40843,N_40129);
or U41846 (N_41846,N_40174,N_40772);
and U41847 (N_41847,N_40103,N_40465);
xor U41848 (N_41848,N_40681,N_40089);
or U41849 (N_41849,N_40998,N_40344);
xnor U41850 (N_41850,N_40408,N_40368);
nor U41851 (N_41851,N_40931,N_40134);
or U41852 (N_41852,N_40699,N_40229);
and U41853 (N_41853,N_40452,N_40460);
nor U41854 (N_41854,N_40941,N_40840);
and U41855 (N_41855,N_40476,N_40932);
and U41856 (N_41856,N_40073,N_40687);
or U41857 (N_41857,N_40111,N_40392);
xor U41858 (N_41858,N_40215,N_40295);
nor U41859 (N_41859,N_40311,N_40026);
nand U41860 (N_41860,N_40644,N_40067);
nand U41861 (N_41861,N_40196,N_40802);
nand U41862 (N_41862,N_40682,N_40644);
nand U41863 (N_41863,N_40339,N_40997);
or U41864 (N_41864,N_40444,N_40829);
nand U41865 (N_41865,N_40272,N_40921);
nor U41866 (N_41866,N_40893,N_40565);
nor U41867 (N_41867,N_40795,N_40929);
or U41868 (N_41868,N_40239,N_40245);
nand U41869 (N_41869,N_40739,N_40732);
or U41870 (N_41870,N_40141,N_40518);
and U41871 (N_41871,N_40760,N_40907);
and U41872 (N_41872,N_40553,N_40924);
nand U41873 (N_41873,N_40204,N_40190);
nor U41874 (N_41874,N_40762,N_40747);
or U41875 (N_41875,N_40862,N_40790);
xor U41876 (N_41876,N_40771,N_40717);
or U41877 (N_41877,N_40980,N_40576);
xor U41878 (N_41878,N_40375,N_40911);
and U41879 (N_41879,N_40715,N_40795);
xnor U41880 (N_41880,N_40830,N_40967);
or U41881 (N_41881,N_40508,N_40269);
or U41882 (N_41882,N_40932,N_40812);
or U41883 (N_41883,N_40744,N_40705);
nand U41884 (N_41884,N_40446,N_40288);
xnor U41885 (N_41885,N_40343,N_40745);
nor U41886 (N_41886,N_40595,N_40092);
nand U41887 (N_41887,N_40898,N_40093);
or U41888 (N_41888,N_40296,N_40421);
nor U41889 (N_41889,N_40759,N_40692);
nor U41890 (N_41890,N_40489,N_40970);
xnor U41891 (N_41891,N_40762,N_40321);
nor U41892 (N_41892,N_40648,N_40083);
and U41893 (N_41893,N_40982,N_40916);
nand U41894 (N_41894,N_40452,N_40323);
nand U41895 (N_41895,N_40019,N_40863);
and U41896 (N_41896,N_40247,N_40771);
xnor U41897 (N_41897,N_40111,N_40623);
and U41898 (N_41898,N_40866,N_40160);
xnor U41899 (N_41899,N_40905,N_40105);
or U41900 (N_41900,N_40406,N_40728);
xnor U41901 (N_41901,N_40838,N_40944);
xnor U41902 (N_41902,N_40633,N_40552);
xor U41903 (N_41903,N_40138,N_40603);
nor U41904 (N_41904,N_40022,N_40303);
and U41905 (N_41905,N_40804,N_40471);
or U41906 (N_41906,N_40766,N_40589);
and U41907 (N_41907,N_40266,N_40609);
xnor U41908 (N_41908,N_40459,N_40315);
or U41909 (N_41909,N_40356,N_40426);
nor U41910 (N_41910,N_40999,N_40576);
nor U41911 (N_41911,N_40956,N_40502);
xnor U41912 (N_41912,N_40438,N_40658);
and U41913 (N_41913,N_40840,N_40663);
nand U41914 (N_41914,N_40202,N_40911);
and U41915 (N_41915,N_40012,N_40024);
and U41916 (N_41916,N_40830,N_40514);
nand U41917 (N_41917,N_40301,N_40991);
xnor U41918 (N_41918,N_40864,N_40164);
xnor U41919 (N_41919,N_40656,N_40965);
and U41920 (N_41920,N_40604,N_40583);
nand U41921 (N_41921,N_40976,N_40485);
xor U41922 (N_41922,N_40224,N_40566);
nor U41923 (N_41923,N_40565,N_40703);
or U41924 (N_41924,N_40438,N_40570);
nand U41925 (N_41925,N_40032,N_40582);
and U41926 (N_41926,N_40623,N_40486);
and U41927 (N_41927,N_40198,N_40953);
xnor U41928 (N_41928,N_40654,N_40647);
or U41929 (N_41929,N_40918,N_40840);
xor U41930 (N_41930,N_40216,N_40985);
nand U41931 (N_41931,N_40680,N_40098);
and U41932 (N_41932,N_40501,N_40682);
and U41933 (N_41933,N_40668,N_40100);
xor U41934 (N_41934,N_40988,N_40196);
or U41935 (N_41935,N_40642,N_40512);
or U41936 (N_41936,N_40987,N_40464);
nand U41937 (N_41937,N_40832,N_40317);
xor U41938 (N_41938,N_40932,N_40853);
nor U41939 (N_41939,N_40207,N_40246);
or U41940 (N_41940,N_40411,N_40318);
xor U41941 (N_41941,N_40614,N_40266);
nor U41942 (N_41942,N_40117,N_40095);
or U41943 (N_41943,N_40589,N_40232);
and U41944 (N_41944,N_40378,N_40249);
or U41945 (N_41945,N_40403,N_40638);
and U41946 (N_41946,N_40578,N_40388);
nor U41947 (N_41947,N_40377,N_40657);
and U41948 (N_41948,N_40297,N_40143);
nand U41949 (N_41949,N_40344,N_40050);
or U41950 (N_41950,N_40780,N_40004);
xor U41951 (N_41951,N_40005,N_40104);
nor U41952 (N_41952,N_40795,N_40001);
or U41953 (N_41953,N_40673,N_40445);
nor U41954 (N_41954,N_40775,N_40233);
and U41955 (N_41955,N_40490,N_40004);
or U41956 (N_41956,N_40837,N_40179);
nand U41957 (N_41957,N_40618,N_40508);
nand U41958 (N_41958,N_40898,N_40753);
xnor U41959 (N_41959,N_40626,N_40781);
xor U41960 (N_41960,N_40957,N_40910);
nand U41961 (N_41961,N_40858,N_40789);
nand U41962 (N_41962,N_40747,N_40966);
nand U41963 (N_41963,N_40106,N_40244);
xnor U41964 (N_41964,N_40321,N_40200);
or U41965 (N_41965,N_40699,N_40579);
nand U41966 (N_41966,N_40714,N_40093);
and U41967 (N_41967,N_40234,N_40570);
or U41968 (N_41968,N_40872,N_40934);
nor U41969 (N_41969,N_40612,N_40190);
nor U41970 (N_41970,N_40676,N_40635);
nand U41971 (N_41971,N_40655,N_40682);
nand U41972 (N_41972,N_40405,N_40389);
and U41973 (N_41973,N_40389,N_40060);
nor U41974 (N_41974,N_40309,N_40879);
and U41975 (N_41975,N_40836,N_40046);
nand U41976 (N_41976,N_40674,N_40873);
xor U41977 (N_41977,N_40344,N_40938);
nor U41978 (N_41978,N_40087,N_40979);
or U41979 (N_41979,N_40024,N_40011);
and U41980 (N_41980,N_40071,N_40610);
xnor U41981 (N_41981,N_40617,N_40997);
nand U41982 (N_41982,N_40458,N_40126);
nor U41983 (N_41983,N_40604,N_40710);
nand U41984 (N_41984,N_40292,N_40609);
nand U41985 (N_41985,N_40769,N_40468);
and U41986 (N_41986,N_40162,N_40812);
nor U41987 (N_41987,N_40948,N_40648);
xor U41988 (N_41988,N_40679,N_40440);
nand U41989 (N_41989,N_40133,N_40870);
nand U41990 (N_41990,N_40806,N_40788);
and U41991 (N_41991,N_40811,N_40906);
nor U41992 (N_41992,N_40154,N_40076);
and U41993 (N_41993,N_40770,N_40918);
or U41994 (N_41994,N_40085,N_40050);
or U41995 (N_41995,N_40140,N_40885);
nor U41996 (N_41996,N_40179,N_40100);
and U41997 (N_41997,N_40349,N_40737);
nand U41998 (N_41998,N_40283,N_40672);
xor U41999 (N_41999,N_40411,N_40354);
and U42000 (N_42000,N_41832,N_41576);
nand U42001 (N_42001,N_41872,N_41676);
or U42002 (N_42002,N_41352,N_41298);
nor U42003 (N_42003,N_41067,N_41121);
xnor U42004 (N_42004,N_41213,N_41010);
nand U42005 (N_42005,N_41146,N_41571);
or U42006 (N_42006,N_41349,N_41488);
nand U42007 (N_42007,N_41995,N_41024);
xor U42008 (N_42008,N_41294,N_41757);
and U42009 (N_42009,N_41268,N_41137);
or U42010 (N_42010,N_41651,N_41749);
xor U42011 (N_42011,N_41653,N_41627);
and U42012 (N_42012,N_41307,N_41562);
xnor U42013 (N_42013,N_41136,N_41492);
and U42014 (N_42014,N_41177,N_41385);
or U42015 (N_42015,N_41343,N_41302);
nand U42016 (N_42016,N_41672,N_41145);
or U42017 (N_42017,N_41109,N_41845);
nand U42018 (N_42018,N_41489,N_41537);
nand U42019 (N_42019,N_41965,N_41120);
and U42020 (N_42020,N_41181,N_41870);
and U42021 (N_42021,N_41310,N_41604);
nand U42022 (N_42022,N_41432,N_41284);
and U42023 (N_42023,N_41303,N_41950);
xnor U42024 (N_42024,N_41191,N_41320);
xnor U42025 (N_42025,N_41457,N_41700);
nand U42026 (N_42026,N_41028,N_41392);
nand U42027 (N_42027,N_41007,N_41732);
xnor U42028 (N_42028,N_41205,N_41463);
nor U42029 (N_42029,N_41591,N_41214);
or U42030 (N_42030,N_41211,N_41923);
xnor U42031 (N_42031,N_41018,N_41776);
and U42032 (N_42032,N_41270,N_41227);
nand U42033 (N_42033,N_41274,N_41476);
and U42034 (N_42034,N_41161,N_41770);
nand U42035 (N_42035,N_41331,N_41056);
and U42036 (N_42036,N_41173,N_41623);
xnor U42037 (N_42037,N_41958,N_41301);
and U42038 (N_42038,N_41053,N_41740);
nor U42039 (N_42039,N_41922,N_41269);
or U42040 (N_42040,N_41397,N_41513);
nand U42041 (N_42041,N_41600,N_41896);
xnor U42042 (N_42042,N_41273,N_41806);
nand U42043 (N_42043,N_41322,N_41708);
nand U42044 (N_42044,N_41547,N_41127);
xnor U42045 (N_42045,N_41663,N_41532);
and U42046 (N_42046,N_41005,N_41744);
and U42047 (N_42047,N_41999,N_41157);
and U42048 (N_42048,N_41012,N_41366);
nor U42049 (N_42049,N_41128,N_41856);
or U42050 (N_42050,N_41855,N_41490);
xnor U42051 (N_42051,N_41761,N_41792);
or U42052 (N_42052,N_41427,N_41168);
xor U42053 (N_42053,N_41854,N_41277);
nand U42054 (N_42054,N_41890,N_41839);
or U42055 (N_42055,N_41686,N_41529);
nand U42056 (N_42056,N_41106,N_41675);
nand U42057 (N_42057,N_41207,N_41802);
and U42058 (N_42058,N_41324,N_41059);
or U42059 (N_42059,N_41011,N_41748);
or U42060 (N_42060,N_41687,N_41539);
nor U42061 (N_42061,N_41071,N_41710);
nand U42062 (N_42062,N_41047,N_41596);
or U42063 (N_42063,N_41875,N_41518);
and U42064 (N_42064,N_41286,N_41643);
nand U42065 (N_42065,N_41479,N_41815);
and U42066 (N_42066,N_41448,N_41200);
or U42067 (N_42067,N_41662,N_41620);
nand U42068 (N_42068,N_41455,N_41008);
or U42069 (N_42069,N_41739,N_41543);
and U42070 (N_42070,N_41674,N_41756);
nor U42071 (N_42071,N_41393,N_41718);
or U42072 (N_42072,N_41658,N_41158);
nor U42073 (N_42073,N_41131,N_41206);
nor U42074 (N_42074,N_41068,N_41225);
and U42075 (N_42075,N_41753,N_41064);
xnor U42076 (N_42076,N_41616,N_41458);
nand U42077 (N_42077,N_41116,N_41791);
and U42078 (N_42078,N_41775,N_41682);
nor U42079 (N_42079,N_41172,N_41678);
or U42080 (N_42080,N_41553,N_41525);
or U42081 (N_42081,N_41486,N_41997);
and U42082 (N_42082,N_41223,N_41696);
and U42083 (N_42083,N_41218,N_41006);
and U42084 (N_42084,N_41783,N_41951);
and U42085 (N_42085,N_41454,N_41669);
nor U42086 (N_42086,N_41926,N_41285);
nand U42087 (N_42087,N_41555,N_41257);
xnor U42088 (N_42088,N_41716,N_41793);
nand U42089 (N_42089,N_41305,N_41849);
xor U42090 (N_42090,N_41969,N_41074);
xor U42091 (N_42091,N_41795,N_41924);
nor U42092 (N_42092,N_41196,N_41641);
nor U42093 (N_42093,N_41626,N_41515);
nor U42094 (N_42094,N_41765,N_41729);
and U42095 (N_42095,N_41557,N_41814);
and U42096 (N_42096,N_41968,N_41750);
or U42097 (N_42097,N_41022,N_41085);
nand U42098 (N_42098,N_41424,N_41873);
xnor U42099 (N_42099,N_41467,N_41735);
or U42100 (N_42100,N_41745,N_41818);
nand U42101 (N_42101,N_41866,N_41099);
and U42102 (N_42102,N_41603,N_41692);
or U42103 (N_42103,N_41523,N_41142);
xor U42104 (N_42104,N_41962,N_41649);
xnor U42105 (N_42105,N_41003,N_41259);
nand U42106 (N_42106,N_41420,N_41434);
nand U42107 (N_42107,N_41703,N_41433);
or U42108 (N_42108,N_41879,N_41248);
or U42109 (N_42109,N_41595,N_41645);
nor U42110 (N_42110,N_41789,N_41988);
and U42111 (N_42111,N_41367,N_41278);
or U42112 (N_42112,N_41378,N_41408);
and U42113 (N_42113,N_41382,N_41138);
nand U42114 (N_42114,N_41607,N_41258);
nor U42115 (N_42115,N_41377,N_41484);
nand U42116 (N_42116,N_41837,N_41981);
or U42117 (N_42117,N_41226,N_41154);
nor U42118 (N_42118,N_41567,N_41833);
and U42119 (N_42119,N_41251,N_41246);
nor U42120 (N_42120,N_41705,N_41544);
and U42121 (N_42121,N_41722,N_41133);
nor U42122 (N_42122,N_41029,N_41334);
nand U42123 (N_42123,N_41185,N_41817);
xnor U42124 (N_42124,N_41400,N_41861);
nand U42125 (N_42125,N_41395,N_41491);
nand U42126 (N_42126,N_41894,N_41994);
or U42127 (N_42127,N_41344,N_41664);
or U42128 (N_42128,N_41680,N_41319);
nand U42129 (N_42129,N_41097,N_41394);
or U42130 (N_42130,N_41572,N_41409);
nor U42131 (N_42131,N_41459,N_41289);
and U42132 (N_42132,N_41528,N_41510);
nand U42133 (N_42133,N_41117,N_41216);
and U42134 (N_42134,N_41465,N_41410);
nand U42135 (N_42135,N_41418,N_41880);
nand U42136 (N_42136,N_41032,N_41501);
or U42137 (N_42137,N_41020,N_41838);
and U42138 (N_42138,N_41220,N_41590);
nor U42139 (N_42139,N_41721,N_41039);
xnor U42140 (N_42140,N_41914,N_41581);
xor U42141 (N_42141,N_41396,N_41611);
xor U42142 (N_42142,N_41940,N_41785);
nand U42143 (N_42143,N_41639,N_41790);
nor U42144 (N_42144,N_41188,N_41704);
or U42145 (N_42145,N_41228,N_41186);
nand U42146 (N_42146,N_41874,N_41497);
xor U42147 (N_42147,N_41964,N_41036);
xor U42148 (N_42148,N_41784,N_41253);
nand U42149 (N_42149,N_41470,N_41862);
nand U42150 (N_42150,N_41435,N_41391);
nand U42151 (N_42151,N_41506,N_41573);
nand U42152 (N_42152,N_41095,N_41564);
xor U42153 (N_42153,N_41473,N_41827);
nand U42154 (N_42154,N_41939,N_41851);
nor U42155 (N_42155,N_41451,N_41925);
nor U42156 (N_42156,N_41709,N_41545);
xnor U42157 (N_42157,N_41163,N_41415);
xnor U42158 (N_42158,N_41612,N_41853);
xnor U42159 (N_42159,N_41916,N_41799);
nand U42160 (N_42160,N_41593,N_41072);
nor U42161 (N_42161,N_41605,N_41934);
nor U42162 (N_42162,N_41453,N_41919);
or U42163 (N_42163,N_41566,N_41149);
nand U42164 (N_42164,N_41941,N_41647);
nor U42165 (N_42165,N_41857,N_41660);
and U42166 (N_42166,N_41671,N_41297);
or U42167 (N_42167,N_41222,N_41265);
and U42168 (N_42168,N_41254,N_41530);
nand U42169 (N_42169,N_41897,N_41909);
or U42170 (N_42170,N_41494,N_41772);
nand U42171 (N_42171,N_41498,N_41824);
nor U42172 (N_42172,N_41483,N_41374);
and U42173 (N_42173,N_41113,N_41014);
and U42174 (N_42174,N_41867,N_41899);
nor U42175 (N_42175,N_41742,N_41780);
or U42176 (N_42176,N_41840,N_41267);
or U42177 (N_42177,N_41670,N_41440);
nand U42178 (N_42178,N_41821,N_41697);
nor U42179 (N_42179,N_41954,N_41130);
and U42180 (N_42180,N_41974,N_41743);
or U42181 (N_42181,N_41438,N_41288);
nand U42182 (N_42182,N_41648,N_41215);
or U42183 (N_42183,N_41192,N_41630);
xor U42184 (N_42184,N_41040,N_41217);
xnor U42185 (N_42185,N_41868,N_41747);
nor U42186 (N_42186,N_41906,N_41579);
xor U42187 (N_42187,N_41235,N_41797);
nor U42188 (N_42188,N_41808,N_41164);
nand U42189 (N_42189,N_41122,N_41715);
nand U42190 (N_42190,N_41401,N_41548);
xor U42191 (N_42191,N_41066,N_41147);
nor U42192 (N_42192,N_41668,N_41758);
or U42193 (N_42193,N_41160,N_41816);
or U42194 (N_42194,N_41930,N_41144);
and U42195 (N_42195,N_41437,N_41842);
nand U42196 (N_42196,N_41339,N_41025);
xnor U42197 (N_42197,N_41688,N_41631);
xnor U42198 (N_42198,N_41293,N_41300);
nor U42199 (N_42199,N_41195,N_41625);
xor U42200 (N_42200,N_41991,N_41464);
and U42201 (N_42201,N_41614,N_41290);
nor U42202 (N_42202,N_41524,N_41610);
nor U42203 (N_42203,N_41657,N_41929);
xnor U42204 (N_42204,N_41000,N_41233);
or U42205 (N_42205,N_41586,N_41738);
nand U42206 (N_42206,N_41460,N_41315);
and U42207 (N_42207,N_41256,N_41520);
and U42208 (N_42208,N_41667,N_41650);
nand U42209 (N_42209,N_41019,N_41219);
xnor U42210 (N_42210,N_41683,N_41993);
xnor U42211 (N_42211,N_41666,N_41264);
and U42212 (N_42212,N_41035,N_41174);
or U42213 (N_42213,N_41013,N_41055);
xor U42214 (N_42214,N_41419,N_41900);
or U42215 (N_42215,N_41159,N_41370);
xor U42216 (N_42216,N_41541,N_41860);
nor U42217 (N_42217,N_41957,N_41504);
and U42218 (N_42218,N_41752,N_41231);
xor U42219 (N_42219,N_41945,N_41794);
and U42220 (N_42220,N_41803,N_41338);
xnor U42221 (N_42221,N_41517,N_41788);
nand U42222 (N_42222,N_41746,N_41632);
or U42223 (N_42223,N_41594,N_41921);
or U42224 (N_42224,N_41684,N_41706);
nand U42225 (N_42225,N_41613,N_41078);
xnor U42226 (N_42226,N_41852,N_41445);
and U42227 (N_42227,N_41111,N_41077);
nor U42228 (N_42228,N_41883,N_41255);
and U42229 (N_42229,N_41920,N_41287);
xnor U42230 (N_42230,N_41076,N_41864);
nand U42231 (N_42231,N_41618,N_41054);
nor U42232 (N_42232,N_41332,N_41058);
and U42233 (N_42233,N_41953,N_41034);
or U42234 (N_42234,N_41977,N_41243);
or U42235 (N_42235,N_41830,N_41110);
nor U42236 (N_42236,N_41903,N_41907);
nor U42237 (N_42237,N_41291,N_41232);
nand U42238 (N_42238,N_41578,N_41328);
or U42239 (N_42239,N_41519,N_41850);
or U42240 (N_42240,N_41779,N_41033);
nor U42241 (N_42241,N_41681,N_41405);
and U42242 (N_42242,N_41351,N_41070);
and U42243 (N_42243,N_41889,N_41182);
or U42244 (N_42244,N_41937,N_41083);
xor U42245 (N_42245,N_41314,N_41597);
and U42246 (N_42246,N_41134,N_41713);
nor U42247 (N_42247,N_41725,N_41026);
or U42248 (N_42248,N_41089,N_41888);
and U42249 (N_42249,N_41598,N_41282);
and U42250 (N_42250,N_41622,N_41183);
and U42251 (N_42251,N_41933,N_41084);
xnor U42252 (N_42252,N_41781,N_41549);
nand U42253 (N_42253,N_41398,N_41534);
or U42254 (N_42254,N_41493,N_41644);
and U42255 (N_42255,N_41296,N_41912);
nor U42256 (N_42256,N_41263,N_41638);
nand U42257 (N_42257,N_41295,N_41364);
and U42258 (N_42258,N_41093,N_41201);
nor U42259 (N_42259,N_41156,N_41987);
nor U42260 (N_42260,N_41998,N_41751);
and U42261 (N_42261,N_41902,N_41325);
nand U42262 (N_42262,N_41221,N_41601);
xor U42263 (N_42263,N_41387,N_41375);
nor U42264 (N_42264,N_41565,N_41811);
and U42265 (N_42265,N_41487,N_41737);
nor U42266 (N_42266,N_41730,N_41475);
and U42267 (N_42267,N_41354,N_41885);
nor U42268 (N_42268,N_41979,N_41826);
and U42269 (N_42269,N_41004,N_41368);
or U42270 (N_42270,N_41384,N_41380);
nand U42271 (N_42271,N_41238,N_41376);
xor U42272 (N_42272,N_41948,N_41234);
xor U42273 (N_42273,N_41661,N_41762);
or U42274 (N_42274,N_41125,N_41834);
xor U42275 (N_42275,N_41119,N_41037);
nand U42276 (N_42276,N_41496,N_41786);
and U42277 (N_42277,N_41240,N_41720);
xnor U42278 (N_42278,N_41043,N_41190);
or U42279 (N_42279,N_41558,N_41984);
or U42280 (N_42280,N_41442,N_41800);
nand U42281 (N_42281,N_41402,N_41150);
nand U42282 (N_42282,N_41098,N_41279);
nand U42283 (N_42283,N_41015,N_41414);
or U42284 (N_42284,N_41229,N_41444);
nor U42285 (N_42285,N_41304,N_41561);
nand U42286 (N_42286,N_41430,N_41989);
nor U42287 (N_42287,N_41313,N_41471);
nor U42288 (N_42288,N_41169,N_41946);
and U42289 (N_42289,N_41973,N_41699);
nand U42290 (N_42290,N_41423,N_41355);
nand U42291 (N_42291,N_41049,N_41373);
or U42292 (N_42292,N_41245,N_41927);
xnor U42293 (N_42293,N_41938,N_41717);
nand U42294 (N_42294,N_41193,N_41166);
nor U42295 (N_42295,N_41139,N_41918);
nand U42296 (N_42296,N_41230,N_41947);
xor U42297 (N_42297,N_41952,N_41412);
nor U42298 (N_42298,N_41508,N_41171);
or U42299 (N_42299,N_41386,N_41416);
xor U42300 (N_42300,N_41411,N_41798);
or U42301 (N_42301,N_41905,N_41642);
or U42302 (N_42302,N_41371,N_41346);
nand U42303 (N_42303,N_41949,N_41353);
or U42304 (N_42304,N_41810,N_41428);
or U42305 (N_42305,N_41091,N_41406);
nor U42306 (N_42306,N_41859,N_41865);
xnor U42307 (N_42307,N_41199,N_41509);
nand U42308 (N_42308,N_41082,N_41820);
or U42309 (N_42309,N_41580,N_41760);
nand U42310 (N_42310,N_41107,N_41863);
nor U42311 (N_42311,N_41970,N_41882);
and U42312 (N_42312,N_41341,N_41679);
and U42313 (N_42313,N_41698,N_41694);
nor U42314 (N_42314,N_41844,N_41503);
nor U42315 (N_42315,N_41990,N_41691);
or U42316 (N_42316,N_41148,N_41809);
xnor U42317 (N_42317,N_41212,N_41407);
or U42318 (N_42318,N_41050,N_41773);
and U42319 (N_42319,N_41321,N_41101);
or U42320 (N_42320,N_41009,N_41726);
nor U42321 (N_42321,N_41724,N_41075);
xor U42322 (N_42322,N_41027,N_41575);
nor U42323 (N_42323,N_41330,N_41847);
and U42324 (N_42324,N_41031,N_41333);
nand U42325 (N_42325,N_41777,N_41335);
or U42326 (N_42326,N_41858,N_41108);
nor U42327 (N_42327,N_41813,N_41249);
nor U42328 (N_42328,N_41659,N_41123);
xor U42329 (N_42329,N_41461,N_41105);
or U42330 (N_42330,N_41309,N_41345);
xnor U42331 (N_42331,N_41702,N_41928);
and U42332 (N_42332,N_41262,N_41224);
xor U42333 (N_42333,N_41250,N_41733);
or U42334 (N_42334,N_41372,N_41546);
nor U42335 (N_42335,N_41568,N_41976);
or U42336 (N_42336,N_41689,N_41425);
and U42337 (N_42337,N_41045,N_41707);
xor U42338 (N_42338,N_41356,N_41589);
nor U42339 (N_42339,N_41961,N_41359);
and U42340 (N_42340,N_41104,N_41090);
xor U42341 (N_42341,N_41980,N_41329);
xnor U42342 (N_42342,N_41271,N_41507);
nor U42343 (N_42343,N_41087,N_41871);
or U42344 (N_42344,N_41311,N_41768);
or U42345 (N_42345,N_41538,N_41540);
nor U42346 (N_42346,N_41363,N_41094);
nor U42347 (N_42347,N_41065,N_41841);
nand U42348 (N_42348,N_41898,N_41472);
and U42349 (N_42349,N_41462,N_41450);
or U42350 (N_42350,N_41646,N_41584);
nor U42351 (N_42351,N_41261,N_41505);
or U42352 (N_42352,N_41426,N_41550);
nor U42353 (N_42353,N_41711,N_41551);
nor U42354 (N_42354,N_41624,N_41609);
and U42355 (N_42355,N_41088,N_41046);
or U42356 (N_42356,N_41061,N_41619);
nand U42357 (N_42357,N_41381,N_41782);
nor U42358 (N_42358,N_41978,N_41588);
nor U42359 (N_42359,N_41244,N_41975);
nor U42360 (N_42360,N_41723,N_41592);
and U42361 (N_42361,N_41560,N_41308);
or U42362 (N_42362,N_41512,N_41996);
xor U42363 (N_42363,N_41983,N_41365);
nand U42364 (N_42364,N_41500,N_41379);
and U42365 (N_42365,N_41608,N_41876);
and U42366 (N_42366,N_41629,N_41469);
nand U42367 (N_42367,N_41347,N_41092);
nand U42368 (N_42368,N_41281,N_41202);
xor U42369 (N_42369,N_41985,N_41892);
xnor U42370 (N_42370,N_41931,N_41362);
and U42371 (N_42371,N_41327,N_41812);
nor U42372 (N_42372,N_41051,N_41100);
nand U42373 (N_42373,N_41252,N_41038);
nand U42374 (N_42374,N_41165,N_41102);
or U42375 (N_42375,N_41485,N_41966);
nor U42376 (N_42376,N_41162,N_41655);
nand U42377 (N_42377,N_41640,N_41570);
nand U42378 (N_42378,N_41153,N_41001);
and U42379 (N_42379,N_41178,N_41474);
nand U42380 (N_42380,N_41348,N_41615);
nand U42381 (N_42381,N_41736,N_41701);
xnor U42382 (N_42382,N_41621,N_41060);
nor U42383 (N_42383,N_41917,N_41413);
or U42384 (N_42384,N_41477,N_41495);
and U42385 (N_42385,N_41714,N_41283);
nand U42386 (N_42386,N_41911,N_41151);
nand U42387 (N_42387,N_41357,N_41441);
and U42388 (N_42388,N_41446,N_41637);
nand U42389 (N_42389,N_41073,N_41326);
or U42390 (N_42390,N_41583,N_41771);
nand U42391 (N_42391,N_41887,N_41533);
xnor U42392 (N_42392,N_41266,N_41960);
and U42393 (N_42393,N_41030,N_41823);
nor U42394 (N_42394,N_41179,N_41439);
or U42395 (N_42395,N_41421,N_41796);
nor U42396 (N_42396,N_41403,N_41901);
xor U42397 (N_42397,N_41468,N_41389);
nand U42398 (N_42398,N_41002,N_41959);
nor U42399 (N_42399,N_41552,N_41982);
xnor U42400 (N_42400,N_41693,N_41187);
nor U42401 (N_42401,N_41831,N_41986);
nor U42402 (N_42402,N_41673,N_41204);
nor U42403 (N_42403,N_41652,N_41239);
nand U42404 (N_42404,N_41801,N_41436);
xor U42405 (N_42405,N_41511,N_41787);
nand U42406 (N_42406,N_41606,N_41023);
xnor U42407 (N_42407,N_41574,N_41677);
xnor U42408 (N_42408,N_41318,N_41086);
nor U42409 (N_42409,N_41276,N_41754);
xor U42410 (N_42410,N_41825,N_41112);
nor U42411 (N_42411,N_41292,N_41340);
or U42412 (N_42412,N_41063,N_41096);
nor U42413 (N_42413,N_41766,N_41728);
nor U42414 (N_42414,N_41526,N_41126);
or U42415 (N_42415,N_41577,N_41358);
and U42416 (N_42416,N_41904,N_41452);
nor U42417 (N_42417,N_41695,N_41778);
or U42418 (N_42418,N_41895,N_41992);
nor U42419 (N_42419,N_41143,N_41635);
or U42420 (N_42420,N_41764,N_41956);
or U42421 (N_42421,N_41198,N_41337);
nor U42422 (N_42422,N_41129,N_41499);
nand U42423 (N_42423,N_41869,N_41967);
and U42424 (N_42424,N_41634,N_41466);
or U42425 (N_42425,N_41942,N_41241);
and U42426 (N_42426,N_41417,N_41654);
nand U42427 (N_42427,N_41361,N_41587);
xor U42428 (N_42428,N_41360,N_41316);
nand U42429 (N_42429,N_41527,N_41388);
nand U42430 (N_42430,N_41114,N_41306);
xnor U42431 (N_42431,N_41848,N_41323);
or U42432 (N_42432,N_41910,N_41633);
and U42433 (N_42433,N_41478,N_41317);
nand U42434 (N_42434,N_41203,N_41843);
and U42435 (N_42435,N_41135,N_41208);
nand U42436 (N_42436,N_41429,N_41514);
nand U42437 (N_42437,N_41480,N_41017);
xnor U42438 (N_42438,N_41052,N_41481);
or U42439 (N_42439,N_41299,N_41963);
xnor U42440 (N_42440,N_41175,N_41774);
and U42441 (N_42441,N_41913,N_41312);
nor U42442 (N_42442,N_41342,N_41554);
nor U42443 (N_42443,N_41390,N_41260);
and U42444 (N_42444,N_41062,N_41665);
and U42445 (N_42445,N_41242,N_41155);
nand U42446 (N_42446,N_41431,N_41456);
and U42447 (N_42447,N_41140,N_41932);
or U42448 (N_42448,N_41828,N_41176);
nand U42449 (N_42449,N_41891,N_41369);
or U42450 (N_42450,N_41184,N_41041);
and U42451 (N_42451,N_41835,N_41908);
nor U42452 (N_42452,N_41124,N_41016);
or U42453 (N_42453,N_41152,N_41690);
and U42454 (N_42454,N_41180,N_41755);
nor U42455 (N_42455,N_41081,N_41422);
and U42456 (N_42456,N_41079,N_41404);
xor U42457 (N_42457,N_41247,N_41103);
or U42458 (N_42458,N_41209,N_41582);
xnor U42459 (N_42459,N_41569,N_41522);
and U42460 (N_42460,N_41599,N_41944);
xor U42461 (N_42461,N_41236,N_41536);
nand U42462 (N_42462,N_41449,N_41819);
nor U42463 (N_42463,N_41915,N_41836);
nand U42464 (N_42464,N_41275,N_41531);
and U42465 (N_42465,N_41057,N_41731);
and U42466 (N_42466,N_41535,N_41189);
and U42467 (N_42467,N_41881,N_41807);
and U42468 (N_42468,N_41482,N_41829);
and U42469 (N_42469,N_41280,N_41712);
nor U42470 (N_42470,N_41936,N_41447);
or U42471 (N_42471,N_41141,N_41822);
or U42472 (N_42472,N_41727,N_41210);
or U42473 (N_42473,N_41197,N_41878);
nor U42474 (N_42474,N_41115,N_41194);
xnor U42475 (N_42475,N_41585,N_41805);
and U42476 (N_42476,N_41118,N_41556);
nor U42477 (N_42477,N_41132,N_41763);
nand U42478 (N_42478,N_41734,N_41237);
xor U42479 (N_42479,N_41846,N_41884);
or U42480 (N_42480,N_41617,N_41972);
xor U42481 (N_42481,N_41170,N_41336);
xnor U42482 (N_42482,N_41048,N_41656);
nor U42483 (N_42483,N_41741,N_41167);
nor U42484 (N_42484,N_41628,N_41804);
xor U42485 (N_42485,N_41521,N_41769);
xor U42486 (N_42486,N_41719,N_41685);
nand U42487 (N_42487,N_41886,N_41021);
xnor U42488 (N_42488,N_41877,N_41636);
nand U42489 (N_42489,N_41443,N_41272);
nand U42490 (N_42490,N_41559,N_41767);
and U42491 (N_42491,N_41935,N_41069);
nor U42492 (N_42492,N_41955,N_41542);
nor U42493 (N_42493,N_41502,N_41042);
or U42494 (N_42494,N_41080,N_41044);
and U42495 (N_42495,N_41563,N_41383);
or U42496 (N_42496,N_41893,N_41516);
nand U42497 (N_42497,N_41943,N_41971);
and U42498 (N_42498,N_41759,N_41602);
nand U42499 (N_42499,N_41350,N_41399);
or U42500 (N_42500,N_41208,N_41261);
nand U42501 (N_42501,N_41478,N_41471);
xor U42502 (N_42502,N_41882,N_41061);
nor U42503 (N_42503,N_41202,N_41521);
nand U42504 (N_42504,N_41815,N_41420);
xor U42505 (N_42505,N_41354,N_41612);
or U42506 (N_42506,N_41722,N_41927);
nor U42507 (N_42507,N_41810,N_41114);
nor U42508 (N_42508,N_41721,N_41429);
nor U42509 (N_42509,N_41098,N_41577);
or U42510 (N_42510,N_41345,N_41849);
and U42511 (N_42511,N_41700,N_41888);
and U42512 (N_42512,N_41036,N_41940);
nor U42513 (N_42513,N_41610,N_41643);
nor U42514 (N_42514,N_41840,N_41355);
xor U42515 (N_42515,N_41573,N_41860);
nand U42516 (N_42516,N_41172,N_41322);
nand U42517 (N_42517,N_41963,N_41768);
and U42518 (N_42518,N_41671,N_41594);
nand U42519 (N_42519,N_41287,N_41836);
and U42520 (N_42520,N_41599,N_41857);
xnor U42521 (N_42521,N_41401,N_41150);
or U42522 (N_42522,N_41794,N_41298);
nor U42523 (N_42523,N_41654,N_41210);
and U42524 (N_42524,N_41135,N_41482);
or U42525 (N_42525,N_41967,N_41643);
and U42526 (N_42526,N_41701,N_41687);
nand U42527 (N_42527,N_41623,N_41338);
xor U42528 (N_42528,N_41815,N_41332);
nor U42529 (N_42529,N_41593,N_41451);
and U42530 (N_42530,N_41796,N_41194);
nor U42531 (N_42531,N_41743,N_41554);
nand U42532 (N_42532,N_41024,N_41039);
or U42533 (N_42533,N_41697,N_41514);
nand U42534 (N_42534,N_41063,N_41738);
nor U42535 (N_42535,N_41308,N_41548);
or U42536 (N_42536,N_41129,N_41534);
nand U42537 (N_42537,N_41748,N_41470);
nor U42538 (N_42538,N_41240,N_41581);
and U42539 (N_42539,N_41472,N_41048);
nor U42540 (N_42540,N_41060,N_41164);
and U42541 (N_42541,N_41216,N_41416);
xor U42542 (N_42542,N_41927,N_41090);
and U42543 (N_42543,N_41326,N_41570);
nand U42544 (N_42544,N_41580,N_41557);
or U42545 (N_42545,N_41944,N_41673);
and U42546 (N_42546,N_41946,N_41064);
xor U42547 (N_42547,N_41707,N_41047);
xnor U42548 (N_42548,N_41787,N_41077);
and U42549 (N_42549,N_41598,N_41532);
xnor U42550 (N_42550,N_41479,N_41748);
or U42551 (N_42551,N_41739,N_41950);
or U42552 (N_42552,N_41864,N_41053);
nor U42553 (N_42553,N_41343,N_41765);
nor U42554 (N_42554,N_41119,N_41601);
and U42555 (N_42555,N_41118,N_41570);
or U42556 (N_42556,N_41648,N_41315);
and U42557 (N_42557,N_41979,N_41487);
xor U42558 (N_42558,N_41607,N_41623);
or U42559 (N_42559,N_41186,N_41206);
or U42560 (N_42560,N_41174,N_41340);
and U42561 (N_42561,N_41871,N_41786);
xnor U42562 (N_42562,N_41724,N_41796);
or U42563 (N_42563,N_41080,N_41154);
nand U42564 (N_42564,N_41431,N_41929);
or U42565 (N_42565,N_41818,N_41034);
and U42566 (N_42566,N_41209,N_41494);
and U42567 (N_42567,N_41166,N_41029);
and U42568 (N_42568,N_41296,N_41176);
or U42569 (N_42569,N_41508,N_41242);
and U42570 (N_42570,N_41823,N_41042);
and U42571 (N_42571,N_41702,N_41225);
or U42572 (N_42572,N_41083,N_41828);
and U42573 (N_42573,N_41277,N_41512);
nand U42574 (N_42574,N_41802,N_41537);
or U42575 (N_42575,N_41119,N_41526);
xnor U42576 (N_42576,N_41546,N_41933);
nor U42577 (N_42577,N_41864,N_41150);
or U42578 (N_42578,N_41273,N_41386);
nor U42579 (N_42579,N_41126,N_41359);
nor U42580 (N_42580,N_41302,N_41958);
xor U42581 (N_42581,N_41602,N_41192);
nand U42582 (N_42582,N_41546,N_41539);
or U42583 (N_42583,N_41257,N_41504);
and U42584 (N_42584,N_41548,N_41945);
xnor U42585 (N_42585,N_41810,N_41397);
nor U42586 (N_42586,N_41143,N_41109);
nand U42587 (N_42587,N_41068,N_41140);
or U42588 (N_42588,N_41774,N_41590);
or U42589 (N_42589,N_41874,N_41062);
and U42590 (N_42590,N_41645,N_41687);
and U42591 (N_42591,N_41849,N_41578);
nor U42592 (N_42592,N_41206,N_41218);
and U42593 (N_42593,N_41670,N_41454);
nand U42594 (N_42594,N_41389,N_41981);
nand U42595 (N_42595,N_41928,N_41996);
nand U42596 (N_42596,N_41220,N_41325);
nor U42597 (N_42597,N_41664,N_41903);
nand U42598 (N_42598,N_41848,N_41235);
nand U42599 (N_42599,N_41938,N_41244);
and U42600 (N_42600,N_41429,N_41988);
nor U42601 (N_42601,N_41180,N_41865);
xor U42602 (N_42602,N_41528,N_41311);
and U42603 (N_42603,N_41521,N_41566);
and U42604 (N_42604,N_41648,N_41304);
and U42605 (N_42605,N_41222,N_41795);
xor U42606 (N_42606,N_41596,N_41442);
xnor U42607 (N_42607,N_41426,N_41705);
and U42608 (N_42608,N_41756,N_41461);
nand U42609 (N_42609,N_41499,N_41375);
nand U42610 (N_42610,N_41379,N_41212);
xor U42611 (N_42611,N_41216,N_41938);
and U42612 (N_42612,N_41169,N_41524);
nor U42613 (N_42613,N_41648,N_41051);
nand U42614 (N_42614,N_41706,N_41594);
nor U42615 (N_42615,N_41009,N_41379);
or U42616 (N_42616,N_41604,N_41440);
nor U42617 (N_42617,N_41872,N_41007);
nor U42618 (N_42618,N_41944,N_41836);
nand U42619 (N_42619,N_41654,N_41847);
and U42620 (N_42620,N_41538,N_41151);
and U42621 (N_42621,N_41984,N_41921);
xnor U42622 (N_42622,N_41004,N_41988);
nor U42623 (N_42623,N_41222,N_41793);
xnor U42624 (N_42624,N_41246,N_41481);
nor U42625 (N_42625,N_41994,N_41950);
nand U42626 (N_42626,N_41226,N_41643);
nand U42627 (N_42627,N_41505,N_41464);
or U42628 (N_42628,N_41890,N_41761);
nor U42629 (N_42629,N_41472,N_41541);
nor U42630 (N_42630,N_41014,N_41667);
or U42631 (N_42631,N_41531,N_41886);
xor U42632 (N_42632,N_41413,N_41231);
nor U42633 (N_42633,N_41260,N_41893);
nand U42634 (N_42634,N_41312,N_41180);
and U42635 (N_42635,N_41514,N_41762);
nor U42636 (N_42636,N_41735,N_41369);
nor U42637 (N_42637,N_41143,N_41953);
or U42638 (N_42638,N_41705,N_41987);
and U42639 (N_42639,N_41465,N_41963);
xor U42640 (N_42640,N_41609,N_41348);
or U42641 (N_42641,N_41492,N_41624);
or U42642 (N_42642,N_41383,N_41710);
xor U42643 (N_42643,N_41060,N_41553);
nor U42644 (N_42644,N_41210,N_41568);
or U42645 (N_42645,N_41021,N_41827);
nand U42646 (N_42646,N_41353,N_41215);
or U42647 (N_42647,N_41514,N_41836);
nand U42648 (N_42648,N_41248,N_41057);
and U42649 (N_42649,N_41721,N_41148);
and U42650 (N_42650,N_41205,N_41030);
nand U42651 (N_42651,N_41589,N_41383);
or U42652 (N_42652,N_41526,N_41106);
nand U42653 (N_42653,N_41689,N_41529);
nand U42654 (N_42654,N_41317,N_41829);
nor U42655 (N_42655,N_41906,N_41796);
xnor U42656 (N_42656,N_41585,N_41987);
and U42657 (N_42657,N_41907,N_41687);
nor U42658 (N_42658,N_41266,N_41627);
nor U42659 (N_42659,N_41953,N_41137);
or U42660 (N_42660,N_41401,N_41635);
or U42661 (N_42661,N_41454,N_41867);
nor U42662 (N_42662,N_41091,N_41202);
nor U42663 (N_42663,N_41579,N_41565);
nor U42664 (N_42664,N_41006,N_41786);
or U42665 (N_42665,N_41518,N_41051);
xnor U42666 (N_42666,N_41851,N_41686);
nand U42667 (N_42667,N_41910,N_41091);
nand U42668 (N_42668,N_41798,N_41747);
and U42669 (N_42669,N_41620,N_41767);
and U42670 (N_42670,N_41430,N_41482);
and U42671 (N_42671,N_41550,N_41503);
nor U42672 (N_42672,N_41855,N_41027);
xor U42673 (N_42673,N_41430,N_41800);
nand U42674 (N_42674,N_41789,N_41337);
nand U42675 (N_42675,N_41902,N_41499);
nand U42676 (N_42676,N_41045,N_41716);
nand U42677 (N_42677,N_41292,N_41397);
nand U42678 (N_42678,N_41821,N_41157);
xor U42679 (N_42679,N_41061,N_41565);
nor U42680 (N_42680,N_41926,N_41315);
nor U42681 (N_42681,N_41895,N_41038);
nand U42682 (N_42682,N_41296,N_41760);
or U42683 (N_42683,N_41311,N_41084);
xor U42684 (N_42684,N_41061,N_41839);
and U42685 (N_42685,N_41979,N_41960);
nor U42686 (N_42686,N_41868,N_41667);
or U42687 (N_42687,N_41128,N_41179);
xnor U42688 (N_42688,N_41475,N_41374);
nor U42689 (N_42689,N_41263,N_41932);
nand U42690 (N_42690,N_41737,N_41701);
nand U42691 (N_42691,N_41685,N_41376);
nand U42692 (N_42692,N_41600,N_41744);
or U42693 (N_42693,N_41883,N_41940);
nand U42694 (N_42694,N_41400,N_41789);
or U42695 (N_42695,N_41051,N_41412);
xnor U42696 (N_42696,N_41919,N_41646);
nand U42697 (N_42697,N_41778,N_41053);
and U42698 (N_42698,N_41249,N_41698);
and U42699 (N_42699,N_41733,N_41791);
nor U42700 (N_42700,N_41947,N_41224);
nor U42701 (N_42701,N_41955,N_41762);
nand U42702 (N_42702,N_41588,N_41976);
or U42703 (N_42703,N_41510,N_41274);
and U42704 (N_42704,N_41544,N_41407);
or U42705 (N_42705,N_41885,N_41056);
nor U42706 (N_42706,N_41654,N_41946);
and U42707 (N_42707,N_41292,N_41850);
xor U42708 (N_42708,N_41540,N_41969);
nor U42709 (N_42709,N_41678,N_41376);
or U42710 (N_42710,N_41908,N_41540);
xor U42711 (N_42711,N_41212,N_41866);
and U42712 (N_42712,N_41664,N_41347);
or U42713 (N_42713,N_41356,N_41901);
xnor U42714 (N_42714,N_41936,N_41232);
nor U42715 (N_42715,N_41124,N_41641);
and U42716 (N_42716,N_41853,N_41537);
nor U42717 (N_42717,N_41425,N_41553);
nor U42718 (N_42718,N_41270,N_41455);
and U42719 (N_42719,N_41113,N_41380);
nand U42720 (N_42720,N_41709,N_41774);
or U42721 (N_42721,N_41993,N_41581);
or U42722 (N_42722,N_41980,N_41276);
or U42723 (N_42723,N_41396,N_41062);
nor U42724 (N_42724,N_41484,N_41585);
or U42725 (N_42725,N_41806,N_41382);
nor U42726 (N_42726,N_41033,N_41448);
and U42727 (N_42727,N_41650,N_41143);
or U42728 (N_42728,N_41746,N_41957);
and U42729 (N_42729,N_41421,N_41021);
nor U42730 (N_42730,N_41101,N_41820);
and U42731 (N_42731,N_41502,N_41170);
nand U42732 (N_42732,N_41231,N_41506);
nand U42733 (N_42733,N_41017,N_41768);
nand U42734 (N_42734,N_41279,N_41211);
and U42735 (N_42735,N_41199,N_41293);
and U42736 (N_42736,N_41849,N_41271);
or U42737 (N_42737,N_41596,N_41727);
or U42738 (N_42738,N_41633,N_41411);
nor U42739 (N_42739,N_41471,N_41122);
xnor U42740 (N_42740,N_41800,N_41149);
nor U42741 (N_42741,N_41566,N_41409);
nand U42742 (N_42742,N_41369,N_41671);
nor U42743 (N_42743,N_41348,N_41610);
nand U42744 (N_42744,N_41094,N_41840);
nand U42745 (N_42745,N_41093,N_41063);
nor U42746 (N_42746,N_41361,N_41126);
nor U42747 (N_42747,N_41136,N_41984);
xor U42748 (N_42748,N_41616,N_41674);
nand U42749 (N_42749,N_41600,N_41682);
nor U42750 (N_42750,N_41859,N_41525);
nand U42751 (N_42751,N_41345,N_41315);
nand U42752 (N_42752,N_41931,N_41973);
and U42753 (N_42753,N_41460,N_41055);
or U42754 (N_42754,N_41200,N_41165);
xor U42755 (N_42755,N_41107,N_41959);
or U42756 (N_42756,N_41526,N_41831);
xor U42757 (N_42757,N_41109,N_41725);
nand U42758 (N_42758,N_41810,N_41570);
nor U42759 (N_42759,N_41046,N_41938);
or U42760 (N_42760,N_41677,N_41018);
and U42761 (N_42761,N_41526,N_41270);
xnor U42762 (N_42762,N_41286,N_41500);
nand U42763 (N_42763,N_41493,N_41376);
and U42764 (N_42764,N_41310,N_41993);
or U42765 (N_42765,N_41318,N_41548);
or U42766 (N_42766,N_41694,N_41837);
xor U42767 (N_42767,N_41365,N_41535);
and U42768 (N_42768,N_41363,N_41502);
or U42769 (N_42769,N_41951,N_41514);
nor U42770 (N_42770,N_41427,N_41859);
and U42771 (N_42771,N_41920,N_41595);
or U42772 (N_42772,N_41678,N_41212);
xor U42773 (N_42773,N_41533,N_41290);
xnor U42774 (N_42774,N_41369,N_41549);
xor U42775 (N_42775,N_41720,N_41171);
xnor U42776 (N_42776,N_41219,N_41015);
xnor U42777 (N_42777,N_41198,N_41887);
or U42778 (N_42778,N_41949,N_41883);
nand U42779 (N_42779,N_41988,N_41986);
xor U42780 (N_42780,N_41251,N_41992);
xnor U42781 (N_42781,N_41017,N_41802);
and U42782 (N_42782,N_41316,N_41378);
nand U42783 (N_42783,N_41255,N_41613);
or U42784 (N_42784,N_41229,N_41688);
or U42785 (N_42785,N_41932,N_41321);
and U42786 (N_42786,N_41193,N_41886);
xnor U42787 (N_42787,N_41639,N_41612);
or U42788 (N_42788,N_41845,N_41865);
or U42789 (N_42789,N_41531,N_41836);
nor U42790 (N_42790,N_41307,N_41184);
nor U42791 (N_42791,N_41205,N_41719);
and U42792 (N_42792,N_41829,N_41600);
nand U42793 (N_42793,N_41607,N_41532);
and U42794 (N_42794,N_41139,N_41605);
nor U42795 (N_42795,N_41378,N_41345);
or U42796 (N_42796,N_41464,N_41121);
and U42797 (N_42797,N_41404,N_41297);
nand U42798 (N_42798,N_41632,N_41537);
and U42799 (N_42799,N_41977,N_41904);
or U42800 (N_42800,N_41107,N_41280);
nor U42801 (N_42801,N_41224,N_41423);
nor U42802 (N_42802,N_41912,N_41206);
nor U42803 (N_42803,N_41383,N_41411);
nand U42804 (N_42804,N_41755,N_41009);
xor U42805 (N_42805,N_41770,N_41172);
and U42806 (N_42806,N_41657,N_41009);
and U42807 (N_42807,N_41543,N_41884);
and U42808 (N_42808,N_41960,N_41809);
nand U42809 (N_42809,N_41908,N_41358);
xor U42810 (N_42810,N_41705,N_41928);
nand U42811 (N_42811,N_41212,N_41231);
nor U42812 (N_42812,N_41796,N_41461);
and U42813 (N_42813,N_41458,N_41359);
nor U42814 (N_42814,N_41358,N_41419);
and U42815 (N_42815,N_41485,N_41869);
nand U42816 (N_42816,N_41747,N_41398);
and U42817 (N_42817,N_41389,N_41707);
nand U42818 (N_42818,N_41990,N_41629);
nand U42819 (N_42819,N_41935,N_41668);
and U42820 (N_42820,N_41246,N_41713);
xnor U42821 (N_42821,N_41273,N_41463);
nand U42822 (N_42822,N_41381,N_41138);
and U42823 (N_42823,N_41937,N_41550);
or U42824 (N_42824,N_41026,N_41749);
and U42825 (N_42825,N_41632,N_41458);
or U42826 (N_42826,N_41463,N_41660);
or U42827 (N_42827,N_41451,N_41083);
or U42828 (N_42828,N_41882,N_41426);
xor U42829 (N_42829,N_41287,N_41094);
or U42830 (N_42830,N_41467,N_41753);
nor U42831 (N_42831,N_41839,N_41467);
nand U42832 (N_42832,N_41998,N_41417);
and U42833 (N_42833,N_41735,N_41312);
and U42834 (N_42834,N_41480,N_41140);
nor U42835 (N_42835,N_41994,N_41322);
nand U42836 (N_42836,N_41253,N_41100);
nor U42837 (N_42837,N_41654,N_41694);
nand U42838 (N_42838,N_41177,N_41695);
and U42839 (N_42839,N_41979,N_41827);
or U42840 (N_42840,N_41639,N_41277);
xor U42841 (N_42841,N_41324,N_41974);
or U42842 (N_42842,N_41279,N_41462);
or U42843 (N_42843,N_41750,N_41978);
nand U42844 (N_42844,N_41526,N_41163);
nor U42845 (N_42845,N_41085,N_41241);
xor U42846 (N_42846,N_41242,N_41184);
nor U42847 (N_42847,N_41400,N_41195);
xnor U42848 (N_42848,N_41225,N_41285);
nand U42849 (N_42849,N_41473,N_41231);
nand U42850 (N_42850,N_41233,N_41527);
and U42851 (N_42851,N_41679,N_41589);
nand U42852 (N_42852,N_41682,N_41411);
nor U42853 (N_42853,N_41595,N_41035);
and U42854 (N_42854,N_41632,N_41820);
or U42855 (N_42855,N_41553,N_41448);
xnor U42856 (N_42856,N_41740,N_41074);
or U42857 (N_42857,N_41741,N_41170);
nor U42858 (N_42858,N_41299,N_41000);
nand U42859 (N_42859,N_41692,N_41568);
and U42860 (N_42860,N_41284,N_41142);
nor U42861 (N_42861,N_41770,N_41420);
nand U42862 (N_42862,N_41885,N_41639);
or U42863 (N_42863,N_41616,N_41539);
nand U42864 (N_42864,N_41016,N_41510);
nand U42865 (N_42865,N_41221,N_41924);
xnor U42866 (N_42866,N_41750,N_41614);
or U42867 (N_42867,N_41907,N_41417);
and U42868 (N_42868,N_41283,N_41899);
xnor U42869 (N_42869,N_41355,N_41136);
nand U42870 (N_42870,N_41708,N_41649);
and U42871 (N_42871,N_41937,N_41435);
and U42872 (N_42872,N_41726,N_41460);
and U42873 (N_42873,N_41531,N_41530);
xor U42874 (N_42874,N_41151,N_41169);
xor U42875 (N_42875,N_41156,N_41020);
and U42876 (N_42876,N_41351,N_41296);
nor U42877 (N_42877,N_41162,N_41606);
or U42878 (N_42878,N_41473,N_41585);
nor U42879 (N_42879,N_41140,N_41239);
nand U42880 (N_42880,N_41702,N_41963);
nand U42881 (N_42881,N_41211,N_41626);
nand U42882 (N_42882,N_41042,N_41690);
nor U42883 (N_42883,N_41882,N_41317);
or U42884 (N_42884,N_41735,N_41424);
or U42885 (N_42885,N_41705,N_41154);
nand U42886 (N_42886,N_41159,N_41652);
and U42887 (N_42887,N_41633,N_41611);
xnor U42888 (N_42888,N_41395,N_41145);
nand U42889 (N_42889,N_41023,N_41864);
nor U42890 (N_42890,N_41855,N_41956);
nand U42891 (N_42891,N_41570,N_41215);
or U42892 (N_42892,N_41954,N_41740);
or U42893 (N_42893,N_41235,N_41530);
nor U42894 (N_42894,N_41163,N_41049);
nor U42895 (N_42895,N_41799,N_41406);
nor U42896 (N_42896,N_41867,N_41296);
xor U42897 (N_42897,N_41367,N_41215);
nor U42898 (N_42898,N_41190,N_41245);
nand U42899 (N_42899,N_41379,N_41629);
xnor U42900 (N_42900,N_41249,N_41399);
xnor U42901 (N_42901,N_41554,N_41106);
nand U42902 (N_42902,N_41979,N_41574);
xnor U42903 (N_42903,N_41539,N_41871);
and U42904 (N_42904,N_41764,N_41390);
nand U42905 (N_42905,N_41449,N_41808);
nor U42906 (N_42906,N_41794,N_41819);
and U42907 (N_42907,N_41665,N_41049);
nand U42908 (N_42908,N_41575,N_41307);
nand U42909 (N_42909,N_41854,N_41527);
nand U42910 (N_42910,N_41155,N_41704);
nand U42911 (N_42911,N_41958,N_41865);
or U42912 (N_42912,N_41828,N_41248);
xor U42913 (N_42913,N_41483,N_41815);
and U42914 (N_42914,N_41465,N_41958);
or U42915 (N_42915,N_41819,N_41458);
nor U42916 (N_42916,N_41089,N_41314);
or U42917 (N_42917,N_41556,N_41474);
nand U42918 (N_42918,N_41484,N_41676);
nor U42919 (N_42919,N_41946,N_41012);
nor U42920 (N_42920,N_41911,N_41442);
and U42921 (N_42921,N_41002,N_41442);
nand U42922 (N_42922,N_41440,N_41409);
nor U42923 (N_42923,N_41325,N_41968);
nor U42924 (N_42924,N_41009,N_41142);
and U42925 (N_42925,N_41715,N_41987);
xor U42926 (N_42926,N_41570,N_41572);
xor U42927 (N_42927,N_41067,N_41501);
nor U42928 (N_42928,N_41513,N_41022);
and U42929 (N_42929,N_41540,N_41500);
and U42930 (N_42930,N_41056,N_41988);
or U42931 (N_42931,N_41446,N_41870);
xor U42932 (N_42932,N_41965,N_41419);
nor U42933 (N_42933,N_41128,N_41320);
nor U42934 (N_42934,N_41811,N_41039);
and U42935 (N_42935,N_41998,N_41398);
nor U42936 (N_42936,N_41187,N_41886);
and U42937 (N_42937,N_41463,N_41365);
and U42938 (N_42938,N_41924,N_41762);
nand U42939 (N_42939,N_41015,N_41880);
or U42940 (N_42940,N_41379,N_41051);
and U42941 (N_42941,N_41943,N_41785);
xnor U42942 (N_42942,N_41840,N_41233);
nand U42943 (N_42943,N_41689,N_41800);
nor U42944 (N_42944,N_41757,N_41335);
nand U42945 (N_42945,N_41520,N_41397);
or U42946 (N_42946,N_41436,N_41586);
nand U42947 (N_42947,N_41166,N_41498);
or U42948 (N_42948,N_41586,N_41334);
nor U42949 (N_42949,N_41407,N_41241);
nand U42950 (N_42950,N_41078,N_41278);
and U42951 (N_42951,N_41961,N_41933);
and U42952 (N_42952,N_41616,N_41499);
nor U42953 (N_42953,N_41171,N_41799);
nor U42954 (N_42954,N_41659,N_41450);
or U42955 (N_42955,N_41807,N_41078);
xor U42956 (N_42956,N_41080,N_41739);
and U42957 (N_42957,N_41523,N_41683);
xnor U42958 (N_42958,N_41384,N_41726);
nor U42959 (N_42959,N_41088,N_41842);
nor U42960 (N_42960,N_41491,N_41641);
or U42961 (N_42961,N_41275,N_41638);
nand U42962 (N_42962,N_41572,N_41869);
nor U42963 (N_42963,N_41854,N_41725);
nand U42964 (N_42964,N_41091,N_41195);
nand U42965 (N_42965,N_41623,N_41276);
nor U42966 (N_42966,N_41591,N_41867);
nand U42967 (N_42967,N_41279,N_41333);
nor U42968 (N_42968,N_41619,N_41849);
and U42969 (N_42969,N_41612,N_41245);
nor U42970 (N_42970,N_41368,N_41130);
nand U42971 (N_42971,N_41499,N_41510);
or U42972 (N_42972,N_41413,N_41474);
and U42973 (N_42973,N_41157,N_41271);
or U42974 (N_42974,N_41320,N_41941);
xor U42975 (N_42975,N_41653,N_41047);
xor U42976 (N_42976,N_41720,N_41922);
or U42977 (N_42977,N_41807,N_41086);
nand U42978 (N_42978,N_41796,N_41292);
and U42979 (N_42979,N_41720,N_41489);
xnor U42980 (N_42980,N_41861,N_41761);
xor U42981 (N_42981,N_41391,N_41268);
and U42982 (N_42982,N_41156,N_41957);
nor U42983 (N_42983,N_41717,N_41787);
or U42984 (N_42984,N_41587,N_41117);
and U42985 (N_42985,N_41937,N_41562);
nor U42986 (N_42986,N_41154,N_41964);
nand U42987 (N_42987,N_41316,N_41069);
nand U42988 (N_42988,N_41031,N_41630);
nor U42989 (N_42989,N_41662,N_41566);
xnor U42990 (N_42990,N_41039,N_41841);
xnor U42991 (N_42991,N_41861,N_41014);
nand U42992 (N_42992,N_41329,N_41121);
and U42993 (N_42993,N_41564,N_41013);
and U42994 (N_42994,N_41978,N_41618);
or U42995 (N_42995,N_41417,N_41238);
nor U42996 (N_42996,N_41907,N_41770);
xor U42997 (N_42997,N_41797,N_41318);
or U42998 (N_42998,N_41905,N_41495);
xor U42999 (N_42999,N_41503,N_41238);
xnor U43000 (N_43000,N_42991,N_42511);
xnor U43001 (N_43001,N_42782,N_42618);
nand U43002 (N_43002,N_42937,N_42243);
nand U43003 (N_43003,N_42377,N_42220);
nand U43004 (N_43004,N_42234,N_42283);
xnor U43005 (N_43005,N_42195,N_42731);
xor U43006 (N_43006,N_42209,N_42280);
or U43007 (N_43007,N_42560,N_42240);
nand U43008 (N_43008,N_42964,N_42295);
nand U43009 (N_43009,N_42325,N_42299);
nor U43010 (N_43010,N_42259,N_42881);
nor U43011 (N_43011,N_42851,N_42887);
nand U43012 (N_43012,N_42126,N_42013);
nand U43013 (N_43013,N_42582,N_42168);
and U43014 (N_43014,N_42064,N_42077);
nor U43015 (N_43015,N_42167,N_42203);
or U43016 (N_43016,N_42027,N_42806);
nand U43017 (N_43017,N_42300,N_42440);
nand U43018 (N_43018,N_42892,N_42778);
xnor U43019 (N_43019,N_42011,N_42174);
or U43020 (N_43020,N_42565,N_42643);
nor U43021 (N_43021,N_42095,N_42099);
nor U43022 (N_43022,N_42375,N_42917);
and U43023 (N_43023,N_42397,N_42951);
xnor U43024 (N_43024,N_42499,N_42121);
xor U43025 (N_43025,N_42670,N_42091);
nand U43026 (N_43026,N_42256,N_42587);
and U43027 (N_43027,N_42182,N_42469);
xnor U43028 (N_43028,N_42625,N_42430);
and U43029 (N_43029,N_42960,N_42974);
xnor U43030 (N_43030,N_42047,N_42854);
and U43031 (N_43031,N_42287,N_42745);
nand U43032 (N_43032,N_42542,N_42196);
nand U43033 (N_43033,N_42119,N_42610);
nor U43034 (N_43034,N_42482,N_42976);
nor U43035 (N_43035,N_42679,N_42031);
nor U43036 (N_43036,N_42012,N_42207);
nor U43037 (N_43037,N_42811,N_42659);
nor U43038 (N_43038,N_42489,N_42224);
xnor U43039 (N_43039,N_42647,N_42003);
nor U43040 (N_43040,N_42836,N_42092);
or U43041 (N_43041,N_42605,N_42164);
and U43042 (N_43042,N_42428,N_42925);
xnor U43043 (N_43043,N_42060,N_42436);
and U43044 (N_43044,N_42297,N_42787);
nor U43045 (N_43045,N_42835,N_42671);
and U43046 (N_43046,N_42304,N_42065);
and U43047 (N_43047,N_42066,N_42739);
or U43048 (N_43048,N_42666,N_42800);
nor U43049 (N_43049,N_42104,N_42574);
or U43050 (N_43050,N_42896,N_42205);
nand U43051 (N_43051,N_42379,N_42691);
xnor U43052 (N_43052,N_42869,N_42050);
xnor U43053 (N_43053,N_42773,N_42563);
and U43054 (N_43054,N_42187,N_42973);
nor U43055 (N_43055,N_42460,N_42353);
nand U43056 (N_43056,N_42197,N_42312);
and U43057 (N_43057,N_42264,N_42798);
xor U43058 (N_43058,N_42999,N_42633);
nor U43059 (N_43059,N_42829,N_42926);
or U43060 (N_43060,N_42330,N_42697);
and U43061 (N_43061,N_42507,N_42941);
nand U43062 (N_43062,N_42635,N_42178);
xnor U43063 (N_43063,N_42970,N_42402);
nor U43064 (N_43064,N_42388,N_42867);
and U43065 (N_43065,N_42438,N_42876);
xnor U43066 (N_43066,N_42911,N_42909);
nor U43067 (N_43067,N_42160,N_42437);
nor U43068 (N_43068,N_42907,N_42626);
xnor U43069 (N_43069,N_42728,N_42744);
nand U43070 (N_43070,N_42023,N_42741);
nor U43071 (N_43071,N_42831,N_42719);
xnor U43072 (N_43072,N_42071,N_42809);
and U43073 (N_43073,N_42766,N_42609);
nand U43074 (N_43074,N_42906,N_42446);
nand U43075 (N_43075,N_42544,N_42775);
xor U43076 (N_43076,N_42162,N_42759);
and U43077 (N_43077,N_42624,N_42943);
xnor U43078 (N_43078,N_42962,N_42746);
or U43079 (N_43079,N_42850,N_42206);
or U43080 (N_43080,N_42229,N_42687);
or U43081 (N_43081,N_42017,N_42459);
or U43082 (N_43082,N_42275,N_42036);
nor U43083 (N_43083,N_42096,N_42281);
or U43084 (N_43084,N_42333,N_42956);
or U43085 (N_43085,N_42871,N_42571);
and U43086 (N_43086,N_42562,N_42588);
xnor U43087 (N_43087,N_42793,N_42005);
nor U43088 (N_43088,N_42302,N_42359);
xnor U43089 (N_43089,N_42703,N_42265);
and U43090 (N_43090,N_42914,N_42037);
or U43091 (N_43091,N_42903,N_42001);
and U43092 (N_43092,N_42645,N_42435);
or U43093 (N_43093,N_42858,N_42891);
and U43094 (N_43094,N_42286,N_42044);
nand U43095 (N_43095,N_42673,N_42586);
or U43096 (N_43096,N_42212,N_42824);
xnor U43097 (N_43097,N_42874,N_42848);
nor U43098 (N_43098,N_42081,N_42232);
nor U43099 (N_43099,N_42805,N_42955);
nor U43100 (N_43100,N_42796,N_42054);
nand U43101 (N_43101,N_42058,N_42268);
nor U43102 (N_43102,N_42525,N_42656);
and U43103 (N_43103,N_42138,N_42153);
or U43104 (N_43104,N_42642,N_42086);
or U43105 (N_43105,N_42788,N_42384);
nor U43106 (N_43106,N_42750,N_42678);
or U43107 (N_43107,N_42710,N_42140);
nand U43108 (N_43108,N_42009,N_42341);
or U43109 (N_43109,N_42331,N_42596);
or U43110 (N_43110,N_42204,N_42238);
nand U43111 (N_43111,N_42087,N_42391);
nor U43112 (N_43112,N_42332,N_42818);
and U43113 (N_43113,N_42905,N_42339);
or U43114 (N_43114,N_42429,N_42315);
xor U43115 (N_43115,N_42105,N_42134);
nand U43116 (N_43116,N_42935,N_42218);
or U43117 (N_43117,N_42704,N_42423);
xor U43118 (N_43118,N_42418,N_42637);
nand U43119 (N_43119,N_42768,N_42825);
nor U43120 (N_43120,N_42715,N_42764);
and U43121 (N_43121,N_42948,N_42466);
and U43122 (N_43122,N_42493,N_42727);
nand U43123 (N_43123,N_42677,N_42711);
xor U43124 (N_43124,N_42405,N_42846);
nand U43125 (N_43125,N_42125,N_42172);
or U43126 (N_43126,N_42815,N_42473);
nor U43127 (N_43127,N_42792,N_42510);
and U43128 (N_43128,N_42061,N_42324);
nand U43129 (N_43129,N_42082,N_42426);
nor U43130 (N_43130,N_42897,N_42658);
xnor U43131 (N_43131,N_42838,N_42602);
and U43132 (N_43132,N_42570,N_42171);
nor U43133 (N_43133,N_42080,N_42404);
nand U43134 (N_43134,N_42409,N_42864);
or U43135 (N_43135,N_42621,N_42709);
nor U43136 (N_43136,N_42736,N_42734);
nor U43137 (N_43137,N_42141,N_42549);
nand U43138 (N_43138,N_42382,N_42120);
nor U43139 (N_43139,N_42564,N_42018);
nand U43140 (N_43140,N_42415,N_42840);
nor U43141 (N_43141,N_42878,N_42716);
nand U43142 (N_43142,N_42479,N_42362);
nor U43143 (N_43143,N_42879,N_42754);
and U43144 (N_43144,N_42462,N_42335);
nand U43145 (N_43145,N_42505,N_42363);
and U43146 (N_43146,N_42398,N_42260);
xnor U43147 (N_43147,N_42093,N_42975);
nand U43148 (N_43148,N_42393,N_42639);
nand U43149 (N_43149,N_42580,N_42445);
and U43150 (N_43150,N_42347,N_42987);
or U43151 (N_43151,N_42180,N_42070);
nor U43152 (N_43152,N_42231,N_42958);
nand U43153 (N_43153,N_42296,N_42517);
and U43154 (N_43154,N_42386,N_42684);
nand U43155 (N_43155,N_42444,N_42557);
or U43156 (N_43156,N_42827,N_42599);
xor U43157 (N_43157,N_42771,N_42233);
nand U43158 (N_43158,N_42757,N_42597);
nor U43159 (N_43159,N_42088,N_42441);
nor U43160 (N_43160,N_42271,N_42947);
nor U43161 (N_43161,N_42250,N_42097);
xor U43162 (N_43162,N_42860,N_42360);
nand U43163 (N_43163,N_42868,N_42450);
nor U43164 (N_43164,N_42569,N_42993);
or U43165 (N_43165,N_42039,N_42213);
nor U43166 (N_43166,N_42048,N_42720);
xor U43167 (N_43167,N_42992,N_42219);
or U43168 (N_43168,N_42116,N_42957);
and U43169 (N_43169,N_42807,N_42814);
nand U43170 (N_43170,N_42900,N_42594);
nand U43171 (N_43171,N_42242,N_42554);
xnor U43172 (N_43172,N_42561,N_42702);
xnor U43173 (N_43173,N_42284,N_42100);
nand U43174 (N_43174,N_42340,N_42261);
and U43175 (N_43175,N_42543,N_42216);
and U43176 (N_43176,N_42593,N_42150);
xor U43177 (N_43177,N_42506,N_42263);
and U43178 (N_43178,N_42713,N_42163);
and U43179 (N_43179,N_42314,N_42457);
xor U43180 (N_43180,N_42726,N_42107);
nand U43181 (N_43181,N_42414,N_42653);
nand U43182 (N_43182,N_42584,N_42244);
xor U43183 (N_43183,N_42456,N_42545);
and U43184 (N_43184,N_42193,N_42354);
and U43185 (N_43185,N_42343,N_42668);
or U43186 (N_43186,N_42342,N_42098);
or U43187 (N_43187,N_42733,N_42274);
xor U43188 (N_43188,N_42756,N_42553);
xor U43189 (N_43189,N_42801,N_42620);
nand U43190 (N_43190,N_42131,N_42755);
xnor U43191 (N_43191,N_42115,N_42680);
or U43192 (N_43192,N_42084,N_42952);
xor U43193 (N_43193,N_42412,N_42063);
or U43194 (N_43194,N_42108,N_42940);
xnor U43195 (N_43195,N_42861,N_42551);
or U43196 (N_43196,N_42660,N_42883);
xor U43197 (N_43197,N_42963,N_42655);
nor U43198 (N_43198,N_42784,N_42454);
or U43199 (N_43199,N_42059,N_42177);
nand U43200 (N_43200,N_42262,N_42309);
or U43201 (N_43201,N_42932,N_42913);
or U43202 (N_43202,N_42581,N_42616);
xnor U43203 (N_43203,N_42631,N_42146);
nand U43204 (N_43204,N_42008,N_42722);
and U43205 (N_43205,N_42531,N_42029);
xnor U43206 (N_43206,N_42695,N_42051);
nand U43207 (N_43207,N_42552,N_42458);
xor U43208 (N_43208,N_42636,N_42361);
nor U43209 (N_43209,N_42664,N_42159);
xnor U43210 (N_43210,N_42950,N_42550);
nor U43211 (N_43211,N_42161,N_42083);
and U43212 (N_43212,N_42303,N_42403);
or U43213 (N_43213,N_42431,N_42420);
nor U43214 (N_43214,N_42498,N_42488);
xor U43215 (N_43215,N_42028,N_42690);
and U43216 (N_43216,N_42394,N_42035);
nor U43217 (N_43217,N_42470,N_42191);
nand U43218 (N_43218,N_42843,N_42133);
and U43219 (N_43219,N_42762,N_42477);
and U43220 (N_43220,N_42129,N_42777);
nor U43221 (N_43221,N_42650,N_42184);
or U43222 (N_43222,N_42540,N_42681);
and U43223 (N_43223,N_42765,N_42345);
nor U43224 (N_43224,N_42122,N_42327);
nor U43225 (N_43225,N_42629,N_42045);
and U43226 (N_43226,N_42533,N_42578);
xor U43227 (N_43227,N_42516,N_42990);
and U43228 (N_43228,N_42057,N_42346);
xnor U43229 (N_43229,N_42451,N_42961);
and U43230 (N_43230,N_42127,N_42984);
xor U43231 (N_43231,N_42856,N_42705);
and U43232 (N_43232,N_42541,N_42165);
or U43233 (N_43233,N_42790,N_42500);
nor U43234 (N_43234,N_42369,N_42701);
nor U43235 (N_43235,N_42461,N_42310);
nor U43236 (N_43236,N_42410,N_42364);
and U43237 (N_43237,N_42714,N_42248);
and U43238 (N_43238,N_42374,N_42538);
or U43239 (N_43239,N_42419,N_42567);
xor U43240 (N_43240,N_42944,N_42712);
nor U43241 (N_43241,N_42024,N_42311);
nand U43242 (N_43242,N_42763,N_42052);
nand U43243 (N_43243,N_42575,N_42251);
nor U43244 (N_43244,N_42724,N_42774);
nand U43245 (N_43245,N_42613,N_42355);
and U43246 (N_43246,N_42021,N_42920);
or U43247 (N_43247,N_42067,N_42845);
nor U43248 (N_43248,N_42615,N_42492);
or U43249 (N_43249,N_42483,N_42137);
and U43250 (N_43250,N_42502,N_42079);
xnor U43251 (N_43251,N_42781,N_42949);
and U43252 (N_43252,N_42202,N_42416);
or U43253 (N_43253,N_42109,N_42748);
nand U43254 (N_43254,N_42534,N_42239);
xor U43255 (N_43255,N_42320,N_42779);
nand U43256 (N_43256,N_42020,N_42548);
and U43257 (N_43257,N_42982,N_42504);
or U43258 (N_43258,N_42558,N_42870);
or U43259 (N_43259,N_42852,N_42676);
nor U43260 (N_43260,N_42532,N_42152);
nor U43261 (N_43261,N_42795,N_42055);
and U43262 (N_43262,N_42518,N_42916);
xor U43263 (N_43263,N_42857,N_42539);
and U43264 (N_43264,N_42901,N_42010);
xnor U43265 (N_43265,N_42767,N_42863);
nor U43266 (N_43266,N_42559,N_42740);
or U43267 (N_43267,N_42529,N_42931);
nor U43268 (N_43268,N_42002,N_42812);
nand U43269 (N_43269,N_42885,N_42923);
or U43270 (N_43270,N_42572,N_42652);
nand U43271 (N_43271,N_42124,N_42761);
nand U43272 (N_43272,N_42252,N_42979);
nor U43273 (N_43273,N_42608,N_42199);
or U43274 (N_43274,N_42322,N_42865);
xnor U43275 (N_43275,N_42844,N_42110);
nand U43276 (N_43276,N_42368,N_42536);
or U43277 (N_43277,N_42972,N_42614);
or U43278 (N_43278,N_42378,N_42237);
nor U43279 (N_43279,N_42693,N_42520);
and U43280 (N_43280,N_42641,N_42953);
xor U43281 (N_43281,N_42481,N_42210);
or U43282 (N_43282,N_42228,N_42357);
xor U43283 (N_43283,N_42434,N_42908);
or U43284 (N_43284,N_42247,N_42094);
nand U43285 (N_43285,N_42804,N_42370);
and U43286 (N_43286,N_42566,N_42634);
nor U43287 (N_43287,N_42185,N_42669);
or U43288 (N_43288,N_42223,N_42279);
or U43289 (N_43289,N_42258,N_42601);
or U43290 (N_43290,N_42758,N_42025);
xnor U43291 (N_43291,N_42503,N_42604);
nand U43292 (N_43292,N_42585,N_42433);
or U43293 (N_43293,N_42826,N_42753);
and U43294 (N_43294,N_42123,N_42285);
and U43295 (N_43295,N_42442,N_42186);
xnor U43296 (N_43296,N_42139,N_42521);
nand U43297 (N_43297,N_42674,N_42336);
nand U43298 (N_43298,N_42524,N_42849);
nand U43299 (N_43299,N_42254,N_42611);
nor U43300 (N_43300,N_42476,N_42074);
and U43301 (N_43301,N_42888,N_42474);
nor U43302 (N_43302,N_42439,N_42073);
xor U43303 (N_43303,N_42241,N_42683);
or U43304 (N_43304,N_42455,N_42808);
nor U43305 (N_43305,N_42249,N_42372);
nand U43306 (N_43306,N_42292,N_42934);
nand U43307 (N_43307,N_42376,N_42270);
and U43308 (N_43308,N_42222,N_42515);
nor U43309 (N_43309,N_42698,N_42034);
and U43310 (N_43310,N_42986,N_42194);
nand U43311 (N_43311,N_42688,N_42007);
nor U43312 (N_43312,N_42118,N_42049);
and U43313 (N_43313,N_42657,N_42735);
and U43314 (N_43314,N_42143,N_42371);
nand U43315 (N_43315,N_42032,N_42873);
nand U43316 (N_43316,N_42910,N_42978);
nand U43317 (N_43317,N_42291,N_42579);
nand U43318 (N_43318,N_42344,N_42519);
or U43319 (N_43319,N_42158,N_42022);
nand U43320 (N_43320,N_42568,N_42667);
nor U43321 (N_43321,N_42069,N_42928);
xor U43322 (N_43322,N_42915,N_42718);
and U43323 (N_43323,N_42307,N_42495);
xnor U43324 (N_43324,N_42833,N_42030);
or U43325 (N_43325,N_42090,N_42425);
nor U43326 (N_43326,N_42780,N_42592);
nor U43327 (N_43327,N_42350,N_42358);
nand U43328 (N_43328,N_42769,N_42338);
xnor U43329 (N_43329,N_42497,N_42789);
and U43330 (N_43330,N_42475,N_42954);
xor U43331 (N_43331,N_42166,N_42623);
nor U43332 (N_43332,N_42465,N_42337);
and U43333 (N_43333,N_42988,N_42149);
or U43334 (N_43334,N_42352,N_42245);
nand U43335 (N_43335,N_42294,N_42959);
and U43336 (N_43336,N_42041,N_42810);
or U43337 (N_43337,N_42484,N_42272);
xor U43338 (N_43338,N_42921,N_42135);
nor U43339 (N_43339,N_42535,N_42799);
and U43340 (N_43340,N_42828,N_42214);
or U43341 (N_43341,N_42390,N_42282);
and U43342 (N_43342,N_42969,N_42000);
xor U43343 (N_43343,N_42649,N_42875);
xnor U43344 (N_43344,N_42929,N_42351);
and U43345 (N_43345,N_42820,N_42772);
or U43346 (N_43346,N_42062,N_42076);
xnor U43347 (N_43347,N_42221,N_42606);
nor U43348 (N_43348,N_42967,N_42743);
nand U43349 (N_43349,N_42924,N_42834);
and U43350 (N_43350,N_42452,N_42101);
xor U43351 (N_43351,N_42556,N_42253);
xnor U43352 (N_43352,N_42385,N_42033);
xor U43353 (N_43353,N_42752,N_42514);
xor U43354 (N_43354,N_42751,N_42513);
and U43355 (N_43355,N_42276,N_42144);
nor U43356 (N_43356,N_42487,N_42406);
xnor U43357 (N_43357,N_42323,N_42760);
xnor U43358 (N_43358,N_42813,N_42496);
nor U43359 (N_43359,N_42103,N_42842);
nand U43360 (N_43360,N_42038,N_42046);
and U43361 (N_43361,N_42056,N_42392);
or U43362 (N_43362,N_42316,N_42890);
or U43363 (N_43363,N_42837,N_42367);
and U43364 (N_43364,N_42053,N_42266);
nand U43365 (N_43365,N_42179,N_42102);
xor U43366 (N_43366,N_42732,N_42821);
nor U43367 (N_43367,N_42306,N_42675);
and U43368 (N_43368,N_42822,N_42922);
and U43369 (N_43369,N_42682,N_42638);
nand U43370 (N_43370,N_42654,N_42942);
nor U43371 (N_43371,N_42816,N_42630);
nor U43372 (N_43372,N_42288,N_42946);
nor U43373 (N_43373,N_42839,N_42464);
nand U43374 (N_43374,N_42523,N_42277);
xnor U43375 (N_43375,N_42068,N_42449);
or U43376 (N_43376,N_42349,N_42236);
or U43377 (N_43377,N_42471,N_42298);
or U43378 (N_43378,N_42694,N_42175);
nand U43379 (N_43379,N_42902,N_42662);
nand U43380 (N_43380,N_42200,N_42128);
and U43381 (N_43381,N_42501,N_42111);
and U43382 (N_43382,N_42389,N_42114);
or U43383 (N_43383,N_42226,N_42453);
xor U43384 (N_43384,N_42188,N_42113);
or U43385 (N_43385,N_42147,N_42075);
nor U43386 (N_43386,N_42154,N_42872);
nand U43387 (N_43387,N_42290,N_42919);
nor U43388 (N_43388,N_42965,N_42512);
and U43389 (N_43389,N_42877,N_42201);
nand U43390 (N_43390,N_42490,N_42491);
nand U43391 (N_43391,N_42886,N_42417);
or U43392 (N_43392,N_42526,N_42904);
nor U43393 (N_43393,N_42015,N_42257);
or U43394 (N_43394,N_42130,N_42617);
nand U43395 (N_43395,N_42721,N_42313);
nor U43396 (N_43396,N_42725,N_42447);
or U43397 (N_43397,N_42547,N_42400);
nand U43398 (N_43398,N_42014,N_42893);
nor U43399 (N_43399,N_42480,N_42573);
nor U43400 (N_43400,N_42467,N_42591);
nand U43401 (N_43401,N_42797,N_42089);
xor U43402 (N_43402,N_42387,N_42329);
or U43403 (N_43403,N_42170,N_42855);
nand U43404 (N_43404,N_42486,N_42365);
and U43405 (N_43405,N_42770,N_42040);
nor U43406 (N_43406,N_42468,N_42427);
nand U43407 (N_43407,N_42472,N_42706);
and U43408 (N_43408,N_42819,N_42269);
nand U43409 (N_43409,N_42401,N_42648);
xor U43410 (N_43410,N_42508,N_42866);
nand U43411 (N_43411,N_42632,N_42072);
xnor U43412 (N_43412,N_42590,N_42612);
xor U43413 (N_43413,N_42527,N_42004);
nand U43414 (N_43414,N_42918,N_42145);
nor U43415 (N_43415,N_42841,N_42348);
nor U43416 (N_43416,N_42085,N_42463);
or U43417 (N_43417,N_42151,N_42696);
or U43418 (N_43418,N_42043,N_42157);
or U43419 (N_43419,N_42577,N_42407);
xor U43420 (N_43420,N_42644,N_42318);
nor U43421 (N_43421,N_42791,N_42383);
and U43422 (N_43422,N_42156,N_42169);
nor U43423 (N_43423,N_42607,N_42555);
nand U43424 (N_43424,N_42832,N_42522);
nand U43425 (N_43425,N_42699,N_42106);
and U43426 (N_43426,N_42155,N_42853);
nor U43427 (N_43427,N_42685,N_42132);
or U43428 (N_43428,N_42308,N_42176);
and U43429 (N_43429,N_42981,N_42830);
xor U43430 (N_43430,N_42847,N_42528);
xnor U43431 (N_43431,N_42912,N_42600);
xnor U43432 (N_43432,N_42708,N_42619);
nand U43433 (N_43433,N_42136,N_42305);
or U43434 (N_43434,N_42859,N_42183);
nor U43435 (N_43435,N_42142,N_42794);
and U43436 (N_43436,N_42783,N_42293);
or U43437 (N_43437,N_42189,N_42895);
xnor U43438 (N_43438,N_42509,N_42945);
nand U43439 (N_43439,N_42665,N_42019);
nor U43440 (N_43440,N_42273,N_42742);
or U43441 (N_43441,N_42889,N_42971);
xnor U43442 (N_43442,N_42933,N_42977);
xnor U43443 (N_43443,N_42983,N_42267);
or U43444 (N_43444,N_42016,N_42968);
or U43445 (N_43445,N_42192,N_42823);
nand U43446 (N_43446,N_42598,N_42989);
and U43447 (N_43447,N_42537,N_42686);
nor U43448 (N_43448,N_42737,N_42939);
nand U43449 (N_43449,N_42700,N_42026);
nand U43450 (N_43450,N_42786,N_42930);
nor U43451 (N_43451,N_42651,N_42227);
or U43452 (N_43452,N_42747,N_42663);
nor U43453 (N_43453,N_42628,N_42707);
nor U43454 (N_43454,N_42994,N_42980);
and U43455 (N_43455,N_42198,N_42424);
and U43456 (N_43456,N_42985,N_42776);
nor U43457 (N_43457,N_42321,N_42730);
or U43458 (N_43458,N_42862,N_42995);
or U43459 (N_43459,N_42803,N_42408);
or U43460 (N_43460,N_42966,N_42817);
or U43461 (N_43461,N_42112,N_42884);
nand U43462 (N_43462,N_42326,N_42661);
nand U43463 (N_43463,N_42785,N_42328);
nor U43464 (N_43464,N_42356,N_42006);
or U43465 (N_43465,N_42230,N_42301);
xor U43466 (N_43466,N_42181,N_42894);
nor U43467 (N_43467,N_42246,N_42289);
xnor U43468 (N_43468,N_42494,N_42432);
or U43469 (N_43469,N_42672,N_42443);
nor U43470 (N_43470,N_42319,N_42927);
or U43471 (N_43471,N_42646,N_42880);
or U43472 (N_43472,N_42255,N_42898);
nand U43473 (N_43473,N_42208,N_42413);
nor U43474 (N_43474,N_42622,N_42899);
and U43475 (N_43475,N_42217,N_42603);
xor U43476 (N_43476,N_42190,N_42576);
or U43477 (N_43477,N_42595,N_42422);
nand U43478 (N_43478,N_42366,N_42448);
nor U43479 (N_43479,N_42411,N_42530);
and U43480 (N_43480,N_42938,N_42749);
or U43481 (N_43481,N_42996,N_42738);
or U43482 (N_43482,N_42334,N_42399);
or U43483 (N_43483,N_42729,N_42148);
nor U43484 (N_43484,N_42215,N_42317);
and U43485 (N_43485,N_42689,N_42485);
or U43486 (N_43486,N_42225,N_42802);
nand U43487 (N_43487,N_42692,N_42396);
and U43488 (N_43488,N_42278,N_42117);
xor U43489 (N_43489,N_42723,N_42173);
xnor U43490 (N_43490,N_42583,N_42211);
nand U43491 (N_43491,N_42998,N_42546);
and U43492 (N_43492,N_42589,N_42936);
nor U43493 (N_43493,N_42395,N_42717);
nand U43494 (N_43494,N_42997,N_42478);
nand U43495 (N_43495,N_42421,N_42627);
and U43496 (N_43496,N_42078,N_42373);
and U43497 (N_43497,N_42042,N_42381);
xnor U43498 (N_43498,N_42640,N_42882);
nor U43499 (N_43499,N_42380,N_42235);
nor U43500 (N_43500,N_42974,N_42219);
nor U43501 (N_43501,N_42852,N_42122);
xnor U43502 (N_43502,N_42868,N_42934);
nor U43503 (N_43503,N_42755,N_42641);
and U43504 (N_43504,N_42104,N_42791);
nand U43505 (N_43505,N_42835,N_42294);
nand U43506 (N_43506,N_42062,N_42853);
and U43507 (N_43507,N_42163,N_42417);
and U43508 (N_43508,N_42795,N_42792);
nand U43509 (N_43509,N_42293,N_42912);
or U43510 (N_43510,N_42226,N_42556);
and U43511 (N_43511,N_42191,N_42148);
and U43512 (N_43512,N_42517,N_42759);
and U43513 (N_43513,N_42262,N_42575);
or U43514 (N_43514,N_42249,N_42549);
and U43515 (N_43515,N_42112,N_42275);
xnor U43516 (N_43516,N_42107,N_42806);
or U43517 (N_43517,N_42585,N_42658);
and U43518 (N_43518,N_42715,N_42052);
or U43519 (N_43519,N_42220,N_42251);
nand U43520 (N_43520,N_42693,N_42954);
or U43521 (N_43521,N_42109,N_42969);
xnor U43522 (N_43522,N_42547,N_42309);
and U43523 (N_43523,N_42836,N_42507);
nand U43524 (N_43524,N_42796,N_42767);
or U43525 (N_43525,N_42683,N_42863);
and U43526 (N_43526,N_42054,N_42248);
xor U43527 (N_43527,N_42848,N_42445);
nand U43528 (N_43528,N_42584,N_42172);
and U43529 (N_43529,N_42233,N_42015);
xnor U43530 (N_43530,N_42158,N_42296);
and U43531 (N_43531,N_42210,N_42035);
xnor U43532 (N_43532,N_42011,N_42669);
nor U43533 (N_43533,N_42170,N_42153);
or U43534 (N_43534,N_42294,N_42379);
or U43535 (N_43535,N_42385,N_42480);
nand U43536 (N_43536,N_42529,N_42478);
nand U43537 (N_43537,N_42100,N_42437);
and U43538 (N_43538,N_42005,N_42162);
and U43539 (N_43539,N_42442,N_42118);
nor U43540 (N_43540,N_42428,N_42571);
and U43541 (N_43541,N_42711,N_42319);
xor U43542 (N_43542,N_42963,N_42912);
and U43543 (N_43543,N_42208,N_42235);
or U43544 (N_43544,N_42640,N_42689);
nor U43545 (N_43545,N_42821,N_42431);
nor U43546 (N_43546,N_42878,N_42964);
xnor U43547 (N_43547,N_42746,N_42812);
xor U43548 (N_43548,N_42817,N_42226);
or U43549 (N_43549,N_42948,N_42956);
or U43550 (N_43550,N_42186,N_42862);
nand U43551 (N_43551,N_42975,N_42259);
nor U43552 (N_43552,N_42857,N_42705);
and U43553 (N_43553,N_42497,N_42443);
nor U43554 (N_43554,N_42491,N_42243);
nor U43555 (N_43555,N_42916,N_42226);
or U43556 (N_43556,N_42414,N_42100);
nand U43557 (N_43557,N_42804,N_42030);
nand U43558 (N_43558,N_42510,N_42500);
xnor U43559 (N_43559,N_42933,N_42380);
xor U43560 (N_43560,N_42981,N_42578);
nand U43561 (N_43561,N_42203,N_42225);
nor U43562 (N_43562,N_42126,N_42642);
nand U43563 (N_43563,N_42341,N_42433);
nor U43564 (N_43564,N_42000,N_42585);
and U43565 (N_43565,N_42489,N_42219);
and U43566 (N_43566,N_42582,N_42965);
and U43567 (N_43567,N_42511,N_42601);
nand U43568 (N_43568,N_42988,N_42796);
or U43569 (N_43569,N_42042,N_42336);
and U43570 (N_43570,N_42801,N_42044);
nand U43571 (N_43571,N_42989,N_42628);
or U43572 (N_43572,N_42275,N_42995);
nand U43573 (N_43573,N_42110,N_42126);
nor U43574 (N_43574,N_42043,N_42013);
nand U43575 (N_43575,N_42450,N_42280);
and U43576 (N_43576,N_42353,N_42202);
nor U43577 (N_43577,N_42656,N_42824);
nand U43578 (N_43578,N_42175,N_42641);
nand U43579 (N_43579,N_42597,N_42935);
nor U43580 (N_43580,N_42544,N_42435);
nor U43581 (N_43581,N_42066,N_42629);
nand U43582 (N_43582,N_42691,N_42987);
or U43583 (N_43583,N_42636,N_42628);
nor U43584 (N_43584,N_42250,N_42365);
or U43585 (N_43585,N_42958,N_42707);
nand U43586 (N_43586,N_42083,N_42451);
nand U43587 (N_43587,N_42154,N_42113);
nor U43588 (N_43588,N_42058,N_42951);
or U43589 (N_43589,N_42993,N_42328);
nor U43590 (N_43590,N_42558,N_42589);
nand U43591 (N_43591,N_42176,N_42996);
and U43592 (N_43592,N_42270,N_42060);
or U43593 (N_43593,N_42801,N_42571);
or U43594 (N_43594,N_42860,N_42063);
or U43595 (N_43595,N_42309,N_42376);
nor U43596 (N_43596,N_42053,N_42290);
and U43597 (N_43597,N_42551,N_42831);
nand U43598 (N_43598,N_42159,N_42202);
nand U43599 (N_43599,N_42130,N_42529);
nor U43600 (N_43600,N_42074,N_42910);
or U43601 (N_43601,N_42694,N_42405);
xor U43602 (N_43602,N_42761,N_42656);
nor U43603 (N_43603,N_42154,N_42948);
nand U43604 (N_43604,N_42080,N_42062);
and U43605 (N_43605,N_42451,N_42787);
nand U43606 (N_43606,N_42416,N_42744);
or U43607 (N_43607,N_42686,N_42317);
or U43608 (N_43608,N_42766,N_42138);
xnor U43609 (N_43609,N_42844,N_42030);
nor U43610 (N_43610,N_42171,N_42181);
and U43611 (N_43611,N_42307,N_42579);
or U43612 (N_43612,N_42483,N_42344);
nand U43613 (N_43613,N_42009,N_42609);
and U43614 (N_43614,N_42919,N_42982);
nor U43615 (N_43615,N_42763,N_42256);
nand U43616 (N_43616,N_42232,N_42082);
nand U43617 (N_43617,N_42587,N_42837);
nor U43618 (N_43618,N_42958,N_42518);
or U43619 (N_43619,N_42266,N_42616);
xnor U43620 (N_43620,N_42278,N_42427);
nand U43621 (N_43621,N_42225,N_42512);
nor U43622 (N_43622,N_42817,N_42912);
xnor U43623 (N_43623,N_42167,N_42196);
nand U43624 (N_43624,N_42268,N_42240);
xnor U43625 (N_43625,N_42771,N_42581);
or U43626 (N_43626,N_42966,N_42386);
nand U43627 (N_43627,N_42726,N_42188);
xnor U43628 (N_43628,N_42618,N_42905);
or U43629 (N_43629,N_42691,N_42835);
nand U43630 (N_43630,N_42026,N_42801);
xor U43631 (N_43631,N_42351,N_42413);
xor U43632 (N_43632,N_42375,N_42446);
and U43633 (N_43633,N_42915,N_42686);
nor U43634 (N_43634,N_42392,N_42478);
nand U43635 (N_43635,N_42200,N_42494);
nor U43636 (N_43636,N_42250,N_42273);
xnor U43637 (N_43637,N_42957,N_42949);
nor U43638 (N_43638,N_42582,N_42149);
xor U43639 (N_43639,N_42632,N_42251);
nand U43640 (N_43640,N_42849,N_42535);
or U43641 (N_43641,N_42566,N_42721);
and U43642 (N_43642,N_42384,N_42427);
or U43643 (N_43643,N_42173,N_42960);
or U43644 (N_43644,N_42885,N_42963);
and U43645 (N_43645,N_42632,N_42900);
nand U43646 (N_43646,N_42462,N_42896);
nand U43647 (N_43647,N_42810,N_42181);
xnor U43648 (N_43648,N_42603,N_42127);
xnor U43649 (N_43649,N_42660,N_42516);
nor U43650 (N_43650,N_42344,N_42667);
and U43651 (N_43651,N_42326,N_42070);
nand U43652 (N_43652,N_42749,N_42976);
and U43653 (N_43653,N_42529,N_42906);
and U43654 (N_43654,N_42897,N_42246);
nand U43655 (N_43655,N_42975,N_42021);
xor U43656 (N_43656,N_42941,N_42819);
nand U43657 (N_43657,N_42320,N_42239);
nor U43658 (N_43658,N_42214,N_42631);
and U43659 (N_43659,N_42462,N_42871);
and U43660 (N_43660,N_42066,N_42074);
and U43661 (N_43661,N_42861,N_42081);
nor U43662 (N_43662,N_42725,N_42034);
or U43663 (N_43663,N_42941,N_42905);
and U43664 (N_43664,N_42744,N_42675);
xnor U43665 (N_43665,N_42423,N_42791);
nand U43666 (N_43666,N_42592,N_42740);
and U43667 (N_43667,N_42683,N_42794);
and U43668 (N_43668,N_42801,N_42158);
or U43669 (N_43669,N_42687,N_42435);
or U43670 (N_43670,N_42803,N_42283);
nand U43671 (N_43671,N_42352,N_42083);
nand U43672 (N_43672,N_42690,N_42625);
or U43673 (N_43673,N_42722,N_42246);
nand U43674 (N_43674,N_42156,N_42771);
nand U43675 (N_43675,N_42691,N_42509);
nor U43676 (N_43676,N_42464,N_42211);
or U43677 (N_43677,N_42428,N_42481);
nor U43678 (N_43678,N_42844,N_42448);
or U43679 (N_43679,N_42811,N_42830);
and U43680 (N_43680,N_42741,N_42515);
xor U43681 (N_43681,N_42635,N_42226);
and U43682 (N_43682,N_42069,N_42475);
nor U43683 (N_43683,N_42386,N_42163);
xnor U43684 (N_43684,N_42919,N_42306);
xnor U43685 (N_43685,N_42433,N_42000);
xor U43686 (N_43686,N_42601,N_42955);
xnor U43687 (N_43687,N_42317,N_42278);
or U43688 (N_43688,N_42877,N_42960);
nand U43689 (N_43689,N_42518,N_42253);
nand U43690 (N_43690,N_42617,N_42719);
or U43691 (N_43691,N_42309,N_42366);
xnor U43692 (N_43692,N_42322,N_42062);
or U43693 (N_43693,N_42709,N_42894);
and U43694 (N_43694,N_42599,N_42159);
xnor U43695 (N_43695,N_42938,N_42046);
xor U43696 (N_43696,N_42159,N_42950);
nor U43697 (N_43697,N_42176,N_42499);
nor U43698 (N_43698,N_42044,N_42419);
or U43699 (N_43699,N_42838,N_42725);
xor U43700 (N_43700,N_42704,N_42447);
and U43701 (N_43701,N_42180,N_42673);
xnor U43702 (N_43702,N_42620,N_42005);
and U43703 (N_43703,N_42657,N_42769);
and U43704 (N_43704,N_42048,N_42486);
nor U43705 (N_43705,N_42997,N_42072);
or U43706 (N_43706,N_42610,N_42400);
nand U43707 (N_43707,N_42074,N_42310);
and U43708 (N_43708,N_42088,N_42732);
nand U43709 (N_43709,N_42880,N_42446);
or U43710 (N_43710,N_42232,N_42327);
and U43711 (N_43711,N_42132,N_42093);
nor U43712 (N_43712,N_42793,N_42750);
xor U43713 (N_43713,N_42229,N_42418);
or U43714 (N_43714,N_42417,N_42824);
nand U43715 (N_43715,N_42316,N_42383);
nand U43716 (N_43716,N_42781,N_42151);
nor U43717 (N_43717,N_42059,N_42361);
and U43718 (N_43718,N_42569,N_42335);
nor U43719 (N_43719,N_42302,N_42506);
and U43720 (N_43720,N_42146,N_42307);
and U43721 (N_43721,N_42026,N_42421);
nor U43722 (N_43722,N_42925,N_42941);
and U43723 (N_43723,N_42527,N_42296);
xor U43724 (N_43724,N_42641,N_42612);
and U43725 (N_43725,N_42479,N_42918);
nand U43726 (N_43726,N_42151,N_42684);
nor U43727 (N_43727,N_42471,N_42500);
nor U43728 (N_43728,N_42499,N_42987);
xor U43729 (N_43729,N_42119,N_42230);
nor U43730 (N_43730,N_42483,N_42524);
xor U43731 (N_43731,N_42976,N_42381);
nand U43732 (N_43732,N_42465,N_42476);
and U43733 (N_43733,N_42686,N_42424);
or U43734 (N_43734,N_42271,N_42538);
xor U43735 (N_43735,N_42248,N_42950);
nor U43736 (N_43736,N_42115,N_42515);
and U43737 (N_43737,N_42966,N_42686);
nand U43738 (N_43738,N_42859,N_42709);
nand U43739 (N_43739,N_42277,N_42415);
and U43740 (N_43740,N_42650,N_42756);
or U43741 (N_43741,N_42986,N_42822);
xnor U43742 (N_43742,N_42670,N_42810);
nand U43743 (N_43743,N_42363,N_42520);
or U43744 (N_43744,N_42917,N_42946);
nand U43745 (N_43745,N_42961,N_42244);
nand U43746 (N_43746,N_42900,N_42745);
and U43747 (N_43747,N_42872,N_42920);
nand U43748 (N_43748,N_42214,N_42819);
nor U43749 (N_43749,N_42482,N_42886);
or U43750 (N_43750,N_42028,N_42990);
nor U43751 (N_43751,N_42249,N_42462);
xor U43752 (N_43752,N_42040,N_42734);
xnor U43753 (N_43753,N_42682,N_42588);
xor U43754 (N_43754,N_42616,N_42286);
nor U43755 (N_43755,N_42031,N_42121);
xor U43756 (N_43756,N_42828,N_42327);
nand U43757 (N_43757,N_42440,N_42724);
or U43758 (N_43758,N_42754,N_42242);
xnor U43759 (N_43759,N_42187,N_42251);
and U43760 (N_43760,N_42610,N_42871);
and U43761 (N_43761,N_42124,N_42855);
nand U43762 (N_43762,N_42333,N_42059);
and U43763 (N_43763,N_42715,N_42373);
nor U43764 (N_43764,N_42919,N_42451);
and U43765 (N_43765,N_42465,N_42585);
nand U43766 (N_43766,N_42446,N_42186);
and U43767 (N_43767,N_42241,N_42800);
and U43768 (N_43768,N_42950,N_42269);
and U43769 (N_43769,N_42381,N_42341);
or U43770 (N_43770,N_42990,N_42356);
nand U43771 (N_43771,N_42507,N_42630);
xnor U43772 (N_43772,N_42682,N_42451);
nor U43773 (N_43773,N_42713,N_42987);
nor U43774 (N_43774,N_42029,N_42779);
and U43775 (N_43775,N_42952,N_42153);
nor U43776 (N_43776,N_42920,N_42363);
xnor U43777 (N_43777,N_42085,N_42618);
nor U43778 (N_43778,N_42583,N_42342);
nand U43779 (N_43779,N_42845,N_42328);
nand U43780 (N_43780,N_42884,N_42882);
nand U43781 (N_43781,N_42534,N_42708);
nor U43782 (N_43782,N_42270,N_42588);
xor U43783 (N_43783,N_42931,N_42489);
or U43784 (N_43784,N_42984,N_42037);
nor U43785 (N_43785,N_42081,N_42269);
xnor U43786 (N_43786,N_42890,N_42667);
and U43787 (N_43787,N_42333,N_42908);
nor U43788 (N_43788,N_42217,N_42721);
nor U43789 (N_43789,N_42965,N_42337);
nor U43790 (N_43790,N_42299,N_42692);
nor U43791 (N_43791,N_42855,N_42366);
nand U43792 (N_43792,N_42592,N_42923);
or U43793 (N_43793,N_42193,N_42973);
nor U43794 (N_43794,N_42316,N_42097);
nor U43795 (N_43795,N_42150,N_42978);
nor U43796 (N_43796,N_42838,N_42969);
nand U43797 (N_43797,N_42729,N_42443);
nand U43798 (N_43798,N_42012,N_42272);
and U43799 (N_43799,N_42186,N_42866);
nand U43800 (N_43800,N_42476,N_42483);
nor U43801 (N_43801,N_42078,N_42860);
and U43802 (N_43802,N_42297,N_42695);
nor U43803 (N_43803,N_42127,N_42031);
nand U43804 (N_43804,N_42879,N_42591);
nand U43805 (N_43805,N_42703,N_42057);
nor U43806 (N_43806,N_42519,N_42466);
or U43807 (N_43807,N_42311,N_42873);
and U43808 (N_43808,N_42330,N_42395);
nor U43809 (N_43809,N_42421,N_42392);
or U43810 (N_43810,N_42139,N_42305);
nand U43811 (N_43811,N_42669,N_42227);
xor U43812 (N_43812,N_42266,N_42120);
and U43813 (N_43813,N_42627,N_42921);
or U43814 (N_43814,N_42356,N_42833);
xor U43815 (N_43815,N_42705,N_42110);
nor U43816 (N_43816,N_42772,N_42305);
and U43817 (N_43817,N_42954,N_42903);
or U43818 (N_43818,N_42599,N_42022);
or U43819 (N_43819,N_42082,N_42845);
and U43820 (N_43820,N_42427,N_42300);
or U43821 (N_43821,N_42862,N_42683);
nor U43822 (N_43822,N_42096,N_42603);
and U43823 (N_43823,N_42660,N_42018);
nand U43824 (N_43824,N_42126,N_42851);
nor U43825 (N_43825,N_42427,N_42877);
or U43826 (N_43826,N_42700,N_42106);
and U43827 (N_43827,N_42040,N_42186);
xnor U43828 (N_43828,N_42111,N_42720);
nand U43829 (N_43829,N_42747,N_42845);
nand U43830 (N_43830,N_42355,N_42413);
nor U43831 (N_43831,N_42657,N_42153);
and U43832 (N_43832,N_42290,N_42789);
and U43833 (N_43833,N_42502,N_42609);
xnor U43834 (N_43834,N_42230,N_42706);
and U43835 (N_43835,N_42140,N_42024);
nor U43836 (N_43836,N_42897,N_42847);
or U43837 (N_43837,N_42806,N_42710);
nor U43838 (N_43838,N_42875,N_42374);
xnor U43839 (N_43839,N_42648,N_42800);
and U43840 (N_43840,N_42940,N_42358);
nand U43841 (N_43841,N_42457,N_42973);
nor U43842 (N_43842,N_42072,N_42537);
nand U43843 (N_43843,N_42193,N_42997);
xor U43844 (N_43844,N_42501,N_42931);
nand U43845 (N_43845,N_42055,N_42111);
and U43846 (N_43846,N_42672,N_42092);
or U43847 (N_43847,N_42222,N_42607);
nand U43848 (N_43848,N_42370,N_42263);
nor U43849 (N_43849,N_42941,N_42161);
xor U43850 (N_43850,N_42610,N_42798);
or U43851 (N_43851,N_42954,N_42762);
xor U43852 (N_43852,N_42719,N_42461);
and U43853 (N_43853,N_42873,N_42628);
and U43854 (N_43854,N_42372,N_42223);
xnor U43855 (N_43855,N_42773,N_42387);
xor U43856 (N_43856,N_42518,N_42495);
nor U43857 (N_43857,N_42403,N_42615);
or U43858 (N_43858,N_42390,N_42134);
or U43859 (N_43859,N_42265,N_42784);
or U43860 (N_43860,N_42133,N_42723);
nor U43861 (N_43861,N_42450,N_42547);
xnor U43862 (N_43862,N_42974,N_42689);
xnor U43863 (N_43863,N_42426,N_42810);
nor U43864 (N_43864,N_42468,N_42952);
xor U43865 (N_43865,N_42270,N_42616);
nand U43866 (N_43866,N_42644,N_42222);
nor U43867 (N_43867,N_42716,N_42008);
nand U43868 (N_43868,N_42750,N_42095);
and U43869 (N_43869,N_42725,N_42828);
nor U43870 (N_43870,N_42201,N_42573);
or U43871 (N_43871,N_42806,N_42824);
and U43872 (N_43872,N_42572,N_42005);
xor U43873 (N_43873,N_42499,N_42281);
and U43874 (N_43874,N_42832,N_42200);
and U43875 (N_43875,N_42317,N_42665);
and U43876 (N_43876,N_42729,N_42702);
nand U43877 (N_43877,N_42151,N_42066);
xnor U43878 (N_43878,N_42127,N_42175);
and U43879 (N_43879,N_42429,N_42949);
xor U43880 (N_43880,N_42560,N_42885);
nand U43881 (N_43881,N_42624,N_42483);
or U43882 (N_43882,N_42863,N_42785);
xor U43883 (N_43883,N_42709,N_42492);
and U43884 (N_43884,N_42200,N_42339);
nand U43885 (N_43885,N_42522,N_42279);
nor U43886 (N_43886,N_42808,N_42807);
or U43887 (N_43887,N_42934,N_42881);
nand U43888 (N_43888,N_42528,N_42908);
and U43889 (N_43889,N_42055,N_42510);
or U43890 (N_43890,N_42192,N_42253);
or U43891 (N_43891,N_42494,N_42050);
or U43892 (N_43892,N_42260,N_42902);
xnor U43893 (N_43893,N_42334,N_42518);
and U43894 (N_43894,N_42519,N_42544);
xor U43895 (N_43895,N_42325,N_42207);
and U43896 (N_43896,N_42669,N_42631);
and U43897 (N_43897,N_42530,N_42602);
nand U43898 (N_43898,N_42715,N_42324);
and U43899 (N_43899,N_42893,N_42734);
nor U43900 (N_43900,N_42632,N_42948);
xnor U43901 (N_43901,N_42205,N_42376);
nor U43902 (N_43902,N_42866,N_42399);
nand U43903 (N_43903,N_42045,N_42360);
or U43904 (N_43904,N_42600,N_42445);
nor U43905 (N_43905,N_42006,N_42909);
nand U43906 (N_43906,N_42670,N_42577);
nand U43907 (N_43907,N_42301,N_42755);
or U43908 (N_43908,N_42416,N_42348);
or U43909 (N_43909,N_42033,N_42973);
nand U43910 (N_43910,N_42717,N_42780);
nand U43911 (N_43911,N_42406,N_42821);
nor U43912 (N_43912,N_42242,N_42795);
or U43913 (N_43913,N_42525,N_42141);
and U43914 (N_43914,N_42423,N_42505);
nor U43915 (N_43915,N_42907,N_42833);
or U43916 (N_43916,N_42620,N_42768);
xnor U43917 (N_43917,N_42894,N_42134);
or U43918 (N_43918,N_42132,N_42332);
or U43919 (N_43919,N_42919,N_42529);
nor U43920 (N_43920,N_42442,N_42613);
xor U43921 (N_43921,N_42119,N_42413);
nor U43922 (N_43922,N_42992,N_42891);
nand U43923 (N_43923,N_42668,N_42065);
xor U43924 (N_43924,N_42715,N_42876);
nand U43925 (N_43925,N_42638,N_42563);
nor U43926 (N_43926,N_42440,N_42923);
or U43927 (N_43927,N_42522,N_42884);
or U43928 (N_43928,N_42637,N_42464);
nand U43929 (N_43929,N_42018,N_42319);
nor U43930 (N_43930,N_42403,N_42673);
or U43931 (N_43931,N_42669,N_42318);
and U43932 (N_43932,N_42988,N_42881);
nor U43933 (N_43933,N_42256,N_42499);
nand U43934 (N_43934,N_42086,N_42622);
nand U43935 (N_43935,N_42713,N_42824);
nor U43936 (N_43936,N_42925,N_42098);
or U43937 (N_43937,N_42309,N_42472);
nand U43938 (N_43938,N_42380,N_42238);
or U43939 (N_43939,N_42901,N_42099);
xnor U43940 (N_43940,N_42392,N_42295);
or U43941 (N_43941,N_42341,N_42041);
nor U43942 (N_43942,N_42009,N_42301);
nand U43943 (N_43943,N_42713,N_42277);
xor U43944 (N_43944,N_42512,N_42517);
nand U43945 (N_43945,N_42861,N_42623);
or U43946 (N_43946,N_42903,N_42873);
nand U43947 (N_43947,N_42982,N_42878);
or U43948 (N_43948,N_42160,N_42876);
nand U43949 (N_43949,N_42198,N_42923);
or U43950 (N_43950,N_42666,N_42763);
nor U43951 (N_43951,N_42836,N_42310);
nor U43952 (N_43952,N_42451,N_42598);
nand U43953 (N_43953,N_42867,N_42259);
xor U43954 (N_43954,N_42247,N_42488);
or U43955 (N_43955,N_42363,N_42387);
xor U43956 (N_43956,N_42430,N_42314);
nand U43957 (N_43957,N_42073,N_42019);
nand U43958 (N_43958,N_42465,N_42183);
and U43959 (N_43959,N_42305,N_42187);
nor U43960 (N_43960,N_42675,N_42482);
nand U43961 (N_43961,N_42002,N_42441);
and U43962 (N_43962,N_42589,N_42142);
nand U43963 (N_43963,N_42711,N_42341);
nand U43964 (N_43964,N_42776,N_42995);
or U43965 (N_43965,N_42905,N_42708);
xor U43966 (N_43966,N_42466,N_42966);
xnor U43967 (N_43967,N_42692,N_42673);
or U43968 (N_43968,N_42188,N_42827);
or U43969 (N_43969,N_42263,N_42426);
nor U43970 (N_43970,N_42778,N_42451);
and U43971 (N_43971,N_42607,N_42754);
nand U43972 (N_43972,N_42828,N_42569);
nand U43973 (N_43973,N_42992,N_42852);
and U43974 (N_43974,N_42026,N_42133);
xnor U43975 (N_43975,N_42449,N_42826);
xor U43976 (N_43976,N_42879,N_42489);
xor U43977 (N_43977,N_42624,N_42034);
and U43978 (N_43978,N_42983,N_42535);
nor U43979 (N_43979,N_42360,N_42121);
xor U43980 (N_43980,N_42442,N_42891);
nand U43981 (N_43981,N_42366,N_42275);
nand U43982 (N_43982,N_42572,N_42320);
and U43983 (N_43983,N_42497,N_42069);
nand U43984 (N_43984,N_42078,N_42831);
and U43985 (N_43985,N_42384,N_42619);
or U43986 (N_43986,N_42430,N_42725);
nand U43987 (N_43987,N_42176,N_42386);
xor U43988 (N_43988,N_42431,N_42008);
or U43989 (N_43989,N_42298,N_42982);
xor U43990 (N_43990,N_42442,N_42225);
xnor U43991 (N_43991,N_42813,N_42304);
and U43992 (N_43992,N_42792,N_42115);
and U43993 (N_43993,N_42929,N_42457);
nand U43994 (N_43994,N_42570,N_42147);
nor U43995 (N_43995,N_42356,N_42117);
nand U43996 (N_43996,N_42217,N_42997);
or U43997 (N_43997,N_42235,N_42743);
nor U43998 (N_43998,N_42575,N_42336);
nor U43999 (N_43999,N_42012,N_42058);
xnor U44000 (N_44000,N_43780,N_43520);
nand U44001 (N_44001,N_43262,N_43135);
nand U44002 (N_44002,N_43014,N_43556);
or U44003 (N_44003,N_43199,N_43862);
xor U44004 (N_44004,N_43063,N_43933);
nand U44005 (N_44005,N_43721,N_43163);
xnor U44006 (N_44006,N_43958,N_43159);
xnor U44007 (N_44007,N_43311,N_43639);
nor U44008 (N_44008,N_43989,N_43422);
nand U44009 (N_44009,N_43859,N_43593);
and U44010 (N_44010,N_43045,N_43632);
and U44011 (N_44011,N_43258,N_43697);
or U44012 (N_44012,N_43146,N_43181);
xnor U44013 (N_44013,N_43255,N_43860);
nand U44014 (N_44014,N_43562,N_43910);
and U44015 (N_44015,N_43162,N_43875);
nand U44016 (N_44016,N_43692,N_43819);
and U44017 (N_44017,N_43242,N_43332);
nor U44018 (N_44018,N_43081,N_43038);
nor U44019 (N_44019,N_43459,N_43726);
nor U44020 (N_44020,N_43441,N_43600);
xor U44021 (N_44021,N_43644,N_43153);
nor U44022 (N_44022,N_43698,N_43306);
xor U44023 (N_44023,N_43013,N_43670);
nand U44024 (N_44024,N_43866,N_43088);
or U44025 (N_44025,N_43288,N_43770);
and U44026 (N_44026,N_43749,N_43265);
xnor U44027 (N_44027,N_43051,N_43517);
nor U44028 (N_44028,N_43673,N_43226);
nand U44029 (N_44029,N_43330,N_43512);
nand U44030 (N_44030,N_43260,N_43050);
xor U44031 (N_44031,N_43779,N_43429);
xnor U44032 (N_44032,N_43508,N_43037);
xor U44033 (N_44033,N_43572,N_43084);
or U44034 (N_44034,N_43083,N_43873);
nor U44035 (N_44035,N_43765,N_43812);
or U44036 (N_44036,N_43060,N_43237);
or U44037 (N_44037,N_43022,N_43233);
nor U44038 (N_44038,N_43743,N_43195);
xor U44039 (N_44039,N_43830,N_43701);
or U44040 (N_44040,N_43884,N_43966);
nor U44041 (N_44041,N_43118,N_43956);
or U44042 (N_44042,N_43164,N_43514);
xor U44043 (N_44043,N_43114,N_43838);
nand U44044 (N_44044,N_43115,N_43753);
nor U44045 (N_44045,N_43229,N_43573);
or U44046 (N_44046,N_43651,N_43519);
xnor U44047 (N_44047,N_43621,N_43494);
xnor U44048 (N_44048,N_43089,N_43535);
nor U44049 (N_44049,N_43827,N_43287);
or U44050 (N_44050,N_43206,N_43559);
or U44051 (N_44051,N_43309,N_43557);
and U44052 (N_44052,N_43348,N_43820);
nand U44053 (N_44053,N_43776,N_43495);
xnor U44054 (N_44054,N_43664,N_43945);
nand U44055 (N_44055,N_43997,N_43683);
nand U44056 (N_44056,N_43406,N_43604);
or U44057 (N_44057,N_43339,N_43205);
and U44058 (N_44058,N_43863,N_43728);
nand U44059 (N_44059,N_43620,N_43546);
nor U44060 (N_44060,N_43794,N_43640);
and U44061 (N_44061,N_43814,N_43847);
and U44062 (N_44062,N_43592,N_43951);
nor U44063 (N_44063,N_43591,N_43035);
or U44064 (N_44064,N_43684,N_43202);
and U44065 (N_44065,N_43053,N_43527);
or U44066 (N_44066,N_43536,N_43563);
and U44067 (N_44067,N_43371,N_43586);
and U44068 (N_44068,N_43104,N_43751);
nand U44069 (N_44069,N_43074,N_43021);
or U44070 (N_44070,N_43361,N_43165);
or U44071 (N_44071,N_43434,N_43221);
and U44072 (N_44072,N_43039,N_43606);
nand U44073 (N_44073,N_43289,N_43445);
and U44074 (N_44074,N_43452,N_43807);
and U44075 (N_44075,N_43950,N_43627);
nor U44076 (N_44076,N_43403,N_43888);
xor U44077 (N_44077,N_43525,N_43842);
or U44078 (N_44078,N_43183,N_43731);
xnor U44079 (N_44079,N_43871,N_43954);
nor U44080 (N_44080,N_43518,N_43451);
xnor U44081 (N_44081,N_43741,N_43688);
nand U44082 (N_44082,N_43388,N_43382);
nor U44083 (N_44083,N_43702,N_43845);
nand U44084 (N_44084,N_43419,N_43856);
and U44085 (N_44085,N_43355,N_43138);
nor U44086 (N_44086,N_43824,N_43170);
nor U44087 (N_44087,N_43674,N_43381);
and U44088 (N_44088,N_43119,N_43669);
or U44089 (N_44089,N_43300,N_43444);
or U44090 (N_44090,N_43178,N_43576);
nand U44091 (N_44091,N_43389,N_43897);
or U44092 (N_44092,N_43618,N_43668);
xor U44093 (N_44093,N_43299,N_43257);
nand U44094 (N_44094,N_43003,N_43048);
or U44095 (N_44095,N_43788,N_43762);
or U44096 (N_44096,N_43052,N_43887);
and U44097 (N_44097,N_43108,N_43077);
and U44098 (N_44098,N_43549,N_43868);
xor U44099 (N_44099,N_43545,N_43432);
nand U44100 (N_44100,N_43764,N_43316);
or U44101 (N_44101,N_43695,N_43009);
and U44102 (N_44102,N_43366,N_43486);
or U44103 (N_44103,N_43786,N_43189);
or U44104 (N_44104,N_43141,N_43948);
nand U44105 (N_44105,N_43942,N_43015);
xnor U44106 (N_44106,N_43658,N_43537);
nor U44107 (N_44107,N_43986,N_43857);
xnor U44108 (N_44108,N_43869,N_43426);
or U44109 (N_44109,N_43338,N_43815);
and U44110 (N_44110,N_43059,N_43811);
nor U44111 (N_44111,N_43047,N_43374);
or U44112 (N_44112,N_43437,N_43369);
nand U44113 (N_44113,N_43107,N_43923);
or U44114 (N_44114,N_43078,N_43589);
nand U44115 (N_44115,N_43921,N_43172);
or U44116 (N_44116,N_43929,N_43372);
xor U44117 (N_44117,N_43346,N_43973);
nand U44118 (N_44118,N_43926,N_43515);
or U44119 (N_44119,N_43666,N_43781);
nand U44120 (N_44120,N_43425,N_43540);
or U44121 (N_44121,N_43511,N_43832);
xnor U44122 (N_44122,N_43342,N_43681);
and U44123 (N_44123,N_43630,N_43924);
nand U44124 (N_44124,N_43834,N_43482);
xnor U44125 (N_44125,N_43131,N_43818);
or U44126 (N_44126,N_43218,N_43200);
and U44127 (N_44127,N_43724,N_43203);
and U44128 (N_44128,N_43803,N_43891);
nand U44129 (N_44129,N_43391,N_43967);
or U44130 (N_44130,N_43358,N_43173);
nor U44131 (N_44131,N_43019,N_43744);
or U44132 (N_44132,N_43392,N_43831);
xor U44133 (N_44133,N_43631,N_43436);
and U44134 (N_44134,N_43828,N_43716);
nand U44135 (N_44135,N_43241,N_43976);
and U44136 (N_44136,N_43784,N_43413);
xnor U44137 (N_44137,N_43882,N_43236);
nand U44138 (N_44138,N_43028,N_43912);
nand U44139 (N_44139,N_43405,N_43217);
nor U44140 (N_44140,N_43072,N_43465);
nor U44141 (N_44141,N_43097,N_43516);
nor U44142 (N_44142,N_43379,N_43182);
xnor U44143 (N_44143,N_43791,N_43944);
xnor U44144 (N_44144,N_43192,N_43808);
xor U44145 (N_44145,N_43416,N_43491);
nand U44146 (N_44146,N_43295,N_43732);
nor U44147 (N_44147,N_43970,N_43583);
nand U44148 (N_44148,N_43715,N_43778);
nand U44149 (N_44149,N_43324,N_43805);
and U44150 (N_44150,N_43936,N_43569);
nand U44151 (N_44151,N_43595,N_43775);
or U44152 (N_44152,N_43499,N_43685);
and U44153 (N_44153,N_43133,N_43602);
nor U44154 (N_44154,N_43801,N_43007);
and U44155 (N_44155,N_43552,N_43030);
nand U44156 (N_44156,N_43325,N_43806);
xnor U44157 (N_44157,N_43132,N_43689);
or U44158 (N_44158,N_43079,N_43106);
and U44159 (N_44159,N_43251,N_43542);
xor U44160 (N_44160,N_43605,N_43817);
nand U44161 (N_44161,N_43064,N_43756);
xor U44162 (N_44162,N_43782,N_43787);
or U44163 (N_44163,N_43949,N_43191);
and U44164 (N_44164,N_43993,N_43964);
and U44165 (N_44165,N_43049,N_43799);
xnor U44166 (N_44166,N_43566,N_43303);
or U44167 (N_44167,N_43027,N_43623);
and U44168 (N_44168,N_43383,N_43718);
or U44169 (N_44169,N_43619,N_43267);
nand U44170 (N_44170,N_43266,N_43872);
nor U44171 (N_44171,N_43550,N_43450);
xnor U44172 (N_44172,N_43087,N_43385);
nor U44173 (N_44173,N_43931,N_43373);
xor U44174 (N_44174,N_43679,N_43755);
or U44175 (N_44175,N_43502,N_43018);
nand U44176 (N_44176,N_43911,N_43171);
and U44177 (N_44177,N_43574,N_43433);
nor U44178 (N_44178,N_43150,N_43328);
or U44179 (N_44179,N_43029,N_43877);
nor U44180 (N_44180,N_43430,N_43895);
and U44181 (N_44181,N_43570,N_43611);
xnor U44182 (N_44182,N_43344,N_43402);
xor U44183 (N_44183,N_43424,N_43941);
nand U44184 (N_44184,N_43657,N_43367);
or U44185 (N_44185,N_43503,N_43228);
or U44186 (N_44186,N_43614,N_43613);
and U44187 (N_44187,N_43365,N_43747);
or U44188 (N_44188,N_43854,N_43472);
xnor U44189 (N_44189,N_43336,N_43323);
nor U44190 (N_44190,N_43759,N_43443);
and U44191 (N_44191,N_43149,N_43905);
and U44192 (N_44192,N_43901,N_43054);
nor U44193 (N_44193,N_43313,N_43748);
nor U44194 (N_44194,N_43634,N_43411);
nor U44195 (N_44195,N_43531,N_43376);
nand U44196 (N_44196,N_43101,N_43560);
nor U44197 (N_44197,N_43547,N_43125);
nand U44198 (N_44198,N_43194,N_43008);
and U44199 (N_44199,N_43678,N_43294);
xor U44200 (N_44200,N_43044,N_43310);
or U44201 (N_44201,N_43913,N_43036);
xor U44202 (N_44202,N_43301,N_43103);
and U44203 (N_44203,N_43487,N_43705);
nand U44204 (N_44204,N_43920,N_43766);
nand U44205 (N_44205,N_43767,N_43588);
nand U44206 (N_44206,N_43709,N_43496);
nor U44207 (N_44207,N_43682,N_43041);
and U44208 (N_44208,N_43963,N_43250);
nor U44209 (N_44209,N_43646,N_43498);
nand U44210 (N_44210,N_43273,N_43160);
nand U44211 (N_44211,N_43675,N_43703);
and U44212 (N_44212,N_43090,N_43031);
and U44213 (N_44213,N_43983,N_43603);
nor U44214 (N_44214,N_43720,N_43220);
or U44215 (N_44215,N_43271,N_43187);
nand U44216 (N_44216,N_43809,N_43354);
and U44217 (N_44217,N_43387,N_43446);
nor U44218 (N_44218,N_43733,N_43186);
and U44219 (N_44219,N_43507,N_43004);
and U44220 (N_44220,N_43057,N_43215);
and U44221 (N_44221,N_43974,N_43408);
nand U44222 (N_44222,N_43211,N_43981);
xor U44223 (N_44223,N_43965,N_43881);
nand U44224 (N_44224,N_43100,N_43687);
nor U44225 (N_44225,N_43501,N_43431);
xor U44226 (N_44226,N_43005,N_43174);
or U44227 (N_44227,N_43399,N_43940);
nand U44228 (N_44228,N_43351,N_43239);
or U44229 (N_44229,N_43151,N_43581);
or U44230 (N_44230,N_43480,N_43633);
nor U44231 (N_44231,N_43719,N_43608);
nand U44232 (N_44232,N_43637,N_43112);
nor U44233 (N_44233,N_43410,N_43461);
xor U44234 (N_44234,N_43340,N_43582);
xnor U44235 (N_44235,N_43175,N_43412);
xor U44236 (N_44236,N_43281,N_43179);
and U44237 (N_44237,N_43243,N_43968);
or U44238 (N_44238,N_43102,N_43925);
xor U44239 (N_44239,N_43326,N_43541);
or U44240 (N_44240,N_43145,N_43398);
and U44241 (N_44241,N_43746,N_43110);
xor U44242 (N_44242,N_43816,N_43427);
and U44243 (N_44243,N_43256,N_43850);
and U44244 (N_44244,N_43626,N_43209);
or U44245 (N_44245,N_43700,N_43774);
xor U44246 (N_44246,N_43990,N_43473);
nand U44247 (N_44247,N_43645,N_43284);
and U44248 (N_44248,N_43065,N_43224);
or U44249 (N_44249,N_43898,N_43699);
xor U44250 (N_44250,N_43717,N_43404);
nand U44251 (N_44251,N_43154,N_43693);
and U44252 (N_44252,N_43609,N_43982);
xnor U44253 (N_44253,N_43418,N_43136);
and U44254 (N_44254,N_43140,N_43972);
nor U44255 (N_44255,N_43423,N_43907);
or U44256 (N_44256,N_43704,N_43095);
nand U44257 (N_44257,N_43977,N_43456);
or U44258 (N_44258,N_43690,N_43772);
nor U44259 (N_44259,N_43971,N_43032);
or U44260 (N_44260,N_43401,N_43393);
and U44261 (N_44261,N_43510,N_43528);
nand U44262 (N_44262,N_43661,N_43016);
xnor U44263 (N_44263,N_43476,N_43522);
nor U44264 (N_44264,N_43488,N_43315);
or U44265 (N_44265,N_43587,N_43909);
xnor U44266 (N_44266,N_43447,N_43353);
and U44267 (N_44267,N_43386,N_43073);
nand U44268 (N_44268,N_43752,N_43865);
nand U44269 (N_44269,N_43580,N_43002);
and U44270 (N_44270,N_43278,N_43396);
xnor U44271 (N_44271,N_43479,N_43290);
nor U44272 (N_44272,N_43335,N_43214);
xor U44273 (N_44273,N_43319,N_43952);
or U44274 (N_44274,N_43046,N_43442);
nand U44275 (N_44275,N_43650,N_43244);
nor U44276 (N_44276,N_43298,N_43467);
nand U44277 (N_44277,N_43708,N_43435);
nor U44278 (N_44278,N_43270,N_43343);
nor U44279 (N_44279,N_43378,N_43852);
xor U44280 (N_44280,N_43493,N_43105);
or U44281 (N_44281,N_43594,N_43204);
xor U44282 (N_44282,N_43252,N_43564);
nor U44283 (N_44283,N_43111,N_43567);
xor U44284 (N_44284,N_43988,N_43185);
nand U44285 (N_44285,N_43919,N_43730);
nand U44286 (N_44286,N_43915,N_43208);
and U44287 (N_44287,N_43397,N_43723);
nand U44288 (N_44288,N_43960,N_43129);
and U44289 (N_44289,N_43616,N_43980);
and U44290 (N_44290,N_43825,N_43795);
or U44291 (N_44291,N_43462,N_43068);
nor U44292 (N_44292,N_43737,N_43835);
nand U44293 (N_44293,N_43883,N_43011);
nand U44294 (N_44294,N_43497,N_43538);
or U44295 (N_44295,N_43622,N_43219);
nor U44296 (N_44296,N_43813,N_43509);
nor U44297 (N_44297,N_43240,N_43978);
nor U44298 (N_44298,N_43984,N_43349);
xor U44299 (N_44299,N_43998,N_43390);
nand U44300 (N_44300,N_43197,N_43238);
nand U44301 (N_44301,N_43802,N_43607);
or U44302 (N_44302,N_43020,N_43272);
xnor U44303 (N_44303,N_43523,N_43790);
xnor U44304 (N_44304,N_43177,N_43777);
nand U44305 (N_44305,N_43357,N_43890);
xor U44306 (N_44306,N_43417,N_43276);
nand U44307 (N_44307,N_43285,N_43122);
nand U44308 (N_44308,N_43846,N_43796);
or U44309 (N_44309,N_43995,N_43946);
nand U44310 (N_44310,N_43554,N_43096);
nor U44311 (N_44311,N_43001,N_43757);
nor U44312 (N_44312,N_43760,N_43449);
and U44313 (N_44313,N_43116,N_43269);
nor U44314 (N_44314,N_43291,N_43076);
or U44315 (N_44315,N_43261,N_43953);
or U44316 (N_44316,N_43286,N_43742);
xor U44317 (N_44317,N_43999,N_43789);
xor U44318 (N_44318,N_43212,N_43568);
xnor U44319 (N_44319,N_43505,N_43829);
and U44320 (N_44320,N_43649,N_43157);
or U44321 (N_44321,N_43320,N_43843);
nand U44322 (N_44322,N_43093,N_43858);
and U44323 (N_44323,N_43394,N_43712);
nand U44324 (N_44324,N_43341,N_43034);
or U44325 (N_44325,N_43484,N_43553);
nand U44326 (N_44326,N_43190,N_43460);
nor U44327 (N_44327,N_43707,N_43892);
nor U44328 (N_44328,N_43066,N_43010);
nand U44329 (N_44329,N_43327,N_43024);
or U44330 (N_44330,N_43263,N_43091);
and U44331 (N_44331,N_43662,N_43414);
nand U44332 (N_44332,N_43277,N_43914);
xor U44333 (N_44333,N_43070,N_43448);
nand U44334 (N_44334,N_43694,N_43302);
or U44335 (N_44335,N_43144,N_43962);
and U44336 (N_44336,N_43996,N_43458);
nor U44337 (N_44337,N_43198,N_43454);
and U44338 (N_44338,N_43653,N_43750);
nand U44339 (N_44339,N_43821,N_43082);
and U44340 (N_44340,N_43822,N_43169);
nand U44341 (N_44341,N_43143,N_43033);
nor U44342 (N_44342,N_43987,N_43483);
xor U44343 (N_44343,N_43314,N_43725);
and U44344 (N_44344,N_43322,N_43099);
nor U44345 (N_44345,N_43025,N_43738);
nor U44346 (N_44346,N_43331,N_43359);
xnor U44347 (N_44347,N_43360,N_43490);
xnor U44348 (N_44348,N_43660,N_43307);
xnor U44349 (N_44349,N_43635,N_43571);
xnor U44350 (N_44350,N_43370,N_43874);
or U44351 (N_44351,N_43994,N_43421);
nor U44352 (N_44352,N_43839,N_43853);
xnor U44353 (N_44353,N_43711,N_43544);
nor U44354 (N_44354,N_43561,N_43478);
nand U44355 (N_44355,N_43642,N_43533);
nor U44356 (N_44356,N_43156,N_43139);
or U44357 (N_44357,N_43530,N_43042);
or U44358 (N_44358,N_43227,N_43565);
and U44359 (N_44359,N_43597,N_43279);
and U44360 (N_44360,N_43513,N_43985);
or U44361 (N_44361,N_43590,N_43245);
and U44362 (N_44362,N_43722,N_43734);
or U44363 (N_44363,N_43475,N_43420);
and U44364 (N_44364,N_43889,N_43641);
xor U44365 (N_44365,N_43268,N_43109);
or U44366 (N_44366,N_43457,N_43826);
nand U44367 (N_44367,N_43648,N_43481);
xor U44368 (N_44368,N_43585,N_43727);
or U44369 (N_44369,N_43686,N_43333);
or U44370 (N_44370,N_43428,N_43006);
or U44371 (N_44371,N_43463,N_43012);
nor U44372 (N_44372,N_43903,N_43155);
xnor U44373 (N_44373,N_43934,N_43833);
or U44374 (N_44374,N_43400,N_43855);
nor U44375 (N_44375,N_43254,N_43293);
nand U44376 (N_44376,N_43375,N_43246);
nand U44377 (N_44377,N_43655,N_43321);
xor U44378 (N_44378,N_43124,N_43955);
nand U44379 (N_44379,N_43283,N_43935);
or U44380 (N_44380,N_43469,N_43026);
nor U44381 (N_44381,N_43017,N_43548);
nor U44382 (N_44382,N_43148,N_43362);
xnor U44383 (N_44383,N_43201,N_43292);
xnor U44384 (N_44384,N_43113,N_43939);
or U44385 (N_44385,N_43761,N_43489);
xor U44386 (N_44386,N_43659,N_43056);
or U44387 (N_44387,N_43395,N_43207);
xor U44388 (N_44388,N_43837,N_43745);
or U44389 (N_44389,N_43848,N_43893);
nand U44390 (N_44390,N_43071,N_43274);
and U44391 (N_44391,N_43928,N_43043);
and U44392 (N_44392,N_43575,N_43851);
nor U44393 (N_44393,N_43067,N_43629);
nor U44394 (N_44394,N_43308,N_43714);
and U44395 (N_44395,N_43961,N_43297);
nand U44396 (N_44396,N_43534,N_43098);
and U44397 (N_44397,N_43235,N_43894);
or U44398 (N_44398,N_43906,N_43213);
xnor U44399 (N_44399,N_43312,N_43532);
nand U44400 (N_44400,N_43176,N_43969);
nor U44401 (N_44401,N_43783,N_43713);
or U44402 (N_44402,N_43232,N_43610);
nand U44403 (N_44403,N_43667,N_43334);
nor U44404 (N_44404,N_43468,N_43729);
and U44405 (N_44405,N_43754,N_43180);
nand U44406 (N_44406,N_43264,N_43407);
and U44407 (N_44407,N_43222,N_43880);
or U44408 (N_44408,N_43652,N_43128);
xnor U44409 (N_44409,N_43638,N_43471);
nor U44410 (N_44410,N_43676,N_43167);
nand U44411 (N_44411,N_43710,N_43647);
nor U44412 (N_44412,N_43317,N_43671);
nor U44413 (N_44413,N_43804,N_43706);
nand U44414 (N_44414,N_43231,N_43477);
or U44415 (N_44415,N_43040,N_43768);
or U44416 (N_44416,N_43696,N_43612);
and U44417 (N_44417,N_43663,N_43259);
nand U44418 (N_44418,N_43885,N_43636);
nor U44419 (N_44419,N_43736,N_43094);
xnor U44420 (N_44420,N_43937,N_43453);
xnor U44421 (N_44421,N_43625,N_43356);
or U44422 (N_44422,N_43793,N_43504);
nand U44423 (N_44423,N_43130,N_43085);
and U44424 (N_44424,N_43474,N_43280);
nand U44425 (N_44425,N_43196,N_43080);
xnor U44426 (N_44426,N_43773,N_43957);
and U44427 (N_44427,N_43922,N_43415);
xnor U44428 (N_44428,N_43492,N_43409);
nor U44429 (N_44429,N_43555,N_43121);
nor U44430 (N_44430,N_43329,N_43943);
nand U44431 (N_44431,N_43296,N_43223);
nor U44432 (N_44432,N_43318,N_43158);
nor U44433 (N_44433,N_43867,N_43543);
xor U44434 (N_44434,N_43364,N_43628);
or U44435 (N_44435,N_43058,N_43677);
nand U44436 (N_44436,N_43529,N_43500);
or U44437 (N_44437,N_43861,N_43282);
nand U44438 (N_44438,N_43879,N_43771);
nor U44439 (N_44439,N_43350,N_43347);
or U44440 (N_44440,N_43485,N_43466);
xnor U44441 (N_44441,N_43142,N_43836);
xnor U44442 (N_44442,N_43584,N_43558);
nand U44443 (N_44443,N_43917,N_43524);
nor U44444 (N_44444,N_43864,N_43377);
xnor U44445 (N_44445,N_43275,N_43598);
nor U44446 (N_44446,N_43384,N_43840);
xnor U44447 (N_44447,N_43184,N_43380);
or U44448 (N_44448,N_43438,N_43916);
xor U44449 (N_44449,N_43680,N_43234);
nand U44450 (N_44450,N_43878,N_43230);
nand U44451 (N_44451,N_43870,N_43769);
nand U44452 (N_44452,N_43470,N_43188);
or U44453 (N_44453,N_43248,N_43740);
xnor U44454 (N_44454,N_43464,N_43932);
and U44455 (N_44455,N_43672,N_43521);
and U44456 (N_44456,N_43643,N_43579);
or U44457 (N_44457,N_43577,N_43127);
or U44458 (N_44458,N_43023,N_43876);
xnor U44459 (N_44459,N_43539,N_43927);
nand U44460 (N_44460,N_43739,N_43120);
nand U44461 (N_44461,N_43691,N_43849);
nand U44462 (N_44462,N_43352,N_43193);
xnor U44463 (N_44463,N_43624,N_43975);
or U44464 (N_44464,N_43304,N_43908);
or U44465 (N_44465,N_43823,N_43798);
or U44466 (N_44466,N_43225,N_43763);
xor U44467 (N_44467,N_43137,N_43249);
nand U44468 (N_44468,N_43117,N_43152);
and U44469 (N_44469,N_43810,N_43938);
or U44470 (N_44470,N_43904,N_43841);
nand U44471 (N_44471,N_43551,N_43455);
xnor U44472 (N_44472,N_43599,N_43918);
nand U44473 (N_44473,N_43844,N_43086);
nand U44474 (N_44474,N_43656,N_43345);
nor U44475 (N_44475,N_43069,N_43126);
nor U44476 (N_44476,N_43596,N_43959);
or U44477 (N_44477,N_43305,N_43253);
nand U44478 (N_44478,N_43991,N_43092);
or U44479 (N_44479,N_43061,N_43440);
xnor U44480 (N_44480,N_43615,N_43210);
nor U44481 (N_44481,N_43896,N_43886);
nor U44482 (N_44482,N_43363,N_43930);
and U44483 (N_44483,N_43062,N_43797);
nor U44484 (N_44484,N_43735,N_43578);
nand U44485 (N_44485,N_43947,N_43134);
nand U44486 (N_44486,N_43785,N_43800);
and U44487 (N_44487,N_43337,N_43123);
nand U44488 (N_44488,N_43055,N_43526);
nor U44489 (N_44489,N_43216,N_43992);
or U44490 (N_44490,N_43168,N_43601);
nand U44491 (N_44491,N_43899,N_43247);
and U44492 (N_44492,N_43665,N_43617);
nand U44493 (N_44493,N_43368,N_43161);
xor U44494 (N_44494,N_43147,N_43902);
or U44495 (N_44495,N_43900,N_43979);
nand U44496 (N_44496,N_43166,N_43506);
and U44497 (N_44497,N_43439,N_43792);
or U44498 (N_44498,N_43654,N_43758);
and U44499 (N_44499,N_43000,N_43075);
nand U44500 (N_44500,N_43865,N_43023);
xor U44501 (N_44501,N_43267,N_43425);
nand U44502 (N_44502,N_43620,N_43133);
xor U44503 (N_44503,N_43657,N_43407);
and U44504 (N_44504,N_43887,N_43453);
xnor U44505 (N_44505,N_43149,N_43613);
and U44506 (N_44506,N_43129,N_43582);
and U44507 (N_44507,N_43523,N_43600);
or U44508 (N_44508,N_43396,N_43169);
or U44509 (N_44509,N_43784,N_43570);
or U44510 (N_44510,N_43855,N_43863);
or U44511 (N_44511,N_43940,N_43775);
or U44512 (N_44512,N_43454,N_43825);
xnor U44513 (N_44513,N_43764,N_43543);
nor U44514 (N_44514,N_43621,N_43998);
nand U44515 (N_44515,N_43066,N_43138);
xor U44516 (N_44516,N_43797,N_43358);
nand U44517 (N_44517,N_43594,N_43272);
or U44518 (N_44518,N_43241,N_43933);
and U44519 (N_44519,N_43862,N_43046);
or U44520 (N_44520,N_43845,N_43398);
xnor U44521 (N_44521,N_43914,N_43334);
nand U44522 (N_44522,N_43773,N_43913);
nand U44523 (N_44523,N_43677,N_43623);
and U44524 (N_44524,N_43742,N_43318);
nor U44525 (N_44525,N_43937,N_43336);
or U44526 (N_44526,N_43285,N_43422);
xor U44527 (N_44527,N_43004,N_43099);
and U44528 (N_44528,N_43665,N_43782);
or U44529 (N_44529,N_43932,N_43792);
and U44530 (N_44530,N_43486,N_43347);
nor U44531 (N_44531,N_43448,N_43059);
nor U44532 (N_44532,N_43554,N_43008);
or U44533 (N_44533,N_43865,N_43192);
or U44534 (N_44534,N_43556,N_43223);
nor U44535 (N_44535,N_43967,N_43383);
nor U44536 (N_44536,N_43793,N_43875);
xor U44537 (N_44537,N_43298,N_43590);
and U44538 (N_44538,N_43612,N_43968);
nand U44539 (N_44539,N_43376,N_43798);
nor U44540 (N_44540,N_43379,N_43313);
or U44541 (N_44541,N_43150,N_43292);
and U44542 (N_44542,N_43055,N_43305);
xnor U44543 (N_44543,N_43050,N_43259);
or U44544 (N_44544,N_43379,N_43023);
nor U44545 (N_44545,N_43079,N_43248);
or U44546 (N_44546,N_43603,N_43548);
nor U44547 (N_44547,N_43193,N_43820);
nand U44548 (N_44548,N_43253,N_43442);
nor U44549 (N_44549,N_43599,N_43910);
nor U44550 (N_44550,N_43525,N_43632);
or U44551 (N_44551,N_43163,N_43715);
and U44552 (N_44552,N_43561,N_43921);
xor U44553 (N_44553,N_43815,N_43551);
xnor U44554 (N_44554,N_43973,N_43652);
and U44555 (N_44555,N_43908,N_43694);
or U44556 (N_44556,N_43696,N_43425);
or U44557 (N_44557,N_43545,N_43275);
nor U44558 (N_44558,N_43737,N_43985);
or U44559 (N_44559,N_43914,N_43567);
and U44560 (N_44560,N_43838,N_43705);
xor U44561 (N_44561,N_43061,N_43828);
or U44562 (N_44562,N_43115,N_43483);
nand U44563 (N_44563,N_43788,N_43716);
xnor U44564 (N_44564,N_43369,N_43502);
nor U44565 (N_44565,N_43180,N_43987);
nand U44566 (N_44566,N_43822,N_43196);
xnor U44567 (N_44567,N_43762,N_43418);
nor U44568 (N_44568,N_43718,N_43138);
or U44569 (N_44569,N_43381,N_43948);
nand U44570 (N_44570,N_43414,N_43581);
and U44571 (N_44571,N_43076,N_43891);
or U44572 (N_44572,N_43971,N_43521);
nand U44573 (N_44573,N_43907,N_43185);
or U44574 (N_44574,N_43446,N_43698);
nor U44575 (N_44575,N_43526,N_43620);
and U44576 (N_44576,N_43671,N_43730);
or U44577 (N_44577,N_43176,N_43777);
and U44578 (N_44578,N_43984,N_43546);
nand U44579 (N_44579,N_43355,N_43233);
or U44580 (N_44580,N_43999,N_43693);
and U44581 (N_44581,N_43344,N_43961);
and U44582 (N_44582,N_43656,N_43349);
and U44583 (N_44583,N_43812,N_43458);
and U44584 (N_44584,N_43336,N_43329);
or U44585 (N_44585,N_43831,N_43177);
and U44586 (N_44586,N_43374,N_43352);
or U44587 (N_44587,N_43227,N_43427);
nor U44588 (N_44588,N_43680,N_43329);
nand U44589 (N_44589,N_43496,N_43708);
nor U44590 (N_44590,N_43337,N_43520);
xor U44591 (N_44591,N_43083,N_43164);
nor U44592 (N_44592,N_43173,N_43047);
or U44593 (N_44593,N_43226,N_43254);
and U44594 (N_44594,N_43735,N_43374);
and U44595 (N_44595,N_43249,N_43638);
nand U44596 (N_44596,N_43655,N_43035);
or U44597 (N_44597,N_43666,N_43762);
or U44598 (N_44598,N_43322,N_43139);
nor U44599 (N_44599,N_43167,N_43731);
and U44600 (N_44600,N_43900,N_43770);
or U44601 (N_44601,N_43399,N_43831);
and U44602 (N_44602,N_43050,N_43513);
nor U44603 (N_44603,N_43578,N_43288);
xnor U44604 (N_44604,N_43426,N_43374);
xnor U44605 (N_44605,N_43540,N_43442);
nor U44606 (N_44606,N_43695,N_43730);
or U44607 (N_44607,N_43711,N_43325);
xor U44608 (N_44608,N_43718,N_43507);
or U44609 (N_44609,N_43236,N_43858);
and U44610 (N_44610,N_43885,N_43137);
and U44611 (N_44611,N_43161,N_43507);
and U44612 (N_44612,N_43153,N_43417);
nand U44613 (N_44613,N_43572,N_43690);
nor U44614 (N_44614,N_43174,N_43273);
nand U44615 (N_44615,N_43188,N_43051);
or U44616 (N_44616,N_43225,N_43610);
or U44617 (N_44617,N_43897,N_43289);
xor U44618 (N_44618,N_43252,N_43024);
or U44619 (N_44619,N_43257,N_43006);
nor U44620 (N_44620,N_43856,N_43204);
nor U44621 (N_44621,N_43176,N_43363);
nand U44622 (N_44622,N_43990,N_43101);
nor U44623 (N_44623,N_43845,N_43425);
nor U44624 (N_44624,N_43051,N_43924);
and U44625 (N_44625,N_43856,N_43057);
or U44626 (N_44626,N_43369,N_43530);
and U44627 (N_44627,N_43990,N_43755);
nand U44628 (N_44628,N_43411,N_43186);
nor U44629 (N_44629,N_43987,N_43474);
nor U44630 (N_44630,N_43573,N_43158);
or U44631 (N_44631,N_43667,N_43753);
and U44632 (N_44632,N_43250,N_43479);
nand U44633 (N_44633,N_43891,N_43198);
xor U44634 (N_44634,N_43039,N_43240);
nor U44635 (N_44635,N_43155,N_43087);
nand U44636 (N_44636,N_43473,N_43033);
or U44637 (N_44637,N_43294,N_43066);
and U44638 (N_44638,N_43834,N_43972);
nand U44639 (N_44639,N_43203,N_43154);
nand U44640 (N_44640,N_43088,N_43656);
nand U44641 (N_44641,N_43665,N_43040);
nand U44642 (N_44642,N_43240,N_43684);
and U44643 (N_44643,N_43632,N_43623);
nand U44644 (N_44644,N_43157,N_43997);
and U44645 (N_44645,N_43667,N_43898);
nor U44646 (N_44646,N_43568,N_43201);
and U44647 (N_44647,N_43954,N_43174);
nand U44648 (N_44648,N_43381,N_43979);
nand U44649 (N_44649,N_43792,N_43134);
and U44650 (N_44650,N_43335,N_43774);
nor U44651 (N_44651,N_43876,N_43083);
nor U44652 (N_44652,N_43300,N_43689);
xnor U44653 (N_44653,N_43377,N_43461);
nand U44654 (N_44654,N_43063,N_43803);
and U44655 (N_44655,N_43038,N_43095);
nor U44656 (N_44656,N_43528,N_43707);
xnor U44657 (N_44657,N_43667,N_43964);
and U44658 (N_44658,N_43503,N_43568);
xor U44659 (N_44659,N_43393,N_43301);
nor U44660 (N_44660,N_43738,N_43264);
or U44661 (N_44661,N_43051,N_43614);
and U44662 (N_44662,N_43124,N_43452);
xnor U44663 (N_44663,N_43106,N_43630);
and U44664 (N_44664,N_43038,N_43707);
and U44665 (N_44665,N_43791,N_43017);
nand U44666 (N_44666,N_43730,N_43267);
xor U44667 (N_44667,N_43338,N_43559);
nor U44668 (N_44668,N_43938,N_43833);
or U44669 (N_44669,N_43397,N_43119);
nor U44670 (N_44670,N_43565,N_43008);
nand U44671 (N_44671,N_43576,N_43435);
and U44672 (N_44672,N_43694,N_43568);
or U44673 (N_44673,N_43687,N_43913);
and U44674 (N_44674,N_43679,N_43164);
and U44675 (N_44675,N_43336,N_43171);
and U44676 (N_44676,N_43221,N_43079);
xor U44677 (N_44677,N_43332,N_43338);
and U44678 (N_44678,N_43517,N_43998);
nand U44679 (N_44679,N_43997,N_43602);
or U44680 (N_44680,N_43935,N_43907);
xnor U44681 (N_44681,N_43299,N_43241);
nand U44682 (N_44682,N_43157,N_43027);
xnor U44683 (N_44683,N_43206,N_43835);
nand U44684 (N_44684,N_43625,N_43378);
or U44685 (N_44685,N_43701,N_43681);
nor U44686 (N_44686,N_43631,N_43098);
xnor U44687 (N_44687,N_43289,N_43384);
or U44688 (N_44688,N_43582,N_43106);
or U44689 (N_44689,N_43792,N_43944);
nor U44690 (N_44690,N_43159,N_43290);
nor U44691 (N_44691,N_43898,N_43499);
nor U44692 (N_44692,N_43269,N_43986);
or U44693 (N_44693,N_43637,N_43191);
nand U44694 (N_44694,N_43577,N_43997);
nand U44695 (N_44695,N_43183,N_43681);
or U44696 (N_44696,N_43355,N_43004);
nand U44697 (N_44697,N_43243,N_43771);
or U44698 (N_44698,N_43411,N_43888);
or U44699 (N_44699,N_43884,N_43182);
nand U44700 (N_44700,N_43918,N_43824);
xnor U44701 (N_44701,N_43270,N_43915);
nor U44702 (N_44702,N_43602,N_43285);
xnor U44703 (N_44703,N_43586,N_43329);
nand U44704 (N_44704,N_43745,N_43538);
nor U44705 (N_44705,N_43856,N_43058);
and U44706 (N_44706,N_43727,N_43305);
nor U44707 (N_44707,N_43156,N_43638);
xor U44708 (N_44708,N_43110,N_43573);
or U44709 (N_44709,N_43709,N_43542);
nand U44710 (N_44710,N_43664,N_43195);
nor U44711 (N_44711,N_43752,N_43244);
and U44712 (N_44712,N_43312,N_43785);
nor U44713 (N_44713,N_43466,N_43243);
and U44714 (N_44714,N_43390,N_43799);
nand U44715 (N_44715,N_43005,N_43869);
xor U44716 (N_44716,N_43170,N_43520);
xor U44717 (N_44717,N_43392,N_43992);
and U44718 (N_44718,N_43735,N_43132);
and U44719 (N_44719,N_43383,N_43696);
nor U44720 (N_44720,N_43484,N_43028);
and U44721 (N_44721,N_43680,N_43936);
and U44722 (N_44722,N_43279,N_43499);
or U44723 (N_44723,N_43194,N_43068);
nor U44724 (N_44724,N_43386,N_43355);
xnor U44725 (N_44725,N_43187,N_43367);
nand U44726 (N_44726,N_43589,N_43400);
xnor U44727 (N_44727,N_43811,N_43969);
and U44728 (N_44728,N_43379,N_43857);
and U44729 (N_44729,N_43577,N_43317);
xnor U44730 (N_44730,N_43702,N_43160);
or U44731 (N_44731,N_43745,N_43236);
xor U44732 (N_44732,N_43483,N_43145);
xnor U44733 (N_44733,N_43387,N_43463);
nor U44734 (N_44734,N_43018,N_43462);
nor U44735 (N_44735,N_43604,N_43413);
nand U44736 (N_44736,N_43832,N_43014);
and U44737 (N_44737,N_43403,N_43341);
nor U44738 (N_44738,N_43993,N_43266);
nor U44739 (N_44739,N_43540,N_43777);
or U44740 (N_44740,N_43249,N_43241);
and U44741 (N_44741,N_43026,N_43430);
nand U44742 (N_44742,N_43259,N_43150);
xor U44743 (N_44743,N_43537,N_43541);
nor U44744 (N_44744,N_43256,N_43794);
or U44745 (N_44745,N_43956,N_43388);
nand U44746 (N_44746,N_43970,N_43039);
nand U44747 (N_44747,N_43866,N_43843);
nor U44748 (N_44748,N_43090,N_43946);
or U44749 (N_44749,N_43889,N_43327);
and U44750 (N_44750,N_43002,N_43635);
nand U44751 (N_44751,N_43290,N_43665);
nor U44752 (N_44752,N_43499,N_43937);
nor U44753 (N_44753,N_43174,N_43069);
nor U44754 (N_44754,N_43387,N_43672);
and U44755 (N_44755,N_43255,N_43742);
or U44756 (N_44756,N_43095,N_43567);
nor U44757 (N_44757,N_43945,N_43392);
xnor U44758 (N_44758,N_43573,N_43328);
and U44759 (N_44759,N_43105,N_43141);
nand U44760 (N_44760,N_43971,N_43257);
or U44761 (N_44761,N_43270,N_43893);
nor U44762 (N_44762,N_43372,N_43321);
nand U44763 (N_44763,N_43777,N_43377);
xnor U44764 (N_44764,N_43003,N_43833);
xnor U44765 (N_44765,N_43327,N_43657);
xor U44766 (N_44766,N_43734,N_43178);
xnor U44767 (N_44767,N_43381,N_43356);
or U44768 (N_44768,N_43095,N_43788);
nor U44769 (N_44769,N_43592,N_43167);
nor U44770 (N_44770,N_43272,N_43616);
and U44771 (N_44771,N_43639,N_43844);
or U44772 (N_44772,N_43504,N_43695);
nand U44773 (N_44773,N_43317,N_43183);
and U44774 (N_44774,N_43249,N_43164);
and U44775 (N_44775,N_43931,N_43225);
xnor U44776 (N_44776,N_43308,N_43491);
and U44777 (N_44777,N_43017,N_43357);
xor U44778 (N_44778,N_43118,N_43930);
or U44779 (N_44779,N_43405,N_43314);
nand U44780 (N_44780,N_43377,N_43824);
or U44781 (N_44781,N_43636,N_43112);
nor U44782 (N_44782,N_43418,N_43360);
nand U44783 (N_44783,N_43510,N_43667);
nor U44784 (N_44784,N_43592,N_43166);
and U44785 (N_44785,N_43936,N_43611);
nor U44786 (N_44786,N_43326,N_43194);
and U44787 (N_44787,N_43569,N_43031);
nor U44788 (N_44788,N_43340,N_43800);
or U44789 (N_44789,N_43207,N_43290);
nor U44790 (N_44790,N_43640,N_43558);
nor U44791 (N_44791,N_43259,N_43762);
xor U44792 (N_44792,N_43756,N_43471);
nor U44793 (N_44793,N_43509,N_43939);
nor U44794 (N_44794,N_43814,N_43790);
nand U44795 (N_44795,N_43940,N_43566);
or U44796 (N_44796,N_43223,N_43606);
and U44797 (N_44797,N_43270,N_43484);
nand U44798 (N_44798,N_43094,N_43661);
and U44799 (N_44799,N_43088,N_43112);
xnor U44800 (N_44800,N_43330,N_43736);
or U44801 (N_44801,N_43807,N_43727);
and U44802 (N_44802,N_43162,N_43429);
or U44803 (N_44803,N_43694,N_43400);
xnor U44804 (N_44804,N_43405,N_43489);
nor U44805 (N_44805,N_43549,N_43940);
nand U44806 (N_44806,N_43249,N_43299);
and U44807 (N_44807,N_43788,N_43384);
nor U44808 (N_44808,N_43285,N_43560);
xnor U44809 (N_44809,N_43498,N_43446);
nor U44810 (N_44810,N_43154,N_43979);
nand U44811 (N_44811,N_43306,N_43962);
xor U44812 (N_44812,N_43155,N_43551);
nor U44813 (N_44813,N_43109,N_43459);
or U44814 (N_44814,N_43306,N_43264);
or U44815 (N_44815,N_43099,N_43589);
or U44816 (N_44816,N_43107,N_43681);
nand U44817 (N_44817,N_43447,N_43279);
or U44818 (N_44818,N_43556,N_43915);
nor U44819 (N_44819,N_43459,N_43129);
xnor U44820 (N_44820,N_43901,N_43700);
nand U44821 (N_44821,N_43280,N_43513);
nand U44822 (N_44822,N_43586,N_43457);
xnor U44823 (N_44823,N_43975,N_43848);
and U44824 (N_44824,N_43105,N_43293);
nand U44825 (N_44825,N_43764,N_43419);
xnor U44826 (N_44826,N_43470,N_43953);
and U44827 (N_44827,N_43386,N_43558);
xnor U44828 (N_44828,N_43873,N_43872);
or U44829 (N_44829,N_43809,N_43493);
or U44830 (N_44830,N_43749,N_43825);
or U44831 (N_44831,N_43260,N_43646);
nand U44832 (N_44832,N_43295,N_43163);
or U44833 (N_44833,N_43027,N_43017);
and U44834 (N_44834,N_43518,N_43844);
nand U44835 (N_44835,N_43870,N_43847);
or U44836 (N_44836,N_43091,N_43782);
xnor U44837 (N_44837,N_43319,N_43889);
or U44838 (N_44838,N_43892,N_43448);
or U44839 (N_44839,N_43310,N_43747);
or U44840 (N_44840,N_43219,N_43949);
nor U44841 (N_44841,N_43170,N_43110);
xor U44842 (N_44842,N_43548,N_43833);
xnor U44843 (N_44843,N_43167,N_43620);
nand U44844 (N_44844,N_43351,N_43164);
nor U44845 (N_44845,N_43792,N_43355);
and U44846 (N_44846,N_43921,N_43747);
nor U44847 (N_44847,N_43155,N_43419);
nor U44848 (N_44848,N_43724,N_43759);
nand U44849 (N_44849,N_43551,N_43884);
xnor U44850 (N_44850,N_43214,N_43846);
xor U44851 (N_44851,N_43528,N_43993);
nor U44852 (N_44852,N_43336,N_43107);
and U44853 (N_44853,N_43308,N_43699);
nand U44854 (N_44854,N_43111,N_43497);
xor U44855 (N_44855,N_43118,N_43218);
xor U44856 (N_44856,N_43050,N_43566);
nand U44857 (N_44857,N_43616,N_43309);
nor U44858 (N_44858,N_43615,N_43064);
nor U44859 (N_44859,N_43708,N_43148);
or U44860 (N_44860,N_43586,N_43680);
nor U44861 (N_44861,N_43895,N_43729);
xor U44862 (N_44862,N_43791,N_43578);
xor U44863 (N_44863,N_43781,N_43654);
or U44864 (N_44864,N_43485,N_43185);
nand U44865 (N_44865,N_43368,N_43141);
and U44866 (N_44866,N_43429,N_43699);
nor U44867 (N_44867,N_43049,N_43475);
nor U44868 (N_44868,N_43296,N_43452);
nand U44869 (N_44869,N_43963,N_43270);
nor U44870 (N_44870,N_43314,N_43686);
nand U44871 (N_44871,N_43834,N_43198);
nor U44872 (N_44872,N_43583,N_43669);
or U44873 (N_44873,N_43620,N_43464);
or U44874 (N_44874,N_43581,N_43355);
or U44875 (N_44875,N_43820,N_43843);
nor U44876 (N_44876,N_43107,N_43248);
xnor U44877 (N_44877,N_43592,N_43191);
xnor U44878 (N_44878,N_43569,N_43103);
xnor U44879 (N_44879,N_43955,N_43728);
nand U44880 (N_44880,N_43876,N_43807);
nor U44881 (N_44881,N_43434,N_43267);
nand U44882 (N_44882,N_43714,N_43444);
nand U44883 (N_44883,N_43738,N_43416);
xnor U44884 (N_44884,N_43398,N_43660);
or U44885 (N_44885,N_43243,N_43443);
nor U44886 (N_44886,N_43303,N_43386);
nor U44887 (N_44887,N_43141,N_43460);
nand U44888 (N_44888,N_43642,N_43886);
nand U44889 (N_44889,N_43208,N_43977);
nor U44890 (N_44890,N_43756,N_43828);
nand U44891 (N_44891,N_43698,N_43083);
and U44892 (N_44892,N_43528,N_43045);
or U44893 (N_44893,N_43816,N_43395);
xor U44894 (N_44894,N_43136,N_43243);
and U44895 (N_44895,N_43152,N_43976);
nor U44896 (N_44896,N_43063,N_43533);
nand U44897 (N_44897,N_43724,N_43211);
or U44898 (N_44898,N_43555,N_43429);
nor U44899 (N_44899,N_43211,N_43663);
xnor U44900 (N_44900,N_43139,N_43292);
nand U44901 (N_44901,N_43267,N_43705);
or U44902 (N_44902,N_43217,N_43893);
and U44903 (N_44903,N_43266,N_43058);
or U44904 (N_44904,N_43048,N_43554);
nor U44905 (N_44905,N_43910,N_43125);
xor U44906 (N_44906,N_43298,N_43338);
and U44907 (N_44907,N_43370,N_43691);
xor U44908 (N_44908,N_43536,N_43662);
or U44909 (N_44909,N_43321,N_43864);
and U44910 (N_44910,N_43933,N_43811);
or U44911 (N_44911,N_43476,N_43981);
nor U44912 (N_44912,N_43197,N_43113);
or U44913 (N_44913,N_43922,N_43645);
xnor U44914 (N_44914,N_43728,N_43412);
nand U44915 (N_44915,N_43951,N_43040);
nor U44916 (N_44916,N_43867,N_43434);
xnor U44917 (N_44917,N_43708,N_43924);
nand U44918 (N_44918,N_43172,N_43807);
or U44919 (N_44919,N_43806,N_43033);
nor U44920 (N_44920,N_43124,N_43294);
nor U44921 (N_44921,N_43696,N_43492);
xnor U44922 (N_44922,N_43266,N_43013);
xnor U44923 (N_44923,N_43121,N_43209);
nor U44924 (N_44924,N_43597,N_43693);
and U44925 (N_44925,N_43221,N_43874);
and U44926 (N_44926,N_43513,N_43773);
or U44927 (N_44927,N_43166,N_43543);
and U44928 (N_44928,N_43154,N_43409);
and U44929 (N_44929,N_43439,N_43910);
and U44930 (N_44930,N_43207,N_43512);
nand U44931 (N_44931,N_43608,N_43205);
nand U44932 (N_44932,N_43497,N_43293);
nand U44933 (N_44933,N_43127,N_43540);
xor U44934 (N_44934,N_43834,N_43098);
and U44935 (N_44935,N_43665,N_43620);
or U44936 (N_44936,N_43418,N_43413);
nor U44937 (N_44937,N_43140,N_43703);
nor U44938 (N_44938,N_43476,N_43158);
and U44939 (N_44939,N_43491,N_43392);
and U44940 (N_44940,N_43733,N_43148);
xor U44941 (N_44941,N_43041,N_43755);
and U44942 (N_44942,N_43353,N_43082);
or U44943 (N_44943,N_43704,N_43681);
and U44944 (N_44944,N_43150,N_43023);
or U44945 (N_44945,N_43184,N_43995);
nand U44946 (N_44946,N_43565,N_43646);
or U44947 (N_44947,N_43275,N_43334);
nand U44948 (N_44948,N_43828,N_43740);
nand U44949 (N_44949,N_43055,N_43428);
or U44950 (N_44950,N_43812,N_43678);
nand U44951 (N_44951,N_43394,N_43799);
xnor U44952 (N_44952,N_43122,N_43656);
and U44953 (N_44953,N_43255,N_43539);
or U44954 (N_44954,N_43287,N_43885);
nor U44955 (N_44955,N_43643,N_43934);
xor U44956 (N_44956,N_43634,N_43933);
or U44957 (N_44957,N_43292,N_43660);
or U44958 (N_44958,N_43862,N_43284);
or U44959 (N_44959,N_43280,N_43255);
nand U44960 (N_44960,N_43246,N_43420);
nor U44961 (N_44961,N_43382,N_43639);
nor U44962 (N_44962,N_43724,N_43969);
nand U44963 (N_44963,N_43071,N_43844);
and U44964 (N_44964,N_43648,N_43697);
nand U44965 (N_44965,N_43791,N_43675);
nand U44966 (N_44966,N_43559,N_43000);
or U44967 (N_44967,N_43123,N_43901);
or U44968 (N_44968,N_43464,N_43057);
xor U44969 (N_44969,N_43713,N_43819);
nor U44970 (N_44970,N_43087,N_43118);
and U44971 (N_44971,N_43036,N_43958);
xnor U44972 (N_44972,N_43471,N_43570);
nand U44973 (N_44973,N_43884,N_43747);
and U44974 (N_44974,N_43090,N_43047);
and U44975 (N_44975,N_43433,N_43825);
nor U44976 (N_44976,N_43928,N_43779);
nand U44977 (N_44977,N_43794,N_43468);
xor U44978 (N_44978,N_43932,N_43415);
or U44979 (N_44979,N_43669,N_43398);
or U44980 (N_44980,N_43007,N_43241);
nand U44981 (N_44981,N_43488,N_43237);
and U44982 (N_44982,N_43415,N_43952);
nor U44983 (N_44983,N_43202,N_43848);
or U44984 (N_44984,N_43983,N_43927);
or U44985 (N_44985,N_43500,N_43162);
nand U44986 (N_44986,N_43950,N_43378);
or U44987 (N_44987,N_43133,N_43352);
nand U44988 (N_44988,N_43232,N_43505);
nand U44989 (N_44989,N_43782,N_43070);
nor U44990 (N_44990,N_43167,N_43705);
nand U44991 (N_44991,N_43590,N_43620);
and U44992 (N_44992,N_43304,N_43740);
and U44993 (N_44993,N_43871,N_43123);
or U44994 (N_44994,N_43987,N_43046);
nor U44995 (N_44995,N_43507,N_43494);
nor U44996 (N_44996,N_43713,N_43562);
nor U44997 (N_44997,N_43507,N_43426);
nor U44998 (N_44998,N_43375,N_43230);
xor U44999 (N_44999,N_43239,N_43074);
and U45000 (N_45000,N_44105,N_44248);
or U45001 (N_45001,N_44309,N_44498);
nor U45002 (N_45002,N_44376,N_44571);
nand U45003 (N_45003,N_44136,N_44311);
xnor U45004 (N_45004,N_44403,N_44122);
or U45005 (N_45005,N_44470,N_44664);
and U45006 (N_45006,N_44493,N_44924);
and U45007 (N_45007,N_44567,N_44942);
and U45008 (N_45008,N_44169,N_44050);
xnor U45009 (N_45009,N_44944,N_44460);
nand U45010 (N_45010,N_44568,N_44476);
nor U45011 (N_45011,N_44831,N_44905);
xor U45012 (N_45012,N_44613,N_44322);
xnor U45013 (N_45013,N_44286,N_44890);
nand U45014 (N_45014,N_44900,N_44653);
or U45015 (N_45015,N_44380,N_44519);
nor U45016 (N_45016,N_44092,N_44920);
or U45017 (N_45017,N_44267,N_44189);
nor U45018 (N_45018,N_44795,N_44171);
nand U45019 (N_45019,N_44006,N_44149);
or U45020 (N_45020,N_44060,N_44718);
nand U45021 (N_45021,N_44885,N_44278);
nor U45022 (N_45022,N_44719,N_44360);
nor U45023 (N_45023,N_44875,N_44121);
xor U45024 (N_45024,N_44689,N_44855);
and U45025 (N_45025,N_44801,N_44787);
xnor U45026 (N_45026,N_44231,N_44504);
xor U45027 (N_45027,N_44912,N_44062);
xnor U45028 (N_45028,N_44454,N_44688);
nand U45029 (N_45029,N_44315,N_44760);
xor U45030 (N_45030,N_44997,N_44371);
and U45031 (N_45031,N_44984,N_44727);
nand U45032 (N_45032,N_44157,N_44946);
or U45033 (N_45033,N_44704,N_44937);
or U45034 (N_45034,N_44178,N_44536);
nand U45035 (N_45035,N_44343,N_44662);
or U45036 (N_45036,N_44175,N_44990);
xor U45037 (N_45037,N_44023,N_44177);
nand U45038 (N_45038,N_44538,N_44856);
nand U45039 (N_45039,N_44846,N_44680);
nand U45040 (N_45040,N_44115,N_44458);
nor U45041 (N_45041,N_44292,N_44180);
nand U45042 (N_45042,N_44008,N_44768);
and U45043 (N_45043,N_44707,N_44961);
nand U45044 (N_45044,N_44948,N_44409);
and U45045 (N_45045,N_44535,N_44017);
and U45046 (N_45046,N_44894,N_44245);
xnor U45047 (N_45047,N_44749,N_44414);
nand U45048 (N_45048,N_44508,N_44031);
nand U45049 (N_45049,N_44975,N_44636);
xnor U45050 (N_45050,N_44250,N_44648);
xnor U45051 (N_45051,N_44235,N_44287);
nor U45052 (N_45052,N_44802,N_44882);
nand U45053 (N_45053,N_44691,N_44510);
nand U45054 (N_45054,N_44502,N_44272);
nor U45055 (N_45055,N_44967,N_44066);
and U45056 (N_45056,N_44971,N_44428);
or U45057 (N_45057,N_44484,N_44154);
xor U45058 (N_45058,N_44084,N_44188);
nor U45059 (N_45059,N_44792,N_44308);
nor U45060 (N_45060,N_44716,N_44012);
nor U45061 (N_45061,N_44466,N_44911);
or U45062 (N_45062,N_44398,N_44399);
nor U45063 (N_45063,N_44133,N_44705);
or U45064 (N_45064,N_44572,N_44767);
nand U45065 (N_45065,N_44629,N_44110);
xor U45066 (N_45066,N_44165,N_44390);
or U45067 (N_45067,N_44565,N_44627);
xnor U45068 (N_45068,N_44268,N_44901);
nand U45069 (N_45069,N_44521,N_44317);
nand U45070 (N_45070,N_44677,N_44168);
nand U45071 (N_45071,N_44468,N_44367);
nor U45072 (N_45072,N_44104,N_44324);
xnor U45073 (N_45073,N_44093,N_44043);
and U45074 (N_45074,N_44439,N_44251);
nand U45075 (N_45075,N_44226,N_44126);
nand U45076 (N_45076,N_44918,N_44992);
xnor U45077 (N_45077,N_44858,N_44745);
and U45078 (N_45078,N_44152,N_44221);
and U45079 (N_45079,N_44878,N_44914);
nor U45080 (N_45080,N_44029,N_44254);
or U45081 (N_45081,N_44244,N_44580);
xnor U45082 (N_45082,N_44533,N_44981);
nor U45083 (N_45083,N_44144,N_44353);
xnor U45084 (N_45084,N_44696,N_44947);
and U45085 (N_45085,N_44421,N_44926);
nor U45086 (N_45086,N_44182,N_44670);
xor U45087 (N_45087,N_44714,N_44257);
or U45088 (N_45088,N_44897,N_44085);
nand U45089 (N_45089,N_44530,N_44055);
nor U45090 (N_45090,N_44892,N_44069);
and U45091 (N_45091,N_44462,N_44668);
or U45092 (N_45092,N_44095,N_44422);
and U45093 (N_45093,N_44867,N_44620);
nor U45094 (N_45094,N_44176,N_44447);
xor U45095 (N_45095,N_44024,N_44067);
nand U45096 (N_45096,N_44578,N_44628);
and U45097 (N_45097,N_44262,N_44819);
nor U45098 (N_45098,N_44539,N_44193);
or U45099 (N_45099,N_44200,N_44326);
nand U45100 (N_45100,N_44587,N_44495);
or U45101 (N_45101,N_44952,N_44228);
or U45102 (N_45102,N_44637,N_44734);
nand U45103 (N_45103,N_44469,N_44475);
nand U45104 (N_45104,N_44387,N_44233);
nand U45105 (N_45105,N_44966,N_44542);
xnor U45106 (N_45106,N_44998,N_44298);
or U45107 (N_45107,N_44342,N_44238);
xnor U45108 (N_45108,N_44687,N_44204);
nand U45109 (N_45109,N_44239,N_44265);
xor U45110 (N_45110,N_44805,N_44640);
nand U45111 (N_45111,N_44957,N_44863);
nand U45112 (N_45112,N_44145,N_44609);
and U45113 (N_45113,N_44988,N_44583);
xnor U45114 (N_45114,N_44592,N_44415);
or U45115 (N_45115,N_44868,N_44137);
nand U45116 (N_45116,N_44797,N_44979);
or U45117 (N_45117,N_44426,N_44321);
xor U45118 (N_45118,N_44903,N_44219);
xor U45119 (N_45119,N_44207,N_44969);
or U45120 (N_45120,N_44773,N_44757);
xor U45121 (N_45121,N_44370,N_44543);
or U45122 (N_45122,N_44974,N_44035);
xnor U45123 (N_45123,N_44943,N_44853);
nor U45124 (N_45124,N_44635,N_44220);
and U45125 (N_45125,N_44611,N_44199);
and U45126 (N_45126,N_44070,N_44741);
nor U45127 (N_45127,N_44005,N_44289);
xor U45128 (N_45128,N_44985,N_44318);
xor U45129 (N_45129,N_44646,N_44818);
or U45130 (N_45130,N_44486,N_44036);
xor U45131 (N_45131,N_44086,N_44927);
and U45132 (N_45132,N_44541,N_44759);
nand U45133 (N_45133,N_44700,N_44123);
xor U45134 (N_45134,N_44563,N_44266);
and U45135 (N_45135,N_44134,N_44162);
xnor U45136 (N_45136,N_44817,N_44340);
or U45137 (N_45137,N_44425,N_44437);
and U45138 (N_45138,N_44566,N_44617);
nor U45139 (N_45139,N_44595,N_44755);
nor U45140 (N_45140,N_44579,N_44828);
nor U45141 (N_45141,N_44044,N_44550);
and U45142 (N_45142,N_44391,N_44601);
nor U45143 (N_45143,N_44939,N_44701);
nand U45144 (N_45144,N_44275,N_44494);
nand U45145 (N_45145,N_44778,N_44660);
or U45146 (N_45146,N_44408,N_44665);
nand U45147 (N_45147,N_44365,N_44283);
xnor U45148 (N_45148,N_44273,N_44499);
xnor U45149 (N_45149,N_44602,N_44038);
or U45150 (N_45150,N_44384,N_44088);
or U45151 (N_45151,N_44872,N_44940);
xnor U45152 (N_45152,N_44980,N_44632);
xor U45153 (N_45153,N_44127,N_44314);
xor U45154 (N_45154,N_44016,N_44658);
xor U45155 (N_45155,N_44837,N_44222);
nand U45156 (N_45156,N_44895,N_44744);
or U45157 (N_45157,N_44747,N_44369);
or U45158 (N_45158,N_44547,N_44101);
xor U45159 (N_45159,N_44335,N_44057);
or U45160 (N_45160,N_44090,N_44331);
nor U45161 (N_45161,N_44772,N_44337);
or U45162 (N_45162,N_44724,N_44783);
and U45163 (N_45163,N_44752,N_44375);
nor U45164 (N_45164,N_44955,N_44982);
nor U45165 (N_45165,N_44514,N_44206);
or U45166 (N_45166,N_44246,N_44652);
nand U45167 (N_45167,N_44896,N_44166);
or U45168 (N_45168,N_44047,N_44443);
xor U45169 (N_45169,N_44794,N_44865);
nand U45170 (N_45170,N_44641,N_44811);
nand U45171 (N_45171,N_44382,N_44366);
nor U45172 (N_45172,N_44803,N_44009);
or U45173 (N_45173,N_44995,N_44761);
and U45174 (N_45174,N_44218,N_44401);
xor U45175 (N_45175,N_44255,N_44518);
nor U45176 (N_45176,N_44113,N_44781);
xnor U45177 (N_45177,N_44073,N_44270);
nand U45178 (N_45178,N_44294,N_44569);
nand U45179 (N_45179,N_44236,N_44779);
nor U45180 (N_45180,N_44622,N_44909);
xor U45181 (N_45181,N_44644,N_44065);
xnor U45182 (N_45182,N_44720,N_44333);
nand U45183 (N_45183,N_44715,N_44284);
or U45184 (N_45184,N_44312,N_44679);
or U45185 (N_45185,N_44824,N_44049);
and U45186 (N_45186,N_44798,N_44832);
and U45187 (N_45187,N_44293,N_44886);
nor U45188 (N_45188,N_44274,N_44938);
or U45189 (N_45189,N_44809,N_44509);
or U45190 (N_45190,N_44698,N_44970);
and U45191 (N_45191,N_44814,N_44338);
nor U45192 (N_45192,N_44842,N_44584);
xor U45193 (N_45193,N_44936,N_44028);
nand U45194 (N_45194,N_44156,N_44789);
and U45195 (N_45195,N_44790,N_44344);
or U45196 (N_45196,N_44537,N_44910);
nand U45197 (N_45197,N_44693,N_44445);
xor U45198 (N_45198,N_44515,N_44619);
or U45199 (N_45199,N_44516,N_44917);
nor U45200 (N_45200,N_44823,N_44280);
and U45201 (N_45201,N_44834,N_44501);
xnor U45202 (N_45202,N_44738,N_44022);
and U45203 (N_45203,N_44520,N_44851);
nand U45204 (N_45204,N_44276,N_44973);
xnor U45205 (N_45205,N_44013,N_44103);
nand U45206 (N_45206,N_44876,N_44362);
nor U45207 (N_45207,N_44585,N_44702);
or U45208 (N_45208,N_44960,N_44756);
nor U45209 (N_45209,N_44850,N_44167);
and U45210 (N_45210,N_44986,N_44135);
or U45211 (N_45211,N_44102,N_44812);
or U45212 (N_45212,N_44094,N_44183);
or U45213 (N_45213,N_44347,N_44302);
or U45214 (N_45214,N_44381,N_44746);
nor U45215 (N_45215,N_44002,N_44925);
and U45216 (N_45216,N_44379,N_44374);
and U45217 (N_45217,N_44305,N_44418);
nand U45218 (N_45218,N_44726,N_44051);
nand U45219 (N_45219,N_44319,N_44526);
xor U45220 (N_45220,N_44299,N_44954);
or U45221 (N_45221,N_44230,N_44849);
and U45222 (N_45222,N_44260,N_44096);
or U45223 (N_45223,N_44959,N_44109);
nor U45224 (N_45224,N_44810,N_44869);
xnor U45225 (N_45225,N_44800,N_44780);
and U45226 (N_45226,N_44282,N_44479);
nand U45227 (N_45227,N_44904,N_44082);
and U45228 (N_45228,N_44999,N_44929);
xnor U45229 (N_45229,N_44068,N_44461);
nor U45230 (N_45230,N_44225,N_44544);
and U45231 (N_45231,N_44359,N_44118);
xor U45232 (N_45232,N_44420,N_44131);
or U45233 (N_45233,N_44472,N_44777);
nand U45234 (N_45234,N_44642,N_44710);
nor U45235 (N_45235,N_44446,N_44160);
nand U45236 (N_45236,N_44643,N_44477);
and U45237 (N_45237,N_44116,N_44582);
or U45238 (N_45238,N_44813,N_44056);
and U45239 (N_45239,N_44424,N_44728);
nand U45240 (N_45240,N_44089,N_44593);
nand U45241 (N_45241,N_44623,N_44120);
or U45242 (N_45242,N_44291,N_44829);
and U45243 (N_45243,N_44913,N_44436);
xnor U45244 (N_45244,N_44108,N_44650);
nor U45245 (N_45245,N_44253,N_44406);
nor U45246 (N_45246,N_44610,N_44383);
xor U45247 (N_45247,N_44862,N_44368);
xnor U45248 (N_45248,N_44881,N_44192);
nand U45249 (N_45249,N_44405,N_44216);
and U45250 (N_45250,N_44467,N_44030);
nor U45251 (N_45251,N_44077,N_44258);
and U45252 (N_45252,N_44978,N_44155);
xor U45253 (N_45253,N_44843,N_44877);
nor U45254 (N_45254,N_44045,N_44923);
nand U45255 (N_45255,N_44485,N_44766);
nor U45256 (N_45256,N_44330,N_44932);
and U45257 (N_45257,N_44861,N_44143);
xnor U45258 (N_45258,N_44279,N_44612);
or U45259 (N_45259,N_44003,N_44483);
nand U45260 (N_45260,N_44296,N_44478);
or U45261 (N_45261,N_44751,N_44845);
xor U45262 (N_45262,N_44473,N_44889);
or U45263 (N_45263,N_44739,N_44796);
xnor U45264 (N_45264,N_44758,N_44722);
and U45265 (N_45265,N_44771,N_44032);
or U45266 (N_45266,N_44654,N_44673);
or U45267 (N_45267,N_44949,N_44667);
nor U45268 (N_45268,N_44329,N_44553);
and U45269 (N_45269,N_44708,N_44763);
or U45270 (N_45270,N_44935,N_44410);
or U45271 (N_45271,N_44211,N_44252);
or U45272 (N_45272,N_44874,N_44678);
or U45273 (N_45273,N_44634,N_44534);
xnor U45274 (N_45274,N_44395,N_44124);
and U45275 (N_45275,N_44586,N_44098);
or U45276 (N_45276,N_44898,N_44733);
nor U45277 (N_45277,N_44825,N_44442);
xnor U45278 (N_45278,N_44902,N_44576);
xor U45279 (N_45279,N_44474,N_44063);
or U45280 (N_45280,N_44799,N_44836);
xnor U45281 (N_45281,N_44240,N_44229);
or U45282 (N_45282,N_44179,N_44916);
xnor U45283 (N_45283,N_44378,N_44621);
xor U45284 (N_45284,N_44243,N_44709);
xor U45285 (N_45285,N_44463,N_44004);
nand U45286 (N_45286,N_44934,N_44804);
and U45287 (N_45287,N_44888,N_44532);
and U45288 (N_45288,N_44316,N_44455);
xnor U45289 (N_45289,N_44844,N_44271);
nand U45290 (N_45290,N_44392,N_44782);
nor U45291 (N_45291,N_44559,N_44857);
or U45292 (N_45292,N_44147,N_44764);
nor U45293 (N_45293,N_44683,N_44681);
xnor U45294 (N_45294,N_44697,N_44491);
or U45295 (N_45295,N_44775,N_44921);
or U45296 (N_45296,N_44968,N_44561);
xnor U45297 (N_45297,N_44300,N_44762);
xnor U45298 (N_45298,N_44020,N_44671);
and U45299 (N_45299,N_44651,N_44061);
nand U45300 (N_45300,N_44303,N_44481);
nor U45301 (N_45301,N_44841,N_44214);
nor U45302 (N_45302,N_44490,N_44721);
nand U45303 (N_45303,N_44033,N_44546);
nor U45304 (N_45304,N_44769,N_44564);
xor U45305 (N_45305,N_44560,N_44164);
and U45306 (N_45306,N_44806,N_44350);
nor U45307 (N_45307,N_44626,N_44264);
and U45308 (N_45308,N_44590,N_44972);
and U45309 (N_45309,N_44600,N_44416);
xor U45310 (N_45310,N_44599,N_44506);
nand U45311 (N_45311,N_44021,N_44125);
or U45312 (N_45312,N_44822,N_44552);
or U45313 (N_45313,N_44010,N_44489);
nand U45314 (N_45314,N_44459,N_44827);
nand U45315 (N_45315,N_44666,N_44996);
and U45316 (N_45316,N_44332,N_44977);
xnor U45317 (N_45317,N_44598,N_44840);
nand U45318 (N_45318,N_44991,N_44694);
nand U45319 (N_45319,N_44496,N_44551);
or U45320 (N_45320,N_44196,N_44336);
or U45321 (N_45321,N_44603,N_44548);
and U45322 (N_45322,N_44306,N_44743);
or U45323 (N_45323,N_44821,N_44776);
nand U45324 (N_45324,N_44633,N_44440);
nand U45325 (N_45325,N_44364,N_44432);
nand U45326 (N_45326,N_44647,N_44041);
nand U45327 (N_45327,N_44277,N_44173);
nor U45328 (N_45328,N_44549,N_44042);
nand U45329 (N_45329,N_44119,N_44618);
nor U45330 (N_45330,N_44419,N_44887);
xnor U45331 (N_45331,N_44497,N_44956);
or U45332 (N_45332,N_44018,N_44430);
and U45333 (N_45333,N_44994,N_44606);
xnor U45334 (N_45334,N_44815,N_44941);
nand U45335 (N_45335,N_44323,N_44597);
or U45336 (N_45336,N_44793,N_44488);
nor U45337 (N_45337,N_44893,N_44570);
nand U45338 (N_45338,N_44327,N_44356);
nand U45339 (N_45339,N_44983,N_44107);
or U45340 (N_45340,N_44608,N_44091);
or U45341 (N_45341,N_44736,N_44117);
and U45342 (N_45342,N_44731,N_44184);
nand U45343 (N_45343,N_44712,N_44181);
xnor U45344 (N_45344,N_44242,N_44607);
or U45345 (N_45345,N_44908,N_44989);
nor U45346 (N_45346,N_44674,N_44423);
and U45347 (N_45347,N_44907,N_44249);
or U45348 (N_45348,N_44269,N_44363);
nor U45349 (N_45349,N_44411,N_44596);
or U45350 (N_45350,N_44870,N_44163);
or U45351 (N_45351,N_44729,N_44774);
nor U45352 (N_45352,N_44449,N_44933);
nand U45353 (N_45353,N_44871,N_44128);
or U45354 (N_45354,N_44523,N_44019);
nor U45355 (N_45355,N_44659,N_44210);
nand U45356 (N_45356,N_44081,N_44099);
nor U45357 (N_45357,N_44754,N_44025);
and U45358 (N_45358,N_44993,N_44187);
nor U45359 (N_45359,N_44170,N_44281);
nand U45360 (N_45360,N_44034,N_44297);
xor U45361 (N_45361,N_44906,N_44361);
or U45362 (N_45362,N_44227,N_44786);
or U45363 (N_45363,N_44573,N_44682);
and U45364 (N_45364,N_44352,N_44208);
or U45365 (N_45365,N_44505,N_44394);
and U45366 (N_45366,N_44725,N_44026);
nor U45367 (N_45367,N_44373,N_44784);
nor U45368 (N_45368,N_44313,N_44295);
nor U45369 (N_45369,N_44638,N_44713);
or U45370 (N_45370,N_44465,N_44830);
nand U45371 (N_45371,N_44212,N_44675);
nor U45372 (N_45372,N_44385,N_44195);
or U45373 (N_45373,N_44431,N_44513);
xor U45374 (N_45374,N_44852,N_44883);
and U45375 (N_45375,N_44205,N_44039);
nor U45376 (N_45376,N_44672,N_44237);
xor U45377 (N_45377,N_44151,N_44232);
and U45378 (N_45378,N_44503,N_44826);
and U45379 (N_45379,N_44630,N_44075);
nor U45380 (N_45380,N_44854,N_44699);
xor U45381 (N_45381,N_44594,N_44146);
and U45382 (N_45382,N_44962,N_44148);
nor U45383 (N_45383,N_44690,N_44080);
nor U45384 (N_45384,N_44873,N_44076);
and U45385 (N_45385,N_44649,N_44788);
and U45386 (N_45386,N_44377,N_44037);
xor U45387 (N_45387,N_44304,N_44111);
xor U45388 (N_45388,N_44083,N_44457);
or U45389 (N_45389,N_44820,N_44150);
nor U45390 (N_45390,N_44577,N_44631);
and U45391 (N_45391,N_44290,N_44197);
nor U45392 (N_45392,N_44528,N_44656);
or U45393 (N_45393,N_44555,N_44000);
or U45394 (N_45394,N_44737,N_44866);
nor U45395 (N_45395,N_44346,N_44334);
xnor U45396 (N_45396,N_44046,N_44616);
nor U45397 (N_45397,N_44791,N_44615);
and U45398 (N_45398,N_44194,N_44357);
and U45399 (N_45399,N_44451,N_44404);
or U45400 (N_45400,N_44706,N_44388);
xnor U45401 (N_45401,N_44203,N_44138);
and U45402 (N_45402,N_44556,N_44015);
and U45403 (N_45403,N_44413,N_44161);
or U45404 (N_45404,N_44581,N_44011);
nor U45405 (N_45405,N_44557,N_44860);
nor U45406 (N_45406,N_44655,N_44201);
and U45407 (N_45407,N_44950,N_44159);
nand U45408 (N_45408,N_44429,N_44614);
nand U45409 (N_45409,N_44433,N_44190);
nand U45410 (N_45410,N_44345,N_44100);
nor U45411 (N_45411,N_44953,N_44574);
xnor U45412 (N_45412,N_44444,N_44964);
nor U45413 (N_45413,N_44864,N_44396);
xor U45414 (N_45414,N_44450,N_44339);
and U45415 (N_45415,N_44711,N_44393);
nor U45416 (N_45416,N_44464,N_44922);
and U45417 (N_45417,N_44217,N_44400);
nand U45418 (N_45418,N_44438,N_44141);
and U45419 (N_45419,N_44919,N_44072);
or U45420 (N_45420,N_44320,N_44604);
xor U45421 (N_45421,N_44527,N_44386);
nand U45422 (N_45422,N_44129,N_44965);
and U45423 (N_45423,N_44130,N_44723);
and U45424 (N_45424,N_44770,N_44328);
nand U45425 (N_45425,N_44517,N_44880);
and U45426 (N_45426,N_44692,N_44202);
or U45427 (N_45427,N_44976,N_44531);
nand U45428 (N_45428,N_44589,N_44562);
or U45429 (N_45429,N_44106,N_44835);
nor U45430 (N_45430,N_44052,N_44234);
nor U45431 (N_45431,N_44512,N_44676);
nand U45432 (N_45432,N_44301,N_44487);
nor U45433 (N_45433,N_44142,N_44372);
and U45434 (N_45434,N_44349,N_44213);
and U45435 (N_45435,N_44402,N_44750);
xor U45436 (N_45436,N_44285,N_44471);
nand U45437 (N_45437,N_44605,N_44735);
nand U45438 (N_45438,N_44007,N_44434);
xnor U45439 (N_45439,N_44307,N_44686);
and U45440 (N_45440,N_44951,N_44753);
nand U45441 (N_45441,N_44351,N_44198);
and U45442 (N_45442,N_44153,N_44669);
xor U45443 (N_45443,N_44412,N_44511);
nand U45444 (N_45444,N_44807,N_44247);
or U45445 (N_45445,N_44740,N_44074);
and U45446 (N_45446,N_44624,N_44808);
nor U45447 (N_45447,N_44891,N_44261);
or U45448 (N_45448,N_44915,N_44112);
or U45449 (N_45449,N_44453,N_44703);
xor U45450 (N_45450,N_44417,N_44931);
and U45451 (N_45451,N_44223,N_44158);
and U45452 (N_45452,N_44684,N_44040);
and U45453 (N_45453,N_44355,N_44174);
xnor U45454 (N_45454,N_44833,N_44838);
nand U45455 (N_45455,N_44078,N_44785);
and U45456 (N_45456,N_44054,N_44191);
xor U45457 (N_45457,N_44140,N_44879);
nor U45458 (N_45458,N_44097,N_44958);
nor U45459 (N_45459,N_44492,N_44456);
xor U45460 (N_45460,N_44087,N_44540);
nand U45461 (N_45461,N_44732,N_44558);
xnor U45462 (N_45462,N_44963,N_44507);
nand U45463 (N_45463,N_44930,N_44452);
xor U45464 (N_45464,N_44256,N_44209);
xor U45465 (N_45465,N_44987,N_44186);
nor U45466 (N_45466,N_44748,N_44064);
and U45467 (N_45467,N_44114,N_44348);
xor U45468 (N_45468,N_44816,N_44132);
nor U45469 (N_45469,N_44522,N_44407);
nand U45470 (N_45470,N_44685,N_44448);
nand U45471 (N_45471,N_44945,N_44441);
nor U45472 (N_45472,N_44730,N_44397);
and U45473 (N_45473,N_44027,N_44482);
nor U45474 (N_45474,N_44215,N_44625);
or U45475 (N_45475,N_44480,N_44742);
nor U45476 (N_45476,N_44657,N_44001);
or U45477 (N_45477,N_44765,N_44661);
or U45478 (N_45478,N_44224,N_44575);
xnor U45479 (N_45479,N_44847,N_44899);
xnor U45480 (N_45480,N_44139,N_44695);
xnor U45481 (N_45481,N_44325,N_44435);
nand U45482 (N_45482,N_44358,N_44053);
nand U45483 (N_45483,N_44354,N_44014);
nor U45484 (N_45484,N_44389,N_44663);
nand U45485 (N_45485,N_44545,N_44172);
and U45486 (N_45486,N_44645,N_44524);
nor U45487 (N_45487,N_44928,N_44554);
xor U45488 (N_45488,N_44263,N_44185);
xnor U45489 (N_45489,N_44525,N_44241);
or U45490 (N_45490,N_44859,N_44310);
nor U45491 (N_45491,N_44588,N_44427);
or U45492 (N_45492,N_44048,N_44717);
or U45493 (N_45493,N_44500,N_44341);
xnor U45494 (N_45494,N_44639,N_44259);
nor U45495 (N_45495,N_44059,N_44839);
nor U45496 (N_45496,N_44288,N_44058);
nor U45497 (N_45497,N_44591,N_44071);
xor U45498 (N_45498,N_44529,N_44848);
and U45499 (N_45499,N_44884,N_44079);
nor U45500 (N_45500,N_44935,N_44145);
xnor U45501 (N_45501,N_44848,N_44664);
xnor U45502 (N_45502,N_44105,N_44976);
nand U45503 (N_45503,N_44014,N_44705);
or U45504 (N_45504,N_44162,N_44020);
nand U45505 (N_45505,N_44526,N_44903);
and U45506 (N_45506,N_44731,N_44346);
nor U45507 (N_45507,N_44118,N_44578);
nand U45508 (N_45508,N_44256,N_44211);
nand U45509 (N_45509,N_44273,N_44000);
nand U45510 (N_45510,N_44227,N_44317);
xnor U45511 (N_45511,N_44563,N_44632);
nor U45512 (N_45512,N_44600,N_44971);
nor U45513 (N_45513,N_44072,N_44374);
and U45514 (N_45514,N_44635,N_44808);
xnor U45515 (N_45515,N_44829,N_44527);
or U45516 (N_45516,N_44420,N_44208);
nor U45517 (N_45517,N_44142,N_44949);
xor U45518 (N_45518,N_44562,N_44022);
or U45519 (N_45519,N_44380,N_44787);
nand U45520 (N_45520,N_44745,N_44238);
or U45521 (N_45521,N_44808,N_44703);
nor U45522 (N_45522,N_44682,N_44008);
nand U45523 (N_45523,N_44566,N_44007);
xor U45524 (N_45524,N_44039,N_44994);
nor U45525 (N_45525,N_44935,N_44710);
nor U45526 (N_45526,N_44206,N_44012);
nand U45527 (N_45527,N_44909,N_44315);
nand U45528 (N_45528,N_44217,N_44571);
xnor U45529 (N_45529,N_44900,N_44785);
nor U45530 (N_45530,N_44417,N_44500);
or U45531 (N_45531,N_44172,N_44600);
nand U45532 (N_45532,N_44935,N_44395);
or U45533 (N_45533,N_44650,N_44327);
and U45534 (N_45534,N_44534,N_44772);
and U45535 (N_45535,N_44577,N_44980);
nor U45536 (N_45536,N_44771,N_44760);
or U45537 (N_45537,N_44765,N_44082);
xnor U45538 (N_45538,N_44111,N_44406);
xor U45539 (N_45539,N_44840,N_44150);
and U45540 (N_45540,N_44708,N_44017);
nand U45541 (N_45541,N_44207,N_44552);
xnor U45542 (N_45542,N_44054,N_44669);
nor U45543 (N_45543,N_44853,N_44002);
nand U45544 (N_45544,N_44197,N_44888);
or U45545 (N_45545,N_44943,N_44082);
and U45546 (N_45546,N_44684,N_44530);
xnor U45547 (N_45547,N_44716,N_44618);
xor U45548 (N_45548,N_44004,N_44709);
and U45549 (N_45549,N_44475,N_44266);
nor U45550 (N_45550,N_44378,N_44140);
and U45551 (N_45551,N_44181,N_44084);
nand U45552 (N_45552,N_44834,N_44723);
and U45553 (N_45553,N_44175,N_44165);
or U45554 (N_45554,N_44004,N_44672);
nor U45555 (N_45555,N_44831,N_44862);
or U45556 (N_45556,N_44453,N_44818);
nor U45557 (N_45557,N_44965,N_44243);
xnor U45558 (N_45558,N_44804,N_44564);
nand U45559 (N_45559,N_44267,N_44565);
xnor U45560 (N_45560,N_44601,N_44683);
xnor U45561 (N_45561,N_44680,N_44686);
and U45562 (N_45562,N_44781,N_44260);
nand U45563 (N_45563,N_44960,N_44741);
or U45564 (N_45564,N_44152,N_44705);
and U45565 (N_45565,N_44072,N_44941);
nor U45566 (N_45566,N_44185,N_44174);
nor U45567 (N_45567,N_44789,N_44361);
and U45568 (N_45568,N_44263,N_44512);
nor U45569 (N_45569,N_44092,N_44298);
and U45570 (N_45570,N_44800,N_44221);
xnor U45571 (N_45571,N_44852,N_44119);
xnor U45572 (N_45572,N_44726,N_44171);
or U45573 (N_45573,N_44524,N_44427);
xor U45574 (N_45574,N_44888,N_44589);
nor U45575 (N_45575,N_44441,N_44461);
or U45576 (N_45576,N_44751,N_44318);
and U45577 (N_45577,N_44505,N_44667);
and U45578 (N_45578,N_44972,N_44373);
and U45579 (N_45579,N_44830,N_44610);
or U45580 (N_45580,N_44015,N_44740);
and U45581 (N_45581,N_44109,N_44199);
xnor U45582 (N_45582,N_44389,N_44415);
nor U45583 (N_45583,N_44624,N_44010);
and U45584 (N_45584,N_44403,N_44315);
and U45585 (N_45585,N_44680,N_44537);
or U45586 (N_45586,N_44843,N_44622);
xnor U45587 (N_45587,N_44501,N_44279);
nand U45588 (N_45588,N_44124,N_44539);
xnor U45589 (N_45589,N_44578,N_44809);
nand U45590 (N_45590,N_44850,N_44948);
and U45591 (N_45591,N_44651,N_44704);
nand U45592 (N_45592,N_44776,N_44107);
xor U45593 (N_45593,N_44973,N_44479);
nor U45594 (N_45594,N_44370,N_44363);
nand U45595 (N_45595,N_44623,N_44363);
xnor U45596 (N_45596,N_44048,N_44890);
or U45597 (N_45597,N_44695,N_44156);
nor U45598 (N_45598,N_44064,N_44263);
nand U45599 (N_45599,N_44926,N_44806);
and U45600 (N_45600,N_44105,N_44636);
nor U45601 (N_45601,N_44001,N_44517);
nor U45602 (N_45602,N_44871,N_44624);
nor U45603 (N_45603,N_44560,N_44504);
or U45604 (N_45604,N_44160,N_44251);
and U45605 (N_45605,N_44325,N_44652);
or U45606 (N_45606,N_44203,N_44146);
and U45607 (N_45607,N_44480,N_44464);
and U45608 (N_45608,N_44501,N_44925);
xnor U45609 (N_45609,N_44658,N_44308);
and U45610 (N_45610,N_44975,N_44820);
nand U45611 (N_45611,N_44173,N_44226);
xor U45612 (N_45612,N_44236,N_44862);
and U45613 (N_45613,N_44062,N_44989);
xnor U45614 (N_45614,N_44611,N_44796);
xnor U45615 (N_45615,N_44286,N_44545);
xnor U45616 (N_45616,N_44262,N_44973);
and U45617 (N_45617,N_44901,N_44507);
nor U45618 (N_45618,N_44248,N_44460);
and U45619 (N_45619,N_44864,N_44136);
or U45620 (N_45620,N_44877,N_44846);
xnor U45621 (N_45621,N_44717,N_44659);
nand U45622 (N_45622,N_44218,N_44426);
nand U45623 (N_45623,N_44207,N_44514);
or U45624 (N_45624,N_44785,N_44216);
nor U45625 (N_45625,N_44321,N_44105);
nand U45626 (N_45626,N_44173,N_44360);
or U45627 (N_45627,N_44696,N_44450);
xor U45628 (N_45628,N_44802,N_44749);
xnor U45629 (N_45629,N_44637,N_44445);
and U45630 (N_45630,N_44257,N_44812);
nand U45631 (N_45631,N_44937,N_44007);
and U45632 (N_45632,N_44219,N_44207);
nand U45633 (N_45633,N_44058,N_44089);
nand U45634 (N_45634,N_44511,N_44605);
xor U45635 (N_45635,N_44661,N_44801);
xor U45636 (N_45636,N_44039,N_44567);
xor U45637 (N_45637,N_44474,N_44585);
xor U45638 (N_45638,N_44573,N_44899);
nor U45639 (N_45639,N_44655,N_44240);
nor U45640 (N_45640,N_44967,N_44515);
and U45641 (N_45641,N_44932,N_44923);
nand U45642 (N_45642,N_44729,N_44225);
and U45643 (N_45643,N_44283,N_44973);
and U45644 (N_45644,N_44480,N_44507);
nor U45645 (N_45645,N_44717,N_44484);
or U45646 (N_45646,N_44294,N_44654);
and U45647 (N_45647,N_44463,N_44118);
nand U45648 (N_45648,N_44204,N_44407);
nand U45649 (N_45649,N_44295,N_44540);
xor U45650 (N_45650,N_44550,N_44652);
nand U45651 (N_45651,N_44186,N_44793);
nor U45652 (N_45652,N_44458,N_44658);
or U45653 (N_45653,N_44610,N_44616);
and U45654 (N_45654,N_44325,N_44906);
nor U45655 (N_45655,N_44967,N_44127);
xnor U45656 (N_45656,N_44253,N_44450);
and U45657 (N_45657,N_44298,N_44490);
or U45658 (N_45658,N_44333,N_44473);
and U45659 (N_45659,N_44454,N_44209);
and U45660 (N_45660,N_44194,N_44847);
nor U45661 (N_45661,N_44765,N_44555);
or U45662 (N_45662,N_44081,N_44697);
and U45663 (N_45663,N_44784,N_44527);
or U45664 (N_45664,N_44654,N_44391);
nand U45665 (N_45665,N_44196,N_44269);
and U45666 (N_45666,N_44845,N_44163);
nor U45667 (N_45667,N_44257,N_44132);
or U45668 (N_45668,N_44139,N_44772);
and U45669 (N_45669,N_44678,N_44927);
and U45670 (N_45670,N_44502,N_44748);
nand U45671 (N_45671,N_44417,N_44418);
nand U45672 (N_45672,N_44774,N_44468);
nand U45673 (N_45673,N_44392,N_44610);
nand U45674 (N_45674,N_44924,N_44738);
and U45675 (N_45675,N_44603,N_44200);
nor U45676 (N_45676,N_44493,N_44224);
xnor U45677 (N_45677,N_44580,N_44437);
nand U45678 (N_45678,N_44254,N_44150);
xor U45679 (N_45679,N_44063,N_44962);
or U45680 (N_45680,N_44917,N_44455);
nor U45681 (N_45681,N_44639,N_44959);
nor U45682 (N_45682,N_44122,N_44499);
xor U45683 (N_45683,N_44453,N_44411);
or U45684 (N_45684,N_44049,N_44436);
nand U45685 (N_45685,N_44015,N_44514);
xor U45686 (N_45686,N_44129,N_44149);
nand U45687 (N_45687,N_44372,N_44599);
and U45688 (N_45688,N_44619,N_44753);
or U45689 (N_45689,N_44015,N_44289);
or U45690 (N_45690,N_44693,N_44887);
xor U45691 (N_45691,N_44397,N_44889);
or U45692 (N_45692,N_44644,N_44310);
or U45693 (N_45693,N_44653,N_44323);
and U45694 (N_45694,N_44830,N_44766);
nand U45695 (N_45695,N_44546,N_44078);
nand U45696 (N_45696,N_44464,N_44564);
and U45697 (N_45697,N_44565,N_44468);
xor U45698 (N_45698,N_44449,N_44591);
xnor U45699 (N_45699,N_44803,N_44752);
or U45700 (N_45700,N_44684,N_44780);
or U45701 (N_45701,N_44853,N_44192);
xor U45702 (N_45702,N_44745,N_44845);
or U45703 (N_45703,N_44568,N_44426);
nor U45704 (N_45704,N_44150,N_44983);
and U45705 (N_45705,N_44956,N_44853);
and U45706 (N_45706,N_44694,N_44602);
or U45707 (N_45707,N_44828,N_44437);
or U45708 (N_45708,N_44294,N_44505);
or U45709 (N_45709,N_44957,N_44472);
or U45710 (N_45710,N_44992,N_44434);
or U45711 (N_45711,N_44316,N_44907);
nor U45712 (N_45712,N_44869,N_44893);
xnor U45713 (N_45713,N_44502,N_44613);
nand U45714 (N_45714,N_44748,N_44681);
or U45715 (N_45715,N_44750,N_44763);
nor U45716 (N_45716,N_44604,N_44844);
or U45717 (N_45717,N_44459,N_44953);
and U45718 (N_45718,N_44583,N_44259);
or U45719 (N_45719,N_44998,N_44333);
nand U45720 (N_45720,N_44736,N_44728);
xor U45721 (N_45721,N_44511,N_44221);
xnor U45722 (N_45722,N_44353,N_44123);
or U45723 (N_45723,N_44109,N_44693);
or U45724 (N_45724,N_44735,N_44949);
nand U45725 (N_45725,N_44128,N_44455);
and U45726 (N_45726,N_44680,N_44216);
xor U45727 (N_45727,N_44814,N_44092);
nand U45728 (N_45728,N_44130,N_44905);
nor U45729 (N_45729,N_44136,N_44304);
nand U45730 (N_45730,N_44460,N_44601);
and U45731 (N_45731,N_44710,N_44582);
nand U45732 (N_45732,N_44827,N_44726);
and U45733 (N_45733,N_44503,N_44763);
and U45734 (N_45734,N_44901,N_44101);
nor U45735 (N_45735,N_44280,N_44043);
or U45736 (N_45736,N_44189,N_44042);
and U45737 (N_45737,N_44315,N_44881);
xor U45738 (N_45738,N_44044,N_44959);
xnor U45739 (N_45739,N_44018,N_44730);
nor U45740 (N_45740,N_44653,N_44814);
and U45741 (N_45741,N_44697,N_44620);
nand U45742 (N_45742,N_44025,N_44291);
or U45743 (N_45743,N_44984,N_44824);
nor U45744 (N_45744,N_44849,N_44745);
xor U45745 (N_45745,N_44149,N_44401);
nor U45746 (N_45746,N_44424,N_44766);
or U45747 (N_45747,N_44735,N_44682);
nand U45748 (N_45748,N_44910,N_44228);
nand U45749 (N_45749,N_44816,N_44636);
nand U45750 (N_45750,N_44630,N_44468);
xor U45751 (N_45751,N_44073,N_44003);
nand U45752 (N_45752,N_44024,N_44003);
or U45753 (N_45753,N_44615,N_44270);
xnor U45754 (N_45754,N_44312,N_44015);
or U45755 (N_45755,N_44609,N_44718);
nor U45756 (N_45756,N_44803,N_44554);
nor U45757 (N_45757,N_44401,N_44719);
or U45758 (N_45758,N_44597,N_44358);
nor U45759 (N_45759,N_44981,N_44095);
xor U45760 (N_45760,N_44705,N_44475);
nor U45761 (N_45761,N_44013,N_44082);
nor U45762 (N_45762,N_44739,N_44867);
and U45763 (N_45763,N_44383,N_44684);
or U45764 (N_45764,N_44434,N_44785);
nand U45765 (N_45765,N_44482,N_44032);
xnor U45766 (N_45766,N_44266,N_44276);
and U45767 (N_45767,N_44878,N_44456);
xor U45768 (N_45768,N_44757,N_44463);
nand U45769 (N_45769,N_44346,N_44571);
and U45770 (N_45770,N_44116,N_44581);
nand U45771 (N_45771,N_44008,N_44373);
and U45772 (N_45772,N_44802,N_44204);
or U45773 (N_45773,N_44107,N_44625);
xnor U45774 (N_45774,N_44732,N_44891);
or U45775 (N_45775,N_44656,N_44382);
or U45776 (N_45776,N_44829,N_44491);
nand U45777 (N_45777,N_44974,N_44298);
xnor U45778 (N_45778,N_44143,N_44344);
xnor U45779 (N_45779,N_44978,N_44667);
nand U45780 (N_45780,N_44048,N_44775);
xor U45781 (N_45781,N_44226,N_44018);
nand U45782 (N_45782,N_44921,N_44369);
and U45783 (N_45783,N_44492,N_44246);
and U45784 (N_45784,N_44716,N_44952);
nand U45785 (N_45785,N_44330,N_44169);
and U45786 (N_45786,N_44612,N_44157);
nand U45787 (N_45787,N_44592,N_44497);
nand U45788 (N_45788,N_44739,N_44057);
nor U45789 (N_45789,N_44135,N_44170);
nor U45790 (N_45790,N_44221,N_44994);
or U45791 (N_45791,N_44811,N_44852);
or U45792 (N_45792,N_44100,N_44453);
nand U45793 (N_45793,N_44925,N_44538);
xnor U45794 (N_45794,N_44889,N_44122);
xnor U45795 (N_45795,N_44714,N_44274);
xor U45796 (N_45796,N_44413,N_44586);
or U45797 (N_45797,N_44454,N_44709);
and U45798 (N_45798,N_44845,N_44204);
and U45799 (N_45799,N_44801,N_44227);
nand U45800 (N_45800,N_44197,N_44045);
and U45801 (N_45801,N_44950,N_44219);
nor U45802 (N_45802,N_44814,N_44740);
nand U45803 (N_45803,N_44431,N_44005);
or U45804 (N_45804,N_44648,N_44345);
xnor U45805 (N_45805,N_44201,N_44397);
nand U45806 (N_45806,N_44547,N_44816);
nand U45807 (N_45807,N_44198,N_44421);
and U45808 (N_45808,N_44378,N_44445);
xor U45809 (N_45809,N_44839,N_44467);
nor U45810 (N_45810,N_44916,N_44336);
and U45811 (N_45811,N_44587,N_44556);
nor U45812 (N_45812,N_44112,N_44146);
and U45813 (N_45813,N_44722,N_44281);
and U45814 (N_45814,N_44915,N_44741);
or U45815 (N_45815,N_44737,N_44436);
or U45816 (N_45816,N_44083,N_44569);
and U45817 (N_45817,N_44789,N_44638);
and U45818 (N_45818,N_44475,N_44302);
nand U45819 (N_45819,N_44096,N_44016);
nand U45820 (N_45820,N_44310,N_44196);
xor U45821 (N_45821,N_44934,N_44360);
and U45822 (N_45822,N_44575,N_44721);
nand U45823 (N_45823,N_44561,N_44265);
xor U45824 (N_45824,N_44792,N_44853);
xnor U45825 (N_45825,N_44295,N_44832);
nand U45826 (N_45826,N_44296,N_44660);
nor U45827 (N_45827,N_44185,N_44361);
or U45828 (N_45828,N_44495,N_44941);
or U45829 (N_45829,N_44402,N_44165);
and U45830 (N_45830,N_44381,N_44242);
xnor U45831 (N_45831,N_44910,N_44249);
or U45832 (N_45832,N_44131,N_44242);
nand U45833 (N_45833,N_44330,N_44345);
and U45834 (N_45834,N_44453,N_44105);
or U45835 (N_45835,N_44378,N_44190);
nand U45836 (N_45836,N_44931,N_44846);
and U45837 (N_45837,N_44763,N_44002);
nor U45838 (N_45838,N_44930,N_44751);
nor U45839 (N_45839,N_44902,N_44464);
nand U45840 (N_45840,N_44234,N_44615);
and U45841 (N_45841,N_44404,N_44909);
or U45842 (N_45842,N_44264,N_44530);
and U45843 (N_45843,N_44244,N_44963);
or U45844 (N_45844,N_44909,N_44756);
or U45845 (N_45845,N_44678,N_44505);
and U45846 (N_45846,N_44336,N_44454);
and U45847 (N_45847,N_44344,N_44719);
nand U45848 (N_45848,N_44728,N_44975);
nand U45849 (N_45849,N_44215,N_44991);
xnor U45850 (N_45850,N_44808,N_44945);
or U45851 (N_45851,N_44407,N_44263);
nand U45852 (N_45852,N_44927,N_44282);
nor U45853 (N_45853,N_44502,N_44470);
nand U45854 (N_45854,N_44601,N_44432);
nor U45855 (N_45855,N_44462,N_44048);
or U45856 (N_45856,N_44768,N_44745);
and U45857 (N_45857,N_44798,N_44805);
or U45858 (N_45858,N_44571,N_44306);
nor U45859 (N_45859,N_44028,N_44679);
xnor U45860 (N_45860,N_44627,N_44992);
xnor U45861 (N_45861,N_44637,N_44481);
and U45862 (N_45862,N_44676,N_44312);
nor U45863 (N_45863,N_44261,N_44410);
nand U45864 (N_45864,N_44787,N_44652);
xor U45865 (N_45865,N_44043,N_44939);
nor U45866 (N_45866,N_44609,N_44067);
and U45867 (N_45867,N_44051,N_44815);
xnor U45868 (N_45868,N_44943,N_44377);
nor U45869 (N_45869,N_44307,N_44533);
or U45870 (N_45870,N_44993,N_44672);
xor U45871 (N_45871,N_44773,N_44869);
and U45872 (N_45872,N_44863,N_44067);
or U45873 (N_45873,N_44204,N_44882);
and U45874 (N_45874,N_44239,N_44978);
or U45875 (N_45875,N_44862,N_44706);
nor U45876 (N_45876,N_44197,N_44056);
nor U45877 (N_45877,N_44459,N_44755);
and U45878 (N_45878,N_44770,N_44630);
and U45879 (N_45879,N_44019,N_44446);
nand U45880 (N_45880,N_44744,N_44039);
nor U45881 (N_45881,N_44272,N_44871);
nor U45882 (N_45882,N_44848,N_44102);
nor U45883 (N_45883,N_44271,N_44357);
and U45884 (N_45884,N_44844,N_44548);
nor U45885 (N_45885,N_44503,N_44698);
nand U45886 (N_45886,N_44045,N_44600);
nor U45887 (N_45887,N_44628,N_44240);
or U45888 (N_45888,N_44723,N_44680);
nor U45889 (N_45889,N_44158,N_44536);
xor U45890 (N_45890,N_44053,N_44803);
and U45891 (N_45891,N_44820,N_44805);
or U45892 (N_45892,N_44684,N_44466);
or U45893 (N_45893,N_44721,N_44678);
or U45894 (N_45894,N_44452,N_44645);
xor U45895 (N_45895,N_44705,N_44716);
nor U45896 (N_45896,N_44464,N_44197);
and U45897 (N_45897,N_44737,N_44582);
xor U45898 (N_45898,N_44923,N_44189);
and U45899 (N_45899,N_44134,N_44022);
nand U45900 (N_45900,N_44140,N_44594);
xnor U45901 (N_45901,N_44373,N_44610);
nand U45902 (N_45902,N_44608,N_44556);
and U45903 (N_45903,N_44551,N_44776);
nand U45904 (N_45904,N_44185,N_44956);
nand U45905 (N_45905,N_44628,N_44655);
xor U45906 (N_45906,N_44962,N_44770);
nand U45907 (N_45907,N_44295,N_44592);
nand U45908 (N_45908,N_44999,N_44845);
nand U45909 (N_45909,N_44429,N_44281);
or U45910 (N_45910,N_44264,N_44142);
and U45911 (N_45911,N_44666,N_44720);
or U45912 (N_45912,N_44381,N_44244);
nand U45913 (N_45913,N_44194,N_44783);
and U45914 (N_45914,N_44932,N_44825);
xor U45915 (N_45915,N_44305,N_44981);
and U45916 (N_45916,N_44963,N_44707);
nand U45917 (N_45917,N_44238,N_44609);
nand U45918 (N_45918,N_44431,N_44064);
or U45919 (N_45919,N_44536,N_44770);
xor U45920 (N_45920,N_44490,N_44864);
and U45921 (N_45921,N_44532,N_44245);
xor U45922 (N_45922,N_44071,N_44718);
or U45923 (N_45923,N_44878,N_44338);
nand U45924 (N_45924,N_44337,N_44215);
nand U45925 (N_45925,N_44159,N_44288);
and U45926 (N_45926,N_44971,N_44326);
and U45927 (N_45927,N_44344,N_44018);
nor U45928 (N_45928,N_44325,N_44953);
and U45929 (N_45929,N_44551,N_44130);
and U45930 (N_45930,N_44641,N_44434);
nor U45931 (N_45931,N_44206,N_44301);
nor U45932 (N_45932,N_44820,N_44764);
xor U45933 (N_45933,N_44445,N_44540);
xnor U45934 (N_45934,N_44951,N_44159);
nand U45935 (N_45935,N_44495,N_44523);
xnor U45936 (N_45936,N_44205,N_44297);
and U45937 (N_45937,N_44964,N_44471);
xor U45938 (N_45938,N_44754,N_44940);
and U45939 (N_45939,N_44464,N_44336);
or U45940 (N_45940,N_44534,N_44482);
or U45941 (N_45941,N_44276,N_44883);
nand U45942 (N_45942,N_44627,N_44489);
xor U45943 (N_45943,N_44064,N_44141);
xnor U45944 (N_45944,N_44623,N_44858);
xnor U45945 (N_45945,N_44254,N_44292);
or U45946 (N_45946,N_44274,N_44869);
or U45947 (N_45947,N_44170,N_44089);
nand U45948 (N_45948,N_44129,N_44662);
xnor U45949 (N_45949,N_44865,N_44250);
and U45950 (N_45950,N_44712,N_44349);
nand U45951 (N_45951,N_44018,N_44114);
xor U45952 (N_45952,N_44399,N_44757);
nand U45953 (N_45953,N_44868,N_44317);
and U45954 (N_45954,N_44758,N_44579);
nand U45955 (N_45955,N_44581,N_44159);
nor U45956 (N_45956,N_44097,N_44194);
nand U45957 (N_45957,N_44327,N_44269);
xnor U45958 (N_45958,N_44902,N_44241);
and U45959 (N_45959,N_44451,N_44252);
or U45960 (N_45960,N_44441,N_44202);
nor U45961 (N_45961,N_44537,N_44521);
xor U45962 (N_45962,N_44790,N_44716);
nor U45963 (N_45963,N_44151,N_44179);
nor U45964 (N_45964,N_44457,N_44697);
and U45965 (N_45965,N_44306,N_44665);
nand U45966 (N_45966,N_44731,N_44646);
or U45967 (N_45967,N_44760,N_44369);
and U45968 (N_45968,N_44492,N_44148);
nor U45969 (N_45969,N_44667,N_44130);
or U45970 (N_45970,N_44177,N_44032);
nand U45971 (N_45971,N_44046,N_44032);
xnor U45972 (N_45972,N_44630,N_44038);
xor U45973 (N_45973,N_44664,N_44150);
or U45974 (N_45974,N_44933,N_44873);
xnor U45975 (N_45975,N_44588,N_44482);
nand U45976 (N_45976,N_44029,N_44373);
nand U45977 (N_45977,N_44242,N_44904);
and U45978 (N_45978,N_44275,N_44663);
or U45979 (N_45979,N_44603,N_44135);
nor U45980 (N_45980,N_44938,N_44875);
xnor U45981 (N_45981,N_44922,N_44135);
and U45982 (N_45982,N_44795,N_44856);
nor U45983 (N_45983,N_44874,N_44092);
or U45984 (N_45984,N_44534,N_44073);
xnor U45985 (N_45985,N_44988,N_44155);
xor U45986 (N_45986,N_44784,N_44753);
nand U45987 (N_45987,N_44924,N_44903);
nand U45988 (N_45988,N_44634,N_44694);
or U45989 (N_45989,N_44257,N_44606);
nand U45990 (N_45990,N_44891,N_44759);
xnor U45991 (N_45991,N_44040,N_44767);
or U45992 (N_45992,N_44486,N_44482);
nor U45993 (N_45993,N_44465,N_44650);
nand U45994 (N_45994,N_44757,N_44384);
and U45995 (N_45995,N_44847,N_44518);
nor U45996 (N_45996,N_44327,N_44855);
nand U45997 (N_45997,N_44850,N_44982);
nand U45998 (N_45998,N_44077,N_44467);
nand U45999 (N_45999,N_44777,N_44080);
nand U46000 (N_46000,N_45202,N_45979);
nor U46001 (N_46001,N_45991,N_45024);
and U46002 (N_46002,N_45925,N_45812);
and U46003 (N_46003,N_45646,N_45769);
xor U46004 (N_46004,N_45149,N_45084);
xnor U46005 (N_46005,N_45474,N_45722);
xor U46006 (N_46006,N_45441,N_45236);
nor U46007 (N_46007,N_45672,N_45189);
nand U46008 (N_46008,N_45679,N_45233);
xor U46009 (N_46009,N_45211,N_45071);
and U46010 (N_46010,N_45250,N_45832);
and U46011 (N_46011,N_45718,N_45675);
nor U46012 (N_46012,N_45124,N_45994);
xnor U46013 (N_46013,N_45207,N_45429);
xnor U46014 (N_46014,N_45428,N_45626);
and U46015 (N_46015,N_45455,N_45651);
or U46016 (N_46016,N_45596,N_45047);
nand U46017 (N_46017,N_45512,N_45362);
nor U46018 (N_46018,N_45475,N_45794);
nand U46019 (N_46019,N_45557,N_45744);
xnor U46020 (N_46020,N_45170,N_45327);
nor U46021 (N_46021,N_45692,N_45637);
nand U46022 (N_46022,N_45385,N_45091);
and U46023 (N_46023,N_45530,N_45868);
or U46024 (N_46024,N_45600,N_45366);
nand U46025 (N_46025,N_45280,N_45048);
or U46026 (N_46026,N_45694,N_45714);
xnor U46027 (N_46027,N_45462,N_45238);
nand U46028 (N_46028,N_45519,N_45396);
nand U46029 (N_46029,N_45373,N_45270);
nor U46030 (N_46030,N_45161,N_45576);
and U46031 (N_46031,N_45405,N_45623);
nor U46032 (N_46032,N_45304,N_45355);
and U46033 (N_46033,N_45768,N_45403);
xnor U46034 (N_46034,N_45864,N_45847);
nor U46035 (N_46035,N_45368,N_45032);
xnor U46036 (N_46036,N_45816,N_45595);
and U46037 (N_46037,N_45805,N_45904);
nor U46038 (N_46038,N_45206,N_45974);
nor U46039 (N_46039,N_45761,N_45518);
nor U46040 (N_46040,N_45825,N_45175);
or U46041 (N_46041,N_45871,N_45743);
and U46042 (N_46042,N_45738,N_45758);
or U46043 (N_46043,N_45398,N_45218);
or U46044 (N_46044,N_45110,N_45147);
or U46045 (N_46045,N_45693,N_45111);
nand U46046 (N_46046,N_45819,N_45547);
nor U46047 (N_46047,N_45815,N_45948);
xor U46048 (N_46048,N_45453,N_45186);
nand U46049 (N_46049,N_45751,N_45906);
or U46050 (N_46050,N_45578,N_45029);
nor U46051 (N_46051,N_45187,N_45099);
nand U46052 (N_46052,N_45687,N_45004);
nor U46053 (N_46053,N_45964,N_45940);
nand U46054 (N_46054,N_45877,N_45570);
or U46055 (N_46055,N_45162,N_45848);
nand U46056 (N_46056,N_45089,N_45747);
nor U46057 (N_46057,N_45840,N_45425);
and U46058 (N_46058,N_45311,N_45834);
xnor U46059 (N_46059,N_45706,N_45021);
xor U46060 (N_46060,N_45484,N_45204);
xnor U46061 (N_46061,N_45305,N_45662);
nor U46062 (N_46062,N_45533,N_45619);
xnor U46063 (N_46063,N_45326,N_45934);
nor U46064 (N_46064,N_45826,N_45513);
nor U46065 (N_46065,N_45856,N_45126);
and U46066 (N_46066,N_45944,N_45440);
nand U46067 (N_46067,N_45583,N_45865);
nand U46068 (N_46068,N_45114,N_45923);
nor U46069 (N_46069,N_45176,N_45836);
nand U46070 (N_46070,N_45508,N_45612);
and U46071 (N_46071,N_45633,N_45433);
or U46072 (N_46072,N_45509,N_45879);
xor U46073 (N_46073,N_45121,N_45157);
xor U46074 (N_46074,N_45230,N_45336);
nand U46075 (N_46075,N_45063,N_45661);
nand U46076 (N_46076,N_45907,N_45846);
and U46077 (N_46077,N_45567,N_45726);
xor U46078 (N_46078,N_45514,N_45750);
xnor U46079 (N_46079,N_45128,N_45655);
xor U46080 (N_46080,N_45688,N_45521);
xor U46081 (N_46081,N_45828,N_45670);
nand U46082 (N_46082,N_45671,N_45381);
nor U46083 (N_46083,N_45835,N_45265);
or U46084 (N_46084,N_45226,N_45892);
nor U46085 (N_46085,N_45494,N_45011);
nor U46086 (N_46086,N_45749,N_45884);
xnor U46087 (N_46087,N_45967,N_45995);
or U46088 (N_46088,N_45763,N_45924);
xor U46089 (N_46089,N_45616,N_45180);
and U46090 (N_46090,N_45215,N_45677);
nand U46091 (N_46091,N_45792,N_45302);
or U46092 (N_46092,N_45787,N_45849);
or U46093 (N_46093,N_45491,N_45650);
and U46094 (N_46094,N_45267,N_45101);
and U46095 (N_46095,N_45057,N_45622);
nor U46096 (N_46096,N_45080,N_45174);
xor U46097 (N_46097,N_45953,N_45807);
nor U46098 (N_46098,N_45083,N_45213);
nand U46099 (N_46099,N_45698,N_45614);
xor U46100 (N_46100,N_45691,N_45275);
and U46101 (N_46101,N_45166,N_45837);
xnor U46102 (N_46102,N_45258,N_45277);
nor U46103 (N_46103,N_45284,N_45724);
and U46104 (N_46104,N_45361,N_45382);
or U46105 (N_46105,N_45801,N_45308);
and U46106 (N_46106,N_45055,N_45190);
nor U46107 (N_46107,N_45467,N_45565);
nand U46108 (N_46108,N_45332,N_45264);
nand U46109 (N_46109,N_45411,N_45862);
xor U46110 (N_46110,N_45005,N_45402);
xor U46111 (N_46111,N_45960,N_45752);
and U46112 (N_46112,N_45127,N_45893);
and U46113 (N_46113,N_45348,N_45607);
and U46114 (N_46114,N_45729,N_45413);
nand U46115 (N_46115,N_45301,N_45818);
nor U46116 (N_46116,N_45129,N_45478);
nor U46117 (N_46117,N_45704,N_45351);
or U46118 (N_46118,N_45375,N_45016);
and U46119 (N_46119,N_45459,N_45120);
nand U46120 (N_46120,N_45782,N_45232);
xor U46121 (N_46121,N_45342,N_45041);
or U46122 (N_46122,N_45423,N_45850);
nand U46123 (N_46123,N_45303,N_45545);
nor U46124 (N_46124,N_45685,N_45417);
xnor U46125 (N_46125,N_45274,N_45842);
and U46126 (N_46126,N_45745,N_45017);
or U46127 (N_46127,N_45860,N_45088);
or U46128 (N_46128,N_45851,N_45605);
or U46129 (N_46129,N_45469,N_45719);
and U46130 (N_46130,N_45081,N_45510);
and U46131 (N_46131,N_45990,N_45598);
nand U46132 (N_46132,N_45422,N_45087);
or U46133 (N_46133,N_45182,N_45771);
and U46134 (N_46134,N_45689,N_45783);
xnor U46135 (N_46135,N_45784,N_45665);
and U46136 (N_46136,N_45324,N_45439);
nand U46137 (N_46137,N_45732,N_45401);
nor U46138 (N_46138,N_45383,N_45989);
nor U46139 (N_46139,N_45167,N_45221);
and U46140 (N_46140,N_45996,N_45905);
xnor U46141 (N_46141,N_45502,N_45171);
and U46142 (N_46142,N_45955,N_45909);
nand U46143 (N_46143,N_45043,N_45014);
xnor U46144 (N_46144,N_45188,N_45086);
xor U46145 (N_46145,N_45552,N_45294);
xor U46146 (N_46146,N_45575,N_45654);
and U46147 (N_46147,N_45058,N_45969);
xnor U46148 (N_46148,N_45555,N_45278);
nor U46149 (N_46149,N_45943,N_45543);
nor U46150 (N_46150,N_45489,N_45483);
nand U46151 (N_46151,N_45701,N_45037);
xor U46152 (N_46152,N_45810,N_45476);
nand U46153 (N_46153,N_45262,N_45659);
and U46154 (N_46154,N_45119,N_45090);
or U46155 (N_46155,N_45485,N_45020);
xor U46156 (N_46156,N_45318,N_45212);
and U46157 (N_46157,N_45939,N_45416);
nor U46158 (N_46158,N_45910,N_45914);
and U46159 (N_46159,N_45635,N_45870);
xor U46160 (N_46160,N_45052,N_45059);
nor U46161 (N_46161,N_45936,N_45921);
nand U46162 (N_46162,N_45730,N_45105);
xnor U46163 (N_46163,N_45388,N_45617);
and U46164 (N_46164,N_45588,N_45611);
and U46165 (N_46165,N_45045,N_45343);
or U46166 (N_46166,N_45959,N_45370);
or U46167 (N_46167,N_45603,N_45448);
nor U46168 (N_46168,N_45299,N_45886);
nand U46169 (N_46169,N_45984,N_45030);
nand U46170 (N_46170,N_45454,N_45293);
and U46171 (N_46171,N_45092,N_45602);
xor U46172 (N_46172,N_45198,N_45261);
nor U46173 (N_46173,N_45900,N_45885);
xnor U46174 (N_46174,N_45673,N_45137);
and U46175 (N_46175,N_45224,N_45337);
xor U46176 (N_46176,N_45173,N_45197);
xor U46177 (N_46177,N_45621,N_45709);
xor U46178 (N_46178,N_45902,N_45103);
nor U46179 (N_46179,N_45060,N_45447);
nor U46180 (N_46180,N_45184,N_45945);
xnor U46181 (N_46181,N_45515,N_45895);
nand U46182 (N_46182,N_45481,N_45279);
and U46183 (N_46183,N_45916,N_45341);
nand U46184 (N_46184,N_45778,N_45775);
or U46185 (N_46185,N_45053,N_45378);
nand U46186 (N_46186,N_45104,N_45855);
xnor U46187 (N_46187,N_45389,N_45859);
and U46188 (N_46188,N_45929,N_45144);
and U46189 (N_46189,N_45424,N_45806);
and U46190 (N_46190,N_45443,N_45431);
xor U46191 (N_46191,N_45898,N_45386);
and U46192 (N_46192,N_45506,N_45070);
xor U46193 (N_46193,N_45479,N_45678);
and U46194 (N_46194,N_45503,N_45820);
and U46195 (N_46195,N_45406,N_45657);
nand U46196 (N_46196,N_45255,N_45920);
nor U46197 (N_46197,N_45501,N_45574);
nand U46198 (N_46198,N_45629,N_45839);
and U46199 (N_46199,N_45106,N_45899);
nor U46200 (N_46200,N_45804,N_45442);
and U46201 (N_46201,N_45572,N_45156);
nor U46202 (N_46202,N_45019,N_45982);
or U46203 (N_46203,N_45432,N_45210);
nor U46204 (N_46204,N_45497,N_45618);
or U46205 (N_46205,N_45050,N_45580);
nor U46206 (N_46206,N_45329,N_45242);
nand U46207 (N_46207,N_45844,N_45998);
nor U46208 (N_46208,N_45272,N_45018);
nand U46209 (N_46209,N_45788,N_45950);
nor U46210 (N_46210,N_45194,N_45528);
xnor U46211 (N_46211,N_45608,N_45643);
xor U46212 (N_46212,N_45781,N_45504);
xnor U46213 (N_46213,N_45590,N_45196);
and U46214 (N_46214,N_45966,N_45134);
xor U46215 (N_46215,N_45115,N_45534);
nor U46216 (N_46216,N_45040,N_45796);
or U46217 (N_46217,N_45937,N_45094);
xor U46218 (N_46218,N_45553,N_45581);
xor U46219 (N_46219,N_45559,N_45875);
nand U46220 (N_46220,N_45241,N_45823);
nor U46221 (N_46221,N_45981,N_45463);
nand U46222 (N_46222,N_45331,N_45068);
or U46223 (N_46223,N_45705,N_45108);
and U46224 (N_46224,N_45122,N_45814);
nand U46225 (N_46225,N_45721,N_45082);
and U46226 (N_46226,N_45027,N_45800);
xnor U46227 (N_46227,N_45680,N_45015);
or U46228 (N_46228,N_45663,N_45951);
xnor U46229 (N_46229,N_45903,N_45644);
xor U46230 (N_46230,N_45142,N_45314);
xnor U46231 (N_46231,N_45395,N_45098);
nand U46232 (N_46232,N_45445,N_45306);
and U46233 (N_46233,N_45252,N_45551);
and U46234 (N_46234,N_45554,N_45291);
or U46235 (N_46235,N_45069,N_45414);
nand U46236 (N_46236,N_45419,N_45740);
nand U46237 (N_46237,N_45728,N_45532);
xor U46238 (N_46238,N_45947,N_45647);
and U46239 (N_46239,N_45296,N_45843);
xor U46240 (N_46240,N_45667,N_45404);
nand U46241 (N_46241,N_45830,N_45880);
nand U46242 (N_46242,N_45977,N_45770);
nand U46243 (N_46243,N_45283,N_45799);
nand U46244 (N_46244,N_45458,N_45878);
nand U46245 (N_46245,N_45708,N_45697);
and U46246 (N_46246,N_45295,N_45539);
nand U46247 (N_46247,N_45472,N_45333);
nand U46248 (N_46248,N_45359,N_45066);
nor U46249 (N_46249,N_45199,N_45606);
nor U46250 (N_46250,N_45913,N_45217);
or U46251 (N_46251,N_45866,N_45102);
nand U46252 (N_46252,N_45713,N_45911);
nand U46253 (N_46253,N_45307,N_45465);
nand U46254 (N_46254,N_45941,N_45408);
and U46255 (N_46255,N_45400,N_45808);
nor U46256 (N_46256,N_45085,N_45789);
nand U46257 (N_46257,N_45584,N_45377);
xor U46258 (N_46258,N_45288,N_45755);
or U46259 (N_46259,N_45821,N_45488);
xnor U46260 (N_46260,N_45035,N_45961);
and U46261 (N_46261,N_45529,N_45263);
nand U46262 (N_46262,N_45310,N_45972);
and U46263 (N_46263,N_45587,N_45702);
and U46264 (N_46264,N_45322,N_45309);
and U46265 (N_46265,N_45109,N_45418);
nand U46266 (N_46266,N_45216,N_45975);
or U46267 (N_46267,N_45407,N_45957);
or U46268 (N_46268,N_45271,N_45649);
and U46269 (N_46269,N_45882,N_45118);
and U46270 (N_46270,N_45610,N_45894);
nand U46271 (N_46271,N_45364,N_45563);
xnor U46272 (N_46272,N_45349,N_45365);
and U46273 (N_46273,N_45560,N_45315);
or U46274 (N_46274,N_45319,N_45410);
or U46275 (N_46275,N_45942,N_45833);
and U46276 (N_46276,N_45461,N_45931);
and U46277 (N_46277,N_45613,N_45181);
nand U46278 (N_46278,N_45867,N_45430);
and U46279 (N_46279,N_45863,N_45131);
and U46280 (N_46280,N_45736,N_45260);
nand U46281 (N_46281,N_45222,N_45193);
nand U46282 (N_46282,N_45550,N_45220);
and U46283 (N_46283,N_45683,N_45927);
or U46284 (N_46284,N_45876,N_45151);
or U46285 (N_46285,N_45785,N_45225);
or U46286 (N_46286,N_45273,N_45434);
or U46287 (N_46287,N_45857,N_45415);
nor U46288 (N_46288,N_45394,N_45988);
xor U46289 (N_46289,N_45592,N_45130);
xnor U46290 (N_46290,N_45568,N_45227);
xnor U46291 (N_46291,N_45379,N_45460);
or U46292 (N_46292,N_45861,N_45505);
xnor U46293 (N_46293,N_45054,N_45451);
or U46294 (N_46294,N_45841,N_45498);
or U46295 (N_46295,N_45527,N_45593);
xor U46296 (N_46296,N_45676,N_45160);
and U46297 (N_46297,N_45079,N_45737);
or U46298 (N_46298,N_45715,N_45253);
nand U46299 (N_46299,N_45970,N_45591);
nor U46300 (N_46300,N_45372,N_45897);
nor U46301 (N_46301,N_45093,N_45511);
nor U46302 (N_46302,N_45872,N_45074);
nor U46303 (N_46303,N_45874,N_45006);
xor U46304 (N_46304,N_45928,N_45962);
nor U46305 (N_46305,N_45746,N_45470);
nor U46306 (N_46306,N_45772,N_45620);
or U46307 (N_46307,N_45625,N_45051);
nor U46308 (N_46308,N_45954,N_45774);
nor U46309 (N_46309,N_45889,N_45486);
xnor U46310 (N_46310,N_45524,N_45711);
xor U46311 (N_46311,N_45240,N_45245);
nor U46312 (N_46312,N_45464,N_45228);
nor U46313 (N_46313,N_45246,N_45642);
xnor U46314 (N_46314,N_45686,N_45496);
nor U46315 (N_46315,N_45450,N_45541);
nand U46316 (N_46316,N_45760,N_45569);
xnor U46317 (N_46317,N_45354,N_45456);
and U46318 (N_46318,N_45231,N_45627);
xor U46319 (N_46319,N_45542,N_45268);
nand U46320 (N_46320,N_45219,N_45468);
nor U46321 (N_46321,N_45997,N_45901);
or U46322 (N_46322,N_45393,N_45630);
nand U46323 (N_46323,N_45535,N_45869);
or U46324 (N_46324,N_45287,N_45168);
nor U46325 (N_46325,N_45531,N_45421);
and U46326 (N_46326,N_45123,N_45699);
nor U46327 (N_46327,N_45695,N_45358);
nor U46328 (N_46328,N_45033,N_45537);
nor U46329 (N_46329,N_45298,N_45457);
or U46330 (N_46330,N_45203,N_45078);
nor U46331 (N_46331,N_45766,N_45922);
nor U46332 (N_46332,N_45640,N_45992);
nand U46333 (N_46333,N_45095,N_45363);
and U46334 (N_46334,N_45132,N_45172);
nor U46335 (N_46335,N_45731,N_45762);
or U46336 (N_46336,N_45237,N_45148);
xor U46337 (N_46337,N_45276,N_45742);
nand U46338 (N_46338,N_45723,N_45684);
or U46339 (N_46339,N_45412,N_45435);
nand U46340 (N_46340,N_45562,N_45759);
or U46341 (N_46341,N_45891,N_45523);
and U46342 (N_46342,N_45538,N_45185);
and U46343 (N_46343,N_45548,N_45656);
or U46344 (N_46344,N_45205,N_45473);
and U46345 (N_46345,N_45077,N_45003);
xnor U46346 (N_46346,N_45838,N_45290);
or U46347 (N_46347,N_45797,N_45338);
xor U46348 (N_46348,N_45000,N_45399);
xnor U46349 (N_46349,N_45624,N_45282);
nand U46350 (N_46350,N_45436,N_45438);
xor U46351 (N_46351,N_45251,N_45201);
or U46352 (N_46352,N_45397,N_45100);
nand U46353 (N_46353,N_45831,N_45437);
nand U46354 (N_46354,N_45500,N_45579);
or U46355 (N_46355,N_45323,N_45480);
xor U46356 (N_46356,N_45717,N_45887);
nor U46357 (N_46357,N_45209,N_45571);
nor U46358 (N_46358,N_45158,N_45036);
nor U46359 (N_46359,N_45072,N_45169);
and U46360 (N_46360,N_45703,N_45163);
xnor U46361 (N_46361,N_45008,N_45281);
nor U46362 (N_46362,N_45813,N_45561);
xor U46363 (N_46363,N_45636,N_45067);
or U46364 (N_46364,N_45653,N_45143);
nor U46365 (N_46365,N_45780,N_45881);
or U46366 (N_46366,N_45499,N_45604);
xnor U46367 (N_46367,N_45609,N_45344);
nand U46368 (N_46368,N_45628,N_45631);
nand U46369 (N_46369,N_45776,N_45845);
xnor U46370 (N_46370,N_45444,N_45556);
nand U46371 (N_46371,N_45392,N_45139);
and U46372 (N_46372,N_45371,N_45525);
and U46373 (N_46373,N_45980,N_45536);
xnor U46374 (N_46374,N_45756,N_45915);
or U46375 (N_46375,N_45764,N_45065);
xor U46376 (N_46376,N_45179,N_45645);
xnor U46377 (N_46377,N_45133,N_45183);
xor U46378 (N_46378,N_45985,N_45492);
and U46379 (N_46379,N_45888,N_45317);
nor U46380 (N_46380,N_45347,N_45648);
or U46381 (N_46381,N_45125,N_45266);
and U46382 (N_46382,N_45652,N_45064);
nand U46383 (N_46383,N_45854,N_45350);
or U46384 (N_46384,N_45321,N_45822);
or U46385 (N_46385,N_45334,N_45155);
nor U46386 (N_46386,N_45013,N_45076);
and U46387 (N_46387,N_45357,N_45919);
nand U46388 (N_46388,N_45352,N_45978);
xor U46389 (N_46389,N_45589,N_45795);
xnor U46390 (N_46390,N_45958,N_45739);
and U46391 (N_46391,N_45248,N_45012);
xnor U46392 (N_46392,N_45135,N_45420);
xor U46393 (N_46393,N_45075,N_45965);
xor U46394 (N_46394,N_45817,N_45757);
xnor U46395 (N_46395,N_45976,N_45917);
or U46396 (N_46396,N_45779,N_45932);
nand U46397 (N_46397,N_45369,N_45986);
nor U46398 (N_46398,N_45446,N_45669);
xnor U46399 (N_46399,N_45269,N_45152);
and U46400 (N_46400,N_45038,N_45259);
or U46401 (N_46401,N_45374,N_45803);
and U46402 (N_46402,N_45912,N_45025);
xor U46403 (N_46403,N_45116,N_45353);
or U46404 (N_46404,N_45001,N_45177);
nand U46405 (N_46405,N_45140,N_45798);
xor U46406 (N_46406,N_45658,N_45582);
xnor U46407 (N_46407,N_45666,N_45968);
and U46408 (N_46408,N_45802,N_45034);
xnor U46409 (N_46409,N_45773,N_45223);
or U46410 (N_46410,N_45192,N_45987);
or U46411 (N_46411,N_45042,N_45520);
or U46412 (N_46412,N_45244,N_45935);
xnor U46413 (N_46413,N_45938,N_45641);
nand U46414 (N_46414,N_45727,N_45056);
and U46415 (N_46415,N_45164,N_45971);
and U46416 (N_46416,N_45022,N_45700);
nor U46417 (N_46417,N_45002,N_45873);
xor U46418 (N_46418,N_45733,N_45009);
or U46419 (N_46419,N_45330,N_45908);
xnor U46420 (N_46420,N_45380,N_45360);
nor U46421 (N_46421,N_45999,N_45487);
nand U46422 (N_46422,N_45564,N_45634);
or U46423 (N_46423,N_45387,N_45026);
or U46424 (N_46424,N_45522,N_45933);
nand U46425 (N_46425,N_45682,N_45716);
or U46426 (N_46426,N_45852,N_45046);
or U46427 (N_46427,N_45956,N_45858);
nand U46428 (N_46428,N_45926,N_45165);
xor U46429 (N_46429,N_45896,N_45320);
nand U46430 (N_46430,N_45039,N_45449);
nor U46431 (N_46431,N_45707,N_45191);
or U46432 (N_46432,N_45356,N_45249);
nor U46433 (N_46433,N_45599,N_45153);
nand U46434 (N_46434,N_45495,N_45159);
nor U46435 (N_46435,N_45061,N_45138);
xor U46436 (N_46436,N_45023,N_45328);
or U46437 (N_46437,N_45044,N_45586);
nand U46438 (N_46438,N_45660,N_45477);
xor U46439 (N_46439,N_45890,N_45777);
nand U46440 (N_46440,N_45674,N_45062);
nand U46441 (N_46441,N_45594,N_45247);
or U46442 (N_46442,N_45946,N_45493);
nor U46443 (N_46443,N_45300,N_45200);
xnor U46444 (N_46444,N_45690,N_45235);
nor U46445 (N_46445,N_45390,N_45010);
nand U46446 (N_46446,N_45313,N_45316);
or U46447 (N_46447,N_45178,N_45681);
nand U46448 (N_46448,N_45516,N_45112);
and U46449 (N_46449,N_45615,N_45577);
xnor U46450 (N_46450,N_45466,N_45113);
nor U46451 (N_46451,N_45208,N_45791);
nor U46452 (N_46452,N_45664,N_45292);
and U46453 (N_46453,N_45829,N_45632);
nand U46454 (N_46454,N_45285,N_45325);
xnor U46455 (N_46455,N_45289,N_45712);
and U46456 (N_46456,N_45725,N_45234);
and U46457 (N_46457,N_45391,N_45507);
or U46458 (N_46458,N_45918,N_45490);
and U46459 (N_46459,N_45214,N_45286);
nand U46460 (N_46460,N_45786,N_45696);
or U46461 (N_46461,N_45811,N_45597);
nor U46462 (N_46462,N_45339,N_45566);
xnor U46463 (N_46463,N_45949,N_45117);
nand U46464 (N_46464,N_45741,N_45993);
nand U46465 (N_46465,N_45601,N_45734);
or U46466 (N_46466,N_45809,N_45638);
and U46467 (N_46467,N_45471,N_45793);
nand U46468 (N_46468,N_45107,N_45376);
xor U46469 (N_46469,N_45312,N_45028);
nand U46470 (N_46470,N_45853,N_45409);
or U46471 (N_46471,N_45753,N_45335);
xnor U46472 (N_46472,N_45735,N_45540);
or U46473 (N_46473,N_45767,N_45983);
or U46474 (N_46474,N_45136,N_45720);
nand U46475 (N_46475,N_45146,N_45141);
nor U46476 (N_46476,N_45426,N_45145);
xor U46477 (N_46477,N_45585,N_45096);
xnor U46478 (N_46478,N_45573,N_45883);
nor U46479 (N_46479,N_45239,N_45963);
and U46480 (N_46480,N_45340,N_45073);
and U46481 (N_46481,N_45254,N_45930);
nor U46482 (N_46482,N_45346,N_45482);
or U46483 (N_46483,N_45710,N_45154);
xnor U46484 (N_46484,N_45297,N_45049);
nand U46485 (N_46485,N_45748,N_45526);
nand U46486 (N_46486,N_45097,N_45546);
or U46487 (N_46487,N_45229,N_45824);
nand U46488 (N_46488,N_45031,N_45549);
xor U46489 (N_46489,N_45790,N_45150);
nand U46490 (N_46490,N_45367,N_45639);
xnor U46491 (N_46491,N_45195,N_45668);
xor U46492 (N_46492,N_45256,N_45765);
and U46493 (N_46493,N_45827,N_45007);
nand U46494 (N_46494,N_45754,N_45952);
and U46495 (N_46495,N_45452,N_45558);
nor U46496 (N_46496,N_45345,N_45257);
or U46497 (N_46497,N_45243,N_45427);
or U46498 (N_46498,N_45384,N_45973);
nor U46499 (N_46499,N_45517,N_45544);
xnor U46500 (N_46500,N_45003,N_45689);
xnor U46501 (N_46501,N_45609,N_45229);
xnor U46502 (N_46502,N_45438,N_45429);
nor U46503 (N_46503,N_45126,N_45863);
nand U46504 (N_46504,N_45805,N_45118);
xnor U46505 (N_46505,N_45333,N_45347);
xnor U46506 (N_46506,N_45414,N_45004);
and U46507 (N_46507,N_45405,N_45398);
nand U46508 (N_46508,N_45827,N_45680);
or U46509 (N_46509,N_45887,N_45201);
nand U46510 (N_46510,N_45055,N_45957);
nand U46511 (N_46511,N_45028,N_45395);
nor U46512 (N_46512,N_45114,N_45547);
nor U46513 (N_46513,N_45525,N_45103);
and U46514 (N_46514,N_45913,N_45720);
or U46515 (N_46515,N_45079,N_45679);
and U46516 (N_46516,N_45973,N_45468);
or U46517 (N_46517,N_45433,N_45528);
nor U46518 (N_46518,N_45226,N_45117);
nand U46519 (N_46519,N_45017,N_45612);
nand U46520 (N_46520,N_45435,N_45486);
xnor U46521 (N_46521,N_45236,N_45327);
nand U46522 (N_46522,N_45148,N_45451);
nor U46523 (N_46523,N_45935,N_45969);
or U46524 (N_46524,N_45295,N_45493);
nand U46525 (N_46525,N_45975,N_45484);
nor U46526 (N_46526,N_45922,N_45588);
and U46527 (N_46527,N_45377,N_45481);
xor U46528 (N_46528,N_45892,N_45609);
nand U46529 (N_46529,N_45927,N_45917);
and U46530 (N_46530,N_45965,N_45770);
nand U46531 (N_46531,N_45733,N_45419);
nor U46532 (N_46532,N_45759,N_45146);
and U46533 (N_46533,N_45963,N_45528);
nand U46534 (N_46534,N_45379,N_45756);
nor U46535 (N_46535,N_45359,N_45567);
nor U46536 (N_46536,N_45937,N_45947);
and U46537 (N_46537,N_45645,N_45406);
or U46538 (N_46538,N_45741,N_45156);
xor U46539 (N_46539,N_45992,N_45854);
xnor U46540 (N_46540,N_45591,N_45385);
xnor U46541 (N_46541,N_45000,N_45101);
or U46542 (N_46542,N_45838,N_45462);
or U46543 (N_46543,N_45345,N_45412);
nand U46544 (N_46544,N_45465,N_45346);
xnor U46545 (N_46545,N_45400,N_45491);
or U46546 (N_46546,N_45219,N_45239);
nor U46547 (N_46547,N_45674,N_45202);
and U46548 (N_46548,N_45581,N_45864);
or U46549 (N_46549,N_45446,N_45812);
xor U46550 (N_46550,N_45270,N_45227);
xor U46551 (N_46551,N_45924,N_45729);
nand U46552 (N_46552,N_45868,N_45911);
and U46553 (N_46553,N_45561,N_45906);
and U46554 (N_46554,N_45067,N_45048);
nand U46555 (N_46555,N_45314,N_45399);
or U46556 (N_46556,N_45263,N_45839);
nor U46557 (N_46557,N_45413,N_45208);
nor U46558 (N_46558,N_45193,N_45810);
xor U46559 (N_46559,N_45513,N_45849);
nor U46560 (N_46560,N_45265,N_45171);
or U46561 (N_46561,N_45508,N_45374);
xor U46562 (N_46562,N_45155,N_45847);
nor U46563 (N_46563,N_45072,N_45997);
and U46564 (N_46564,N_45711,N_45733);
and U46565 (N_46565,N_45613,N_45893);
or U46566 (N_46566,N_45524,N_45205);
nor U46567 (N_46567,N_45354,N_45994);
nor U46568 (N_46568,N_45815,N_45536);
nand U46569 (N_46569,N_45203,N_45129);
nand U46570 (N_46570,N_45985,N_45520);
nand U46571 (N_46571,N_45093,N_45251);
or U46572 (N_46572,N_45734,N_45967);
nand U46573 (N_46573,N_45241,N_45001);
and U46574 (N_46574,N_45112,N_45591);
nand U46575 (N_46575,N_45057,N_45121);
or U46576 (N_46576,N_45746,N_45135);
nor U46577 (N_46577,N_45000,N_45551);
nand U46578 (N_46578,N_45522,N_45422);
xor U46579 (N_46579,N_45749,N_45385);
xnor U46580 (N_46580,N_45554,N_45903);
xor U46581 (N_46581,N_45883,N_45624);
or U46582 (N_46582,N_45510,N_45644);
or U46583 (N_46583,N_45930,N_45589);
nand U46584 (N_46584,N_45459,N_45571);
nand U46585 (N_46585,N_45182,N_45892);
and U46586 (N_46586,N_45358,N_45356);
xor U46587 (N_46587,N_45732,N_45425);
nor U46588 (N_46588,N_45178,N_45907);
and U46589 (N_46589,N_45196,N_45044);
and U46590 (N_46590,N_45589,N_45375);
xnor U46591 (N_46591,N_45647,N_45756);
or U46592 (N_46592,N_45704,N_45160);
xor U46593 (N_46593,N_45564,N_45918);
nand U46594 (N_46594,N_45751,N_45244);
or U46595 (N_46595,N_45541,N_45979);
nor U46596 (N_46596,N_45928,N_45959);
and U46597 (N_46597,N_45501,N_45414);
and U46598 (N_46598,N_45263,N_45646);
nor U46599 (N_46599,N_45272,N_45246);
nor U46600 (N_46600,N_45907,N_45640);
and U46601 (N_46601,N_45053,N_45264);
nand U46602 (N_46602,N_45794,N_45267);
xor U46603 (N_46603,N_45359,N_45617);
or U46604 (N_46604,N_45899,N_45132);
or U46605 (N_46605,N_45625,N_45647);
xnor U46606 (N_46606,N_45478,N_45724);
and U46607 (N_46607,N_45959,N_45431);
nor U46608 (N_46608,N_45340,N_45782);
xnor U46609 (N_46609,N_45984,N_45489);
nor U46610 (N_46610,N_45583,N_45097);
nand U46611 (N_46611,N_45382,N_45926);
and U46612 (N_46612,N_45636,N_45997);
xor U46613 (N_46613,N_45072,N_45704);
nand U46614 (N_46614,N_45586,N_45832);
or U46615 (N_46615,N_45962,N_45025);
nand U46616 (N_46616,N_45880,N_45916);
nor U46617 (N_46617,N_45936,N_45089);
nand U46618 (N_46618,N_45360,N_45373);
xor U46619 (N_46619,N_45719,N_45308);
and U46620 (N_46620,N_45452,N_45586);
xor U46621 (N_46621,N_45541,N_45861);
and U46622 (N_46622,N_45105,N_45929);
or U46623 (N_46623,N_45193,N_45611);
xor U46624 (N_46624,N_45578,N_45883);
xnor U46625 (N_46625,N_45880,N_45240);
and U46626 (N_46626,N_45206,N_45991);
xnor U46627 (N_46627,N_45826,N_45302);
and U46628 (N_46628,N_45785,N_45236);
nor U46629 (N_46629,N_45543,N_45211);
or U46630 (N_46630,N_45768,N_45794);
nand U46631 (N_46631,N_45493,N_45153);
nor U46632 (N_46632,N_45766,N_45089);
and U46633 (N_46633,N_45064,N_45406);
xnor U46634 (N_46634,N_45494,N_45653);
nand U46635 (N_46635,N_45283,N_45120);
or U46636 (N_46636,N_45101,N_45111);
nor U46637 (N_46637,N_45978,N_45807);
or U46638 (N_46638,N_45442,N_45426);
and U46639 (N_46639,N_45600,N_45930);
and U46640 (N_46640,N_45161,N_45333);
xnor U46641 (N_46641,N_45320,N_45700);
nand U46642 (N_46642,N_45506,N_45411);
and U46643 (N_46643,N_45925,N_45172);
and U46644 (N_46644,N_45463,N_45362);
or U46645 (N_46645,N_45663,N_45738);
or U46646 (N_46646,N_45358,N_45008);
xnor U46647 (N_46647,N_45221,N_45096);
and U46648 (N_46648,N_45112,N_45729);
nand U46649 (N_46649,N_45746,N_45725);
nand U46650 (N_46650,N_45984,N_45994);
nor U46651 (N_46651,N_45492,N_45388);
or U46652 (N_46652,N_45519,N_45891);
xor U46653 (N_46653,N_45319,N_45961);
or U46654 (N_46654,N_45983,N_45737);
or U46655 (N_46655,N_45199,N_45131);
nor U46656 (N_46656,N_45910,N_45421);
xor U46657 (N_46657,N_45738,N_45129);
or U46658 (N_46658,N_45229,N_45372);
nand U46659 (N_46659,N_45854,N_45683);
or U46660 (N_46660,N_45491,N_45606);
or U46661 (N_46661,N_45585,N_45903);
nand U46662 (N_46662,N_45375,N_45034);
nand U46663 (N_46663,N_45701,N_45541);
or U46664 (N_46664,N_45038,N_45778);
nor U46665 (N_46665,N_45378,N_45777);
xnor U46666 (N_46666,N_45219,N_45442);
nand U46667 (N_46667,N_45137,N_45987);
nor U46668 (N_46668,N_45652,N_45091);
xor U46669 (N_46669,N_45681,N_45461);
and U46670 (N_46670,N_45822,N_45756);
xnor U46671 (N_46671,N_45719,N_45501);
xor U46672 (N_46672,N_45897,N_45514);
and U46673 (N_46673,N_45921,N_45095);
xnor U46674 (N_46674,N_45333,N_45815);
nand U46675 (N_46675,N_45876,N_45271);
nor U46676 (N_46676,N_45954,N_45676);
and U46677 (N_46677,N_45706,N_45806);
nand U46678 (N_46678,N_45260,N_45022);
and U46679 (N_46679,N_45543,N_45554);
xor U46680 (N_46680,N_45718,N_45884);
nor U46681 (N_46681,N_45756,N_45411);
nand U46682 (N_46682,N_45111,N_45298);
or U46683 (N_46683,N_45869,N_45463);
nand U46684 (N_46684,N_45160,N_45183);
nand U46685 (N_46685,N_45499,N_45306);
nor U46686 (N_46686,N_45768,N_45185);
or U46687 (N_46687,N_45090,N_45805);
nor U46688 (N_46688,N_45912,N_45633);
or U46689 (N_46689,N_45549,N_45386);
or U46690 (N_46690,N_45294,N_45069);
or U46691 (N_46691,N_45986,N_45943);
and U46692 (N_46692,N_45614,N_45396);
or U46693 (N_46693,N_45564,N_45761);
nand U46694 (N_46694,N_45856,N_45805);
xnor U46695 (N_46695,N_45249,N_45740);
nand U46696 (N_46696,N_45002,N_45656);
nor U46697 (N_46697,N_45759,N_45394);
nor U46698 (N_46698,N_45715,N_45033);
nor U46699 (N_46699,N_45203,N_45887);
nor U46700 (N_46700,N_45554,N_45273);
nand U46701 (N_46701,N_45379,N_45120);
nor U46702 (N_46702,N_45570,N_45678);
or U46703 (N_46703,N_45130,N_45457);
and U46704 (N_46704,N_45241,N_45531);
or U46705 (N_46705,N_45319,N_45706);
nand U46706 (N_46706,N_45985,N_45015);
xnor U46707 (N_46707,N_45483,N_45427);
and U46708 (N_46708,N_45507,N_45152);
or U46709 (N_46709,N_45876,N_45708);
xor U46710 (N_46710,N_45096,N_45432);
or U46711 (N_46711,N_45301,N_45504);
and U46712 (N_46712,N_45286,N_45041);
nand U46713 (N_46713,N_45721,N_45466);
nand U46714 (N_46714,N_45368,N_45995);
nand U46715 (N_46715,N_45003,N_45329);
nand U46716 (N_46716,N_45709,N_45151);
and U46717 (N_46717,N_45071,N_45330);
and U46718 (N_46718,N_45834,N_45526);
and U46719 (N_46719,N_45058,N_45803);
and U46720 (N_46720,N_45287,N_45927);
and U46721 (N_46721,N_45671,N_45087);
xor U46722 (N_46722,N_45398,N_45763);
and U46723 (N_46723,N_45322,N_45299);
and U46724 (N_46724,N_45767,N_45903);
or U46725 (N_46725,N_45307,N_45346);
xnor U46726 (N_46726,N_45671,N_45174);
or U46727 (N_46727,N_45139,N_45029);
xor U46728 (N_46728,N_45130,N_45710);
xnor U46729 (N_46729,N_45440,N_45320);
nor U46730 (N_46730,N_45821,N_45981);
nor U46731 (N_46731,N_45427,N_45771);
or U46732 (N_46732,N_45044,N_45906);
or U46733 (N_46733,N_45428,N_45066);
nand U46734 (N_46734,N_45320,N_45130);
nand U46735 (N_46735,N_45444,N_45824);
or U46736 (N_46736,N_45245,N_45252);
nand U46737 (N_46737,N_45674,N_45280);
or U46738 (N_46738,N_45800,N_45352);
nor U46739 (N_46739,N_45365,N_45453);
nand U46740 (N_46740,N_45881,N_45412);
or U46741 (N_46741,N_45447,N_45911);
nor U46742 (N_46742,N_45032,N_45392);
nand U46743 (N_46743,N_45634,N_45397);
nor U46744 (N_46744,N_45756,N_45264);
nor U46745 (N_46745,N_45047,N_45248);
or U46746 (N_46746,N_45502,N_45169);
nor U46747 (N_46747,N_45442,N_45679);
or U46748 (N_46748,N_45143,N_45096);
xor U46749 (N_46749,N_45618,N_45883);
xor U46750 (N_46750,N_45303,N_45083);
and U46751 (N_46751,N_45488,N_45988);
nand U46752 (N_46752,N_45739,N_45112);
nand U46753 (N_46753,N_45044,N_45721);
xnor U46754 (N_46754,N_45359,N_45206);
and U46755 (N_46755,N_45380,N_45645);
or U46756 (N_46756,N_45425,N_45265);
nor U46757 (N_46757,N_45031,N_45481);
nand U46758 (N_46758,N_45209,N_45115);
nand U46759 (N_46759,N_45099,N_45158);
and U46760 (N_46760,N_45594,N_45941);
and U46761 (N_46761,N_45248,N_45485);
nand U46762 (N_46762,N_45902,N_45490);
and U46763 (N_46763,N_45428,N_45406);
nor U46764 (N_46764,N_45585,N_45252);
nor U46765 (N_46765,N_45891,N_45870);
and U46766 (N_46766,N_45042,N_45480);
or U46767 (N_46767,N_45904,N_45960);
nand U46768 (N_46768,N_45875,N_45599);
or U46769 (N_46769,N_45452,N_45109);
nor U46770 (N_46770,N_45528,N_45873);
and U46771 (N_46771,N_45757,N_45224);
nand U46772 (N_46772,N_45980,N_45848);
and U46773 (N_46773,N_45862,N_45009);
nand U46774 (N_46774,N_45189,N_45719);
nor U46775 (N_46775,N_45101,N_45957);
xor U46776 (N_46776,N_45803,N_45599);
or U46777 (N_46777,N_45841,N_45561);
nor U46778 (N_46778,N_45037,N_45664);
nand U46779 (N_46779,N_45534,N_45218);
nor U46780 (N_46780,N_45960,N_45793);
or U46781 (N_46781,N_45747,N_45333);
nor U46782 (N_46782,N_45335,N_45901);
xor U46783 (N_46783,N_45987,N_45044);
nor U46784 (N_46784,N_45219,N_45183);
or U46785 (N_46785,N_45713,N_45562);
nor U46786 (N_46786,N_45609,N_45182);
nor U46787 (N_46787,N_45634,N_45234);
nand U46788 (N_46788,N_45875,N_45260);
and U46789 (N_46789,N_45962,N_45813);
xnor U46790 (N_46790,N_45062,N_45620);
xnor U46791 (N_46791,N_45363,N_45312);
and U46792 (N_46792,N_45424,N_45708);
xor U46793 (N_46793,N_45443,N_45594);
xor U46794 (N_46794,N_45728,N_45758);
and U46795 (N_46795,N_45214,N_45836);
nand U46796 (N_46796,N_45504,N_45955);
and U46797 (N_46797,N_45659,N_45275);
xor U46798 (N_46798,N_45006,N_45788);
and U46799 (N_46799,N_45848,N_45657);
xor U46800 (N_46800,N_45839,N_45843);
nand U46801 (N_46801,N_45937,N_45235);
xor U46802 (N_46802,N_45201,N_45124);
nor U46803 (N_46803,N_45706,N_45619);
xor U46804 (N_46804,N_45444,N_45841);
xor U46805 (N_46805,N_45381,N_45777);
xnor U46806 (N_46806,N_45237,N_45209);
or U46807 (N_46807,N_45024,N_45726);
and U46808 (N_46808,N_45721,N_45055);
nor U46809 (N_46809,N_45468,N_45850);
nor U46810 (N_46810,N_45937,N_45791);
xor U46811 (N_46811,N_45264,N_45069);
nor U46812 (N_46812,N_45090,N_45064);
nand U46813 (N_46813,N_45452,N_45378);
nor U46814 (N_46814,N_45768,N_45124);
nor U46815 (N_46815,N_45756,N_45876);
and U46816 (N_46816,N_45262,N_45864);
or U46817 (N_46817,N_45109,N_45038);
or U46818 (N_46818,N_45095,N_45307);
nand U46819 (N_46819,N_45656,N_45926);
nand U46820 (N_46820,N_45058,N_45822);
and U46821 (N_46821,N_45682,N_45501);
nor U46822 (N_46822,N_45952,N_45792);
and U46823 (N_46823,N_45652,N_45043);
nand U46824 (N_46824,N_45087,N_45190);
nor U46825 (N_46825,N_45984,N_45601);
and U46826 (N_46826,N_45396,N_45027);
and U46827 (N_46827,N_45791,N_45377);
and U46828 (N_46828,N_45929,N_45680);
and U46829 (N_46829,N_45798,N_45575);
nor U46830 (N_46830,N_45043,N_45919);
or U46831 (N_46831,N_45915,N_45318);
nor U46832 (N_46832,N_45235,N_45878);
xnor U46833 (N_46833,N_45993,N_45453);
and U46834 (N_46834,N_45183,N_45904);
and U46835 (N_46835,N_45359,N_45971);
xor U46836 (N_46836,N_45379,N_45812);
xnor U46837 (N_46837,N_45659,N_45546);
nand U46838 (N_46838,N_45181,N_45874);
nor U46839 (N_46839,N_45093,N_45237);
xnor U46840 (N_46840,N_45268,N_45533);
nand U46841 (N_46841,N_45744,N_45698);
or U46842 (N_46842,N_45710,N_45209);
xnor U46843 (N_46843,N_45716,N_45668);
xor U46844 (N_46844,N_45144,N_45122);
or U46845 (N_46845,N_45935,N_45123);
nor U46846 (N_46846,N_45955,N_45255);
nand U46847 (N_46847,N_45016,N_45983);
nand U46848 (N_46848,N_45280,N_45092);
and U46849 (N_46849,N_45198,N_45416);
or U46850 (N_46850,N_45309,N_45370);
xor U46851 (N_46851,N_45710,N_45277);
or U46852 (N_46852,N_45154,N_45985);
or U46853 (N_46853,N_45431,N_45919);
or U46854 (N_46854,N_45941,N_45971);
and U46855 (N_46855,N_45867,N_45032);
and U46856 (N_46856,N_45837,N_45628);
xnor U46857 (N_46857,N_45101,N_45753);
or U46858 (N_46858,N_45940,N_45760);
nor U46859 (N_46859,N_45397,N_45685);
nand U46860 (N_46860,N_45955,N_45805);
xor U46861 (N_46861,N_45067,N_45120);
xor U46862 (N_46862,N_45442,N_45092);
and U46863 (N_46863,N_45680,N_45420);
nand U46864 (N_46864,N_45870,N_45652);
xnor U46865 (N_46865,N_45923,N_45504);
nand U46866 (N_46866,N_45022,N_45148);
xor U46867 (N_46867,N_45769,N_45429);
nor U46868 (N_46868,N_45191,N_45171);
and U46869 (N_46869,N_45502,N_45072);
or U46870 (N_46870,N_45767,N_45848);
nand U46871 (N_46871,N_45112,N_45079);
nor U46872 (N_46872,N_45742,N_45647);
nand U46873 (N_46873,N_45910,N_45726);
nand U46874 (N_46874,N_45008,N_45244);
nand U46875 (N_46875,N_45809,N_45992);
nand U46876 (N_46876,N_45440,N_45638);
and U46877 (N_46877,N_45529,N_45202);
nor U46878 (N_46878,N_45320,N_45911);
nor U46879 (N_46879,N_45900,N_45499);
xor U46880 (N_46880,N_45247,N_45525);
or U46881 (N_46881,N_45264,N_45224);
or U46882 (N_46882,N_45995,N_45577);
or U46883 (N_46883,N_45724,N_45666);
nand U46884 (N_46884,N_45011,N_45598);
nor U46885 (N_46885,N_45651,N_45988);
nor U46886 (N_46886,N_45825,N_45278);
nor U46887 (N_46887,N_45270,N_45430);
or U46888 (N_46888,N_45845,N_45769);
and U46889 (N_46889,N_45352,N_45660);
or U46890 (N_46890,N_45046,N_45016);
nand U46891 (N_46891,N_45216,N_45736);
and U46892 (N_46892,N_45643,N_45789);
or U46893 (N_46893,N_45159,N_45983);
xor U46894 (N_46894,N_45694,N_45233);
and U46895 (N_46895,N_45861,N_45094);
and U46896 (N_46896,N_45307,N_45137);
xnor U46897 (N_46897,N_45699,N_45287);
nor U46898 (N_46898,N_45663,N_45373);
xor U46899 (N_46899,N_45135,N_45712);
xnor U46900 (N_46900,N_45394,N_45899);
and U46901 (N_46901,N_45306,N_45803);
nor U46902 (N_46902,N_45709,N_45723);
or U46903 (N_46903,N_45612,N_45849);
xor U46904 (N_46904,N_45999,N_45954);
and U46905 (N_46905,N_45446,N_45941);
nor U46906 (N_46906,N_45067,N_45728);
xor U46907 (N_46907,N_45324,N_45068);
and U46908 (N_46908,N_45604,N_45326);
and U46909 (N_46909,N_45885,N_45884);
and U46910 (N_46910,N_45689,N_45054);
and U46911 (N_46911,N_45054,N_45442);
nand U46912 (N_46912,N_45086,N_45129);
nor U46913 (N_46913,N_45753,N_45283);
nor U46914 (N_46914,N_45692,N_45192);
nor U46915 (N_46915,N_45076,N_45305);
xnor U46916 (N_46916,N_45640,N_45954);
nor U46917 (N_46917,N_45184,N_45419);
and U46918 (N_46918,N_45764,N_45085);
xnor U46919 (N_46919,N_45669,N_45922);
nand U46920 (N_46920,N_45727,N_45191);
nor U46921 (N_46921,N_45339,N_45375);
xor U46922 (N_46922,N_45730,N_45247);
xor U46923 (N_46923,N_45056,N_45927);
or U46924 (N_46924,N_45092,N_45450);
and U46925 (N_46925,N_45951,N_45461);
nand U46926 (N_46926,N_45767,N_45517);
nand U46927 (N_46927,N_45328,N_45407);
nor U46928 (N_46928,N_45221,N_45639);
nor U46929 (N_46929,N_45479,N_45713);
or U46930 (N_46930,N_45226,N_45028);
nor U46931 (N_46931,N_45714,N_45706);
and U46932 (N_46932,N_45592,N_45188);
nor U46933 (N_46933,N_45559,N_45610);
nor U46934 (N_46934,N_45830,N_45911);
nand U46935 (N_46935,N_45842,N_45474);
nor U46936 (N_46936,N_45302,N_45379);
nor U46937 (N_46937,N_45161,N_45627);
xor U46938 (N_46938,N_45742,N_45118);
xnor U46939 (N_46939,N_45366,N_45443);
xnor U46940 (N_46940,N_45127,N_45129);
and U46941 (N_46941,N_45069,N_45140);
nand U46942 (N_46942,N_45192,N_45330);
or U46943 (N_46943,N_45935,N_45087);
xnor U46944 (N_46944,N_45955,N_45713);
and U46945 (N_46945,N_45201,N_45238);
nor U46946 (N_46946,N_45712,N_45599);
xor U46947 (N_46947,N_45929,N_45413);
or U46948 (N_46948,N_45342,N_45705);
nor U46949 (N_46949,N_45347,N_45025);
nor U46950 (N_46950,N_45580,N_45733);
nand U46951 (N_46951,N_45829,N_45876);
nand U46952 (N_46952,N_45303,N_45420);
nand U46953 (N_46953,N_45211,N_45123);
xor U46954 (N_46954,N_45592,N_45639);
nand U46955 (N_46955,N_45214,N_45507);
and U46956 (N_46956,N_45134,N_45536);
nor U46957 (N_46957,N_45085,N_45634);
or U46958 (N_46958,N_45449,N_45664);
or U46959 (N_46959,N_45286,N_45749);
and U46960 (N_46960,N_45628,N_45055);
nand U46961 (N_46961,N_45737,N_45902);
nor U46962 (N_46962,N_45502,N_45057);
xor U46963 (N_46963,N_45577,N_45912);
and U46964 (N_46964,N_45611,N_45756);
and U46965 (N_46965,N_45482,N_45487);
or U46966 (N_46966,N_45279,N_45630);
nor U46967 (N_46967,N_45584,N_45672);
nor U46968 (N_46968,N_45430,N_45946);
and U46969 (N_46969,N_45458,N_45325);
or U46970 (N_46970,N_45190,N_45759);
nand U46971 (N_46971,N_45147,N_45137);
nand U46972 (N_46972,N_45201,N_45510);
and U46973 (N_46973,N_45655,N_45661);
xnor U46974 (N_46974,N_45190,N_45287);
nand U46975 (N_46975,N_45621,N_45970);
xnor U46976 (N_46976,N_45980,N_45285);
and U46977 (N_46977,N_45956,N_45023);
xor U46978 (N_46978,N_45125,N_45762);
nor U46979 (N_46979,N_45925,N_45376);
and U46980 (N_46980,N_45600,N_45303);
and U46981 (N_46981,N_45595,N_45850);
and U46982 (N_46982,N_45029,N_45241);
and U46983 (N_46983,N_45318,N_45073);
nand U46984 (N_46984,N_45024,N_45001);
or U46985 (N_46985,N_45021,N_45119);
nor U46986 (N_46986,N_45043,N_45547);
xnor U46987 (N_46987,N_45263,N_45673);
or U46988 (N_46988,N_45511,N_45288);
or U46989 (N_46989,N_45171,N_45322);
xnor U46990 (N_46990,N_45074,N_45314);
nor U46991 (N_46991,N_45108,N_45829);
or U46992 (N_46992,N_45469,N_45051);
xor U46993 (N_46993,N_45513,N_45679);
nor U46994 (N_46994,N_45674,N_45050);
or U46995 (N_46995,N_45630,N_45830);
xor U46996 (N_46996,N_45746,N_45281);
or U46997 (N_46997,N_45291,N_45863);
nor U46998 (N_46998,N_45486,N_45971);
nor U46999 (N_46999,N_45100,N_45429);
nor U47000 (N_47000,N_46520,N_46475);
or U47001 (N_47001,N_46359,N_46511);
nor U47002 (N_47002,N_46514,N_46190);
xnor U47003 (N_47003,N_46193,N_46168);
nor U47004 (N_47004,N_46509,N_46479);
or U47005 (N_47005,N_46568,N_46563);
or U47006 (N_47006,N_46839,N_46334);
nand U47007 (N_47007,N_46480,N_46277);
nor U47008 (N_47008,N_46517,N_46717);
nor U47009 (N_47009,N_46855,N_46536);
xor U47010 (N_47010,N_46543,N_46130);
xnor U47011 (N_47011,N_46247,N_46437);
or U47012 (N_47012,N_46605,N_46036);
nor U47013 (N_47013,N_46306,N_46452);
nand U47014 (N_47014,N_46987,N_46411);
nor U47015 (N_47015,N_46267,N_46080);
nor U47016 (N_47016,N_46675,N_46676);
nor U47017 (N_47017,N_46912,N_46670);
nor U47018 (N_47018,N_46027,N_46117);
nand U47019 (N_47019,N_46995,N_46524);
or U47020 (N_47020,N_46488,N_46991);
and U47021 (N_47021,N_46200,N_46115);
or U47022 (N_47022,N_46952,N_46460);
xnor U47023 (N_47023,N_46575,N_46063);
or U47024 (N_47024,N_46097,N_46091);
or U47025 (N_47025,N_46899,N_46803);
or U47026 (N_47026,N_46988,N_46639);
nor U47027 (N_47027,N_46137,N_46029);
xor U47028 (N_47028,N_46463,N_46999);
and U47029 (N_47029,N_46667,N_46573);
nor U47030 (N_47030,N_46729,N_46501);
xnor U47031 (N_47031,N_46816,N_46651);
and U47032 (N_47032,N_46406,N_46963);
or U47033 (N_47033,N_46278,N_46449);
nor U47034 (N_47034,N_46333,N_46169);
nor U47035 (N_47035,N_46533,N_46262);
nand U47036 (N_47036,N_46099,N_46045);
nor U47037 (N_47037,N_46645,N_46177);
nor U47038 (N_47038,N_46268,N_46019);
nand U47039 (N_47039,N_46841,N_46212);
or U47040 (N_47040,N_46873,N_46923);
nand U47041 (N_47041,N_46931,N_46018);
xnor U47042 (N_47042,N_46461,N_46287);
xnor U47043 (N_47043,N_46409,N_46219);
and U47044 (N_47044,N_46310,N_46496);
xor U47045 (N_47045,N_46064,N_46060);
or U47046 (N_47046,N_46955,N_46805);
and U47047 (N_47047,N_46625,N_46769);
xnor U47048 (N_47048,N_46489,N_46614);
nand U47049 (N_47049,N_46562,N_46736);
and U47050 (N_47050,N_46565,N_46884);
xor U47051 (N_47051,N_46753,N_46728);
nand U47052 (N_47052,N_46726,N_46210);
xor U47053 (N_47053,N_46126,N_46497);
and U47054 (N_47054,N_46096,N_46281);
xnor U47055 (N_47055,N_46922,N_46879);
xor U47056 (N_47056,N_46778,N_46217);
nor U47057 (N_47057,N_46684,N_46840);
or U47058 (N_47058,N_46085,N_46551);
xnor U47059 (N_47059,N_46171,N_46188);
xor U47060 (N_47060,N_46697,N_46040);
nand U47061 (N_47061,N_46415,N_46288);
nor U47062 (N_47062,N_46900,N_46601);
or U47063 (N_47063,N_46905,N_46291);
nor U47064 (N_47064,N_46612,N_46853);
xor U47065 (N_47065,N_46673,N_46478);
nand U47066 (N_47066,N_46054,N_46748);
or U47067 (N_47067,N_46237,N_46066);
or U47068 (N_47068,N_46035,N_46484);
xnor U47069 (N_47069,N_46048,N_46861);
xor U47070 (N_47070,N_46081,N_46597);
nor U47071 (N_47071,N_46567,N_46631);
nand U47072 (N_47072,N_46093,N_46882);
nor U47073 (N_47073,N_46549,N_46733);
and U47074 (N_47074,N_46227,N_46579);
and U47075 (N_47075,N_46968,N_46438);
nor U47076 (N_47076,N_46499,N_46062);
nor U47077 (N_47077,N_46176,N_46745);
nand U47078 (N_47078,N_46621,N_46155);
and U47079 (N_47079,N_46011,N_46704);
nand U47080 (N_47080,N_46896,N_46980);
xnor U47081 (N_47081,N_46604,N_46957);
and U47082 (N_47082,N_46958,N_46146);
and U47083 (N_47083,N_46355,N_46930);
or U47084 (N_47084,N_46934,N_46807);
xor U47085 (N_47085,N_46413,N_46088);
xnor U47086 (N_47086,N_46820,N_46300);
or U47087 (N_47087,N_46053,N_46788);
nor U47088 (N_47088,N_46809,N_46077);
or U47089 (N_47089,N_46456,N_46588);
nor U47090 (N_47090,N_46919,N_46644);
xor U47091 (N_47091,N_46860,N_46388);
or U47092 (N_47092,N_46215,N_46358);
nand U47093 (N_47093,N_46347,N_46434);
nand U47094 (N_47094,N_46948,N_46867);
nand U47095 (N_47095,N_46638,N_46619);
and U47096 (N_47096,N_46342,N_46608);
xor U47097 (N_47097,N_46422,N_46668);
and U47098 (N_47098,N_46458,N_46251);
nor U47099 (N_47099,N_46942,N_46205);
xor U47100 (N_47100,N_46441,N_46302);
and U47101 (N_47101,N_46823,N_46838);
and U47102 (N_47102,N_46233,N_46801);
nor U47103 (N_47103,N_46365,N_46771);
nand U47104 (N_47104,N_46381,N_46180);
xnor U47105 (N_47105,N_46401,N_46314);
and U47106 (N_47106,N_46510,N_46239);
nor U47107 (N_47107,N_46910,N_46174);
nor U47108 (N_47108,N_46785,N_46556);
nand U47109 (N_47109,N_46775,N_46364);
nor U47110 (N_47110,N_46725,N_46106);
and U47111 (N_47111,N_46353,N_46653);
xnor U47112 (N_47112,N_46741,N_46954);
xor U47113 (N_47113,N_46537,N_46634);
and U47114 (N_47114,N_46050,N_46256);
nor U47115 (N_47115,N_46476,N_46010);
xnor U47116 (N_47116,N_46167,N_46089);
nor U47117 (N_47117,N_46028,N_46553);
nand U47118 (N_47118,N_46084,N_46777);
xnor U47119 (N_47119,N_46315,N_46026);
nor U47120 (N_47120,N_46731,N_46890);
nand U47121 (N_47121,N_46122,N_46003);
or U47122 (N_47122,N_46574,N_46802);
or U47123 (N_47123,N_46373,N_46317);
xnor U47124 (N_47124,N_46844,N_46477);
nand U47125 (N_47125,N_46014,N_46742);
and U47126 (N_47126,N_46285,N_46038);
or U47127 (N_47127,N_46787,N_46301);
xnor U47128 (N_47128,N_46603,N_46711);
and U47129 (N_47129,N_46503,N_46184);
and U47130 (N_47130,N_46012,N_46746);
xnor U47131 (N_47131,N_46786,N_46120);
nand U47132 (N_47132,N_46420,N_46044);
nor U47133 (N_47133,N_46362,N_46135);
nand U47134 (N_47134,N_46490,N_46783);
or U47135 (N_47135,N_46751,N_46542);
or U47136 (N_47136,N_46566,N_46620);
nand U47137 (N_47137,N_46072,N_46580);
nand U47138 (N_47138,N_46328,N_46981);
or U47139 (N_47139,N_46990,N_46749);
nor U47140 (N_47140,N_46664,N_46245);
nand U47141 (N_47141,N_46204,N_46055);
or U47142 (N_47142,N_46795,N_46435);
nand U47143 (N_47143,N_46720,N_46747);
and U47144 (N_47144,N_46858,N_46114);
nor U47145 (N_47145,N_46544,N_46624);
xor U47146 (N_47146,N_46383,N_46444);
and U47147 (N_47147,N_46074,N_46175);
xnor U47148 (N_47148,N_46109,N_46796);
nor U47149 (N_47149,N_46033,N_46623);
nor U47150 (N_47150,N_46655,N_46304);
or U47151 (N_47151,N_46221,N_46815);
nand U47152 (N_47152,N_46945,N_46518);
or U47153 (N_47153,N_46056,N_46230);
xor U47154 (N_47154,N_46756,N_46630);
nand U47155 (N_47155,N_46375,N_46973);
nor U47156 (N_47156,N_46862,N_46471);
or U47157 (N_47157,N_46782,N_46405);
xnor U47158 (N_47158,N_46241,N_46762);
nand U47159 (N_47159,N_46031,N_46454);
nor U47160 (N_47160,N_46195,N_46739);
nor U47161 (N_47161,N_46618,N_46352);
nor U47162 (N_47162,N_46760,N_46020);
or U47163 (N_47163,N_46164,N_46951);
and U47164 (N_47164,N_46323,N_46886);
and U47165 (N_47165,N_46545,N_46107);
nor U47166 (N_47166,N_46332,N_46558);
xor U47167 (N_47167,N_46279,N_46552);
nor U47168 (N_47168,N_46687,N_46829);
xnor U47169 (N_47169,N_46773,N_46198);
nor U47170 (N_47170,N_46357,N_46067);
nand U47171 (N_47171,N_46234,N_46207);
nand U47172 (N_47172,N_46439,N_46292);
or U47173 (N_47173,N_46800,N_46997);
nand U47174 (N_47174,N_46859,N_46242);
xnor U47175 (N_47175,N_46863,N_46585);
or U47176 (N_47176,N_46978,N_46949);
or U47177 (N_47177,N_46395,N_46560);
nor U47178 (N_47178,N_46340,N_46335);
or U47179 (N_47179,N_46700,N_46271);
xnor U47180 (N_47180,N_46950,N_46123);
nor U47181 (N_47181,N_46308,N_46436);
or U47182 (N_47182,N_46901,N_46136);
nand U47183 (N_47183,N_46424,N_46034);
xnor U47184 (N_47184,N_46400,N_46290);
nor U47185 (N_47185,N_46376,N_46979);
or U47186 (N_47186,N_46992,N_46133);
and U47187 (N_47187,N_46070,N_46540);
xor U47188 (N_47188,N_46804,N_46532);
nand U47189 (N_47189,N_46069,N_46068);
and U47190 (N_47190,N_46962,N_46160);
xor U47191 (N_47191,N_46734,N_46904);
nor U47192 (N_47192,N_46329,N_46776);
nor U47193 (N_47193,N_46892,N_46913);
and U47194 (N_47194,N_46309,N_46508);
nand U47195 (N_47195,N_46345,N_46535);
xor U47196 (N_47196,N_46691,N_46094);
xnor U47197 (N_47197,N_46289,N_46525);
or U47198 (N_47198,N_46921,N_46286);
nand U47199 (N_47199,N_46681,N_46004);
and U47200 (N_47200,N_46512,N_46276);
xor U47201 (N_47201,N_46534,N_46513);
nand U47202 (N_47202,N_46702,N_46421);
and U47203 (N_47203,N_46893,N_46946);
and U47204 (N_47204,N_46455,N_46515);
and U47205 (N_47205,N_46961,N_46548);
nor U47206 (N_47206,N_46390,N_46875);
nor U47207 (N_47207,N_46522,N_46235);
and U47208 (N_47208,N_46170,N_46825);
and U47209 (N_47209,N_46743,N_46214);
nor U47210 (N_47210,N_46633,N_46025);
and U47211 (N_47211,N_46482,N_46417);
nand U47212 (N_47212,N_46147,N_46819);
xnor U47213 (N_47213,N_46822,N_46626);
nand U47214 (N_47214,N_46008,N_46039);
nor U47215 (N_47215,N_46927,N_46849);
or U47216 (N_47216,N_46337,N_46685);
or U47217 (N_47217,N_46557,N_46131);
or U47218 (N_47218,N_46985,N_46346);
nand U47219 (N_47219,N_46216,N_46648);
nand U47220 (N_47220,N_46000,N_46202);
nor U47221 (N_47221,N_46453,N_46758);
and U47222 (N_47222,N_46102,N_46022);
xor U47223 (N_47223,N_46470,N_46403);
or U47224 (N_47224,N_46850,N_46678);
xor U47225 (N_47225,N_46159,N_46158);
nand U47226 (N_47226,N_46236,N_46928);
xnor U47227 (N_47227,N_46370,N_46794);
nand U47228 (N_47228,N_46977,N_46495);
nand U47229 (N_47229,N_46095,N_46582);
xnor U47230 (N_47230,N_46492,N_46935);
xor U47231 (N_47231,N_46843,N_46464);
and U47232 (N_47232,N_46732,N_46764);
nand U47233 (N_47233,N_46766,N_46847);
nor U47234 (N_47234,N_46688,N_46172);
and U47235 (N_47235,N_46058,N_46888);
xor U47236 (N_47236,N_46663,N_46113);
or U47237 (N_47237,N_46087,N_46701);
and U47238 (N_47238,N_46763,N_46692);
xor U47239 (N_47239,N_46600,N_46294);
nand U47240 (N_47240,N_46752,N_46516);
or U47241 (N_47241,N_46658,N_46918);
nand U47242 (N_47242,N_46791,N_46360);
nor U47243 (N_47243,N_46336,N_46679);
nor U47244 (N_47244,N_46361,N_46299);
nand U47245 (N_47245,N_46396,N_46821);
nand U47246 (N_47246,N_46683,N_46939);
nor U47247 (N_47247,N_46715,N_46468);
or U47248 (N_47248,N_46419,N_46295);
nand U47249 (N_47249,N_46866,N_46249);
nand U47250 (N_47250,N_46827,N_46589);
nor U47251 (N_47251,N_46322,N_46937);
xnor U47252 (N_47252,N_46628,N_46143);
nor U47253 (N_47253,N_46369,N_46491);
nand U47254 (N_47254,N_46153,N_46940);
nand U47255 (N_47255,N_46924,N_46851);
or U47256 (N_47256,N_46206,N_46293);
or U47257 (N_47257,N_46706,N_46920);
nor U47258 (N_47258,N_46964,N_46248);
nand U47259 (N_47259,N_46616,N_46569);
xnor U47260 (N_47260,N_46989,N_46982);
nor U47261 (N_47261,N_46727,N_46041);
or U47262 (N_47262,N_46561,N_46057);
and U47263 (N_47263,N_46909,N_46713);
nand U47264 (N_47264,N_46870,N_46666);
nor U47265 (N_47265,N_46680,N_46211);
or U47266 (N_47266,N_46046,N_46016);
nor U47267 (N_47267,N_46166,N_46194);
nand U47268 (N_47268,N_46349,N_46694);
xor U47269 (N_47269,N_46654,N_46152);
or U47270 (N_47270,N_46142,N_46721);
xnor U47271 (N_47271,N_46469,N_46779);
nor U47272 (N_47272,N_46015,N_46538);
and U47273 (N_47273,N_46149,N_46103);
nand U47274 (N_47274,N_46897,N_46223);
nor U47275 (N_47275,N_46090,N_46933);
nand U47276 (N_47276,N_46554,N_46986);
and U47277 (N_47277,N_46772,N_46643);
or U47278 (N_47278,N_46865,N_46264);
nand U47279 (N_47279,N_46790,N_46002);
and U47280 (N_47280,N_46864,N_46440);
or U47281 (N_47281,N_46891,N_46459);
xnor U47282 (N_47282,N_46494,N_46425);
and U47283 (N_47283,N_46877,N_46723);
nand U47284 (N_47284,N_46972,N_46876);
or U47285 (N_47285,N_46208,N_46363);
nor U47286 (N_47286,N_46521,N_46856);
xor U47287 (N_47287,N_46757,N_46124);
or U47288 (N_47288,N_46075,N_46627);
or U47289 (N_47289,N_46367,N_46254);
or U47290 (N_47290,N_46784,N_46344);
nand U47291 (N_47291,N_46707,N_46156);
nand U47292 (N_47292,N_46504,N_46086);
nand U47293 (N_47293,N_46652,N_46507);
xor U47294 (N_47294,N_46065,N_46854);
nor U47295 (N_47295,N_46483,N_46399);
nor U47296 (N_47296,N_46646,N_46082);
and U47297 (N_47297,N_46813,N_46793);
nor U47298 (N_47298,N_46564,N_46593);
or U47299 (N_47299,N_46837,N_46780);
nand U47300 (N_47300,N_46970,N_46996);
and U47301 (N_47301,N_46209,N_46023);
nor U47302 (N_47302,N_46445,N_46830);
nand U47303 (N_47303,N_46686,N_46914);
nor U47304 (N_47304,N_46519,N_46178);
nor U47305 (N_47305,N_46049,N_46586);
nor U47306 (N_47306,N_46885,N_46283);
nor U47307 (N_47307,N_46530,N_46881);
xnor U47308 (N_47308,N_46781,N_46872);
nand U47309 (N_47309,N_46179,N_46547);
or U47310 (N_47310,N_46374,N_46125);
xnor U47311 (N_47311,N_46611,N_46581);
or U47312 (N_47312,N_46319,N_46774);
nor U47313 (N_47313,N_46737,N_46959);
xor U47314 (N_47314,N_46121,N_46157);
xor U47315 (N_47315,N_46541,N_46220);
and U47316 (N_47316,N_46690,N_46141);
xnor U47317 (N_47317,N_46506,N_46637);
or U47318 (N_47318,N_46472,N_46100);
and U47319 (N_47319,N_46189,N_46810);
xor U47320 (N_47320,N_46001,N_46154);
nand U47321 (N_47321,N_46682,N_46331);
xor U47322 (N_47322,N_46908,N_46523);
and U47323 (N_47323,N_46321,N_46442);
nand U47324 (N_47324,N_46284,N_46971);
and U47325 (N_47325,N_46430,N_46273);
xnor U47326 (N_47326,N_46831,N_46826);
nand U47327 (N_47327,N_46938,N_46559);
nand U47328 (N_47328,N_46325,N_46378);
and U47329 (N_47329,N_46426,N_46428);
and U47330 (N_47330,N_46186,N_46042);
and U47331 (N_47331,N_46339,N_46635);
and U47332 (N_47332,N_46185,N_46665);
and U47333 (N_47333,N_46274,N_46410);
and U47334 (N_47334,N_46030,N_46591);
nor U47335 (N_47335,N_46974,N_46894);
and U47336 (N_47336,N_46228,N_46191);
nor U47337 (N_47337,N_46138,N_46465);
xor U47338 (N_47338,N_46578,N_46017);
or U47339 (N_47339,N_46151,N_46696);
xor U47340 (N_47340,N_46052,N_46709);
or U47341 (N_47341,N_46617,N_46032);
xor U47342 (N_47342,N_46719,N_46916);
and U47343 (N_47343,N_46832,N_46258);
and U47344 (N_47344,N_46660,N_46671);
xor U47345 (N_47345,N_46051,N_46842);
nor U47346 (N_47346,N_46225,N_46669);
nand U47347 (N_47347,N_46485,N_46338);
nor U47348 (N_47348,N_46622,N_46371);
and U47349 (N_47349,N_46481,N_46526);
nand U47350 (N_47350,N_46078,N_46705);
xnor U47351 (N_47351,N_46350,N_46493);
xnor U47352 (N_47352,N_46457,N_46163);
and U47353 (N_47353,N_46183,N_46698);
nor U47354 (N_47354,N_46555,N_46275);
xor U47355 (N_47355,N_46226,N_46379);
xnor U47356 (N_47356,N_46104,N_46712);
nor U47357 (N_47357,N_46993,N_46738);
xor U47358 (N_47358,N_46699,N_46451);
nor U47359 (N_47359,N_46505,N_46730);
xor U47360 (N_47360,N_46351,N_46944);
nand U47361 (N_47361,N_46474,N_46570);
or U47362 (N_47362,N_46735,N_46929);
nor U47363 (N_47363,N_46119,N_46768);
xor U47364 (N_47364,N_46812,N_46139);
nor U47365 (N_47365,N_46953,N_46083);
or U47366 (N_47366,N_46848,N_46203);
xnor U47367 (N_47367,N_46714,N_46043);
nand U47368 (N_47368,N_46609,N_46677);
nor U47369 (N_47369,N_46594,N_46129);
nor U47370 (N_47370,N_46744,N_46936);
nor U47371 (N_47371,N_46710,N_46969);
nand U47372 (N_47372,N_46009,N_46253);
or U47373 (N_47373,N_46037,N_46846);
xor U47374 (N_47374,N_46059,N_46213);
or U47375 (N_47375,N_46145,N_46318);
and U47376 (N_47376,N_46956,N_46240);
or U47377 (N_47377,N_46531,N_46498);
or U47378 (N_47378,N_46834,N_46161);
and U47379 (N_47379,N_46947,N_46391);
or U47380 (N_47380,N_46407,N_46836);
nor U47381 (N_47381,N_46577,N_46173);
xnor U47382 (N_47382,N_46380,N_46602);
nand U47383 (N_47383,N_46433,N_46528);
nor U47384 (N_47384,N_46368,N_46659);
or U47385 (N_47385,N_46201,N_46414);
xor U47386 (N_47386,N_46320,N_46326);
and U47387 (N_47387,N_46404,N_46382);
or U47388 (N_47388,N_46389,N_46789);
xor U47389 (N_47389,N_46222,N_46307);
nor U47390 (N_47390,N_46366,N_46500);
and U47391 (N_47391,N_46615,N_46148);
or U47392 (N_47392,N_46312,N_46427);
and U47393 (N_47393,N_46606,N_46250);
nor U47394 (N_47394,N_46792,N_46845);
or U47395 (N_47395,N_46806,N_46898);
or U47396 (N_47396,N_46874,N_46903);
nor U47397 (N_47397,N_46192,N_46047);
or U47398 (N_47398,N_46243,N_46402);
nor U47399 (N_47399,N_46599,N_46007);
xor U47400 (N_47400,N_46895,N_46572);
or U47401 (N_47401,N_46252,N_46112);
or U47402 (N_47402,N_46754,N_46828);
and U47403 (N_47403,N_46116,N_46079);
xnor U47404 (N_47404,N_46348,N_46984);
xor U47405 (N_47405,N_46656,N_46224);
or U47406 (N_47406,N_46887,N_46101);
nand U47407 (N_47407,N_46811,N_46718);
xnor U47408 (N_47408,N_46943,N_46313);
xnor U47409 (N_47409,N_46466,N_46649);
or U47410 (N_47410,N_46661,N_46182);
nor U47411 (N_47411,N_46994,N_46906);
and U47412 (N_47412,N_46755,N_46181);
or U47413 (N_47413,N_46632,N_46767);
nand U47414 (N_47414,N_46443,N_46871);
xor U47415 (N_47415,N_46196,N_46006);
nor U47416 (N_47416,N_46911,N_46932);
xor U47417 (N_47417,N_46423,N_46377);
and U47418 (N_47418,N_46467,N_46965);
or U47419 (N_47419,N_46394,N_46610);
or U47420 (N_47420,N_46765,N_46132);
nand U47421 (N_47421,N_46393,N_46397);
xor U47422 (N_47422,N_46587,N_46447);
or U47423 (N_47423,N_46613,N_46590);
xnor U47424 (N_47424,N_46398,N_46092);
nand U47425 (N_47425,N_46689,N_46833);
or U47426 (N_47426,N_46462,N_46797);
and U47427 (N_47427,N_46657,N_46257);
or U47428 (N_47428,N_46356,N_46061);
nand U47429 (N_47429,N_46798,N_46761);
nor U47430 (N_47430,N_46595,N_46502);
xor U47431 (N_47431,N_46473,N_46641);
and U47432 (N_47432,N_46280,N_46303);
nor U47433 (N_47433,N_46372,N_46546);
xor U47434 (N_47434,N_46118,N_46265);
and U47435 (N_47435,N_46330,N_46907);
nand U47436 (N_47436,N_46311,N_46592);
and U47437 (N_47437,N_46387,N_46197);
nand U47438 (N_47438,N_46005,N_46386);
or U47439 (N_47439,N_46868,N_46218);
nor U47440 (N_47440,N_46770,N_46024);
and U47441 (N_47441,N_46297,N_46835);
xnor U47442 (N_47442,N_46571,N_46244);
and U47443 (N_47443,N_46576,N_46127);
or U47444 (N_47444,N_46917,N_46238);
nor U47445 (N_47445,N_46385,N_46607);
xnor U47446 (N_47446,N_46108,N_46298);
nor U47447 (N_47447,N_46246,N_46162);
and U47448 (N_47448,N_46598,N_46740);
or U47449 (N_47449,N_46799,N_46134);
nor U47450 (N_47450,N_46596,N_46071);
and U47451 (N_47451,N_46976,N_46429);
nand U47452 (N_47452,N_46724,N_46967);
and U47453 (N_47453,N_46269,N_46111);
or U47454 (N_47454,N_46925,N_46674);
nor U47455 (N_47455,N_46431,N_46232);
nand U47456 (N_47456,N_46527,N_46529);
nand U47457 (N_47457,N_46384,N_46880);
nor U47458 (N_47458,N_46708,N_46266);
xor U47459 (N_47459,N_46392,N_46642);
nor U47460 (N_47460,N_46324,N_46889);
or U47461 (N_47461,N_46105,N_46305);
nand U47462 (N_47462,N_46231,N_46255);
and U47463 (N_47463,N_46817,N_46341);
or U47464 (N_47464,N_46128,N_46703);
nor U47465 (N_47465,N_46539,N_46941);
or U47466 (N_47466,N_46261,N_46960);
or U47467 (N_47467,N_46750,N_46550);
and U47468 (N_47468,N_46966,N_46327);
or U47469 (N_47469,N_46814,N_46636);
xnor U47470 (N_47470,N_46165,N_46076);
and U47471 (N_47471,N_46448,N_46926);
nand U47472 (N_47472,N_46647,N_46073);
nor U47473 (N_47473,N_46412,N_46693);
and U47474 (N_47474,N_46316,N_46650);
and U47475 (N_47475,N_46354,N_46110);
or U47476 (N_47476,N_46695,N_46487);
and U47477 (N_47477,N_46983,N_46878);
and U47478 (N_47478,N_46282,N_46013);
or U47479 (N_47479,N_46260,N_46263);
nor U47480 (N_47480,N_46824,N_46486);
nand U47481 (N_47481,N_46446,N_46199);
xor U47482 (N_47482,N_46140,N_46021);
nor U47483 (N_47483,N_46716,N_46808);
nor U47484 (N_47484,N_46998,N_46902);
nor U47485 (N_47485,N_46640,N_46584);
and U47486 (N_47486,N_46270,N_46432);
nor U47487 (N_47487,N_46975,N_46144);
and U47488 (N_47488,N_46759,N_46883);
nor U47489 (N_47489,N_46098,N_46852);
xor U47490 (N_47490,N_46187,N_46343);
xnor U47491 (N_47491,N_46869,N_46408);
xor U47492 (N_47492,N_46583,N_46272);
nand U47493 (N_47493,N_46915,N_46672);
nand U47494 (N_47494,N_46150,N_46857);
xnor U47495 (N_47495,N_46450,N_46259);
nand U47496 (N_47496,N_46629,N_46722);
or U47497 (N_47497,N_46416,N_46229);
xor U47498 (N_47498,N_46818,N_46296);
xor U47499 (N_47499,N_46662,N_46418);
nand U47500 (N_47500,N_46536,N_46607);
or U47501 (N_47501,N_46378,N_46763);
nor U47502 (N_47502,N_46391,N_46909);
xnor U47503 (N_47503,N_46430,N_46177);
nand U47504 (N_47504,N_46152,N_46122);
nand U47505 (N_47505,N_46633,N_46851);
nand U47506 (N_47506,N_46887,N_46167);
nand U47507 (N_47507,N_46263,N_46902);
nand U47508 (N_47508,N_46361,N_46382);
and U47509 (N_47509,N_46903,N_46648);
and U47510 (N_47510,N_46916,N_46348);
or U47511 (N_47511,N_46970,N_46104);
and U47512 (N_47512,N_46095,N_46868);
nand U47513 (N_47513,N_46007,N_46482);
and U47514 (N_47514,N_46771,N_46850);
or U47515 (N_47515,N_46931,N_46657);
nand U47516 (N_47516,N_46570,N_46309);
nor U47517 (N_47517,N_46504,N_46030);
and U47518 (N_47518,N_46343,N_46712);
and U47519 (N_47519,N_46171,N_46691);
xor U47520 (N_47520,N_46095,N_46475);
or U47521 (N_47521,N_46335,N_46367);
xnor U47522 (N_47522,N_46359,N_46603);
nor U47523 (N_47523,N_46046,N_46143);
nor U47524 (N_47524,N_46586,N_46274);
nand U47525 (N_47525,N_46110,N_46961);
xor U47526 (N_47526,N_46690,N_46461);
nand U47527 (N_47527,N_46393,N_46360);
nand U47528 (N_47528,N_46760,N_46402);
nand U47529 (N_47529,N_46582,N_46886);
and U47530 (N_47530,N_46943,N_46937);
nand U47531 (N_47531,N_46990,N_46877);
nor U47532 (N_47532,N_46578,N_46548);
nor U47533 (N_47533,N_46067,N_46211);
xnor U47534 (N_47534,N_46029,N_46753);
nor U47535 (N_47535,N_46408,N_46710);
nand U47536 (N_47536,N_46366,N_46729);
nor U47537 (N_47537,N_46597,N_46121);
nand U47538 (N_47538,N_46586,N_46214);
nor U47539 (N_47539,N_46029,N_46525);
or U47540 (N_47540,N_46212,N_46613);
or U47541 (N_47541,N_46242,N_46784);
nor U47542 (N_47542,N_46669,N_46989);
and U47543 (N_47543,N_46414,N_46081);
or U47544 (N_47544,N_46898,N_46467);
xnor U47545 (N_47545,N_46395,N_46633);
nor U47546 (N_47546,N_46784,N_46318);
or U47547 (N_47547,N_46962,N_46404);
and U47548 (N_47548,N_46585,N_46934);
and U47549 (N_47549,N_46919,N_46142);
and U47550 (N_47550,N_46654,N_46103);
xor U47551 (N_47551,N_46390,N_46525);
and U47552 (N_47552,N_46173,N_46931);
and U47553 (N_47553,N_46487,N_46617);
xnor U47554 (N_47554,N_46043,N_46217);
nand U47555 (N_47555,N_46625,N_46916);
or U47556 (N_47556,N_46672,N_46096);
nor U47557 (N_47557,N_46700,N_46518);
or U47558 (N_47558,N_46001,N_46461);
or U47559 (N_47559,N_46588,N_46789);
xor U47560 (N_47560,N_46030,N_46615);
xor U47561 (N_47561,N_46830,N_46481);
or U47562 (N_47562,N_46357,N_46310);
and U47563 (N_47563,N_46831,N_46539);
and U47564 (N_47564,N_46271,N_46348);
or U47565 (N_47565,N_46792,N_46385);
xor U47566 (N_47566,N_46863,N_46503);
xnor U47567 (N_47567,N_46526,N_46440);
and U47568 (N_47568,N_46352,N_46968);
and U47569 (N_47569,N_46316,N_46976);
and U47570 (N_47570,N_46005,N_46935);
nand U47571 (N_47571,N_46890,N_46764);
or U47572 (N_47572,N_46235,N_46599);
xor U47573 (N_47573,N_46044,N_46992);
nor U47574 (N_47574,N_46627,N_46338);
xnor U47575 (N_47575,N_46168,N_46230);
or U47576 (N_47576,N_46098,N_46908);
nand U47577 (N_47577,N_46042,N_46091);
xnor U47578 (N_47578,N_46690,N_46334);
nand U47579 (N_47579,N_46621,N_46098);
xnor U47580 (N_47580,N_46295,N_46186);
or U47581 (N_47581,N_46829,N_46445);
or U47582 (N_47582,N_46488,N_46914);
nor U47583 (N_47583,N_46700,N_46623);
and U47584 (N_47584,N_46568,N_46880);
nand U47585 (N_47585,N_46868,N_46940);
xor U47586 (N_47586,N_46323,N_46652);
and U47587 (N_47587,N_46553,N_46979);
nor U47588 (N_47588,N_46491,N_46179);
xnor U47589 (N_47589,N_46147,N_46201);
nor U47590 (N_47590,N_46772,N_46668);
xor U47591 (N_47591,N_46923,N_46175);
and U47592 (N_47592,N_46952,N_46942);
and U47593 (N_47593,N_46543,N_46136);
xor U47594 (N_47594,N_46384,N_46841);
nand U47595 (N_47595,N_46268,N_46207);
or U47596 (N_47596,N_46538,N_46026);
nor U47597 (N_47597,N_46501,N_46943);
xor U47598 (N_47598,N_46963,N_46667);
nor U47599 (N_47599,N_46445,N_46245);
nor U47600 (N_47600,N_46971,N_46926);
or U47601 (N_47601,N_46759,N_46430);
xor U47602 (N_47602,N_46708,N_46220);
nor U47603 (N_47603,N_46360,N_46747);
or U47604 (N_47604,N_46563,N_46633);
nor U47605 (N_47605,N_46161,N_46805);
nor U47606 (N_47606,N_46235,N_46486);
nor U47607 (N_47607,N_46748,N_46735);
or U47608 (N_47608,N_46007,N_46073);
or U47609 (N_47609,N_46047,N_46388);
xor U47610 (N_47610,N_46600,N_46346);
xnor U47611 (N_47611,N_46603,N_46636);
nor U47612 (N_47612,N_46358,N_46809);
xor U47613 (N_47613,N_46497,N_46858);
xnor U47614 (N_47614,N_46747,N_46147);
xor U47615 (N_47615,N_46895,N_46300);
xnor U47616 (N_47616,N_46718,N_46461);
xor U47617 (N_47617,N_46468,N_46872);
nand U47618 (N_47618,N_46290,N_46327);
or U47619 (N_47619,N_46930,N_46913);
nor U47620 (N_47620,N_46280,N_46017);
xnor U47621 (N_47621,N_46627,N_46341);
nand U47622 (N_47622,N_46446,N_46366);
nand U47623 (N_47623,N_46947,N_46312);
nand U47624 (N_47624,N_46270,N_46448);
or U47625 (N_47625,N_46962,N_46784);
xnor U47626 (N_47626,N_46387,N_46865);
or U47627 (N_47627,N_46719,N_46501);
xor U47628 (N_47628,N_46473,N_46785);
nor U47629 (N_47629,N_46999,N_46036);
and U47630 (N_47630,N_46394,N_46581);
and U47631 (N_47631,N_46954,N_46228);
nand U47632 (N_47632,N_46908,N_46683);
xnor U47633 (N_47633,N_46867,N_46158);
xor U47634 (N_47634,N_46444,N_46882);
xnor U47635 (N_47635,N_46235,N_46751);
and U47636 (N_47636,N_46806,N_46182);
or U47637 (N_47637,N_46984,N_46206);
and U47638 (N_47638,N_46071,N_46646);
xor U47639 (N_47639,N_46444,N_46321);
or U47640 (N_47640,N_46425,N_46041);
nor U47641 (N_47641,N_46637,N_46682);
and U47642 (N_47642,N_46957,N_46906);
and U47643 (N_47643,N_46493,N_46715);
nand U47644 (N_47644,N_46644,N_46623);
and U47645 (N_47645,N_46787,N_46456);
nand U47646 (N_47646,N_46253,N_46332);
nor U47647 (N_47647,N_46241,N_46033);
nand U47648 (N_47648,N_46272,N_46171);
nand U47649 (N_47649,N_46479,N_46318);
xnor U47650 (N_47650,N_46184,N_46066);
nand U47651 (N_47651,N_46046,N_46801);
or U47652 (N_47652,N_46066,N_46189);
xnor U47653 (N_47653,N_46617,N_46661);
xor U47654 (N_47654,N_46029,N_46499);
nor U47655 (N_47655,N_46379,N_46487);
and U47656 (N_47656,N_46327,N_46161);
and U47657 (N_47657,N_46522,N_46463);
and U47658 (N_47658,N_46022,N_46803);
nor U47659 (N_47659,N_46468,N_46233);
and U47660 (N_47660,N_46008,N_46978);
nand U47661 (N_47661,N_46361,N_46506);
nand U47662 (N_47662,N_46980,N_46101);
nor U47663 (N_47663,N_46014,N_46588);
nor U47664 (N_47664,N_46639,N_46641);
nor U47665 (N_47665,N_46878,N_46484);
xnor U47666 (N_47666,N_46588,N_46970);
and U47667 (N_47667,N_46454,N_46758);
and U47668 (N_47668,N_46676,N_46424);
or U47669 (N_47669,N_46101,N_46340);
nand U47670 (N_47670,N_46225,N_46841);
xnor U47671 (N_47671,N_46378,N_46100);
nor U47672 (N_47672,N_46824,N_46869);
or U47673 (N_47673,N_46351,N_46748);
or U47674 (N_47674,N_46159,N_46722);
xor U47675 (N_47675,N_46431,N_46372);
and U47676 (N_47676,N_46997,N_46072);
nor U47677 (N_47677,N_46212,N_46894);
and U47678 (N_47678,N_46023,N_46898);
nor U47679 (N_47679,N_46196,N_46203);
nand U47680 (N_47680,N_46379,N_46097);
and U47681 (N_47681,N_46117,N_46515);
and U47682 (N_47682,N_46991,N_46314);
xor U47683 (N_47683,N_46012,N_46009);
nor U47684 (N_47684,N_46799,N_46368);
nand U47685 (N_47685,N_46334,N_46799);
xor U47686 (N_47686,N_46966,N_46072);
xnor U47687 (N_47687,N_46984,N_46745);
xor U47688 (N_47688,N_46602,N_46295);
or U47689 (N_47689,N_46443,N_46336);
and U47690 (N_47690,N_46540,N_46752);
nand U47691 (N_47691,N_46069,N_46603);
or U47692 (N_47692,N_46954,N_46414);
or U47693 (N_47693,N_46600,N_46979);
nor U47694 (N_47694,N_46239,N_46603);
xnor U47695 (N_47695,N_46263,N_46786);
or U47696 (N_47696,N_46271,N_46275);
nor U47697 (N_47697,N_46231,N_46165);
xnor U47698 (N_47698,N_46229,N_46485);
or U47699 (N_47699,N_46378,N_46039);
or U47700 (N_47700,N_46372,N_46151);
and U47701 (N_47701,N_46027,N_46279);
nand U47702 (N_47702,N_46595,N_46654);
or U47703 (N_47703,N_46961,N_46135);
xnor U47704 (N_47704,N_46266,N_46589);
nand U47705 (N_47705,N_46076,N_46845);
or U47706 (N_47706,N_46184,N_46438);
or U47707 (N_47707,N_46258,N_46967);
xnor U47708 (N_47708,N_46677,N_46633);
xnor U47709 (N_47709,N_46195,N_46411);
xnor U47710 (N_47710,N_46797,N_46461);
nor U47711 (N_47711,N_46598,N_46928);
xor U47712 (N_47712,N_46345,N_46885);
or U47713 (N_47713,N_46223,N_46035);
nand U47714 (N_47714,N_46097,N_46622);
xnor U47715 (N_47715,N_46259,N_46441);
and U47716 (N_47716,N_46913,N_46780);
and U47717 (N_47717,N_46444,N_46900);
nand U47718 (N_47718,N_46943,N_46115);
or U47719 (N_47719,N_46078,N_46381);
nor U47720 (N_47720,N_46587,N_46571);
and U47721 (N_47721,N_46056,N_46677);
xnor U47722 (N_47722,N_46495,N_46613);
xnor U47723 (N_47723,N_46842,N_46589);
and U47724 (N_47724,N_46894,N_46541);
and U47725 (N_47725,N_46302,N_46700);
nor U47726 (N_47726,N_46375,N_46413);
or U47727 (N_47727,N_46339,N_46593);
xnor U47728 (N_47728,N_46525,N_46889);
xor U47729 (N_47729,N_46004,N_46161);
xnor U47730 (N_47730,N_46974,N_46149);
nor U47731 (N_47731,N_46126,N_46377);
or U47732 (N_47732,N_46286,N_46903);
and U47733 (N_47733,N_46733,N_46993);
nand U47734 (N_47734,N_46962,N_46917);
nor U47735 (N_47735,N_46494,N_46513);
xnor U47736 (N_47736,N_46942,N_46252);
nor U47737 (N_47737,N_46198,N_46744);
nand U47738 (N_47738,N_46165,N_46506);
or U47739 (N_47739,N_46447,N_46657);
nor U47740 (N_47740,N_46121,N_46780);
nand U47741 (N_47741,N_46478,N_46613);
or U47742 (N_47742,N_46469,N_46098);
or U47743 (N_47743,N_46391,N_46793);
or U47744 (N_47744,N_46000,N_46352);
xnor U47745 (N_47745,N_46232,N_46531);
nand U47746 (N_47746,N_46786,N_46918);
or U47747 (N_47747,N_46566,N_46389);
nand U47748 (N_47748,N_46376,N_46686);
nor U47749 (N_47749,N_46263,N_46759);
or U47750 (N_47750,N_46576,N_46441);
xnor U47751 (N_47751,N_46699,N_46455);
xnor U47752 (N_47752,N_46742,N_46787);
nor U47753 (N_47753,N_46873,N_46115);
and U47754 (N_47754,N_46540,N_46759);
nor U47755 (N_47755,N_46381,N_46839);
nand U47756 (N_47756,N_46568,N_46399);
and U47757 (N_47757,N_46625,N_46257);
nand U47758 (N_47758,N_46419,N_46169);
nand U47759 (N_47759,N_46568,N_46977);
nand U47760 (N_47760,N_46316,N_46356);
xor U47761 (N_47761,N_46429,N_46458);
or U47762 (N_47762,N_46035,N_46482);
xnor U47763 (N_47763,N_46347,N_46952);
nor U47764 (N_47764,N_46631,N_46274);
nor U47765 (N_47765,N_46294,N_46457);
nand U47766 (N_47766,N_46870,N_46269);
nand U47767 (N_47767,N_46101,N_46069);
nor U47768 (N_47768,N_46536,N_46819);
or U47769 (N_47769,N_46255,N_46156);
xnor U47770 (N_47770,N_46065,N_46732);
and U47771 (N_47771,N_46645,N_46847);
nor U47772 (N_47772,N_46663,N_46027);
nor U47773 (N_47773,N_46671,N_46225);
xor U47774 (N_47774,N_46878,N_46809);
or U47775 (N_47775,N_46743,N_46219);
and U47776 (N_47776,N_46810,N_46556);
and U47777 (N_47777,N_46446,N_46591);
nand U47778 (N_47778,N_46176,N_46188);
and U47779 (N_47779,N_46387,N_46680);
nor U47780 (N_47780,N_46144,N_46434);
xnor U47781 (N_47781,N_46386,N_46451);
or U47782 (N_47782,N_46028,N_46431);
xnor U47783 (N_47783,N_46075,N_46972);
or U47784 (N_47784,N_46140,N_46146);
and U47785 (N_47785,N_46874,N_46891);
or U47786 (N_47786,N_46781,N_46457);
nand U47787 (N_47787,N_46907,N_46908);
nand U47788 (N_47788,N_46395,N_46607);
or U47789 (N_47789,N_46117,N_46917);
nor U47790 (N_47790,N_46084,N_46975);
nand U47791 (N_47791,N_46734,N_46221);
and U47792 (N_47792,N_46029,N_46838);
nand U47793 (N_47793,N_46789,N_46243);
nor U47794 (N_47794,N_46896,N_46233);
nor U47795 (N_47795,N_46257,N_46084);
nand U47796 (N_47796,N_46265,N_46612);
or U47797 (N_47797,N_46422,N_46429);
and U47798 (N_47798,N_46124,N_46701);
or U47799 (N_47799,N_46419,N_46616);
nor U47800 (N_47800,N_46036,N_46311);
and U47801 (N_47801,N_46447,N_46802);
xnor U47802 (N_47802,N_46588,N_46294);
nor U47803 (N_47803,N_46998,N_46159);
nand U47804 (N_47804,N_46217,N_46261);
xor U47805 (N_47805,N_46740,N_46431);
xor U47806 (N_47806,N_46393,N_46057);
nor U47807 (N_47807,N_46852,N_46536);
and U47808 (N_47808,N_46008,N_46081);
and U47809 (N_47809,N_46490,N_46092);
or U47810 (N_47810,N_46769,N_46715);
xnor U47811 (N_47811,N_46425,N_46969);
nand U47812 (N_47812,N_46980,N_46160);
or U47813 (N_47813,N_46167,N_46737);
xnor U47814 (N_47814,N_46161,N_46945);
and U47815 (N_47815,N_46458,N_46023);
or U47816 (N_47816,N_46833,N_46182);
or U47817 (N_47817,N_46222,N_46672);
and U47818 (N_47818,N_46452,N_46986);
nand U47819 (N_47819,N_46888,N_46369);
xnor U47820 (N_47820,N_46109,N_46954);
xnor U47821 (N_47821,N_46605,N_46743);
nand U47822 (N_47822,N_46204,N_46943);
nand U47823 (N_47823,N_46296,N_46506);
or U47824 (N_47824,N_46378,N_46147);
and U47825 (N_47825,N_46289,N_46625);
nand U47826 (N_47826,N_46603,N_46676);
or U47827 (N_47827,N_46594,N_46394);
nor U47828 (N_47828,N_46722,N_46730);
xor U47829 (N_47829,N_46891,N_46399);
or U47830 (N_47830,N_46552,N_46866);
xor U47831 (N_47831,N_46793,N_46609);
and U47832 (N_47832,N_46728,N_46605);
nand U47833 (N_47833,N_46975,N_46414);
nand U47834 (N_47834,N_46426,N_46063);
nor U47835 (N_47835,N_46641,N_46709);
nand U47836 (N_47836,N_46328,N_46206);
or U47837 (N_47837,N_46135,N_46558);
and U47838 (N_47838,N_46299,N_46056);
or U47839 (N_47839,N_46420,N_46748);
nand U47840 (N_47840,N_46473,N_46008);
xnor U47841 (N_47841,N_46182,N_46475);
and U47842 (N_47842,N_46537,N_46327);
nand U47843 (N_47843,N_46592,N_46009);
or U47844 (N_47844,N_46733,N_46316);
nand U47845 (N_47845,N_46481,N_46573);
xor U47846 (N_47846,N_46180,N_46839);
nor U47847 (N_47847,N_46547,N_46555);
nor U47848 (N_47848,N_46602,N_46102);
and U47849 (N_47849,N_46978,N_46396);
and U47850 (N_47850,N_46734,N_46078);
nand U47851 (N_47851,N_46389,N_46031);
or U47852 (N_47852,N_46990,N_46289);
xnor U47853 (N_47853,N_46699,N_46323);
and U47854 (N_47854,N_46067,N_46317);
xor U47855 (N_47855,N_46210,N_46148);
or U47856 (N_47856,N_46338,N_46377);
xor U47857 (N_47857,N_46326,N_46142);
xnor U47858 (N_47858,N_46613,N_46248);
nand U47859 (N_47859,N_46180,N_46060);
nand U47860 (N_47860,N_46347,N_46055);
or U47861 (N_47861,N_46284,N_46794);
nor U47862 (N_47862,N_46214,N_46847);
nand U47863 (N_47863,N_46130,N_46180);
xor U47864 (N_47864,N_46359,N_46915);
or U47865 (N_47865,N_46481,N_46879);
xnor U47866 (N_47866,N_46674,N_46809);
or U47867 (N_47867,N_46638,N_46700);
nand U47868 (N_47868,N_46822,N_46662);
nand U47869 (N_47869,N_46890,N_46772);
or U47870 (N_47870,N_46262,N_46405);
nor U47871 (N_47871,N_46529,N_46847);
and U47872 (N_47872,N_46640,N_46663);
xnor U47873 (N_47873,N_46635,N_46040);
nor U47874 (N_47874,N_46973,N_46197);
xnor U47875 (N_47875,N_46539,N_46417);
nor U47876 (N_47876,N_46300,N_46909);
and U47877 (N_47877,N_46633,N_46491);
nand U47878 (N_47878,N_46404,N_46715);
xor U47879 (N_47879,N_46921,N_46653);
nand U47880 (N_47880,N_46993,N_46030);
nand U47881 (N_47881,N_46715,N_46842);
and U47882 (N_47882,N_46675,N_46819);
and U47883 (N_47883,N_46570,N_46278);
or U47884 (N_47884,N_46176,N_46292);
or U47885 (N_47885,N_46380,N_46785);
and U47886 (N_47886,N_46187,N_46416);
or U47887 (N_47887,N_46614,N_46080);
xnor U47888 (N_47888,N_46960,N_46958);
and U47889 (N_47889,N_46013,N_46628);
xnor U47890 (N_47890,N_46814,N_46409);
nor U47891 (N_47891,N_46118,N_46334);
nor U47892 (N_47892,N_46373,N_46654);
nand U47893 (N_47893,N_46841,N_46181);
nand U47894 (N_47894,N_46375,N_46583);
or U47895 (N_47895,N_46639,N_46003);
nand U47896 (N_47896,N_46562,N_46787);
nor U47897 (N_47897,N_46300,N_46484);
nand U47898 (N_47898,N_46139,N_46495);
or U47899 (N_47899,N_46152,N_46307);
nor U47900 (N_47900,N_46313,N_46222);
nand U47901 (N_47901,N_46979,N_46214);
nand U47902 (N_47902,N_46932,N_46241);
nand U47903 (N_47903,N_46773,N_46135);
xor U47904 (N_47904,N_46096,N_46070);
nor U47905 (N_47905,N_46710,N_46483);
or U47906 (N_47906,N_46477,N_46351);
nor U47907 (N_47907,N_46886,N_46572);
nand U47908 (N_47908,N_46123,N_46638);
and U47909 (N_47909,N_46691,N_46331);
nor U47910 (N_47910,N_46715,N_46627);
or U47911 (N_47911,N_46712,N_46044);
nor U47912 (N_47912,N_46557,N_46974);
nor U47913 (N_47913,N_46499,N_46616);
and U47914 (N_47914,N_46698,N_46560);
nor U47915 (N_47915,N_46770,N_46155);
nand U47916 (N_47916,N_46791,N_46497);
nand U47917 (N_47917,N_46077,N_46156);
xor U47918 (N_47918,N_46392,N_46387);
nor U47919 (N_47919,N_46395,N_46179);
xor U47920 (N_47920,N_46834,N_46148);
and U47921 (N_47921,N_46155,N_46321);
nor U47922 (N_47922,N_46714,N_46876);
xor U47923 (N_47923,N_46699,N_46607);
and U47924 (N_47924,N_46003,N_46540);
and U47925 (N_47925,N_46937,N_46941);
and U47926 (N_47926,N_46269,N_46288);
xor U47927 (N_47927,N_46986,N_46174);
nor U47928 (N_47928,N_46075,N_46061);
xnor U47929 (N_47929,N_46628,N_46218);
nand U47930 (N_47930,N_46919,N_46048);
nor U47931 (N_47931,N_46303,N_46681);
or U47932 (N_47932,N_46910,N_46242);
nand U47933 (N_47933,N_46108,N_46099);
and U47934 (N_47934,N_46742,N_46999);
and U47935 (N_47935,N_46123,N_46247);
or U47936 (N_47936,N_46652,N_46641);
and U47937 (N_47937,N_46434,N_46568);
and U47938 (N_47938,N_46872,N_46209);
and U47939 (N_47939,N_46004,N_46789);
xnor U47940 (N_47940,N_46864,N_46574);
nor U47941 (N_47941,N_46796,N_46935);
or U47942 (N_47942,N_46097,N_46574);
and U47943 (N_47943,N_46292,N_46453);
and U47944 (N_47944,N_46744,N_46973);
and U47945 (N_47945,N_46544,N_46106);
xnor U47946 (N_47946,N_46476,N_46280);
and U47947 (N_47947,N_46519,N_46706);
nor U47948 (N_47948,N_46565,N_46114);
and U47949 (N_47949,N_46631,N_46568);
nand U47950 (N_47950,N_46967,N_46974);
nand U47951 (N_47951,N_46705,N_46743);
and U47952 (N_47952,N_46725,N_46859);
xor U47953 (N_47953,N_46407,N_46031);
and U47954 (N_47954,N_46670,N_46889);
nor U47955 (N_47955,N_46816,N_46028);
and U47956 (N_47956,N_46540,N_46570);
nor U47957 (N_47957,N_46884,N_46321);
xnor U47958 (N_47958,N_46179,N_46948);
nand U47959 (N_47959,N_46789,N_46981);
nor U47960 (N_47960,N_46022,N_46347);
nor U47961 (N_47961,N_46366,N_46529);
nand U47962 (N_47962,N_46740,N_46146);
and U47963 (N_47963,N_46235,N_46346);
nand U47964 (N_47964,N_46383,N_46542);
and U47965 (N_47965,N_46470,N_46973);
nand U47966 (N_47966,N_46608,N_46950);
or U47967 (N_47967,N_46252,N_46389);
and U47968 (N_47968,N_46116,N_46334);
xnor U47969 (N_47969,N_46867,N_46188);
nor U47970 (N_47970,N_46535,N_46096);
or U47971 (N_47971,N_46126,N_46634);
nor U47972 (N_47972,N_46849,N_46253);
nor U47973 (N_47973,N_46375,N_46887);
and U47974 (N_47974,N_46330,N_46428);
xnor U47975 (N_47975,N_46259,N_46548);
or U47976 (N_47976,N_46117,N_46796);
xor U47977 (N_47977,N_46136,N_46708);
or U47978 (N_47978,N_46859,N_46036);
nand U47979 (N_47979,N_46153,N_46528);
xor U47980 (N_47980,N_46481,N_46093);
and U47981 (N_47981,N_46124,N_46636);
nand U47982 (N_47982,N_46602,N_46440);
or U47983 (N_47983,N_46079,N_46892);
nor U47984 (N_47984,N_46691,N_46166);
nor U47985 (N_47985,N_46610,N_46766);
or U47986 (N_47986,N_46204,N_46537);
or U47987 (N_47987,N_46263,N_46874);
or U47988 (N_47988,N_46416,N_46029);
and U47989 (N_47989,N_46571,N_46855);
and U47990 (N_47990,N_46253,N_46271);
and U47991 (N_47991,N_46830,N_46897);
xnor U47992 (N_47992,N_46964,N_46597);
nand U47993 (N_47993,N_46050,N_46729);
nand U47994 (N_47994,N_46209,N_46600);
and U47995 (N_47995,N_46235,N_46655);
nand U47996 (N_47996,N_46060,N_46828);
nor U47997 (N_47997,N_46228,N_46846);
nor U47998 (N_47998,N_46687,N_46429);
and U47999 (N_47999,N_46969,N_46372);
nor U48000 (N_48000,N_47916,N_47016);
nand U48001 (N_48001,N_47523,N_47542);
nand U48002 (N_48002,N_47330,N_47602);
and U48003 (N_48003,N_47613,N_47652);
or U48004 (N_48004,N_47486,N_47809);
xor U48005 (N_48005,N_47707,N_47969);
or U48006 (N_48006,N_47792,N_47252);
nand U48007 (N_48007,N_47197,N_47596);
nor U48008 (N_48008,N_47152,N_47996);
or U48009 (N_48009,N_47189,N_47585);
nand U48010 (N_48010,N_47991,N_47510);
xor U48011 (N_48011,N_47636,N_47227);
or U48012 (N_48012,N_47888,N_47056);
or U48013 (N_48013,N_47306,N_47644);
and U48014 (N_48014,N_47610,N_47989);
nor U48015 (N_48015,N_47417,N_47354);
nor U48016 (N_48016,N_47900,N_47304);
and U48017 (N_48017,N_47750,N_47063);
and U48018 (N_48018,N_47032,N_47090);
and U48019 (N_48019,N_47679,N_47935);
nor U48020 (N_48020,N_47084,N_47563);
nor U48021 (N_48021,N_47774,N_47908);
nand U48022 (N_48022,N_47008,N_47919);
and U48023 (N_48023,N_47011,N_47479);
and U48024 (N_48024,N_47561,N_47415);
or U48025 (N_48025,N_47203,N_47641);
xor U48026 (N_48026,N_47493,N_47348);
and U48027 (N_48027,N_47529,N_47349);
or U48028 (N_48028,N_47757,N_47733);
xnor U48029 (N_48029,N_47003,N_47570);
nor U48030 (N_48030,N_47424,N_47307);
and U48031 (N_48031,N_47836,N_47783);
or U48032 (N_48032,N_47186,N_47590);
nand U48033 (N_48033,N_47877,N_47778);
nand U48034 (N_48034,N_47369,N_47393);
nor U48035 (N_48035,N_47817,N_47873);
xor U48036 (N_48036,N_47154,N_47949);
xnor U48037 (N_48037,N_47476,N_47403);
or U48038 (N_48038,N_47893,N_47168);
nand U48039 (N_48039,N_47494,N_47437);
or U48040 (N_48040,N_47970,N_47869);
or U48041 (N_48041,N_47193,N_47030);
xor U48042 (N_48042,N_47866,N_47638);
and U48043 (N_48043,N_47045,N_47279);
nor U48044 (N_48044,N_47519,N_47210);
nor U48045 (N_48045,N_47243,N_47767);
nand U48046 (N_48046,N_47364,N_47997);
or U48047 (N_48047,N_47994,N_47961);
xor U48048 (N_48048,N_47853,N_47628);
nand U48049 (N_48049,N_47847,N_47093);
nand U48050 (N_48050,N_47018,N_47591);
or U48051 (N_48051,N_47400,N_47426);
nor U48052 (N_48052,N_47691,N_47109);
xnor U48053 (N_48053,N_47839,N_47823);
or U48054 (N_48054,N_47301,N_47451);
or U48055 (N_48055,N_47124,N_47050);
nor U48056 (N_48056,N_47717,N_47571);
or U48057 (N_48057,N_47162,N_47594);
nor U48058 (N_48058,N_47785,N_47512);
nand U48059 (N_48059,N_47943,N_47864);
nor U48060 (N_48060,N_47868,N_47879);
or U48061 (N_48061,N_47047,N_47734);
xnor U48062 (N_48062,N_47072,N_47020);
or U48063 (N_48063,N_47959,N_47661);
or U48064 (N_48064,N_47262,N_47577);
nor U48065 (N_48065,N_47067,N_47153);
xnor U48066 (N_48066,N_47752,N_47917);
or U48067 (N_48067,N_47000,N_47681);
or U48068 (N_48068,N_47421,N_47600);
nand U48069 (N_48069,N_47697,N_47356);
nor U48070 (N_48070,N_47956,N_47492);
nand U48071 (N_48071,N_47608,N_47946);
nor U48072 (N_48072,N_47657,N_47992);
nor U48073 (N_48073,N_47040,N_47378);
nor U48074 (N_48074,N_47736,N_47578);
nand U48075 (N_48075,N_47155,N_47553);
nand U48076 (N_48076,N_47719,N_47414);
nor U48077 (N_48077,N_47850,N_47339);
or U48078 (N_48078,N_47901,N_47503);
or U48079 (N_48079,N_47548,N_47222);
or U48080 (N_48080,N_47345,N_47945);
and U48081 (N_48081,N_47801,N_47024);
xor U48082 (N_48082,N_47278,N_47118);
xor U48083 (N_48083,N_47998,N_47704);
nor U48084 (N_48084,N_47208,N_47245);
nor U48085 (N_48085,N_47397,N_47232);
and U48086 (N_48086,N_47485,N_47845);
or U48087 (N_48087,N_47782,N_47293);
or U48088 (N_48088,N_47899,N_47137);
or U48089 (N_48089,N_47722,N_47713);
xnor U48090 (N_48090,N_47487,N_47226);
nand U48091 (N_48091,N_47588,N_47502);
or U48092 (N_48092,N_47972,N_47267);
nor U48093 (N_48093,N_47347,N_47974);
nand U48094 (N_48094,N_47199,N_47151);
nand U48095 (N_48095,N_47004,N_47688);
xor U48096 (N_48096,N_47754,N_47312);
xor U48097 (N_48097,N_47927,N_47676);
nand U48098 (N_48098,N_47743,N_47568);
or U48099 (N_48099,N_47423,N_47791);
nand U48100 (N_48100,N_47834,N_47036);
and U48101 (N_48101,N_47854,N_47457);
or U48102 (N_48102,N_47445,N_47584);
nor U48103 (N_48103,N_47179,N_47240);
nand U48104 (N_48104,N_47844,N_47675);
and U48105 (N_48105,N_47574,N_47695);
nor U48106 (N_48106,N_47357,N_47618);
nand U48107 (N_48107,N_47382,N_47611);
and U48108 (N_48108,N_47058,N_47896);
and U48109 (N_48109,N_47496,N_47670);
nor U48110 (N_48110,N_47526,N_47601);
nor U48111 (N_48111,N_47773,N_47143);
and U48112 (N_48112,N_47883,N_47073);
or U48113 (N_48113,N_47701,N_47291);
and U48114 (N_48114,N_47089,N_47172);
or U48115 (N_48115,N_47119,N_47550);
or U48116 (N_48116,N_47887,N_47790);
nand U48117 (N_48117,N_47039,N_47101);
nor U48118 (N_48118,N_47727,N_47206);
nand U48119 (N_48119,N_47721,N_47474);
xor U48120 (N_48120,N_47022,N_47205);
nand U48121 (N_48121,N_47374,N_47187);
nand U48122 (N_48122,N_47131,N_47082);
or U48123 (N_48123,N_47544,N_47086);
or U48124 (N_48124,N_47122,N_47117);
nand U48125 (N_48125,N_47560,N_47068);
and U48126 (N_48126,N_47800,N_47559);
nor U48127 (N_48127,N_47287,N_47256);
and U48128 (N_48128,N_47764,N_47284);
and U48129 (N_48129,N_47698,N_47121);
or U48130 (N_48130,N_47448,N_47668);
xor U48131 (N_48131,N_47795,N_47753);
or U48132 (N_48132,N_47453,N_47202);
or U48133 (N_48133,N_47066,N_47564);
nor U48134 (N_48134,N_47858,N_47925);
or U48135 (N_48135,N_47371,N_47833);
nor U48136 (N_48136,N_47141,N_47724);
or U48137 (N_48137,N_47219,N_47504);
or U48138 (N_48138,N_47280,N_47111);
and U48139 (N_48139,N_47696,N_47904);
nor U48140 (N_48140,N_47430,N_47516);
nand U48141 (N_48141,N_47412,N_47391);
nor U48142 (N_48142,N_47021,N_47471);
xnor U48143 (N_48143,N_47182,N_47805);
xor U48144 (N_48144,N_47979,N_47178);
and U48145 (N_48145,N_47741,N_47133);
nand U48146 (N_48146,N_47147,N_47110);
or U48147 (N_48147,N_47663,N_47295);
nor U48148 (N_48148,N_47258,N_47837);
nor U48149 (N_48149,N_47087,N_47060);
nor U48150 (N_48150,N_47038,N_47432);
xor U48151 (N_48151,N_47346,N_47710);
xnor U48152 (N_48152,N_47402,N_47007);
or U48153 (N_48153,N_47181,N_47288);
and U48154 (N_48154,N_47253,N_47229);
or U48155 (N_48155,N_47338,N_47742);
xnor U48156 (N_48156,N_47798,N_47794);
nand U48157 (N_48157,N_47239,N_47083);
nand U48158 (N_48158,N_47351,N_47265);
or U48159 (N_48159,N_47880,N_47650);
nor U48160 (N_48160,N_47468,N_47929);
or U48161 (N_48161,N_47127,N_47438);
xnor U48162 (N_48162,N_47419,N_47576);
or U48163 (N_48163,N_47069,N_47300);
and U48164 (N_48164,N_47209,N_47751);
nor U48165 (N_48165,N_47405,N_47687);
nand U48166 (N_48166,N_47454,N_47936);
or U48167 (N_48167,N_47740,N_47671);
nor U48168 (N_48168,N_47748,N_47861);
xor U48169 (N_48169,N_47664,N_47302);
nand U48170 (N_48170,N_47520,N_47034);
and U48171 (N_48171,N_47843,N_47055);
or U48172 (N_48172,N_47455,N_47720);
xor U48173 (N_48173,N_47669,N_47499);
nand U48174 (N_48174,N_47370,N_47480);
nand U48175 (N_48175,N_47612,N_47418);
nor U48176 (N_48176,N_47938,N_47729);
and U48177 (N_48177,N_47857,N_47627);
xnor U48178 (N_48178,N_47379,N_47250);
and U48179 (N_48179,N_47749,N_47971);
or U48180 (N_48180,N_47035,N_47409);
xnor U48181 (N_48181,N_47940,N_47174);
and U48182 (N_48182,N_47260,N_47025);
xor U48183 (N_48183,N_47501,N_47876);
nor U48184 (N_48184,N_47064,N_47048);
and U48185 (N_48185,N_47715,N_47198);
or U48186 (N_48186,N_47614,N_47142);
nor U48187 (N_48187,N_47170,N_47188);
or U48188 (N_48188,N_47184,N_47283);
nor U48189 (N_48189,N_47158,N_47218);
and U48190 (N_48190,N_47659,N_47065);
or U48191 (N_48191,N_47814,N_47120);
xor U48192 (N_48192,N_47275,N_47842);
nor U48193 (N_48193,N_47408,N_47102);
nor U48194 (N_48194,N_47116,N_47760);
xnor U48195 (N_48195,N_47286,N_47460);
or U48196 (N_48196,N_47231,N_47694);
xnor U48197 (N_48197,N_47123,N_47993);
nand U48198 (N_48198,N_47973,N_47770);
or U48199 (N_48199,N_47732,N_47350);
or U48200 (N_48200,N_47268,N_47665);
xor U48201 (N_48201,N_47930,N_47806);
and U48202 (N_48202,N_47881,N_47104);
and U48203 (N_48203,N_47822,N_47728);
nand U48204 (N_48204,N_47075,N_47237);
nand U48205 (N_48205,N_47595,N_47355);
nand U48206 (N_48206,N_47684,N_47091);
xor U48207 (N_48207,N_47508,N_47248);
nor U48208 (N_48208,N_47326,N_47939);
and U48209 (N_48209,N_47603,N_47871);
xnor U48210 (N_48210,N_47952,N_47017);
xnor U48211 (N_48211,N_47289,N_47813);
nand U48212 (N_48212,N_47944,N_47098);
xnor U48213 (N_48213,N_47324,N_47950);
xnor U48214 (N_48214,N_47634,N_47582);
and U48215 (N_48215,N_47921,N_47316);
xnor U48216 (N_48216,N_47495,N_47846);
xnor U48217 (N_48217,N_47658,N_47700);
nor U48218 (N_48218,N_47815,N_47140);
and U48219 (N_48219,N_47551,N_47489);
nand U48220 (N_48220,N_47948,N_47277);
xnor U48221 (N_48221,N_47238,N_47322);
and U48222 (N_48222,N_47201,N_47292);
and U48223 (N_48223,N_47735,N_47463);
and U48224 (N_48224,N_47818,N_47885);
nand U48225 (N_48225,N_47699,N_47444);
nand U48226 (N_48226,N_47129,N_47768);
nor U48227 (N_48227,N_47890,N_47976);
nand U48228 (N_48228,N_47213,N_47458);
or U48229 (N_48229,N_47076,N_47848);
xnor U48230 (N_48230,N_47867,N_47294);
and U48231 (N_48231,N_47865,N_47088);
or U48232 (N_48232,N_47290,N_47894);
or U48233 (N_48233,N_47359,N_47583);
and U48234 (N_48234,N_47318,N_47255);
or U48235 (N_48235,N_47870,N_47281);
nor U48236 (N_48236,N_47144,N_47953);
and U48237 (N_48237,N_47539,N_47235);
or U48238 (N_48238,N_47130,N_47459);
or U48239 (N_48239,N_47183,N_47106);
nor U48240 (N_48240,N_47808,N_47317);
or U48241 (N_48241,N_47505,N_47363);
xor U48242 (N_48242,N_47149,N_47175);
and U48243 (N_48243,N_47525,N_47014);
and U48244 (N_48244,N_47990,N_47545);
and U48245 (N_48245,N_47171,N_47466);
xor U48246 (N_48246,N_47766,N_47367);
and U48247 (N_48247,N_47725,N_47532);
nand U48248 (N_48248,N_47759,N_47984);
xnor U48249 (N_48249,N_47630,N_47625);
xnor U48250 (N_48250,N_47744,N_47620);
and U48251 (N_48251,N_47673,N_47788);
or U48252 (N_48252,N_47257,N_47562);
and U48253 (N_48253,N_47010,N_47856);
xor U48254 (N_48254,N_47597,N_47401);
xnor U48255 (N_48255,N_47233,N_47763);
or U48256 (N_48256,N_47924,N_47810);
and U48257 (N_48257,N_47540,N_47282);
xnor U48258 (N_48258,N_47926,N_47266);
and U48259 (N_48259,N_47598,N_47207);
and U48260 (N_48260,N_47467,N_47737);
and U48261 (N_48261,N_47534,N_47196);
xnor U48262 (N_48262,N_47113,N_47261);
or U48263 (N_48263,N_47321,N_47860);
nor U48264 (N_48264,N_47537,N_47366);
or U48265 (N_48265,N_47947,N_47125);
xnor U48266 (N_48266,N_47506,N_47731);
and U48267 (N_48267,N_47811,N_47033);
or U48268 (N_48268,N_47965,N_47452);
or U48269 (N_48269,N_47392,N_47518);
xnor U48270 (N_48270,N_47019,N_47821);
nand U48271 (N_48271,N_47156,N_47706);
nand U48272 (N_48272,N_47828,N_47365);
nand U48273 (N_48273,N_47450,N_47762);
or U48274 (N_48274,N_47384,N_47928);
nor U48275 (N_48275,N_47541,N_47580);
nand U48276 (N_48276,N_47862,N_47422);
or U48277 (N_48277,N_47703,N_47490);
nor U48278 (N_48278,N_47434,N_47249);
xor U48279 (N_48279,N_47566,N_47986);
nand U48280 (N_48280,N_47380,N_47830);
and U48281 (N_48281,N_47875,N_47522);
xor U48282 (N_48282,N_47332,N_47957);
and U48283 (N_48283,N_47962,N_47647);
or U48284 (N_48284,N_47730,N_47236);
xnor U48285 (N_48285,N_47884,N_47646);
nand U48286 (N_48286,N_47889,N_47922);
xnor U48287 (N_48287,N_47655,N_47586);
or U48288 (N_48288,N_47254,N_47096);
or U48289 (N_48289,N_47159,N_47746);
nor U48290 (N_48290,N_47361,N_47407);
xnor U48291 (N_48291,N_47672,N_47319);
and U48292 (N_48292,N_47745,N_47772);
or U48293 (N_48293,N_47078,N_47711);
and U48294 (N_48294,N_47642,N_47648);
nor U48295 (N_48295,N_47639,N_47824);
nor U48296 (N_48296,N_47395,N_47473);
or U48297 (N_48297,N_47826,N_47211);
nor U48298 (N_48298,N_47941,N_47524);
or U48299 (N_48299,N_47194,N_47427);
or U48300 (N_48300,N_47500,N_47978);
xnor U48301 (N_48301,N_47139,N_47368);
and U48302 (N_48302,N_47934,N_47225);
xnor U48303 (N_48303,N_47832,N_47220);
and U48304 (N_48304,N_47593,N_47755);
or U48305 (N_48305,N_47816,N_47398);
xnor U48306 (N_48306,N_47413,N_47579);
or U48307 (N_48307,N_47388,N_47891);
nand U48308 (N_48308,N_47488,N_47776);
nand U48309 (N_48309,N_47079,N_47263);
nand U48310 (N_48310,N_47975,N_47053);
and U48311 (N_48311,N_47484,N_47299);
nand U48312 (N_48312,N_47352,N_47204);
and U48313 (N_48313,N_47689,N_47533);
nand U48314 (N_48314,N_47342,N_47799);
and U48315 (N_48315,N_47340,N_47624);
or U48316 (N_48316,N_47827,N_47416);
nor U48317 (N_48317,N_47954,N_47999);
or U48318 (N_48318,N_47464,N_47114);
and U48319 (N_48319,N_47910,N_47386);
and U48320 (N_48320,N_47276,N_47581);
nand U48321 (N_48321,N_47645,N_47191);
or U48322 (N_48322,N_47680,N_47511);
and U48323 (N_48323,N_47399,N_47052);
nor U48324 (N_48324,N_47331,N_47726);
nor U48325 (N_48325,N_47977,N_47166);
nand U48326 (N_48326,N_47797,N_47469);
nand U48327 (N_48327,N_47062,N_47164);
xor U48328 (N_48328,N_47146,N_47376);
nor U48329 (N_48329,N_47966,N_47536);
nor U48330 (N_48330,N_47425,N_47223);
nand U48331 (N_48331,N_47920,N_47538);
xnor U48332 (N_48332,N_47041,N_47712);
or U48333 (N_48333,N_47554,N_47043);
xor U48334 (N_48334,N_47851,N_47136);
or U48335 (N_48335,N_47431,N_47428);
or U48336 (N_48336,N_47514,N_47988);
nor U48337 (N_48337,N_47214,N_47377);
or U48338 (N_48338,N_47677,N_47042);
nor U48339 (N_48339,N_47622,N_47441);
xor U48340 (N_48340,N_47360,N_47132);
nor U48341 (N_48341,N_47607,N_47528);
nor U48342 (N_48342,N_47874,N_47796);
or U48343 (N_48343,N_47892,N_47535);
nand U48344 (N_48344,N_47491,N_47200);
and U48345 (N_48345,N_47012,N_47433);
nand U48346 (N_48346,N_47100,N_47002);
nand U48347 (N_48347,N_47557,N_47789);
nor U48348 (N_48348,N_47631,N_47802);
xor U48349 (N_48349,N_47604,N_47309);
xor U48350 (N_48350,N_47353,N_47738);
and U48351 (N_48351,N_47080,N_47558);
or U48352 (N_48352,N_47898,N_47006);
xnor U48353 (N_48353,N_47678,N_47094);
and U48354 (N_48354,N_47835,N_47343);
nand U48355 (N_48355,N_47411,N_47333);
nand U48356 (N_48356,N_47981,N_47656);
nand U48357 (N_48357,N_47660,N_47297);
nand U48358 (N_48358,N_47643,N_47446);
xnor U48359 (N_48359,N_47325,N_47314);
or U48360 (N_48360,N_47148,N_47247);
and U48361 (N_48361,N_47160,N_47362);
xnor U48362 (N_48362,N_47552,N_47264);
xor U48363 (N_48363,N_47115,N_47784);
and U48364 (N_48364,N_47462,N_47420);
xnor U48365 (N_48365,N_47633,N_47305);
nand U48366 (N_48366,N_47057,N_47666);
nor U48367 (N_48367,N_47138,N_47872);
xnor U48368 (N_48368,N_47327,N_47176);
and U48369 (N_48369,N_47215,N_47410);
and U48370 (N_48370,N_47013,N_47481);
nor U48371 (N_48371,N_47244,N_47859);
nand U48372 (N_48372,N_47902,N_47394);
and U48373 (N_48373,N_47819,N_47897);
nor U48374 (N_48374,N_47180,N_47841);
xor U48375 (N_48375,N_47831,N_47313);
or U48376 (N_48376,N_47621,N_47009);
or U48377 (N_48377,N_47112,N_47640);
nand U48378 (N_48378,N_47716,N_47081);
or U48379 (N_48379,N_47723,N_47095);
or U48380 (N_48380,N_47995,N_47190);
xnor U48381 (N_48381,N_47456,N_47224);
nor U48382 (N_48382,N_47906,N_47165);
xor U48383 (N_48383,N_47383,N_47498);
or U48384 (N_48384,N_47787,N_47573);
and U48385 (N_48385,N_47311,N_47054);
xor U48386 (N_48386,N_47549,N_47543);
nor U48387 (N_48387,N_47335,N_47037);
and U48388 (N_48388,N_47027,N_47029);
and U48389 (N_48389,N_47912,N_47482);
nand U48390 (N_48390,N_47105,N_47777);
xor U48391 (N_48391,N_47807,N_47829);
xnor U48392 (N_48392,N_47686,N_47023);
xnor U48393 (N_48393,N_47128,N_47517);
xnor U48394 (N_48394,N_47780,N_47527);
nand U48395 (N_48395,N_47337,N_47513);
or U48396 (N_48396,N_47372,N_47163);
nand U48397 (N_48397,N_47221,N_47216);
xnor U48398 (N_48398,N_47964,N_47389);
and U48399 (N_48399,N_47592,N_47271);
or U48400 (N_48400,N_47982,N_47521);
xnor U48401 (N_48401,N_47274,N_47103);
xnor U48402 (N_48402,N_47708,N_47968);
nor U48403 (N_48403,N_47077,N_47909);
or U48404 (N_48404,N_47623,N_47509);
xnor U48405 (N_48405,N_47135,N_47531);
and U48406 (N_48406,N_47958,N_47031);
or U48407 (N_48407,N_47569,N_47028);
and U48408 (N_48408,N_47985,N_47983);
and U48409 (N_48409,N_47477,N_47882);
xnor U48410 (N_48410,N_47185,N_47878);
nor U48411 (N_48411,N_47606,N_47246);
or U48412 (N_48412,N_47387,N_47914);
or U48413 (N_48413,N_47587,N_47635);
or U48414 (N_48414,N_47615,N_47886);
and U48415 (N_48415,N_47195,N_47515);
nor U48416 (N_48416,N_47242,N_47771);
xnor U48417 (N_48417,N_47739,N_47567);
and U48418 (N_48418,N_47905,N_47918);
nor U48419 (N_48419,N_47461,N_47692);
nand U48420 (N_48420,N_47059,N_47269);
xnor U48421 (N_48421,N_47329,N_47960);
and U48422 (N_48422,N_47609,N_47396);
or U48423 (N_48423,N_47440,N_47097);
xor U48424 (N_48424,N_47475,N_47234);
and U48425 (N_48425,N_47915,N_47980);
or U48426 (N_48426,N_47649,N_47507);
nand U48427 (N_48427,N_47336,N_47617);
or U48428 (N_48428,N_47803,N_47344);
and U48429 (N_48429,N_47272,N_47328);
xor U48430 (N_48430,N_47323,N_47126);
and U48431 (N_48431,N_47942,N_47161);
xor U48432 (N_48432,N_47820,N_47765);
xor U48433 (N_48433,N_47406,N_47756);
nor U48434 (N_48434,N_47632,N_47913);
nand U48435 (N_48435,N_47718,N_47169);
and U48436 (N_48436,N_47044,N_47085);
and U48437 (N_48437,N_47478,N_47967);
and U48438 (N_48438,N_47472,N_47026);
or U48439 (N_48439,N_47070,N_47804);
or U48440 (N_48440,N_47682,N_47605);
xnor U48441 (N_48441,N_47556,N_47439);
xor U48442 (N_48442,N_47217,N_47907);
nand U48443 (N_48443,N_47310,N_47092);
nand U48444 (N_48444,N_47911,N_47761);
nand U48445 (N_48445,N_47390,N_47442);
nand U48446 (N_48446,N_47951,N_47049);
xor U48447 (N_48447,N_47385,N_47546);
and U48448 (N_48448,N_47685,N_47690);
xor U48449 (N_48449,N_47555,N_47449);
nor U48450 (N_48450,N_47812,N_47150);
nor U48451 (N_48451,N_47589,N_47134);
or U48452 (N_48452,N_47145,N_47547);
nand U48453 (N_48453,N_47616,N_47320);
or U48454 (N_48454,N_47099,N_47572);
xor U48455 (N_48455,N_47987,N_47296);
and U48456 (N_48456,N_47933,N_47963);
nor U48457 (N_48457,N_47167,N_47107);
and U48458 (N_48458,N_47470,N_47705);
xnor U48459 (N_48459,N_47825,N_47212);
and U48460 (N_48460,N_47575,N_47775);
nor U48461 (N_48461,N_47447,N_47637);
and U48462 (N_48462,N_47626,N_47937);
nor U48463 (N_48463,N_47483,N_47758);
and U48464 (N_48464,N_47662,N_47334);
or U48465 (N_48465,N_47667,N_47855);
nand U48466 (N_48466,N_47015,N_47903);
and U48467 (N_48467,N_47849,N_47838);
and U48468 (N_48468,N_47157,N_47443);
and U48469 (N_48469,N_47779,N_47619);
xor U48470 (N_48470,N_47683,N_47341);
or U48471 (N_48471,N_47173,N_47714);
or U48472 (N_48472,N_47259,N_47273);
xor U48473 (N_48473,N_47436,N_47654);
and U48474 (N_48474,N_47955,N_47404);
nand U48475 (N_48475,N_47793,N_47251);
or U48476 (N_48476,N_47315,N_47435);
and U48477 (N_48477,N_47923,N_47465);
nand U48478 (N_48478,N_47565,N_47298);
xnor U48479 (N_48479,N_47241,N_47228);
nor U48480 (N_48480,N_47381,N_47358);
or U48481 (N_48481,N_47599,N_47429);
xnor U48482 (N_48482,N_47530,N_47074);
nor U48483 (N_48483,N_47108,N_47895);
xor U48484 (N_48484,N_47071,N_47852);
and U48485 (N_48485,N_47375,N_47653);
nor U48486 (N_48486,N_47769,N_47674);
nand U48487 (N_48487,N_47192,N_47061);
xor U48488 (N_48488,N_47046,N_47270);
or U48489 (N_48489,N_47005,N_47931);
xnor U48490 (N_48490,N_47709,N_47303);
and U48491 (N_48491,N_47177,N_47629);
or U48492 (N_48492,N_47693,N_47863);
xor U48493 (N_48493,N_47308,N_47786);
or U48494 (N_48494,N_47702,N_47230);
nand U48495 (N_48495,N_47051,N_47001);
or U48496 (N_48496,N_47747,N_47840);
nor U48497 (N_48497,N_47373,N_47781);
and U48498 (N_48498,N_47285,N_47932);
nor U48499 (N_48499,N_47497,N_47651);
xnor U48500 (N_48500,N_47729,N_47174);
and U48501 (N_48501,N_47379,N_47634);
or U48502 (N_48502,N_47917,N_47024);
or U48503 (N_48503,N_47700,N_47887);
xnor U48504 (N_48504,N_47214,N_47688);
nand U48505 (N_48505,N_47420,N_47730);
or U48506 (N_48506,N_47028,N_47119);
xnor U48507 (N_48507,N_47694,N_47349);
nor U48508 (N_48508,N_47850,N_47858);
or U48509 (N_48509,N_47365,N_47127);
or U48510 (N_48510,N_47427,N_47372);
xnor U48511 (N_48511,N_47336,N_47430);
xnor U48512 (N_48512,N_47845,N_47577);
nor U48513 (N_48513,N_47055,N_47878);
and U48514 (N_48514,N_47547,N_47812);
xnor U48515 (N_48515,N_47460,N_47495);
nor U48516 (N_48516,N_47826,N_47788);
and U48517 (N_48517,N_47443,N_47509);
nand U48518 (N_48518,N_47210,N_47397);
and U48519 (N_48519,N_47568,N_47723);
xor U48520 (N_48520,N_47430,N_47904);
nor U48521 (N_48521,N_47312,N_47256);
nor U48522 (N_48522,N_47907,N_47588);
nand U48523 (N_48523,N_47809,N_47741);
and U48524 (N_48524,N_47281,N_47148);
and U48525 (N_48525,N_47915,N_47793);
nand U48526 (N_48526,N_47831,N_47022);
nand U48527 (N_48527,N_47730,N_47617);
nand U48528 (N_48528,N_47591,N_47990);
nor U48529 (N_48529,N_47555,N_47397);
or U48530 (N_48530,N_47839,N_47447);
or U48531 (N_48531,N_47464,N_47668);
nand U48532 (N_48532,N_47867,N_47017);
xnor U48533 (N_48533,N_47626,N_47464);
xnor U48534 (N_48534,N_47774,N_47602);
nand U48535 (N_48535,N_47869,N_47928);
and U48536 (N_48536,N_47468,N_47737);
nor U48537 (N_48537,N_47519,N_47596);
xnor U48538 (N_48538,N_47649,N_47326);
nor U48539 (N_48539,N_47251,N_47179);
or U48540 (N_48540,N_47473,N_47783);
and U48541 (N_48541,N_47215,N_47897);
xor U48542 (N_48542,N_47007,N_47318);
nand U48543 (N_48543,N_47039,N_47572);
xnor U48544 (N_48544,N_47209,N_47681);
xnor U48545 (N_48545,N_47772,N_47229);
and U48546 (N_48546,N_47975,N_47840);
or U48547 (N_48547,N_47496,N_47601);
and U48548 (N_48548,N_47922,N_47892);
nor U48549 (N_48549,N_47338,N_47507);
nor U48550 (N_48550,N_47940,N_47154);
and U48551 (N_48551,N_47956,N_47035);
or U48552 (N_48552,N_47435,N_47928);
nor U48553 (N_48553,N_47888,N_47957);
nand U48554 (N_48554,N_47646,N_47299);
and U48555 (N_48555,N_47277,N_47437);
nor U48556 (N_48556,N_47946,N_47068);
nand U48557 (N_48557,N_47971,N_47645);
xnor U48558 (N_48558,N_47084,N_47173);
nand U48559 (N_48559,N_47679,N_47013);
nor U48560 (N_48560,N_47932,N_47486);
and U48561 (N_48561,N_47891,N_47100);
nor U48562 (N_48562,N_47811,N_47359);
nand U48563 (N_48563,N_47484,N_47149);
nand U48564 (N_48564,N_47530,N_47023);
or U48565 (N_48565,N_47271,N_47008);
nand U48566 (N_48566,N_47850,N_47723);
and U48567 (N_48567,N_47939,N_47171);
nor U48568 (N_48568,N_47959,N_47349);
and U48569 (N_48569,N_47964,N_47687);
or U48570 (N_48570,N_47388,N_47252);
nor U48571 (N_48571,N_47935,N_47841);
nor U48572 (N_48572,N_47009,N_47064);
and U48573 (N_48573,N_47416,N_47792);
or U48574 (N_48574,N_47565,N_47931);
nor U48575 (N_48575,N_47740,N_47281);
nand U48576 (N_48576,N_47067,N_47667);
xor U48577 (N_48577,N_47847,N_47493);
xnor U48578 (N_48578,N_47572,N_47875);
nor U48579 (N_48579,N_47818,N_47668);
and U48580 (N_48580,N_47893,N_47445);
or U48581 (N_48581,N_47352,N_47454);
nand U48582 (N_48582,N_47005,N_47738);
and U48583 (N_48583,N_47336,N_47531);
or U48584 (N_48584,N_47150,N_47653);
xnor U48585 (N_48585,N_47718,N_47132);
and U48586 (N_48586,N_47914,N_47665);
and U48587 (N_48587,N_47950,N_47768);
nor U48588 (N_48588,N_47680,N_47239);
or U48589 (N_48589,N_47942,N_47493);
nand U48590 (N_48590,N_47772,N_47990);
nor U48591 (N_48591,N_47101,N_47938);
nor U48592 (N_48592,N_47479,N_47012);
nand U48593 (N_48593,N_47311,N_47950);
nor U48594 (N_48594,N_47493,N_47014);
and U48595 (N_48595,N_47492,N_47908);
nand U48596 (N_48596,N_47065,N_47221);
nand U48597 (N_48597,N_47302,N_47537);
xnor U48598 (N_48598,N_47021,N_47269);
or U48599 (N_48599,N_47297,N_47588);
xnor U48600 (N_48600,N_47434,N_47844);
nor U48601 (N_48601,N_47961,N_47942);
nand U48602 (N_48602,N_47822,N_47197);
xnor U48603 (N_48603,N_47801,N_47845);
nand U48604 (N_48604,N_47157,N_47468);
and U48605 (N_48605,N_47809,N_47225);
and U48606 (N_48606,N_47921,N_47544);
xnor U48607 (N_48607,N_47620,N_47600);
xnor U48608 (N_48608,N_47409,N_47315);
nand U48609 (N_48609,N_47795,N_47889);
nor U48610 (N_48610,N_47730,N_47674);
nor U48611 (N_48611,N_47106,N_47893);
or U48612 (N_48612,N_47876,N_47779);
nor U48613 (N_48613,N_47940,N_47048);
and U48614 (N_48614,N_47120,N_47285);
nor U48615 (N_48615,N_47593,N_47321);
nor U48616 (N_48616,N_47997,N_47414);
nand U48617 (N_48617,N_47599,N_47551);
nor U48618 (N_48618,N_47818,N_47889);
xnor U48619 (N_48619,N_47154,N_47114);
and U48620 (N_48620,N_47578,N_47961);
nor U48621 (N_48621,N_47177,N_47662);
nor U48622 (N_48622,N_47984,N_47838);
and U48623 (N_48623,N_47795,N_47258);
xnor U48624 (N_48624,N_47801,N_47037);
nor U48625 (N_48625,N_47184,N_47192);
or U48626 (N_48626,N_47857,N_47497);
or U48627 (N_48627,N_47100,N_47162);
nand U48628 (N_48628,N_47386,N_47643);
nor U48629 (N_48629,N_47845,N_47128);
nor U48630 (N_48630,N_47241,N_47651);
and U48631 (N_48631,N_47668,N_47732);
xor U48632 (N_48632,N_47039,N_47224);
and U48633 (N_48633,N_47925,N_47281);
and U48634 (N_48634,N_47817,N_47934);
and U48635 (N_48635,N_47823,N_47673);
or U48636 (N_48636,N_47481,N_47359);
or U48637 (N_48637,N_47681,N_47511);
nand U48638 (N_48638,N_47544,N_47414);
xnor U48639 (N_48639,N_47832,N_47244);
or U48640 (N_48640,N_47253,N_47734);
and U48641 (N_48641,N_47398,N_47049);
and U48642 (N_48642,N_47857,N_47784);
nor U48643 (N_48643,N_47109,N_47830);
nand U48644 (N_48644,N_47217,N_47673);
xnor U48645 (N_48645,N_47160,N_47001);
nand U48646 (N_48646,N_47312,N_47460);
xnor U48647 (N_48647,N_47715,N_47952);
or U48648 (N_48648,N_47651,N_47844);
xor U48649 (N_48649,N_47124,N_47938);
and U48650 (N_48650,N_47522,N_47925);
nor U48651 (N_48651,N_47669,N_47668);
nor U48652 (N_48652,N_47167,N_47442);
and U48653 (N_48653,N_47165,N_47101);
nand U48654 (N_48654,N_47025,N_47389);
nor U48655 (N_48655,N_47881,N_47445);
or U48656 (N_48656,N_47374,N_47626);
and U48657 (N_48657,N_47451,N_47591);
nand U48658 (N_48658,N_47130,N_47961);
and U48659 (N_48659,N_47802,N_47924);
xnor U48660 (N_48660,N_47692,N_47697);
nand U48661 (N_48661,N_47725,N_47752);
or U48662 (N_48662,N_47560,N_47123);
nor U48663 (N_48663,N_47709,N_47866);
or U48664 (N_48664,N_47025,N_47292);
nor U48665 (N_48665,N_47800,N_47357);
or U48666 (N_48666,N_47870,N_47540);
nor U48667 (N_48667,N_47072,N_47901);
or U48668 (N_48668,N_47858,N_47133);
nor U48669 (N_48669,N_47989,N_47442);
nor U48670 (N_48670,N_47674,N_47204);
xnor U48671 (N_48671,N_47031,N_47580);
xor U48672 (N_48672,N_47340,N_47864);
or U48673 (N_48673,N_47046,N_47484);
and U48674 (N_48674,N_47327,N_47335);
nand U48675 (N_48675,N_47234,N_47741);
nand U48676 (N_48676,N_47363,N_47717);
or U48677 (N_48677,N_47109,N_47475);
xor U48678 (N_48678,N_47587,N_47973);
and U48679 (N_48679,N_47932,N_47997);
and U48680 (N_48680,N_47553,N_47537);
and U48681 (N_48681,N_47259,N_47080);
xor U48682 (N_48682,N_47088,N_47118);
nor U48683 (N_48683,N_47525,N_47174);
nor U48684 (N_48684,N_47556,N_47152);
and U48685 (N_48685,N_47491,N_47390);
nand U48686 (N_48686,N_47231,N_47860);
and U48687 (N_48687,N_47277,N_47898);
nand U48688 (N_48688,N_47931,N_47469);
and U48689 (N_48689,N_47333,N_47469);
xnor U48690 (N_48690,N_47308,N_47163);
nor U48691 (N_48691,N_47608,N_47182);
nand U48692 (N_48692,N_47813,N_47521);
xor U48693 (N_48693,N_47310,N_47877);
xnor U48694 (N_48694,N_47933,N_47192);
or U48695 (N_48695,N_47718,N_47353);
and U48696 (N_48696,N_47941,N_47670);
nand U48697 (N_48697,N_47736,N_47826);
nor U48698 (N_48698,N_47331,N_47958);
xor U48699 (N_48699,N_47132,N_47698);
nor U48700 (N_48700,N_47274,N_47731);
xnor U48701 (N_48701,N_47078,N_47492);
xor U48702 (N_48702,N_47961,N_47394);
nand U48703 (N_48703,N_47357,N_47297);
and U48704 (N_48704,N_47109,N_47680);
xnor U48705 (N_48705,N_47332,N_47238);
xnor U48706 (N_48706,N_47560,N_47580);
xor U48707 (N_48707,N_47615,N_47892);
xor U48708 (N_48708,N_47911,N_47734);
nand U48709 (N_48709,N_47610,N_47615);
nand U48710 (N_48710,N_47889,N_47694);
xor U48711 (N_48711,N_47142,N_47240);
xnor U48712 (N_48712,N_47547,N_47581);
nand U48713 (N_48713,N_47516,N_47673);
and U48714 (N_48714,N_47691,N_47181);
nand U48715 (N_48715,N_47049,N_47816);
nand U48716 (N_48716,N_47816,N_47301);
or U48717 (N_48717,N_47035,N_47256);
xor U48718 (N_48718,N_47743,N_47116);
or U48719 (N_48719,N_47944,N_47894);
or U48720 (N_48720,N_47036,N_47621);
and U48721 (N_48721,N_47107,N_47882);
nor U48722 (N_48722,N_47282,N_47676);
nand U48723 (N_48723,N_47201,N_47404);
or U48724 (N_48724,N_47419,N_47848);
and U48725 (N_48725,N_47146,N_47588);
or U48726 (N_48726,N_47158,N_47302);
or U48727 (N_48727,N_47960,N_47799);
nor U48728 (N_48728,N_47287,N_47548);
xor U48729 (N_48729,N_47549,N_47370);
nand U48730 (N_48730,N_47232,N_47169);
xor U48731 (N_48731,N_47003,N_47390);
and U48732 (N_48732,N_47930,N_47061);
nor U48733 (N_48733,N_47730,N_47720);
nor U48734 (N_48734,N_47125,N_47842);
nor U48735 (N_48735,N_47119,N_47399);
xnor U48736 (N_48736,N_47773,N_47450);
nand U48737 (N_48737,N_47629,N_47938);
xor U48738 (N_48738,N_47083,N_47818);
nand U48739 (N_48739,N_47584,N_47556);
nand U48740 (N_48740,N_47080,N_47654);
nor U48741 (N_48741,N_47826,N_47428);
or U48742 (N_48742,N_47428,N_47637);
nor U48743 (N_48743,N_47423,N_47906);
nand U48744 (N_48744,N_47827,N_47073);
nor U48745 (N_48745,N_47253,N_47087);
or U48746 (N_48746,N_47688,N_47124);
nand U48747 (N_48747,N_47189,N_47889);
nor U48748 (N_48748,N_47766,N_47287);
nand U48749 (N_48749,N_47368,N_47225);
nor U48750 (N_48750,N_47658,N_47850);
nand U48751 (N_48751,N_47741,N_47852);
xnor U48752 (N_48752,N_47257,N_47657);
and U48753 (N_48753,N_47670,N_47330);
and U48754 (N_48754,N_47485,N_47255);
xnor U48755 (N_48755,N_47079,N_47560);
nand U48756 (N_48756,N_47993,N_47668);
or U48757 (N_48757,N_47793,N_47043);
or U48758 (N_48758,N_47036,N_47920);
and U48759 (N_48759,N_47438,N_47142);
nand U48760 (N_48760,N_47329,N_47383);
or U48761 (N_48761,N_47226,N_47522);
xor U48762 (N_48762,N_47041,N_47738);
and U48763 (N_48763,N_47231,N_47734);
nand U48764 (N_48764,N_47106,N_47585);
and U48765 (N_48765,N_47568,N_47837);
xor U48766 (N_48766,N_47250,N_47242);
or U48767 (N_48767,N_47738,N_47873);
nor U48768 (N_48768,N_47292,N_47464);
and U48769 (N_48769,N_47484,N_47985);
nand U48770 (N_48770,N_47372,N_47473);
xor U48771 (N_48771,N_47892,N_47734);
nor U48772 (N_48772,N_47518,N_47710);
and U48773 (N_48773,N_47529,N_47736);
or U48774 (N_48774,N_47288,N_47323);
and U48775 (N_48775,N_47775,N_47342);
nand U48776 (N_48776,N_47174,N_47465);
nand U48777 (N_48777,N_47189,N_47988);
and U48778 (N_48778,N_47410,N_47010);
xor U48779 (N_48779,N_47109,N_47579);
xnor U48780 (N_48780,N_47525,N_47925);
and U48781 (N_48781,N_47822,N_47347);
nand U48782 (N_48782,N_47140,N_47762);
nor U48783 (N_48783,N_47776,N_47652);
nand U48784 (N_48784,N_47464,N_47854);
nor U48785 (N_48785,N_47290,N_47688);
xor U48786 (N_48786,N_47425,N_47196);
and U48787 (N_48787,N_47630,N_47513);
nor U48788 (N_48788,N_47692,N_47537);
nor U48789 (N_48789,N_47047,N_47892);
nand U48790 (N_48790,N_47749,N_47004);
xnor U48791 (N_48791,N_47648,N_47199);
or U48792 (N_48792,N_47498,N_47359);
nand U48793 (N_48793,N_47742,N_47832);
nor U48794 (N_48794,N_47506,N_47816);
nor U48795 (N_48795,N_47774,N_47620);
nor U48796 (N_48796,N_47817,N_47383);
and U48797 (N_48797,N_47143,N_47122);
nand U48798 (N_48798,N_47412,N_47935);
and U48799 (N_48799,N_47188,N_47796);
nand U48800 (N_48800,N_47215,N_47127);
nor U48801 (N_48801,N_47811,N_47750);
xnor U48802 (N_48802,N_47708,N_47004);
nor U48803 (N_48803,N_47604,N_47686);
nand U48804 (N_48804,N_47078,N_47240);
or U48805 (N_48805,N_47439,N_47755);
or U48806 (N_48806,N_47645,N_47711);
and U48807 (N_48807,N_47941,N_47077);
or U48808 (N_48808,N_47935,N_47394);
nor U48809 (N_48809,N_47237,N_47189);
and U48810 (N_48810,N_47618,N_47286);
nand U48811 (N_48811,N_47922,N_47728);
or U48812 (N_48812,N_47687,N_47977);
or U48813 (N_48813,N_47451,N_47231);
xnor U48814 (N_48814,N_47187,N_47748);
and U48815 (N_48815,N_47822,N_47587);
nand U48816 (N_48816,N_47989,N_47305);
or U48817 (N_48817,N_47030,N_47153);
nand U48818 (N_48818,N_47627,N_47934);
nor U48819 (N_48819,N_47630,N_47416);
nor U48820 (N_48820,N_47746,N_47895);
nand U48821 (N_48821,N_47654,N_47689);
nor U48822 (N_48822,N_47922,N_47134);
xor U48823 (N_48823,N_47215,N_47233);
nor U48824 (N_48824,N_47633,N_47717);
nand U48825 (N_48825,N_47800,N_47925);
nor U48826 (N_48826,N_47589,N_47888);
nand U48827 (N_48827,N_47384,N_47619);
and U48828 (N_48828,N_47979,N_47394);
xnor U48829 (N_48829,N_47941,N_47982);
and U48830 (N_48830,N_47274,N_47576);
nor U48831 (N_48831,N_47810,N_47132);
or U48832 (N_48832,N_47917,N_47827);
or U48833 (N_48833,N_47871,N_47395);
nor U48834 (N_48834,N_47893,N_47160);
nand U48835 (N_48835,N_47322,N_47835);
nand U48836 (N_48836,N_47315,N_47237);
and U48837 (N_48837,N_47539,N_47491);
xor U48838 (N_48838,N_47351,N_47111);
or U48839 (N_48839,N_47353,N_47992);
and U48840 (N_48840,N_47648,N_47222);
or U48841 (N_48841,N_47501,N_47775);
xor U48842 (N_48842,N_47282,N_47326);
nor U48843 (N_48843,N_47811,N_47201);
nor U48844 (N_48844,N_47785,N_47702);
xnor U48845 (N_48845,N_47036,N_47176);
xor U48846 (N_48846,N_47084,N_47051);
or U48847 (N_48847,N_47255,N_47565);
nor U48848 (N_48848,N_47849,N_47142);
xor U48849 (N_48849,N_47255,N_47544);
xnor U48850 (N_48850,N_47773,N_47622);
nand U48851 (N_48851,N_47133,N_47495);
xnor U48852 (N_48852,N_47435,N_47762);
xor U48853 (N_48853,N_47132,N_47916);
nor U48854 (N_48854,N_47412,N_47896);
or U48855 (N_48855,N_47349,N_47742);
xor U48856 (N_48856,N_47903,N_47374);
xor U48857 (N_48857,N_47105,N_47547);
nor U48858 (N_48858,N_47342,N_47092);
nor U48859 (N_48859,N_47064,N_47626);
and U48860 (N_48860,N_47193,N_47890);
and U48861 (N_48861,N_47293,N_47949);
nor U48862 (N_48862,N_47415,N_47169);
or U48863 (N_48863,N_47779,N_47815);
or U48864 (N_48864,N_47388,N_47357);
nand U48865 (N_48865,N_47784,N_47344);
nand U48866 (N_48866,N_47704,N_47904);
nand U48867 (N_48867,N_47464,N_47411);
or U48868 (N_48868,N_47153,N_47657);
or U48869 (N_48869,N_47273,N_47961);
nand U48870 (N_48870,N_47270,N_47695);
nor U48871 (N_48871,N_47876,N_47665);
and U48872 (N_48872,N_47331,N_47038);
or U48873 (N_48873,N_47421,N_47689);
nor U48874 (N_48874,N_47045,N_47187);
nor U48875 (N_48875,N_47940,N_47868);
or U48876 (N_48876,N_47175,N_47101);
nor U48877 (N_48877,N_47874,N_47767);
xnor U48878 (N_48878,N_47392,N_47932);
or U48879 (N_48879,N_47609,N_47999);
or U48880 (N_48880,N_47001,N_47607);
or U48881 (N_48881,N_47642,N_47734);
nand U48882 (N_48882,N_47703,N_47957);
and U48883 (N_48883,N_47600,N_47035);
xnor U48884 (N_48884,N_47297,N_47711);
xor U48885 (N_48885,N_47584,N_47118);
or U48886 (N_48886,N_47104,N_47926);
and U48887 (N_48887,N_47545,N_47101);
xor U48888 (N_48888,N_47856,N_47756);
xnor U48889 (N_48889,N_47387,N_47574);
nor U48890 (N_48890,N_47754,N_47217);
nand U48891 (N_48891,N_47067,N_47996);
or U48892 (N_48892,N_47792,N_47046);
xnor U48893 (N_48893,N_47973,N_47055);
and U48894 (N_48894,N_47944,N_47734);
and U48895 (N_48895,N_47531,N_47063);
xnor U48896 (N_48896,N_47847,N_47619);
and U48897 (N_48897,N_47734,N_47422);
nor U48898 (N_48898,N_47208,N_47572);
nand U48899 (N_48899,N_47821,N_47482);
nor U48900 (N_48900,N_47111,N_47712);
and U48901 (N_48901,N_47766,N_47750);
or U48902 (N_48902,N_47520,N_47947);
and U48903 (N_48903,N_47606,N_47715);
or U48904 (N_48904,N_47623,N_47661);
nor U48905 (N_48905,N_47443,N_47481);
nand U48906 (N_48906,N_47593,N_47154);
and U48907 (N_48907,N_47695,N_47085);
or U48908 (N_48908,N_47036,N_47885);
nor U48909 (N_48909,N_47455,N_47296);
nand U48910 (N_48910,N_47480,N_47983);
nor U48911 (N_48911,N_47022,N_47602);
xor U48912 (N_48912,N_47454,N_47167);
or U48913 (N_48913,N_47104,N_47010);
xnor U48914 (N_48914,N_47225,N_47924);
and U48915 (N_48915,N_47139,N_47906);
or U48916 (N_48916,N_47284,N_47609);
or U48917 (N_48917,N_47182,N_47711);
and U48918 (N_48918,N_47641,N_47577);
or U48919 (N_48919,N_47896,N_47871);
and U48920 (N_48920,N_47142,N_47073);
nor U48921 (N_48921,N_47367,N_47819);
nor U48922 (N_48922,N_47648,N_47287);
nand U48923 (N_48923,N_47498,N_47649);
xor U48924 (N_48924,N_47355,N_47910);
and U48925 (N_48925,N_47667,N_47081);
xor U48926 (N_48926,N_47400,N_47133);
xnor U48927 (N_48927,N_47949,N_47766);
nor U48928 (N_48928,N_47216,N_47301);
and U48929 (N_48929,N_47988,N_47479);
nand U48930 (N_48930,N_47163,N_47483);
nor U48931 (N_48931,N_47009,N_47574);
and U48932 (N_48932,N_47051,N_47859);
and U48933 (N_48933,N_47233,N_47694);
and U48934 (N_48934,N_47424,N_47860);
nand U48935 (N_48935,N_47606,N_47796);
nor U48936 (N_48936,N_47006,N_47373);
xnor U48937 (N_48937,N_47814,N_47921);
and U48938 (N_48938,N_47592,N_47739);
or U48939 (N_48939,N_47189,N_47762);
xnor U48940 (N_48940,N_47794,N_47585);
or U48941 (N_48941,N_47140,N_47787);
nor U48942 (N_48942,N_47514,N_47702);
nor U48943 (N_48943,N_47359,N_47859);
nand U48944 (N_48944,N_47605,N_47845);
xor U48945 (N_48945,N_47350,N_47896);
xor U48946 (N_48946,N_47156,N_47545);
nor U48947 (N_48947,N_47658,N_47138);
xor U48948 (N_48948,N_47616,N_47716);
nor U48949 (N_48949,N_47333,N_47452);
nor U48950 (N_48950,N_47670,N_47803);
or U48951 (N_48951,N_47203,N_47923);
nand U48952 (N_48952,N_47858,N_47507);
or U48953 (N_48953,N_47501,N_47196);
xnor U48954 (N_48954,N_47975,N_47115);
nor U48955 (N_48955,N_47081,N_47990);
nand U48956 (N_48956,N_47394,N_47366);
nor U48957 (N_48957,N_47920,N_47973);
xor U48958 (N_48958,N_47690,N_47532);
xnor U48959 (N_48959,N_47499,N_47850);
nor U48960 (N_48960,N_47839,N_47043);
xor U48961 (N_48961,N_47726,N_47027);
nand U48962 (N_48962,N_47158,N_47896);
nand U48963 (N_48963,N_47212,N_47651);
and U48964 (N_48964,N_47561,N_47592);
xnor U48965 (N_48965,N_47379,N_47077);
and U48966 (N_48966,N_47196,N_47663);
or U48967 (N_48967,N_47684,N_47093);
and U48968 (N_48968,N_47077,N_47183);
and U48969 (N_48969,N_47385,N_47167);
or U48970 (N_48970,N_47654,N_47583);
xnor U48971 (N_48971,N_47567,N_47737);
nand U48972 (N_48972,N_47749,N_47197);
and U48973 (N_48973,N_47081,N_47861);
xnor U48974 (N_48974,N_47808,N_47076);
and U48975 (N_48975,N_47036,N_47059);
and U48976 (N_48976,N_47865,N_47231);
or U48977 (N_48977,N_47471,N_47935);
nand U48978 (N_48978,N_47738,N_47975);
and U48979 (N_48979,N_47167,N_47870);
nor U48980 (N_48980,N_47971,N_47347);
or U48981 (N_48981,N_47636,N_47656);
xor U48982 (N_48982,N_47469,N_47352);
or U48983 (N_48983,N_47775,N_47336);
xor U48984 (N_48984,N_47202,N_47131);
nor U48985 (N_48985,N_47035,N_47433);
or U48986 (N_48986,N_47636,N_47986);
or U48987 (N_48987,N_47549,N_47747);
nor U48988 (N_48988,N_47249,N_47784);
nand U48989 (N_48989,N_47856,N_47558);
and U48990 (N_48990,N_47237,N_47553);
nand U48991 (N_48991,N_47055,N_47305);
or U48992 (N_48992,N_47732,N_47121);
and U48993 (N_48993,N_47033,N_47918);
or U48994 (N_48994,N_47868,N_47610);
or U48995 (N_48995,N_47470,N_47627);
xnor U48996 (N_48996,N_47424,N_47534);
or U48997 (N_48997,N_47826,N_47919);
nor U48998 (N_48998,N_47317,N_47444);
nand U48999 (N_48999,N_47263,N_47793);
nor U49000 (N_49000,N_48720,N_48361);
nand U49001 (N_49001,N_48200,N_48255);
nand U49002 (N_49002,N_48191,N_48382);
or U49003 (N_49003,N_48489,N_48176);
and U49004 (N_49004,N_48126,N_48083);
and U49005 (N_49005,N_48692,N_48063);
nor U49006 (N_49006,N_48783,N_48959);
and U49007 (N_49007,N_48181,N_48015);
or U49008 (N_49008,N_48158,N_48195);
xor U49009 (N_49009,N_48823,N_48930);
nor U49010 (N_49010,N_48673,N_48737);
and U49011 (N_49011,N_48171,N_48254);
nor U49012 (N_49012,N_48035,N_48584);
xor U49013 (N_49013,N_48424,N_48731);
nand U49014 (N_49014,N_48793,N_48051);
or U49015 (N_49015,N_48878,N_48236);
or U49016 (N_49016,N_48658,N_48438);
nor U49017 (N_49017,N_48198,N_48706);
xnor U49018 (N_49018,N_48767,N_48145);
nand U49019 (N_49019,N_48134,N_48306);
nand U49020 (N_49020,N_48066,N_48642);
nor U49021 (N_49021,N_48507,N_48550);
or U49022 (N_49022,N_48443,N_48968);
or U49023 (N_49023,N_48407,N_48984);
nor U49024 (N_49024,N_48087,N_48262);
and U49025 (N_49025,N_48179,N_48451);
nor U49026 (N_49026,N_48116,N_48532);
or U49027 (N_49027,N_48841,N_48009);
nand U49028 (N_49028,N_48399,N_48142);
nor U49029 (N_49029,N_48265,N_48644);
nor U49030 (N_49030,N_48909,N_48531);
xor U49031 (N_49031,N_48515,N_48668);
nor U49032 (N_49032,N_48359,N_48848);
and U49033 (N_49033,N_48989,N_48798);
nand U49034 (N_49034,N_48659,N_48026);
nor U49035 (N_49035,N_48953,N_48711);
and U49036 (N_49036,N_48772,N_48098);
or U49037 (N_49037,N_48303,N_48390);
or U49038 (N_49038,N_48334,N_48699);
nand U49039 (N_49039,N_48514,N_48824);
and U49040 (N_49040,N_48010,N_48726);
and U49041 (N_49041,N_48627,N_48843);
and U49042 (N_49042,N_48863,N_48937);
xor U49043 (N_49043,N_48712,N_48392);
and U49044 (N_49044,N_48694,N_48975);
or U49045 (N_49045,N_48539,N_48773);
nor U49046 (N_49046,N_48441,N_48394);
nand U49047 (N_49047,N_48639,N_48470);
nand U49048 (N_49048,N_48974,N_48908);
or U49049 (N_49049,N_48876,N_48131);
nor U49050 (N_49050,N_48247,N_48887);
nor U49051 (N_49051,N_48415,N_48319);
nor U49052 (N_49052,N_48840,N_48282);
nor U49053 (N_49053,N_48916,N_48224);
nor U49054 (N_49054,N_48956,N_48913);
nor U49055 (N_49055,N_48799,N_48256);
nor U49056 (N_49056,N_48226,N_48881);
nor U49057 (N_49057,N_48425,N_48696);
nor U49058 (N_49058,N_48803,N_48329);
nor U49059 (N_49059,N_48091,N_48251);
nand U49060 (N_49060,N_48951,N_48853);
xor U49061 (N_49061,N_48914,N_48092);
and U49062 (N_49062,N_48463,N_48095);
xnor U49063 (N_49063,N_48367,N_48419);
xor U49064 (N_49064,N_48014,N_48175);
or U49065 (N_49065,N_48002,N_48194);
nor U49066 (N_49066,N_48442,N_48779);
nand U49067 (N_49067,N_48429,N_48990);
and U49068 (N_49068,N_48704,N_48384);
nand U49069 (N_49069,N_48374,N_48548);
and U49070 (N_49070,N_48789,N_48741);
and U49071 (N_49071,N_48048,N_48343);
xor U49072 (N_49072,N_48237,N_48202);
or U49073 (N_49073,N_48437,N_48647);
nor U49074 (N_49074,N_48906,N_48148);
or U49075 (N_49075,N_48447,N_48743);
or U49076 (N_49076,N_48894,N_48184);
or U49077 (N_49077,N_48677,N_48089);
xnor U49078 (N_49078,N_48345,N_48635);
nand U49079 (N_49079,N_48431,N_48593);
and U49080 (N_49080,N_48983,N_48925);
nand U49081 (N_49081,N_48121,N_48307);
xor U49082 (N_49082,N_48378,N_48281);
and U49083 (N_49083,N_48756,N_48153);
and U49084 (N_49084,N_48457,N_48551);
and U49085 (N_49085,N_48868,N_48032);
or U49086 (N_49086,N_48228,N_48041);
or U49087 (N_49087,N_48820,N_48729);
nand U49088 (N_49088,N_48701,N_48280);
xnor U49089 (N_49089,N_48341,N_48004);
xnor U49090 (N_49090,N_48948,N_48498);
nand U49091 (N_49091,N_48263,N_48864);
or U49092 (N_49092,N_48826,N_48537);
xnor U49093 (N_49093,N_48398,N_48420);
or U49094 (N_49094,N_48664,N_48033);
nand U49095 (N_49095,N_48613,N_48269);
nand U49096 (N_49096,N_48223,N_48490);
xor U49097 (N_49097,N_48193,N_48240);
nand U49098 (N_49098,N_48053,N_48751);
and U49099 (N_49099,N_48060,N_48935);
xnor U49100 (N_49100,N_48558,N_48369);
or U49101 (N_49101,N_48244,N_48528);
and U49102 (N_49102,N_48735,N_48318);
nand U49103 (N_49103,N_48112,N_48533);
and U49104 (N_49104,N_48631,N_48513);
xor U49105 (N_49105,N_48534,N_48747);
and U49106 (N_49106,N_48172,N_48596);
or U49107 (N_49107,N_48745,N_48574);
xor U49108 (N_49108,N_48468,N_48554);
nor U49109 (N_49109,N_48454,N_48999);
nor U49110 (N_49110,N_48353,N_48402);
nand U49111 (N_49111,N_48527,N_48671);
and U49112 (N_49112,N_48233,N_48589);
nand U49113 (N_49113,N_48972,N_48072);
nand U49114 (N_49114,N_48362,N_48922);
nand U49115 (N_49115,N_48850,N_48595);
or U49116 (N_49116,N_48872,N_48510);
nor U49117 (N_49117,N_48070,N_48225);
nor U49118 (N_49118,N_48466,N_48620);
and U49119 (N_49119,N_48117,N_48727);
nand U49120 (N_49120,N_48264,N_48844);
nor U49121 (N_49121,N_48765,N_48292);
and U49122 (N_49122,N_48942,N_48832);
or U49123 (N_49123,N_48414,N_48078);
nor U49124 (N_49124,N_48366,N_48499);
or U49125 (N_49125,N_48340,N_48312);
or U49126 (N_49126,N_48884,N_48757);
and U49127 (N_49127,N_48350,N_48276);
xor U49128 (N_49128,N_48649,N_48025);
nor U49129 (N_49129,N_48376,N_48006);
or U49130 (N_49130,N_48617,N_48661);
and U49131 (N_49131,N_48128,N_48849);
and U49132 (N_49132,N_48847,N_48991);
and U49133 (N_49133,N_48569,N_48001);
nand U49134 (N_49134,N_48188,N_48234);
nor U49135 (N_49135,N_48215,N_48963);
nor U49136 (N_49136,N_48971,N_48081);
nand U49137 (N_49137,N_48260,N_48064);
or U49138 (N_49138,N_48640,N_48875);
nand U49139 (N_49139,N_48055,N_48150);
and U49140 (N_49140,N_48509,N_48748);
nand U49141 (N_49141,N_48337,N_48433);
xnor U49142 (N_49142,N_48903,N_48713);
and U49143 (N_49143,N_48855,N_48688);
or U49144 (N_49144,N_48401,N_48759);
xnor U49145 (N_49145,N_48493,N_48090);
or U49146 (N_49146,N_48299,N_48427);
or U49147 (N_49147,N_48812,N_48829);
and U49148 (N_49148,N_48612,N_48780);
nand U49149 (N_49149,N_48452,N_48594);
or U49150 (N_49150,N_48607,N_48143);
and U49151 (N_49151,N_48185,N_48119);
or U49152 (N_49152,N_48039,N_48506);
xnor U49153 (N_49153,N_48173,N_48679);
and U49154 (N_49154,N_48600,N_48159);
nand U49155 (N_49155,N_48921,N_48544);
nand U49156 (N_49156,N_48183,N_48027);
xor U49157 (N_49157,N_48615,N_48710);
nand U49158 (N_49158,N_48044,N_48007);
and U49159 (N_49159,N_48208,N_48725);
nand U49160 (N_49160,N_48705,N_48118);
or U49161 (N_49161,N_48302,N_48245);
nor U49162 (N_49162,N_48439,N_48397);
or U49163 (N_49163,N_48738,N_48178);
nand U49164 (N_49164,N_48106,N_48568);
nand U49165 (N_49165,N_48858,N_48645);
and U49166 (N_49166,N_48272,N_48124);
nand U49167 (N_49167,N_48651,N_48152);
nor U49168 (N_49168,N_48683,N_48634);
xnor U49169 (N_49169,N_48180,N_48213);
nor U49170 (N_49170,N_48034,N_48235);
or U49171 (N_49171,N_48348,N_48444);
xor U49172 (N_49172,N_48491,N_48804);
nor U49173 (N_49173,N_48132,N_48721);
nor U49174 (N_49174,N_48416,N_48549);
or U49175 (N_49175,N_48708,N_48286);
nor U49176 (N_49176,N_48831,N_48502);
or U49177 (N_49177,N_48943,N_48949);
nand U49178 (N_49178,N_48723,N_48603);
nand U49179 (N_49179,N_48771,N_48834);
nand U49180 (N_49180,N_48564,N_48088);
and U49181 (N_49181,N_48845,N_48981);
xor U49182 (N_49182,N_48022,N_48579);
xor U49183 (N_49183,N_48786,N_48618);
or U49184 (N_49184,N_48811,N_48776);
and U49185 (N_49185,N_48883,N_48998);
nor U49186 (N_49186,N_48562,N_48879);
nand U49187 (N_49187,N_48209,N_48573);
nand U49188 (N_49188,N_48426,N_48859);
or U49189 (N_49189,N_48516,N_48403);
and U49190 (N_49190,N_48870,N_48258);
and U49191 (N_49191,N_48626,N_48717);
nor U49192 (N_49192,N_48216,N_48962);
and U49193 (N_49193,N_48332,N_48144);
nand U49194 (N_49194,N_48604,N_48151);
nand U49195 (N_49195,N_48952,N_48763);
xor U49196 (N_49196,N_48842,N_48321);
xnor U49197 (N_49197,N_48471,N_48678);
or U49198 (N_49198,N_48339,N_48459);
nor U49199 (N_49199,N_48475,N_48838);
nor U49200 (N_49200,N_48917,N_48702);
nand U49201 (N_49201,N_48630,N_48775);
xnor U49202 (N_49202,N_48120,N_48156);
and U49203 (N_49203,N_48028,N_48524);
and U49204 (N_49204,N_48781,N_48016);
nor U49205 (N_49205,N_48555,N_48650);
or U49206 (N_49206,N_48000,N_48423);
or U49207 (N_49207,N_48168,N_48581);
and U49208 (N_49208,N_48774,N_48778);
xnor U49209 (N_49209,N_48129,N_48375);
nand U49210 (N_49210,N_48421,N_48695);
and U49211 (N_49211,N_48076,N_48800);
xnor U49212 (N_49212,N_48816,N_48289);
nor U49213 (N_49213,N_48483,N_48389);
and U49214 (N_49214,N_48099,N_48291);
or U49215 (N_49215,N_48261,N_48749);
and U49216 (N_49216,N_48199,N_48163);
or U49217 (N_49217,N_48586,N_48204);
nor U49218 (N_49218,N_48703,N_48744);
and U49219 (N_49219,N_48785,N_48123);
xor U49220 (N_49220,N_48283,N_48485);
nor U49221 (N_49221,N_48391,N_48995);
nor U49222 (N_49222,N_48680,N_48525);
nand U49223 (N_49223,N_48760,N_48246);
and U49224 (N_49224,N_48685,N_48154);
or U49225 (N_49225,N_48297,N_48212);
xor U49226 (N_49226,N_48050,N_48986);
nor U49227 (N_49227,N_48249,N_48395);
or U49228 (N_49228,N_48857,N_48895);
or U49229 (N_49229,N_48275,N_48988);
nand U49230 (N_49230,N_48632,N_48082);
or U49231 (N_49231,N_48764,N_48753);
or U49232 (N_49232,N_48157,N_48492);
or U49233 (N_49233,N_48886,N_48500);
and U49234 (N_49234,N_48363,N_48461);
or U49235 (N_49235,N_48977,N_48540);
nor U49236 (N_49236,N_48349,N_48802);
nand U49237 (N_49237,N_48381,N_48325);
xor U49238 (N_49238,N_48924,N_48357);
nand U49239 (N_49239,N_48517,N_48961);
or U49240 (N_49240,N_48578,N_48323);
xor U49241 (N_49241,N_48835,N_48274);
and U49242 (N_49242,N_48238,N_48370);
or U49243 (N_49243,N_48206,N_48149);
nor U49244 (N_49244,N_48239,N_48700);
nand U49245 (N_49245,N_48970,N_48445);
and U49246 (N_49246,N_48583,N_48522);
nor U49247 (N_49247,N_48122,N_48130);
or U49248 (N_49248,N_48428,N_48511);
xnor U49249 (N_49249,N_48331,N_48590);
nand U49250 (N_49250,N_48690,N_48587);
nand U49251 (N_49251,N_48455,N_48839);
and U49252 (N_49252,N_48681,N_48293);
xor U49253 (N_49253,N_48890,N_48371);
or U49254 (N_49254,N_48993,N_48309);
and U49255 (N_49255,N_48766,N_48203);
nor U49256 (N_49256,N_48477,N_48792);
nand U49257 (N_49257,N_48567,N_48487);
nand U49258 (N_49258,N_48248,N_48285);
or U49259 (N_49259,N_48755,N_48065);
or U49260 (N_49260,N_48020,N_48571);
nand U49261 (N_49261,N_48746,N_48434);
nor U49262 (N_49262,N_48563,N_48788);
nand U49263 (N_49263,N_48967,N_48611);
nor U49264 (N_49264,N_48787,N_48432);
nand U49265 (N_49265,N_48217,N_48889);
nand U49266 (N_49266,N_48404,N_48655);
and U49267 (N_49267,N_48197,N_48139);
xnor U49268 (N_49268,N_48556,N_48624);
and U49269 (N_49269,N_48410,N_48494);
or U49270 (N_49270,N_48547,N_48067);
xnor U49271 (N_49271,N_48104,N_48724);
nor U49272 (N_49272,N_48453,N_48231);
nor U49273 (N_49273,N_48030,N_48940);
xor U49274 (N_49274,N_48059,N_48958);
nand U49275 (N_49275,N_48526,N_48733);
xnor U49276 (N_49276,N_48480,N_48268);
nor U49277 (N_49277,N_48330,N_48808);
and U49278 (N_49278,N_48818,N_48017);
nand U49279 (N_49279,N_48941,N_48406);
nor U49280 (N_49280,N_48114,N_48657);
or U49281 (N_49281,N_48865,N_48662);
nand U49282 (N_49282,N_48653,N_48311);
nand U49283 (N_49283,N_48504,N_48221);
nand U49284 (N_49284,N_48460,N_48828);
nor U49285 (N_49285,N_48997,N_48242);
xnor U49286 (N_49286,N_48021,N_48687);
and U49287 (N_49287,N_48777,N_48230);
xor U49288 (N_49288,N_48086,N_48458);
and U49289 (N_49289,N_48669,N_48011);
and U49290 (N_49290,N_48807,N_48270);
nor U49291 (N_49291,N_48597,N_48310);
and U49292 (N_49292,N_48201,N_48898);
or U49293 (N_49293,N_48938,N_48575);
and U49294 (N_49294,N_48546,N_48521);
and U49295 (N_49295,N_48503,N_48978);
and U49296 (N_49296,N_48638,N_48322);
or U49297 (N_49297,N_48388,N_48486);
nor U49298 (N_49298,N_48969,N_48902);
nor U49299 (N_49299,N_48137,N_48608);
xnor U49300 (N_49300,N_48982,N_48417);
nor U49301 (N_49301,N_48385,N_48860);
or U49302 (N_49302,N_48582,N_48005);
nor U49303 (N_49303,N_48170,N_48147);
and U49304 (N_49304,N_48085,N_48656);
and U49305 (N_49305,N_48232,N_48609);
or U49306 (N_49306,N_48797,N_48430);
nor U49307 (N_49307,N_48979,N_48162);
nand U49308 (N_49308,N_48739,N_48365);
and U49309 (N_49309,N_48450,N_48932);
nand U49310 (N_49310,N_48177,N_48167);
xor U49311 (N_49311,N_48387,N_48934);
nand U49312 (N_49312,N_48919,N_48891);
and U49313 (N_49313,N_48073,N_48610);
and U49314 (N_49314,N_48707,N_48869);
nor U49315 (N_49315,N_48253,N_48192);
nor U49316 (N_49316,N_48880,N_48512);
xnor U49317 (N_49317,N_48619,N_48189);
or U49318 (N_49318,N_48825,N_48409);
and U49319 (N_49319,N_48565,N_48164);
xnor U49320 (N_49320,N_48716,N_48377);
or U49321 (N_49321,N_48910,N_48125);
nand U49322 (N_49322,N_48698,N_48408);
xor U49323 (N_49323,N_48520,N_48623);
xor U49324 (N_49324,N_48740,N_48346);
and U49325 (N_49325,N_48791,N_48637);
xor U49326 (N_49326,N_48046,N_48071);
xnor U49327 (N_49327,N_48304,N_48852);
or U49328 (N_49328,N_48750,N_48560);
nand U49329 (N_49329,N_48393,N_48396);
and U49330 (N_49330,N_48052,N_48300);
or U49331 (N_49331,N_48873,N_48538);
xnor U49332 (N_49332,N_48056,N_48628);
and U49333 (N_49333,N_48945,N_48160);
xor U49334 (N_49334,N_48043,N_48557);
or U49335 (N_49335,N_48418,N_48742);
or U49336 (N_49336,N_48219,N_48572);
nor U49337 (N_49337,N_48278,N_48994);
nor U49338 (N_49338,N_48317,N_48355);
and U49339 (N_49339,N_48874,N_48328);
xnor U49340 (N_49340,N_48709,N_48354);
nand U49341 (N_49341,N_48287,N_48905);
xnor U49342 (N_49342,N_48205,N_48097);
xor U49343 (N_49343,N_48271,N_48758);
and U49344 (N_49344,N_48279,N_48728);
and U49345 (N_49345,N_48754,N_48008);
xor U49346 (N_49346,N_48190,N_48241);
or U49347 (N_49347,N_48652,N_48508);
nand U49348 (N_49348,N_48629,N_48140);
and U49349 (N_49349,N_48599,N_48096);
nand U49350 (N_49350,N_48676,N_48079);
nor U49351 (N_49351,N_48080,N_48057);
or U49352 (N_49352,N_48862,N_48900);
nand U49353 (N_49353,N_48012,N_48102);
xnor U49354 (N_49354,N_48166,N_48111);
nor U49355 (N_49355,N_48719,N_48915);
and U49356 (N_49356,N_48405,N_48411);
and U49357 (N_49357,N_48795,N_48294);
or U49358 (N_49358,N_48288,N_48383);
or U49359 (N_49359,N_48769,N_48936);
nor U49360 (N_49360,N_48552,N_48187);
and U49361 (N_49361,N_48037,N_48955);
or U49362 (N_49362,N_48481,N_48259);
or U49363 (N_49363,N_48062,N_48752);
and U49364 (N_49364,N_48333,N_48672);
nor U49365 (N_49365,N_48069,N_48155);
nand U49366 (N_49366,N_48976,N_48666);
xnor U49367 (N_49367,N_48926,N_48636);
xor U49368 (N_49368,N_48031,N_48602);
xnor U49369 (N_49369,N_48243,N_48836);
nor U49370 (N_49370,N_48736,N_48592);
nand U49371 (N_49371,N_48146,N_48127);
or U49372 (N_49372,N_48290,N_48229);
nor U49373 (N_49373,N_48136,N_48267);
nor U49374 (N_49374,N_48856,N_48478);
or U49375 (N_49375,N_48013,N_48308);
nand U49376 (N_49376,N_48049,N_48686);
or U49377 (N_49377,N_48214,N_48084);
or U49378 (N_49378,N_48985,N_48561);
or U49379 (N_49379,N_48358,N_48211);
nor U49380 (N_49380,N_48591,N_48024);
or U49381 (N_49381,N_48115,N_48058);
xnor U49382 (N_49382,N_48944,N_48814);
xnor U49383 (N_49383,N_48074,N_48622);
xor U49384 (N_49384,N_48135,N_48472);
xnor U49385 (N_49385,N_48412,N_48161);
nor U49386 (N_49386,N_48356,N_48827);
nor U49387 (N_49387,N_48950,N_48250);
nor U49388 (N_49388,N_48380,N_48964);
or U49389 (N_49389,N_48316,N_48360);
xor U49390 (N_49390,N_48833,N_48019);
nor U49391 (N_49391,N_48576,N_48505);
nor U49392 (N_49392,N_48109,N_48815);
xor U49393 (N_49393,N_48851,N_48911);
xnor U49394 (N_49394,N_48641,N_48496);
nor U49395 (N_49395,N_48036,N_48957);
xnor U49396 (N_49396,N_48822,N_48368);
nor U49397 (N_49397,N_48497,N_48542);
xnor U49398 (N_49398,N_48761,N_48675);
xor U49399 (N_49399,N_48456,N_48169);
or U49400 (N_49400,N_48897,N_48352);
and U49401 (N_49401,N_48580,N_48422);
nor U49402 (N_49402,N_48440,N_48061);
or U49403 (N_49403,N_48138,N_48810);
nand U49404 (N_49404,N_48435,N_48042);
xor U49405 (N_49405,N_48519,N_48682);
nand U49406 (N_49406,N_48448,N_48813);
xnor U49407 (N_49407,N_48113,N_48616);
and U49408 (N_49408,N_48819,N_48805);
nor U49409 (N_49409,N_48386,N_48809);
nand U49410 (N_49410,N_48794,N_48186);
xor U49411 (N_49411,N_48877,N_48689);
nor U49412 (N_49412,N_48697,N_48722);
xor U49413 (N_49413,N_48110,N_48347);
nor U49414 (N_49414,N_48469,N_48518);
nor U49415 (N_49415,N_48535,N_48488);
or U49416 (N_49416,N_48830,N_48501);
nand U49417 (N_49417,N_48553,N_48684);
xnor U49418 (N_49418,N_48559,N_48133);
xnor U49419 (N_49419,N_48373,N_48182);
nor U49420 (N_49420,N_48536,N_48482);
nor U49421 (N_49421,N_48654,N_48606);
nand U49422 (N_49422,N_48817,N_48023);
and U49423 (N_49423,N_48077,N_48674);
nand U49424 (N_49424,N_48996,N_48648);
or U49425 (N_49425,N_48670,N_48734);
and U49426 (N_49426,N_48992,N_48577);
xor U49427 (N_49427,N_48108,N_48693);
and U49428 (N_49428,N_48313,N_48837);
nand U49429 (N_49429,N_48888,N_48530);
or U49430 (N_49430,N_48296,N_48326);
or U49431 (N_49431,N_48927,N_48207);
and U49432 (N_49432,N_48920,N_48165);
or U49433 (N_49433,N_48105,N_48342);
nand U49434 (N_49434,N_48107,N_48449);
nor U49435 (N_49435,N_48901,N_48301);
or U49436 (N_49436,N_48933,N_48436);
and U49437 (N_49437,N_48801,N_48273);
and U49438 (N_49438,N_48643,N_48315);
xor U49439 (N_49439,N_48923,N_48103);
or U49440 (N_49440,N_48614,N_48732);
and U49441 (N_49441,N_48464,N_48018);
or U49442 (N_49442,N_48625,N_48196);
nand U49443 (N_49443,N_48529,N_48585);
xor U49444 (N_49444,N_48338,N_48284);
and U49445 (N_49445,N_48954,N_48474);
xor U49446 (N_49446,N_48523,N_48045);
nand U49447 (N_49447,N_48899,N_48928);
xnor U49448 (N_49448,N_48960,N_48227);
and U49449 (N_49449,N_48364,N_48093);
nand U49450 (N_49450,N_48210,N_48413);
nand U49451 (N_49451,N_48570,N_48861);
xnor U49452 (N_49452,N_48854,N_48462);
or U49453 (N_49453,N_48295,N_48598);
and U49454 (N_49454,N_48715,N_48047);
nor U49455 (N_49455,N_48846,N_48896);
and U49456 (N_49456,N_48588,N_48327);
nand U49457 (N_49457,N_48912,N_48479);
and U49458 (N_49458,N_48907,N_48980);
or U49459 (N_49459,N_48040,N_48476);
xor U49460 (N_49460,N_48473,N_48484);
nand U49461 (N_49461,N_48277,N_48029);
nand U49462 (N_49462,N_48467,N_48633);
nor U49463 (N_49463,N_48796,N_48946);
nand U49464 (N_49464,N_48973,N_48621);
or U49465 (N_49465,N_48336,N_48101);
nand U49466 (N_49466,N_48252,N_48893);
nand U49467 (N_49467,N_48714,N_48545);
nor U49468 (N_49468,N_48038,N_48730);
nand U49469 (N_49469,N_48667,N_48324);
nor U49470 (N_49470,N_48446,N_48566);
or U49471 (N_49471,N_48762,N_48965);
nor U49472 (N_49472,N_48821,N_48605);
nor U49473 (N_49473,N_48929,N_48400);
nor U49474 (N_49474,N_48663,N_48174);
nand U49475 (N_49475,N_48100,N_48495);
xnor U49476 (N_49476,N_48314,N_48784);
nor U49477 (N_49477,N_48298,N_48068);
or U49478 (N_49478,N_48885,N_48882);
xnor U49479 (N_49479,N_48351,N_48665);
nand U49480 (N_49480,N_48220,N_48344);
and U49481 (N_49481,N_48871,N_48075);
xor U49482 (N_49482,N_48465,N_48305);
nor U49483 (N_49483,N_48660,N_48904);
or U49484 (N_49484,N_48918,N_48718);
or U49485 (N_49485,N_48222,N_48003);
and U49486 (N_49486,N_48543,N_48379);
xnor U49487 (N_49487,N_48266,N_48867);
or U49488 (N_49488,N_48335,N_48691);
and U49489 (N_49489,N_48866,N_48541);
xor U49490 (N_49490,N_48947,N_48141);
or U49491 (N_49491,N_48806,N_48770);
nand U49492 (N_49492,N_48372,N_48094);
and U49493 (N_49493,N_48966,N_48939);
nor U49494 (N_49494,N_48218,N_48892);
xnor U49495 (N_49495,N_48768,N_48646);
nand U49496 (N_49496,N_48601,N_48790);
nand U49497 (N_49497,N_48054,N_48931);
or U49498 (N_49498,N_48320,N_48782);
xnor U49499 (N_49499,N_48987,N_48257);
xor U49500 (N_49500,N_48863,N_48454);
nand U49501 (N_49501,N_48854,N_48454);
nand U49502 (N_49502,N_48834,N_48283);
xor U49503 (N_49503,N_48725,N_48516);
nand U49504 (N_49504,N_48135,N_48590);
and U49505 (N_49505,N_48706,N_48959);
xor U49506 (N_49506,N_48048,N_48483);
nand U49507 (N_49507,N_48475,N_48266);
xor U49508 (N_49508,N_48177,N_48127);
xnor U49509 (N_49509,N_48860,N_48347);
or U49510 (N_49510,N_48616,N_48264);
or U49511 (N_49511,N_48390,N_48891);
or U49512 (N_49512,N_48415,N_48709);
nor U49513 (N_49513,N_48846,N_48378);
or U49514 (N_49514,N_48638,N_48062);
or U49515 (N_49515,N_48326,N_48758);
xnor U49516 (N_49516,N_48575,N_48524);
or U49517 (N_49517,N_48734,N_48934);
nand U49518 (N_49518,N_48547,N_48518);
xnor U49519 (N_49519,N_48241,N_48322);
or U49520 (N_49520,N_48194,N_48001);
xor U49521 (N_49521,N_48437,N_48312);
and U49522 (N_49522,N_48181,N_48652);
nand U49523 (N_49523,N_48634,N_48033);
nand U49524 (N_49524,N_48786,N_48114);
nor U49525 (N_49525,N_48841,N_48755);
or U49526 (N_49526,N_48754,N_48950);
nand U49527 (N_49527,N_48116,N_48918);
xor U49528 (N_49528,N_48531,N_48291);
or U49529 (N_49529,N_48161,N_48192);
or U49530 (N_49530,N_48198,N_48783);
nor U49531 (N_49531,N_48410,N_48646);
nand U49532 (N_49532,N_48046,N_48604);
xor U49533 (N_49533,N_48811,N_48629);
xor U49534 (N_49534,N_48831,N_48361);
xnor U49535 (N_49535,N_48762,N_48331);
nand U49536 (N_49536,N_48200,N_48363);
and U49537 (N_49537,N_48759,N_48002);
and U49538 (N_49538,N_48590,N_48205);
and U49539 (N_49539,N_48866,N_48922);
and U49540 (N_49540,N_48512,N_48877);
nor U49541 (N_49541,N_48878,N_48050);
nand U49542 (N_49542,N_48735,N_48079);
and U49543 (N_49543,N_48917,N_48468);
nand U49544 (N_49544,N_48631,N_48957);
or U49545 (N_49545,N_48339,N_48746);
or U49546 (N_49546,N_48572,N_48707);
or U49547 (N_49547,N_48956,N_48844);
xor U49548 (N_49548,N_48819,N_48453);
or U49549 (N_49549,N_48732,N_48837);
nand U49550 (N_49550,N_48665,N_48321);
xnor U49551 (N_49551,N_48806,N_48445);
nor U49552 (N_49552,N_48181,N_48776);
xnor U49553 (N_49553,N_48354,N_48815);
nor U49554 (N_49554,N_48687,N_48417);
nand U49555 (N_49555,N_48115,N_48863);
nand U49556 (N_49556,N_48737,N_48547);
xor U49557 (N_49557,N_48713,N_48649);
nand U49558 (N_49558,N_48799,N_48735);
or U49559 (N_49559,N_48644,N_48606);
nand U49560 (N_49560,N_48338,N_48782);
xnor U49561 (N_49561,N_48457,N_48729);
nand U49562 (N_49562,N_48804,N_48409);
and U49563 (N_49563,N_48422,N_48628);
or U49564 (N_49564,N_48374,N_48801);
xnor U49565 (N_49565,N_48029,N_48235);
and U49566 (N_49566,N_48205,N_48698);
or U49567 (N_49567,N_48705,N_48254);
nor U49568 (N_49568,N_48882,N_48368);
nor U49569 (N_49569,N_48552,N_48348);
and U49570 (N_49570,N_48703,N_48556);
nor U49571 (N_49571,N_48645,N_48968);
or U49572 (N_49572,N_48815,N_48168);
xnor U49573 (N_49573,N_48442,N_48679);
and U49574 (N_49574,N_48076,N_48359);
xnor U49575 (N_49575,N_48637,N_48798);
nand U49576 (N_49576,N_48247,N_48134);
nand U49577 (N_49577,N_48048,N_48394);
nand U49578 (N_49578,N_48576,N_48256);
nand U49579 (N_49579,N_48877,N_48702);
nor U49580 (N_49580,N_48610,N_48080);
nand U49581 (N_49581,N_48755,N_48449);
nor U49582 (N_49582,N_48317,N_48168);
nand U49583 (N_49583,N_48448,N_48037);
nor U49584 (N_49584,N_48292,N_48505);
nor U49585 (N_49585,N_48314,N_48220);
xnor U49586 (N_49586,N_48107,N_48550);
xnor U49587 (N_49587,N_48980,N_48357);
or U49588 (N_49588,N_48511,N_48304);
xor U49589 (N_49589,N_48500,N_48281);
xor U49590 (N_49590,N_48575,N_48778);
xor U49591 (N_49591,N_48492,N_48279);
nor U49592 (N_49592,N_48186,N_48065);
or U49593 (N_49593,N_48556,N_48773);
nand U49594 (N_49594,N_48388,N_48977);
nand U49595 (N_49595,N_48645,N_48695);
xor U49596 (N_49596,N_48764,N_48903);
nor U49597 (N_49597,N_48398,N_48315);
and U49598 (N_49598,N_48082,N_48122);
and U49599 (N_49599,N_48449,N_48453);
nor U49600 (N_49600,N_48313,N_48274);
nor U49601 (N_49601,N_48569,N_48821);
xor U49602 (N_49602,N_48104,N_48441);
and U49603 (N_49603,N_48319,N_48174);
and U49604 (N_49604,N_48060,N_48420);
xnor U49605 (N_49605,N_48743,N_48755);
nand U49606 (N_49606,N_48463,N_48265);
and U49607 (N_49607,N_48275,N_48649);
xor U49608 (N_49608,N_48227,N_48467);
nand U49609 (N_49609,N_48475,N_48409);
xnor U49610 (N_49610,N_48521,N_48204);
nand U49611 (N_49611,N_48949,N_48475);
xor U49612 (N_49612,N_48109,N_48618);
or U49613 (N_49613,N_48428,N_48798);
nand U49614 (N_49614,N_48416,N_48402);
nand U49615 (N_49615,N_48987,N_48067);
or U49616 (N_49616,N_48481,N_48625);
nand U49617 (N_49617,N_48613,N_48621);
nand U49618 (N_49618,N_48599,N_48021);
and U49619 (N_49619,N_48093,N_48679);
and U49620 (N_49620,N_48612,N_48818);
or U49621 (N_49621,N_48744,N_48574);
nor U49622 (N_49622,N_48701,N_48149);
nor U49623 (N_49623,N_48066,N_48713);
or U49624 (N_49624,N_48897,N_48771);
nand U49625 (N_49625,N_48784,N_48454);
nand U49626 (N_49626,N_48778,N_48843);
and U49627 (N_49627,N_48018,N_48108);
xor U49628 (N_49628,N_48779,N_48147);
nor U49629 (N_49629,N_48908,N_48756);
xor U49630 (N_49630,N_48166,N_48790);
xor U49631 (N_49631,N_48716,N_48899);
nor U49632 (N_49632,N_48152,N_48371);
nor U49633 (N_49633,N_48462,N_48289);
nand U49634 (N_49634,N_48512,N_48030);
nor U49635 (N_49635,N_48480,N_48279);
nand U49636 (N_49636,N_48987,N_48461);
or U49637 (N_49637,N_48016,N_48160);
and U49638 (N_49638,N_48872,N_48169);
or U49639 (N_49639,N_48003,N_48846);
or U49640 (N_49640,N_48333,N_48979);
nand U49641 (N_49641,N_48808,N_48718);
xor U49642 (N_49642,N_48600,N_48169);
or U49643 (N_49643,N_48202,N_48821);
xor U49644 (N_49644,N_48672,N_48937);
xor U49645 (N_49645,N_48494,N_48268);
nand U49646 (N_49646,N_48050,N_48423);
nand U49647 (N_49647,N_48566,N_48215);
xnor U49648 (N_49648,N_48000,N_48037);
nand U49649 (N_49649,N_48602,N_48088);
xnor U49650 (N_49650,N_48917,N_48387);
xnor U49651 (N_49651,N_48321,N_48179);
xnor U49652 (N_49652,N_48416,N_48107);
nand U49653 (N_49653,N_48106,N_48396);
or U49654 (N_49654,N_48656,N_48451);
or U49655 (N_49655,N_48259,N_48562);
nand U49656 (N_49656,N_48333,N_48776);
and U49657 (N_49657,N_48737,N_48589);
xor U49658 (N_49658,N_48894,N_48402);
nor U49659 (N_49659,N_48361,N_48964);
nand U49660 (N_49660,N_48982,N_48051);
xor U49661 (N_49661,N_48099,N_48059);
and U49662 (N_49662,N_48832,N_48770);
xor U49663 (N_49663,N_48107,N_48658);
and U49664 (N_49664,N_48023,N_48375);
nand U49665 (N_49665,N_48318,N_48420);
xnor U49666 (N_49666,N_48585,N_48146);
xor U49667 (N_49667,N_48868,N_48641);
xor U49668 (N_49668,N_48971,N_48104);
xnor U49669 (N_49669,N_48768,N_48016);
nand U49670 (N_49670,N_48670,N_48198);
and U49671 (N_49671,N_48933,N_48356);
nor U49672 (N_49672,N_48507,N_48427);
nor U49673 (N_49673,N_48309,N_48969);
xnor U49674 (N_49674,N_48441,N_48579);
nand U49675 (N_49675,N_48468,N_48119);
nor U49676 (N_49676,N_48145,N_48964);
xnor U49677 (N_49677,N_48061,N_48408);
nand U49678 (N_49678,N_48335,N_48032);
xnor U49679 (N_49679,N_48646,N_48487);
or U49680 (N_49680,N_48395,N_48954);
or U49681 (N_49681,N_48208,N_48764);
nor U49682 (N_49682,N_48873,N_48189);
nand U49683 (N_49683,N_48475,N_48017);
or U49684 (N_49684,N_48723,N_48530);
xor U49685 (N_49685,N_48092,N_48137);
or U49686 (N_49686,N_48005,N_48662);
nor U49687 (N_49687,N_48180,N_48761);
nand U49688 (N_49688,N_48222,N_48164);
and U49689 (N_49689,N_48361,N_48740);
or U49690 (N_49690,N_48187,N_48558);
and U49691 (N_49691,N_48508,N_48932);
or U49692 (N_49692,N_48659,N_48151);
and U49693 (N_49693,N_48374,N_48757);
nand U49694 (N_49694,N_48940,N_48488);
and U49695 (N_49695,N_48755,N_48709);
and U49696 (N_49696,N_48596,N_48592);
nor U49697 (N_49697,N_48875,N_48719);
xor U49698 (N_49698,N_48184,N_48681);
nand U49699 (N_49699,N_48860,N_48548);
nor U49700 (N_49700,N_48050,N_48864);
nand U49701 (N_49701,N_48378,N_48150);
nand U49702 (N_49702,N_48777,N_48131);
or U49703 (N_49703,N_48387,N_48540);
nor U49704 (N_49704,N_48646,N_48389);
and U49705 (N_49705,N_48376,N_48418);
nand U49706 (N_49706,N_48518,N_48673);
and U49707 (N_49707,N_48628,N_48615);
nand U49708 (N_49708,N_48991,N_48886);
or U49709 (N_49709,N_48195,N_48978);
nand U49710 (N_49710,N_48745,N_48836);
nand U49711 (N_49711,N_48954,N_48603);
nand U49712 (N_49712,N_48492,N_48381);
nand U49713 (N_49713,N_48955,N_48779);
xor U49714 (N_49714,N_48686,N_48598);
or U49715 (N_49715,N_48470,N_48739);
nand U49716 (N_49716,N_48747,N_48231);
or U49717 (N_49717,N_48529,N_48395);
nor U49718 (N_49718,N_48088,N_48631);
nand U49719 (N_49719,N_48991,N_48647);
xnor U49720 (N_49720,N_48078,N_48927);
or U49721 (N_49721,N_48647,N_48277);
nand U49722 (N_49722,N_48607,N_48007);
nand U49723 (N_49723,N_48573,N_48777);
nand U49724 (N_49724,N_48057,N_48019);
nand U49725 (N_49725,N_48963,N_48454);
and U49726 (N_49726,N_48887,N_48617);
nor U49727 (N_49727,N_48162,N_48103);
nand U49728 (N_49728,N_48866,N_48247);
and U49729 (N_49729,N_48688,N_48490);
or U49730 (N_49730,N_48259,N_48353);
or U49731 (N_49731,N_48593,N_48308);
nor U49732 (N_49732,N_48794,N_48738);
nor U49733 (N_49733,N_48352,N_48142);
or U49734 (N_49734,N_48830,N_48351);
xor U49735 (N_49735,N_48194,N_48739);
or U49736 (N_49736,N_48180,N_48880);
nor U49737 (N_49737,N_48852,N_48500);
nor U49738 (N_49738,N_48513,N_48374);
nor U49739 (N_49739,N_48782,N_48471);
or U49740 (N_49740,N_48017,N_48131);
nor U49741 (N_49741,N_48962,N_48603);
and U49742 (N_49742,N_48800,N_48356);
or U49743 (N_49743,N_48125,N_48572);
xnor U49744 (N_49744,N_48151,N_48710);
and U49745 (N_49745,N_48783,N_48832);
xnor U49746 (N_49746,N_48533,N_48308);
nor U49747 (N_49747,N_48297,N_48505);
and U49748 (N_49748,N_48690,N_48442);
or U49749 (N_49749,N_48669,N_48526);
and U49750 (N_49750,N_48981,N_48759);
or U49751 (N_49751,N_48919,N_48571);
nor U49752 (N_49752,N_48017,N_48672);
nor U49753 (N_49753,N_48460,N_48601);
and U49754 (N_49754,N_48410,N_48061);
or U49755 (N_49755,N_48130,N_48808);
nand U49756 (N_49756,N_48166,N_48003);
nand U49757 (N_49757,N_48184,N_48382);
or U49758 (N_49758,N_48726,N_48672);
nor U49759 (N_49759,N_48179,N_48777);
and U49760 (N_49760,N_48101,N_48655);
xnor U49761 (N_49761,N_48795,N_48639);
xor U49762 (N_49762,N_48739,N_48967);
nand U49763 (N_49763,N_48266,N_48529);
nor U49764 (N_49764,N_48835,N_48934);
nand U49765 (N_49765,N_48820,N_48424);
xor U49766 (N_49766,N_48425,N_48051);
xor U49767 (N_49767,N_48708,N_48196);
and U49768 (N_49768,N_48057,N_48071);
nand U49769 (N_49769,N_48687,N_48627);
and U49770 (N_49770,N_48450,N_48867);
nand U49771 (N_49771,N_48766,N_48952);
nor U49772 (N_49772,N_48600,N_48337);
nor U49773 (N_49773,N_48588,N_48448);
nor U49774 (N_49774,N_48807,N_48055);
and U49775 (N_49775,N_48245,N_48747);
and U49776 (N_49776,N_48332,N_48620);
xor U49777 (N_49777,N_48007,N_48618);
and U49778 (N_49778,N_48023,N_48998);
xor U49779 (N_49779,N_48440,N_48809);
and U49780 (N_49780,N_48863,N_48942);
or U49781 (N_49781,N_48113,N_48719);
nor U49782 (N_49782,N_48629,N_48322);
nand U49783 (N_49783,N_48052,N_48433);
nand U49784 (N_49784,N_48530,N_48330);
and U49785 (N_49785,N_48389,N_48310);
xor U49786 (N_49786,N_48312,N_48346);
nor U49787 (N_49787,N_48596,N_48988);
or U49788 (N_49788,N_48483,N_48711);
and U49789 (N_49789,N_48416,N_48163);
nand U49790 (N_49790,N_48647,N_48975);
nor U49791 (N_49791,N_48413,N_48103);
nand U49792 (N_49792,N_48833,N_48082);
or U49793 (N_49793,N_48486,N_48635);
xor U49794 (N_49794,N_48054,N_48179);
xor U49795 (N_49795,N_48716,N_48458);
nor U49796 (N_49796,N_48059,N_48768);
nand U49797 (N_49797,N_48432,N_48198);
or U49798 (N_49798,N_48374,N_48161);
nor U49799 (N_49799,N_48217,N_48864);
nor U49800 (N_49800,N_48041,N_48096);
and U49801 (N_49801,N_48943,N_48781);
xor U49802 (N_49802,N_48399,N_48061);
xnor U49803 (N_49803,N_48325,N_48277);
and U49804 (N_49804,N_48427,N_48125);
xnor U49805 (N_49805,N_48870,N_48660);
xnor U49806 (N_49806,N_48373,N_48206);
or U49807 (N_49807,N_48126,N_48741);
nand U49808 (N_49808,N_48445,N_48102);
or U49809 (N_49809,N_48604,N_48881);
nor U49810 (N_49810,N_48487,N_48819);
xor U49811 (N_49811,N_48235,N_48485);
nand U49812 (N_49812,N_48959,N_48504);
nor U49813 (N_49813,N_48680,N_48779);
xor U49814 (N_49814,N_48995,N_48304);
or U49815 (N_49815,N_48863,N_48243);
nor U49816 (N_49816,N_48763,N_48971);
xnor U49817 (N_49817,N_48972,N_48991);
nor U49818 (N_49818,N_48627,N_48626);
or U49819 (N_49819,N_48251,N_48616);
nand U49820 (N_49820,N_48167,N_48661);
or U49821 (N_49821,N_48590,N_48551);
nand U49822 (N_49822,N_48870,N_48836);
nor U49823 (N_49823,N_48286,N_48728);
or U49824 (N_49824,N_48504,N_48194);
or U49825 (N_49825,N_48803,N_48517);
or U49826 (N_49826,N_48841,N_48109);
xnor U49827 (N_49827,N_48769,N_48456);
and U49828 (N_49828,N_48335,N_48152);
nand U49829 (N_49829,N_48519,N_48140);
or U49830 (N_49830,N_48637,N_48542);
nand U49831 (N_49831,N_48111,N_48607);
and U49832 (N_49832,N_48030,N_48297);
nor U49833 (N_49833,N_48421,N_48541);
xnor U49834 (N_49834,N_48459,N_48530);
and U49835 (N_49835,N_48057,N_48689);
nor U49836 (N_49836,N_48696,N_48382);
nor U49837 (N_49837,N_48000,N_48440);
xnor U49838 (N_49838,N_48315,N_48027);
nand U49839 (N_49839,N_48720,N_48829);
or U49840 (N_49840,N_48559,N_48007);
or U49841 (N_49841,N_48488,N_48599);
xor U49842 (N_49842,N_48550,N_48471);
or U49843 (N_49843,N_48112,N_48292);
nand U49844 (N_49844,N_48284,N_48633);
or U49845 (N_49845,N_48890,N_48455);
or U49846 (N_49846,N_48645,N_48680);
xor U49847 (N_49847,N_48480,N_48273);
and U49848 (N_49848,N_48861,N_48768);
or U49849 (N_49849,N_48766,N_48217);
and U49850 (N_49850,N_48251,N_48246);
nand U49851 (N_49851,N_48527,N_48296);
and U49852 (N_49852,N_48053,N_48171);
or U49853 (N_49853,N_48354,N_48953);
nor U49854 (N_49854,N_48501,N_48700);
xor U49855 (N_49855,N_48279,N_48339);
nor U49856 (N_49856,N_48384,N_48021);
and U49857 (N_49857,N_48387,N_48221);
nor U49858 (N_49858,N_48915,N_48921);
and U49859 (N_49859,N_48970,N_48687);
and U49860 (N_49860,N_48958,N_48776);
nand U49861 (N_49861,N_48594,N_48089);
xor U49862 (N_49862,N_48200,N_48631);
and U49863 (N_49863,N_48322,N_48656);
and U49864 (N_49864,N_48848,N_48453);
or U49865 (N_49865,N_48256,N_48746);
xnor U49866 (N_49866,N_48333,N_48731);
or U49867 (N_49867,N_48774,N_48714);
nand U49868 (N_49868,N_48995,N_48400);
xnor U49869 (N_49869,N_48244,N_48826);
nor U49870 (N_49870,N_48801,N_48054);
nand U49871 (N_49871,N_48954,N_48353);
nor U49872 (N_49872,N_48550,N_48830);
or U49873 (N_49873,N_48087,N_48767);
nand U49874 (N_49874,N_48210,N_48516);
xor U49875 (N_49875,N_48787,N_48840);
nor U49876 (N_49876,N_48228,N_48492);
nor U49877 (N_49877,N_48095,N_48028);
nor U49878 (N_49878,N_48532,N_48147);
xnor U49879 (N_49879,N_48686,N_48559);
or U49880 (N_49880,N_48596,N_48223);
nor U49881 (N_49881,N_48585,N_48704);
xnor U49882 (N_49882,N_48021,N_48964);
xor U49883 (N_49883,N_48658,N_48610);
or U49884 (N_49884,N_48443,N_48786);
or U49885 (N_49885,N_48479,N_48568);
or U49886 (N_49886,N_48085,N_48615);
xnor U49887 (N_49887,N_48342,N_48120);
nand U49888 (N_49888,N_48047,N_48089);
nor U49889 (N_49889,N_48310,N_48063);
and U49890 (N_49890,N_48896,N_48898);
nor U49891 (N_49891,N_48168,N_48452);
xor U49892 (N_49892,N_48819,N_48695);
or U49893 (N_49893,N_48568,N_48264);
nor U49894 (N_49894,N_48049,N_48112);
or U49895 (N_49895,N_48658,N_48969);
and U49896 (N_49896,N_48739,N_48119);
nand U49897 (N_49897,N_48757,N_48067);
xor U49898 (N_49898,N_48899,N_48307);
nor U49899 (N_49899,N_48195,N_48516);
nor U49900 (N_49900,N_48561,N_48508);
nor U49901 (N_49901,N_48337,N_48081);
nand U49902 (N_49902,N_48481,N_48327);
or U49903 (N_49903,N_48414,N_48816);
nand U49904 (N_49904,N_48883,N_48369);
nand U49905 (N_49905,N_48725,N_48497);
and U49906 (N_49906,N_48379,N_48984);
nand U49907 (N_49907,N_48728,N_48339);
nand U49908 (N_49908,N_48193,N_48216);
xor U49909 (N_49909,N_48453,N_48560);
or U49910 (N_49910,N_48463,N_48484);
xnor U49911 (N_49911,N_48321,N_48404);
xor U49912 (N_49912,N_48910,N_48757);
or U49913 (N_49913,N_48054,N_48024);
or U49914 (N_49914,N_48530,N_48754);
and U49915 (N_49915,N_48411,N_48703);
xor U49916 (N_49916,N_48356,N_48473);
nand U49917 (N_49917,N_48828,N_48036);
xnor U49918 (N_49918,N_48016,N_48796);
xnor U49919 (N_49919,N_48261,N_48152);
nor U49920 (N_49920,N_48376,N_48094);
xor U49921 (N_49921,N_48322,N_48580);
nand U49922 (N_49922,N_48797,N_48664);
xor U49923 (N_49923,N_48863,N_48457);
nor U49924 (N_49924,N_48284,N_48549);
nor U49925 (N_49925,N_48681,N_48585);
and U49926 (N_49926,N_48981,N_48615);
and U49927 (N_49927,N_48875,N_48743);
or U49928 (N_49928,N_48572,N_48320);
nand U49929 (N_49929,N_48201,N_48553);
xnor U49930 (N_49930,N_48990,N_48248);
xnor U49931 (N_49931,N_48510,N_48024);
xor U49932 (N_49932,N_48271,N_48413);
nor U49933 (N_49933,N_48746,N_48950);
xor U49934 (N_49934,N_48878,N_48629);
and U49935 (N_49935,N_48850,N_48354);
nand U49936 (N_49936,N_48153,N_48902);
and U49937 (N_49937,N_48112,N_48216);
or U49938 (N_49938,N_48810,N_48740);
nor U49939 (N_49939,N_48863,N_48313);
xor U49940 (N_49940,N_48944,N_48872);
and U49941 (N_49941,N_48741,N_48124);
nand U49942 (N_49942,N_48288,N_48240);
or U49943 (N_49943,N_48762,N_48599);
xor U49944 (N_49944,N_48222,N_48779);
nor U49945 (N_49945,N_48440,N_48711);
and U49946 (N_49946,N_48868,N_48483);
and U49947 (N_49947,N_48291,N_48901);
nand U49948 (N_49948,N_48244,N_48619);
xnor U49949 (N_49949,N_48256,N_48533);
nor U49950 (N_49950,N_48507,N_48927);
nand U49951 (N_49951,N_48157,N_48347);
or U49952 (N_49952,N_48335,N_48395);
and U49953 (N_49953,N_48685,N_48297);
nor U49954 (N_49954,N_48749,N_48901);
xnor U49955 (N_49955,N_48901,N_48578);
xor U49956 (N_49956,N_48431,N_48814);
and U49957 (N_49957,N_48711,N_48522);
nand U49958 (N_49958,N_48241,N_48960);
nor U49959 (N_49959,N_48260,N_48143);
xnor U49960 (N_49960,N_48489,N_48837);
or U49961 (N_49961,N_48335,N_48024);
or U49962 (N_49962,N_48230,N_48168);
or U49963 (N_49963,N_48880,N_48531);
nand U49964 (N_49964,N_48501,N_48783);
and U49965 (N_49965,N_48394,N_48943);
xor U49966 (N_49966,N_48698,N_48217);
or U49967 (N_49967,N_48538,N_48147);
or U49968 (N_49968,N_48247,N_48343);
and U49969 (N_49969,N_48457,N_48546);
or U49970 (N_49970,N_48088,N_48194);
and U49971 (N_49971,N_48826,N_48883);
nor U49972 (N_49972,N_48951,N_48281);
xnor U49973 (N_49973,N_48042,N_48111);
and U49974 (N_49974,N_48315,N_48481);
xor U49975 (N_49975,N_48224,N_48960);
nand U49976 (N_49976,N_48705,N_48900);
or U49977 (N_49977,N_48503,N_48493);
and U49978 (N_49978,N_48806,N_48815);
and U49979 (N_49979,N_48307,N_48138);
nand U49980 (N_49980,N_48966,N_48786);
or U49981 (N_49981,N_48516,N_48878);
nor U49982 (N_49982,N_48482,N_48627);
nand U49983 (N_49983,N_48823,N_48563);
nand U49984 (N_49984,N_48356,N_48772);
xor U49985 (N_49985,N_48929,N_48726);
and U49986 (N_49986,N_48482,N_48336);
nor U49987 (N_49987,N_48121,N_48394);
xor U49988 (N_49988,N_48506,N_48573);
nor U49989 (N_49989,N_48177,N_48103);
or U49990 (N_49990,N_48008,N_48832);
xnor U49991 (N_49991,N_48003,N_48604);
and U49992 (N_49992,N_48835,N_48100);
and U49993 (N_49993,N_48326,N_48515);
and U49994 (N_49994,N_48243,N_48214);
and U49995 (N_49995,N_48463,N_48991);
or U49996 (N_49996,N_48148,N_48215);
or U49997 (N_49997,N_48046,N_48083);
and U49998 (N_49998,N_48065,N_48264);
nand U49999 (N_49999,N_48292,N_48141);
and UO_0 (O_0,N_49790,N_49274);
or UO_1 (O_1,N_49179,N_49898);
or UO_2 (O_2,N_49391,N_49389);
nand UO_3 (O_3,N_49710,N_49417);
nand UO_4 (O_4,N_49143,N_49090);
nor UO_5 (O_5,N_49257,N_49494);
nand UO_6 (O_6,N_49893,N_49138);
and UO_7 (O_7,N_49980,N_49131);
nand UO_8 (O_8,N_49248,N_49992);
or UO_9 (O_9,N_49217,N_49250);
nor UO_10 (O_10,N_49962,N_49644);
or UO_11 (O_11,N_49024,N_49434);
nor UO_12 (O_12,N_49146,N_49570);
nand UO_13 (O_13,N_49709,N_49142);
and UO_14 (O_14,N_49552,N_49587);
or UO_15 (O_15,N_49205,N_49484);
xor UO_16 (O_16,N_49188,N_49464);
or UO_17 (O_17,N_49707,N_49376);
and UO_18 (O_18,N_49934,N_49214);
or UO_19 (O_19,N_49503,N_49746);
nand UO_20 (O_20,N_49974,N_49492);
xor UO_21 (O_21,N_49774,N_49816);
nor UO_22 (O_22,N_49115,N_49286);
or UO_23 (O_23,N_49043,N_49581);
or UO_24 (O_24,N_49760,N_49148);
nor UO_25 (O_25,N_49845,N_49254);
or UO_26 (O_26,N_49378,N_49442);
or UO_27 (O_27,N_49030,N_49575);
and UO_28 (O_28,N_49813,N_49914);
or UO_29 (O_29,N_49358,N_49667);
nor UO_30 (O_30,N_49907,N_49824);
nand UO_31 (O_31,N_49366,N_49008);
nor UO_32 (O_32,N_49216,N_49732);
nand UO_33 (O_33,N_49921,N_49226);
nand UO_34 (O_34,N_49461,N_49384);
or UO_35 (O_35,N_49505,N_49791);
xor UO_36 (O_36,N_49363,N_49512);
or UO_37 (O_37,N_49322,N_49764);
xnor UO_38 (O_38,N_49556,N_49046);
or UO_39 (O_39,N_49308,N_49802);
nor UO_40 (O_40,N_49261,N_49475);
xnor UO_41 (O_41,N_49441,N_49811);
and UO_42 (O_42,N_49691,N_49862);
nand UO_43 (O_43,N_49999,N_49271);
or UO_44 (O_44,N_49749,N_49809);
nor UO_45 (O_45,N_49496,N_49177);
nor UO_46 (O_46,N_49868,N_49565);
nor UO_47 (O_47,N_49941,N_49814);
xnor UO_48 (O_48,N_49601,N_49643);
xnor UO_49 (O_49,N_49078,N_49620);
or UO_50 (O_50,N_49989,N_49653);
nand UO_51 (O_51,N_49616,N_49443);
nand UO_52 (O_52,N_49285,N_49852);
xor UO_53 (O_53,N_49237,N_49338);
or UO_54 (O_54,N_49310,N_49804);
nor UO_55 (O_55,N_49471,N_49950);
nand UO_56 (O_56,N_49943,N_49435);
and UO_57 (O_57,N_49121,N_49932);
or UO_58 (O_58,N_49299,N_49798);
nand UO_59 (O_59,N_49208,N_49438);
xnor UO_60 (O_60,N_49354,N_49977);
nor UO_61 (O_61,N_49718,N_49042);
or UO_62 (O_62,N_49678,N_49806);
nor UO_63 (O_63,N_49132,N_49053);
nand UO_64 (O_64,N_49327,N_49113);
or UO_65 (O_65,N_49976,N_49087);
or UO_66 (O_66,N_49083,N_49129);
nor UO_67 (O_67,N_49057,N_49031);
and UO_68 (O_68,N_49243,N_49199);
xor UO_69 (O_69,N_49164,N_49733);
or UO_70 (O_70,N_49096,N_49022);
nand UO_71 (O_71,N_49750,N_49149);
or UO_72 (O_72,N_49101,N_49987);
or UO_73 (O_73,N_49882,N_49972);
and UO_74 (O_74,N_49588,N_49696);
nor UO_75 (O_75,N_49652,N_49045);
xnor UO_76 (O_76,N_49770,N_49965);
or UO_77 (O_77,N_49896,N_49831);
nor UO_78 (O_78,N_49986,N_49162);
and UO_79 (O_79,N_49547,N_49719);
nand UO_80 (O_80,N_49597,N_49544);
or UO_81 (O_81,N_49320,N_49541);
and UO_82 (O_82,N_49383,N_49298);
nand UO_83 (O_83,N_49326,N_49283);
or UO_84 (O_84,N_49223,N_49751);
nor UO_85 (O_85,N_49721,N_49938);
nor UO_86 (O_86,N_49036,N_49903);
nor UO_87 (O_87,N_49676,N_49268);
nand UO_88 (O_88,N_49398,N_49228);
and UO_89 (O_89,N_49571,N_49742);
nor UO_90 (O_90,N_49507,N_49170);
nand UO_91 (O_91,N_49230,N_49841);
xnor UO_92 (O_92,N_49004,N_49215);
or UO_93 (O_93,N_49945,N_49404);
nand UO_94 (O_94,N_49161,N_49483);
nand UO_95 (O_95,N_49100,N_49933);
or UO_96 (O_96,N_49917,N_49669);
xor UO_97 (O_97,N_49604,N_49970);
or UO_98 (O_98,N_49879,N_49263);
and UO_99 (O_99,N_49075,N_49624);
or UO_100 (O_100,N_49850,N_49614);
and UO_101 (O_101,N_49960,N_49954);
nor UO_102 (O_102,N_49682,N_49655);
xor UO_103 (O_103,N_49531,N_49516);
or UO_104 (O_104,N_49866,N_49032);
or UO_105 (O_105,N_49886,N_49446);
and UO_106 (O_106,N_49532,N_49679);
nor UO_107 (O_107,N_49108,N_49387);
nor UO_108 (O_108,N_49489,N_49830);
nor UO_109 (O_109,N_49399,N_49756);
or UO_110 (O_110,N_49787,N_49041);
nor UO_111 (O_111,N_49474,N_49018);
or UO_112 (O_112,N_49955,N_49777);
or UO_113 (O_113,N_49797,N_49175);
xor UO_114 (O_114,N_49325,N_49603);
and UO_115 (O_115,N_49003,N_49858);
and UO_116 (O_116,N_49346,N_49002);
or UO_117 (O_117,N_49488,N_49712);
nor UO_118 (O_118,N_49069,N_49685);
and UO_119 (O_119,N_49379,N_49273);
nand UO_120 (O_120,N_49854,N_49540);
nor UO_121 (O_121,N_49135,N_49740);
nor UO_122 (O_122,N_49688,N_49559);
and UO_123 (O_123,N_49582,N_49887);
or UO_124 (O_124,N_49224,N_49159);
and UO_125 (O_125,N_49528,N_49805);
xnor UO_126 (O_126,N_49680,N_49996);
xnor UO_127 (O_127,N_49715,N_49585);
nand UO_128 (O_128,N_49744,N_49572);
nor UO_129 (O_129,N_49517,N_49659);
and UO_130 (O_130,N_49234,N_49073);
nor UO_131 (O_131,N_49463,N_49419);
nand UO_132 (O_132,N_49009,N_49686);
or UO_133 (O_133,N_49763,N_49807);
nand UO_134 (O_134,N_49984,N_49748);
xnor UO_135 (O_135,N_49364,N_49859);
xnor UO_136 (O_136,N_49197,N_49029);
nor UO_137 (O_137,N_49178,N_49481);
or UO_138 (O_138,N_49819,N_49079);
and UO_139 (O_139,N_49842,N_49510);
and UO_140 (O_140,N_49506,N_49448);
nor UO_141 (O_141,N_49044,N_49875);
xnor UO_142 (O_142,N_49453,N_49826);
xor UO_143 (O_143,N_49698,N_49759);
and UO_144 (O_144,N_49877,N_49640);
nand UO_145 (O_145,N_49281,N_49220);
nor UO_146 (O_146,N_49180,N_49037);
and UO_147 (O_147,N_49277,N_49410);
xor UO_148 (O_148,N_49204,N_49344);
nand UO_149 (O_149,N_49059,N_49232);
and UO_150 (O_150,N_49985,N_49247);
and UO_151 (O_151,N_49625,N_49158);
nand UO_152 (O_152,N_49118,N_49077);
xor UO_153 (O_153,N_49975,N_49521);
xnor UO_154 (O_154,N_49219,N_49181);
nor UO_155 (O_155,N_49818,N_49820);
nor UO_156 (O_156,N_49776,N_49892);
nor UO_157 (O_157,N_49618,N_49752);
nor UO_158 (O_158,N_49602,N_49632);
nand UO_159 (O_159,N_49373,N_49035);
or UO_160 (O_160,N_49315,N_49705);
xnor UO_161 (O_161,N_49757,N_49339);
nand UO_162 (O_162,N_49983,N_49971);
nand UO_163 (O_163,N_49051,N_49104);
nand UO_164 (O_164,N_49596,N_49392);
nor UO_165 (O_165,N_49287,N_49425);
and UO_166 (O_166,N_49949,N_49773);
xnor UO_167 (O_167,N_49335,N_49309);
nand UO_168 (O_168,N_49677,N_49169);
xnor UO_169 (O_169,N_49594,N_49871);
nor UO_170 (O_170,N_49660,N_49076);
nand UO_171 (O_171,N_49401,N_49103);
and UO_172 (O_172,N_49539,N_49846);
xor UO_173 (O_173,N_49658,N_49249);
nand UO_174 (O_174,N_49926,N_49106);
nand UO_175 (O_175,N_49737,N_49393);
nand UO_176 (O_176,N_49167,N_49951);
xnor UO_177 (O_177,N_49490,N_49340);
xor UO_178 (O_178,N_49405,N_49470);
nor UO_179 (O_179,N_49068,N_49125);
and UO_180 (O_180,N_49317,N_49613);
nand UO_181 (O_181,N_49525,N_49551);
nand UO_182 (O_182,N_49988,N_49049);
and UO_183 (O_183,N_49380,N_49110);
nand UO_184 (O_184,N_49671,N_49112);
or UO_185 (O_185,N_49642,N_49687);
nand UO_186 (O_186,N_49120,N_49935);
nor UO_187 (O_187,N_49562,N_49156);
nand UO_188 (O_188,N_49833,N_49005);
xor UO_189 (O_189,N_49873,N_49360);
nor UO_190 (O_190,N_49743,N_49089);
and UO_191 (O_191,N_49174,N_49947);
nand UO_192 (O_192,N_49145,N_49140);
or UO_193 (O_193,N_49421,N_49176);
and UO_194 (O_194,N_49206,N_49825);
and UO_195 (O_195,N_49792,N_49229);
nor UO_196 (O_196,N_49072,N_49981);
and UO_197 (O_197,N_49568,N_49088);
and UO_198 (O_198,N_49674,N_49487);
xnor UO_199 (O_199,N_49429,N_49840);
nand UO_200 (O_200,N_49406,N_49646);
nand UO_201 (O_201,N_49353,N_49351);
xor UO_202 (O_202,N_49692,N_49323);
and UO_203 (O_203,N_49504,N_49593);
xor UO_204 (O_204,N_49134,N_49105);
nor UO_205 (O_205,N_49966,N_49781);
or UO_206 (O_206,N_49063,N_49447);
nor UO_207 (O_207,N_49246,N_49296);
nand UO_208 (O_208,N_49708,N_49221);
xnor UO_209 (O_209,N_49662,N_49400);
and UO_210 (O_210,N_49333,N_49319);
or UO_211 (O_211,N_49194,N_49827);
and UO_212 (O_212,N_49193,N_49675);
nand UO_213 (O_213,N_49227,N_49835);
or UO_214 (O_214,N_49796,N_49650);
or UO_215 (O_215,N_49923,N_49838);
or UO_216 (O_216,N_49297,N_49994);
nand UO_217 (O_217,N_49538,N_49055);
nand UO_218 (O_218,N_49374,N_49012);
or UO_219 (O_219,N_49520,N_49573);
or UO_220 (O_220,N_49280,N_49902);
and UO_221 (O_221,N_49124,N_49092);
nor UO_222 (O_222,N_49225,N_49722);
or UO_223 (O_223,N_49395,N_49067);
nand UO_224 (O_224,N_49166,N_49300);
nor UO_225 (O_225,N_49458,N_49924);
or UO_226 (O_226,N_49386,N_49634);
nor UO_227 (O_227,N_49244,N_49165);
xnor UO_228 (O_228,N_49304,N_49745);
nor UO_229 (O_229,N_49431,N_49245);
xor UO_230 (O_230,N_49302,N_49548);
or UO_231 (O_231,N_49359,N_49959);
and UO_232 (O_232,N_49665,N_49969);
nor UO_233 (O_233,N_49729,N_49497);
and UO_234 (O_234,N_49252,N_49656);
nand UO_235 (O_235,N_49592,N_49785);
or UO_236 (O_236,N_49198,N_49058);
xnor UO_237 (O_237,N_49390,N_49670);
nor UO_238 (O_238,N_49576,N_49313);
xnor UO_239 (O_239,N_49612,N_49714);
or UO_240 (O_240,N_49433,N_49615);
nand UO_241 (O_241,N_49080,N_49352);
nor UO_242 (O_242,N_49127,N_49154);
or UO_243 (O_243,N_49098,N_49953);
or UO_244 (O_244,N_49734,N_49210);
nor UO_245 (O_245,N_49038,N_49948);
and UO_246 (O_246,N_49524,N_49645);
and UO_247 (O_247,N_49253,N_49681);
nand UO_248 (O_248,N_49895,N_49451);
nand UO_249 (O_249,N_49196,N_49855);
nand UO_250 (O_250,N_49266,N_49535);
or UO_251 (O_251,N_49242,N_49288);
or UO_252 (O_252,N_49093,N_49716);
xor UO_253 (O_253,N_49367,N_49881);
nand UO_254 (O_254,N_49514,N_49851);
nor UO_255 (O_255,N_49459,N_49084);
and UO_256 (O_256,N_49622,N_49839);
and UO_257 (O_257,N_49269,N_49815);
nand UO_258 (O_258,N_49466,N_49526);
and UO_259 (O_259,N_49025,N_49119);
xor UO_260 (O_260,N_49258,N_49095);
xor UO_261 (O_261,N_49201,N_49578);
nand UO_262 (O_262,N_49753,N_49284);
xor UO_263 (O_263,N_49728,N_49689);
xnor UO_264 (O_264,N_49810,N_49017);
nor UO_265 (O_265,N_49761,N_49369);
nor UO_266 (O_266,N_49856,N_49889);
nand UO_267 (O_267,N_49307,N_49884);
xor UO_268 (O_268,N_49872,N_49978);
xnor UO_269 (O_269,N_49995,N_49457);
nand UO_270 (O_270,N_49522,N_49537);
or UO_271 (O_271,N_49928,N_49701);
and UO_272 (O_272,N_49991,N_49626);
xor UO_273 (O_273,N_49305,N_49021);
xnor UO_274 (O_274,N_49292,N_49607);
or UO_275 (O_275,N_49717,N_49704);
nor UO_276 (O_276,N_49420,N_49929);
xnor UO_277 (O_277,N_49937,N_49808);
nor UO_278 (O_278,N_49337,N_49589);
and UO_279 (O_279,N_49040,N_49793);
xor UO_280 (O_280,N_49412,N_49783);
and UO_281 (O_281,N_49621,N_49595);
and UO_282 (O_282,N_49086,N_49880);
or UO_283 (O_283,N_49428,N_49385);
or UO_284 (O_284,N_49747,N_49515);
and UO_285 (O_285,N_49894,N_49560);
or UO_286 (O_286,N_49890,N_49111);
nand UO_287 (O_287,N_49906,N_49725);
or UO_288 (O_288,N_49649,N_49766);
xnor UO_289 (O_289,N_49136,N_49543);
and UO_290 (O_290,N_49736,N_49312);
or UO_291 (O_291,N_49182,N_49913);
nor UO_292 (O_292,N_49306,N_49303);
or UO_293 (O_293,N_49486,N_49109);
nor UO_294 (O_294,N_49654,N_49699);
nor UO_295 (O_295,N_49262,N_49979);
and UO_296 (O_296,N_49927,N_49508);
or UO_297 (O_297,N_49065,N_49343);
nand UO_298 (O_298,N_49278,N_49255);
xor UO_299 (O_299,N_49114,N_49657);
nand UO_300 (O_300,N_49795,N_49860);
or UO_301 (O_301,N_49186,N_49758);
xnor UO_302 (O_302,N_49415,N_49545);
nand UO_303 (O_303,N_49735,N_49509);
nor UO_304 (O_304,N_49173,N_49117);
or UO_305 (O_305,N_49282,N_49579);
nor UO_306 (O_306,N_49402,N_49563);
and UO_307 (O_307,N_49861,N_49289);
and UO_308 (O_308,N_49047,N_49240);
nor UO_309 (O_309,N_49048,N_49342);
nand UO_310 (O_310,N_49799,N_49925);
nor UO_311 (O_311,N_49014,N_49207);
or UO_312 (O_312,N_49368,N_49432);
and UO_313 (O_313,N_49910,N_49518);
nor UO_314 (O_314,N_49627,N_49328);
nor UO_315 (O_315,N_49122,N_49445);
nand UO_316 (O_316,N_49967,N_49794);
nor UO_317 (O_317,N_49511,N_49836);
xor UO_318 (O_318,N_49946,N_49424);
and UO_319 (O_319,N_49430,N_49301);
and UO_320 (O_320,N_49534,N_49097);
or UO_321 (O_321,N_49423,N_49473);
nor UO_322 (O_322,N_49452,N_49469);
and UO_323 (O_323,N_49973,N_49332);
or UO_324 (O_324,N_49911,N_49623);
or UO_325 (O_325,N_49553,N_49265);
or UO_326 (O_326,N_49062,N_49739);
nand UO_327 (O_327,N_49519,N_49638);
nand UO_328 (O_328,N_49754,N_49316);
nor UO_329 (O_329,N_49741,N_49381);
nor UO_330 (O_330,N_49187,N_49370);
nand UO_331 (O_331,N_49418,N_49817);
nand UO_332 (O_332,N_49812,N_49844);
or UO_333 (O_333,N_49026,N_49144);
nor UO_334 (O_334,N_49591,N_49775);
nor UO_335 (O_335,N_49664,N_49347);
nand UO_336 (O_336,N_49546,N_49956);
or UO_337 (O_337,N_49211,N_49784);
nor UO_338 (O_338,N_49372,N_49908);
nand UO_339 (O_339,N_49139,N_49130);
or UO_340 (O_340,N_49542,N_49336);
nand UO_341 (O_341,N_49789,N_49082);
and UO_342 (O_342,N_49414,N_49891);
or UO_343 (O_343,N_49648,N_49788);
nand UO_344 (O_344,N_49183,N_49467);
or UO_345 (O_345,N_49918,N_49061);
or UO_346 (O_346,N_49912,N_49800);
nor UO_347 (O_347,N_49500,N_49081);
nor UO_348 (O_348,N_49867,N_49480);
nor UO_349 (O_349,N_49064,N_49456);
nor UO_350 (O_350,N_49961,N_49264);
nand UO_351 (O_351,N_49608,N_49905);
nor UO_352 (O_352,N_49609,N_49666);
or UO_353 (O_353,N_49377,N_49157);
or UO_354 (O_354,N_49998,N_49102);
and UO_355 (O_355,N_49189,N_49450);
and UO_356 (O_356,N_49293,N_49993);
and UO_357 (O_357,N_49931,N_49356);
or UO_358 (O_358,N_49606,N_49290);
xnor UO_359 (O_359,N_49171,N_49202);
nor UO_360 (O_360,N_49413,N_49056);
and UO_361 (O_361,N_49922,N_49876);
or UO_362 (O_362,N_49408,N_49028);
nand UO_363 (O_363,N_49772,N_49066);
or UO_364 (O_364,N_49899,N_49116);
and UO_365 (O_365,N_49034,N_49629);
or UO_366 (O_366,N_49324,N_49590);
or UO_367 (O_367,N_49697,N_49060);
nand UO_368 (O_368,N_49628,N_49703);
or UO_369 (O_369,N_49279,N_49863);
nor UO_370 (O_370,N_49437,N_49371);
nor UO_371 (O_371,N_49222,N_49555);
or UO_372 (O_372,N_49865,N_49633);
or UO_373 (O_373,N_49444,N_49690);
nand UO_374 (O_374,N_49878,N_49416);
xor UO_375 (O_375,N_49530,N_49864);
nand UO_376 (O_376,N_49153,N_49847);
nor UO_377 (O_377,N_49997,N_49476);
nor UO_378 (O_378,N_49672,N_49557);
nand UO_379 (O_379,N_49190,N_49731);
nand UO_380 (O_380,N_49663,N_49554);
or UO_381 (O_381,N_49726,N_49334);
nand UO_382 (O_382,N_49501,N_49888);
nor UO_383 (O_383,N_49683,N_49837);
nand UO_384 (O_384,N_49397,N_49779);
nor UO_385 (O_385,N_49270,N_49231);
or UO_386 (O_386,N_49567,N_49673);
or UO_387 (O_387,N_49455,N_49027);
or UO_388 (O_388,N_49449,N_49832);
xor UO_389 (O_389,N_49584,N_49874);
and UO_390 (O_390,N_49765,N_49276);
nor UO_391 (O_391,N_49610,N_49550);
or UO_392 (O_392,N_49155,N_49963);
nor UO_393 (O_393,N_49599,N_49786);
and UO_394 (O_394,N_49409,N_49314);
xnor UO_395 (O_395,N_49151,N_49163);
nor UO_396 (O_396,N_49256,N_49684);
xor UO_397 (O_397,N_49828,N_49050);
or UO_398 (O_398,N_49006,N_49936);
nor UO_399 (O_399,N_49583,N_49070);
or UO_400 (O_400,N_49958,N_49382);
xnor UO_401 (O_401,N_49771,N_49611);
and UO_402 (O_402,N_49168,N_49485);
and UO_403 (O_403,N_49702,N_49407);
xor UO_404 (O_404,N_49426,N_49849);
nor UO_405 (O_405,N_49085,N_49651);
and UO_406 (O_406,N_49235,N_49605);
or UO_407 (O_407,N_49904,N_49126);
nand UO_408 (O_408,N_49272,N_49357);
and UO_409 (O_409,N_49020,N_49493);
nor UO_410 (O_410,N_49823,N_49782);
xor UO_411 (O_411,N_49502,N_49803);
and UO_412 (O_412,N_49598,N_49636);
nor UO_413 (O_413,N_49637,N_49071);
or UO_414 (O_414,N_49239,N_49561);
nor UO_415 (O_415,N_49647,N_49586);
or UO_416 (O_416,N_49780,N_49919);
and UO_417 (O_417,N_49185,N_49128);
nor UO_418 (O_418,N_49236,N_49834);
nand UO_419 (O_419,N_49074,N_49498);
nor UO_420 (O_420,N_49920,N_49693);
nand UO_421 (O_421,N_49990,N_49713);
nand UO_422 (O_422,N_49730,N_49191);
nor UO_423 (O_423,N_49007,N_49821);
nand UO_424 (O_424,N_49259,N_49439);
or UO_425 (O_425,N_49694,N_49465);
nand UO_426 (O_426,N_49123,N_49019);
and UO_427 (O_427,N_49150,N_49010);
nand UO_428 (O_428,N_49212,N_49982);
xor UO_429 (O_429,N_49388,N_49801);
and UO_430 (O_430,N_49957,N_49440);
or UO_431 (O_431,N_49362,N_49460);
or UO_432 (O_432,N_49052,N_49695);
or UO_433 (O_433,N_49952,N_49011);
xnor UO_434 (O_434,N_49513,N_49462);
and UO_435 (O_435,N_49478,N_49291);
or UO_436 (O_436,N_49039,N_49968);
nand UO_437 (O_437,N_49900,N_49099);
nand UO_438 (O_438,N_49141,N_49499);
or UO_439 (O_439,N_49857,N_49706);
nand UO_440 (O_440,N_49574,N_49001);
and UO_441 (O_441,N_49213,N_49762);
and UO_442 (O_442,N_49491,N_49152);
xor UO_443 (O_443,N_49639,N_49238);
nor UO_444 (O_444,N_49311,N_49533);
xnor UO_445 (O_445,N_49482,N_49013);
and UO_446 (O_446,N_49641,N_49137);
nand UO_447 (O_447,N_49427,N_49436);
and UO_448 (O_448,N_49023,N_49355);
nor UO_449 (O_449,N_49885,N_49822);
xnor UO_450 (O_450,N_49909,N_49348);
xor UO_451 (O_451,N_49184,N_49349);
and UO_452 (O_452,N_49295,N_49403);
nand UO_453 (O_453,N_49897,N_49192);
and UO_454 (O_454,N_49233,N_49422);
or UO_455 (O_455,N_49454,N_49558);
xnor UO_456 (O_456,N_49321,N_49345);
nand UO_457 (O_457,N_49394,N_49870);
and UO_458 (O_458,N_49600,N_49549);
or UO_459 (O_459,N_49564,N_49727);
or UO_460 (O_460,N_49195,N_49330);
and UO_461 (O_461,N_49769,N_49630);
and UO_462 (O_462,N_49341,N_49853);
nand UO_463 (O_463,N_49209,N_49203);
or UO_464 (O_464,N_49350,N_49755);
nor UO_465 (O_465,N_49091,N_49711);
and UO_466 (O_466,N_49094,N_49329);
nand UO_467 (O_467,N_49631,N_49767);
and UO_468 (O_468,N_49361,N_49015);
nor UO_469 (O_469,N_49619,N_49869);
nand UO_470 (O_470,N_49720,N_49107);
xnor UO_471 (O_471,N_49529,N_49523);
nor UO_472 (O_472,N_49218,N_49724);
or UO_473 (O_473,N_49318,N_49723);
xor UO_474 (O_474,N_49964,N_49661);
nor UO_475 (O_475,N_49778,N_49133);
or UO_476 (O_476,N_49331,N_49883);
xor UO_477 (O_477,N_49365,N_49251);
nand UO_478 (O_478,N_49527,N_49411);
and UO_479 (O_479,N_49375,N_49275);
nor UO_480 (O_480,N_49700,N_49939);
nand UO_481 (O_481,N_49396,N_49200);
nand UO_482 (O_482,N_49054,N_49942);
xnor UO_483 (O_483,N_49479,N_49577);
nand UO_484 (O_484,N_49580,N_49901);
or UO_485 (O_485,N_49738,N_49944);
xor UO_486 (O_486,N_49260,N_49916);
nor UO_487 (O_487,N_49915,N_49848);
nor UO_488 (O_488,N_49294,N_49940);
nor UO_489 (O_489,N_49033,N_49172);
nand UO_490 (O_490,N_49241,N_49635);
xor UO_491 (O_491,N_49536,N_49617);
nor UO_492 (O_492,N_49930,N_49495);
and UO_493 (O_493,N_49472,N_49843);
nand UO_494 (O_494,N_49829,N_49768);
nor UO_495 (O_495,N_49477,N_49468);
nand UO_496 (O_496,N_49569,N_49160);
xnor UO_497 (O_497,N_49267,N_49566);
nor UO_498 (O_498,N_49668,N_49000);
or UO_499 (O_499,N_49147,N_49016);
nand UO_500 (O_500,N_49571,N_49568);
nor UO_501 (O_501,N_49207,N_49375);
xnor UO_502 (O_502,N_49801,N_49539);
and UO_503 (O_503,N_49032,N_49302);
xnor UO_504 (O_504,N_49533,N_49066);
nor UO_505 (O_505,N_49792,N_49592);
or UO_506 (O_506,N_49911,N_49386);
xnor UO_507 (O_507,N_49987,N_49351);
nand UO_508 (O_508,N_49706,N_49542);
xor UO_509 (O_509,N_49139,N_49095);
xor UO_510 (O_510,N_49857,N_49966);
or UO_511 (O_511,N_49128,N_49494);
or UO_512 (O_512,N_49106,N_49305);
nor UO_513 (O_513,N_49561,N_49949);
or UO_514 (O_514,N_49437,N_49761);
nor UO_515 (O_515,N_49352,N_49022);
xnor UO_516 (O_516,N_49315,N_49897);
or UO_517 (O_517,N_49571,N_49640);
xor UO_518 (O_518,N_49161,N_49004);
nor UO_519 (O_519,N_49348,N_49440);
nand UO_520 (O_520,N_49390,N_49664);
nor UO_521 (O_521,N_49187,N_49769);
or UO_522 (O_522,N_49207,N_49182);
xnor UO_523 (O_523,N_49416,N_49273);
or UO_524 (O_524,N_49559,N_49110);
nand UO_525 (O_525,N_49339,N_49095);
xor UO_526 (O_526,N_49357,N_49662);
nand UO_527 (O_527,N_49074,N_49680);
xor UO_528 (O_528,N_49621,N_49683);
xor UO_529 (O_529,N_49498,N_49418);
nor UO_530 (O_530,N_49886,N_49144);
and UO_531 (O_531,N_49860,N_49140);
nor UO_532 (O_532,N_49734,N_49855);
nor UO_533 (O_533,N_49496,N_49543);
nand UO_534 (O_534,N_49393,N_49543);
xnor UO_535 (O_535,N_49813,N_49901);
and UO_536 (O_536,N_49508,N_49964);
and UO_537 (O_537,N_49256,N_49736);
xnor UO_538 (O_538,N_49275,N_49365);
and UO_539 (O_539,N_49474,N_49734);
nand UO_540 (O_540,N_49524,N_49177);
or UO_541 (O_541,N_49045,N_49894);
xnor UO_542 (O_542,N_49534,N_49340);
nor UO_543 (O_543,N_49527,N_49795);
xor UO_544 (O_544,N_49252,N_49335);
nand UO_545 (O_545,N_49813,N_49240);
nor UO_546 (O_546,N_49825,N_49333);
nor UO_547 (O_547,N_49990,N_49392);
or UO_548 (O_548,N_49134,N_49873);
nand UO_549 (O_549,N_49008,N_49589);
nand UO_550 (O_550,N_49855,N_49147);
xnor UO_551 (O_551,N_49676,N_49938);
xnor UO_552 (O_552,N_49427,N_49452);
nand UO_553 (O_553,N_49656,N_49550);
or UO_554 (O_554,N_49281,N_49994);
xnor UO_555 (O_555,N_49367,N_49088);
nor UO_556 (O_556,N_49324,N_49940);
xor UO_557 (O_557,N_49503,N_49322);
nand UO_558 (O_558,N_49537,N_49761);
or UO_559 (O_559,N_49354,N_49583);
xor UO_560 (O_560,N_49823,N_49405);
xor UO_561 (O_561,N_49441,N_49034);
nand UO_562 (O_562,N_49739,N_49524);
and UO_563 (O_563,N_49085,N_49375);
nand UO_564 (O_564,N_49673,N_49339);
xor UO_565 (O_565,N_49024,N_49548);
or UO_566 (O_566,N_49193,N_49439);
nand UO_567 (O_567,N_49007,N_49021);
or UO_568 (O_568,N_49388,N_49076);
nand UO_569 (O_569,N_49332,N_49856);
xnor UO_570 (O_570,N_49053,N_49304);
or UO_571 (O_571,N_49401,N_49999);
nand UO_572 (O_572,N_49666,N_49989);
or UO_573 (O_573,N_49665,N_49475);
and UO_574 (O_574,N_49045,N_49451);
xor UO_575 (O_575,N_49525,N_49560);
nor UO_576 (O_576,N_49357,N_49945);
and UO_577 (O_577,N_49626,N_49361);
nor UO_578 (O_578,N_49315,N_49706);
nor UO_579 (O_579,N_49636,N_49811);
and UO_580 (O_580,N_49770,N_49473);
or UO_581 (O_581,N_49446,N_49010);
xor UO_582 (O_582,N_49247,N_49554);
nor UO_583 (O_583,N_49370,N_49260);
or UO_584 (O_584,N_49850,N_49939);
nor UO_585 (O_585,N_49106,N_49148);
or UO_586 (O_586,N_49607,N_49989);
nor UO_587 (O_587,N_49922,N_49440);
nand UO_588 (O_588,N_49531,N_49289);
or UO_589 (O_589,N_49154,N_49776);
nand UO_590 (O_590,N_49663,N_49629);
and UO_591 (O_591,N_49078,N_49029);
or UO_592 (O_592,N_49045,N_49789);
nand UO_593 (O_593,N_49631,N_49009);
or UO_594 (O_594,N_49664,N_49201);
and UO_595 (O_595,N_49947,N_49500);
xor UO_596 (O_596,N_49509,N_49103);
nor UO_597 (O_597,N_49088,N_49343);
xor UO_598 (O_598,N_49779,N_49552);
nand UO_599 (O_599,N_49037,N_49560);
or UO_600 (O_600,N_49164,N_49858);
nor UO_601 (O_601,N_49397,N_49465);
nor UO_602 (O_602,N_49678,N_49454);
or UO_603 (O_603,N_49651,N_49424);
nand UO_604 (O_604,N_49499,N_49073);
nor UO_605 (O_605,N_49074,N_49234);
or UO_606 (O_606,N_49276,N_49073);
and UO_607 (O_607,N_49559,N_49738);
and UO_608 (O_608,N_49374,N_49101);
or UO_609 (O_609,N_49579,N_49562);
or UO_610 (O_610,N_49295,N_49060);
nor UO_611 (O_611,N_49564,N_49329);
nand UO_612 (O_612,N_49992,N_49112);
xnor UO_613 (O_613,N_49237,N_49661);
or UO_614 (O_614,N_49387,N_49854);
and UO_615 (O_615,N_49670,N_49971);
xnor UO_616 (O_616,N_49645,N_49339);
nand UO_617 (O_617,N_49713,N_49133);
and UO_618 (O_618,N_49564,N_49926);
and UO_619 (O_619,N_49186,N_49823);
and UO_620 (O_620,N_49793,N_49644);
nand UO_621 (O_621,N_49386,N_49763);
or UO_622 (O_622,N_49331,N_49025);
nand UO_623 (O_623,N_49865,N_49065);
nand UO_624 (O_624,N_49292,N_49959);
nor UO_625 (O_625,N_49500,N_49580);
nand UO_626 (O_626,N_49383,N_49003);
xnor UO_627 (O_627,N_49430,N_49387);
xnor UO_628 (O_628,N_49892,N_49084);
nand UO_629 (O_629,N_49365,N_49253);
and UO_630 (O_630,N_49494,N_49036);
or UO_631 (O_631,N_49438,N_49331);
or UO_632 (O_632,N_49764,N_49804);
nor UO_633 (O_633,N_49472,N_49556);
nand UO_634 (O_634,N_49822,N_49170);
and UO_635 (O_635,N_49713,N_49122);
nor UO_636 (O_636,N_49279,N_49178);
nand UO_637 (O_637,N_49666,N_49505);
nor UO_638 (O_638,N_49673,N_49561);
and UO_639 (O_639,N_49663,N_49154);
and UO_640 (O_640,N_49646,N_49925);
nor UO_641 (O_641,N_49614,N_49978);
nand UO_642 (O_642,N_49590,N_49870);
xnor UO_643 (O_643,N_49165,N_49334);
nand UO_644 (O_644,N_49802,N_49734);
xor UO_645 (O_645,N_49419,N_49591);
nand UO_646 (O_646,N_49571,N_49534);
or UO_647 (O_647,N_49737,N_49953);
and UO_648 (O_648,N_49637,N_49436);
nor UO_649 (O_649,N_49816,N_49842);
xnor UO_650 (O_650,N_49326,N_49482);
nor UO_651 (O_651,N_49416,N_49200);
or UO_652 (O_652,N_49843,N_49105);
xor UO_653 (O_653,N_49631,N_49044);
nand UO_654 (O_654,N_49578,N_49027);
or UO_655 (O_655,N_49810,N_49356);
and UO_656 (O_656,N_49650,N_49022);
and UO_657 (O_657,N_49023,N_49811);
nor UO_658 (O_658,N_49908,N_49029);
or UO_659 (O_659,N_49690,N_49591);
and UO_660 (O_660,N_49938,N_49023);
xor UO_661 (O_661,N_49734,N_49584);
xnor UO_662 (O_662,N_49927,N_49254);
nand UO_663 (O_663,N_49796,N_49845);
and UO_664 (O_664,N_49097,N_49695);
and UO_665 (O_665,N_49858,N_49361);
or UO_666 (O_666,N_49637,N_49629);
xnor UO_667 (O_667,N_49096,N_49320);
nor UO_668 (O_668,N_49502,N_49688);
or UO_669 (O_669,N_49325,N_49619);
and UO_670 (O_670,N_49287,N_49506);
xor UO_671 (O_671,N_49691,N_49094);
nor UO_672 (O_672,N_49967,N_49438);
nor UO_673 (O_673,N_49780,N_49477);
xnor UO_674 (O_674,N_49376,N_49810);
and UO_675 (O_675,N_49223,N_49086);
nand UO_676 (O_676,N_49187,N_49403);
and UO_677 (O_677,N_49535,N_49716);
and UO_678 (O_678,N_49376,N_49005);
nand UO_679 (O_679,N_49643,N_49132);
or UO_680 (O_680,N_49377,N_49996);
and UO_681 (O_681,N_49340,N_49815);
or UO_682 (O_682,N_49371,N_49630);
xor UO_683 (O_683,N_49562,N_49818);
and UO_684 (O_684,N_49526,N_49553);
or UO_685 (O_685,N_49399,N_49496);
xor UO_686 (O_686,N_49177,N_49979);
and UO_687 (O_687,N_49773,N_49963);
nor UO_688 (O_688,N_49129,N_49417);
xor UO_689 (O_689,N_49300,N_49485);
nor UO_690 (O_690,N_49952,N_49219);
and UO_691 (O_691,N_49453,N_49748);
nand UO_692 (O_692,N_49423,N_49886);
nor UO_693 (O_693,N_49615,N_49691);
or UO_694 (O_694,N_49267,N_49940);
and UO_695 (O_695,N_49466,N_49271);
xor UO_696 (O_696,N_49791,N_49769);
or UO_697 (O_697,N_49481,N_49337);
nor UO_698 (O_698,N_49107,N_49131);
and UO_699 (O_699,N_49791,N_49336);
nor UO_700 (O_700,N_49807,N_49165);
nand UO_701 (O_701,N_49028,N_49275);
nand UO_702 (O_702,N_49607,N_49566);
and UO_703 (O_703,N_49615,N_49976);
nor UO_704 (O_704,N_49023,N_49104);
nand UO_705 (O_705,N_49046,N_49306);
nand UO_706 (O_706,N_49065,N_49158);
or UO_707 (O_707,N_49823,N_49431);
or UO_708 (O_708,N_49444,N_49470);
xor UO_709 (O_709,N_49389,N_49656);
and UO_710 (O_710,N_49530,N_49080);
xnor UO_711 (O_711,N_49030,N_49639);
or UO_712 (O_712,N_49871,N_49175);
xnor UO_713 (O_713,N_49933,N_49820);
or UO_714 (O_714,N_49327,N_49948);
nor UO_715 (O_715,N_49482,N_49599);
or UO_716 (O_716,N_49387,N_49194);
nand UO_717 (O_717,N_49493,N_49843);
or UO_718 (O_718,N_49703,N_49600);
and UO_719 (O_719,N_49426,N_49742);
or UO_720 (O_720,N_49827,N_49439);
or UO_721 (O_721,N_49237,N_49179);
or UO_722 (O_722,N_49979,N_49163);
nand UO_723 (O_723,N_49387,N_49617);
nand UO_724 (O_724,N_49558,N_49593);
xnor UO_725 (O_725,N_49804,N_49224);
nand UO_726 (O_726,N_49226,N_49330);
and UO_727 (O_727,N_49880,N_49770);
nand UO_728 (O_728,N_49033,N_49902);
and UO_729 (O_729,N_49537,N_49333);
xor UO_730 (O_730,N_49994,N_49094);
or UO_731 (O_731,N_49750,N_49101);
nor UO_732 (O_732,N_49941,N_49794);
nand UO_733 (O_733,N_49989,N_49739);
or UO_734 (O_734,N_49417,N_49827);
and UO_735 (O_735,N_49628,N_49621);
and UO_736 (O_736,N_49439,N_49693);
or UO_737 (O_737,N_49158,N_49408);
and UO_738 (O_738,N_49207,N_49189);
nand UO_739 (O_739,N_49517,N_49487);
nand UO_740 (O_740,N_49766,N_49393);
nand UO_741 (O_741,N_49730,N_49133);
nand UO_742 (O_742,N_49747,N_49854);
nor UO_743 (O_743,N_49099,N_49503);
and UO_744 (O_744,N_49224,N_49269);
or UO_745 (O_745,N_49764,N_49597);
xnor UO_746 (O_746,N_49117,N_49228);
or UO_747 (O_747,N_49177,N_49323);
nor UO_748 (O_748,N_49457,N_49907);
nor UO_749 (O_749,N_49266,N_49529);
or UO_750 (O_750,N_49519,N_49159);
nor UO_751 (O_751,N_49814,N_49241);
or UO_752 (O_752,N_49109,N_49474);
or UO_753 (O_753,N_49842,N_49040);
or UO_754 (O_754,N_49219,N_49518);
nor UO_755 (O_755,N_49381,N_49684);
or UO_756 (O_756,N_49419,N_49056);
xor UO_757 (O_757,N_49909,N_49889);
or UO_758 (O_758,N_49439,N_49832);
or UO_759 (O_759,N_49575,N_49456);
nor UO_760 (O_760,N_49880,N_49700);
or UO_761 (O_761,N_49488,N_49105);
and UO_762 (O_762,N_49057,N_49759);
nand UO_763 (O_763,N_49310,N_49326);
nand UO_764 (O_764,N_49302,N_49440);
and UO_765 (O_765,N_49831,N_49161);
xnor UO_766 (O_766,N_49911,N_49491);
or UO_767 (O_767,N_49493,N_49781);
nor UO_768 (O_768,N_49738,N_49494);
nor UO_769 (O_769,N_49964,N_49043);
nor UO_770 (O_770,N_49839,N_49918);
and UO_771 (O_771,N_49137,N_49888);
nor UO_772 (O_772,N_49642,N_49123);
or UO_773 (O_773,N_49869,N_49601);
nor UO_774 (O_774,N_49211,N_49032);
nand UO_775 (O_775,N_49953,N_49537);
and UO_776 (O_776,N_49781,N_49512);
xnor UO_777 (O_777,N_49685,N_49191);
or UO_778 (O_778,N_49261,N_49848);
nand UO_779 (O_779,N_49371,N_49133);
nor UO_780 (O_780,N_49765,N_49481);
nor UO_781 (O_781,N_49176,N_49360);
xor UO_782 (O_782,N_49273,N_49024);
or UO_783 (O_783,N_49757,N_49253);
or UO_784 (O_784,N_49070,N_49954);
nor UO_785 (O_785,N_49691,N_49988);
nand UO_786 (O_786,N_49796,N_49462);
nand UO_787 (O_787,N_49105,N_49603);
nand UO_788 (O_788,N_49980,N_49209);
and UO_789 (O_789,N_49737,N_49003);
xnor UO_790 (O_790,N_49170,N_49106);
nor UO_791 (O_791,N_49259,N_49572);
nand UO_792 (O_792,N_49685,N_49953);
and UO_793 (O_793,N_49337,N_49491);
nor UO_794 (O_794,N_49826,N_49577);
xnor UO_795 (O_795,N_49582,N_49827);
or UO_796 (O_796,N_49857,N_49309);
and UO_797 (O_797,N_49142,N_49029);
and UO_798 (O_798,N_49953,N_49599);
nor UO_799 (O_799,N_49859,N_49564);
nand UO_800 (O_800,N_49551,N_49942);
nor UO_801 (O_801,N_49652,N_49593);
and UO_802 (O_802,N_49276,N_49853);
or UO_803 (O_803,N_49263,N_49379);
xor UO_804 (O_804,N_49169,N_49125);
or UO_805 (O_805,N_49470,N_49788);
nor UO_806 (O_806,N_49035,N_49834);
nand UO_807 (O_807,N_49061,N_49046);
or UO_808 (O_808,N_49531,N_49708);
nor UO_809 (O_809,N_49636,N_49996);
and UO_810 (O_810,N_49571,N_49849);
or UO_811 (O_811,N_49649,N_49012);
and UO_812 (O_812,N_49353,N_49714);
nor UO_813 (O_813,N_49050,N_49756);
and UO_814 (O_814,N_49122,N_49228);
nor UO_815 (O_815,N_49568,N_49657);
nand UO_816 (O_816,N_49003,N_49647);
nor UO_817 (O_817,N_49091,N_49586);
or UO_818 (O_818,N_49112,N_49855);
nand UO_819 (O_819,N_49134,N_49916);
xor UO_820 (O_820,N_49626,N_49920);
and UO_821 (O_821,N_49211,N_49639);
or UO_822 (O_822,N_49047,N_49435);
xor UO_823 (O_823,N_49211,N_49029);
xnor UO_824 (O_824,N_49533,N_49041);
and UO_825 (O_825,N_49091,N_49865);
xor UO_826 (O_826,N_49707,N_49375);
or UO_827 (O_827,N_49775,N_49687);
or UO_828 (O_828,N_49662,N_49978);
nor UO_829 (O_829,N_49272,N_49748);
nor UO_830 (O_830,N_49640,N_49023);
nor UO_831 (O_831,N_49851,N_49613);
xor UO_832 (O_832,N_49922,N_49776);
and UO_833 (O_833,N_49148,N_49543);
or UO_834 (O_834,N_49933,N_49212);
nor UO_835 (O_835,N_49403,N_49484);
xnor UO_836 (O_836,N_49490,N_49067);
nand UO_837 (O_837,N_49234,N_49785);
nand UO_838 (O_838,N_49487,N_49349);
and UO_839 (O_839,N_49309,N_49867);
or UO_840 (O_840,N_49326,N_49410);
nand UO_841 (O_841,N_49515,N_49940);
xnor UO_842 (O_842,N_49213,N_49745);
and UO_843 (O_843,N_49967,N_49491);
or UO_844 (O_844,N_49238,N_49224);
and UO_845 (O_845,N_49018,N_49386);
nand UO_846 (O_846,N_49609,N_49329);
xor UO_847 (O_847,N_49049,N_49487);
nand UO_848 (O_848,N_49332,N_49336);
nor UO_849 (O_849,N_49696,N_49381);
and UO_850 (O_850,N_49694,N_49516);
and UO_851 (O_851,N_49500,N_49218);
xnor UO_852 (O_852,N_49264,N_49482);
nand UO_853 (O_853,N_49117,N_49779);
and UO_854 (O_854,N_49013,N_49153);
and UO_855 (O_855,N_49425,N_49958);
nand UO_856 (O_856,N_49374,N_49358);
xnor UO_857 (O_857,N_49824,N_49768);
or UO_858 (O_858,N_49109,N_49724);
nand UO_859 (O_859,N_49107,N_49628);
nand UO_860 (O_860,N_49866,N_49897);
or UO_861 (O_861,N_49922,N_49836);
xnor UO_862 (O_862,N_49834,N_49209);
nor UO_863 (O_863,N_49584,N_49062);
and UO_864 (O_864,N_49855,N_49412);
xor UO_865 (O_865,N_49753,N_49325);
or UO_866 (O_866,N_49841,N_49174);
xor UO_867 (O_867,N_49972,N_49913);
or UO_868 (O_868,N_49336,N_49625);
or UO_869 (O_869,N_49030,N_49210);
xor UO_870 (O_870,N_49042,N_49857);
or UO_871 (O_871,N_49269,N_49023);
or UO_872 (O_872,N_49684,N_49881);
or UO_873 (O_873,N_49231,N_49366);
and UO_874 (O_874,N_49861,N_49804);
xnor UO_875 (O_875,N_49809,N_49573);
nand UO_876 (O_876,N_49046,N_49742);
nor UO_877 (O_877,N_49969,N_49342);
or UO_878 (O_878,N_49827,N_49960);
xnor UO_879 (O_879,N_49017,N_49246);
and UO_880 (O_880,N_49564,N_49040);
nand UO_881 (O_881,N_49569,N_49137);
nor UO_882 (O_882,N_49459,N_49931);
nor UO_883 (O_883,N_49883,N_49566);
or UO_884 (O_884,N_49506,N_49909);
nand UO_885 (O_885,N_49129,N_49125);
nor UO_886 (O_886,N_49306,N_49279);
xnor UO_887 (O_887,N_49279,N_49952);
or UO_888 (O_888,N_49766,N_49208);
xor UO_889 (O_889,N_49621,N_49816);
and UO_890 (O_890,N_49730,N_49986);
xor UO_891 (O_891,N_49925,N_49841);
nor UO_892 (O_892,N_49687,N_49652);
xnor UO_893 (O_893,N_49468,N_49557);
or UO_894 (O_894,N_49758,N_49322);
and UO_895 (O_895,N_49940,N_49371);
nand UO_896 (O_896,N_49562,N_49464);
and UO_897 (O_897,N_49880,N_49954);
and UO_898 (O_898,N_49821,N_49584);
nor UO_899 (O_899,N_49410,N_49567);
and UO_900 (O_900,N_49356,N_49214);
nor UO_901 (O_901,N_49449,N_49896);
xor UO_902 (O_902,N_49732,N_49020);
nand UO_903 (O_903,N_49194,N_49588);
nand UO_904 (O_904,N_49398,N_49015);
and UO_905 (O_905,N_49950,N_49502);
or UO_906 (O_906,N_49164,N_49806);
and UO_907 (O_907,N_49840,N_49934);
nor UO_908 (O_908,N_49152,N_49595);
nand UO_909 (O_909,N_49477,N_49377);
nor UO_910 (O_910,N_49247,N_49660);
xnor UO_911 (O_911,N_49604,N_49948);
and UO_912 (O_912,N_49455,N_49996);
xor UO_913 (O_913,N_49587,N_49675);
xnor UO_914 (O_914,N_49641,N_49324);
xor UO_915 (O_915,N_49229,N_49406);
nand UO_916 (O_916,N_49557,N_49346);
xnor UO_917 (O_917,N_49214,N_49640);
xor UO_918 (O_918,N_49886,N_49103);
nand UO_919 (O_919,N_49009,N_49310);
or UO_920 (O_920,N_49521,N_49195);
or UO_921 (O_921,N_49930,N_49646);
nor UO_922 (O_922,N_49321,N_49979);
nand UO_923 (O_923,N_49247,N_49674);
nor UO_924 (O_924,N_49878,N_49710);
nor UO_925 (O_925,N_49631,N_49334);
nor UO_926 (O_926,N_49180,N_49556);
and UO_927 (O_927,N_49918,N_49400);
or UO_928 (O_928,N_49302,N_49468);
xor UO_929 (O_929,N_49064,N_49864);
xnor UO_930 (O_930,N_49708,N_49178);
xor UO_931 (O_931,N_49804,N_49083);
nand UO_932 (O_932,N_49975,N_49277);
or UO_933 (O_933,N_49719,N_49026);
nand UO_934 (O_934,N_49734,N_49582);
or UO_935 (O_935,N_49433,N_49603);
nor UO_936 (O_936,N_49661,N_49293);
nor UO_937 (O_937,N_49153,N_49264);
nor UO_938 (O_938,N_49904,N_49484);
xnor UO_939 (O_939,N_49475,N_49791);
xnor UO_940 (O_940,N_49556,N_49641);
or UO_941 (O_941,N_49438,N_49985);
or UO_942 (O_942,N_49718,N_49114);
nand UO_943 (O_943,N_49324,N_49604);
or UO_944 (O_944,N_49545,N_49803);
or UO_945 (O_945,N_49061,N_49621);
and UO_946 (O_946,N_49991,N_49413);
or UO_947 (O_947,N_49295,N_49766);
and UO_948 (O_948,N_49917,N_49901);
nor UO_949 (O_949,N_49460,N_49788);
nand UO_950 (O_950,N_49291,N_49820);
nor UO_951 (O_951,N_49006,N_49267);
nor UO_952 (O_952,N_49072,N_49896);
xor UO_953 (O_953,N_49086,N_49923);
or UO_954 (O_954,N_49598,N_49529);
nand UO_955 (O_955,N_49335,N_49330);
or UO_956 (O_956,N_49754,N_49159);
and UO_957 (O_957,N_49624,N_49863);
xnor UO_958 (O_958,N_49902,N_49963);
xnor UO_959 (O_959,N_49613,N_49329);
nor UO_960 (O_960,N_49401,N_49998);
nand UO_961 (O_961,N_49558,N_49598);
nor UO_962 (O_962,N_49900,N_49515);
and UO_963 (O_963,N_49465,N_49128);
xor UO_964 (O_964,N_49143,N_49535);
xor UO_965 (O_965,N_49656,N_49213);
and UO_966 (O_966,N_49066,N_49249);
xor UO_967 (O_967,N_49415,N_49956);
or UO_968 (O_968,N_49334,N_49364);
or UO_969 (O_969,N_49881,N_49992);
or UO_970 (O_970,N_49797,N_49599);
nand UO_971 (O_971,N_49827,N_49636);
or UO_972 (O_972,N_49767,N_49040);
nand UO_973 (O_973,N_49964,N_49004);
or UO_974 (O_974,N_49593,N_49535);
nand UO_975 (O_975,N_49535,N_49243);
nand UO_976 (O_976,N_49959,N_49527);
and UO_977 (O_977,N_49363,N_49642);
xnor UO_978 (O_978,N_49744,N_49035);
nand UO_979 (O_979,N_49745,N_49826);
or UO_980 (O_980,N_49678,N_49850);
xnor UO_981 (O_981,N_49681,N_49276);
nand UO_982 (O_982,N_49584,N_49525);
xor UO_983 (O_983,N_49998,N_49083);
xnor UO_984 (O_984,N_49749,N_49006);
nor UO_985 (O_985,N_49283,N_49363);
or UO_986 (O_986,N_49465,N_49353);
xor UO_987 (O_987,N_49341,N_49322);
and UO_988 (O_988,N_49431,N_49002);
nand UO_989 (O_989,N_49494,N_49294);
xnor UO_990 (O_990,N_49414,N_49942);
xor UO_991 (O_991,N_49447,N_49491);
or UO_992 (O_992,N_49346,N_49985);
nand UO_993 (O_993,N_49702,N_49821);
and UO_994 (O_994,N_49844,N_49760);
and UO_995 (O_995,N_49966,N_49771);
or UO_996 (O_996,N_49796,N_49619);
or UO_997 (O_997,N_49413,N_49319);
nand UO_998 (O_998,N_49469,N_49623);
xor UO_999 (O_999,N_49440,N_49946);
nand UO_1000 (O_1000,N_49124,N_49708);
xnor UO_1001 (O_1001,N_49192,N_49798);
nor UO_1002 (O_1002,N_49402,N_49109);
and UO_1003 (O_1003,N_49508,N_49205);
xor UO_1004 (O_1004,N_49322,N_49014);
nand UO_1005 (O_1005,N_49065,N_49464);
or UO_1006 (O_1006,N_49995,N_49846);
xor UO_1007 (O_1007,N_49540,N_49390);
and UO_1008 (O_1008,N_49836,N_49167);
xnor UO_1009 (O_1009,N_49483,N_49496);
nor UO_1010 (O_1010,N_49084,N_49443);
and UO_1011 (O_1011,N_49099,N_49955);
xor UO_1012 (O_1012,N_49779,N_49217);
xnor UO_1013 (O_1013,N_49076,N_49675);
nor UO_1014 (O_1014,N_49797,N_49815);
nand UO_1015 (O_1015,N_49004,N_49227);
or UO_1016 (O_1016,N_49460,N_49938);
or UO_1017 (O_1017,N_49882,N_49012);
xnor UO_1018 (O_1018,N_49832,N_49239);
nor UO_1019 (O_1019,N_49794,N_49618);
and UO_1020 (O_1020,N_49108,N_49069);
nor UO_1021 (O_1021,N_49515,N_49021);
or UO_1022 (O_1022,N_49785,N_49565);
nor UO_1023 (O_1023,N_49777,N_49696);
or UO_1024 (O_1024,N_49460,N_49798);
or UO_1025 (O_1025,N_49921,N_49616);
and UO_1026 (O_1026,N_49508,N_49628);
nor UO_1027 (O_1027,N_49504,N_49353);
nand UO_1028 (O_1028,N_49742,N_49512);
xor UO_1029 (O_1029,N_49300,N_49554);
or UO_1030 (O_1030,N_49444,N_49911);
nand UO_1031 (O_1031,N_49854,N_49224);
nand UO_1032 (O_1032,N_49457,N_49313);
or UO_1033 (O_1033,N_49651,N_49603);
xor UO_1034 (O_1034,N_49152,N_49084);
and UO_1035 (O_1035,N_49162,N_49309);
and UO_1036 (O_1036,N_49259,N_49743);
nor UO_1037 (O_1037,N_49593,N_49934);
nor UO_1038 (O_1038,N_49334,N_49079);
or UO_1039 (O_1039,N_49532,N_49460);
and UO_1040 (O_1040,N_49210,N_49278);
and UO_1041 (O_1041,N_49530,N_49624);
xor UO_1042 (O_1042,N_49574,N_49839);
xnor UO_1043 (O_1043,N_49587,N_49306);
and UO_1044 (O_1044,N_49504,N_49839);
nor UO_1045 (O_1045,N_49795,N_49685);
and UO_1046 (O_1046,N_49460,N_49596);
or UO_1047 (O_1047,N_49072,N_49912);
xnor UO_1048 (O_1048,N_49750,N_49110);
and UO_1049 (O_1049,N_49388,N_49613);
nor UO_1050 (O_1050,N_49639,N_49341);
and UO_1051 (O_1051,N_49588,N_49744);
and UO_1052 (O_1052,N_49110,N_49278);
and UO_1053 (O_1053,N_49951,N_49392);
and UO_1054 (O_1054,N_49705,N_49799);
nor UO_1055 (O_1055,N_49946,N_49998);
or UO_1056 (O_1056,N_49690,N_49956);
nand UO_1057 (O_1057,N_49965,N_49344);
and UO_1058 (O_1058,N_49746,N_49352);
nand UO_1059 (O_1059,N_49978,N_49987);
or UO_1060 (O_1060,N_49077,N_49496);
nor UO_1061 (O_1061,N_49855,N_49744);
and UO_1062 (O_1062,N_49471,N_49209);
nor UO_1063 (O_1063,N_49144,N_49084);
and UO_1064 (O_1064,N_49300,N_49039);
or UO_1065 (O_1065,N_49949,N_49113);
nor UO_1066 (O_1066,N_49228,N_49867);
xor UO_1067 (O_1067,N_49813,N_49365);
and UO_1068 (O_1068,N_49602,N_49364);
nor UO_1069 (O_1069,N_49162,N_49623);
xor UO_1070 (O_1070,N_49271,N_49616);
nand UO_1071 (O_1071,N_49867,N_49333);
or UO_1072 (O_1072,N_49116,N_49007);
and UO_1073 (O_1073,N_49668,N_49438);
and UO_1074 (O_1074,N_49975,N_49819);
nand UO_1075 (O_1075,N_49901,N_49046);
xnor UO_1076 (O_1076,N_49269,N_49495);
nand UO_1077 (O_1077,N_49594,N_49784);
nor UO_1078 (O_1078,N_49050,N_49839);
xor UO_1079 (O_1079,N_49326,N_49367);
or UO_1080 (O_1080,N_49737,N_49186);
or UO_1081 (O_1081,N_49093,N_49882);
nand UO_1082 (O_1082,N_49725,N_49463);
xnor UO_1083 (O_1083,N_49149,N_49922);
xor UO_1084 (O_1084,N_49554,N_49079);
xnor UO_1085 (O_1085,N_49843,N_49217);
nand UO_1086 (O_1086,N_49055,N_49702);
nand UO_1087 (O_1087,N_49909,N_49618);
xnor UO_1088 (O_1088,N_49676,N_49953);
and UO_1089 (O_1089,N_49288,N_49830);
nand UO_1090 (O_1090,N_49192,N_49693);
or UO_1091 (O_1091,N_49742,N_49770);
and UO_1092 (O_1092,N_49599,N_49011);
xnor UO_1093 (O_1093,N_49589,N_49677);
nand UO_1094 (O_1094,N_49580,N_49992);
xnor UO_1095 (O_1095,N_49922,N_49505);
and UO_1096 (O_1096,N_49193,N_49287);
or UO_1097 (O_1097,N_49276,N_49963);
nand UO_1098 (O_1098,N_49305,N_49230);
and UO_1099 (O_1099,N_49060,N_49800);
nor UO_1100 (O_1100,N_49981,N_49172);
nor UO_1101 (O_1101,N_49578,N_49959);
xor UO_1102 (O_1102,N_49481,N_49871);
xnor UO_1103 (O_1103,N_49391,N_49387);
or UO_1104 (O_1104,N_49722,N_49432);
nor UO_1105 (O_1105,N_49711,N_49997);
and UO_1106 (O_1106,N_49625,N_49606);
and UO_1107 (O_1107,N_49144,N_49518);
xnor UO_1108 (O_1108,N_49444,N_49736);
nand UO_1109 (O_1109,N_49540,N_49442);
and UO_1110 (O_1110,N_49389,N_49207);
nor UO_1111 (O_1111,N_49805,N_49473);
or UO_1112 (O_1112,N_49943,N_49450);
or UO_1113 (O_1113,N_49883,N_49546);
xor UO_1114 (O_1114,N_49978,N_49603);
xor UO_1115 (O_1115,N_49907,N_49060);
xor UO_1116 (O_1116,N_49543,N_49546);
xnor UO_1117 (O_1117,N_49409,N_49887);
nor UO_1118 (O_1118,N_49397,N_49509);
nor UO_1119 (O_1119,N_49155,N_49456);
or UO_1120 (O_1120,N_49554,N_49796);
and UO_1121 (O_1121,N_49297,N_49995);
nor UO_1122 (O_1122,N_49907,N_49999);
xor UO_1123 (O_1123,N_49292,N_49300);
nand UO_1124 (O_1124,N_49046,N_49127);
nand UO_1125 (O_1125,N_49703,N_49511);
and UO_1126 (O_1126,N_49921,N_49314);
or UO_1127 (O_1127,N_49747,N_49612);
nor UO_1128 (O_1128,N_49826,N_49776);
nor UO_1129 (O_1129,N_49819,N_49038);
nor UO_1130 (O_1130,N_49307,N_49051);
and UO_1131 (O_1131,N_49497,N_49827);
xnor UO_1132 (O_1132,N_49592,N_49608);
nor UO_1133 (O_1133,N_49709,N_49766);
nor UO_1134 (O_1134,N_49201,N_49659);
xnor UO_1135 (O_1135,N_49404,N_49631);
nand UO_1136 (O_1136,N_49010,N_49833);
or UO_1137 (O_1137,N_49451,N_49352);
and UO_1138 (O_1138,N_49383,N_49263);
nand UO_1139 (O_1139,N_49110,N_49306);
nor UO_1140 (O_1140,N_49872,N_49238);
and UO_1141 (O_1141,N_49097,N_49552);
nor UO_1142 (O_1142,N_49620,N_49832);
or UO_1143 (O_1143,N_49254,N_49514);
and UO_1144 (O_1144,N_49682,N_49658);
nand UO_1145 (O_1145,N_49137,N_49451);
or UO_1146 (O_1146,N_49207,N_49964);
and UO_1147 (O_1147,N_49819,N_49244);
or UO_1148 (O_1148,N_49904,N_49423);
and UO_1149 (O_1149,N_49782,N_49603);
nor UO_1150 (O_1150,N_49166,N_49502);
or UO_1151 (O_1151,N_49995,N_49435);
nor UO_1152 (O_1152,N_49103,N_49477);
nand UO_1153 (O_1153,N_49345,N_49837);
nor UO_1154 (O_1154,N_49380,N_49870);
xor UO_1155 (O_1155,N_49394,N_49999);
nor UO_1156 (O_1156,N_49693,N_49800);
xnor UO_1157 (O_1157,N_49360,N_49264);
xnor UO_1158 (O_1158,N_49306,N_49996);
and UO_1159 (O_1159,N_49708,N_49300);
or UO_1160 (O_1160,N_49081,N_49337);
nor UO_1161 (O_1161,N_49757,N_49594);
nand UO_1162 (O_1162,N_49869,N_49908);
and UO_1163 (O_1163,N_49961,N_49480);
and UO_1164 (O_1164,N_49719,N_49191);
nand UO_1165 (O_1165,N_49329,N_49391);
and UO_1166 (O_1166,N_49164,N_49761);
and UO_1167 (O_1167,N_49549,N_49464);
nand UO_1168 (O_1168,N_49785,N_49668);
or UO_1169 (O_1169,N_49128,N_49481);
or UO_1170 (O_1170,N_49258,N_49217);
and UO_1171 (O_1171,N_49281,N_49548);
nor UO_1172 (O_1172,N_49953,N_49893);
and UO_1173 (O_1173,N_49189,N_49077);
or UO_1174 (O_1174,N_49413,N_49762);
xnor UO_1175 (O_1175,N_49678,N_49504);
or UO_1176 (O_1176,N_49953,N_49759);
xnor UO_1177 (O_1177,N_49827,N_49640);
xnor UO_1178 (O_1178,N_49247,N_49621);
nand UO_1179 (O_1179,N_49145,N_49966);
nand UO_1180 (O_1180,N_49011,N_49557);
nor UO_1181 (O_1181,N_49285,N_49922);
and UO_1182 (O_1182,N_49432,N_49366);
xnor UO_1183 (O_1183,N_49746,N_49357);
or UO_1184 (O_1184,N_49847,N_49887);
nand UO_1185 (O_1185,N_49707,N_49968);
nor UO_1186 (O_1186,N_49478,N_49537);
nor UO_1187 (O_1187,N_49222,N_49549);
nand UO_1188 (O_1188,N_49425,N_49461);
nand UO_1189 (O_1189,N_49106,N_49910);
nor UO_1190 (O_1190,N_49182,N_49869);
nor UO_1191 (O_1191,N_49934,N_49931);
nor UO_1192 (O_1192,N_49223,N_49649);
xnor UO_1193 (O_1193,N_49249,N_49379);
xor UO_1194 (O_1194,N_49451,N_49995);
and UO_1195 (O_1195,N_49496,N_49732);
nor UO_1196 (O_1196,N_49360,N_49440);
and UO_1197 (O_1197,N_49211,N_49317);
nand UO_1198 (O_1198,N_49102,N_49128);
nand UO_1199 (O_1199,N_49323,N_49306);
nor UO_1200 (O_1200,N_49615,N_49393);
and UO_1201 (O_1201,N_49928,N_49908);
nor UO_1202 (O_1202,N_49483,N_49947);
xor UO_1203 (O_1203,N_49893,N_49022);
nor UO_1204 (O_1204,N_49110,N_49654);
xnor UO_1205 (O_1205,N_49048,N_49230);
xnor UO_1206 (O_1206,N_49528,N_49647);
and UO_1207 (O_1207,N_49483,N_49452);
or UO_1208 (O_1208,N_49013,N_49343);
and UO_1209 (O_1209,N_49644,N_49953);
nor UO_1210 (O_1210,N_49959,N_49182);
nand UO_1211 (O_1211,N_49704,N_49911);
and UO_1212 (O_1212,N_49431,N_49433);
xor UO_1213 (O_1213,N_49742,N_49082);
xor UO_1214 (O_1214,N_49769,N_49379);
xor UO_1215 (O_1215,N_49711,N_49490);
nor UO_1216 (O_1216,N_49853,N_49406);
or UO_1217 (O_1217,N_49746,N_49452);
or UO_1218 (O_1218,N_49056,N_49777);
nand UO_1219 (O_1219,N_49339,N_49144);
nor UO_1220 (O_1220,N_49046,N_49446);
nor UO_1221 (O_1221,N_49975,N_49279);
or UO_1222 (O_1222,N_49664,N_49330);
or UO_1223 (O_1223,N_49904,N_49281);
nand UO_1224 (O_1224,N_49619,N_49447);
and UO_1225 (O_1225,N_49532,N_49981);
or UO_1226 (O_1226,N_49516,N_49148);
nor UO_1227 (O_1227,N_49053,N_49365);
nand UO_1228 (O_1228,N_49469,N_49195);
xor UO_1229 (O_1229,N_49746,N_49741);
and UO_1230 (O_1230,N_49212,N_49927);
nor UO_1231 (O_1231,N_49299,N_49580);
or UO_1232 (O_1232,N_49381,N_49241);
and UO_1233 (O_1233,N_49022,N_49161);
nand UO_1234 (O_1234,N_49774,N_49787);
xnor UO_1235 (O_1235,N_49649,N_49293);
nand UO_1236 (O_1236,N_49814,N_49570);
and UO_1237 (O_1237,N_49834,N_49868);
nand UO_1238 (O_1238,N_49994,N_49881);
and UO_1239 (O_1239,N_49191,N_49479);
nand UO_1240 (O_1240,N_49922,N_49800);
nand UO_1241 (O_1241,N_49342,N_49642);
nor UO_1242 (O_1242,N_49044,N_49090);
nand UO_1243 (O_1243,N_49845,N_49350);
xnor UO_1244 (O_1244,N_49832,N_49928);
and UO_1245 (O_1245,N_49685,N_49386);
nor UO_1246 (O_1246,N_49630,N_49499);
xor UO_1247 (O_1247,N_49514,N_49149);
or UO_1248 (O_1248,N_49211,N_49084);
and UO_1249 (O_1249,N_49612,N_49243);
or UO_1250 (O_1250,N_49139,N_49006);
or UO_1251 (O_1251,N_49302,N_49606);
nor UO_1252 (O_1252,N_49654,N_49200);
nand UO_1253 (O_1253,N_49149,N_49659);
nand UO_1254 (O_1254,N_49125,N_49117);
nor UO_1255 (O_1255,N_49579,N_49954);
xor UO_1256 (O_1256,N_49007,N_49535);
or UO_1257 (O_1257,N_49512,N_49485);
xnor UO_1258 (O_1258,N_49421,N_49126);
and UO_1259 (O_1259,N_49037,N_49428);
xnor UO_1260 (O_1260,N_49849,N_49203);
and UO_1261 (O_1261,N_49896,N_49120);
nand UO_1262 (O_1262,N_49639,N_49129);
xnor UO_1263 (O_1263,N_49417,N_49185);
nand UO_1264 (O_1264,N_49733,N_49428);
or UO_1265 (O_1265,N_49264,N_49267);
nor UO_1266 (O_1266,N_49425,N_49243);
nand UO_1267 (O_1267,N_49985,N_49904);
xor UO_1268 (O_1268,N_49270,N_49927);
xnor UO_1269 (O_1269,N_49245,N_49141);
nor UO_1270 (O_1270,N_49149,N_49051);
or UO_1271 (O_1271,N_49421,N_49975);
xnor UO_1272 (O_1272,N_49749,N_49060);
and UO_1273 (O_1273,N_49354,N_49591);
nor UO_1274 (O_1274,N_49675,N_49706);
nand UO_1275 (O_1275,N_49126,N_49855);
and UO_1276 (O_1276,N_49574,N_49230);
xnor UO_1277 (O_1277,N_49473,N_49158);
or UO_1278 (O_1278,N_49749,N_49433);
nand UO_1279 (O_1279,N_49699,N_49453);
nand UO_1280 (O_1280,N_49183,N_49180);
xor UO_1281 (O_1281,N_49924,N_49562);
xor UO_1282 (O_1282,N_49040,N_49452);
nor UO_1283 (O_1283,N_49864,N_49723);
and UO_1284 (O_1284,N_49934,N_49091);
or UO_1285 (O_1285,N_49566,N_49793);
nor UO_1286 (O_1286,N_49281,N_49258);
xnor UO_1287 (O_1287,N_49875,N_49769);
nand UO_1288 (O_1288,N_49415,N_49371);
and UO_1289 (O_1289,N_49024,N_49949);
or UO_1290 (O_1290,N_49088,N_49902);
nand UO_1291 (O_1291,N_49987,N_49354);
or UO_1292 (O_1292,N_49733,N_49666);
and UO_1293 (O_1293,N_49927,N_49352);
and UO_1294 (O_1294,N_49709,N_49707);
and UO_1295 (O_1295,N_49105,N_49370);
nand UO_1296 (O_1296,N_49855,N_49859);
or UO_1297 (O_1297,N_49719,N_49246);
and UO_1298 (O_1298,N_49562,N_49642);
xnor UO_1299 (O_1299,N_49679,N_49572);
and UO_1300 (O_1300,N_49596,N_49515);
nor UO_1301 (O_1301,N_49479,N_49098);
xor UO_1302 (O_1302,N_49962,N_49454);
nor UO_1303 (O_1303,N_49041,N_49071);
and UO_1304 (O_1304,N_49816,N_49790);
and UO_1305 (O_1305,N_49581,N_49746);
and UO_1306 (O_1306,N_49346,N_49455);
or UO_1307 (O_1307,N_49253,N_49399);
or UO_1308 (O_1308,N_49513,N_49657);
nor UO_1309 (O_1309,N_49382,N_49695);
nand UO_1310 (O_1310,N_49646,N_49583);
nand UO_1311 (O_1311,N_49364,N_49162);
or UO_1312 (O_1312,N_49003,N_49818);
nor UO_1313 (O_1313,N_49866,N_49586);
and UO_1314 (O_1314,N_49788,N_49856);
xor UO_1315 (O_1315,N_49550,N_49055);
xnor UO_1316 (O_1316,N_49926,N_49321);
nor UO_1317 (O_1317,N_49075,N_49271);
and UO_1318 (O_1318,N_49483,N_49968);
and UO_1319 (O_1319,N_49870,N_49035);
nor UO_1320 (O_1320,N_49962,N_49832);
nand UO_1321 (O_1321,N_49426,N_49838);
nand UO_1322 (O_1322,N_49645,N_49306);
and UO_1323 (O_1323,N_49466,N_49398);
xor UO_1324 (O_1324,N_49022,N_49919);
nor UO_1325 (O_1325,N_49587,N_49941);
xor UO_1326 (O_1326,N_49684,N_49136);
xnor UO_1327 (O_1327,N_49465,N_49585);
xor UO_1328 (O_1328,N_49499,N_49801);
nand UO_1329 (O_1329,N_49138,N_49004);
nand UO_1330 (O_1330,N_49087,N_49968);
and UO_1331 (O_1331,N_49215,N_49127);
nor UO_1332 (O_1332,N_49322,N_49598);
nand UO_1333 (O_1333,N_49387,N_49128);
nand UO_1334 (O_1334,N_49472,N_49389);
nor UO_1335 (O_1335,N_49454,N_49083);
and UO_1336 (O_1336,N_49232,N_49668);
and UO_1337 (O_1337,N_49151,N_49447);
nor UO_1338 (O_1338,N_49194,N_49133);
nand UO_1339 (O_1339,N_49594,N_49979);
or UO_1340 (O_1340,N_49261,N_49732);
and UO_1341 (O_1341,N_49258,N_49765);
nand UO_1342 (O_1342,N_49219,N_49289);
xor UO_1343 (O_1343,N_49798,N_49172);
xor UO_1344 (O_1344,N_49640,N_49314);
nand UO_1345 (O_1345,N_49467,N_49560);
nor UO_1346 (O_1346,N_49307,N_49867);
nand UO_1347 (O_1347,N_49587,N_49316);
xor UO_1348 (O_1348,N_49313,N_49492);
nand UO_1349 (O_1349,N_49041,N_49350);
or UO_1350 (O_1350,N_49687,N_49122);
nor UO_1351 (O_1351,N_49687,N_49751);
nor UO_1352 (O_1352,N_49328,N_49185);
nor UO_1353 (O_1353,N_49077,N_49967);
nor UO_1354 (O_1354,N_49127,N_49178);
and UO_1355 (O_1355,N_49766,N_49147);
or UO_1356 (O_1356,N_49172,N_49852);
nand UO_1357 (O_1357,N_49455,N_49459);
xor UO_1358 (O_1358,N_49262,N_49208);
nand UO_1359 (O_1359,N_49047,N_49359);
and UO_1360 (O_1360,N_49577,N_49333);
and UO_1361 (O_1361,N_49866,N_49985);
nor UO_1362 (O_1362,N_49327,N_49705);
nor UO_1363 (O_1363,N_49509,N_49611);
nor UO_1364 (O_1364,N_49185,N_49459);
and UO_1365 (O_1365,N_49228,N_49698);
nor UO_1366 (O_1366,N_49706,N_49761);
nand UO_1367 (O_1367,N_49839,N_49051);
or UO_1368 (O_1368,N_49201,N_49500);
nand UO_1369 (O_1369,N_49527,N_49879);
or UO_1370 (O_1370,N_49164,N_49646);
nor UO_1371 (O_1371,N_49925,N_49053);
nor UO_1372 (O_1372,N_49067,N_49549);
xnor UO_1373 (O_1373,N_49458,N_49085);
nor UO_1374 (O_1374,N_49494,N_49968);
and UO_1375 (O_1375,N_49109,N_49246);
or UO_1376 (O_1376,N_49419,N_49535);
or UO_1377 (O_1377,N_49225,N_49754);
and UO_1378 (O_1378,N_49858,N_49444);
and UO_1379 (O_1379,N_49517,N_49929);
nor UO_1380 (O_1380,N_49030,N_49188);
nor UO_1381 (O_1381,N_49677,N_49253);
nand UO_1382 (O_1382,N_49392,N_49714);
nor UO_1383 (O_1383,N_49003,N_49472);
nor UO_1384 (O_1384,N_49678,N_49360);
nand UO_1385 (O_1385,N_49598,N_49908);
xnor UO_1386 (O_1386,N_49437,N_49875);
nor UO_1387 (O_1387,N_49161,N_49680);
or UO_1388 (O_1388,N_49696,N_49389);
nand UO_1389 (O_1389,N_49409,N_49173);
and UO_1390 (O_1390,N_49107,N_49813);
or UO_1391 (O_1391,N_49590,N_49543);
xor UO_1392 (O_1392,N_49521,N_49862);
or UO_1393 (O_1393,N_49778,N_49578);
xnor UO_1394 (O_1394,N_49880,N_49957);
or UO_1395 (O_1395,N_49209,N_49197);
nor UO_1396 (O_1396,N_49628,N_49414);
nor UO_1397 (O_1397,N_49656,N_49306);
or UO_1398 (O_1398,N_49123,N_49709);
and UO_1399 (O_1399,N_49547,N_49531);
and UO_1400 (O_1400,N_49011,N_49641);
or UO_1401 (O_1401,N_49939,N_49009);
nand UO_1402 (O_1402,N_49131,N_49560);
or UO_1403 (O_1403,N_49727,N_49692);
and UO_1404 (O_1404,N_49203,N_49877);
and UO_1405 (O_1405,N_49780,N_49465);
xnor UO_1406 (O_1406,N_49809,N_49377);
and UO_1407 (O_1407,N_49760,N_49944);
and UO_1408 (O_1408,N_49281,N_49421);
xnor UO_1409 (O_1409,N_49015,N_49107);
nor UO_1410 (O_1410,N_49274,N_49409);
nor UO_1411 (O_1411,N_49666,N_49598);
nand UO_1412 (O_1412,N_49097,N_49034);
xor UO_1413 (O_1413,N_49040,N_49583);
and UO_1414 (O_1414,N_49402,N_49759);
xnor UO_1415 (O_1415,N_49212,N_49988);
and UO_1416 (O_1416,N_49434,N_49063);
xor UO_1417 (O_1417,N_49588,N_49156);
and UO_1418 (O_1418,N_49497,N_49612);
and UO_1419 (O_1419,N_49904,N_49457);
nor UO_1420 (O_1420,N_49625,N_49938);
xor UO_1421 (O_1421,N_49833,N_49900);
xor UO_1422 (O_1422,N_49683,N_49939);
and UO_1423 (O_1423,N_49972,N_49721);
and UO_1424 (O_1424,N_49581,N_49189);
and UO_1425 (O_1425,N_49567,N_49400);
nand UO_1426 (O_1426,N_49949,N_49635);
and UO_1427 (O_1427,N_49659,N_49343);
and UO_1428 (O_1428,N_49757,N_49529);
and UO_1429 (O_1429,N_49250,N_49681);
nand UO_1430 (O_1430,N_49384,N_49843);
xor UO_1431 (O_1431,N_49383,N_49087);
xnor UO_1432 (O_1432,N_49508,N_49718);
or UO_1433 (O_1433,N_49434,N_49326);
and UO_1434 (O_1434,N_49249,N_49822);
nor UO_1435 (O_1435,N_49247,N_49229);
nor UO_1436 (O_1436,N_49784,N_49933);
nand UO_1437 (O_1437,N_49615,N_49224);
xor UO_1438 (O_1438,N_49067,N_49258);
or UO_1439 (O_1439,N_49479,N_49523);
and UO_1440 (O_1440,N_49533,N_49027);
nor UO_1441 (O_1441,N_49513,N_49795);
nor UO_1442 (O_1442,N_49814,N_49579);
or UO_1443 (O_1443,N_49948,N_49196);
and UO_1444 (O_1444,N_49600,N_49422);
or UO_1445 (O_1445,N_49746,N_49781);
and UO_1446 (O_1446,N_49484,N_49704);
nand UO_1447 (O_1447,N_49414,N_49596);
nand UO_1448 (O_1448,N_49521,N_49190);
nand UO_1449 (O_1449,N_49900,N_49818);
nand UO_1450 (O_1450,N_49809,N_49215);
and UO_1451 (O_1451,N_49019,N_49264);
xor UO_1452 (O_1452,N_49956,N_49372);
and UO_1453 (O_1453,N_49919,N_49467);
and UO_1454 (O_1454,N_49152,N_49939);
nor UO_1455 (O_1455,N_49540,N_49234);
xor UO_1456 (O_1456,N_49180,N_49334);
nand UO_1457 (O_1457,N_49744,N_49103);
nand UO_1458 (O_1458,N_49194,N_49349);
and UO_1459 (O_1459,N_49329,N_49265);
and UO_1460 (O_1460,N_49919,N_49543);
nand UO_1461 (O_1461,N_49497,N_49614);
and UO_1462 (O_1462,N_49978,N_49604);
xnor UO_1463 (O_1463,N_49710,N_49022);
xnor UO_1464 (O_1464,N_49309,N_49936);
nand UO_1465 (O_1465,N_49180,N_49473);
or UO_1466 (O_1466,N_49306,N_49559);
nand UO_1467 (O_1467,N_49437,N_49083);
nor UO_1468 (O_1468,N_49208,N_49972);
or UO_1469 (O_1469,N_49504,N_49020);
or UO_1470 (O_1470,N_49068,N_49304);
nand UO_1471 (O_1471,N_49085,N_49023);
nand UO_1472 (O_1472,N_49367,N_49350);
xor UO_1473 (O_1473,N_49594,N_49812);
xnor UO_1474 (O_1474,N_49625,N_49479);
nand UO_1475 (O_1475,N_49782,N_49385);
xnor UO_1476 (O_1476,N_49145,N_49310);
nand UO_1477 (O_1477,N_49787,N_49002);
and UO_1478 (O_1478,N_49887,N_49484);
nand UO_1479 (O_1479,N_49288,N_49558);
xor UO_1480 (O_1480,N_49396,N_49794);
xor UO_1481 (O_1481,N_49852,N_49558);
nor UO_1482 (O_1482,N_49806,N_49859);
xnor UO_1483 (O_1483,N_49153,N_49452);
and UO_1484 (O_1484,N_49333,N_49314);
nor UO_1485 (O_1485,N_49937,N_49278);
or UO_1486 (O_1486,N_49962,N_49789);
or UO_1487 (O_1487,N_49288,N_49722);
xor UO_1488 (O_1488,N_49089,N_49740);
xnor UO_1489 (O_1489,N_49287,N_49025);
nand UO_1490 (O_1490,N_49026,N_49357);
or UO_1491 (O_1491,N_49223,N_49345);
nor UO_1492 (O_1492,N_49598,N_49361);
or UO_1493 (O_1493,N_49192,N_49784);
and UO_1494 (O_1494,N_49284,N_49095);
xnor UO_1495 (O_1495,N_49803,N_49027);
xor UO_1496 (O_1496,N_49472,N_49483);
nor UO_1497 (O_1497,N_49395,N_49118);
and UO_1498 (O_1498,N_49922,N_49630);
or UO_1499 (O_1499,N_49064,N_49379);
nand UO_1500 (O_1500,N_49108,N_49392);
or UO_1501 (O_1501,N_49496,N_49634);
and UO_1502 (O_1502,N_49120,N_49254);
nor UO_1503 (O_1503,N_49635,N_49851);
nor UO_1504 (O_1504,N_49134,N_49333);
and UO_1505 (O_1505,N_49902,N_49196);
or UO_1506 (O_1506,N_49776,N_49761);
nand UO_1507 (O_1507,N_49172,N_49880);
or UO_1508 (O_1508,N_49897,N_49875);
and UO_1509 (O_1509,N_49230,N_49837);
nor UO_1510 (O_1510,N_49857,N_49391);
nor UO_1511 (O_1511,N_49911,N_49211);
xnor UO_1512 (O_1512,N_49346,N_49480);
xor UO_1513 (O_1513,N_49132,N_49579);
or UO_1514 (O_1514,N_49754,N_49868);
xor UO_1515 (O_1515,N_49924,N_49035);
or UO_1516 (O_1516,N_49758,N_49965);
xor UO_1517 (O_1517,N_49497,N_49809);
or UO_1518 (O_1518,N_49144,N_49192);
nand UO_1519 (O_1519,N_49486,N_49838);
nand UO_1520 (O_1520,N_49660,N_49741);
nor UO_1521 (O_1521,N_49069,N_49804);
and UO_1522 (O_1522,N_49182,N_49735);
or UO_1523 (O_1523,N_49793,N_49391);
and UO_1524 (O_1524,N_49050,N_49853);
and UO_1525 (O_1525,N_49353,N_49851);
xor UO_1526 (O_1526,N_49031,N_49711);
or UO_1527 (O_1527,N_49808,N_49391);
xnor UO_1528 (O_1528,N_49386,N_49850);
nand UO_1529 (O_1529,N_49328,N_49184);
nor UO_1530 (O_1530,N_49110,N_49941);
nand UO_1531 (O_1531,N_49167,N_49049);
and UO_1532 (O_1532,N_49125,N_49079);
or UO_1533 (O_1533,N_49834,N_49163);
or UO_1534 (O_1534,N_49835,N_49953);
nor UO_1535 (O_1535,N_49630,N_49286);
and UO_1536 (O_1536,N_49549,N_49571);
nor UO_1537 (O_1537,N_49231,N_49668);
nand UO_1538 (O_1538,N_49347,N_49486);
and UO_1539 (O_1539,N_49566,N_49053);
nor UO_1540 (O_1540,N_49627,N_49555);
or UO_1541 (O_1541,N_49862,N_49069);
or UO_1542 (O_1542,N_49899,N_49657);
and UO_1543 (O_1543,N_49644,N_49450);
xor UO_1544 (O_1544,N_49787,N_49181);
xor UO_1545 (O_1545,N_49321,N_49180);
xor UO_1546 (O_1546,N_49099,N_49068);
nand UO_1547 (O_1547,N_49599,N_49615);
and UO_1548 (O_1548,N_49115,N_49685);
and UO_1549 (O_1549,N_49856,N_49100);
or UO_1550 (O_1550,N_49169,N_49987);
nor UO_1551 (O_1551,N_49201,N_49709);
or UO_1552 (O_1552,N_49880,N_49259);
nor UO_1553 (O_1553,N_49433,N_49545);
xor UO_1554 (O_1554,N_49305,N_49679);
nand UO_1555 (O_1555,N_49291,N_49617);
nor UO_1556 (O_1556,N_49225,N_49282);
nand UO_1557 (O_1557,N_49259,N_49675);
nand UO_1558 (O_1558,N_49486,N_49296);
nand UO_1559 (O_1559,N_49813,N_49665);
nand UO_1560 (O_1560,N_49854,N_49428);
and UO_1561 (O_1561,N_49799,N_49777);
and UO_1562 (O_1562,N_49546,N_49803);
and UO_1563 (O_1563,N_49258,N_49568);
nor UO_1564 (O_1564,N_49975,N_49284);
nor UO_1565 (O_1565,N_49695,N_49098);
nand UO_1566 (O_1566,N_49452,N_49771);
nand UO_1567 (O_1567,N_49178,N_49325);
and UO_1568 (O_1568,N_49680,N_49473);
nand UO_1569 (O_1569,N_49535,N_49715);
nor UO_1570 (O_1570,N_49247,N_49174);
nor UO_1571 (O_1571,N_49097,N_49730);
nor UO_1572 (O_1572,N_49868,N_49705);
xnor UO_1573 (O_1573,N_49945,N_49495);
xor UO_1574 (O_1574,N_49349,N_49735);
and UO_1575 (O_1575,N_49456,N_49897);
xor UO_1576 (O_1576,N_49287,N_49501);
nand UO_1577 (O_1577,N_49875,N_49878);
or UO_1578 (O_1578,N_49696,N_49592);
and UO_1579 (O_1579,N_49430,N_49948);
nor UO_1580 (O_1580,N_49504,N_49470);
nor UO_1581 (O_1581,N_49202,N_49639);
nor UO_1582 (O_1582,N_49763,N_49817);
or UO_1583 (O_1583,N_49029,N_49659);
nor UO_1584 (O_1584,N_49528,N_49108);
or UO_1585 (O_1585,N_49693,N_49121);
nand UO_1586 (O_1586,N_49530,N_49638);
nand UO_1587 (O_1587,N_49726,N_49290);
nor UO_1588 (O_1588,N_49717,N_49440);
nand UO_1589 (O_1589,N_49803,N_49732);
and UO_1590 (O_1590,N_49326,N_49844);
or UO_1591 (O_1591,N_49366,N_49139);
xnor UO_1592 (O_1592,N_49712,N_49833);
or UO_1593 (O_1593,N_49948,N_49966);
xnor UO_1594 (O_1594,N_49447,N_49120);
xnor UO_1595 (O_1595,N_49997,N_49634);
xor UO_1596 (O_1596,N_49789,N_49234);
or UO_1597 (O_1597,N_49879,N_49798);
nor UO_1598 (O_1598,N_49844,N_49537);
nand UO_1599 (O_1599,N_49745,N_49794);
nand UO_1600 (O_1600,N_49662,N_49081);
xnor UO_1601 (O_1601,N_49012,N_49183);
nor UO_1602 (O_1602,N_49721,N_49284);
or UO_1603 (O_1603,N_49611,N_49831);
xor UO_1604 (O_1604,N_49233,N_49911);
nor UO_1605 (O_1605,N_49335,N_49283);
and UO_1606 (O_1606,N_49706,N_49461);
nand UO_1607 (O_1607,N_49412,N_49224);
and UO_1608 (O_1608,N_49543,N_49588);
and UO_1609 (O_1609,N_49341,N_49735);
nor UO_1610 (O_1610,N_49238,N_49474);
xnor UO_1611 (O_1611,N_49806,N_49652);
nand UO_1612 (O_1612,N_49208,N_49384);
or UO_1613 (O_1613,N_49047,N_49390);
nand UO_1614 (O_1614,N_49135,N_49780);
or UO_1615 (O_1615,N_49117,N_49535);
and UO_1616 (O_1616,N_49678,N_49722);
or UO_1617 (O_1617,N_49772,N_49576);
and UO_1618 (O_1618,N_49122,N_49555);
nand UO_1619 (O_1619,N_49228,N_49442);
or UO_1620 (O_1620,N_49387,N_49997);
nand UO_1621 (O_1621,N_49726,N_49810);
nand UO_1622 (O_1622,N_49244,N_49699);
and UO_1623 (O_1623,N_49792,N_49672);
and UO_1624 (O_1624,N_49998,N_49934);
nand UO_1625 (O_1625,N_49520,N_49792);
or UO_1626 (O_1626,N_49040,N_49788);
and UO_1627 (O_1627,N_49245,N_49397);
and UO_1628 (O_1628,N_49730,N_49983);
nor UO_1629 (O_1629,N_49632,N_49331);
xnor UO_1630 (O_1630,N_49629,N_49402);
nand UO_1631 (O_1631,N_49370,N_49234);
and UO_1632 (O_1632,N_49784,N_49456);
nand UO_1633 (O_1633,N_49998,N_49751);
nor UO_1634 (O_1634,N_49496,N_49796);
and UO_1635 (O_1635,N_49386,N_49710);
nor UO_1636 (O_1636,N_49351,N_49747);
nor UO_1637 (O_1637,N_49512,N_49739);
or UO_1638 (O_1638,N_49993,N_49694);
or UO_1639 (O_1639,N_49391,N_49824);
nand UO_1640 (O_1640,N_49325,N_49245);
and UO_1641 (O_1641,N_49324,N_49615);
nand UO_1642 (O_1642,N_49502,N_49170);
or UO_1643 (O_1643,N_49480,N_49711);
nand UO_1644 (O_1644,N_49344,N_49867);
and UO_1645 (O_1645,N_49002,N_49049);
xnor UO_1646 (O_1646,N_49951,N_49675);
xnor UO_1647 (O_1647,N_49825,N_49411);
nor UO_1648 (O_1648,N_49897,N_49470);
nor UO_1649 (O_1649,N_49206,N_49398);
or UO_1650 (O_1650,N_49756,N_49503);
nand UO_1651 (O_1651,N_49021,N_49338);
or UO_1652 (O_1652,N_49033,N_49618);
nor UO_1653 (O_1653,N_49484,N_49169);
nand UO_1654 (O_1654,N_49504,N_49331);
xnor UO_1655 (O_1655,N_49396,N_49361);
and UO_1656 (O_1656,N_49590,N_49366);
xnor UO_1657 (O_1657,N_49412,N_49352);
and UO_1658 (O_1658,N_49114,N_49709);
xor UO_1659 (O_1659,N_49288,N_49673);
or UO_1660 (O_1660,N_49247,N_49688);
nor UO_1661 (O_1661,N_49762,N_49868);
nand UO_1662 (O_1662,N_49902,N_49276);
nand UO_1663 (O_1663,N_49059,N_49534);
xor UO_1664 (O_1664,N_49233,N_49590);
and UO_1665 (O_1665,N_49596,N_49938);
nor UO_1666 (O_1666,N_49246,N_49645);
nor UO_1667 (O_1667,N_49726,N_49558);
or UO_1668 (O_1668,N_49809,N_49767);
nand UO_1669 (O_1669,N_49272,N_49452);
xnor UO_1670 (O_1670,N_49820,N_49975);
nand UO_1671 (O_1671,N_49580,N_49517);
and UO_1672 (O_1672,N_49687,N_49283);
nor UO_1673 (O_1673,N_49676,N_49271);
nand UO_1674 (O_1674,N_49505,N_49539);
and UO_1675 (O_1675,N_49449,N_49620);
nand UO_1676 (O_1676,N_49508,N_49298);
nor UO_1677 (O_1677,N_49735,N_49068);
and UO_1678 (O_1678,N_49499,N_49320);
and UO_1679 (O_1679,N_49457,N_49791);
nand UO_1680 (O_1680,N_49445,N_49489);
nand UO_1681 (O_1681,N_49949,N_49239);
and UO_1682 (O_1682,N_49927,N_49433);
nor UO_1683 (O_1683,N_49828,N_49799);
xnor UO_1684 (O_1684,N_49317,N_49885);
xor UO_1685 (O_1685,N_49852,N_49567);
nand UO_1686 (O_1686,N_49053,N_49881);
or UO_1687 (O_1687,N_49142,N_49734);
nor UO_1688 (O_1688,N_49412,N_49419);
or UO_1689 (O_1689,N_49261,N_49489);
or UO_1690 (O_1690,N_49131,N_49716);
and UO_1691 (O_1691,N_49880,N_49325);
nor UO_1692 (O_1692,N_49790,N_49709);
nand UO_1693 (O_1693,N_49206,N_49755);
nand UO_1694 (O_1694,N_49641,N_49294);
xor UO_1695 (O_1695,N_49024,N_49853);
or UO_1696 (O_1696,N_49485,N_49372);
xor UO_1697 (O_1697,N_49062,N_49571);
nor UO_1698 (O_1698,N_49537,N_49327);
nor UO_1699 (O_1699,N_49178,N_49573);
nor UO_1700 (O_1700,N_49451,N_49543);
nand UO_1701 (O_1701,N_49426,N_49511);
xor UO_1702 (O_1702,N_49178,N_49828);
and UO_1703 (O_1703,N_49839,N_49092);
nand UO_1704 (O_1704,N_49946,N_49773);
nand UO_1705 (O_1705,N_49844,N_49701);
nor UO_1706 (O_1706,N_49236,N_49507);
and UO_1707 (O_1707,N_49720,N_49372);
and UO_1708 (O_1708,N_49724,N_49906);
or UO_1709 (O_1709,N_49087,N_49545);
nor UO_1710 (O_1710,N_49142,N_49038);
and UO_1711 (O_1711,N_49015,N_49023);
and UO_1712 (O_1712,N_49944,N_49691);
nor UO_1713 (O_1713,N_49682,N_49683);
and UO_1714 (O_1714,N_49585,N_49073);
and UO_1715 (O_1715,N_49585,N_49188);
and UO_1716 (O_1716,N_49747,N_49936);
or UO_1717 (O_1717,N_49265,N_49575);
and UO_1718 (O_1718,N_49130,N_49317);
or UO_1719 (O_1719,N_49016,N_49551);
xor UO_1720 (O_1720,N_49692,N_49591);
nand UO_1721 (O_1721,N_49211,N_49406);
and UO_1722 (O_1722,N_49253,N_49280);
xor UO_1723 (O_1723,N_49387,N_49428);
or UO_1724 (O_1724,N_49660,N_49886);
or UO_1725 (O_1725,N_49162,N_49203);
nand UO_1726 (O_1726,N_49370,N_49140);
xor UO_1727 (O_1727,N_49078,N_49499);
and UO_1728 (O_1728,N_49946,N_49446);
nor UO_1729 (O_1729,N_49498,N_49288);
nor UO_1730 (O_1730,N_49227,N_49695);
nor UO_1731 (O_1731,N_49034,N_49969);
nand UO_1732 (O_1732,N_49911,N_49159);
and UO_1733 (O_1733,N_49286,N_49746);
xor UO_1734 (O_1734,N_49301,N_49193);
nor UO_1735 (O_1735,N_49859,N_49179);
xnor UO_1736 (O_1736,N_49181,N_49024);
nor UO_1737 (O_1737,N_49370,N_49232);
nor UO_1738 (O_1738,N_49733,N_49058);
nor UO_1739 (O_1739,N_49070,N_49725);
nor UO_1740 (O_1740,N_49323,N_49607);
or UO_1741 (O_1741,N_49852,N_49551);
or UO_1742 (O_1742,N_49034,N_49045);
xnor UO_1743 (O_1743,N_49580,N_49040);
or UO_1744 (O_1744,N_49476,N_49003);
nor UO_1745 (O_1745,N_49168,N_49877);
xor UO_1746 (O_1746,N_49088,N_49955);
and UO_1747 (O_1747,N_49454,N_49107);
or UO_1748 (O_1748,N_49386,N_49205);
or UO_1749 (O_1749,N_49322,N_49713);
nor UO_1750 (O_1750,N_49798,N_49301);
or UO_1751 (O_1751,N_49620,N_49913);
xor UO_1752 (O_1752,N_49728,N_49834);
or UO_1753 (O_1753,N_49964,N_49473);
or UO_1754 (O_1754,N_49239,N_49102);
xor UO_1755 (O_1755,N_49037,N_49996);
nand UO_1756 (O_1756,N_49664,N_49538);
nand UO_1757 (O_1757,N_49443,N_49407);
nor UO_1758 (O_1758,N_49587,N_49151);
or UO_1759 (O_1759,N_49324,N_49561);
nand UO_1760 (O_1760,N_49769,N_49313);
or UO_1761 (O_1761,N_49940,N_49592);
nor UO_1762 (O_1762,N_49152,N_49525);
and UO_1763 (O_1763,N_49971,N_49551);
nand UO_1764 (O_1764,N_49616,N_49709);
nor UO_1765 (O_1765,N_49351,N_49058);
xor UO_1766 (O_1766,N_49230,N_49304);
nor UO_1767 (O_1767,N_49296,N_49005);
nor UO_1768 (O_1768,N_49834,N_49393);
xor UO_1769 (O_1769,N_49913,N_49585);
nor UO_1770 (O_1770,N_49274,N_49820);
or UO_1771 (O_1771,N_49665,N_49336);
or UO_1772 (O_1772,N_49002,N_49043);
nor UO_1773 (O_1773,N_49371,N_49378);
or UO_1774 (O_1774,N_49875,N_49846);
and UO_1775 (O_1775,N_49461,N_49529);
and UO_1776 (O_1776,N_49891,N_49690);
and UO_1777 (O_1777,N_49989,N_49879);
and UO_1778 (O_1778,N_49065,N_49127);
nor UO_1779 (O_1779,N_49906,N_49558);
nor UO_1780 (O_1780,N_49348,N_49443);
nand UO_1781 (O_1781,N_49249,N_49208);
xnor UO_1782 (O_1782,N_49879,N_49167);
nand UO_1783 (O_1783,N_49022,N_49145);
nand UO_1784 (O_1784,N_49566,N_49118);
or UO_1785 (O_1785,N_49104,N_49292);
xnor UO_1786 (O_1786,N_49149,N_49160);
nand UO_1787 (O_1787,N_49176,N_49054);
xor UO_1788 (O_1788,N_49179,N_49378);
or UO_1789 (O_1789,N_49206,N_49351);
and UO_1790 (O_1790,N_49503,N_49285);
and UO_1791 (O_1791,N_49517,N_49032);
nor UO_1792 (O_1792,N_49288,N_49844);
nor UO_1793 (O_1793,N_49154,N_49915);
nor UO_1794 (O_1794,N_49736,N_49904);
and UO_1795 (O_1795,N_49231,N_49634);
xnor UO_1796 (O_1796,N_49879,N_49189);
xnor UO_1797 (O_1797,N_49481,N_49505);
nor UO_1798 (O_1798,N_49694,N_49566);
and UO_1799 (O_1799,N_49306,N_49908);
and UO_1800 (O_1800,N_49296,N_49148);
nor UO_1801 (O_1801,N_49480,N_49876);
nand UO_1802 (O_1802,N_49944,N_49359);
and UO_1803 (O_1803,N_49096,N_49500);
or UO_1804 (O_1804,N_49760,N_49657);
nand UO_1805 (O_1805,N_49147,N_49877);
nor UO_1806 (O_1806,N_49481,N_49312);
and UO_1807 (O_1807,N_49213,N_49625);
nor UO_1808 (O_1808,N_49540,N_49361);
or UO_1809 (O_1809,N_49366,N_49713);
nand UO_1810 (O_1810,N_49972,N_49031);
nor UO_1811 (O_1811,N_49009,N_49644);
xnor UO_1812 (O_1812,N_49610,N_49849);
nand UO_1813 (O_1813,N_49850,N_49076);
xnor UO_1814 (O_1814,N_49664,N_49511);
nor UO_1815 (O_1815,N_49808,N_49349);
nor UO_1816 (O_1816,N_49598,N_49579);
nand UO_1817 (O_1817,N_49554,N_49042);
xnor UO_1818 (O_1818,N_49384,N_49694);
nor UO_1819 (O_1819,N_49944,N_49786);
and UO_1820 (O_1820,N_49709,N_49816);
nor UO_1821 (O_1821,N_49127,N_49561);
or UO_1822 (O_1822,N_49143,N_49871);
nand UO_1823 (O_1823,N_49087,N_49917);
xor UO_1824 (O_1824,N_49187,N_49180);
or UO_1825 (O_1825,N_49124,N_49429);
nor UO_1826 (O_1826,N_49739,N_49749);
or UO_1827 (O_1827,N_49943,N_49559);
and UO_1828 (O_1828,N_49796,N_49117);
xnor UO_1829 (O_1829,N_49084,N_49795);
or UO_1830 (O_1830,N_49942,N_49940);
xnor UO_1831 (O_1831,N_49483,N_49850);
nand UO_1832 (O_1832,N_49148,N_49936);
or UO_1833 (O_1833,N_49626,N_49001);
nor UO_1834 (O_1834,N_49233,N_49296);
xor UO_1835 (O_1835,N_49540,N_49414);
and UO_1836 (O_1836,N_49678,N_49871);
and UO_1837 (O_1837,N_49447,N_49095);
xnor UO_1838 (O_1838,N_49654,N_49691);
nand UO_1839 (O_1839,N_49575,N_49249);
nand UO_1840 (O_1840,N_49059,N_49074);
xnor UO_1841 (O_1841,N_49245,N_49494);
nor UO_1842 (O_1842,N_49559,N_49242);
nor UO_1843 (O_1843,N_49833,N_49310);
xnor UO_1844 (O_1844,N_49545,N_49221);
xor UO_1845 (O_1845,N_49522,N_49793);
or UO_1846 (O_1846,N_49508,N_49637);
or UO_1847 (O_1847,N_49648,N_49106);
and UO_1848 (O_1848,N_49969,N_49256);
xor UO_1849 (O_1849,N_49091,N_49569);
nand UO_1850 (O_1850,N_49821,N_49877);
nand UO_1851 (O_1851,N_49070,N_49612);
nand UO_1852 (O_1852,N_49057,N_49369);
nand UO_1853 (O_1853,N_49795,N_49025);
xnor UO_1854 (O_1854,N_49535,N_49969);
nand UO_1855 (O_1855,N_49538,N_49094);
and UO_1856 (O_1856,N_49149,N_49796);
nand UO_1857 (O_1857,N_49103,N_49878);
and UO_1858 (O_1858,N_49200,N_49594);
nor UO_1859 (O_1859,N_49973,N_49872);
and UO_1860 (O_1860,N_49188,N_49708);
xor UO_1861 (O_1861,N_49744,N_49111);
or UO_1862 (O_1862,N_49810,N_49807);
or UO_1863 (O_1863,N_49315,N_49559);
xnor UO_1864 (O_1864,N_49919,N_49757);
nor UO_1865 (O_1865,N_49943,N_49693);
and UO_1866 (O_1866,N_49578,N_49723);
xnor UO_1867 (O_1867,N_49318,N_49989);
xnor UO_1868 (O_1868,N_49629,N_49319);
nor UO_1869 (O_1869,N_49757,N_49786);
nand UO_1870 (O_1870,N_49311,N_49892);
nand UO_1871 (O_1871,N_49719,N_49030);
nor UO_1872 (O_1872,N_49735,N_49520);
xnor UO_1873 (O_1873,N_49404,N_49869);
nand UO_1874 (O_1874,N_49114,N_49636);
xor UO_1875 (O_1875,N_49215,N_49381);
or UO_1876 (O_1876,N_49684,N_49988);
nand UO_1877 (O_1877,N_49131,N_49220);
nand UO_1878 (O_1878,N_49437,N_49613);
or UO_1879 (O_1879,N_49401,N_49159);
xnor UO_1880 (O_1880,N_49833,N_49081);
nand UO_1881 (O_1881,N_49398,N_49813);
and UO_1882 (O_1882,N_49730,N_49036);
nand UO_1883 (O_1883,N_49561,N_49383);
nand UO_1884 (O_1884,N_49818,N_49561);
nor UO_1885 (O_1885,N_49644,N_49429);
and UO_1886 (O_1886,N_49466,N_49149);
and UO_1887 (O_1887,N_49474,N_49561);
and UO_1888 (O_1888,N_49752,N_49027);
and UO_1889 (O_1889,N_49214,N_49816);
xor UO_1890 (O_1890,N_49217,N_49412);
nand UO_1891 (O_1891,N_49904,N_49078);
xnor UO_1892 (O_1892,N_49596,N_49588);
xnor UO_1893 (O_1893,N_49250,N_49991);
xor UO_1894 (O_1894,N_49788,N_49270);
or UO_1895 (O_1895,N_49462,N_49556);
and UO_1896 (O_1896,N_49083,N_49985);
nand UO_1897 (O_1897,N_49179,N_49918);
nand UO_1898 (O_1898,N_49473,N_49668);
and UO_1899 (O_1899,N_49972,N_49598);
nand UO_1900 (O_1900,N_49272,N_49526);
xnor UO_1901 (O_1901,N_49383,N_49423);
and UO_1902 (O_1902,N_49103,N_49238);
or UO_1903 (O_1903,N_49034,N_49141);
nor UO_1904 (O_1904,N_49299,N_49751);
and UO_1905 (O_1905,N_49322,N_49772);
nor UO_1906 (O_1906,N_49243,N_49620);
nor UO_1907 (O_1907,N_49033,N_49822);
xor UO_1908 (O_1908,N_49053,N_49006);
xnor UO_1909 (O_1909,N_49021,N_49027);
nand UO_1910 (O_1910,N_49540,N_49826);
and UO_1911 (O_1911,N_49118,N_49599);
nor UO_1912 (O_1912,N_49119,N_49488);
nand UO_1913 (O_1913,N_49594,N_49093);
or UO_1914 (O_1914,N_49685,N_49970);
or UO_1915 (O_1915,N_49236,N_49866);
and UO_1916 (O_1916,N_49546,N_49557);
nor UO_1917 (O_1917,N_49684,N_49724);
nor UO_1918 (O_1918,N_49979,N_49459);
nand UO_1919 (O_1919,N_49659,N_49189);
nand UO_1920 (O_1920,N_49687,N_49047);
and UO_1921 (O_1921,N_49410,N_49834);
and UO_1922 (O_1922,N_49308,N_49456);
xnor UO_1923 (O_1923,N_49127,N_49758);
or UO_1924 (O_1924,N_49696,N_49394);
and UO_1925 (O_1925,N_49867,N_49800);
nand UO_1926 (O_1926,N_49234,N_49458);
xor UO_1927 (O_1927,N_49107,N_49946);
nand UO_1928 (O_1928,N_49489,N_49251);
nand UO_1929 (O_1929,N_49752,N_49212);
nand UO_1930 (O_1930,N_49989,N_49719);
or UO_1931 (O_1931,N_49580,N_49270);
nand UO_1932 (O_1932,N_49173,N_49931);
nor UO_1933 (O_1933,N_49641,N_49779);
and UO_1934 (O_1934,N_49476,N_49589);
nand UO_1935 (O_1935,N_49275,N_49052);
and UO_1936 (O_1936,N_49871,N_49550);
or UO_1937 (O_1937,N_49717,N_49793);
xor UO_1938 (O_1938,N_49058,N_49310);
and UO_1939 (O_1939,N_49803,N_49553);
or UO_1940 (O_1940,N_49227,N_49489);
nor UO_1941 (O_1941,N_49882,N_49459);
or UO_1942 (O_1942,N_49897,N_49465);
and UO_1943 (O_1943,N_49891,N_49590);
nand UO_1944 (O_1944,N_49425,N_49568);
and UO_1945 (O_1945,N_49871,N_49789);
xor UO_1946 (O_1946,N_49554,N_49594);
nor UO_1947 (O_1947,N_49662,N_49102);
nor UO_1948 (O_1948,N_49745,N_49968);
or UO_1949 (O_1949,N_49482,N_49676);
xnor UO_1950 (O_1950,N_49365,N_49445);
xor UO_1951 (O_1951,N_49951,N_49336);
nand UO_1952 (O_1952,N_49228,N_49569);
xor UO_1953 (O_1953,N_49176,N_49779);
nand UO_1954 (O_1954,N_49275,N_49521);
nand UO_1955 (O_1955,N_49721,N_49032);
xnor UO_1956 (O_1956,N_49613,N_49212);
and UO_1957 (O_1957,N_49722,N_49263);
nor UO_1958 (O_1958,N_49231,N_49963);
xor UO_1959 (O_1959,N_49161,N_49422);
and UO_1960 (O_1960,N_49630,N_49118);
nor UO_1961 (O_1961,N_49839,N_49033);
nor UO_1962 (O_1962,N_49568,N_49806);
xnor UO_1963 (O_1963,N_49782,N_49303);
nor UO_1964 (O_1964,N_49211,N_49501);
or UO_1965 (O_1965,N_49681,N_49402);
and UO_1966 (O_1966,N_49442,N_49550);
or UO_1967 (O_1967,N_49750,N_49368);
xor UO_1968 (O_1968,N_49436,N_49705);
xor UO_1969 (O_1969,N_49653,N_49420);
nor UO_1970 (O_1970,N_49758,N_49491);
nand UO_1971 (O_1971,N_49507,N_49813);
xor UO_1972 (O_1972,N_49763,N_49180);
nand UO_1973 (O_1973,N_49953,N_49889);
nor UO_1974 (O_1974,N_49272,N_49360);
nand UO_1975 (O_1975,N_49441,N_49317);
nor UO_1976 (O_1976,N_49041,N_49287);
and UO_1977 (O_1977,N_49850,N_49455);
or UO_1978 (O_1978,N_49869,N_49296);
and UO_1979 (O_1979,N_49889,N_49580);
and UO_1980 (O_1980,N_49234,N_49143);
or UO_1981 (O_1981,N_49355,N_49826);
or UO_1982 (O_1982,N_49834,N_49014);
and UO_1983 (O_1983,N_49489,N_49236);
nor UO_1984 (O_1984,N_49502,N_49462);
nand UO_1985 (O_1985,N_49903,N_49366);
or UO_1986 (O_1986,N_49315,N_49095);
or UO_1987 (O_1987,N_49312,N_49175);
xnor UO_1988 (O_1988,N_49664,N_49603);
nor UO_1989 (O_1989,N_49733,N_49933);
or UO_1990 (O_1990,N_49994,N_49463);
or UO_1991 (O_1991,N_49038,N_49093);
or UO_1992 (O_1992,N_49367,N_49508);
and UO_1993 (O_1993,N_49342,N_49027);
nor UO_1994 (O_1994,N_49024,N_49406);
xnor UO_1995 (O_1995,N_49855,N_49722);
and UO_1996 (O_1996,N_49087,N_49884);
nand UO_1997 (O_1997,N_49070,N_49734);
nor UO_1998 (O_1998,N_49827,N_49090);
xor UO_1999 (O_1999,N_49829,N_49360);
xor UO_2000 (O_2000,N_49029,N_49847);
and UO_2001 (O_2001,N_49866,N_49426);
or UO_2002 (O_2002,N_49697,N_49540);
nand UO_2003 (O_2003,N_49759,N_49262);
xor UO_2004 (O_2004,N_49442,N_49532);
and UO_2005 (O_2005,N_49867,N_49259);
and UO_2006 (O_2006,N_49931,N_49340);
or UO_2007 (O_2007,N_49851,N_49179);
or UO_2008 (O_2008,N_49907,N_49758);
or UO_2009 (O_2009,N_49698,N_49651);
nor UO_2010 (O_2010,N_49504,N_49324);
nand UO_2011 (O_2011,N_49359,N_49162);
nor UO_2012 (O_2012,N_49235,N_49247);
and UO_2013 (O_2013,N_49861,N_49227);
nor UO_2014 (O_2014,N_49032,N_49209);
nand UO_2015 (O_2015,N_49380,N_49096);
xnor UO_2016 (O_2016,N_49987,N_49131);
nor UO_2017 (O_2017,N_49837,N_49197);
or UO_2018 (O_2018,N_49295,N_49948);
nor UO_2019 (O_2019,N_49607,N_49871);
nor UO_2020 (O_2020,N_49805,N_49399);
nor UO_2021 (O_2021,N_49446,N_49401);
or UO_2022 (O_2022,N_49194,N_49957);
nand UO_2023 (O_2023,N_49310,N_49798);
nor UO_2024 (O_2024,N_49508,N_49831);
or UO_2025 (O_2025,N_49136,N_49293);
nor UO_2026 (O_2026,N_49559,N_49252);
nor UO_2027 (O_2027,N_49121,N_49864);
nor UO_2028 (O_2028,N_49629,N_49127);
and UO_2029 (O_2029,N_49633,N_49516);
xor UO_2030 (O_2030,N_49336,N_49613);
xor UO_2031 (O_2031,N_49232,N_49413);
nand UO_2032 (O_2032,N_49772,N_49828);
or UO_2033 (O_2033,N_49400,N_49632);
and UO_2034 (O_2034,N_49123,N_49721);
or UO_2035 (O_2035,N_49917,N_49619);
xor UO_2036 (O_2036,N_49349,N_49315);
nor UO_2037 (O_2037,N_49755,N_49088);
nand UO_2038 (O_2038,N_49851,N_49383);
or UO_2039 (O_2039,N_49381,N_49484);
or UO_2040 (O_2040,N_49941,N_49867);
and UO_2041 (O_2041,N_49346,N_49765);
and UO_2042 (O_2042,N_49250,N_49475);
or UO_2043 (O_2043,N_49153,N_49093);
or UO_2044 (O_2044,N_49956,N_49820);
nor UO_2045 (O_2045,N_49491,N_49140);
nor UO_2046 (O_2046,N_49216,N_49123);
nand UO_2047 (O_2047,N_49594,N_49231);
and UO_2048 (O_2048,N_49406,N_49480);
nand UO_2049 (O_2049,N_49588,N_49282);
or UO_2050 (O_2050,N_49708,N_49514);
xor UO_2051 (O_2051,N_49318,N_49456);
nor UO_2052 (O_2052,N_49695,N_49888);
and UO_2053 (O_2053,N_49051,N_49775);
nand UO_2054 (O_2054,N_49447,N_49501);
xor UO_2055 (O_2055,N_49511,N_49256);
xnor UO_2056 (O_2056,N_49946,N_49826);
and UO_2057 (O_2057,N_49618,N_49569);
nand UO_2058 (O_2058,N_49831,N_49727);
and UO_2059 (O_2059,N_49453,N_49002);
xor UO_2060 (O_2060,N_49515,N_49791);
nor UO_2061 (O_2061,N_49938,N_49714);
nor UO_2062 (O_2062,N_49617,N_49126);
or UO_2063 (O_2063,N_49591,N_49873);
nor UO_2064 (O_2064,N_49433,N_49499);
or UO_2065 (O_2065,N_49999,N_49617);
nand UO_2066 (O_2066,N_49463,N_49567);
nand UO_2067 (O_2067,N_49320,N_49180);
nor UO_2068 (O_2068,N_49353,N_49354);
nand UO_2069 (O_2069,N_49377,N_49727);
xnor UO_2070 (O_2070,N_49166,N_49290);
nand UO_2071 (O_2071,N_49641,N_49856);
or UO_2072 (O_2072,N_49656,N_49860);
nor UO_2073 (O_2073,N_49337,N_49923);
xnor UO_2074 (O_2074,N_49290,N_49209);
and UO_2075 (O_2075,N_49032,N_49736);
xnor UO_2076 (O_2076,N_49306,N_49204);
xor UO_2077 (O_2077,N_49303,N_49397);
nor UO_2078 (O_2078,N_49966,N_49236);
and UO_2079 (O_2079,N_49004,N_49145);
nor UO_2080 (O_2080,N_49888,N_49739);
or UO_2081 (O_2081,N_49307,N_49395);
and UO_2082 (O_2082,N_49754,N_49901);
nand UO_2083 (O_2083,N_49271,N_49459);
or UO_2084 (O_2084,N_49446,N_49364);
xor UO_2085 (O_2085,N_49076,N_49156);
nand UO_2086 (O_2086,N_49836,N_49239);
and UO_2087 (O_2087,N_49092,N_49511);
nor UO_2088 (O_2088,N_49844,N_49557);
nor UO_2089 (O_2089,N_49464,N_49845);
or UO_2090 (O_2090,N_49888,N_49597);
xor UO_2091 (O_2091,N_49196,N_49572);
or UO_2092 (O_2092,N_49236,N_49296);
nand UO_2093 (O_2093,N_49661,N_49831);
nor UO_2094 (O_2094,N_49618,N_49231);
xor UO_2095 (O_2095,N_49314,N_49130);
and UO_2096 (O_2096,N_49958,N_49072);
nand UO_2097 (O_2097,N_49415,N_49684);
xnor UO_2098 (O_2098,N_49475,N_49887);
nand UO_2099 (O_2099,N_49475,N_49546);
nor UO_2100 (O_2100,N_49515,N_49647);
or UO_2101 (O_2101,N_49754,N_49281);
xnor UO_2102 (O_2102,N_49662,N_49135);
and UO_2103 (O_2103,N_49964,N_49476);
or UO_2104 (O_2104,N_49157,N_49875);
nand UO_2105 (O_2105,N_49713,N_49998);
or UO_2106 (O_2106,N_49009,N_49504);
nor UO_2107 (O_2107,N_49165,N_49936);
or UO_2108 (O_2108,N_49535,N_49860);
xor UO_2109 (O_2109,N_49076,N_49037);
and UO_2110 (O_2110,N_49345,N_49206);
and UO_2111 (O_2111,N_49398,N_49833);
xnor UO_2112 (O_2112,N_49381,N_49778);
xor UO_2113 (O_2113,N_49721,N_49078);
or UO_2114 (O_2114,N_49817,N_49518);
and UO_2115 (O_2115,N_49723,N_49080);
nand UO_2116 (O_2116,N_49064,N_49476);
or UO_2117 (O_2117,N_49403,N_49832);
nand UO_2118 (O_2118,N_49626,N_49192);
xnor UO_2119 (O_2119,N_49058,N_49299);
or UO_2120 (O_2120,N_49497,N_49914);
or UO_2121 (O_2121,N_49946,N_49251);
nor UO_2122 (O_2122,N_49026,N_49985);
nand UO_2123 (O_2123,N_49991,N_49365);
or UO_2124 (O_2124,N_49973,N_49363);
nand UO_2125 (O_2125,N_49753,N_49308);
or UO_2126 (O_2126,N_49007,N_49583);
and UO_2127 (O_2127,N_49687,N_49768);
or UO_2128 (O_2128,N_49949,N_49017);
xnor UO_2129 (O_2129,N_49190,N_49000);
nor UO_2130 (O_2130,N_49223,N_49072);
nor UO_2131 (O_2131,N_49759,N_49301);
xor UO_2132 (O_2132,N_49337,N_49704);
nand UO_2133 (O_2133,N_49811,N_49819);
nand UO_2134 (O_2134,N_49032,N_49222);
nand UO_2135 (O_2135,N_49746,N_49592);
nor UO_2136 (O_2136,N_49092,N_49697);
nand UO_2137 (O_2137,N_49026,N_49377);
nand UO_2138 (O_2138,N_49070,N_49856);
nor UO_2139 (O_2139,N_49248,N_49080);
and UO_2140 (O_2140,N_49167,N_49903);
xor UO_2141 (O_2141,N_49343,N_49801);
and UO_2142 (O_2142,N_49643,N_49726);
or UO_2143 (O_2143,N_49729,N_49604);
and UO_2144 (O_2144,N_49909,N_49708);
and UO_2145 (O_2145,N_49921,N_49733);
xnor UO_2146 (O_2146,N_49196,N_49554);
or UO_2147 (O_2147,N_49643,N_49065);
and UO_2148 (O_2148,N_49393,N_49268);
and UO_2149 (O_2149,N_49563,N_49228);
or UO_2150 (O_2150,N_49703,N_49507);
nor UO_2151 (O_2151,N_49614,N_49569);
and UO_2152 (O_2152,N_49604,N_49746);
and UO_2153 (O_2153,N_49975,N_49057);
or UO_2154 (O_2154,N_49805,N_49103);
and UO_2155 (O_2155,N_49741,N_49710);
xor UO_2156 (O_2156,N_49277,N_49557);
or UO_2157 (O_2157,N_49373,N_49876);
and UO_2158 (O_2158,N_49068,N_49537);
xnor UO_2159 (O_2159,N_49359,N_49464);
and UO_2160 (O_2160,N_49374,N_49154);
xnor UO_2161 (O_2161,N_49365,N_49464);
or UO_2162 (O_2162,N_49095,N_49123);
and UO_2163 (O_2163,N_49470,N_49713);
and UO_2164 (O_2164,N_49685,N_49584);
nand UO_2165 (O_2165,N_49996,N_49047);
nor UO_2166 (O_2166,N_49602,N_49366);
and UO_2167 (O_2167,N_49864,N_49671);
or UO_2168 (O_2168,N_49266,N_49862);
nor UO_2169 (O_2169,N_49495,N_49783);
xnor UO_2170 (O_2170,N_49513,N_49026);
nand UO_2171 (O_2171,N_49268,N_49059);
and UO_2172 (O_2172,N_49830,N_49753);
and UO_2173 (O_2173,N_49667,N_49582);
nor UO_2174 (O_2174,N_49487,N_49708);
xor UO_2175 (O_2175,N_49410,N_49658);
or UO_2176 (O_2176,N_49749,N_49643);
or UO_2177 (O_2177,N_49061,N_49571);
nand UO_2178 (O_2178,N_49251,N_49597);
or UO_2179 (O_2179,N_49205,N_49928);
xor UO_2180 (O_2180,N_49254,N_49173);
nand UO_2181 (O_2181,N_49010,N_49376);
and UO_2182 (O_2182,N_49771,N_49197);
nand UO_2183 (O_2183,N_49562,N_49401);
and UO_2184 (O_2184,N_49595,N_49472);
xnor UO_2185 (O_2185,N_49818,N_49201);
nand UO_2186 (O_2186,N_49398,N_49866);
nor UO_2187 (O_2187,N_49699,N_49985);
or UO_2188 (O_2188,N_49581,N_49288);
and UO_2189 (O_2189,N_49045,N_49418);
xnor UO_2190 (O_2190,N_49042,N_49995);
xnor UO_2191 (O_2191,N_49665,N_49887);
xnor UO_2192 (O_2192,N_49749,N_49588);
nor UO_2193 (O_2193,N_49843,N_49853);
xnor UO_2194 (O_2194,N_49049,N_49327);
or UO_2195 (O_2195,N_49130,N_49377);
nand UO_2196 (O_2196,N_49935,N_49422);
nand UO_2197 (O_2197,N_49915,N_49639);
nor UO_2198 (O_2198,N_49001,N_49579);
and UO_2199 (O_2199,N_49244,N_49385);
or UO_2200 (O_2200,N_49793,N_49714);
nand UO_2201 (O_2201,N_49699,N_49168);
or UO_2202 (O_2202,N_49584,N_49975);
nand UO_2203 (O_2203,N_49531,N_49975);
xnor UO_2204 (O_2204,N_49427,N_49234);
xor UO_2205 (O_2205,N_49210,N_49576);
nor UO_2206 (O_2206,N_49936,N_49876);
xor UO_2207 (O_2207,N_49161,N_49531);
nor UO_2208 (O_2208,N_49199,N_49644);
or UO_2209 (O_2209,N_49144,N_49010);
nand UO_2210 (O_2210,N_49798,N_49812);
and UO_2211 (O_2211,N_49745,N_49400);
xnor UO_2212 (O_2212,N_49628,N_49786);
or UO_2213 (O_2213,N_49719,N_49604);
xnor UO_2214 (O_2214,N_49757,N_49205);
nand UO_2215 (O_2215,N_49146,N_49977);
nor UO_2216 (O_2216,N_49304,N_49458);
nor UO_2217 (O_2217,N_49375,N_49700);
and UO_2218 (O_2218,N_49933,N_49134);
or UO_2219 (O_2219,N_49237,N_49098);
xor UO_2220 (O_2220,N_49855,N_49903);
nor UO_2221 (O_2221,N_49856,N_49252);
and UO_2222 (O_2222,N_49509,N_49067);
nand UO_2223 (O_2223,N_49312,N_49332);
and UO_2224 (O_2224,N_49478,N_49918);
nor UO_2225 (O_2225,N_49301,N_49041);
or UO_2226 (O_2226,N_49299,N_49383);
nand UO_2227 (O_2227,N_49620,N_49730);
nand UO_2228 (O_2228,N_49126,N_49972);
xnor UO_2229 (O_2229,N_49274,N_49689);
or UO_2230 (O_2230,N_49402,N_49002);
nand UO_2231 (O_2231,N_49559,N_49208);
and UO_2232 (O_2232,N_49554,N_49928);
nor UO_2233 (O_2233,N_49410,N_49817);
nor UO_2234 (O_2234,N_49640,N_49618);
and UO_2235 (O_2235,N_49847,N_49692);
xor UO_2236 (O_2236,N_49447,N_49802);
nor UO_2237 (O_2237,N_49718,N_49774);
nand UO_2238 (O_2238,N_49344,N_49007);
nand UO_2239 (O_2239,N_49104,N_49972);
nand UO_2240 (O_2240,N_49045,N_49021);
nor UO_2241 (O_2241,N_49868,N_49477);
nor UO_2242 (O_2242,N_49550,N_49710);
nor UO_2243 (O_2243,N_49995,N_49280);
xnor UO_2244 (O_2244,N_49689,N_49155);
or UO_2245 (O_2245,N_49279,N_49537);
nor UO_2246 (O_2246,N_49104,N_49780);
nand UO_2247 (O_2247,N_49392,N_49322);
and UO_2248 (O_2248,N_49600,N_49109);
or UO_2249 (O_2249,N_49672,N_49003);
and UO_2250 (O_2250,N_49746,N_49987);
xor UO_2251 (O_2251,N_49683,N_49720);
xnor UO_2252 (O_2252,N_49239,N_49461);
nand UO_2253 (O_2253,N_49461,N_49535);
nand UO_2254 (O_2254,N_49707,N_49313);
and UO_2255 (O_2255,N_49362,N_49669);
and UO_2256 (O_2256,N_49324,N_49430);
and UO_2257 (O_2257,N_49266,N_49414);
nor UO_2258 (O_2258,N_49121,N_49960);
and UO_2259 (O_2259,N_49785,N_49210);
nor UO_2260 (O_2260,N_49132,N_49465);
nor UO_2261 (O_2261,N_49810,N_49968);
nand UO_2262 (O_2262,N_49381,N_49005);
and UO_2263 (O_2263,N_49413,N_49965);
or UO_2264 (O_2264,N_49774,N_49250);
nand UO_2265 (O_2265,N_49798,N_49178);
xnor UO_2266 (O_2266,N_49681,N_49852);
and UO_2267 (O_2267,N_49846,N_49907);
and UO_2268 (O_2268,N_49241,N_49714);
xnor UO_2269 (O_2269,N_49902,N_49029);
nor UO_2270 (O_2270,N_49819,N_49945);
nand UO_2271 (O_2271,N_49871,N_49145);
and UO_2272 (O_2272,N_49677,N_49615);
nand UO_2273 (O_2273,N_49995,N_49271);
nor UO_2274 (O_2274,N_49827,N_49464);
and UO_2275 (O_2275,N_49076,N_49984);
or UO_2276 (O_2276,N_49488,N_49541);
xor UO_2277 (O_2277,N_49038,N_49659);
and UO_2278 (O_2278,N_49859,N_49014);
nand UO_2279 (O_2279,N_49616,N_49012);
and UO_2280 (O_2280,N_49209,N_49463);
nor UO_2281 (O_2281,N_49105,N_49405);
xnor UO_2282 (O_2282,N_49871,N_49281);
and UO_2283 (O_2283,N_49382,N_49779);
xnor UO_2284 (O_2284,N_49693,N_49134);
and UO_2285 (O_2285,N_49549,N_49306);
nor UO_2286 (O_2286,N_49160,N_49562);
xor UO_2287 (O_2287,N_49964,N_49179);
or UO_2288 (O_2288,N_49755,N_49107);
nor UO_2289 (O_2289,N_49217,N_49691);
nand UO_2290 (O_2290,N_49518,N_49354);
nor UO_2291 (O_2291,N_49508,N_49751);
nand UO_2292 (O_2292,N_49412,N_49008);
xnor UO_2293 (O_2293,N_49195,N_49779);
and UO_2294 (O_2294,N_49512,N_49835);
or UO_2295 (O_2295,N_49387,N_49423);
xor UO_2296 (O_2296,N_49297,N_49916);
or UO_2297 (O_2297,N_49708,N_49196);
nand UO_2298 (O_2298,N_49656,N_49716);
xnor UO_2299 (O_2299,N_49839,N_49221);
or UO_2300 (O_2300,N_49628,N_49213);
xnor UO_2301 (O_2301,N_49877,N_49107);
nand UO_2302 (O_2302,N_49810,N_49157);
xnor UO_2303 (O_2303,N_49880,N_49068);
and UO_2304 (O_2304,N_49374,N_49767);
or UO_2305 (O_2305,N_49304,N_49725);
nand UO_2306 (O_2306,N_49734,N_49058);
xor UO_2307 (O_2307,N_49476,N_49921);
nor UO_2308 (O_2308,N_49339,N_49618);
and UO_2309 (O_2309,N_49362,N_49231);
nand UO_2310 (O_2310,N_49664,N_49843);
and UO_2311 (O_2311,N_49917,N_49661);
xnor UO_2312 (O_2312,N_49455,N_49846);
or UO_2313 (O_2313,N_49988,N_49281);
or UO_2314 (O_2314,N_49011,N_49303);
xor UO_2315 (O_2315,N_49173,N_49211);
or UO_2316 (O_2316,N_49571,N_49067);
nand UO_2317 (O_2317,N_49746,N_49296);
or UO_2318 (O_2318,N_49730,N_49731);
nor UO_2319 (O_2319,N_49902,N_49807);
xnor UO_2320 (O_2320,N_49597,N_49092);
nor UO_2321 (O_2321,N_49332,N_49838);
nand UO_2322 (O_2322,N_49713,N_49778);
nor UO_2323 (O_2323,N_49851,N_49307);
and UO_2324 (O_2324,N_49958,N_49667);
nand UO_2325 (O_2325,N_49800,N_49834);
nor UO_2326 (O_2326,N_49964,N_49867);
xor UO_2327 (O_2327,N_49568,N_49619);
and UO_2328 (O_2328,N_49684,N_49739);
xnor UO_2329 (O_2329,N_49786,N_49737);
or UO_2330 (O_2330,N_49682,N_49159);
nand UO_2331 (O_2331,N_49200,N_49156);
nor UO_2332 (O_2332,N_49615,N_49552);
or UO_2333 (O_2333,N_49837,N_49139);
nor UO_2334 (O_2334,N_49277,N_49165);
nor UO_2335 (O_2335,N_49098,N_49346);
nand UO_2336 (O_2336,N_49025,N_49829);
xnor UO_2337 (O_2337,N_49004,N_49186);
xor UO_2338 (O_2338,N_49492,N_49131);
and UO_2339 (O_2339,N_49470,N_49656);
nand UO_2340 (O_2340,N_49679,N_49614);
nand UO_2341 (O_2341,N_49200,N_49044);
nor UO_2342 (O_2342,N_49948,N_49576);
and UO_2343 (O_2343,N_49260,N_49638);
or UO_2344 (O_2344,N_49315,N_49607);
nor UO_2345 (O_2345,N_49602,N_49898);
or UO_2346 (O_2346,N_49383,N_49464);
nand UO_2347 (O_2347,N_49940,N_49259);
xnor UO_2348 (O_2348,N_49773,N_49974);
nor UO_2349 (O_2349,N_49604,N_49160);
or UO_2350 (O_2350,N_49392,N_49531);
xor UO_2351 (O_2351,N_49636,N_49493);
nand UO_2352 (O_2352,N_49678,N_49838);
nand UO_2353 (O_2353,N_49031,N_49237);
nor UO_2354 (O_2354,N_49638,N_49149);
xnor UO_2355 (O_2355,N_49293,N_49120);
and UO_2356 (O_2356,N_49162,N_49423);
xor UO_2357 (O_2357,N_49674,N_49645);
xnor UO_2358 (O_2358,N_49596,N_49554);
or UO_2359 (O_2359,N_49505,N_49065);
nor UO_2360 (O_2360,N_49011,N_49265);
xnor UO_2361 (O_2361,N_49897,N_49168);
nor UO_2362 (O_2362,N_49011,N_49827);
and UO_2363 (O_2363,N_49072,N_49906);
and UO_2364 (O_2364,N_49004,N_49333);
nor UO_2365 (O_2365,N_49994,N_49721);
and UO_2366 (O_2366,N_49216,N_49410);
nand UO_2367 (O_2367,N_49315,N_49177);
xor UO_2368 (O_2368,N_49451,N_49088);
nor UO_2369 (O_2369,N_49744,N_49646);
xor UO_2370 (O_2370,N_49169,N_49502);
xnor UO_2371 (O_2371,N_49497,N_49658);
or UO_2372 (O_2372,N_49351,N_49315);
xnor UO_2373 (O_2373,N_49575,N_49576);
and UO_2374 (O_2374,N_49787,N_49937);
nor UO_2375 (O_2375,N_49902,N_49612);
or UO_2376 (O_2376,N_49563,N_49940);
nor UO_2377 (O_2377,N_49785,N_49339);
nor UO_2378 (O_2378,N_49867,N_49289);
or UO_2379 (O_2379,N_49252,N_49239);
or UO_2380 (O_2380,N_49215,N_49301);
xnor UO_2381 (O_2381,N_49285,N_49335);
or UO_2382 (O_2382,N_49355,N_49104);
and UO_2383 (O_2383,N_49340,N_49197);
or UO_2384 (O_2384,N_49304,N_49785);
nor UO_2385 (O_2385,N_49839,N_49901);
nand UO_2386 (O_2386,N_49375,N_49304);
or UO_2387 (O_2387,N_49342,N_49870);
and UO_2388 (O_2388,N_49040,N_49701);
or UO_2389 (O_2389,N_49752,N_49728);
nor UO_2390 (O_2390,N_49994,N_49826);
or UO_2391 (O_2391,N_49850,N_49774);
nor UO_2392 (O_2392,N_49292,N_49067);
xor UO_2393 (O_2393,N_49034,N_49513);
nor UO_2394 (O_2394,N_49029,N_49593);
or UO_2395 (O_2395,N_49688,N_49294);
nand UO_2396 (O_2396,N_49714,N_49958);
nor UO_2397 (O_2397,N_49593,N_49816);
nand UO_2398 (O_2398,N_49096,N_49016);
nor UO_2399 (O_2399,N_49637,N_49665);
nand UO_2400 (O_2400,N_49648,N_49808);
nor UO_2401 (O_2401,N_49784,N_49599);
or UO_2402 (O_2402,N_49019,N_49304);
xor UO_2403 (O_2403,N_49681,N_49586);
nand UO_2404 (O_2404,N_49524,N_49126);
xor UO_2405 (O_2405,N_49553,N_49708);
and UO_2406 (O_2406,N_49671,N_49827);
nand UO_2407 (O_2407,N_49323,N_49286);
and UO_2408 (O_2408,N_49684,N_49554);
xor UO_2409 (O_2409,N_49653,N_49256);
nand UO_2410 (O_2410,N_49474,N_49675);
and UO_2411 (O_2411,N_49285,N_49485);
xnor UO_2412 (O_2412,N_49734,N_49384);
nand UO_2413 (O_2413,N_49468,N_49464);
or UO_2414 (O_2414,N_49853,N_49173);
nor UO_2415 (O_2415,N_49316,N_49976);
nand UO_2416 (O_2416,N_49460,N_49305);
xor UO_2417 (O_2417,N_49595,N_49962);
xnor UO_2418 (O_2418,N_49814,N_49688);
nor UO_2419 (O_2419,N_49843,N_49425);
nand UO_2420 (O_2420,N_49490,N_49558);
xnor UO_2421 (O_2421,N_49042,N_49242);
and UO_2422 (O_2422,N_49963,N_49762);
nor UO_2423 (O_2423,N_49442,N_49559);
and UO_2424 (O_2424,N_49112,N_49049);
nand UO_2425 (O_2425,N_49566,N_49172);
nand UO_2426 (O_2426,N_49074,N_49112);
nor UO_2427 (O_2427,N_49515,N_49695);
nand UO_2428 (O_2428,N_49189,N_49739);
and UO_2429 (O_2429,N_49023,N_49367);
xnor UO_2430 (O_2430,N_49630,N_49645);
xnor UO_2431 (O_2431,N_49886,N_49608);
nor UO_2432 (O_2432,N_49691,N_49445);
nor UO_2433 (O_2433,N_49622,N_49548);
and UO_2434 (O_2434,N_49306,N_49833);
and UO_2435 (O_2435,N_49445,N_49263);
xor UO_2436 (O_2436,N_49556,N_49336);
or UO_2437 (O_2437,N_49265,N_49201);
nand UO_2438 (O_2438,N_49056,N_49816);
nand UO_2439 (O_2439,N_49293,N_49358);
and UO_2440 (O_2440,N_49212,N_49196);
and UO_2441 (O_2441,N_49248,N_49901);
nand UO_2442 (O_2442,N_49543,N_49531);
nor UO_2443 (O_2443,N_49103,N_49341);
or UO_2444 (O_2444,N_49892,N_49086);
nand UO_2445 (O_2445,N_49818,N_49806);
nand UO_2446 (O_2446,N_49711,N_49436);
xnor UO_2447 (O_2447,N_49951,N_49579);
and UO_2448 (O_2448,N_49330,N_49323);
nor UO_2449 (O_2449,N_49656,N_49394);
or UO_2450 (O_2450,N_49184,N_49769);
nor UO_2451 (O_2451,N_49359,N_49051);
nor UO_2452 (O_2452,N_49079,N_49859);
nand UO_2453 (O_2453,N_49290,N_49370);
xor UO_2454 (O_2454,N_49011,N_49099);
or UO_2455 (O_2455,N_49010,N_49316);
nor UO_2456 (O_2456,N_49528,N_49447);
nor UO_2457 (O_2457,N_49647,N_49438);
or UO_2458 (O_2458,N_49291,N_49449);
and UO_2459 (O_2459,N_49484,N_49101);
nand UO_2460 (O_2460,N_49889,N_49537);
or UO_2461 (O_2461,N_49212,N_49092);
or UO_2462 (O_2462,N_49915,N_49412);
nand UO_2463 (O_2463,N_49189,N_49002);
or UO_2464 (O_2464,N_49902,N_49702);
xnor UO_2465 (O_2465,N_49816,N_49950);
and UO_2466 (O_2466,N_49822,N_49155);
or UO_2467 (O_2467,N_49561,N_49387);
or UO_2468 (O_2468,N_49401,N_49489);
and UO_2469 (O_2469,N_49919,N_49236);
nor UO_2470 (O_2470,N_49855,N_49548);
and UO_2471 (O_2471,N_49114,N_49664);
xnor UO_2472 (O_2472,N_49638,N_49076);
and UO_2473 (O_2473,N_49030,N_49458);
xor UO_2474 (O_2474,N_49191,N_49517);
or UO_2475 (O_2475,N_49117,N_49619);
xnor UO_2476 (O_2476,N_49582,N_49392);
nand UO_2477 (O_2477,N_49974,N_49920);
nand UO_2478 (O_2478,N_49582,N_49360);
xor UO_2479 (O_2479,N_49412,N_49079);
or UO_2480 (O_2480,N_49467,N_49963);
xnor UO_2481 (O_2481,N_49140,N_49907);
or UO_2482 (O_2482,N_49834,N_49462);
or UO_2483 (O_2483,N_49158,N_49341);
xnor UO_2484 (O_2484,N_49439,N_49111);
and UO_2485 (O_2485,N_49573,N_49599);
and UO_2486 (O_2486,N_49609,N_49346);
or UO_2487 (O_2487,N_49372,N_49902);
xor UO_2488 (O_2488,N_49873,N_49906);
nor UO_2489 (O_2489,N_49363,N_49814);
xnor UO_2490 (O_2490,N_49354,N_49497);
and UO_2491 (O_2491,N_49657,N_49107);
nand UO_2492 (O_2492,N_49700,N_49259);
or UO_2493 (O_2493,N_49100,N_49481);
xor UO_2494 (O_2494,N_49674,N_49507);
or UO_2495 (O_2495,N_49518,N_49283);
or UO_2496 (O_2496,N_49942,N_49473);
nor UO_2497 (O_2497,N_49044,N_49318);
and UO_2498 (O_2498,N_49970,N_49294);
or UO_2499 (O_2499,N_49425,N_49135);
xor UO_2500 (O_2500,N_49225,N_49133);
or UO_2501 (O_2501,N_49667,N_49255);
or UO_2502 (O_2502,N_49640,N_49373);
nand UO_2503 (O_2503,N_49334,N_49201);
nor UO_2504 (O_2504,N_49358,N_49978);
nor UO_2505 (O_2505,N_49829,N_49897);
xnor UO_2506 (O_2506,N_49810,N_49136);
or UO_2507 (O_2507,N_49282,N_49322);
nor UO_2508 (O_2508,N_49303,N_49807);
nor UO_2509 (O_2509,N_49520,N_49208);
nand UO_2510 (O_2510,N_49886,N_49793);
xor UO_2511 (O_2511,N_49812,N_49705);
or UO_2512 (O_2512,N_49434,N_49183);
or UO_2513 (O_2513,N_49357,N_49450);
nand UO_2514 (O_2514,N_49990,N_49873);
or UO_2515 (O_2515,N_49666,N_49061);
nor UO_2516 (O_2516,N_49168,N_49162);
nor UO_2517 (O_2517,N_49694,N_49988);
or UO_2518 (O_2518,N_49780,N_49626);
xnor UO_2519 (O_2519,N_49140,N_49473);
xor UO_2520 (O_2520,N_49220,N_49009);
nor UO_2521 (O_2521,N_49774,N_49475);
and UO_2522 (O_2522,N_49882,N_49330);
nor UO_2523 (O_2523,N_49634,N_49954);
xor UO_2524 (O_2524,N_49247,N_49702);
or UO_2525 (O_2525,N_49648,N_49468);
or UO_2526 (O_2526,N_49885,N_49235);
nor UO_2527 (O_2527,N_49206,N_49121);
xnor UO_2528 (O_2528,N_49136,N_49988);
nand UO_2529 (O_2529,N_49232,N_49173);
xor UO_2530 (O_2530,N_49017,N_49309);
and UO_2531 (O_2531,N_49095,N_49871);
xnor UO_2532 (O_2532,N_49681,N_49767);
or UO_2533 (O_2533,N_49122,N_49790);
nor UO_2534 (O_2534,N_49542,N_49993);
nand UO_2535 (O_2535,N_49736,N_49404);
nor UO_2536 (O_2536,N_49318,N_49699);
nor UO_2537 (O_2537,N_49227,N_49072);
xnor UO_2538 (O_2538,N_49468,N_49526);
nor UO_2539 (O_2539,N_49155,N_49355);
and UO_2540 (O_2540,N_49978,N_49901);
nor UO_2541 (O_2541,N_49374,N_49874);
nand UO_2542 (O_2542,N_49478,N_49220);
and UO_2543 (O_2543,N_49441,N_49975);
nand UO_2544 (O_2544,N_49312,N_49692);
and UO_2545 (O_2545,N_49032,N_49746);
xor UO_2546 (O_2546,N_49949,N_49419);
and UO_2547 (O_2547,N_49636,N_49380);
nand UO_2548 (O_2548,N_49717,N_49915);
xnor UO_2549 (O_2549,N_49479,N_49183);
and UO_2550 (O_2550,N_49722,N_49759);
or UO_2551 (O_2551,N_49586,N_49793);
xor UO_2552 (O_2552,N_49987,N_49430);
nor UO_2553 (O_2553,N_49266,N_49001);
nand UO_2554 (O_2554,N_49532,N_49951);
nor UO_2555 (O_2555,N_49407,N_49020);
nand UO_2556 (O_2556,N_49769,N_49734);
and UO_2557 (O_2557,N_49241,N_49684);
and UO_2558 (O_2558,N_49103,N_49870);
nand UO_2559 (O_2559,N_49897,N_49352);
xnor UO_2560 (O_2560,N_49228,N_49196);
or UO_2561 (O_2561,N_49211,N_49357);
or UO_2562 (O_2562,N_49601,N_49152);
xor UO_2563 (O_2563,N_49895,N_49994);
and UO_2564 (O_2564,N_49643,N_49508);
xnor UO_2565 (O_2565,N_49878,N_49943);
nand UO_2566 (O_2566,N_49810,N_49327);
and UO_2567 (O_2567,N_49447,N_49207);
nor UO_2568 (O_2568,N_49596,N_49927);
or UO_2569 (O_2569,N_49861,N_49642);
and UO_2570 (O_2570,N_49150,N_49330);
nor UO_2571 (O_2571,N_49676,N_49329);
nand UO_2572 (O_2572,N_49496,N_49311);
nand UO_2573 (O_2573,N_49942,N_49971);
xnor UO_2574 (O_2574,N_49124,N_49922);
nor UO_2575 (O_2575,N_49933,N_49201);
or UO_2576 (O_2576,N_49747,N_49632);
or UO_2577 (O_2577,N_49606,N_49426);
nor UO_2578 (O_2578,N_49761,N_49009);
or UO_2579 (O_2579,N_49269,N_49375);
nand UO_2580 (O_2580,N_49483,N_49201);
and UO_2581 (O_2581,N_49119,N_49292);
and UO_2582 (O_2582,N_49858,N_49648);
nor UO_2583 (O_2583,N_49393,N_49776);
and UO_2584 (O_2584,N_49752,N_49977);
nor UO_2585 (O_2585,N_49533,N_49452);
xnor UO_2586 (O_2586,N_49686,N_49024);
or UO_2587 (O_2587,N_49603,N_49827);
or UO_2588 (O_2588,N_49368,N_49761);
and UO_2589 (O_2589,N_49097,N_49675);
or UO_2590 (O_2590,N_49553,N_49751);
xnor UO_2591 (O_2591,N_49204,N_49600);
or UO_2592 (O_2592,N_49219,N_49321);
nand UO_2593 (O_2593,N_49957,N_49008);
nand UO_2594 (O_2594,N_49005,N_49717);
nor UO_2595 (O_2595,N_49010,N_49626);
or UO_2596 (O_2596,N_49497,N_49483);
and UO_2597 (O_2597,N_49105,N_49371);
or UO_2598 (O_2598,N_49228,N_49784);
and UO_2599 (O_2599,N_49679,N_49963);
xor UO_2600 (O_2600,N_49061,N_49335);
xnor UO_2601 (O_2601,N_49380,N_49223);
nor UO_2602 (O_2602,N_49810,N_49857);
and UO_2603 (O_2603,N_49845,N_49974);
nor UO_2604 (O_2604,N_49490,N_49635);
nand UO_2605 (O_2605,N_49575,N_49847);
nand UO_2606 (O_2606,N_49442,N_49405);
and UO_2607 (O_2607,N_49820,N_49784);
nor UO_2608 (O_2608,N_49059,N_49589);
nand UO_2609 (O_2609,N_49349,N_49749);
nand UO_2610 (O_2610,N_49237,N_49962);
xor UO_2611 (O_2611,N_49911,N_49806);
or UO_2612 (O_2612,N_49141,N_49899);
nand UO_2613 (O_2613,N_49499,N_49886);
nor UO_2614 (O_2614,N_49405,N_49864);
and UO_2615 (O_2615,N_49523,N_49391);
nor UO_2616 (O_2616,N_49290,N_49732);
nor UO_2617 (O_2617,N_49660,N_49992);
or UO_2618 (O_2618,N_49983,N_49406);
nand UO_2619 (O_2619,N_49716,N_49280);
or UO_2620 (O_2620,N_49299,N_49635);
and UO_2621 (O_2621,N_49448,N_49753);
nand UO_2622 (O_2622,N_49854,N_49382);
nand UO_2623 (O_2623,N_49330,N_49593);
and UO_2624 (O_2624,N_49740,N_49260);
xnor UO_2625 (O_2625,N_49653,N_49364);
nand UO_2626 (O_2626,N_49062,N_49362);
nor UO_2627 (O_2627,N_49345,N_49334);
and UO_2628 (O_2628,N_49836,N_49226);
nand UO_2629 (O_2629,N_49860,N_49829);
nand UO_2630 (O_2630,N_49986,N_49813);
nand UO_2631 (O_2631,N_49223,N_49021);
and UO_2632 (O_2632,N_49729,N_49882);
xnor UO_2633 (O_2633,N_49104,N_49901);
xnor UO_2634 (O_2634,N_49763,N_49703);
and UO_2635 (O_2635,N_49999,N_49564);
xnor UO_2636 (O_2636,N_49796,N_49710);
nor UO_2637 (O_2637,N_49908,N_49320);
nand UO_2638 (O_2638,N_49073,N_49127);
and UO_2639 (O_2639,N_49749,N_49556);
nand UO_2640 (O_2640,N_49959,N_49950);
nand UO_2641 (O_2641,N_49685,N_49482);
or UO_2642 (O_2642,N_49666,N_49411);
nor UO_2643 (O_2643,N_49934,N_49834);
and UO_2644 (O_2644,N_49233,N_49204);
and UO_2645 (O_2645,N_49495,N_49701);
nand UO_2646 (O_2646,N_49172,N_49642);
and UO_2647 (O_2647,N_49081,N_49171);
or UO_2648 (O_2648,N_49675,N_49342);
xnor UO_2649 (O_2649,N_49164,N_49701);
xor UO_2650 (O_2650,N_49059,N_49847);
and UO_2651 (O_2651,N_49495,N_49567);
and UO_2652 (O_2652,N_49159,N_49993);
or UO_2653 (O_2653,N_49398,N_49283);
or UO_2654 (O_2654,N_49101,N_49919);
nor UO_2655 (O_2655,N_49471,N_49230);
or UO_2656 (O_2656,N_49680,N_49059);
nand UO_2657 (O_2657,N_49735,N_49415);
or UO_2658 (O_2658,N_49313,N_49485);
and UO_2659 (O_2659,N_49044,N_49602);
nor UO_2660 (O_2660,N_49567,N_49998);
nor UO_2661 (O_2661,N_49077,N_49696);
and UO_2662 (O_2662,N_49487,N_49493);
xnor UO_2663 (O_2663,N_49673,N_49951);
nand UO_2664 (O_2664,N_49396,N_49383);
xnor UO_2665 (O_2665,N_49387,N_49386);
nor UO_2666 (O_2666,N_49674,N_49535);
and UO_2667 (O_2667,N_49656,N_49895);
nor UO_2668 (O_2668,N_49857,N_49313);
and UO_2669 (O_2669,N_49592,N_49662);
or UO_2670 (O_2670,N_49840,N_49073);
or UO_2671 (O_2671,N_49848,N_49895);
or UO_2672 (O_2672,N_49872,N_49509);
nand UO_2673 (O_2673,N_49708,N_49972);
nand UO_2674 (O_2674,N_49079,N_49140);
and UO_2675 (O_2675,N_49785,N_49039);
xor UO_2676 (O_2676,N_49620,N_49818);
and UO_2677 (O_2677,N_49258,N_49331);
and UO_2678 (O_2678,N_49199,N_49385);
xor UO_2679 (O_2679,N_49198,N_49517);
xnor UO_2680 (O_2680,N_49951,N_49830);
nor UO_2681 (O_2681,N_49216,N_49699);
or UO_2682 (O_2682,N_49094,N_49299);
nand UO_2683 (O_2683,N_49389,N_49646);
nor UO_2684 (O_2684,N_49667,N_49412);
nand UO_2685 (O_2685,N_49071,N_49483);
and UO_2686 (O_2686,N_49711,N_49235);
xor UO_2687 (O_2687,N_49079,N_49376);
nand UO_2688 (O_2688,N_49471,N_49678);
xor UO_2689 (O_2689,N_49067,N_49070);
nand UO_2690 (O_2690,N_49568,N_49542);
nand UO_2691 (O_2691,N_49404,N_49179);
and UO_2692 (O_2692,N_49542,N_49159);
xnor UO_2693 (O_2693,N_49553,N_49103);
and UO_2694 (O_2694,N_49699,N_49292);
nand UO_2695 (O_2695,N_49449,N_49117);
nor UO_2696 (O_2696,N_49216,N_49416);
nand UO_2697 (O_2697,N_49372,N_49369);
and UO_2698 (O_2698,N_49177,N_49630);
nand UO_2699 (O_2699,N_49545,N_49129);
nor UO_2700 (O_2700,N_49205,N_49518);
nor UO_2701 (O_2701,N_49419,N_49537);
and UO_2702 (O_2702,N_49101,N_49245);
nand UO_2703 (O_2703,N_49777,N_49022);
and UO_2704 (O_2704,N_49746,N_49841);
nor UO_2705 (O_2705,N_49211,N_49351);
and UO_2706 (O_2706,N_49352,N_49354);
nor UO_2707 (O_2707,N_49685,N_49491);
nor UO_2708 (O_2708,N_49203,N_49575);
or UO_2709 (O_2709,N_49309,N_49800);
and UO_2710 (O_2710,N_49926,N_49622);
xor UO_2711 (O_2711,N_49603,N_49314);
nor UO_2712 (O_2712,N_49920,N_49814);
nand UO_2713 (O_2713,N_49188,N_49599);
nand UO_2714 (O_2714,N_49624,N_49385);
nor UO_2715 (O_2715,N_49570,N_49712);
and UO_2716 (O_2716,N_49070,N_49393);
nand UO_2717 (O_2717,N_49217,N_49123);
xor UO_2718 (O_2718,N_49791,N_49248);
nor UO_2719 (O_2719,N_49073,N_49304);
nor UO_2720 (O_2720,N_49037,N_49363);
xor UO_2721 (O_2721,N_49486,N_49462);
and UO_2722 (O_2722,N_49814,N_49879);
xnor UO_2723 (O_2723,N_49324,N_49287);
or UO_2724 (O_2724,N_49196,N_49509);
nand UO_2725 (O_2725,N_49368,N_49982);
xor UO_2726 (O_2726,N_49559,N_49933);
or UO_2727 (O_2727,N_49125,N_49178);
and UO_2728 (O_2728,N_49313,N_49902);
xor UO_2729 (O_2729,N_49469,N_49840);
nor UO_2730 (O_2730,N_49209,N_49379);
and UO_2731 (O_2731,N_49065,N_49072);
or UO_2732 (O_2732,N_49858,N_49787);
nand UO_2733 (O_2733,N_49215,N_49780);
nor UO_2734 (O_2734,N_49646,N_49644);
and UO_2735 (O_2735,N_49409,N_49622);
xnor UO_2736 (O_2736,N_49948,N_49034);
nor UO_2737 (O_2737,N_49433,N_49686);
xnor UO_2738 (O_2738,N_49325,N_49608);
nor UO_2739 (O_2739,N_49792,N_49635);
nand UO_2740 (O_2740,N_49278,N_49509);
xnor UO_2741 (O_2741,N_49192,N_49993);
nor UO_2742 (O_2742,N_49742,N_49465);
xor UO_2743 (O_2743,N_49101,N_49441);
and UO_2744 (O_2744,N_49191,N_49802);
nor UO_2745 (O_2745,N_49356,N_49218);
xnor UO_2746 (O_2746,N_49451,N_49414);
xor UO_2747 (O_2747,N_49113,N_49911);
nand UO_2748 (O_2748,N_49657,N_49631);
xnor UO_2749 (O_2749,N_49568,N_49750);
nand UO_2750 (O_2750,N_49704,N_49835);
xor UO_2751 (O_2751,N_49167,N_49742);
or UO_2752 (O_2752,N_49449,N_49311);
and UO_2753 (O_2753,N_49990,N_49811);
xor UO_2754 (O_2754,N_49586,N_49713);
nor UO_2755 (O_2755,N_49010,N_49547);
xor UO_2756 (O_2756,N_49297,N_49001);
nand UO_2757 (O_2757,N_49333,N_49512);
nand UO_2758 (O_2758,N_49409,N_49605);
and UO_2759 (O_2759,N_49208,N_49566);
and UO_2760 (O_2760,N_49778,N_49096);
nand UO_2761 (O_2761,N_49221,N_49024);
and UO_2762 (O_2762,N_49952,N_49920);
nor UO_2763 (O_2763,N_49418,N_49515);
nor UO_2764 (O_2764,N_49323,N_49867);
and UO_2765 (O_2765,N_49902,N_49349);
or UO_2766 (O_2766,N_49913,N_49430);
xor UO_2767 (O_2767,N_49241,N_49853);
nor UO_2768 (O_2768,N_49947,N_49242);
nand UO_2769 (O_2769,N_49295,N_49463);
nor UO_2770 (O_2770,N_49207,N_49698);
or UO_2771 (O_2771,N_49652,N_49901);
or UO_2772 (O_2772,N_49503,N_49192);
nor UO_2773 (O_2773,N_49412,N_49369);
or UO_2774 (O_2774,N_49650,N_49341);
nand UO_2775 (O_2775,N_49285,N_49899);
nand UO_2776 (O_2776,N_49777,N_49759);
and UO_2777 (O_2777,N_49336,N_49661);
and UO_2778 (O_2778,N_49865,N_49945);
nor UO_2779 (O_2779,N_49377,N_49955);
nor UO_2780 (O_2780,N_49647,N_49652);
nand UO_2781 (O_2781,N_49489,N_49410);
nand UO_2782 (O_2782,N_49404,N_49315);
or UO_2783 (O_2783,N_49365,N_49866);
and UO_2784 (O_2784,N_49633,N_49222);
nor UO_2785 (O_2785,N_49063,N_49610);
nor UO_2786 (O_2786,N_49686,N_49602);
nand UO_2787 (O_2787,N_49582,N_49871);
or UO_2788 (O_2788,N_49459,N_49457);
or UO_2789 (O_2789,N_49573,N_49529);
or UO_2790 (O_2790,N_49793,N_49970);
or UO_2791 (O_2791,N_49473,N_49202);
nand UO_2792 (O_2792,N_49531,N_49445);
and UO_2793 (O_2793,N_49326,N_49232);
xnor UO_2794 (O_2794,N_49046,N_49012);
xor UO_2795 (O_2795,N_49319,N_49501);
and UO_2796 (O_2796,N_49708,N_49377);
xnor UO_2797 (O_2797,N_49629,N_49427);
or UO_2798 (O_2798,N_49723,N_49581);
nand UO_2799 (O_2799,N_49161,N_49007);
or UO_2800 (O_2800,N_49140,N_49505);
xnor UO_2801 (O_2801,N_49964,N_49906);
or UO_2802 (O_2802,N_49893,N_49419);
nand UO_2803 (O_2803,N_49469,N_49513);
and UO_2804 (O_2804,N_49967,N_49645);
nor UO_2805 (O_2805,N_49806,N_49661);
or UO_2806 (O_2806,N_49436,N_49278);
xor UO_2807 (O_2807,N_49504,N_49013);
xor UO_2808 (O_2808,N_49658,N_49592);
or UO_2809 (O_2809,N_49139,N_49408);
nand UO_2810 (O_2810,N_49754,N_49482);
and UO_2811 (O_2811,N_49465,N_49016);
or UO_2812 (O_2812,N_49032,N_49971);
nor UO_2813 (O_2813,N_49914,N_49313);
nand UO_2814 (O_2814,N_49005,N_49272);
or UO_2815 (O_2815,N_49354,N_49725);
and UO_2816 (O_2816,N_49324,N_49246);
and UO_2817 (O_2817,N_49574,N_49659);
xor UO_2818 (O_2818,N_49669,N_49596);
nor UO_2819 (O_2819,N_49097,N_49850);
or UO_2820 (O_2820,N_49758,N_49463);
and UO_2821 (O_2821,N_49607,N_49234);
or UO_2822 (O_2822,N_49830,N_49680);
or UO_2823 (O_2823,N_49700,N_49118);
nand UO_2824 (O_2824,N_49853,N_49871);
and UO_2825 (O_2825,N_49040,N_49068);
nand UO_2826 (O_2826,N_49508,N_49056);
xnor UO_2827 (O_2827,N_49714,N_49237);
or UO_2828 (O_2828,N_49894,N_49489);
or UO_2829 (O_2829,N_49221,N_49022);
and UO_2830 (O_2830,N_49895,N_49202);
and UO_2831 (O_2831,N_49478,N_49498);
nand UO_2832 (O_2832,N_49511,N_49717);
or UO_2833 (O_2833,N_49924,N_49474);
or UO_2834 (O_2834,N_49124,N_49108);
nor UO_2835 (O_2835,N_49173,N_49754);
nand UO_2836 (O_2836,N_49066,N_49729);
xor UO_2837 (O_2837,N_49791,N_49640);
or UO_2838 (O_2838,N_49229,N_49913);
and UO_2839 (O_2839,N_49242,N_49936);
xor UO_2840 (O_2840,N_49523,N_49238);
xnor UO_2841 (O_2841,N_49058,N_49110);
nand UO_2842 (O_2842,N_49800,N_49080);
or UO_2843 (O_2843,N_49123,N_49923);
xor UO_2844 (O_2844,N_49064,N_49151);
nand UO_2845 (O_2845,N_49314,N_49196);
and UO_2846 (O_2846,N_49045,N_49892);
nor UO_2847 (O_2847,N_49617,N_49182);
or UO_2848 (O_2848,N_49564,N_49673);
nor UO_2849 (O_2849,N_49826,N_49146);
or UO_2850 (O_2850,N_49893,N_49731);
or UO_2851 (O_2851,N_49941,N_49984);
nand UO_2852 (O_2852,N_49586,N_49906);
nor UO_2853 (O_2853,N_49283,N_49748);
or UO_2854 (O_2854,N_49946,N_49123);
nor UO_2855 (O_2855,N_49444,N_49842);
nor UO_2856 (O_2856,N_49044,N_49932);
or UO_2857 (O_2857,N_49361,N_49658);
or UO_2858 (O_2858,N_49115,N_49242);
nand UO_2859 (O_2859,N_49526,N_49986);
or UO_2860 (O_2860,N_49717,N_49342);
nor UO_2861 (O_2861,N_49213,N_49379);
and UO_2862 (O_2862,N_49507,N_49407);
nor UO_2863 (O_2863,N_49170,N_49320);
nand UO_2864 (O_2864,N_49367,N_49924);
xor UO_2865 (O_2865,N_49898,N_49434);
nand UO_2866 (O_2866,N_49627,N_49620);
and UO_2867 (O_2867,N_49250,N_49981);
nor UO_2868 (O_2868,N_49516,N_49489);
nand UO_2869 (O_2869,N_49508,N_49134);
xnor UO_2870 (O_2870,N_49290,N_49571);
xnor UO_2871 (O_2871,N_49577,N_49518);
and UO_2872 (O_2872,N_49422,N_49176);
xor UO_2873 (O_2873,N_49804,N_49030);
nand UO_2874 (O_2874,N_49843,N_49109);
nor UO_2875 (O_2875,N_49693,N_49668);
nor UO_2876 (O_2876,N_49569,N_49608);
nand UO_2877 (O_2877,N_49690,N_49405);
nor UO_2878 (O_2878,N_49780,N_49180);
or UO_2879 (O_2879,N_49459,N_49223);
xnor UO_2880 (O_2880,N_49750,N_49974);
nor UO_2881 (O_2881,N_49546,N_49837);
or UO_2882 (O_2882,N_49781,N_49808);
xnor UO_2883 (O_2883,N_49930,N_49011);
or UO_2884 (O_2884,N_49051,N_49531);
and UO_2885 (O_2885,N_49700,N_49962);
and UO_2886 (O_2886,N_49577,N_49281);
or UO_2887 (O_2887,N_49719,N_49393);
xor UO_2888 (O_2888,N_49931,N_49136);
nand UO_2889 (O_2889,N_49217,N_49784);
nor UO_2890 (O_2890,N_49891,N_49926);
nand UO_2891 (O_2891,N_49067,N_49485);
nor UO_2892 (O_2892,N_49137,N_49307);
and UO_2893 (O_2893,N_49223,N_49050);
or UO_2894 (O_2894,N_49363,N_49740);
nand UO_2895 (O_2895,N_49421,N_49711);
and UO_2896 (O_2896,N_49679,N_49618);
and UO_2897 (O_2897,N_49397,N_49089);
or UO_2898 (O_2898,N_49009,N_49498);
nor UO_2899 (O_2899,N_49635,N_49889);
nor UO_2900 (O_2900,N_49328,N_49327);
nand UO_2901 (O_2901,N_49859,N_49472);
xor UO_2902 (O_2902,N_49156,N_49610);
xnor UO_2903 (O_2903,N_49574,N_49221);
xor UO_2904 (O_2904,N_49524,N_49234);
or UO_2905 (O_2905,N_49195,N_49735);
nand UO_2906 (O_2906,N_49943,N_49051);
and UO_2907 (O_2907,N_49525,N_49587);
nor UO_2908 (O_2908,N_49257,N_49402);
or UO_2909 (O_2909,N_49452,N_49664);
nor UO_2910 (O_2910,N_49369,N_49117);
nand UO_2911 (O_2911,N_49863,N_49981);
nor UO_2912 (O_2912,N_49653,N_49976);
nor UO_2913 (O_2913,N_49678,N_49361);
and UO_2914 (O_2914,N_49326,N_49976);
nand UO_2915 (O_2915,N_49528,N_49433);
nor UO_2916 (O_2916,N_49758,N_49909);
and UO_2917 (O_2917,N_49580,N_49586);
xnor UO_2918 (O_2918,N_49439,N_49967);
nor UO_2919 (O_2919,N_49327,N_49016);
or UO_2920 (O_2920,N_49276,N_49651);
xor UO_2921 (O_2921,N_49286,N_49003);
or UO_2922 (O_2922,N_49154,N_49035);
or UO_2923 (O_2923,N_49445,N_49689);
nand UO_2924 (O_2924,N_49243,N_49993);
nor UO_2925 (O_2925,N_49016,N_49184);
and UO_2926 (O_2926,N_49653,N_49623);
or UO_2927 (O_2927,N_49354,N_49197);
nor UO_2928 (O_2928,N_49623,N_49166);
xnor UO_2929 (O_2929,N_49698,N_49729);
nor UO_2930 (O_2930,N_49477,N_49458);
and UO_2931 (O_2931,N_49334,N_49362);
and UO_2932 (O_2932,N_49691,N_49019);
and UO_2933 (O_2933,N_49345,N_49664);
and UO_2934 (O_2934,N_49847,N_49097);
or UO_2935 (O_2935,N_49860,N_49864);
or UO_2936 (O_2936,N_49173,N_49286);
xor UO_2937 (O_2937,N_49385,N_49240);
nor UO_2938 (O_2938,N_49831,N_49728);
and UO_2939 (O_2939,N_49622,N_49996);
nor UO_2940 (O_2940,N_49321,N_49241);
nor UO_2941 (O_2941,N_49476,N_49770);
xor UO_2942 (O_2942,N_49608,N_49806);
and UO_2943 (O_2943,N_49368,N_49080);
nand UO_2944 (O_2944,N_49687,N_49322);
xnor UO_2945 (O_2945,N_49378,N_49670);
xnor UO_2946 (O_2946,N_49140,N_49158);
nor UO_2947 (O_2947,N_49458,N_49855);
and UO_2948 (O_2948,N_49518,N_49634);
nor UO_2949 (O_2949,N_49568,N_49851);
xor UO_2950 (O_2950,N_49261,N_49675);
nor UO_2951 (O_2951,N_49385,N_49109);
xnor UO_2952 (O_2952,N_49016,N_49494);
nand UO_2953 (O_2953,N_49404,N_49498);
nand UO_2954 (O_2954,N_49453,N_49996);
xor UO_2955 (O_2955,N_49121,N_49185);
nand UO_2956 (O_2956,N_49065,N_49258);
or UO_2957 (O_2957,N_49227,N_49530);
and UO_2958 (O_2958,N_49547,N_49490);
xor UO_2959 (O_2959,N_49587,N_49120);
xor UO_2960 (O_2960,N_49888,N_49267);
and UO_2961 (O_2961,N_49581,N_49280);
and UO_2962 (O_2962,N_49860,N_49985);
and UO_2963 (O_2963,N_49647,N_49701);
and UO_2964 (O_2964,N_49377,N_49405);
nand UO_2965 (O_2965,N_49900,N_49878);
and UO_2966 (O_2966,N_49453,N_49217);
xor UO_2967 (O_2967,N_49499,N_49207);
nand UO_2968 (O_2968,N_49540,N_49898);
or UO_2969 (O_2969,N_49076,N_49309);
nor UO_2970 (O_2970,N_49074,N_49329);
or UO_2971 (O_2971,N_49030,N_49479);
or UO_2972 (O_2972,N_49356,N_49880);
xor UO_2973 (O_2973,N_49943,N_49492);
or UO_2974 (O_2974,N_49241,N_49544);
nand UO_2975 (O_2975,N_49355,N_49844);
and UO_2976 (O_2976,N_49621,N_49254);
or UO_2977 (O_2977,N_49491,N_49889);
nor UO_2978 (O_2978,N_49412,N_49175);
or UO_2979 (O_2979,N_49775,N_49638);
and UO_2980 (O_2980,N_49665,N_49820);
xor UO_2981 (O_2981,N_49035,N_49917);
xnor UO_2982 (O_2982,N_49470,N_49208);
or UO_2983 (O_2983,N_49576,N_49435);
and UO_2984 (O_2984,N_49380,N_49896);
and UO_2985 (O_2985,N_49938,N_49122);
nor UO_2986 (O_2986,N_49698,N_49915);
or UO_2987 (O_2987,N_49361,N_49635);
nor UO_2988 (O_2988,N_49888,N_49077);
or UO_2989 (O_2989,N_49746,N_49595);
and UO_2990 (O_2990,N_49004,N_49746);
xnor UO_2991 (O_2991,N_49253,N_49845);
nand UO_2992 (O_2992,N_49444,N_49546);
xnor UO_2993 (O_2993,N_49144,N_49940);
nand UO_2994 (O_2994,N_49295,N_49019);
xnor UO_2995 (O_2995,N_49213,N_49514);
nand UO_2996 (O_2996,N_49569,N_49665);
xor UO_2997 (O_2997,N_49233,N_49507);
xor UO_2998 (O_2998,N_49185,N_49880);
nand UO_2999 (O_2999,N_49170,N_49598);
and UO_3000 (O_3000,N_49078,N_49024);
nand UO_3001 (O_3001,N_49906,N_49499);
xnor UO_3002 (O_3002,N_49532,N_49158);
nor UO_3003 (O_3003,N_49169,N_49150);
and UO_3004 (O_3004,N_49483,N_49655);
and UO_3005 (O_3005,N_49888,N_49770);
xor UO_3006 (O_3006,N_49293,N_49447);
and UO_3007 (O_3007,N_49430,N_49699);
xor UO_3008 (O_3008,N_49770,N_49417);
xnor UO_3009 (O_3009,N_49096,N_49568);
nand UO_3010 (O_3010,N_49319,N_49262);
xnor UO_3011 (O_3011,N_49196,N_49372);
nor UO_3012 (O_3012,N_49447,N_49573);
and UO_3013 (O_3013,N_49472,N_49618);
nand UO_3014 (O_3014,N_49964,N_49892);
nand UO_3015 (O_3015,N_49725,N_49530);
nand UO_3016 (O_3016,N_49591,N_49656);
or UO_3017 (O_3017,N_49848,N_49495);
xor UO_3018 (O_3018,N_49585,N_49578);
and UO_3019 (O_3019,N_49680,N_49200);
and UO_3020 (O_3020,N_49322,N_49343);
or UO_3021 (O_3021,N_49967,N_49608);
or UO_3022 (O_3022,N_49237,N_49955);
xnor UO_3023 (O_3023,N_49960,N_49269);
nand UO_3024 (O_3024,N_49729,N_49612);
nand UO_3025 (O_3025,N_49754,N_49303);
xor UO_3026 (O_3026,N_49481,N_49793);
xor UO_3027 (O_3027,N_49938,N_49699);
or UO_3028 (O_3028,N_49487,N_49611);
or UO_3029 (O_3029,N_49746,N_49567);
nand UO_3030 (O_3030,N_49593,N_49879);
nor UO_3031 (O_3031,N_49195,N_49583);
or UO_3032 (O_3032,N_49969,N_49973);
and UO_3033 (O_3033,N_49802,N_49352);
and UO_3034 (O_3034,N_49177,N_49165);
nor UO_3035 (O_3035,N_49378,N_49490);
nand UO_3036 (O_3036,N_49903,N_49184);
nand UO_3037 (O_3037,N_49949,N_49022);
xor UO_3038 (O_3038,N_49939,N_49254);
or UO_3039 (O_3039,N_49191,N_49591);
nor UO_3040 (O_3040,N_49554,N_49906);
xnor UO_3041 (O_3041,N_49051,N_49291);
nand UO_3042 (O_3042,N_49025,N_49704);
or UO_3043 (O_3043,N_49376,N_49959);
nor UO_3044 (O_3044,N_49399,N_49461);
or UO_3045 (O_3045,N_49080,N_49976);
xor UO_3046 (O_3046,N_49927,N_49121);
nor UO_3047 (O_3047,N_49230,N_49033);
xnor UO_3048 (O_3048,N_49151,N_49742);
nor UO_3049 (O_3049,N_49464,N_49964);
nand UO_3050 (O_3050,N_49362,N_49491);
xor UO_3051 (O_3051,N_49463,N_49199);
and UO_3052 (O_3052,N_49305,N_49967);
nor UO_3053 (O_3053,N_49976,N_49882);
or UO_3054 (O_3054,N_49249,N_49566);
or UO_3055 (O_3055,N_49811,N_49592);
nand UO_3056 (O_3056,N_49939,N_49326);
nor UO_3057 (O_3057,N_49590,N_49962);
or UO_3058 (O_3058,N_49773,N_49480);
nand UO_3059 (O_3059,N_49993,N_49587);
nor UO_3060 (O_3060,N_49052,N_49711);
xnor UO_3061 (O_3061,N_49738,N_49516);
nor UO_3062 (O_3062,N_49913,N_49299);
nand UO_3063 (O_3063,N_49843,N_49808);
and UO_3064 (O_3064,N_49621,N_49665);
or UO_3065 (O_3065,N_49452,N_49352);
nor UO_3066 (O_3066,N_49479,N_49487);
nand UO_3067 (O_3067,N_49344,N_49073);
nand UO_3068 (O_3068,N_49857,N_49994);
xor UO_3069 (O_3069,N_49102,N_49508);
xnor UO_3070 (O_3070,N_49780,N_49313);
nand UO_3071 (O_3071,N_49506,N_49553);
and UO_3072 (O_3072,N_49119,N_49964);
and UO_3073 (O_3073,N_49614,N_49426);
or UO_3074 (O_3074,N_49177,N_49907);
xor UO_3075 (O_3075,N_49622,N_49731);
nor UO_3076 (O_3076,N_49332,N_49901);
nand UO_3077 (O_3077,N_49619,N_49959);
or UO_3078 (O_3078,N_49507,N_49073);
xor UO_3079 (O_3079,N_49714,N_49042);
and UO_3080 (O_3080,N_49582,N_49646);
and UO_3081 (O_3081,N_49812,N_49589);
or UO_3082 (O_3082,N_49086,N_49083);
or UO_3083 (O_3083,N_49843,N_49306);
nand UO_3084 (O_3084,N_49578,N_49451);
nor UO_3085 (O_3085,N_49259,N_49611);
nor UO_3086 (O_3086,N_49704,N_49559);
nor UO_3087 (O_3087,N_49822,N_49556);
or UO_3088 (O_3088,N_49945,N_49276);
nor UO_3089 (O_3089,N_49542,N_49686);
nor UO_3090 (O_3090,N_49840,N_49774);
or UO_3091 (O_3091,N_49022,N_49248);
nor UO_3092 (O_3092,N_49187,N_49735);
and UO_3093 (O_3093,N_49205,N_49660);
nand UO_3094 (O_3094,N_49989,N_49763);
nand UO_3095 (O_3095,N_49353,N_49727);
and UO_3096 (O_3096,N_49293,N_49576);
xor UO_3097 (O_3097,N_49463,N_49324);
nor UO_3098 (O_3098,N_49483,N_49390);
nand UO_3099 (O_3099,N_49000,N_49809);
or UO_3100 (O_3100,N_49079,N_49818);
and UO_3101 (O_3101,N_49796,N_49928);
or UO_3102 (O_3102,N_49795,N_49592);
nand UO_3103 (O_3103,N_49426,N_49079);
nor UO_3104 (O_3104,N_49580,N_49288);
nor UO_3105 (O_3105,N_49175,N_49582);
nor UO_3106 (O_3106,N_49305,N_49978);
xor UO_3107 (O_3107,N_49297,N_49254);
nand UO_3108 (O_3108,N_49905,N_49197);
or UO_3109 (O_3109,N_49043,N_49413);
nor UO_3110 (O_3110,N_49821,N_49539);
or UO_3111 (O_3111,N_49837,N_49171);
and UO_3112 (O_3112,N_49510,N_49833);
nand UO_3113 (O_3113,N_49671,N_49878);
or UO_3114 (O_3114,N_49700,N_49709);
nand UO_3115 (O_3115,N_49810,N_49971);
xor UO_3116 (O_3116,N_49893,N_49576);
xor UO_3117 (O_3117,N_49216,N_49605);
nor UO_3118 (O_3118,N_49911,N_49692);
xor UO_3119 (O_3119,N_49165,N_49098);
and UO_3120 (O_3120,N_49789,N_49643);
and UO_3121 (O_3121,N_49354,N_49862);
and UO_3122 (O_3122,N_49564,N_49184);
or UO_3123 (O_3123,N_49985,N_49281);
or UO_3124 (O_3124,N_49620,N_49099);
or UO_3125 (O_3125,N_49899,N_49350);
nand UO_3126 (O_3126,N_49110,N_49068);
and UO_3127 (O_3127,N_49506,N_49326);
xor UO_3128 (O_3128,N_49514,N_49264);
and UO_3129 (O_3129,N_49838,N_49774);
nand UO_3130 (O_3130,N_49866,N_49355);
or UO_3131 (O_3131,N_49433,N_49865);
and UO_3132 (O_3132,N_49921,N_49193);
xor UO_3133 (O_3133,N_49988,N_49997);
nand UO_3134 (O_3134,N_49252,N_49189);
xor UO_3135 (O_3135,N_49593,N_49529);
xor UO_3136 (O_3136,N_49452,N_49347);
or UO_3137 (O_3137,N_49186,N_49837);
nand UO_3138 (O_3138,N_49873,N_49178);
nand UO_3139 (O_3139,N_49883,N_49781);
nand UO_3140 (O_3140,N_49772,N_49184);
nand UO_3141 (O_3141,N_49477,N_49530);
nor UO_3142 (O_3142,N_49537,N_49818);
or UO_3143 (O_3143,N_49487,N_49734);
xnor UO_3144 (O_3144,N_49764,N_49876);
nand UO_3145 (O_3145,N_49797,N_49417);
nor UO_3146 (O_3146,N_49143,N_49757);
or UO_3147 (O_3147,N_49010,N_49061);
xnor UO_3148 (O_3148,N_49266,N_49597);
or UO_3149 (O_3149,N_49771,N_49954);
and UO_3150 (O_3150,N_49053,N_49938);
nand UO_3151 (O_3151,N_49306,N_49380);
and UO_3152 (O_3152,N_49273,N_49956);
and UO_3153 (O_3153,N_49176,N_49383);
nand UO_3154 (O_3154,N_49044,N_49021);
or UO_3155 (O_3155,N_49021,N_49502);
xnor UO_3156 (O_3156,N_49976,N_49825);
and UO_3157 (O_3157,N_49506,N_49712);
nand UO_3158 (O_3158,N_49059,N_49490);
nor UO_3159 (O_3159,N_49984,N_49600);
and UO_3160 (O_3160,N_49065,N_49021);
xor UO_3161 (O_3161,N_49150,N_49849);
xnor UO_3162 (O_3162,N_49821,N_49263);
xnor UO_3163 (O_3163,N_49244,N_49343);
nor UO_3164 (O_3164,N_49900,N_49371);
and UO_3165 (O_3165,N_49730,N_49031);
or UO_3166 (O_3166,N_49875,N_49268);
xnor UO_3167 (O_3167,N_49131,N_49873);
or UO_3168 (O_3168,N_49155,N_49426);
nor UO_3169 (O_3169,N_49074,N_49802);
nand UO_3170 (O_3170,N_49539,N_49357);
or UO_3171 (O_3171,N_49568,N_49559);
nand UO_3172 (O_3172,N_49635,N_49742);
and UO_3173 (O_3173,N_49305,N_49953);
xor UO_3174 (O_3174,N_49457,N_49492);
and UO_3175 (O_3175,N_49739,N_49052);
xor UO_3176 (O_3176,N_49630,N_49570);
and UO_3177 (O_3177,N_49178,N_49497);
nand UO_3178 (O_3178,N_49012,N_49152);
and UO_3179 (O_3179,N_49740,N_49417);
nor UO_3180 (O_3180,N_49700,N_49533);
or UO_3181 (O_3181,N_49100,N_49207);
xnor UO_3182 (O_3182,N_49404,N_49728);
nor UO_3183 (O_3183,N_49084,N_49270);
nand UO_3184 (O_3184,N_49406,N_49274);
nand UO_3185 (O_3185,N_49987,N_49469);
nor UO_3186 (O_3186,N_49325,N_49989);
and UO_3187 (O_3187,N_49498,N_49638);
xnor UO_3188 (O_3188,N_49383,N_49835);
nand UO_3189 (O_3189,N_49657,N_49273);
or UO_3190 (O_3190,N_49909,N_49158);
nor UO_3191 (O_3191,N_49440,N_49678);
and UO_3192 (O_3192,N_49252,N_49133);
nand UO_3193 (O_3193,N_49941,N_49811);
xnor UO_3194 (O_3194,N_49886,N_49211);
nor UO_3195 (O_3195,N_49055,N_49172);
and UO_3196 (O_3196,N_49465,N_49302);
nand UO_3197 (O_3197,N_49217,N_49468);
nand UO_3198 (O_3198,N_49466,N_49511);
and UO_3199 (O_3199,N_49522,N_49317);
nand UO_3200 (O_3200,N_49233,N_49194);
nand UO_3201 (O_3201,N_49354,N_49038);
nor UO_3202 (O_3202,N_49648,N_49889);
xnor UO_3203 (O_3203,N_49716,N_49461);
nand UO_3204 (O_3204,N_49860,N_49593);
nor UO_3205 (O_3205,N_49771,N_49980);
nor UO_3206 (O_3206,N_49983,N_49448);
and UO_3207 (O_3207,N_49694,N_49912);
or UO_3208 (O_3208,N_49331,N_49004);
xor UO_3209 (O_3209,N_49194,N_49624);
nand UO_3210 (O_3210,N_49271,N_49718);
or UO_3211 (O_3211,N_49122,N_49329);
or UO_3212 (O_3212,N_49162,N_49372);
nand UO_3213 (O_3213,N_49209,N_49605);
nand UO_3214 (O_3214,N_49257,N_49606);
xnor UO_3215 (O_3215,N_49545,N_49655);
xnor UO_3216 (O_3216,N_49929,N_49710);
nand UO_3217 (O_3217,N_49339,N_49898);
nand UO_3218 (O_3218,N_49181,N_49176);
or UO_3219 (O_3219,N_49128,N_49286);
and UO_3220 (O_3220,N_49535,N_49536);
nand UO_3221 (O_3221,N_49889,N_49800);
nand UO_3222 (O_3222,N_49542,N_49448);
or UO_3223 (O_3223,N_49061,N_49232);
nand UO_3224 (O_3224,N_49417,N_49840);
xnor UO_3225 (O_3225,N_49136,N_49196);
xnor UO_3226 (O_3226,N_49817,N_49006);
nor UO_3227 (O_3227,N_49832,N_49525);
nor UO_3228 (O_3228,N_49052,N_49322);
and UO_3229 (O_3229,N_49660,N_49289);
xor UO_3230 (O_3230,N_49314,N_49105);
or UO_3231 (O_3231,N_49716,N_49622);
xnor UO_3232 (O_3232,N_49738,N_49041);
and UO_3233 (O_3233,N_49364,N_49310);
nor UO_3234 (O_3234,N_49765,N_49254);
nor UO_3235 (O_3235,N_49626,N_49257);
xnor UO_3236 (O_3236,N_49354,N_49081);
nand UO_3237 (O_3237,N_49773,N_49860);
and UO_3238 (O_3238,N_49886,N_49792);
nand UO_3239 (O_3239,N_49058,N_49373);
xor UO_3240 (O_3240,N_49414,N_49742);
nor UO_3241 (O_3241,N_49227,N_49456);
nand UO_3242 (O_3242,N_49883,N_49441);
and UO_3243 (O_3243,N_49453,N_49036);
nor UO_3244 (O_3244,N_49166,N_49705);
and UO_3245 (O_3245,N_49067,N_49323);
xnor UO_3246 (O_3246,N_49948,N_49388);
xnor UO_3247 (O_3247,N_49598,N_49342);
and UO_3248 (O_3248,N_49812,N_49325);
nor UO_3249 (O_3249,N_49477,N_49106);
nor UO_3250 (O_3250,N_49153,N_49691);
or UO_3251 (O_3251,N_49915,N_49449);
and UO_3252 (O_3252,N_49789,N_49403);
and UO_3253 (O_3253,N_49587,N_49541);
xor UO_3254 (O_3254,N_49380,N_49818);
nand UO_3255 (O_3255,N_49258,N_49485);
and UO_3256 (O_3256,N_49146,N_49426);
or UO_3257 (O_3257,N_49170,N_49956);
and UO_3258 (O_3258,N_49818,N_49335);
nor UO_3259 (O_3259,N_49244,N_49101);
nor UO_3260 (O_3260,N_49229,N_49737);
and UO_3261 (O_3261,N_49475,N_49493);
nor UO_3262 (O_3262,N_49783,N_49108);
or UO_3263 (O_3263,N_49512,N_49364);
and UO_3264 (O_3264,N_49843,N_49035);
xor UO_3265 (O_3265,N_49091,N_49574);
nor UO_3266 (O_3266,N_49948,N_49091);
nor UO_3267 (O_3267,N_49487,N_49206);
and UO_3268 (O_3268,N_49130,N_49119);
or UO_3269 (O_3269,N_49695,N_49800);
nor UO_3270 (O_3270,N_49567,N_49202);
or UO_3271 (O_3271,N_49259,N_49996);
nor UO_3272 (O_3272,N_49874,N_49525);
and UO_3273 (O_3273,N_49870,N_49285);
xnor UO_3274 (O_3274,N_49497,N_49962);
nand UO_3275 (O_3275,N_49052,N_49404);
nor UO_3276 (O_3276,N_49404,N_49561);
xnor UO_3277 (O_3277,N_49452,N_49907);
nor UO_3278 (O_3278,N_49613,N_49847);
or UO_3279 (O_3279,N_49636,N_49539);
and UO_3280 (O_3280,N_49566,N_49499);
and UO_3281 (O_3281,N_49066,N_49354);
nand UO_3282 (O_3282,N_49624,N_49751);
or UO_3283 (O_3283,N_49706,N_49449);
xor UO_3284 (O_3284,N_49002,N_49574);
and UO_3285 (O_3285,N_49455,N_49943);
or UO_3286 (O_3286,N_49627,N_49261);
nand UO_3287 (O_3287,N_49632,N_49495);
and UO_3288 (O_3288,N_49379,N_49550);
and UO_3289 (O_3289,N_49568,N_49620);
xor UO_3290 (O_3290,N_49494,N_49662);
xnor UO_3291 (O_3291,N_49623,N_49271);
xor UO_3292 (O_3292,N_49238,N_49796);
nor UO_3293 (O_3293,N_49881,N_49069);
and UO_3294 (O_3294,N_49159,N_49283);
and UO_3295 (O_3295,N_49063,N_49733);
or UO_3296 (O_3296,N_49523,N_49113);
nor UO_3297 (O_3297,N_49708,N_49433);
xor UO_3298 (O_3298,N_49969,N_49738);
nor UO_3299 (O_3299,N_49759,N_49776);
nor UO_3300 (O_3300,N_49264,N_49725);
xnor UO_3301 (O_3301,N_49775,N_49268);
or UO_3302 (O_3302,N_49369,N_49167);
xnor UO_3303 (O_3303,N_49430,N_49905);
or UO_3304 (O_3304,N_49166,N_49882);
nor UO_3305 (O_3305,N_49443,N_49164);
nor UO_3306 (O_3306,N_49216,N_49960);
xor UO_3307 (O_3307,N_49935,N_49751);
or UO_3308 (O_3308,N_49307,N_49335);
or UO_3309 (O_3309,N_49977,N_49543);
or UO_3310 (O_3310,N_49123,N_49785);
nor UO_3311 (O_3311,N_49720,N_49584);
nor UO_3312 (O_3312,N_49913,N_49595);
or UO_3313 (O_3313,N_49222,N_49238);
and UO_3314 (O_3314,N_49694,N_49056);
nand UO_3315 (O_3315,N_49591,N_49627);
or UO_3316 (O_3316,N_49538,N_49701);
xnor UO_3317 (O_3317,N_49304,N_49376);
or UO_3318 (O_3318,N_49861,N_49990);
xor UO_3319 (O_3319,N_49755,N_49548);
nor UO_3320 (O_3320,N_49929,N_49694);
nor UO_3321 (O_3321,N_49267,N_49218);
nand UO_3322 (O_3322,N_49573,N_49673);
nor UO_3323 (O_3323,N_49462,N_49494);
and UO_3324 (O_3324,N_49273,N_49249);
nand UO_3325 (O_3325,N_49331,N_49700);
or UO_3326 (O_3326,N_49091,N_49491);
nand UO_3327 (O_3327,N_49420,N_49579);
or UO_3328 (O_3328,N_49664,N_49825);
xor UO_3329 (O_3329,N_49345,N_49032);
nor UO_3330 (O_3330,N_49461,N_49942);
nor UO_3331 (O_3331,N_49474,N_49763);
nand UO_3332 (O_3332,N_49572,N_49108);
nand UO_3333 (O_3333,N_49881,N_49840);
nor UO_3334 (O_3334,N_49909,N_49284);
and UO_3335 (O_3335,N_49743,N_49264);
and UO_3336 (O_3336,N_49527,N_49335);
nor UO_3337 (O_3337,N_49577,N_49819);
or UO_3338 (O_3338,N_49640,N_49558);
or UO_3339 (O_3339,N_49373,N_49820);
and UO_3340 (O_3340,N_49703,N_49854);
nor UO_3341 (O_3341,N_49020,N_49476);
nand UO_3342 (O_3342,N_49014,N_49416);
and UO_3343 (O_3343,N_49169,N_49383);
and UO_3344 (O_3344,N_49410,N_49054);
or UO_3345 (O_3345,N_49352,N_49329);
nor UO_3346 (O_3346,N_49612,N_49102);
nor UO_3347 (O_3347,N_49425,N_49641);
and UO_3348 (O_3348,N_49174,N_49430);
and UO_3349 (O_3349,N_49300,N_49268);
or UO_3350 (O_3350,N_49899,N_49405);
xnor UO_3351 (O_3351,N_49597,N_49404);
nand UO_3352 (O_3352,N_49237,N_49986);
or UO_3353 (O_3353,N_49474,N_49608);
xnor UO_3354 (O_3354,N_49796,N_49726);
or UO_3355 (O_3355,N_49038,N_49623);
nor UO_3356 (O_3356,N_49031,N_49598);
xor UO_3357 (O_3357,N_49948,N_49235);
xor UO_3358 (O_3358,N_49704,N_49369);
and UO_3359 (O_3359,N_49094,N_49268);
nand UO_3360 (O_3360,N_49938,N_49639);
nand UO_3361 (O_3361,N_49022,N_49939);
nand UO_3362 (O_3362,N_49954,N_49142);
or UO_3363 (O_3363,N_49826,N_49938);
nand UO_3364 (O_3364,N_49476,N_49311);
nand UO_3365 (O_3365,N_49630,N_49646);
or UO_3366 (O_3366,N_49008,N_49012);
and UO_3367 (O_3367,N_49283,N_49131);
nor UO_3368 (O_3368,N_49688,N_49270);
or UO_3369 (O_3369,N_49130,N_49227);
nand UO_3370 (O_3370,N_49965,N_49707);
nor UO_3371 (O_3371,N_49314,N_49516);
nor UO_3372 (O_3372,N_49074,N_49454);
and UO_3373 (O_3373,N_49015,N_49065);
xnor UO_3374 (O_3374,N_49956,N_49494);
or UO_3375 (O_3375,N_49233,N_49606);
and UO_3376 (O_3376,N_49590,N_49569);
nor UO_3377 (O_3377,N_49831,N_49473);
or UO_3378 (O_3378,N_49366,N_49358);
and UO_3379 (O_3379,N_49558,N_49685);
or UO_3380 (O_3380,N_49654,N_49866);
and UO_3381 (O_3381,N_49361,N_49898);
nand UO_3382 (O_3382,N_49154,N_49978);
and UO_3383 (O_3383,N_49959,N_49459);
nor UO_3384 (O_3384,N_49370,N_49340);
nor UO_3385 (O_3385,N_49426,N_49275);
nor UO_3386 (O_3386,N_49827,N_49898);
and UO_3387 (O_3387,N_49716,N_49390);
nor UO_3388 (O_3388,N_49202,N_49802);
xnor UO_3389 (O_3389,N_49781,N_49551);
xor UO_3390 (O_3390,N_49117,N_49033);
and UO_3391 (O_3391,N_49917,N_49837);
and UO_3392 (O_3392,N_49320,N_49087);
xor UO_3393 (O_3393,N_49702,N_49154);
nor UO_3394 (O_3394,N_49040,N_49466);
or UO_3395 (O_3395,N_49419,N_49802);
and UO_3396 (O_3396,N_49827,N_49789);
xor UO_3397 (O_3397,N_49108,N_49354);
nor UO_3398 (O_3398,N_49951,N_49659);
nor UO_3399 (O_3399,N_49510,N_49575);
or UO_3400 (O_3400,N_49928,N_49183);
xnor UO_3401 (O_3401,N_49926,N_49770);
and UO_3402 (O_3402,N_49210,N_49109);
and UO_3403 (O_3403,N_49957,N_49113);
and UO_3404 (O_3404,N_49828,N_49852);
xnor UO_3405 (O_3405,N_49806,N_49437);
or UO_3406 (O_3406,N_49471,N_49613);
nand UO_3407 (O_3407,N_49070,N_49268);
nand UO_3408 (O_3408,N_49944,N_49701);
nor UO_3409 (O_3409,N_49910,N_49389);
nand UO_3410 (O_3410,N_49099,N_49110);
and UO_3411 (O_3411,N_49411,N_49131);
or UO_3412 (O_3412,N_49218,N_49462);
xnor UO_3413 (O_3413,N_49406,N_49711);
nand UO_3414 (O_3414,N_49598,N_49642);
nor UO_3415 (O_3415,N_49104,N_49031);
nor UO_3416 (O_3416,N_49954,N_49988);
or UO_3417 (O_3417,N_49296,N_49368);
or UO_3418 (O_3418,N_49881,N_49997);
nor UO_3419 (O_3419,N_49774,N_49900);
and UO_3420 (O_3420,N_49880,N_49240);
nor UO_3421 (O_3421,N_49701,N_49929);
or UO_3422 (O_3422,N_49341,N_49830);
and UO_3423 (O_3423,N_49474,N_49046);
nor UO_3424 (O_3424,N_49939,N_49314);
or UO_3425 (O_3425,N_49966,N_49908);
or UO_3426 (O_3426,N_49390,N_49317);
nand UO_3427 (O_3427,N_49576,N_49112);
or UO_3428 (O_3428,N_49323,N_49715);
or UO_3429 (O_3429,N_49219,N_49940);
xor UO_3430 (O_3430,N_49641,N_49711);
nor UO_3431 (O_3431,N_49683,N_49003);
nand UO_3432 (O_3432,N_49123,N_49738);
nand UO_3433 (O_3433,N_49597,N_49964);
nand UO_3434 (O_3434,N_49569,N_49370);
nor UO_3435 (O_3435,N_49883,N_49471);
or UO_3436 (O_3436,N_49902,N_49857);
and UO_3437 (O_3437,N_49767,N_49648);
and UO_3438 (O_3438,N_49132,N_49469);
or UO_3439 (O_3439,N_49094,N_49902);
or UO_3440 (O_3440,N_49605,N_49938);
nor UO_3441 (O_3441,N_49106,N_49003);
nand UO_3442 (O_3442,N_49609,N_49007);
nor UO_3443 (O_3443,N_49516,N_49162);
nor UO_3444 (O_3444,N_49860,N_49247);
xnor UO_3445 (O_3445,N_49529,N_49077);
xnor UO_3446 (O_3446,N_49829,N_49863);
nand UO_3447 (O_3447,N_49595,N_49375);
nand UO_3448 (O_3448,N_49475,N_49320);
xnor UO_3449 (O_3449,N_49039,N_49001);
nand UO_3450 (O_3450,N_49766,N_49027);
nand UO_3451 (O_3451,N_49973,N_49530);
and UO_3452 (O_3452,N_49365,N_49974);
xnor UO_3453 (O_3453,N_49332,N_49798);
xnor UO_3454 (O_3454,N_49723,N_49210);
xnor UO_3455 (O_3455,N_49080,N_49011);
or UO_3456 (O_3456,N_49904,N_49517);
xnor UO_3457 (O_3457,N_49447,N_49400);
nor UO_3458 (O_3458,N_49507,N_49920);
or UO_3459 (O_3459,N_49307,N_49331);
xor UO_3460 (O_3460,N_49266,N_49854);
nor UO_3461 (O_3461,N_49892,N_49846);
nor UO_3462 (O_3462,N_49069,N_49360);
and UO_3463 (O_3463,N_49375,N_49515);
nand UO_3464 (O_3464,N_49705,N_49302);
and UO_3465 (O_3465,N_49720,N_49894);
nand UO_3466 (O_3466,N_49613,N_49612);
and UO_3467 (O_3467,N_49816,N_49389);
nand UO_3468 (O_3468,N_49834,N_49560);
nor UO_3469 (O_3469,N_49641,N_49404);
nand UO_3470 (O_3470,N_49156,N_49955);
or UO_3471 (O_3471,N_49690,N_49193);
xor UO_3472 (O_3472,N_49609,N_49348);
and UO_3473 (O_3473,N_49152,N_49944);
nand UO_3474 (O_3474,N_49237,N_49740);
nand UO_3475 (O_3475,N_49860,N_49239);
nand UO_3476 (O_3476,N_49859,N_49561);
and UO_3477 (O_3477,N_49577,N_49803);
nand UO_3478 (O_3478,N_49687,N_49225);
and UO_3479 (O_3479,N_49952,N_49406);
nand UO_3480 (O_3480,N_49870,N_49798);
nor UO_3481 (O_3481,N_49388,N_49180);
or UO_3482 (O_3482,N_49949,N_49814);
and UO_3483 (O_3483,N_49371,N_49171);
and UO_3484 (O_3484,N_49431,N_49643);
nand UO_3485 (O_3485,N_49379,N_49025);
nand UO_3486 (O_3486,N_49926,N_49454);
nand UO_3487 (O_3487,N_49376,N_49088);
nor UO_3488 (O_3488,N_49029,N_49101);
nand UO_3489 (O_3489,N_49444,N_49091);
nand UO_3490 (O_3490,N_49027,N_49264);
nor UO_3491 (O_3491,N_49482,N_49374);
or UO_3492 (O_3492,N_49526,N_49977);
and UO_3493 (O_3493,N_49755,N_49857);
and UO_3494 (O_3494,N_49116,N_49569);
xnor UO_3495 (O_3495,N_49293,N_49717);
nor UO_3496 (O_3496,N_49160,N_49835);
nand UO_3497 (O_3497,N_49530,N_49878);
nand UO_3498 (O_3498,N_49049,N_49317);
and UO_3499 (O_3499,N_49536,N_49210);
or UO_3500 (O_3500,N_49484,N_49823);
or UO_3501 (O_3501,N_49047,N_49704);
nand UO_3502 (O_3502,N_49992,N_49278);
xor UO_3503 (O_3503,N_49695,N_49280);
nor UO_3504 (O_3504,N_49767,N_49495);
xnor UO_3505 (O_3505,N_49530,N_49194);
nand UO_3506 (O_3506,N_49098,N_49271);
or UO_3507 (O_3507,N_49753,N_49751);
nor UO_3508 (O_3508,N_49735,N_49862);
nand UO_3509 (O_3509,N_49701,N_49882);
and UO_3510 (O_3510,N_49200,N_49166);
and UO_3511 (O_3511,N_49218,N_49020);
and UO_3512 (O_3512,N_49620,N_49729);
nor UO_3513 (O_3513,N_49601,N_49391);
xnor UO_3514 (O_3514,N_49637,N_49658);
or UO_3515 (O_3515,N_49255,N_49005);
or UO_3516 (O_3516,N_49033,N_49768);
nand UO_3517 (O_3517,N_49605,N_49145);
or UO_3518 (O_3518,N_49826,N_49128);
xnor UO_3519 (O_3519,N_49480,N_49595);
or UO_3520 (O_3520,N_49877,N_49177);
nand UO_3521 (O_3521,N_49621,N_49108);
nor UO_3522 (O_3522,N_49672,N_49948);
and UO_3523 (O_3523,N_49388,N_49126);
or UO_3524 (O_3524,N_49181,N_49966);
nand UO_3525 (O_3525,N_49716,N_49673);
or UO_3526 (O_3526,N_49301,N_49220);
and UO_3527 (O_3527,N_49620,N_49760);
and UO_3528 (O_3528,N_49906,N_49581);
and UO_3529 (O_3529,N_49153,N_49447);
nor UO_3530 (O_3530,N_49900,N_49756);
and UO_3531 (O_3531,N_49747,N_49958);
or UO_3532 (O_3532,N_49509,N_49218);
and UO_3533 (O_3533,N_49995,N_49467);
xor UO_3534 (O_3534,N_49143,N_49685);
xnor UO_3535 (O_3535,N_49772,N_49745);
or UO_3536 (O_3536,N_49952,N_49852);
nor UO_3537 (O_3537,N_49806,N_49333);
nor UO_3538 (O_3538,N_49159,N_49088);
nor UO_3539 (O_3539,N_49247,N_49406);
xor UO_3540 (O_3540,N_49272,N_49483);
xor UO_3541 (O_3541,N_49822,N_49704);
and UO_3542 (O_3542,N_49621,N_49470);
nand UO_3543 (O_3543,N_49001,N_49975);
nor UO_3544 (O_3544,N_49016,N_49453);
xor UO_3545 (O_3545,N_49947,N_49909);
nand UO_3546 (O_3546,N_49436,N_49737);
xor UO_3547 (O_3547,N_49792,N_49232);
nor UO_3548 (O_3548,N_49797,N_49011);
xor UO_3549 (O_3549,N_49106,N_49122);
or UO_3550 (O_3550,N_49050,N_49454);
nand UO_3551 (O_3551,N_49965,N_49808);
nand UO_3552 (O_3552,N_49004,N_49734);
nor UO_3553 (O_3553,N_49486,N_49375);
or UO_3554 (O_3554,N_49987,N_49811);
xor UO_3555 (O_3555,N_49802,N_49643);
nand UO_3556 (O_3556,N_49654,N_49696);
xnor UO_3557 (O_3557,N_49049,N_49397);
nand UO_3558 (O_3558,N_49502,N_49135);
and UO_3559 (O_3559,N_49947,N_49993);
xnor UO_3560 (O_3560,N_49448,N_49046);
or UO_3561 (O_3561,N_49236,N_49534);
xnor UO_3562 (O_3562,N_49462,N_49211);
nor UO_3563 (O_3563,N_49556,N_49354);
nor UO_3564 (O_3564,N_49058,N_49343);
nand UO_3565 (O_3565,N_49554,N_49784);
xor UO_3566 (O_3566,N_49949,N_49996);
or UO_3567 (O_3567,N_49422,N_49590);
xnor UO_3568 (O_3568,N_49464,N_49105);
nand UO_3569 (O_3569,N_49055,N_49000);
or UO_3570 (O_3570,N_49704,N_49121);
nand UO_3571 (O_3571,N_49170,N_49933);
nor UO_3572 (O_3572,N_49891,N_49798);
nand UO_3573 (O_3573,N_49932,N_49579);
nor UO_3574 (O_3574,N_49739,N_49511);
nand UO_3575 (O_3575,N_49502,N_49565);
and UO_3576 (O_3576,N_49544,N_49064);
nand UO_3577 (O_3577,N_49450,N_49626);
nand UO_3578 (O_3578,N_49764,N_49397);
nand UO_3579 (O_3579,N_49295,N_49187);
and UO_3580 (O_3580,N_49306,N_49502);
xor UO_3581 (O_3581,N_49413,N_49275);
and UO_3582 (O_3582,N_49184,N_49768);
xnor UO_3583 (O_3583,N_49373,N_49314);
xnor UO_3584 (O_3584,N_49625,N_49913);
and UO_3585 (O_3585,N_49906,N_49636);
nand UO_3586 (O_3586,N_49489,N_49501);
nand UO_3587 (O_3587,N_49323,N_49655);
nand UO_3588 (O_3588,N_49854,N_49181);
xnor UO_3589 (O_3589,N_49596,N_49827);
or UO_3590 (O_3590,N_49635,N_49338);
nor UO_3591 (O_3591,N_49434,N_49446);
and UO_3592 (O_3592,N_49064,N_49950);
and UO_3593 (O_3593,N_49694,N_49534);
nand UO_3594 (O_3594,N_49298,N_49401);
or UO_3595 (O_3595,N_49482,N_49708);
and UO_3596 (O_3596,N_49113,N_49940);
nand UO_3597 (O_3597,N_49469,N_49930);
and UO_3598 (O_3598,N_49392,N_49085);
and UO_3599 (O_3599,N_49886,N_49945);
nand UO_3600 (O_3600,N_49774,N_49914);
nand UO_3601 (O_3601,N_49190,N_49852);
and UO_3602 (O_3602,N_49828,N_49482);
or UO_3603 (O_3603,N_49049,N_49749);
or UO_3604 (O_3604,N_49540,N_49985);
nand UO_3605 (O_3605,N_49251,N_49529);
nand UO_3606 (O_3606,N_49742,N_49606);
and UO_3607 (O_3607,N_49489,N_49681);
nor UO_3608 (O_3608,N_49141,N_49481);
xor UO_3609 (O_3609,N_49836,N_49064);
and UO_3610 (O_3610,N_49258,N_49371);
or UO_3611 (O_3611,N_49226,N_49263);
or UO_3612 (O_3612,N_49591,N_49102);
or UO_3613 (O_3613,N_49188,N_49804);
nand UO_3614 (O_3614,N_49476,N_49480);
nand UO_3615 (O_3615,N_49072,N_49387);
nor UO_3616 (O_3616,N_49440,N_49963);
nand UO_3617 (O_3617,N_49239,N_49207);
xnor UO_3618 (O_3618,N_49946,N_49491);
and UO_3619 (O_3619,N_49062,N_49420);
nand UO_3620 (O_3620,N_49237,N_49650);
nor UO_3621 (O_3621,N_49734,N_49093);
nor UO_3622 (O_3622,N_49263,N_49828);
and UO_3623 (O_3623,N_49571,N_49823);
and UO_3624 (O_3624,N_49050,N_49392);
and UO_3625 (O_3625,N_49688,N_49631);
xor UO_3626 (O_3626,N_49540,N_49868);
and UO_3627 (O_3627,N_49752,N_49202);
xnor UO_3628 (O_3628,N_49932,N_49603);
nand UO_3629 (O_3629,N_49829,N_49115);
and UO_3630 (O_3630,N_49257,N_49580);
nor UO_3631 (O_3631,N_49904,N_49097);
nor UO_3632 (O_3632,N_49357,N_49599);
nor UO_3633 (O_3633,N_49185,N_49260);
or UO_3634 (O_3634,N_49092,N_49144);
nand UO_3635 (O_3635,N_49471,N_49705);
and UO_3636 (O_3636,N_49297,N_49608);
or UO_3637 (O_3637,N_49976,N_49148);
nor UO_3638 (O_3638,N_49291,N_49030);
nor UO_3639 (O_3639,N_49401,N_49969);
nand UO_3640 (O_3640,N_49899,N_49531);
xor UO_3641 (O_3641,N_49530,N_49138);
and UO_3642 (O_3642,N_49705,N_49797);
or UO_3643 (O_3643,N_49663,N_49278);
nor UO_3644 (O_3644,N_49965,N_49325);
or UO_3645 (O_3645,N_49115,N_49593);
nand UO_3646 (O_3646,N_49253,N_49443);
nand UO_3647 (O_3647,N_49745,N_49311);
xnor UO_3648 (O_3648,N_49196,N_49635);
xnor UO_3649 (O_3649,N_49058,N_49846);
nor UO_3650 (O_3650,N_49691,N_49473);
or UO_3651 (O_3651,N_49910,N_49492);
nor UO_3652 (O_3652,N_49575,N_49340);
xnor UO_3653 (O_3653,N_49925,N_49519);
nor UO_3654 (O_3654,N_49653,N_49967);
nor UO_3655 (O_3655,N_49537,N_49513);
nor UO_3656 (O_3656,N_49895,N_49934);
and UO_3657 (O_3657,N_49749,N_49216);
or UO_3658 (O_3658,N_49533,N_49473);
nor UO_3659 (O_3659,N_49705,N_49176);
xor UO_3660 (O_3660,N_49447,N_49467);
and UO_3661 (O_3661,N_49977,N_49996);
nand UO_3662 (O_3662,N_49138,N_49702);
nand UO_3663 (O_3663,N_49756,N_49146);
nor UO_3664 (O_3664,N_49801,N_49112);
nand UO_3665 (O_3665,N_49289,N_49802);
xor UO_3666 (O_3666,N_49011,N_49889);
or UO_3667 (O_3667,N_49137,N_49367);
or UO_3668 (O_3668,N_49459,N_49248);
or UO_3669 (O_3669,N_49806,N_49515);
xor UO_3670 (O_3670,N_49790,N_49282);
nor UO_3671 (O_3671,N_49783,N_49310);
and UO_3672 (O_3672,N_49212,N_49543);
xnor UO_3673 (O_3673,N_49557,N_49787);
or UO_3674 (O_3674,N_49870,N_49506);
nand UO_3675 (O_3675,N_49257,N_49371);
nand UO_3676 (O_3676,N_49392,N_49028);
and UO_3677 (O_3677,N_49791,N_49895);
nand UO_3678 (O_3678,N_49622,N_49880);
xor UO_3679 (O_3679,N_49335,N_49111);
and UO_3680 (O_3680,N_49785,N_49613);
nor UO_3681 (O_3681,N_49469,N_49386);
and UO_3682 (O_3682,N_49027,N_49256);
xor UO_3683 (O_3683,N_49074,N_49206);
nor UO_3684 (O_3684,N_49728,N_49012);
or UO_3685 (O_3685,N_49097,N_49804);
and UO_3686 (O_3686,N_49062,N_49135);
and UO_3687 (O_3687,N_49262,N_49386);
xnor UO_3688 (O_3688,N_49183,N_49887);
nor UO_3689 (O_3689,N_49944,N_49427);
xor UO_3690 (O_3690,N_49816,N_49135);
xnor UO_3691 (O_3691,N_49113,N_49383);
nor UO_3692 (O_3692,N_49245,N_49782);
and UO_3693 (O_3693,N_49838,N_49768);
xnor UO_3694 (O_3694,N_49704,N_49512);
nand UO_3695 (O_3695,N_49726,N_49146);
xor UO_3696 (O_3696,N_49222,N_49556);
or UO_3697 (O_3697,N_49807,N_49812);
nand UO_3698 (O_3698,N_49358,N_49845);
and UO_3699 (O_3699,N_49450,N_49761);
nand UO_3700 (O_3700,N_49696,N_49857);
xnor UO_3701 (O_3701,N_49764,N_49895);
nor UO_3702 (O_3702,N_49033,N_49159);
and UO_3703 (O_3703,N_49895,N_49705);
nor UO_3704 (O_3704,N_49114,N_49725);
or UO_3705 (O_3705,N_49053,N_49102);
nor UO_3706 (O_3706,N_49989,N_49619);
or UO_3707 (O_3707,N_49832,N_49461);
xnor UO_3708 (O_3708,N_49433,N_49573);
nand UO_3709 (O_3709,N_49550,N_49229);
xnor UO_3710 (O_3710,N_49379,N_49512);
and UO_3711 (O_3711,N_49596,N_49266);
or UO_3712 (O_3712,N_49362,N_49429);
and UO_3713 (O_3713,N_49002,N_49080);
nor UO_3714 (O_3714,N_49881,N_49816);
nand UO_3715 (O_3715,N_49053,N_49538);
nor UO_3716 (O_3716,N_49697,N_49478);
and UO_3717 (O_3717,N_49405,N_49244);
xnor UO_3718 (O_3718,N_49942,N_49055);
or UO_3719 (O_3719,N_49134,N_49373);
nand UO_3720 (O_3720,N_49636,N_49359);
nand UO_3721 (O_3721,N_49853,N_49365);
or UO_3722 (O_3722,N_49638,N_49859);
and UO_3723 (O_3723,N_49367,N_49537);
xor UO_3724 (O_3724,N_49930,N_49843);
xor UO_3725 (O_3725,N_49090,N_49875);
or UO_3726 (O_3726,N_49615,N_49534);
or UO_3727 (O_3727,N_49286,N_49398);
nand UO_3728 (O_3728,N_49611,N_49804);
and UO_3729 (O_3729,N_49470,N_49270);
xnor UO_3730 (O_3730,N_49287,N_49033);
and UO_3731 (O_3731,N_49515,N_49150);
nor UO_3732 (O_3732,N_49410,N_49456);
nor UO_3733 (O_3733,N_49297,N_49128);
xnor UO_3734 (O_3734,N_49798,N_49946);
nand UO_3735 (O_3735,N_49963,N_49702);
nand UO_3736 (O_3736,N_49561,N_49083);
xnor UO_3737 (O_3737,N_49436,N_49564);
xor UO_3738 (O_3738,N_49911,N_49983);
and UO_3739 (O_3739,N_49670,N_49179);
xnor UO_3740 (O_3740,N_49819,N_49364);
or UO_3741 (O_3741,N_49395,N_49088);
nand UO_3742 (O_3742,N_49525,N_49665);
and UO_3743 (O_3743,N_49532,N_49440);
nand UO_3744 (O_3744,N_49762,N_49382);
and UO_3745 (O_3745,N_49569,N_49251);
or UO_3746 (O_3746,N_49975,N_49536);
xnor UO_3747 (O_3747,N_49434,N_49018);
xor UO_3748 (O_3748,N_49816,N_49296);
or UO_3749 (O_3749,N_49087,N_49277);
nand UO_3750 (O_3750,N_49412,N_49499);
or UO_3751 (O_3751,N_49881,N_49738);
nand UO_3752 (O_3752,N_49100,N_49820);
xnor UO_3753 (O_3753,N_49176,N_49018);
nand UO_3754 (O_3754,N_49921,N_49159);
nand UO_3755 (O_3755,N_49597,N_49926);
or UO_3756 (O_3756,N_49431,N_49653);
nor UO_3757 (O_3757,N_49887,N_49735);
and UO_3758 (O_3758,N_49997,N_49332);
and UO_3759 (O_3759,N_49631,N_49853);
and UO_3760 (O_3760,N_49318,N_49413);
nand UO_3761 (O_3761,N_49126,N_49841);
or UO_3762 (O_3762,N_49281,N_49141);
nand UO_3763 (O_3763,N_49423,N_49171);
nand UO_3764 (O_3764,N_49842,N_49118);
or UO_3765 (O_3765,N_49429,N_49214);
or UO_3766 (O_3766,N_49427,N_49949);
xnor UO_3767 (O_3767,N_49969,N_49061);
xor UO_3768 (O_3768,N_49333,N_49819);
or UO_3769 (O_3769,N_49522,N_49169);
xnor UO_3770 (O_3770,N_49019,N_49741);
or UO_3771 (O_3771,N_49235,N_49368);
nor UO_3772 (O_3772,N_49877,N_49932);
nand UO_3773 (O_3773,N_49410,N_49895);
nor UO_3774 (O_3774,N_49531,N_49782);
and UO_3775 (O_3775,N_49299,N_49203);
or UO_3776 (O_3776,N_49244,N_49809);
nor UO_3777 (O_3777,N_49617,N_49420);
nand UO_3778 (O_3778,N_49795,N_49198);
nand UO_3779 (O_3779,N_49457,N_49106);
nor UO_3780 (O_3780,N_49307,N_49513);
and UO_3781 (O_3781,N_49409,N_49125);
or UO_3782 (O_3782,N_49014,N_49487);
xor UO_3783 (O_3783,N_49232,N_49071);
xnor UO_3784 (O_3784,N_49940,N_49741);
nor UO_3785 (O_3785,N_49562,N_49140);
xor UO_3786 (O_3786,N_49105,N_49399);
nor UO_3787 (O_3787,N_49316,N_49542);
or UO_3788 (O_3788,N_49586,N_49106);
or UO_3789 (O_3789,N_49625,N_49212);
xnor UO_3790 (O_3790,N_49076,N_49400);
xor UO_3791 (O_3791,N_49031,N_49690);
xnor UO_3792 (O_3792,N_49447,N_49452);
or UO_3793 (O_3793,N_49400,N_49311);
or UO_3794 (O_3794,N_49774,N_49704);
nand UO_3795 (O_3795,N_49832,N_49786);
or UO_3796 (O_3796,N_49901,N_49957);
xor UO_3797 (O_3797,N_49568,N_49927);
xnor UO_3798 (O_3798,N_49942,N_49031);
xnor UO_3799 (O_3799,N_49919,N_49170);
nand UO_3800 (O_3800,N_49750,N_49937);
nand UO_3801 (O_3801,N_49145,N_49210);
or UO_3802 (O_3802,N_49892,N_49651);
nand UO_3803 (O_3803,N_49409,N_49110);
xor UO_3804 (O_3804,N_49445,N_49554);
and UO_3805 (O_3805,N_49720,N_49114);
xor UO_3806 (O_3806,N_49668,N_49897);
or UO_3807 (O_3807,N_49555,N_49078);
nor UO_3808 (O_3808,N_49573,N_49596);
xnor UO_3809 (O_3809,N_49175,N_49149);
xor UO_3810 (O_3810,N_49997,N_49279);
or UO_3811 (O_3811,N_49835,N_49606);
and UO_3812 (O_3812,N_49273,N_49590);
and UO_3813 (O_3813,N_49502,N_49380);
and UO_3814 (O_3814,N_49953,N_49740);
or UO_3815 (O_3815,N_49875,N_49662);
nor UO_3816 (O_3816,N_49144,N_49835);
nor UO_3817 (O_3817,N_49317,N_49235);
and UO_3818 (O_3818,N_49036,N_49923);
nor UO_3819 (O_3819,N_49728,N_49864);
and UO_3820 (O_3820,N_49923,N_49732);
nand UO_3821 (O_3821,N_49227,N_49415);
nor UO_3822 (O_3822,N_49324,N_49999);
nor UO_3823 (O_3823,N_49168,N_49563);
nand UO_3824 (O_3824,N_49751,N_49963);
or UO_3825 (O_3825,N_49549,N_49776);
xor UO_3826 (O_3826,N_49865,N_49845);
nand UO_3827 (O_3827,N_49712,N_49899);
nor UO_3828 (O_3828,N_49015,N_49634);
nor UO_3829 (O_3829,N_49291,N_49091);
nor UO_3830 (O_3830,N_49010,N_49761);
or UO_3831 (O_3831,N_49851,N_49014);
nand UO_3832 (O_3832,N_49462,N_49729);
xor UO_3833 (O_3833,N_49265,N_49958);
or UO_3834 (O_3834,N_49809,N_49487);
nand UO_3835 (O_3835,N_49547,N_49484);
and UO_3836 (O_3836,N_49748,N_49795);
xnor UO_3837 (O_3837,N_49361,N_49175);
nand UO_3838 (O_3838,N_49325,N_49390);
nand UO_3839 (O_3839,N_49864,N_49754);
xnor UO_3840 (O_3840,N_49892,N_49119);
or UO_3841 (O_3841,N_49891,N_49000);
xor UO_3842 (O_3842,N_49874,N_49978);
xor UO_3843 (O_3843,N_49818,N_49057);
nand UO_3844 (O_3844,N_49298,N_49021);
or UO_3845 (O_3845,N_49623,N_49898);
or UO_3846 (O_3846,N_49282,N_49382);
and UO_3847 (O_3847,N_49260,N_49691);
xor UO_3848 (O_3848,N_49766,N_49591);
nand UO_3849 (O_3849,N_49221,N_49268);
nor UO_3850 (O_3850,N_49626,N_49743);
xnor UO_3851 (O_3851,N_49174,N_49541);
xor UO_3852 (O_3852,N_49880,N_49491);
xor UO_3853 (O_3853,N_49523,N_49546);
nand UO_3854 (O_3854,N_49233,N_49268);
xor UO_3855 (O_3855,N_49661,N_49956);
nor UO_3856 (O_3856,N_49306,N_49002);
nor UO_3857 (O_3857,N_49743,N_49008);
or UO_3858 (O_3858,N_49329,N_49532);
nand UO_3859 (O_3859,N_49266,N_49264);
xnor UO_3860 (O_3860,N_49281,N_49135);
xnor UO_3861 (O_3861,N_49492,N_49260);
and UO_3862 (O_3862,N_49018,N_49649);
nand UO_3863 (O_3863,N_49548,N_49937);
or UO_3864 (O_3864,N_49574,N_49815);
and UO_3865 (O_3865,N_49905,N_49798);
xnor UO_3866 (O_3866,N_49011,N_49331);
and UO_3867 (O_3867,N_49972,N_49040);
xnor UO_3868 (O_3868,N_49938,N_49269);
nand UO_3869 (O_3869,N_49925,N_49736);
nor UO_3870 (O_3870,N_49312,N_49684);
and UO_3871 (O_3871,N_49851,N_49729);
nand UO_3872 (O_3872,N_49140,N_49066);
and UO_3873 (O_3873,N_49008,N_49195);
nand UO_3874 (O_3874,N_49022,N_49677);
and UO_3875 (O_3875,N_49292,N_49420);
nor UO_3876 (O_3876,N_49623,N_49677);
nor UO_3877 (O_3877,N_49511,N_49351);
or UO_3878 (O_3878,N_49761,N_49092);
nor UO_3879 (O_3879,N_49998,N_49480);
or UO_3880 (O_3880,N_49144,N_49106);
and UO_3881 (O_3881,N_49167,N_49193);
or UO_3882 (O_3882,N_49792,N_49647);
and UO_3883 (O_3883,N_49122,N_49819);
nor UO_3884 (O_3884,N_49255,N_49421);
or UO_3885 (O_3885,N_49071,N_49173);
or UO_3886 (O_3886,N_49333,N_49132);
and UO_3887 (O_3887,N_49458,N_49395);
nand UO_3888 (O_3888,N_49530,N_49772);
nor UO_3889 (O_3889,N_49576,N_49295);
or UO_3890 (O_3890,N_49497,N_49293);
xor UO_3891 (O_3891,N_49914,N_49477);
or UO_3892 (O_3892,N_49451,N_49747);
or UO_3893 (O_3893,N_49332,N_49645);
nor UO_3894 (O_3894,N_49032,N_49862);
nor UO_3895 (O_3895,N_49540,N_49729);
xnor UO_3896 (O_3896,N_49897,N_49723);
and UO_3897 (O_3897,N_49967,N_49021);
xor UO_3898 (O_3898,N_49994,N_49434);
or UO_3899 (O_3899,N_49204,N_49815);
nor UO_3900 (O_3900,N_49323,N_49646);
xnor UO_3901 (O_3901,N_49226,N_49440);
or UO_3902 (O_3902,N_49569,N_49075);
nor UO_3903 (O_3903,N_49546,N_49767);
and UO_3904 (O_3904,N_49337,N_49837);
or UO_3905 (O_3905,N_49172,N_49454);
nand UO_3906 (O_3906,N_49155,N_49947);
nor UO_3907 (O_3907,N_49569,N_49438);
or UO_3908 (O_3908,N_49652,N_49725);
nand UO_3909 (O_3909,N_49187,N_49907);
xor UO_3910 (O_3910,N_49802,N_49899);
nand UO_3911 (O_3911,N_49307,N_49902);
or UO_3912 (O_3912,N_49901,N_49818);
and UO_3913 (O_3913,N_49262,N_49973);
xnor UO_3914 (O_3914,N_49440,N_49640);
xor UO_3915 (O_3915,N_49224,N_49537);
and UO_3916 (O_3916,N_49909,N_49439);
nand UO_3917 (O_3917,N_49516,N_49985);
nand UO_3918 (O_3918,N_49643,N_49606);
xor UO_3919 (O_3919,N_49654,N_49065);
and UO_3920 (O_3920,N_49552,N_49988);
xnor UO_3921 (O_3921,N_49300,N_49918);
and UO_3922 (O_3922,N_49884,N_49071);
or UO_3923 (O_3923,N_49181,N_49192);
and UO_3924 (O_3924,N_49214,N_49121);
nand UO_3925 (O_3925,N_49061,N_49291);
xnor UO_3926 (O_3926,N_49856,N_49843);
nor UO_3927 (O_3927,N_49634,N_49811);
or UO_3928 (O_3928,N_49513,N_49405);
nand UO_3929 (O_3929,N_49642,N_49011);
nor UO_3930 (O_3930,N_49961,N_49550);
nor UO_3931 (O_3931,N_49281,N_49630);
nand UO_3932 (O_3932,N_49333,N_49463);
xnor UO_3933 (O_3933,N_49275,N_49571);
and UO_3934 (O_3934,N_49478,N_49841);
nor UO_3935 (O_3935,N_49624,N_49839);
xnor UO_3936 (O_3936,N_49099,N_49268);
nand UO_3937 (O_3937,N_49522,N_49299);
and UO_3938 (O_3938,N_49953,N_49993);
xnor UO_3939 (O_3939,N_49540,N_49310);
xnor UO_3940 (O_3940,N_49027,N_49870);
and UO_3941 (O_3941,N_49868,N_49599);
or UO_3942 (O_3942,N_49275,N_49897);
and UO_3943 (O_3943,N_49188,N_49954);
nand UO_3944 (O_3944,N_49054,N_49317);
or UO_3945 (O_3945,N_49147,N_49874);
or UO_3946 (O_3946,N_49195,N_49658);
and UO_3947 (O_3947,N_49505,N_49792);
nand UO_3948 (O_3948,N_49984,N_49958);
nor UO_3949 (O_3949,N_49422,N_49082);
and UO_3950 (O_3950,N_49380,N_49839);
and UO_3951 (O_3951,N_49656,N_49163);
xor UO_3952 (O_3952,N_49676,N_49869);
xnor UO_3953 (O_3953,N_49269,N_49596);
and UO_3954 (O_3954,N_49575,N_49587);
nor UO_3955 (O_3955,N_49676,N_49088);
nand UO_3956 (O_3956,N_49103,N_49955);
or UO_3957 (O_3957,N_49918,N_49972);
xor UO_3958 (O_3958,N_49331,N_49280);
nor UO_3959 (O_3959,N_49232,N_49843);
nand UO_3960 (O_3960,N_49738,N_49989);
nand UO_3961 (O_3961,N_49140,N_49396);
or UO_3962 (O_3962,N_49450,N_49577);
xnor UO_3963 (O_3963,N_49541,N_49144);
or UO_3964 (O_3964,N_49742,N_49978);
and UO_3965 (O_3965,N_49711,N_49622);
xor UO_3966 (O_3966,N_49911,N_49077);
or UO_3967 (O_3967,N_49852,N_49158);
nor UO_3968 (O_3968,N_49329,N_49709);
and UO_3969 (O_3969,N_49324,N_49267);
nand UO_3970 (O_3970,N_49180,N_49603);
nand UO_3971 (O_3971,N_49941,N_49930);
or UO_3972 (O_3972,N_49463,N_49905);
and UO_3973 (O_3973,N_49863,N_49679);
nor UO_3974 (O_3974,N_49618,N_49603);
nand UO_3975 (O_3975,N_49898,N_49604);
and UO_3976 (O_3976,N_49018,N_49333);
and UO_3977 (O_3977,N_49952,N_49940);
or UO_3978 (O_3978,N_49840,N_49600);
and UO_3979 (O_3979,N_49141,N_49417);
nand UO_3980 (O_3980,N_49649,N_49931);
xnor UO_3981 (O_3981,N_49742,N_49006);
nand UO_3982 (O_3982,N_49584,N_49851);
nor UO_3983 (O_3983,N_49894,N_49186);
and UO_3984 (O_3984,N_49362,N_49043);
xor UO_3985 (O_3985,N_49327,N_49544);
nor UO_3986 (O_3986,N_49201,N_49878);
nand UO_3987 (O_3987,N_49091,N_49089);
xnor UO_3988 (O_3988,N_49954,N_49867);
nor UO_3989 (O_3989,N_49340,N_49798);
xnor UO_3990 (O_3990,N_49058,N_49741);
nor UO_3991 (O_3991,N_49206,N_49368);
and UO_3992 (O_3992,N_49486,N_49945);
and UO_3993 (O_3993,N_49635,N_49936);
and UO_3994 (O_3994,N_49553,N_49438);
xor UO_3995 (O_3995,N_49493,N_49578);
or UO_3996 (O_3996,N_49373,N_49523);
or UO_3997 (O_3997,N_49648,N_49352);
and UO_3998 (O_3998,N_49764,N_49655);
nand UO_3999 (O_3999,N_49982,N_49523);
or UO_4000 (O_4000,N_49459,N_49131);
nand UO_4001 (O_4001,N_49250,N_49451);
nand UO_4002 (O_4002,N_49892,N_49567);
and UO_4003 (O_4003,N_49992,N_49605);
nor UO_4004 (O_4004,N_49342,N_49414);
xor UO_4005 (O_4005,N_49568,N_49432);
or UO_4006 (O_4006,N_49372,N_49205);
xnor UO_4007 (O_4007,N_49474,N_49460);
and UO_4008 (O_4008,N_49035,N_49719);
or UO_4009 (O_4009,N_49286,N_49647);
nor UO_4010 (O_4010,N_49261,N_49571);
or UO_4011 (O_4011,N_49009,N_49323);
nand UO_4012 (O_4012,N_49651,N_49710);
nor UO_4013 (O_4013,N_49342,N_49443);
or UO_4014 (O_4014,N_49991,N_49952);
nand UO_4015 (O_4015,N_49618,N_49015);
or UO_4016 (O_4016,N_49040,N_49909);
nand UO_4017 (O_4017,N_49012,N_49592);
or UO_4018 (O_4018,N_49880,N_49221);
nor UO_4019 (O_4019,N_49650,N_49402);
nand UO_4020 (O_4020,N_49346,N_49967);
and UO_4021 (O_4021,N_49384,N_49283);
nor UO_4022 (O_4022,N_49113,N_49664);
or UO_4023 (O_4023,N_49647,N_49153);
and UO_4024 (O_4024,N_49133,N_49803);
xor UO_4025 (O_4025,N_49778,N_49677);
xnor UO_4026 (O_4026,N_49681,N_49444);
or UO_4027 (O_4027,N_49542,N_49730);
nor UO_4028 (O_4028,N_49397,N_49583);
xor UO_4029 (O_4029,N_49476,N_49364);
or UO_4030 (O_4030,N_49239,N_49245);
nand UO_4031 (O_4031,N_49992,N_49016);
nor UO_4032 (O_4032,N_49527,N_49032);
or UO_4033 (O_4033,N_49706,N_49179);
xnor UO_4034 (O_4034,N_49988,N_49537);
or UO_4035 (O_4035,N_49061,N_49970);
or UO_4036 (O_4036,N_49795,N_49356);
nand UO_4037 (O_4037,N_49670,N_49357);
and UO_4038 (O_4038,N_49729,N_49274);
nand UO_4039 (O_4039,N_49135,N_49870);
nor UO_4040 (O_4040,N_49233,N_49458);
nor UO_4041 (O_4041,N_49473,N_49045);
nand UO_4042 (O_4042,N_49110,N_49794);
xor UO_4043 (O_4043,N_49479,N_49268);
nor UO_4044 (O_4044,N_49815,N_49944);
and UO_4045 (O_4045,N_49782,N_49770);
nor UO_4046 (O_4046,N_49573,N_49746);
or UO_4047 (O_4047,N_49397,N_49749);
and UO_4048 (O_4048,N_49299,N_49136);
and UO_4049 (O_4049,N_49925,N_49914);
nand UO_4050 (O_4050,N_49336,N_49430);
nor UO_4051 (O_4051,N_49820,N_49312);
nor UO_4052 (O_4052,N_49538,N_49605);
xor UO_4053 (O_4053,N_49180,N_49383);
or UO_4054 (O_4054,N_49360,N_49316);
nand UO_4055 (O_4055,N_49832,N_49803);
and UO_4056 (O_4056,N_49093,N_49559);
nor UO_4057 (O_4057,N_49161,N_49574);
and UO_4058 (O_4058,N_49159,N_49749);
nor UO_4059 (O_4059,N_49202,N_49930);
xor UO_4060 (O_4060,N_49947,N_49470);
or UO_4061 (O_4061,N_49801,N_49428);
xnor UO_4062 (O_4062,N_49490,N_49965);
or UO_4063 (O_4063,N_49581,N_49607);
nand UO_4064 (O_4064,N_49799,N_49003);
or UO_4065 (O_4065,N_49706,N_49653);
and UO_4066 (O_4066,N_49780,N_49430);
nand UO_4067 (O_4067,N_49586,N_49006);
and UO_4068 (O_4068,N_49935,N_49066);
or UO_4069 (O_4069,N_49820,N_49363);
or UO_4070 (O_4070,N_49563,N_49885);
nand UO_4071 (O_4071,N_49672,N_49842);
or UO_4072 (O_4072,N_49664,N_49413);
nor UO_4073 (O_4073,N_49350,N_49868);
or UO_4074 (O_4074,N_49377,N_49773);
and UO_4075 (O_4075,N_49748,N_49990);
and UO_4076 (O_4076,N_49012,N_49664);
and UO_4077 (O_4077,N_49248,N_49129);
and UO_4078 (O_4078,N_49151,N_49939);
xnor UO_4079 (O_4079,N_49052,N_49813);
nor UO_4080 (O_4080,N_49866,N_49581);
xor UO_4081 (O_4081,N_49521,N_49748);
or UO_4082 (O_4082,N_49126,N_49174);
nand UO_4083 (O_4083,N_49412,N_49238);
xnor UO_4084 (O_4084,N_49742,N_49735);
nand UO_4085 (O_4085,N_49343,N_49546);
nand UO_4086 (O_4086,N_49011,N_49163);
and UO_4087 (O_4087,N_49852,N_49820);
and UO_4088 (O_4088,N_49600,N_49494);
or UO_4089 (O_4089,N_49461,N_49957);
and UO_4090 (O_4090,N_49382,N_49912);
and UO_4091 (O_4091,N_49818,N_49101);
nor UO_4092 (O_4092,N_49141,N_49277);
and UO_4093 (O_4093,N_49353,N_49514);
nor UO_4094 (O_4094,N_49963,N_49986);
xnor UO_4095 (O_4095,N_49453,N_49308);
and UO_4096 (O_4096,N_49115,N_49325);
and UO_4097 (O_4097,N_49060,N_49219);
nand UO_4098 (O_4098,N_49997,N_49941);
or UO_4099 (O_4099,N_49005,N_49159);
or UO_4100 (O_4100,N_49737,N_49831);
nor UO_4101 (O_4101,N_49841,N_49640);
or UO_4102 (O_4102,N_49260,N_49239);
nor UO_4103 (O_4103,N_49831,N_49950);
or UO_4104 (O_4104,N_49681,N_49258);
xnor UO_4105 (O_4105,N_49014,N_49627);
and UO_4106 (O_4106,N_49829,N_49410);
xor UO_4107 (O_4107,N_49962,N_49006);
and UO_4108 (O_4108,N_49264,N_49469);
or UO_4109 (O_4109,N_49872,N_49488);
and UO_4110 (O_4110,N_49228,N_49056);
or UO_4111 (O_4111,N_49998,N_49923);
and UO_4112 (O_4112,N_49234,N_49148);
or UO_4113 (O_4113,N_49732,N_49887);
nand UO_4114 (O_4114,N_49948,N_49356);
xor UO_4115 (O_4115,N_49785,N_49551);
nor UO_4116 (O_4116,N_49061,N_49971);
nand UO_4117 (O_4117,N_49999,N_49867);
and UO_4118 (O_4118,N_49277,N_49148);
nand UO_4119 (O_4119,N_49827,N_49357);
nor UO_4120 (O_4120,N_49395,N_49391);
xor UO_4121 (O_4121,N_49540,N_49915);
nand UO_4122 (O_4122,N_49639,N_49406);
and UO_4123 (O_4123,N_49536,N_49292);
xnor UO_4124 (O_4124,N_49053,N_49755);
nor UO_4125 (O_4125,N_49247,N_49375);
nor UO_4126 (O_4126,N_49541,N_49358);
nor UO_4127 (O_4127,N_49603,N_49037);
and UO_4128 (O_4128,N_49871,N_49733);
nor UO_4129 (O_4129,N_49809,N_49495);
nand UO_4130 (O_4130,N_49368,N_49957);
nor UO_4131 (O_4131,N_49492,N_49382);
or UO_4132 (O_4132,N_49369,N_49999);
or UO_4133 (O_4133,N_49829,N_49084);
and UO_4134 (O_4134,N_49150,N_49053);
or UO_4135 (O_4135,N_49911,N_49822);
or UO_4136 (O_4136,N_49145,N_49648);
nor UO_4137 (O_4137,N_49800,N_49137);
or UO_4138 (O_4138,N_49617,N_49656);
or UO_4139 (O_4139,N_49329,N_49192);
nand UO_4140 (O_4140,N_49340,N_49666);
xnor UO_4141 (O_4141,N_49487,N_49269);
and UO_4142 (O_4142,N_49331,N_49826);
and UO_4143 (O_4143,N_49956,N_49176);
xor UO_4144 (O_4144,N_49384,N_49888);
nand UO_4145 (O_4145,N_49496,N_49965);
xor UO_4146 (O_4146,N_49403,N_49464);
nor UO_4147 (O_4147,N_49284,N_49848);
nand UO_4148 (O_4148,N_49744,N_49946);
or UO_4149 (O_4149,N_49277,N_49259);
nor UO_4150 (O_4150,N_49235,N_49030);
and UO_4151 (O_4151,N_49589,N_49665);
nor UO_4152 (O_4152,N_49365,N_49142);
and UO_4153 (O_4153,N_49694,N_49706);
nand UO_4154 (O_4154,N_49210,N_49929);
xor UO_4155 (O_4155,N_49033,N_49717);
nor UO_4156 (O_4156,N_49338,N_49320);
nor UO_4157 (O_4157,N_49982,N_49373);
and UO_4158 (O_4158,N_49623,N_49500);
and UO_4159 (O_4159,N_49890,N_49416);
nor UO_4160 (O_4160,N_49499,N_49727);
and UO_4161 (O_4161,N_49665,N_49064);
nand UO_4162 (O_4162,N_49919,N_49770);
nor UO_4163 (O_4163,N_49038,N_49980);
or UO_4164 (O_4164,N_49959,N_49745);
nand UO_4165 (O_4165,N_49357,N_49325);
or UO_4166 (O_4166,N_49830,N_49716);
nand UO_4167 (O_4167,N_49323,N_49999);
nor UO_4168 (O_4168,N_49870,N_49363);
or UO_4169 (O_4169,N_49866,N_49821);
nor UO_4170 (O_4170,N_49018,N_49340);
nand UO_4171 (O_4171,N_49227,N_49416);
nor UO_4172 (O_4172,N_49858,N_49166);
or UO_4173 (O_4173,N_49333,N_49209);
or UO_4174 (O_4174,N_49391,N_49753);
xnor UO_4175 (O_4175,N_49360,N_49933);
nor UO_4176 (O_4176,N_49606,N_49070);
or UO_4177 (O_4177,N_49068,N_49450);
xor UO_4178 (O_4178,N_49970,N_49772);
or UO_4179 (O_4179,N_49460,N_49373);
xor UO_4180 (O_4180,N_49343,N_49661);
nand UO_4181 (O_4181,N_49657,N_49894);
nand UO_4182 (O_4182,N_49029,N_49726);
nand UO_4183 (O_4183,N_49323,N_49084);
and UO_4184 (O_4184,N_49968,N_49104);
xor UO_4185 (O_4185,N_49712,N_49240);
nor UO_4186 (O_4186,N_49869,N_49221);
xnor UO_4187 (O_4187,N_49415,N_49813);
nand UO_4188 (O_4188,N_49859,N_49058);
nor UO_4189 (O_4189,N_49357,N_49563);
or UO_4190 (O_4190,N_49694,N_49287);
and UO_4191 (O_4191,N_49179,N_49438);
nand UO_4192 (O_4192,N_49986,N_49998);
xnor UO_4193 (O_4193,N_49211,N_49099);
and UO_4194 (O_4194,N_49216,N_49268);
nand UO_4195 (O_4195,N_49142,N_49611);
xnor UO_4196 (O_4196,N_49518,N_49176);
and UO_4197 (O_4197,N_49086,N_49527);
or UO_4198 (O_4198,N_49506,N_49040);
nand UO_4199 (O_4199,N_49939,N_49029);
and UO_4200 (O_4200,N_49771,N_49936);
nor UO_4201 (O_4201,N_49267,N_49053);
nand UO_4202 (O_4202,N_49696,N_49104);
or UO_4203 (O_4203,N_49057,N_49972);
and UO_4204 (O_4204,N_49235,N_49398);
nand UO_4205 (O_4205,N_49883,N_49134);
and UO_4206 (O_4206,N_49469,N_49599);
nand UO_4207 (O_4207,N_49048,N_49540);
nor UO_4208 (O_4208,N_49354,N_49544);
or UO_4209 (O_4209,N_49589,N_49782);
nor UO_4210 (O_4210,N_49173,N_49029);
and UO_4211 (O_4211,N_49086,N_49471);
xor UO_4212 (O_4212,N_49929,N_49533);
nor UO_4213 (O_4213,N_49480,N_49147);
nor UO_4214 (O_4214,N_49230,N_49377);
or UO_4215 (O_4215,N_49601,N_49740);
or UO_4216 (O_4216,N_49484,N_49273);
nand UO_4217 (O_4217,N_49390,N_49429);
and UO_4218 (O_4218,N_49078,N_49149);
or UO_4219 (O_4219,N_49330,N_49181);
nand UO_4220 (O_4220,N_49008,N_49567);
nor UO_4221 (O_4221,N_49612,N_49604);
or UO_4222 (O_4222,N_49195,N_49592);
and UO_4223 (O_4223,N_49498,N_49265);
nor UO_4224 (O_4224,N_49681,N_49094);
nor UO_4225 (O_4225,N_49763,N_49531);
and UO_4226 (O_4226,N_49588,N_49205);
nand UO_4227 (O_4227,N_49100,N_49081);
or UO_4228 (O_4228,N_49126,N_49345);
nor UO_4229 (O_4229,N_49568,N_49852);
and UO_4230 (O_4230,N_49178,N_49909);
nand UO_4231 (O_4231,N_49721,N_49315);
nor UO_4232 (O_4232,N_49060,N_49604);
xor UO_4233 (O_4233,N_49638,N_49131);
nor UO_4234 (O_4234,N_49749,N_49995);
nor UO_4235 (O_4235,N_49600,N_49986);
or UO_4236 (O_4236,N_49872,N_49595);
nor UO_4237 (O_4237,N_49639,N_49420);
or UO_4238 (O_4238,N_49119,N_49987);
or UO_4239 (O_4239,N_49632,N_49102);
xor UO_4240 (O_4240,N_49207,N_49814);
and UO_4241 (O_4241,N_49524,N_49964);
xnor UO_4242 (O_4242,N_49707,N_49828);
xnor UO_4243 (O_4243,N_49016,N_49867);
nor UO_4244 (O_4244,N_49795,N_49362);
nor UO_4245 (O_4245,N_49318,N_49127);
nand UO_4246 (O_4246,N_49509,N_49194);
or UO_4247 (O_4247,N_49906,N_49314);
nand UO_4248 (O_4248,N_49720,N_49969);
nor UO_4249 (O_4249,N_49729,N_49824);
or UO_4250 (O_4250,N_49615,N_49230);
nand UO_4251 (O_4251,N_49561,N_49217);
and UO_4252 (O_4252,N_49536,N_49999);
nor UO_4253 (O_4253,N_49670,N_49914);
nand UO_4254 (O_4254,N_49902,N_49856);
nor UO_4255 (O_4255,N_49532,N_49628);
nor UO_4256 (O_4256,N_49066,N_49661);
xor UO_4257 (O_4257,N_49874,N_49607);
nor UO_4258 (O_4258,N_49590,N_49191);
or UO_4259 (O_4259,N_49652,N_49566);
or UO_4260 (O_4260,N_49033,N_49640);
nor UO_4261 (O_4261,N_49516,N_49885);
xor UO_4262 (O_4262,N_49868,N_49243);
nor UO_4263 (O_4263,N_49274,N_49346);
nor UO_4264 (O_4264,N_49248,N_49073);
nor UO_4265 (O_4265,N_49040,N_49880);
and UO_4266 (O_4266,N_49806,N_49166);
and UO_4267 (O_4267,N_49690,N_49021);
and UO_4268 (O_4268,N_49756,N_49852);
xnor UO_4269 (O_4269,N_49195,N_49609);
xor UO_4270 (O_4270,N_49076,N_49814);
or UO_4271 (O_4271,N_49129,N_49897);
xor UO_4272 (O_4272,N_49692,N_49024);
and UO_4273 (O_4273,N_49706,N_49089);
xor UO_4274 (O_4274,N_49783,N_49559);
xor UO_4275 (O_4275,N_49233,N_49542);
or UO_4276 (O_4276,N_49506,N_49120);
nor UO_4277 (O_4277,N_49597,N_49285);
or UO_4278 (O_4278,N_49764,N_49412);
xor UO_4279 (O_4279,N_49295,N_49357);
xor UO_4280 (O_4280,N_49247,N_49970);
and UO_4281 (O_4281,N_49400,N_49247);
nand UO_4282 (O_4282,N_49543,N_49901);
and UO_4283 (O_4283,N_49901,N_49886);
or UO_4284 (O_4284,N_49667,N_49779);
nor UO_4285 (O_4285,N_49619,N_49783);
nor UO_4286 (O_4286,N_49561,N_49218);
nand UO_4287 (O_4287,N_49022,N_49173);
nor UO_4288 (O_4288,N_49519,N_49402);
or UO_4289 (O_4289,N_49786,N_49650);
and UO_4290 (O_4290,N_49590,N_49243);
or UO_4291 (O_4291,N_49933,N_49940);
nor UO_4292 (O_4292,N_49913,N_49739);
nor UO_4293 (O_4293,N_49892,N_49012);
nor UO_4294 (O_4294,N_49912,N_49900);
xnor UO_4295 (O_4295,N_49532,N_49840);
xor UO_4296 (O_4296,N_49785,N_49591);
nand UO_4297 (O_4297,N_49374,N_49527);
nor UO_4298 (O_4298,N_49707,N_49713);
nand UO_4299 (O_4299,N_49203,N_49847);
nor UO_4300 (O_4300,N_49975,N_49289);
nor UO_4301 (O_4301,N_49943,N_49989);
and UO_4302 (O_4302,N_49115,N_49661);
and UO_4303 (O_4303,N_49498,N_49272);
nand UO_4304 (O_4304,N_49166,N_49569);
or UO_4305 (O_4305,N_49316,N_49813);
and UO_4306 (O_4306,N_49384,N_49139);
nand UO_4307 (O_4307,N_49959,N_49500);
xor UO_4308 (O_4308,N_49090,N_49015);
and UO_4309 (O_4309,N_49674,N_49382);
or UO_4310 (O_4310,N_49670,N_49581);
and UO_4311 (O_4311,N_49213,N_49635);
xnor UO_4312 (O_4312,N_49123,N_49355);
nand UO_4313 (O_4313,N_49411,N_49294);
or UO_4314 (O_4314,N_49243,N_49214);
nand UO_4315 (O_4315,N_49275,N_49477);
nand UO_4316 (O_4316,N_49698,N_49178);
nand UO_4317 (O_4317,N_49973,N_49579);
nand UO_4318 (O_4318,N_49070,N_49704);
and UO_4319 (O_4319,N_49796,N_49497);
xnor UO_4320 (O_4320,N_49203,N_49386);
xnor UO_4321 (O_4321,N_49194,N_49749);
and UO_4322 (O_4322,N_49648,N_49185);
xnor UO_4323 (O_4323,N_49852,N_49945);
or UO_4324 (O_4324,N_49509,N_49494);
or UO_4325 (O_4325,N_49327,N_49696);
nand UO_4326 (O_4326,N_49091,N_49304);
xor UO_4327 (O_4327,N_49851,N_49852);
nor UO_4328 (O_4328,N_49288,N_49210);
or UO_4329 (O_4329,N_49813,N_49683);
and UO_4330 (O_4330,N_49094,N_49434);
nand UO_4331 (O_4331,N_49689,N_49494);
nor UO_4332 (O_4332,N_49252,N_49113);
nor UO_4333 (O_4333,N_49773,N_49721);
or UO_4334 (O_4334,N_49092,N_49898);
or UO_4335 (O_4335,N_49724,N_49630);
or UO_4336 (O_4336,N_49280,N_49188);
or UO_4337 (O_4337,N_49562,N_49169);
nor UO_4338 (O_4338,N_49002,N_49691);
nand UO_4339 (O_4339,N_49863,N_49295);
nand UO_4340 (O_4340,N_49705,N_49929);
xnor UO_4341 (O_4341,N_49060,N_49304);
and UO_4342 (O_4342,N_49446,N_49084);
and UO_4343 (O_4343,N_49400,N_49369);
or UO_4344 (O_4344,N_49965,N_49270);
and UO_4345 (O_4345,N_49481,N_49985);
nand UO_4346 (O_4346,N_49939,N_49121);
xor UO_4347 (O_4347,N_49917,N_49665);
and UO_4348 (O_4348,N_49189,N_49241);
nor UO_4349 (O_4349,N_49461,N_49485);
or UO_4350 (O_4350,N_49010,N_49733);
xor UO_4351 (O_4351,N_49949,N_49636);
and UO_4352 (O_4352,N_49924,N_49454);
and UO_4353 (O_4353,N_49657,N_49239);
xnor UO_4354 (O_4354,N_49969,N_49914);
nor UO_4355 (O_4355,N_49881,N_49707);
xnor UO_4356 (O_4356,N_49369,N_49962);
nand UO_4357 (O_4357,N_49741,N_49633);
or UO_4358 (O_4358,N_49153,N_49949);
nor UO_4359 (O_4359,N_49699,N_49532);
nor UO_4360 (O_4360,N_49766,N_49341);
xor UO_4361 (O_4361,N_49139,N_49443);
nor UO_4362 (O_4362,N_49124,N_49229);
xnor UO_4363 (O_4363,N_49176,N_49327);
nor UO_4364 (O_4364,N_49842,N_49825);
xor UO_4365 (O_4365,N_49978,N_49937);
nand UO_4366 (O_4366,N_49909,N_49671);
and UO_4367 (O_4367,N_49989,N_49506);
and UO_4368 (O_4368,N_49999,N_49794);
nor UO_4369 (O_4369,N_49680,N_49063);
nand UO_4370 (O_4370,N_49785,N_49239);
nand UO_4371 (O_4371,N_49405,N_49863);
nor UO_4372 (O_4372,N_49353,N_49444);
and UO_4373 (O_4373,N_49918,N_49862);
and UO_4374 (O_4374,N_49759,N_49284);
and UO_4375 (O_4375,N_49192,N_49107);
or UO_4376 (O_4376,N_49548,N_49347);
and UO_4377 (O_4377,N_49076,N_49061);
and UO_4378 (O_4378,N_49714,N_49542);
or UO_4379 (O_4379,N_49865,N_49694);
and UO_4380 (O_4380,N_49482,N_49362);
xor UO_4381 (O_4381,N_49035,N_49867);
nor UO_4382 (O_4382,N_49754,N_49831);
or UO_4383 (O_4383,N_49598,N_49974);
xor UO_4384 (O_4384,N_49669,N_49736);
and UO_4385 (O_4385,N_49874,N_49286);
and UO_4386 (O_4386,N_49121,N_49935);
xnor UO_4387 (O_4387,N_49171,N_49201);
nor UO_4388 (O_4388,N_49549,N_49045);
xor UO_4389 (O_4389,N_49553,N_49316);
nand UO_4390 (O_4390,N_49528,N_49884);
nor UO_4391 (O_4391,N_49844,N_49162);
or UO_4392 (O_4392,N_49103,N_49838);
nor UO_4393 (O_4393,N_49929,N_49078);
nor UO_4394 (O_4394,N_49086,N_49123);
nor UO_4395 (O_4395,N_49178,N_49287);
or UO_4396 (O_4396,N_49288,N_49583);
xor UO_4397 (O_4397,N_49341,N_49718);
xor UO_4398 (O_4398,N_49081,N_49227);
xor UO_4399 (O_4399,N_49702,N_49557);
xor UO_4400 (O_4400,N_49028,N_49066);
and UO_4401 (O_4401,N_49705,N_49381);
and UO_4402 (O_4402,N_49196,N_49570);
and UO_4403 (O_4403,N_49849,N_49477);
nand UO_4404 (O_4404,N_49921,N_49540);
or UO_4405 (O_4405,N_49256,N_49531);
or UO_4406 (O_4406,N_49764,N_49292);
or UO_4407 (O_4407,N_49461,N_49554);
or UO_4408 (O_4408,N_49496,N_49473);
nand UO_4409 (O_4409,N_49311,N_49652);
xor UO_4410 (O_4410,N_49990,N_49084);
xor UO_4411 (O_4411,N_49918,N_49206);
nand UO_4412 (O_4412,N_49149,N_49157);
nand UO_4413 (O_4413,N_49431,N_49642);
xor UO_4414 (O_4414,N_49835,N_49538);
nand UO_4415 (O_4415,N_49842,N_49462);
nand UO_4416 (O_4416,N_49748,N_49250);
and UO_4417 (O_4417,N_49616,N_49198);
nor UO_4418 (O_4418,N_49684,N_49798);
and UO_4419 (O_4419,N_49578,N_49666);
nand UO_4420 (O_4420,N_49495,N_49010);
nand UO_4421 (O_4421,N_49020,N_49372);
xnor UO_4422 (O_4422,N_49865,N_49884);
nand UO_4423 (O_4423,N_49395,N_49838);
nor UO_4424 (O_4424,N_49861,N_49284);
and UO_4425 (O_4425,N_49732,N_49420);
xnor UO_4426 (O_4426,N_49847,N_49212);
or UO_4427 (O_4427,N_49442,N_49328);
and UO_4428 (O_4428,N_49954,N_49515);
and UO_4429 (O_4429,N_49168,N_49718);
nor UO_4430 (O_4430,N_49173,N_49583);
and UO_4431 (O_4431,N_49014,N_49526);
nor UO_4432 (O_4432,N_49707,N_49736);
and UO_4433 (O_4433,N_49948,N_49276);
nor UO_4434 (O_4434,N_49290,N_49004);
or UO_4435 (O_4435,N_49269,N_49306);
nand UO_4436 (O_4436,N_49027,N_49611);
or UO_4437 (O_4437,N_49911,N_49754);
and UO_4438 (O_4438,N_49351,N_49475);
nand UO_4439 (O_4439,N_49546,N_49698);
xor UO_4440 (O_4440,N_49990,N_49504);
nand UO_4441 (O_4441,N_49962,N_49695);
nor UO_4442 (O_4442,N_49930,N_49761);
nand UO_4443 (O_4443,N_49940,N_49674);
and UO_4444 (O_4444,N_49665,N_49954);
nor UO_4445 (O_4445,N_49343,N_49610);
or UO_4446 (O_4446,N_49299,N_49341);
and UO_4447 (O_4447,N_49659,N_49015);
nand UO_4448 (O_4448,N_49038,N_49104);
nor UO_4449 (O_4449,N_49449,N_49719);
or UO_4450 (O_4450,N_49864,N_49355);
or UO_4451 (O_4451,N_49534,N_49365);
or UO_4452 (O_4452,N_49070,N_49936);
nand UO_4453 (O_4453,N_49001,N_49808);
nor UO_4454 (O_4454,N_49918,N_49263);
and UO_4455 (O_4455,N_49546,N_49408);
xor UO_4456 (O_4456,N_49891,N_49823);
and UO_4457 (O_4457,N_49853,N_49700);
nor UO_4458 (O_4458,N_49689,N_49362);
nand UO_4459 (O_4459,N_49114,N_49462);
xnor UO_4460 (O_4460,N_49515,N_49836);
and UO_4461 (O_4461,N_49521,N_49615);
nand UO_4462 (O_4462,N_49787,N_49162);
or UO_4463 (O_4463,N_49296,N_49495);
or UO_4464 (O_4464,N_49612,N_49649);
nand UO_4465 (O_4465,N_49787,N_49292);
or UO_4466 (O_4466,N_49230,N_49770);
and UO_4467 (O_4467,N_49010,N_49481);
nor UO_4468 (O_4468,N_49293,N_49716);
xor UO_4469 (O_4469,N_49702,N_49057);
or UO_4470 (O_4470,N_49780,N_49137);
and UO_4471 (O_4471,N_49597,N_49069);
nor UO_4472 (O_4472,N_49103,N_49394);
nor UO_4473 (O_4473,N_49609,N_49787);
xnor UO_4474 (O_4474,N_49629,N_49615);
or UO_4475 (O_4475,N_49652,N_49910);
xor UO_4476 (O_4476,N_49370,N_49464);
and UO_4477 (O_4477,N_49480,N_49959);
nand UO_4478 (O_4478,N_49132,N_49786);
nand UO_4479 (O_4479,N_49963,N_49703);
and UO_4480 (O_4480,N_49965,N_49523);
nand UO_4481 (O_4481,N_49632,N_49062);
or UO_4482 (O_4482,N_49298,N_49694);
or UO_4483 (O_4483,N_49877,N_49089);
or UO_4484 (O_4484,N_49742,N_49887);
nand UO_4485 (O_4485,N_49976,N_49952);
and UO_4486 (O_4486,N_49068,N_49887);
and UO_4487 (O_4487,N_49801,N_49171);
nand UO_4488 (O_4488,N_49228,N_49399);
nand UO_4489 (O_4489,N_49415,N_49935);
nor UO_4490 (O_4490,N_49265,N_49319);
and UO_4491 (O_4491,N_49401,N_49553);
xnor UO_4492 (O_4492,N_49112,N_49301);
xnor UO_4493 (O_4493,N_49688,N_49397);
and UO_4494 (O_4494,N_49090,N_49711);
xnor UO_4495 (O_4495,N_49696,N_49343);
nand UO_4496 (O_4496,N_49250,N_49764);
and UO_4497 (O_4497,N_49064,N_49058);
nand UO_4498 (O_4498,N_49030,N_49263);
nand UO_4499 (O_4499,N_49031,N_49929);
nor UO_4500 (O_4500,N_49638,N_49215);
nand UO_4501 (O_4501,N_49753,N_49726);
and UO_4502 (O_4502,N_49856,N_49937);
nor UO_4503 (O_4503,N_49133,N_49723);
and UO_4504 (O_4504,N_49908,N_49150);
or UO_4505 (O_4505,N_49235,N_49727);
or UO_4506 (O_4506,N_49733,N_49524);
or UO_4507 (O_4507,N_49733,N_49082);
xor UO_4508 (O_4508,N_49983,N_49109);
nor UO_4509 (O_4509,N_49354,N_49251);
nand UO_4510 (O_4510,N_49474,N_49492);
nor UO_4511 (O_4511,N_49820,N_49512);
or UO_4512 (O_4512,N_49717,N_49486);
nand UO_4513 (O_4513,N_49137,N_49528);
nor UO_4514 (O_4514,N_49945,N_49104);
nor UO_4515 (O_4515,N_49066,N_49245);
and UO_4516 (O_4516,N_49349,N_49129);
xnor UO_4517 (O_4517,N_49367,N_49314);
xnor UO_4518 (O_4518,N_49859,N_49159);
or UO_4519 (O_4519,N_49744,N_49488);
nand UO_4520 (O_4520,N_49468,N_49120);
nor UO_4521 (O_4521,N_49878,N_49719);
nand UO_4522 (O_4522,N_49169,N_49496);
xnor UO_4523 (O_4523,N_49863,N_49903);
nand UO_4524 (O_4524,N_49541,N_49635);
and UO_4525 (O_4525,N_49961,N_49930);
xor UO_4526 (O_4526,N_49946,N_49338);
xor UO_4527 (O_4527,N_49356,N_49765);
and UO_4528 (O_4528,N_49524,N_49336);
and UO_4529 (O_4529,N_49823,N_49867);
nor UO_4530 (O_4530,N_49241,N_49308);
nand UO_4531 (O_4531,N_49454,N_49180);
xnor UO_4532 (O_4532,N_49667,N_49218);
and UO_4533 (O_4533,N_49071,N_49484);
xnor UO_4534 (O_4534,N_49623,N_49933);
xnor UO_4535 (O_4535,N_49655,N_49552);
nor UO_4536 (O_4536,N_49185,N_49403);
or UO_4537 (O_4537,N_49936,N_49482);
xnor UO_4538 (O_4538,N_49465,N_49849);
nor UO_4539 (O_4539,N_49677,N_49906);
nand UO_4540 (O_4540,N_49773,N_49551);
nand UO_4541 (O_4541,N_49477,N_49720);
and UO_4542 (O_4542,N_49887,N_49817);
or UO_4543 (O_4543,N_49566,N_49219);
nor UO_4544 (O_4544,N_49745,N_49808);
nor UO_4545 (O_4545,N_49092,N_49553);
nor UO_4546 (O_4546,N_49060,N_49794);
or UO_4547 (O_4547,N_49762,N_49545);
nor UO_4548 (O_4548,N_49289,N_49105);
or UO_4549 (O_4549,N_49129,N_49673);
or UO_4550 (O_4550,N_49685,N_49263);
or UO_4551 (O_4551,N_49270,N_49557);
and UO_4552 (O_4552,N_49788,N_49342);
xnor UO_4553 (O_4553,N_49663,N_49229);
nand UO_4554 (O_4554,N_49598,N_49340);
xnor UO_4555 (O_4555,N_49554,N_49803);
xnor UO_4556 (O_4556,N_49775,N_49375);
or UO_4557 (O_4557,N_49173,N_49469);
xor UO_4558 (O_4558,N_49167,N_49269);
nand UO_4559 (O_4559,N_49423,N_49947);
or UO_4560 (O_4560,N_49705,N_49435);
xnor UO_4561 (O_4561,N_49238,N_49539);
nor UO_4562 (O_4562,N_49910,N_49161);
nand UO_4563 (O_4563,N_49708,N_49021);
nor UO_4564 (O_4564,N_49411,N_49726);
xor UO_4565 (O_4565,N_49795,N_49241);
and UO_4566 (O_4566,N_49461,N_49471);
nor UO_4567 (O_4567,N_49140,N_49785);
nor UO_4568 (O_4568,N_49943,N_49806);
and UO_4569 (O_4569,N_49996,N_49810);
and UO_4570 (O_4570,N_49147,N_49786);
and UO_4571 (O_4571,N_49975,N_49543);
xnor UO_4572 (O_4572,N_49439,N_49897);
nor UO_4573 (O_4573,N_49748,N_49444);
xor UO_4574 (O_4574,N_49632,N_49614);
xnor UO_4575 (O_4575,N_49381,N_49153);
xor UO_4576 (O_4576,N_49883,N_49184);
and UO_4577 (O_4577,N_49625,N_49926);
nand UO_4578 (O_4578,N_49872,N_49417);
or UO_4579 (O_4579,N_49776,N_49704);
nor UO_4580 (O_4580,N_49873,N_49175);
xor UO_4581 (O_4581,N_49254,N_49883);
or UO_4582 (O_4582,N_49482,N_49704);
and UO_4583 (O_4583,N_49467,N_49255);
and UO_4584 (O_4584,N_49107,N_49386);
or UO_4585 (O_4585,N_49018,N_49959);
or UO_4586 (O_4586,N_49089,N_49626);
xnor UO_4587 (O_4587,N_49378,N_49036);
nand UO_4588 (O_4588,N_49195,N_49011);
or UO_4589 (O_4589,N_49864,N_49497);
xnor UO_4590 (O_4590,N_49066,N_49043);
and UO_4591 (O_4591,N_49628,N_49139);
and UO_4592 (O_4592,N_49104,N_49314);
or UO_4593 (O_4593,N_49469,N_49038);
xor UO_4594 (O_4594,N_49199,N_49927);
xnor UO_4595 (O_4595,N_49531,N_49400);
xor UO_4596 (O_4596,N_49033,N_49987);
nor UO_4597 (O_4597,N_49070,N_49347);
nand UO_4598 (O_4598,N_49272,N_49218);
or UO_4599 (O_4599,N_49172,N_49832);
or UO_4600 (O_4600,N_49488,N_49483);
or UO_4601 (O_4601,N_49267,N_49769);
nor UO_4602 (O_4602,N_49815,N_49892);
or UO_4603 (O_4603,N_49977,N_49927);
and UO_4604 (O_4604,N_49569,N_49537);
xnor UO_4605 (O_4605,N_49905,N_49018);
nand UO_4606 (O_4606,N_49140,N_49069);
nand UO_4607 (O_4607,N_49289,N_49472);
nand UO_4608 (O_4608,N_49343,N_49762);
nor UO_4609 (O_4609,N_49238,N_49836);
and UO_4610 (O_4610,N_49895,N_49296);
or UO_4611 (O_4611,N_49263,N_49991);
or UO_4612 (O_4612,N_49171,N_49998);
or UO_4613 (O_4613,N_49444,N_49980);
xnor UO_4614 (O_4614,N_49578,N_49511);
nor UO_4615 (O_4615,N_49325,N_49417);
and UO_4616 (O_4616,N_49959,N_49764);
or UO_4617 (O_4617,N_49446,N_49457);
and UO_4618 (O_4618,N_49617,N_49871);
nor UO_4619 (O_4619,N_49138,N_49991);
xnor UO_4620 (O_4620,N_49068,N_49804);
nand UO_4621 (O_4621,N_49422,N_49187);
nor UO_4622 (O_4622,N_49350,N_49015);
and UO_4623 (O_4623,N_49737,N_49126);
xor UO_4624 (O_4624,N_49809,N_49309);
or UO_4625 (O_4625,N_49681,N_49650);
nand UO_4626 (O_4626,N_49266,N_49772);
nor UO_4627 (O_4627,N_49238,N_49983);
or UO_4628 (O_4628,N_49286,N_49283);
or UO_4629 (O_4629,N_49517,N_49694);
nor UO_4630 (O_4630,N_49989,N_49838);
nand UO_4631 (O_4631,N_49301,N_49799);
nor UO_4632 (O_4632,N_49450,N_49043);
and UO_4633 (O_4633,N_49524,N_49067);
and UO_4634 (O_4634,N_49398,N_49387);
nor UO_4635 (O_4635,N_49232,N_49438);
nor UO_4636 (O_4636,N_49433,N_49959);
and UO_4637 (O_4637,N_49239,N_49241);
or UO_4638 (O_4638,N_49682,N_49955);
nor UO_4639 (O_4639,N_49003,N_49065);
nand UO_4640 (O_4640,N_49033,N_49816);
nand UO_4641 (O_4641,N_49592,N_49031);
xor UO_4642 (O_4642,N_49808,N_49544);
nand UO_4643 (O_4643,N_49537,N_49207);
xnor UO_4644 (O_4644,N_49354,N_49561);
nor UO_4645 (O_4645,N_49637,N_49512);
nor UO_4646 (O_4646,N_49874,N_49130);
nor UO_4647 (O_4647,N_49932,N_49938);
xor UO_4648 (O_4648,N_49190,N_49621);
or UO_4649 (O_4649,N_49326,N_49679);
or UO_4650 (O_4650,N_49675,N_49673);
and UO_4651 (O_4651,N_49969,N_49070);
nand UO_4652 (O_4652,N_49532,N_49359);
and UO_4653 (O_4653,N_49138,N_49713);
and UO_4654 (O_4654,N_49042,N_49430);
nor UO_4655 (O_4655,N_49811,N_49082);
nand UO_4656 (O_4656,N_49976,N_49680);
xor UO_4657 (O_4657,N_49906,N_49682);
xor UO_4658 (O_4658,N_49675,N_49378);
or UO_4659 (O_4659,N_49055,N_49761);
nand UO_4660 (O_4660,N_49410,N_49231);
xor UO_4661 (O_4661,N_49615,N_49538);
or UO_4662 (O_4662,N_49677,N_49309);
or UO_4663 (O_4663,N_49832,N_49196);
xor UO_4664 (O_4664,N_49448,N_49885);
nand UO_4665 (O_4665,N_49999,N_49950);
xor UO_4666 (O_4666,N_49230,N_49119);
and UO_4667 (O_4667,N_49473,N_49731);
nand UO_4668 (O_4668,N_49482,N_49657);
xnor UO_4669 (O_4669,N_49194,N_49027);
nor UO_4670 (O_4670,N_49035,N_49126);
and UO_4671 (O_4671,N_49204,N_49431);
or UO_4672 (O_4672,N_49783,N_49143);
and UO_4673 (O_4673,N_49079,N_49755);
or UO_4674 (O_4674,N_49478,N_49767);
nor UO_4675 (O_4675,N_49488,N_49504);
nand UO_4676 (O_4676,N_49378,N_49341);
and UO_4677 (O_4677,N_49552,N_49510);
and UO_4678 (O_4678,N_49364,N_49963);
and UO_4679 (O_4679,N_49372,N_49561);
xnor UO_4680 (O_4680,N_49375,N_49873);
and UO_4681 (O_4681,N_49810,N_49793);
xnor UO_4682 (O_4682,N_49440,N_49084);
nand UO_4683 (O_4683,N_49733,N_49490);
or UO_4684 (O_4684,N_49733,N_49977);
xor UO_4685 (O_4685,N_49888,N_49595);
nand UO_4686 (O_4686,N_49968,N_49128);
nor UO_4687 (O_4687,N_49200,N_49639);
and UO_4688 (O_4688,N_49760,N_49991);
or UO_4689 (O_4689,N_49082,N_49079);
and UO_4690 (O_4690,N_49102,N_49183);
nor UO_4691 (O_4691,N_49737,N_49984);
or UO_4692 (O_4692,N_49549,N_49614);
or UO_4693 (O_4693,N_49378,N_49913);
nor UO_4694 (O_4694,N_49613,N_49688);
nor UO_4695 (O_4695,N_49883,N_49357);
and UO_4696 (O_4696,N_49827,N_49004);
and UO_4697 (O_4697,N_49820,N_49382);
xor UO_4698 (O_4698,N_49253,N_49528);
xor UO_4699 (O_4699,N_49747,N_49954);
nor UO_4700 (O_4700,N_49232,N_49268);
nor UO_4701 (O_4701,N_49760,N_49019);
xor UO_4702 (O_4702,N_49367,N_49701);
nand UO_4703 (O_4703,N_49774,N_49647);
or UO_4704 (O_4704,N_49432,N_49653);
xor UO_4705 (O_4705,N_49062,N_49263);
nor UO_4706 (O_4706,N_49072,N_49560);
nor UO_4707 (O_4707,N_49537,N_49737);
nor UO_4708 (O_4708,N_49355,N_49422);
or UO_4709 (O_4709,N_49696,N_49326);
or UO_4710 (O_4710,N_49333,N_49223);
xor UO_4711 (O_4711,N_49832,N_49875);
nor UO_4712 (O_4712,N_49543,N_49818);
xnor UO_4713 (O_4713,N_49612,N_49273);
and UO_4714 (O_4714,N_49161,N_49796);
nor UO_4715 (O_4715,N_49020,N_49804);
or UO_4716 (O_4716,N_49029,N_49348);
and UO_4717 (O_4717,N_49785,N_49055);
nand UO_4718 (O_4718,N_49360,N_49910);
and UO_4719 (O_4719,N_49725,N_49217);
and UO_4720 (O_4720,N_49689,N_49459);
nor UO_4721 (O_4721,N_49755,N_49718);
nand UO_4722 (O_4722,N_49056,N_49384);
xnor UO_4723 (O_4723,N_49906,N_49644);
or UO_4724 (O_4724,N_49708,N_49717);
and UO_4725 (O_4725,N_49229,N_49157);
xnor UO_4726 (O_4726,N_49743,N_49460);
xnor UO_4727 (O_4727,N_49484,N_49514);
nor UO_4728 (O_4728,N_49506,N_49442);
nand UO_4729 (O_4729,N_49391,N_49910);
or UO_4730 (O_4730,N_49829,N_49246);
or UO_4731 (O_4731,N_49699,N_49766);
and UO_4732 (O_4732,N_49739,N_49356);
or UO_4733 (O_4733,N_49087,N_49929);
nor UO_4734 (O_4734,N_49535,N_49250);
xnor UO_4735 (O_4735,N_49457,N_49466);
or UO_4736 (O_4736,N_49027,N_49237);
nand UO_4737 (O_4737,N_49207,N_49791);
or UO_4738 (O_4738,N_49187,N_49314);
and UO_4739 (O_4739,N_49358,N_49683);
and UO_4740 (O_4740,N_49844,N_49890);
or UO_4741 (O_4741,N_49125,N_49777);
nor UO_4742 (O_4742,N_49977,N_49192);
xnor UO_4743 (O_4743,N_49970,N_49527);
nor UO_4744 (O_4744,N_49720,N_49940);
nor UO_4745 (O_4745,N_49254,N_49962);
or UO_4746 (O_4746,N_49835,N_49479);
and UO_4747 (O_4747,N_49260,N_49504);
and UO_4748 (O_4748,N_49031,N_49769);
nor UO_4749 (O_4749,N_49957,N_49623);
xnor UO_4750 (O_4750,N_49354,N_49582);
nand UO_4751 (O_4751,N_49554,N_49985);
nor UO_4752 (O_4752,N_49039,N_49946);
nand UO_4753 (O_4753,N_49483,N_49528);
and UO_4754 (O_4754,N_49603,N_49761);
xnor UO_4755 (O_4755,N_49693,N_49935);
or UO_4756 (O_4756,N_49590,N_49095);
xnor UO_4757 (O_4757,N_49065,N_49231);
or UO_4758 (O_4758,N_49519,N_49860);
nand UO_4759 (O_4759,N_49392,N_49830);
xnor UO_4760 (O_4760,N_49192,N_49577);
or UO_4761 (O_4761,N_49980,N_49364);
or UO_4762 (O_4762,N_49996,N_49456);
and UO_4763 (O_4763,N_49476,N_49411);
and UO_4764 (O_4764,N_49965,N_49054);
xor UO_4765 (O_4765,N_49991,N_49609);
xor UO_4766 (O_4766,N_49744,N_49193);
or UO_4767 (O_4767,N_49250,N_49695);
and UO_4768 (O_4768,N_49296,N_49596);
nand UO_4769 (O_4769,N_49019,N_49415);
xnor UO_4770 (O_4770,N_49882,N_49622);
or UO_4771 (O_4771,N_49854,N_49095);
xor UO_4772 (O_4772,N_49014,N_49391);
nand UO_4773 (O_4773,N_49652,N_49398);
and UO_4774 (O_4774,N_49186,N_49753);
and UO_4775 (O_4775,N_49788,N_49810);
and UO_4776 (O_4776,N_49142,N_49114);
nand UO_4777 (O_4777,N_49834,N_49962);
xor UO_4778 (O_4778,N_49102,N_49008);
nor UO_4779 (O_4779,N_49306,N_49657);
xnor UO_4780 (O_4780,N_49965,N_49301);
and UO_4781 (O_4781,N_49818,N_49092);
nor UO_4782 (O_4782,N_49137,N_49824);
nor UO_4783 (O_4783,N_49811,N_49980);
nor UO_4784 (O_4784,N_49828,N_49903);
xor UO_4785 (O_4785,N_49162,N_49506);
nand UO_4786 (O_4786,N_49683,N_49763);
nand UO_4787 (O_4787,N_49224,N_49435);
xor UO_4788 (O_4788,N_49614,N_49005);
nand UO_4789 (O_4789,N_49854,N_49109);
nand UO_4790 (O_4790,N_49102,N_49724);
xnor UO_4791 (O_4791,N_49030,N_49214);
or UO_4792 (O_4792,N_49395,N_49173);
xnor UO_4793 (O_4793,N_49458,N_49843);
nand UO_4794 (O_4794,N_49392,N_49139);
nand UO_4795 (O_4795,N_49686,N_49468);
and UO_4796 (O_4796,N_49382,N_49334);
or UO_4797 (O_4797,N_49201,N_49540);
xnor UO_4798 (O_4798,N_49278,N_49172);
xor UO_4799 (O_4799,N_49477,N_49820);
xor UO_4800 (O_4800,N_49956,N_49618);
nor UO_4801 (O_4801,N_49519,N_49480);
nand UO_4802 (O_4802,N_49528,N_49080);
and UO_4803 (O_4803,N_49448,N_49294);
xnor UO_4804 (O_4804,N_49140,N_49519);
xnor UO_4805 (O_4805,N_49633,N_49490);
nand UO_4806 (O_4806,N_49325,N_49997);
nor UO_4807 (O_4807,N_49345,N_49119);
and UO_4808 (O_4808,N_49129,N_49995);
or UO_4809 (O_4809,N_49923,N_49891);
and UO_4810 (O_4810,N_49470,N_49019);
and UO_4811 (O_4811,N_49518,N_49209);
nand UO_4812 (O_4812,N_49938,N_49397);
or UO_4813 (O_4813,N_49308,N_49704);
or UO_4814 (O_4814,N_49810,N_49547);
and UO_4815 (O_4815,N_49556,N_49253);
nand UO_4816 (O_4816,N_49619,N_49803);
nor UO_4817 (O_4817,N_49397,N_49555);
or UO_4818 (O_4818,N_49545,N_49660);
and UO_4819 (O_4819,N_49880,N_49304);
nand UO_4820 (O_4820,N_49746,N_49523);
nand UO_4821 (O_4821,N_49550,N_49031);
nor UO_4822 (O_4822,N_49422,N_49281);
or UO_4823 (O_4823,N_49688,N_49352);
xnor UO_4824 (O_4824,N_49590,N_49664);
xnor UO_4825 (O_4825,N_49953,N_49898);
nor UO_4826 (O_4826,N_49057,N_49530);
and UO_4827 (O_4827,N_49359,N_49582);
and UO_4828 (O_4828,N_49891,N_49636);
or UO_4829 (O_4829,N_49534,N_49067);
or UO_4830 (O_4830,N_49507,N_49052);
or UO_4831 (O_4831,N_49215,N_49860);
xnor UO_4832 (O_4832,N_49656,N_49456);
nor UO_4833 (O_4833,N_49642,N_49669);
and UO_4834 (O_4834,N_49652,N_49370);
nand UO_4835 (O_4835,N_49804,N_49950);
nand UO_4836 (O_4836,N_49742,N_49229);
xor UO_4837 (O_4837,N_49419,N_49109);
nand UO_4838 (O_4838,N_49460,N_49039);
and UO_4839 (O_4839,N_49987,N_49880);
nand UO_4840 (O_4840,N_49922,N_49442);
nand UO_4841 (O_4841,N_49471,N_49674);
xnor UO_4842 (O_4842,N_49502,N_49223);
or UO_4843 (O_4843,N_49892,N_49337);
nand UO_4844 (O_4844,N_49684,N_49058);
and UO_4845 (O_4845,N_49351,N_49108);
xnor UO_4846 (O_4846,N_49839,N_49740);
nor UO_4847 (O_4847,N_49548,N_49492);
and UO_4848 (O_4848,N_49632,N_49676);
or UO_4849 (O_4849,N_49920,N_49844);
or UO_4850 (O_4850,N_49769,N_49839);
nand UO_4851 (O_4851,N_49184,N_49589);
and UO_4852 (O_4852,N_49394,N_49597);
xor UO_4853 (O_4853,N_49255,N_49476);
xnor UO_4854 (O_4854,N_49454,N_49054);
xnor UO_4855 (O_4855,N_49698,N_49978);
xnor UO_4856 (O_4856,N_49853,N_49309);
or UO_4857 (O_4857,N_49195,N_49443);
or UO_4858 (O_4858,N_49400,N_49936);
nor UO_4859 (O_4859,N_49711,N_49857);
nand UO_4860 (O_4860,N_49868,N_49446);
xnor UO_4861 (O_4861,N_49991,N_49030);
xnor UO_4862 (O_4862,N_49637,N_49916);
nand UO_4863 (O_4863,N_49617,N_49056);
or UO_4864 (O_4864,N_49481,N_49862);
and UO_4865 (O_4865,N_49311,N_49221);
and UO_4866 (O_4866,N_49117,N_49251);
and UO_4867 (O_4867,N_49241,N_49326);
and UO_4868 (O_4868,N_49953,N_49397);
and UO_4869 (O_4869,N_49585,N_49989);
xnor UO_4870 (O_4870,N_49611,N_49835);
nand UO_4871 (O_4871,N_49195,N_49978);
xnor UO_4872 (O_4872,N_49616,N_49998);
xor UO_4873 (O_4873,N_49851,N_49396);
or UO_4874 (O_4874,N_49029,N_49619);
or UO_4875 (O_4875,N_49103,N_49237);
and UO_4876 (O_4876,N_49048,N_49218);
xor UO_4877 (O_4877,N_49596,N_49462);
xor UO_4878 (O_4878,N_49966,N_49515);
and UO_4879 (O_4879,N_49422,N_49941);
xor UO_4880 (O_4880,N_49102,N_49544);
or UO_4881 (O_4881,N_49234,N_49829);
and UO_4882 (O_4882,N_49806,N_49502);
nor UO_4883 (O_4883,N_49824,N_49979);
and UO_4884 (O_4884,N_49489,N_49038);
or UO_4885 (O_4885,N_49930,N_49995);
xnor UO_4886 (O_4886,N_49923,N_49596);
xnor UO_4887 (O_4887,N_49587,N_49066);
nand UO_4888 (O_4888,N_49666,N_49520);
nor UO_4889 (O_4889,N_49255,N_49713);
and UO_4890 (O_4890,N_49650,N_49283);
or UO_4891 (O_4891,N_49019,N_49187);
xnor UO_4892 (O_4892,N_49381,N_49220);
or UO_4893 (O_4893,N_49559,N_49662);
nand UO_4894 (O_4894,N_49907,N_49605);
xor UO_4895 (O_4895,N_49875,N_49189);
nand UO_4896 (O_4896,N_49743,N_49904);
nand UO_4897 (O_4897,N_49985,N_49057);
or UO_4898 (O_4898,N_49625,N_49321);
and UO_4899 (O_4899,N_49043,N_49894);
xor UO_4900 (O_4900,N_49953,N_49136);
xor UO_4901 (O_4901,N_49057,N_49291);
nor UO_4902 (O_4902,N_49530,N_49497);
and UO_4903 (O_4903,N_49772,N_49097);
nor UO_4904 (O_4904,N_49226,N_49526);
and UO_4905 (O_4905,N_49766,N_49305);
xnor UO_4906 (O_4906,N_49443,N_49489);
xnor UO_4907 (O_4907,N_49739,N_49015);
nor UO_4908 (O_4908,N_49307,N_49172);
nor UO_4909 (O_4909,N_49915,N_49672);
nand UO_4910 (O_4910,N_49084,N_49891);
and UO_4911 (O_4911,N_49785,N_49469);
xnor UO_4912 (O_4912,N_49835,N_49630);
xnor UO_4913 (O_4913,N_49594,N_49386);
nor UO_4914 (O_4914,N_49715,N_49910);
and UO_4915 (O_4915,N_49385,N_49598);
xor UO_4916 (O_4916,N_49080,N_49056);
nand UO_4917 (O_4917,N_49414,N_49681);
xnor UO_4918 (O_4918,N_49438,N_49322);
xor UO_4919 (O_4919,N_49351,N_49243);
and UO_4920 (O_4920,N_49625,N_49207);
xor UO_4921 (O_4921,N_49064,N_49276);
and UO_4922 (O_4922,N_49085,N_49800);
nor UO_4923 (O_4923,N_49084,N_49785);
nand UO_4924 (O_4924,N_49038,N_49363);
nand UO_4925 (O_4925,N_49410,N_49544);
nand UO_4926 (O_4926,N_49697,N_49405);
xor UO_4927 (O_4927,N_49369,N_49324);
or UO_4928 (O_4928,N_49239,N_49402);
nor UO_4929 (O_4929,N_49099,N_49778);
xor UO_4930 (O_4930,N_49945,N_49035);
nor UO_4931 (O_4931,N_49409,N_49771);
or UO_4932 (O_4932,N_49625,N_49225);
nor UO_4933 (O_4933,N_49375,N_49186);
nand UO_4934 (O_4934,N_49309,N_49582);
xor UO_4935 (O_4935,N_49252,N_49881);
or UO_4936 (O_4936,N_49901,N_49303);
nor UO_4937 (O_4937,N_49400,N_49972);
nor UO_4938 (O_4938,N_49562,N_49922);
nor UO_4939 (O_4939,N_49718,N_49078);
or UO_4940 (O_4940,N_49352,N_49743);
nor UO_4941 (O_4941,N_49546,N_49102);
and UO_4942 (O_4942,N_49168,N_49171);
xnor UO_4943 (O_4943,N_49801,N_49266);
nor UO_4944 (O_4944,N_49769,N_49304);
xnor UO_4945 (O_4945,N_49607,N_49822);
xnor UO_4946 (O_4946,N_49111,N_49591);
and UO_4947 (O_4947,N_49789,N_49187);
nand UO_4948 (O_4948,N_49582,N_49951);
xnor UO_4949 (O_4949,N_49815,N_49933);
nor UO_4950 (O_4950,N_49078,N_49519);
and UO_4951 (O_4951,N_49390,N_49200);
or UO_4952 (O_4952,N_49775,N_49174);
nor UO_4953 (O_4953,N_49004,N_49782);
and UO_4954 (O_4954,N_49129,N_49176);
xnor UO_4955 (O_4955,N_49304,N_49310);
xor UO_4956 (O_4956,N_49598,N_49458);
or UO_4957 (O_4957,N_49766,N_49011);
xnor UO_4958 (O_4958,N_49971,N_49407);
nor UO_4959 (O_4959,N_49670,N_49308);
xnor UO_4960 (O_4960,N_49900,N_49959);
and UO_4961 (O_4961,N_49813,N_49164);
nand UO_4962 (O_4962,N_49819,N_49428);
xnor UO_4963 (O_4963,N_49760,N_49157);
nor UO_4964 (O_4964,N_49555,N_49435);
or UO_4965 (O_4965,N_49930,N_49018);
nand UO_4966 (O_4966,N_49686,N_49370);
xor UO_4967 (O_4967,N_49902,N_49368);
xor UO_4968 (O_4968,N_49003,N_49206);
nor UO_4969 (O_4969,N_49900,N_49851);
and UO_4970 (O_4970,N_49606,N_49712);
or UO_4971 (O_4971,N_49020,N_49776);
nand UO_4972 (O_4972,N_49666,N_49768);
nand UO_4973 (O_4973,N_49427,N_49458);
nand UO_4974 (O_4974,N_49007,N_49637);
nand UO_4975 (O_4975,N_49069,N_49072);
or UO_4976 (O_4976,N_49976,N_49122);
or UO_4977 (O_4977,N_49285,N_49049);
and UO_4978 (O_4978,N_49866,N_49729);
xor UO_4979 (O_4979,N_49156,N_49366);
or UO_4980 (O_4980,N_49049,N_49689);
nand UO_4981 (O_4981,N_49072,N_49335);
nand UO_4982 (O_4982,N_49656,N_49882);
and UO_4983 (O_4983,N_49176,N_49505);
nor UO_4984 (O_4984,N_49926,N_49868);
or UO_4985 (O_4985,N_49564,N_49594);
xnor UO_4986 (O_4986,N_49649,N_49007);
xor UO_4987 (O_4987,N_49730,N_49676);
and UO_4988 (O_4988,N_49819,N_49615);
nor UO_4989 (O_4989,N_49083,N_49520);
nor UO_4990 (O_4990,N_49728,N_49950);
nor UO_4991 (O_4991,N_49475,N_49425);
nand UO_4992 (O_4992,N_49192,N_49312);
nor UO_4993 (O_4993,N_49247,N_49825);
and UO_4994 (O_4994,N_49574,N_49689);
and UO_4995 (O_4995,N_49008,N_49654);
or UO_4996 (O_4996,N_49742,N_49001);
nand UO_4997 (O_4997,N_49321,N_49038);
nand UO_4998 (O_4998,N_49906,N_49213);
and UO_4999 (O_4999,N_49567,N_49761);
endmodule