module basic_2000_20000_2500_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1379,In_1923);
nor U1 (N_1,In_392,In_578);
or U2 (N_2,In_594,In_1238);
nand U3 (N_3,In_583,In_845);
or U4 (N_4,In_1431,In_1943);
nand U5 (N_5,In_27,In_1003);
or U6 (N_6,In_1051,In_225);
or U7 (N_7,In_401,In_1066);
or U8 (N_8,In_1504,In_1600);
nand U9 (N_9,In_1150,In_308);
nand U10 (N_10,In_551,In_1561);
nand U11 (N_11,In_610,In_772);
nor U12 (N_12,In_321,In_1632);
and U13 (N_13,In_1472,In_75);
or U14 (N_14,In_524,In_967);
xnor U15 (N_15,In_329,In_188);
nand U16 (N_16,In_1221,In_474);
nand U17 (N_17,In_86,In_1851);
or U18 (N_18,In_160,In_1217);
and U19 (N_19,In_1081,In_1102);
nor U20 (N_20,In_52,In_1772);
nand U21 (N_21,In_1018,In_390);
or U22 (N_22,In_1073,In_1760);
and U23 (N_23,In_1307,In_30);
or U24 (N_24,In_1695,In_1161);
xor U25 (N_25,In_1998,In_489);
xnor U26 (N_26,In_1854,In_97);
and U27 (N_27,In_289,In_1512);
and U28 (N_28,In_1718,In_332);
or U29 (N_29,In_1913,In_196);
xnor U30 (N_30,In_1162,In_1730);
and U31 (N_31,In_912,In_1176);
nor U32 (N_32,In_1787,In_1380);
nor U33 (N_33,In_436,In_1319);
nor U34 (N_34,In_1287,In_1000);
and U35 (N_35,In_848,In_1711);
or U36 (N_36,In_90,In_71);
or U37 (N_37,In_876,In_643);
and U38 (N_38,In_1311,In_701);
nand U39 (N_39,In_1761,In_1643);
or U40 (N_40,In_1402,In_693);
or U41 (N_41,In_1118,In_17);
nor U42 (N_42,In_1139,In_1870);
nor U43 (N_43,In_1293,In_1327);
nand U44 (N_44,In_975,In_310);
nor U45 (N_45,In_1346,In_1853);
or U46 (N_46,In_928,In_1029);
nand U47 (N_47,In_341,In_124);
nor U48 (N_48,In_507,In_1861);
xor U49 (N_49,In_800,In_414);
xor U50 (N_50,In_1507,In_349);
xnor U51 (N_51,In_900,In_103);
nor U52 (N_52,In_295,In_1734);
or U53 (N_53,In_1912,In_477);
nor U54 (N_54,In_1664,In_1275);
or U55 (N_55,In_627,In_1849);
and U56 (N_56,In_860,In_1631);
nand U57 (N_57,In_304,In_847);
and U58 (N_58,In_810,In_1929);
xnor U59 (N_59,In_731,In_363);
or U60 (N_60,In_842,In_1628);
xor U61 (N_61,In_1814,In_81);
nand U62 (N_62,In_151,In_1147);
and U63 (N_63,In_797,In_495);
xor U64 (N_64,In_1426,In_1336);
nor U65 (N_65,In_1850,In_1758);
xnor U66 (N_66,In_1676,In_1501);
nor U67 (N_67,In_290,In_770);
xor U68 (N_68,In_286,In_443);
nor U69 (N_69,In_1422,In_1973);
and U70 (N_70,In_77,In_1776);
or U71 (N_71,In_1441,In_650);
or U72 (N_72,In_587,In_107);
nand U73 (N_73,In_128,In_1617);
and U74 (N_74,In_665,In_1585);
xnor U75 (N_75,In_155,In_1403);
or U76 (N_76,In_1612,In_1484);
nor U77 (N_77,In_1188,In_316);
xnor U78 (N_78,In_98,In_624);
nand U79 (N_79,In_490,In_1658);
nand U80 (N_80,In_827,In_790);
xnor U81 (N_81,In_1198,In_742);
nand U82 (N_82,In_1526,In_1947);
nand U83 (N_83,In_512,In_1322);
or U84 (N_84,In_408,In_994);
nor U85 (N_85,In_194,In_210);
and U86 (N_86,In_1439,In_419);
xor U87 (N_87,In_33,In_461);
or U88 (N_88,In_616,In_13);
xnor U89 (N_89,In_139,In_1265);
nor U90 (N_90,In_230,In_1562);
and U91 (N_91,In_1595,In_428);
or U92 (N_92,In_1412,In_1341);
and U93 (N_93,In_240,In_1009);
or U94 (N_94,In_1707,In_792);
xor U95 (N_95,In_1520,In_862);
nor U96 (N_96,In_169,In_1078);
xor U97 (N_97,In_1185,In_325);
xnor U98 (N_98,In_360,In_1087);
nor U99 (N_99,In_161,In_266);
and U100 (N_100,In_434,In_1358);
or U101 (N_101,In_1822,In_1661);
nand U102 (N_102,In_924,In_1563);
nand U103 (N_103,In_1685,In_809);
and U104 (N_104,In_1729,In_949);
nor U105 (N_105,In_1032,In_406);
and U106 (N_106,In_1012,In_1510);
and U107 (N_107,In_1249,In_785);
or U108 (N_108,In_1765,In_1682);
nand U109 (N_109,In_754,In_121);
nand U110 (N_110,In_700,In_1572);
xor U111 (N_111,In_1714,In_181);
and U112 (N_112,In_41,In_1424);
and U113 (N_113,In_233,In_762);
xor U114 (N_114,In_1283,In_226);
nand U115 (N_115,In_599,In_714);
and U116 (N_116,In_555,In_1590);
or U117 (N_117,In_1039,In_966);
or U118 (N_118,In_447,In_1928);
and U119 (N_119,In_1976,In_1392);
nand U120 (N_120,In_1946,In_1114);
nand U121 (N_121,In_560,In_856);
nand U122 (N_122,In_898,In_576);
xnor U123 (N_123,In_1037,In_1187);
xnor U124 (N_124,In_1253,In_386);
or U125 (N_125,In_683,In_1212);
xnor U126 (N_126,In_1807,In_276);
nor U127 (N_127,In_1706,In_268);
or U128 (N_128,In_1309,In_1663);
or U129 (N_129,In_1724,In_1206);
and U130 (N_130,In_1789,In_905);
nand U131 (N_131,In_844,In_697);
nor U132 (N_132,In_1337,In_1317);
nor U133 (N_133,In_351,In_1015);
xor U134 (N_134,In_147,In_106);
xnor U135 (N_135,In_821,In_305);
or U136 (N_136,In_1074,In_618);
or U137 (N_137,In_1404,In_1677);
nor U138 (N_138,In_1038,In_93);
and U139 (N_139,In_620,In_273);
or U140 (N_140,In_1517,In_942);
nand U141 (N_141,In_116,In_277);
and U142 (N_142,In_1136,In_1497);
or U143 (N_143,In_167,In_1108);
nand U144 (N_144,In_1483,In_202);
xor U145 (N_145,In_1732,In_192);
xor U146 (N_146,In_958,In_1480);
nand U147 (N_147,In_868,In_562);
xor U148 (N_148,In_1615,In_1021);
or U149 (N_149,In_1812,In_1644);
nand U150 (N_150,In_750,In_1027);
xor U151 (N_151,In_982,In_874);
xnor U152 (N_152,In_945,In_1826);
nor U153 (N_153,In_1276,In_365);
and U154 (N_154,In_1836,In_866);
or U155 (N_155,In_1802,In_66);
nor U156 (N_156,In_981,In_342);
and U157 (N_157,In_1626,In_1171);
nor U158 (N_158,In_1531,In_270);
and U159 (N_159,In_424,In_1816);
or U160 (N_160,In_872,In_374);
xnor U161 (N_161,In_398,In_539);
nand U162 (N_162,In_1268,In_659);
or U163 (N_163,In_119,In_1377);
or U164 (N_164,In_483,In_435);
and U165 (N_165,In_1475,In_1057);
and U166 (N_166,In_972,In_1214);
and U167 (N_167,In_193,In_645);
nor U168 (N_168,In_499,In_1951);
and U169 (N_169,In_1020,In_10);
and U170 (N_170,In_777,In_1623);
nand U171 (N_171,In_550,In_937);
or U172 (N_172,In_1,In_669);
and U173 (N_173,In_300,In_1264);
nand U174 (N_174,In_29,In_122);
nand U175 (N_175,In_1479,In_1825);
nor U176 (N_176,In_1324,In_999);
and U177 (N_177,In_470,In_707);
and U178 (N_178,In_1454,In_350);
and U179 (N_179,In_317,In_1558);
or U180 (N_180,In_1827,In_246);
nor U181 (N_181,In_702,In_32);
and U182 (N_182,In_664,In_1602);
xor U183 (N_183,In_1005,In_244);
nor U184 (N_184,In_1984,In_1399);
nor U185 (N_185,In_1613,In_1725);
nand U186 (N_186,In_1914,In_138);
xor U187 (N_187,In_1616,In_698);
or U188 (N_188,In_783,In_852);
and U189 (N_189,In_1149,In_1524);
nand U190 (N_190,In_1806,In_239);
nand U191 (N_191,In_347,In_55);
nor U192 (N_192,In_1058,In_1965);
nand U193 (N_193,In_454,In_563);
xor U194 (N_194,In_82,In_796);
nand U195 (N_195,In_123,In_1476);
nand U196 (N_196,In_168,In_186);
xnor U197 (N_197,In_1292,In_1222);
or U198 (N_198,In_726,In_48);
nand U199 (N_199,In_1937,In_156);
and U200 (N_200,In_1838,In_1941);
and U201 (N_201,In_484,In_1077);
nand U202 (N_202,In_1314,In_888);
xor U203 (N_203,In_915,In_387);
or U204 (N_204,In_590,In_1873);
nor U205 (N_205,In_553,In_430);
xor U206 (N_206,In_1556,In_765);
nand U207 (N_207,In_815,In_1641);
nand U208 (N_208,In_1678,In_871);
nand U209 (N_209,In_1331,In_298);
or U210 (N_210,In_913,In_1462);
nand U211 (N_211,In_120,In_1306);
and U212 (N_212,In_1902,In_1587);
nand U213 (N_213,In_200,In_884);
and U214 (N_214,In_1508,In_1353);
and U215 (N_215,In_1071,In_385);
nor U216 (N_216,In_965,In_154);
nand U217 (N_217,In_1376,In_1178);
nand U218 (N_218,In_1609,In_1796);
or U219 (N_219,In_1938,In_1375);
nor U220 (N_220,In_545,In_838);
xnor U221 (N_221,In_222,In_1408);
xnor U222 (N_222,In_1614,In_1843);
or U223 (N_223,In_1239,In_37);
or U224 (N_224,In_279,In_996);
nor U225 (N_225,In_1667,In_1112);
nand U226 (N_226,In_330,In_536);
nor U227 (N_227,In_117,In_541);
or U228 (N_228,In_1304,In_251);
nand U229 (N_229,In_1095,In_1487);
xor U230 (N_230,In_1285,In_1592);
and U231 (N_231,In_1895,In_780);
or U232 (N_232,In_1415,In_1271);
nand U233 (N_233,In_699,In_1876);
nor U234 (N_234,In_1633,In_1908);
nor U235 (N_235,In_493,In_991);
xnor U236 (N_236,In_1719,In_1611);
xor U237 (N_237,In_198,In_1605);
nor U238 (N_238,In_1897,In_203);
xor U239 (N_239,In_899,In_311);
and U240 (N_240,In_1430,In_1061);
or U241 (N_241,In_944,In_668);
nand U242 (N_242,In_1330,In_486);
xor U243 (N_243,In_1260,In_1781);
nor U244 (N_244,In_1799,In_1269);
nand U245 (N_245,In_1753,In_444);
xnor U246 (N_246,In_1298,In_1192);
nand U247 (N_247,In_1429,In_508);
or U248 (N_248,In_1859,In_1553);
or U249 (N_249,In_1817,In_1010);
nor U250 (N_250,In_849,In_1294);
or U251 (N_251,In_811,In_150);
nand U252 (N_252,In_1247,In_736);
or U253 (N_253,In_453,In_1208);
nor U254 (N_254,In_172,In_1181);
xnor U255 (N_255,In_509,In_729);
nand U256 (N_256,In_165,In_1344);
xor U257 (N_257,In_1210,In_109);
or U258 (N_258,In_1554,In_397);
nand U259 (N_259,In_175,In_463);
nand U260 (N_260,In_719,In_1156);
nand U261 (N_261,In_1014,In_974);
xnor U262 (N_262,In_189,In_565);
and U263 (N_263,In_1154,In_1205);
nand U264 (N_264,In_1026,In_812);
nand U265 (N_265,In_696,In_1991);
xnor U266 (N_266,In_923,In_1601);
nor U267 (N_267,In_1608,In_920);
xnor U268 (N_268,In_1352,In_1803);
xor U269 (N_269,In_721,In_326);
nand U270 (N_270,In_813,In_1070);
nor U271 (N_271,In_208,In_191);
or U272 (N_272,In_1362,In_1235);
xnor U273 (N_273,In_376,In_1278);
nand U274 (N_274,In_88,In_802);
nor U275 (N_275,In_1373,In_104);
and U276 (N_276,In_243,In_609);
and U277 (N_277,In_1668,In_980);
nor U278 (N_278,In_1444,In_1215);
and U279 (N_279,In_893,In_788);
xor U280 (N_280,In_47,In_1700);
nand U281 (N_281,In_1610,In_955);
nand U282 (N_282,In_672,In_904);
or U283 (N_283,In_80,In_1939);
nor U284 (N_284,In_1469,In_262);
nor U285 (N_285,In_652,In_85);
nand U286 (N_286,In_759,In_25);
xor U287 (N_287,In_766,In_585);
or U288 (N_288,In_677,In_673);
nor U289 (N_289,In_1801,In_348);
or U290 (N_290,In_1140,In_218);
nor U291 (N_291,In_1420,In_1202);
xnor U292 (N_292,In_223,In_1457);
nand U293 (N_293,In_241,In_598);
xnor U294 (N_294,In_205,In_603);
nand U295 (N_295,In_1548,In_1721);
nand U296 (N_296,In_1654,In_1717);
and U297 (N_297,In_53,In_640);
or U298 (N_298,In_1871,In_658);
nor U299 (N_299,In_666,In_1693);
nand U300 (N_300,In_684,In_1131);
xor U301 (N_301,In_1440,In_1323);
or U302 (N_302,In_1433,In_144);
or U303 (N_303,In_703,In_378);
nand U304 (N_304,In_1523,In_1972);
or U305 (N_305,In_1999,In_481);
and U306 (N_306,In_1153,In_70);
or U307 (N_307,In_889,In_38);
or U308 (N_308,In_1751,In_778);
xnor U309 (N_309,In_709,In_1931);
nor U310 (N_310,In_1922,In_1930);
or U311 (N_311,In_1257,In_817);
xnor U312 (N_312,In_569,In_1279);
nor U313 (N_313,In_581,In_1863);
and U314 (N_314,In_543,In_83);
xnor U315 (N_315,In_1907,In_695);
nand U316 (N_316,In_739,In_857);
and U317 (N_317,In_769,In_34);
and U318 (N_318,In_1582,In_1833);
and U319 (N_319,In_1478,In_79);
and U320 (N_320,In_1123,In_1115);
xor U321 (N_321,In_275,In_1398);
xnor U322 (N_322,In_67,In_1233);
nor U323 (N_323,In_1715,In_1088);
nand U324 (N_324,In_1918,In_1967);
or U325 (N_325,In_779,In_918);
and U326 (N_326,In_929,In_1974);
nand U327 (N_327,In_1637,In_630);
or U328 (N_328,In_1190,In_671);
or U329 (N_329,In_548,In_1446);
and U330 (N_330,In_1213,In_328);
nor U331 (N_331,In_1167,In_356);
or U332 (N_332,In_1409,In_1227);
and U333 (N_333,In_1735,In_213);
nor U334 (N_334,In_1818,In_511);
xnor U335 (N_335,In_1391,In_588);
and U336 (N_336,In_1418,In_1840);
and U337 (N_337,In_1726,In_1129);
nand U338 (N_338,In_320,In_1086);
nand U339 (N_339,In_331,In_897);
or U340 (N_340,In_61,In_1072);
or U341 (N_341,In_694,In_663);
nor U342 (N_342,In_220,In_657);
nand U343 (N_343,In_256,In_201);
and U344 (N_344,In_1727,In_1366);
nor U345 (N_345,In_1211,In_629);
xor U346 (N_346,In_7,In_1017);
nand U347 (N_347,In_1450,In_16);
nor U348 (N_348,In_1107,In_396);
or U349 (N_349,In_1228,In_76);
and U350 (N_350,In_1485,In_1442);
xnor U351 (N_351,In_322,In_1891);
or U352 (N_352,In_132,In_1704);
xor U353 (N_353,In_1852,In_1993);
nor U354 (N_354,In_628,In_1569);
nand U355 (N_355,In_1223,In_110);
nand U356 (N_356,In_1195,In_114);
nand U357 (N_357,In_494,In_1094);
xnor U358 (N_358,In_1680,In_840);
nand U359 (N_359,In_1622,In_1575);
nor U360 (N_360,In_992,In_960);
or U361 (N_361,In_1350,In_1688);
nor U362 (N_362,In_971,In_854);
or U363 (N_363,In_1522,In_1675);
or U364 (N_364,In_1845,In_1924);
and U365 (N_365,In_1552,In_1369);
or U366 (N_366,In_505,In_1437);
or U367 (N_367,In_724,In_727);
and U368 (N_368,In_1097,In_6);
nor U369 (N_369,In_87,In_559);
xor U370 (N_370,In_1542,In_1494);
xor U371 (N_371,In_916,In_1339);
or U372 (N_372,In_823,In_1477);
or U373 (N_373,In_1964,In_1525);
nor U374 (N_374,In_1085,In_102);
or U375 (N_375,In_140,In_1823);
nand U376 (N_376,In_936,In_1745);
xnor U377 (N_377,In_1425,In_834);
nor U378 (N_378,In_1829,In_1981);
nand U379 (N_379,In_312,In_1056);
and U380 (N_380,In_850,In_1839);
and U381 (N_381,In_1988,In_1573);
nand U382 (N_382,In_451,In_43);
xnor U383 (N_383,In_460,In_1906);
and U384 (N_384,In_1465,In_748);
nand U385 (N_385,In_1579,In_1694);
nor U386 (N_386,In_299,In_1541);
nand U387 (N_387,In_1888,In_125);
xor U388 (N_388,In_1428,In_1042);
nand U389 (N_389,In_1992,In_688);
nand U390 (N_390,In_1461,In_283);
or U391 (N_391,In_1259,In_1499);
nor U392 (N_392,In_814,In_23);
nor U393 (N_393,In_626,In_1496);
nand U394 (N_394,In_527,In_957);
and U395 (N_395,In_1019,In_987);
nand U396 (N_396,In_1646,In_735);
nor U397 (N_397,In_492,In_1098);
nor U398 (N_398,In_1246,In_743);
and U399 (N_399,In_925,In_1400);
xor U400 (N_400,In_1200,In_1917);
xor U401 (N_401,In_864,In_1084);
nor U402 (N_402,In_1968,In_1957);
xor U403 (N_403,In_285,In_366);
or U404 (N_404,In_549,In_1657);
xnor U405 (N_405,In_831,In_951);
or U406 (N_406,In_1248,In_1093);
xor U407 (N_407,In_1242,In_795);
nor U408 (N_408,In_501,In_523);
nor U409 (N_409,In_1756,In_28);
and U410 (N_410,In_1893,In_361);
and U411 (N_411,In_1024,In_896);
nor U412 (N_412,In_642,In_45);
nand U413 (N_413,In_336,In_1388);
nor U414 (N_414,In_1049,In_1495);
and U415 (N_415,In_1881,In_728);
or U416 (N_416,In_1830,In_863);
xnor U417 (N_417,In_962,In_605);
or U418 (N_418,In_1696,In_1125);
nand U419 (N_419,In_1180,In_441);
xor U420 (N_420,In_614,In_934);
or U421 (N_421,In_529,In_1759);
or U422 (N_422,In_782,In_660);
and U423 (N_423,In_717,In_1831);
nor U424 (N_424,In_1218,In_1263);
nor U425 (N_425,In_1673,In_1251);
nor U426 (N_426,In_180,In_1326);
xor U427 (N_427,In_1464,In_1280);
nor U428 (N_428,In_1349,In_961);
and U429 (N_429,In_1564,In_415);
xnor U430 (N_430,In_1557,In_1396);
and U431 (N_431,In_1133,In_1703);
nor U432 (N_432,In_1148,In_1945);
and U433 (N_433,In_877,In_1354);
nor U434 (N_434,In_464,In_1518);
and U435 (N_435,In_1173,In_1624);
or U436 (N_436,In_1090,In_1410);
or U437 (N_437,In_458,In_1004);
xnor U438 (N_438,In_1124,In_740);
nand U439 (N_439,In_163,In_323);
nor U440 (N_440,In_177,In_998);
nand U441 (N_441,In_1193,In_1141);
xor U442 (N_442,In_14,In_467);
xor U443 (N_443,In_1513,In_1539);
and U444 (N_444,In_540,In_989);
or U445 (N_445,In_1597,In_1889);
xor U446 (N_446,In_1785,In_1357);
or U447 (N_447,In_655,In_259);
nand U448 (N_448,In_1954,In_1545);
or U449 (N_449,In_1069,In_1750);
nand U450 (N_450,In_1030,In_1808);
nand U451 (N_451,In_1295,In_1079);
and U452 (N_452,In_439,In_1417);
xor U453 (N_453,In_1768,In_1064);
and U454 (N_454,In_1698,In_1325);
nor U455 (N_455,In_1137,In_1255);
xor U456 (N_456,In_973,In_153);
nand U457 (N_457,In_9,In_12);
and U458 (N_458,In_602,In_1463);
xor U459 (N_459,In_1033,In_1791);
nor U460 (N_460,In_339,In_1747);
and U461 (N_461,In_1713,In_1184);
or U462 (N_462,In_713,In_1560);
or U463 (N_463,In_1231,In_1671);
nor U464 (N_464,In_1219,In_568);
and U465 (N_465,In_1013,In_1697);
or U466 (N_466,In_1532,In_134);
and U467 (N_467,In_1674,In_446);
xnor U468 (N_468,In_1708,In_438);
xor U469 (N_469,In_113,In_1647);
and U470 (N_470,In_522,In_836);
or U471 (N_471,In_654,In_195);
or U472 (N_472,In_1313,In_1782);
or U473 (N_473,In_338,In_1355);
nand U474 (N_474,In_786,In_1862);
nor U475 (N_475,In_636,In_263);
nand U476 (N_476,In_1864,In_1958);
and U477 (N_477,In_1456,In_1048);
nand U478 (N_478,In_725,In_1363);
nand U479 (N_479,In_1393,In_1683);
xor U480 (N_480,In_1896,In_418);
nor U481 (N_481,In_364,In_1530);
and U482 (N_482,In_274,In_1145);
and U483 (N_483,In_1467,In_681);
or U484 (N_484,In_1963,In_1712);
and U485 (N_485,In_411,In_370);
or U486 (N_486,In_1925,In_1686);
and U487 (N_487,In_557,In_1529);
or U488 (N_488,In_1565,In_1284);
nand U489 (N_489,In_1634,In_517);
nor U490 (N_490,In_1949,In_1333);
nand U491 (N_491,In_1691,In_15);
nor U492 (N_492,In_1296,In_440);
and U493 (N_493,In_1911,In_741);
nor U494 (N_494,In_142,In_1509);
xnor U495 (N_495,In_288,In_1250);
nand U496 (N_496,In_1288,In_1043);
and U497 (N_497,In_5,In_1394);
or U498 (N_498,In_885,In_1122);
or U499 (N_499,In_1533,In_1502);
and U500 (N_500,In_1687,In_395);
nor U501 (N_501,In_1890,In_373);
xnor U502 (N_502,In_948,In_216);
xnor U503 (N_503,In_352,In_18);
or U504 (N_504,In_1977,In_1128);
xor U505 (N_505,In_20,In_1411);
nand U506 (N_506,In_1550,In_1075);
and U507 (N_507,In_1733,In_1774);
and U508 (N_508,In_711,In_1743);
nor U509 (N_509,In_1920,In_841);
and U510 (N_510,In_1356,In_404);
and U511 (N_511,In_917,In_1471);
and U512 (N_512,In_405,In_215);
and U513 (N_513,In_1535,In_1544);
nor U514 (N_514,In_1299,In_1577);
xnor U515 (N_515,In_462,In_1291);
nand U516 (N_516,In_1621,In_1942);
nor U517 (N_517,In_789,In_1655);
and U518 (N_518,In_1316,In_737);
xor U519 (N_519,In_1382,In_1979);
and U520 (N_520,In_799,In_612);
or U521 (N_521,In_1910,In_344);
nor U522 (N_522,In_1104,In_1220);
and U523 (N_523,In_580,In_1121);
nand U524 (N_524,In_1879,In_280);
nand U525 (N_525,In_1679,In_1230);
and U526 (N_526,In_1819,In_248);
nand U527 (N_527,In_426,In_1488);
or U528 (N_528,In_1025,In_1254);
xor U529 (N_529,In_145,In_738);
xnor U530 (N_530,In_1491,In_1948);
xnor U531 (N_531,In_591,In_372);
nor U532 (N_532,In_648,In_384);
or U533 (N_533,In_260,In_829);
nor U534 (N_534,In_1361,In_1741);
nor U535 (N_535,In_1865,In_1877);
nand U536 (N_536,In_324,In_959);
nor U537 (N_537,In_531,In_1194);
nor U538 (N_538,In_1842,In_678);
and U539 (N_539,In_675,In_136);
nor U540 (N_540,In_257,In_1728);
nor U541 (N_541,In_985,In_940);
xnor U542 (N_542,In_1978,In_1652);
nor U543 (N_543,In_471,In_689);
nand U544 (N_544,In_1868,In_837);
xor U545 (N_545,In_89,In_1581);
and U546 (N_546,In_1427,In_1944);
nand U547 (N_547,In_1568,In_534);
xnor U548 (N_548,In_57,In_1875);
nor U549 (N_549,In_1639,In_1932);
nor U550 (N_550,In_1470,In_391);
and U551 (N_551,In_319,In_865);
and U552 (N_552,In_1297,In_1482);
nand U553 (N_553,In_1594,In_1528);
and U554 (N_554,In_519,In_1878);
or U555 (N_555,In_1882,In_853);
and U556 (N_556,In_927,In_127);
and U557 (N_557,In_633,In_410);
xnor U558 (N_558,In_264,In_1068);
nor U559 (N_559,In_833,In_625);
and U560 (N_560,In_152,In_1282);
xnor U561 (N_561,In_421,In_46);
nand U562 (N_562,In_1289,In_561);
nor U563 (N_563,In_1340,In_1742);
and U564 (N_564,In_977,In_808);
nor U565 (N_565,In_212,In_1809);
nor U566 (N_566,In_1351,In_1549);
xor U567 (N_567,In_296,In_126);
nor U568 (N_568,In_1383,In_108);
nor U569 (N_569,In_733,In_1082);
and U570 (N_570,In_1236,In_807);
and U571 (N_571,In_1448,In_1046);
xnor U572 (N_572,In_556,In_498);
nor U573 (N_573,In_1045,In_422);
xnor U574 (N_574,In_1312,In_1489);
xnor U575 (N_575,In_747,In_528);
xnor U576 (N_576,In_1604,In_1002);
nand U577 (N_577,In_281,In_1837);
or U578 (N_578,In_761,In_1723);
nor U579 (N_579,In_1901,In_1884);
xnor U580 (N_580,In_635,In_1303);
xnor U581 (N_581,In_1933,In_1245);
nor U582 (N_582,In_1434,In_1599);
nor U583 (N_583,In_1731,In_516);
and U584 (N_584,In_1387,In_986);
and U585 (N_585,In_383,In_963);
or U586 (N_586,In_798,In_525);
or U587 (N_587,In_1055,In_318);
or U588 (N_588,In_595,In_869);
xor U589 (N_589,In_258,In_1053);
nor U590 (N_590,In_1047,In_639);
nand U591 (N_591,In_375,In_513);
nand U592 (N_592,In_1405,In_1035);
nor U593 (N_593,In_1113,In_661);
xor U594 (N_594,In_1335,In_825);
or U595 (N_595,In_1065,In_1659);
nor U596 (N_596,In_1754,In_1905);
and U597 (N_597,In_26,In_1770);
nor U598 (N_598,In_1261,In_306);
and U599 (N_599,In_503,In_1744);
nand U600 (N_600,In_1537,In_1815);
nand U601 (N_601,In_219,In_979);
nor U602 (N_602,In_1040,In_1769);
nand U603 (N_603,In_1169,In_1321);
or U604 (N_604,In_1407,In_990);
and U605 (N_605,In_333,In_1790);
xnor U606 (N_606,In_72,In_1580);
nand U607 (N_607,In_452,In_692);
and U608 (N_608,In_1701,In_1916);
nor U609 (N_609,In_1567,In_101);
xor U610 (N_610,In_1665,In_84);
and U611 (N_611,In_892,In_939);
nor U612 (N_612,In_1459,In_941);
and U613 (N_613,In_880,In_1710);
nor U614 (N_614,In_1159,In_1486);
xor U615 (N_615,In_932,In_1736);
or U616 (N_616,In_362,In_623);
or U617 (N_617,In_488,In_343);
and U618 (N_618,In_1500,In_1174);
and U619 (N_619,In_267,In_1225);
nand U620 (N_620,In_1551,In_1503);
nand U621 (N_621,In_1971,In_1083);
nor U622 (N_622,In_1950,In_781);
and U623 (N_623,In_1143,In_674);
and U624 (N_624,In_1996,In_1034);
xor U625 (N_625,In_207,In_632);
nor U626 (N_626,In_1648,In_969);
or U627 (N_627,In_170,In_749);
xnor U628 (N_628,In_11,In_575);
xnor U629 (N_629,In_157,In_1468);
or U630 (N_630,In_644,In_1546);
and U631 (N_631,In_997,In_173);
xnor U632 (N_632,In_459,In_716);
nor U633 (N_633,In_1226,In_1574);
nor U634 (N_634,In_956,In_943);
and U635 (N_635,In_1460,In_935);
xnor U636 (N_636,In_1709,In_1385);
and U637 (N_637,In_1099,In_855);
and U638 (N_638,In_255,In_954);
xnor U639 (N_639,In_582,In_64);
or U640 (N_640,In_882,In_953);
or U641 (N_641,In_1956,In_171);
xor U642 (N_642,In_1940,In_231);
xnor U643 (N_643,In_1305,In_1767);
xor U644 (N_644,In_1894,In_1584);
or U645 (N_645,In_606,In_137);
or U646 (N_646,In_574,In_647);
nand U647 (N_647,In_1752,In_1669);
xnor U648 (N_648,In_1466,In_1120);
nand U649 (N_649,In_1256,In_984);
and U650 (N_650,In_357,In_978);
xnor U651 (N_651,In_1273,In_1771);
xnor U652 (N_652,In_400,In_1059);
or U653 (N_653,In_402,In_78);
nand U654 (N_654,In_1959,In_773);
and U655 (N_655,In_1052,In_1089);
or U656 (N_656,In_1880,In_1347);
nor U657 (N_657,In_1915,In_879);
and U658 (N_658,In_73,In_820);
nand U659 (N_659,In_787,In_1438);
and U660 (N_660,In_537,In_1234);
nand U661 (N_661,In_634,In_302);
or U662 (N_662,In_804,In_1142);
xor U663 (N_663,In_1378,In_615);
and U664 (N_664,In_345,In_1490);
or U665 (N_665,In_1847,In_756);
xnor U666 (N_666,In_775,In_1886);
nand U667 (N_667,In_403,In_229);
nand U668 (N_668,In_1559,In_313);
or U669 (N_669,In_682,In_571);
xor U670 (N_670,In_1821,In_1684);
or U671 (N_671,In_526,In_19);
and U672 (N_672,In_250,In_554);
nor U673 (N_673,In_1797,In_1386);
nor U674 (N_674,In_111,In_174);
nand U675 (N_675,In_1435,In_619);
xnor U676 (N_676,In_1534,In_63);
xor U677 (N_677,In_1343,In_1705);
xor U678 (N_678,In_496,In_468);
nand U679 (N_679,In_952,In_1738);
nor U680 (N_680,In_950,In_221);
and U681 (N_681,In_760,In_679);
nor U682 (N_682,In_1885,In_1370);
and U683 (N_683,In_1764,In_1994);
nor U684 (N_684,In_1995,In_91);
nor U685 (N_685,In_1207,In_710);
xnor U686 (N_686,In_287,In_1635);
nor U687 (N_687,In_242,In_1091);
nand U688 (N_688,In_141,In_1636);
nor U689 (N_689,In_1315,In_1989);
nand U690 (N_690,In_819,In_1638);
xnor U691 (N_691,In_607,In_1739);
nand U692 (N_692,In_1903,In_469);
xnor U693 (N_693,In_449,In_1160);
or U694 (N_694,In_922,In_1151);
xor U695 (N_695,In_294,In_1997);
and U696 (N_696,In_1054,In_1779);
nor U697 (N_697,In_1062,In_1164);
and U698 (N_698,In_1505,In_1578);
nor U699 (N_699,In_429,In_1170);
or U700 (N_700,In_500,In_757);
xor U701 (N_701,In_455,In_497);
xor U702 (N_702,In_518,In_1955);
nand U703 (N_703,In_676,In_1252);
nand U704 (N_704,In_40,In_340);
and U705 (N_705,In_1824,In_292);
nand U706 (N_706,In_1146,In_1372);
and U707 (N_707,In_1919,In_297);
xnor U708 (N_708,In_204,In_1720);
xnor U709 (N_709,In_1445,In_1041);
nor U710 (N_710,In_1328,In_1898);
xnor U711 (N_711,In_1866,In_1755);
nor U712 (N_712,In_768,In_1650);
xor U713 (N_713,In_1540,In_1975);
nand U714 (N_714,In_1571,In_1591);
nand U715 (N_715,In_1926,In_1762);
nand U716 (N_716,In_826,In_1310);
nor U717 (N_717,In_1447,In_478);
nor U718 (N_718,In_976,In_970);
xor U719 (N_719,In_1547,In_1381);
nor U720 (N_720,In_1130,In_846);
nor U721 (N_721,In_793,In_722);
nand U722 (N_722,In_1241,In_1342);
xor U723 (N_723,In_926,In_1811);
xor U724 (N_724,In_431,In_1199);
and U725 (N_725,In_50,In_909);
or U726 (N_726,In_197,In_1419);
nand U727 (N_727,In_662,In_261);
nor U728 (N_728,In_1196,In_919);
nand U729 (N_729,In_309,In_708);
and U730 (N_730,In_35,In_354);
xnor U731 (N_731,In_1302,In_510);
or U732 (N_732,In_1474,In_1166);
xor U733 (N_733,In_506,In_1001);
nand U734 (N_734,In_1793,In_1023);
and U735 (N_735,In_1784,In_1191);
and U736 (N_736,In_670,In_1649);
nor U737 (N_737,In_254,In_1105);
xnor U738 (N_738,In_303,In_427);
xnor U739 (N_739,In_1277,In_1936);
nor U740 (N_740,In_1555,In_146);
nor U741 (N_741,In_907,In_611);
nor U742 (N_742,In_1927,In_69);
xor U743 (N_743,In_886,In_1716);
nand U744 (N_744,In_1301,In_214);
nand U745 (N_745,In_767,In_227);
nand U746 (N_746,In_485,In_1566);
nor U747 (N_747,In_1209,In_867);
nand U748 (N_748,In_1692,In_1101);
xor U749 (N_749,In_335,In_24);
or U750 (N_750,In_100,In_931);
nand U751 (N_751,In_1670,In_1748);
nor U752 (N_752,In_65,In_1498);
nor U753 (N_753,In_1583,In_1892);
xnor U754 (N_754,In_1134,In_74);
and U755 (N_755,In_49,In_1022);
xor U756 (N_756,In_521,In_1186);
nor U757 (N_757,In_1966,In_1813);
nand U758 (N_758,In_1157,In_236);
or U759 (N_759,In_1274,In_407);
nand U760 (N_760,In_1835,In_1778);
xor U761 (N_761,In_130,In_448);
nor U762 (N_762,In_465,In_622);
and U763 (N_763,In_1028,In_1792);
and U764 (N_764,In_1063,In_830);
nand U765 (N_765,In_558,In_228);
xnor U766 (N_766,In_613,In_1365);
and U767 (N_767,In_1395,In_1834);
or U768 (N_768,In_491,In_353);
or U769 (N_769,In_269,In_199);
and U770 (N_770,In_389,In_475);
and U771 (N_771,In_54,In_22);
nor U772 (N_772,In_1521,In_377);
nand U773 (N_773,In_445,In_995);
and U774 (N_774,In_564,In_1934);
nand U775 (N_775,In_479,In_51);
and U776 (N_776,In_394,In_1627);
nor U777 (N_777,In_593,In_58);
or U778 (N_778,In_1406,In_149);
and U779 (N_779,In_252,In_1783);
nor U780 (N_780,In_1067,In_938);
or U781 (N_781,In_178,In_1961);
or U782 (N_782,In_1458,In_1921);
and U783 (N_783,In_1506,In_903);
nor U784 (N_784,In_891,In_608);
nand U785 (N_785,In_906,In_806);
xor U786 (N_786,In_68,In_1364);
nand U787 (N_787,In_1266,In_1773);
nand U788 (N_788,In_1775,In_1848);
xor U789 (N_789,In_805,In_822);
or U790 (N_790,In_1952,In_1869);
nor U791 (N_791,In_301,In_176);
nor U792 (N_792,In_367,In_895);
or U793 (N_793,In_1857,In_1389);
nand U794 (N_794,In_579,In_1983);
xnor U795 (N_795,In_247,In_1589);
or U796 (N_796,In_1281,In_476);
and U797 (N_797,In_96,In_1629);
xor U798 (N_798,In_118,In_946);
nor U799 (N_799,In_1270,In_803);
or U800 (N_800,In_99,In_933);
or U801 (N_801,In_835,In_1432);
nor U802 (N_802,In_423,In_382);
xnor U803 (N_803,In_1401,In_504);
nor U804 (N_804,In_148,In_753);
xor U805 (N_805,In_1421,In_638);
nand U806 (N_806,In_1990,In_894);
xor U807 (N_807,In_1116,In_1100);
nor U808 (N_808,In_1258,In_1740);
nor U809 (N_809,In_265,In_1374);
nor U810 (N_810,In_1986,In_570);
nor U811 (N_811,In_1413,In_1182);
or U812 (N_812,In_480,In_1656);
xnor U813 (N_813,In_1980,In_327);
xor U814 (N_814,In_245,In_315);
or U815 (N_815,In_1110,In_1511);
xnor U816 (N_816,In_1846,In_487);
xnor U817 (N_817,In_159,In_1662);
or U818 (N_818,In_573,In_1858);
or U819 (N_819,In_1338,In_420);
or U820 (N_820,In_1883,In_1320);
nand U821 (N_821,In_1653,In_732);
nor U822 (N_822,In_166,In_39);
or U823 (N_823,In_457,In_187);
and U824 (N_824,In_1262,In_1794);
nand U825 (N_825,In_1619,In_993);
or U826 (N_826,In_94,In_604);
and U827 (N_827,In_3,In_235);
nand U828 (N_828,In_1138,In_1844);
xor U829 (N_829,In_1119,In_914);
xor U830 (N_830,In_232,In_1642);
nand U831 (N_831,In_278,In_369);
xnor U832 (N_832,In_1514,In_1900);
and U833 (N_833,In_234,In_1345);
nor U834 (N_834,In_1780,In_1860);
nand U835 (N_835,In_1452,In_1493);
xnor U836 (N_836,In_653,In_502);
xor U837 (N_837,In_1103,In_1872);
nor U838 (N_838,In_631,In_237);
or U839 (N_839,In_600,In_515);
and U840 (N_840,In_1007,In_687);
nor U841 (N_841,In_1982,In_1588);
or U842 (N_842,In_1874,In_291);
xor U843 (N_843,In_964,In_1371);
or U844 (N_844,In_1516,In_1237);
nand U845 (N_845,In_1473,In_1286);
or U846 (N_846,In_1127,In_95);
nor U847 (N_847,In_744,In_158);
xor U848 (N_848,In_1536,In_1126);
nand U849 (N_849,In_1576,In_425);
nand U850 (N_850,In_1443,In_745);
or U851 (N_851,In_1423,In_92);
nor U852 (N_852,In_718,In_1031);
nor U853 (N_853,In_432,In_1593);
and U854 (N_854,In_1737,In_1300);
nor U855 (N_855,In_1144,In_746);
and U856 (N_856,In_1766,In_115);
nand U857 (N_857,In_908,In_755);
and U858 (N_858,In_538,In_1763);
or U859 (N_859,In_712,In_1080);
or U860 (N_860,In_861,In_433);
xor U861 (N_861,In_1689,In_238);
and U862 (N_862,In_649,In_758);
nand U863 (N_863,In_680,In_535);
and U864 (N_864,In_1384,In_544);
nor U865 (N_865,In_314,In_1165);
nand U866 (N_866,In_1596,In_1367);
nor U867 (N_867,In_776,In_1232);
nor U868 (N_868,In_1969,In_44);
or U869 (N_869,In_930,In_646);
nor U870 (N_870,In_1935,In_1777);
and U871 (N_871,In_715,In_706);
or U872 (N_872,In_162,In_705);
xnor U873 (N_873,In_482,In_1543);
xnor U874 (N_874,In_368,In_4);
nand U875 (N_875,In_1179,In_1359);
nor U876 (N_876,In_1096,In_1640);
and U877 (N_877,In_520,In_1092);
or U878 (N_878,In_1189,In_31);
and U879 (N_879,In_1855,In_667);
xor U880 (N_880,In_1828,In_184);
and U881 (N_881,In_1152,In_206);
or U882 (N_882,In_1625,In_542);
xnor U883 (N_883,In_1607,In_1229);
or U884 (N_884,In_730,In_1820);
xnor U885 (N_885,In_851,In_1436);
nand U886 (N_886,In_1008,In_380);
xnor U887 (N_887,In_129,In_1368);
nor U888 (N_888,In_8,In_843);
xnor U889 (N_889,In_881,In_1453);
nor U890 (N_890,In_1172,In_566);
and U891 (N_891,In_1416,In_224);
and U892 (N_892,In_1183,In_472);
nor U893 (N_893,In_1390,In_1224);
xnor U894 (N_894,In_514,In_1449);
nand U895 (N_895,In_413,In_143);
nand U896 (N_896,In_1666,In_752);
xnor U897 (N_897,In_1016,In_1201);
xnor U898 (N_898,In_968,In_1109);
nand U899 (N_899,In_1805,In_359);
xnor U900 (N_900,In_1244,In_1538);
or U901 (N_901,In_60,In_1690);
nor U902 (N_902,In_824,In_1798);
xnor U903 (N_903,In_1348,In_983);
xor U904 (N_904,In_1749,In_473);
nor U905 (N_905,In_1117,In_801);
nor U906 (N_906,In_828,In_371);
nor U907 (N_907,In_774,In_416);
xnor U908 (N_908,In_1618,In_293);
and U909 (N_909,In_1243,In_1011);
nor U910 (N_910,In_1620,In_211);
or U911 (N_911,In_393,In_1672);
and U912 (N_912,In_1603,In_921);
nand U913 (N_913,In_272,In_1804);
xor U914 (N_914,In_704,In_1329);
and U915 (N_915,In_346,In_1106);
xor U916 (N_916,In_1414,In_1216);
or U917 (N_917,In_641,In_209);
or U918 (N_918,In_597,In_437);
or U919 (N_919,In_1519,In_567);
xnor U920 (N_920,In_1290,In_890);
and U921 (N_921,In_1163,In_337);
nor U922 (N_922,In_1985,In_1515);
nand U923 (N_923,In_164,In_442);
or U924 (N_924,In_217,In_1899);
or U925 (N_925,In_685,In_1960);
nand U926 (N_926,In_589,In_911);
xor U927 (N_927,In_771,In_183);
xnor U928 (N_928,In_1962,In_1135);
nand U929 (N_929,In_1050,In_1197);
or U930 (N_930,In_901,In_1175);
and U931 (N_931,In_734,In_1036);
and U932 (N_932,In_1660,In_530);
or U933 (N_933,In_592,In_858);
xor U934 (N_934,In_1570,In_794);
nor U935 (N_935,In_1746,In_883);
nand U936 (N_936,In_1795,In_1481);
or U937 (N_937,In_1788,In_875);
nor U938 (N_938,In_686,In_182);
nor U939 (N_939,In_1451,In_56);
nand U940 (N_940,In_358,In_839);
xor U941 (N_941,In_910,In_617);
nand U942 (N_942,In_832,In_859);
nor U943 (N_943,In_59,In_1240);
and U944 (N_944,In_1111,In_271);
xor U945 (N_945,In_0,In_764);
or U946 (N_946,In_887,In_1586);
and U947 (N_947,In_947,In_412);
and U948 (N_948,In_1177,In_1887);
and U949 (N_949,In_36,In_1832);
and U950 (N_950,In_1132,In_105);
nand U951 (N_951,In_1856,In_388);
or U952 (N_952,In_1987,In_873);
nor U953 (N_953,In_1527,In_334);
xnor U954 (N_954,In_1334,In_586);
xor U955 (N_955,In_1044,In_112);
and U956 (N_956,In_1267,In_1722);
xnor U957 (N_957,In_62,In_1630);
or U958 (N_958,In_450,In_135);
xor U959 (N_959,In_651,In_1006);
or U960 (N_960,In_1492,In_2);
nand U961 (N_961,In_1272,In_533);
or U962 (N_962,In_988,In_185);
or U963 (N_963,In_1909,In_21);
nor U964 (N_964,In_1757,In_546);
nand U965 (N_965,In_417,In_1645);
nand U966 (N_966,In_355,In_1867);
nand U967 (N_967,In_1332,In_1606);
xor U968 (N_968,In_1904,In_751);
and U969 (N_969,In_1204,In_1076);
nand U970 (N_970,In_249,In_690);
xnor U971 (N_971,In_596,In_284);
and U972 (N_972,In_1651,In_547);
and U973 (N_973,In_379,In_572);
or U974 (N_974,In_466,In_818);
nand U975 (N_975,In_1702,In_1308);
or U976 (N_976,In_1455,In_691);
and U977 (N_977,In_282,In_456);
nor U978 (N_978,In_1800,In_179);
nand U979 (N_979,In_791,In_1786);
xnor U980 (N_980,In_656,In_532);
or U981 (N_981,In_381,In_1155);
nor U982 (N_982,In_190,In_637);
nand U983 (N_983,In_763,In_1158);
nand U984 (N_984,In_1681,In_584);
nand U985 (N_985,In_878,In_621);
nand U986 (N_986,In_399,In_601);
xnor U987 (N_987,In_720,In_816);
and U988 (N_988,In_1970,In_1318);
and U989 (N_989,In_902,In_131);
nor U990 (N_990,In_552,In_1841);
or U991 (N_991,In_133,In_1203);
nand U992 (N_992,In_1699,In_1810);
and U993 (N_993,In_1168,In_409);
and U994 (N_994,In_577,In_1360);
xnor U995 (N_995,In_870,In_1598);
nand U996 (N_996,In_1953,In_42);
xnor U997 (N_997,In_253,In_723);
nor U998 (N_998,In_307,In_784);
and U999 (N_999,In_1060,In_1397);
and U1000 (N_1000,In_390,In_483);
xnor U1001 (N_1001,In_1785,In_1123);
nor U1002 (N_1002,In_1971,In_21);
nand U1003 (N_1003,In_125,In_1579);
nor U1004 (N_1004,In_913,In_528);
or U1005 (N_1005,In_258,In_1737);
nor U1006 (N_1006,In_294,In_1615);
or U1007 (N_1007,In_1697,In_1456);
nand U1008 (N_1008,In_1335,In_1456);
and U1009 (N_1009,In_1086,In_661);
nand U1010 (N_1010,In_207,In_134);
nand U1011 (N_1011,In_1015,In_1801);
nand U1012 (N_1012,In_42,In_47);
xor U1013 (N_1013,In_1830,In_706);
or U1014 (N_1014,In_935,In_124);
xnor U1015 (N_1015,In_54,In_1097);
or U1016 (N_1016,In_1999,In_365);
xor U1017 (N_1017,In_1380,In_1177);
nand U1018 (N_1018,In_386,In_1706);
and U1019 (N_1019,In_21,In_1867);
and U1020 (N_1020,In_853,In_1472);
and U1021 (N_1021,In_305,In_1175);
or U1022 (N_1022,In_1025,In_1357);
nand U1023 (N_1023,In_490,In_1237);
or U1024 (N_1024,In_812,In_1584);
or U1025 (N_1025,In_1787,In_1712);
xor U1026 (N_1026,In_1851,In_381);
or U1027 (N_1027,In_68,In_1865);
and U1028 (N_1028,In_1059,In_1755);
nor U1029 (N_1029,In_849,In_655);
and U1030 (N_1030,In_1825,In_1584);
or U1031 (N_1031,In_1580,In_594);
and U1032 (N_1032,In_1295,In_906);
nor U1033 (N_1033,In_715,In_789);
or U1034 (N_1034,In_467,In_843);
or U1035 (N_1035,In_1962,In_1014);
nand U1036 (N_1036,In_1291,In_44);
or U1037 (N_1037,In_551,In_1109);
and U1038 (N_1038,In_1152,In_1268);
and U1039 (N_1039,In_143,In_1211);
xnor U1040 (N_1040,In_1189,In_996);
xor U1041 (N_1041,In_472,In_528);
xnor U1042 (N_1042,In_678,In_1823);
nand U1043 (N_1043,In_740,In_1525);
xnor U1044 (N_1044,In_569,In_637);
nand U1045 (N_1045,In_900,In_318);
or U1046 (N_1046,In_1929,In_511);
or U1047 (N_1047,In_1521,In_1417);
xor U1048 (N_1048,In_1844,In_981);
nor U1049 (N_1049,In_1083,In_344);
and U1050 (N_1050,In_81,In_1311);
and U1051 (N_1051,In_329,In_1279);
nand U1052 (N_1052,In_1843,In_1089);
nand U1053 (N_1053,In_1866,In_676);
nand U1054 (N_1054,In_78,In_222);
and U1055 (N_1055,In_46,In_1227);
and U1056 (N_1056,In_711,In_556);
or U1057 (N_1057,In_1698,In_431);
nor U1058 (N_1058,In_540,In_123);
or U1059 (N_1059,In_1906,In_1986);
nor U1060 (N_1060,In_195,In_1273);
nor U1061 (N_1061,In_1749,In_1340);
or U1062 (N_1062,In_386,In_205);
and U1063 (N_1063,In_1207,In_1648);
and U1064 (N_1064,In_1296,In_340);
nand U1065 (N_1065,In_940,In_180);
nor U1066 (N_1066,In_822,In_1270);
xnor U1067 (N_1067,In_923,In_1758);
xnor U1068 (N_1068,In_1096,In_1262);
xnor U1069 (N_1069,In_1478,In_245);
and U1070 (N_1070,In_1194,In_642);
xnor U1071 (N_1071,In_1426,In_414);
nand U1072 (N_1072,In_1459,In_1718);
or U1073 (N_1073,In_507,In_1008);
or U1074 (N_1074,In_1134,In_1427);
xnor U1075 (N_1075,In_1493,In_1000);
and U1076 (N_1076,In_1341,In_1672);
xor U1077 (N_1077,In_1700,In_1210);
and U1078 (N_1078,In_733,In_54);
and U1079 (N_1079,In_713,In_523);
nor U1080 (N_1080,In_564,In_218);
and U1081 (N_1081,In_325,In_1663);
xnor U1082 (N_1082,In_1747,In_1005);
nand U1083 (N_1083,In_942,In_1786);
and U1084 (N_1084,In_380,In_698);
nand U1085 (N_1085,In_653,In_801);
xnor U1086 (N_1086,In_1949,In_1753);
xnor U1087 (N_1087,In_888,In_1583);
and U1088 (N_1088,In_1956,In_1502);
xor U1089 (N_1089,In_53,In_556);
xnor U1090 (N_1090,In_1497,In_719);
nand U1091 (N_1091,In_1538,In_1362);
nor U1092 (N_1092,In_1908,In_1685);
nor U1093 (N_1093,In_1203,In_1718);
nand U1094 (N_1094,In_492,In_1157);
nand U1095 (N_1095,In_1418,In_1229);
xnor U1096 (N_1096,In_438,In_1698);
xor U1097 (N_1097,In_144,In_447);
and U1098 (N_1098,In_1569,In_1416);
and U1099 (N_1099,In_116,In_1929);
and U1100 (N_1100,In_1624,In_1744);
nand U1101 (N_1101,In_1823,In_1409);
nor U1102 (N_1102,In_1871,In_1716);
nor U1103 (N_1103,In_1343,In_1002);
xor U1104 (N_1104,In_1625,In_1794);
xnor U1105 (N_1105,In_1130,In_1088);
nand U1106 (N_1106,In_1937,In_955);
xor U1107 (N_1107,In_1002,In_218);
or U1108 (N_1108,In_1226,In_1425);
and U1109 (N_1109,In_634,In_1588);
or U1110 (N_1110,In_1744,In_936);
nand U1111 (N_1111,In_1017,In_1780);
nor U1112 (N_1112,In_1839,In_69);
or U1113 (N_1113,In_599,In_897);
or U1114 (N_1114,In_290,In_164);
xor U1115 (N_1115,In_759,In_1491);
nand U1116 (N_1116,In_861,In_533);
nor U1117 (N_1117,In_1028,In_1013);
nand U1118 (N_1118,In_1670,In_1976);
xor U1119 (N_1119,In_1122,In_783);
nand U1120 (N_1120,In_485,In_561);
or U1121 (N_1121,In_255,In_296);
nor U1122 (N_1122,In_224,In_826);
or U1123 (N_1123,In_855,In_1849);
xnor U1124 (N_1124,In_861,In_893);
xor U1125 (N_1125,In_247,In_745);
nor U1126 (N_1126,In_1676,In_1475);
nor U1127 (N_1127,In_1058,In_1238);
xnor U1128 (N_1128,In_323,In_351);
or U1129 (N_1129,In_825,In_667);
nand U1130 (N_1130,In_1901,In_1996);
nand U1131 (N_1131,In_902,In_1513);
or U1132 (N_1132,In_708,In_432);
or U1133 (N_1133,In_1755,In_586);
or U1134 (N_1134,In_977,In_505);
nor U1135 (N_1135,In_581,In_1810);
nand U1136 (N_1136,In_1358,In_107);
xnor U1137 (N_1137,In_618,In_30);
nand U1138 (N_1138,In_853,In_1419);
xor U1139 (N_1139,In_1675,In_1599);
nand U1140 (N_1140,In_125,In_510);
nor U1141 (N_1141,In_1618,In_1877);
nor U1142 (N_1142,In_578,In_1211);
nand U1143 (N_1143,In_780,In_1523);
nand U1144 (N_1144,In_978,In_236);
nand U1145 (N_1145,In_520,In_1575);
nand U1146 (N_1146,In_973,In_1991);
nand U1147 (N_1147,In_778,In_1871);
or U1148 (N_1148,In_15,In_1239);
nor U1149 (N_1149,In_167,In_1223);
nand U1150 (N_1150,In_828,In_348);
nor U1151 (N_1151,In_779,In_1476);
nand U1152 (N_1152,In_395,In_607);
nand U1153 (N_1153,In_837,In_912);
nand U1154 (N_1154,In_757,In_1001);
xnor U1155 (N_1155,In_1863,In_227);
or U1156 (N_1156,In_890,In_523);
and U1157 (N_1157,In_1041,In_1833);
or U1158 (N_1158,In_443,In_447);
nand U1159 (N_1159,In_1376,In_347);
and U1160 (N_1160,In_1557,In_430);
xnor U1161 (N_1161,In_266,In_1736);
xor U1162 (N_1162,In_1009,In_709);
or U1163 (N_1163,In_1653,In_1814);
and U1164 (N_1164,In_1641,In_523);
and U1165 (N_1165,In_353,In_1392);
and U1166 (N_1166,In_1291,In_1955);
nor U1167 (N_1167,In_1329,In_645);
nand U1168 (N_1168,In_532,In_38);
or U1169 (N_1169,In_490,In_1198);
nand U1170 (N_1170,In_429,In_749);
and U1171 (N_1171,In_1183,In_1584);
or U1172 (N_1172,In_1813,In_108);
and U1173 (N_1173,In_1464,In_818);
xor U1174 (N_1174,In_1160,In_1234);
or U1175 (N_1175,In_682,In_121);
or U1176 (N_1176,In_695,In_201);
nor U1177 (N_1177,In_355,In_1252);
or U1178 (N_1178,In_243,In_1306);
nand U1179 (N_1179,In_821,In_1569);
and U1180 (N_1180,In_1680,In_728);
xnor U1181 (N_1181,In_1619,In_1372);
and U1182 (N_1182,In_1463,In_412);
nand U1183 (N_1183,In_645,In_1308);
nand U1184 (N_1184,In_86,In_1102);
and U1185 (N_1185,In_426,In_654);
nand U1186 (N_1186,In_1917,In_1457);
xnor U1187 (N_1187,In_674,In_1793);
nor U1188 (N_1188,In_1500,In_1877);
and U1189 (N_1189,In_906,In_976);
and U1190 (N_1190,In_1256,In_1551);
nand U1191 (N_1191,In_1359,In_1296);
nand U1192 (N_1192,In_124,In_1864);
nor U1193 (N_1193,In_1142,In_440);
or U1194 (N_1194,In_888,In_127);
or U1195 (N_1195,In_1865,In_1087);
or U1196 (N_1196,In_1426,In_1356);
or U1197 (N_1197,In_939,In_1214);
nand U1198 (N_1198,In_1755,In_329);
xor U1199 (N_1199,In_427,In_1230);
and U1200 (N_1200,In_1400,In_924);
and U1201 (N_1201,In_574,In_1968);
and U1202 (N_1202,In_755,In_1438);
nor U1203 (N_1203,In_1916,In_1547);
nand U1204 (N_1204,In_1957,In_1120);
and U1205 (N_1205,In_1173,In_229);
xnor U1206 (N_1206,In_1549,In_1648);
nor U1207 (N_1207,In_887,In_1654);
or U1208 (N_1208,In_641,In_1771);
xor U1209 (N_1209,In_1565,In_1903);
nand U1210 (N_1210,In_1391,In_757);
or U1211 (N_1211,In_109,In_1866);
nand U1212 (N_1212,In_1615,In_776);
and U1213 (N_1213,In_1969,In_384);
xnor U1214 (N_1214,In_1461,In_1545);
and U1215 (N_1215,In_546,In_1416);
xor U1216 (N_1216,In_1509,In_87);
and U1217 (N_1217,In_1496,In_438);
xor U1218 (N_1218,In_823,In_221);
nor U1219 (N_1219,In_956,In_878);
and U1220 (N_1220,In_1109,In_1471);
nand U1221 (N_1221,In_1394,In_1918);
or U1222 (N_1222,In_263,In_1576);
nand U1223 (N_1223,In_1806,In_1177);
or U1224 (N_1224,In_670,In_1054);
xor U1225 (N_1225,In_372,In_1814);
or U1226 (N_1226,In_1799,In_205);
and U1227 (N_1227,In_416,In_722);
and U1228 (N_1228,In_363,In_1897);
nand U1229 (N_1229,In_1699,In_402);
and U1230 (N_1230,In_1082,In_533);
nor U1231 (N_1231,In_18,In_1077);
nor U1232 (N_1232,In_684,In_873);
or U1233 (N_1233,In_1318,In_37);
nor U1234 (N_1234,In_1289,In_986);
or U1235 (N_1235,In_1313,In_1417);
nor U1236 (N_1236,In_1186,In_282);
or U1237 (N_1237,In_1316,In_1283);
nor U1238 (N_1238,In_929,In_958);
xnor U1239 (N_1239,In_1368,In_1429);
nand U1240 (N_1240,In_1183,In_540);
and U1241 (N_1241,In_1964,In_1316);
and U1242 (N_1242,In_1067,In_96);
and U1243 (N_1243,In_1241,In_157);
xor U1244 (N_1244,In_935,In_383);
nand U1245 (N_1245,In_1003,In_310);
xor U1246 (N_1246,In_936,In_1977);
and U1247 (N_1247,In_172,In_439);
nor U1248 (N_1248,In_375,In_464);
nor U1249 (N_1249,In_1254,In_838);
nand U1250 (N_1250,In_1497,In_571);
xor U1251 (N_1251,In_610,In_264);
and U1252 (N_1252,In_687,In_1552);
and U1253 (N_1253,In_504,In_1968);
nor U1254 (N_1254,In_10,In_547);
xnor U1255 (N_1255,In_55,In_235);
xor U1256 (N_1256,In_765,In_1347);
xnor U1257 (N_1257,In_397,In_305);
nor U1258 (N_1258,In_1440,In_1225);
xor U1259 (N_1259,In_1594,In_1680);
nand U1260 (N_1260,In_1796,In_828);
nand U1261 (N_1261,In_58,In_1952);
nand U1262 (N_1262,In_1309,In_1994);
and U1263 (N_1263,In_1966,In_1239);
or U1264 (N_1264,In_878,In_1391);
xor U1265 (N_1265,In_330,In_1726);
nor U1266 (N_1266,In_523,In_13);
nor U1267 (N_1267,In_270,In_1611);
nand U1268 (N_1268,In_1716,In_275);
or U1269 (N_1269,In_145,In_63);
nor U1270 (N_1270,In_1860,In_284);
xor U1271 (N_1271,In_792,In_1094);
xor U1272 (N_1272,In_1500,In_1612);
xor U1273 (N_1273,In_1773,In_1092);
nand U1274 (N_1274,In_571,In_192);
xor U1275 (N_1275,In_965,In_784);
and U1276 (N_1276,In_1928,In_1872);
and U1277 (N_1277,In_280,In_1024);
nor U1278 (N_1278,In_1031,In_1506);
xnor U1279 (N_1279,In_901,In_1617);
xor U1280 (N_1280,In_1508,In_514);
nand U1281 (N_1281,In_623,In_767);
nor U1282 (N_1282,In_1591,In_428);
or U1283 (N_1283,In_1701,In_1619);
nand U1284 (N_1284,In_1317,In_132);
nor U1285 (N_1285,In_412,In_1460);
or U1286 (N_1286,In_1964,In_222);
and U1287 (N_1287,In_1726,In_1899);
xor U1288 (N_1288,In_1925,In_163);
nor U1289 (N_1289,In_1318,In_1657);
nand U1290 (N_1290,In_162,In_1872);
or U1291 (N_1291,In_1434,In_1338);
and U1292 (N_1292,In_986,In_1867);
nor U1293 (N_1293,In_1659,In_25);
or U1294 (N_1294,In_1402,In_1099);
nand U1295 (N_1295,In_640,In_269);
nand U1296 (N_1296,In_1289,In_1754);
xnor U1297 (N_1297,In_1452,In_837);
and U1298 (N_1298,In_595,In_708);
and U1299 (N_1299,In_837,In_1877);
and U1300 (N_1300,In_703,In_1969);
or U1301 (N_1301,In_1653,In_1214);
or U1302 (N_1302,In_362,In_1655);
nand U1303 (N_1303,In_794,In_530);
xor U1304 (N_1304,In_1606,In_625);
and U1305 (N_1305,In_385,In_1031);
xor U1306 (N_1306,In_1420,In_1480);
and U1307 (N_1307,In_463,In_171);
and U1308 (N_1308,In_653,In_1005);
nand U1309 (N_1309,In_1904,In_1285);
nand U1310 (N_1310,In_1995,In_1177);
nand U1311 (N_1311,In_1503,In_1281);
and U1312 (N_1312,In_1453,In_1501);
nand U1313 (N_1313,In_111,In_1655);
nand U1314 (N_1314,In_442,In_1641);
or U1315 (N_1315,In_1620,In_305);
nor U1316 (N_1316,In_919,In_872);
nand U1317 (N_1317,In_1953,In_1539);
nor U1318 (N_1318,In_1723,In_1901);
and U1319 (N_1319,In_0,In_1834);
nand U1320 (N_1320,In_362,In_95);
and U1321 (N_1321,In_1308,In_1798);
and U1322 (N_1322,In_156,In_1477);
xor U1323 (N_1323,In_332,In_828);
and U1324 (N_1324,In_74,In_1091);
xnor U1325 (N_1325,In_1032,In_1436);
nand U1326 (N_1326,In_1250,In_468);
xnor U1327 (N_1327,In_889,In_1542);
and U1328 (N_1328,In_197,In_1664);
nor U1329 (N_1329,In_502,In_1395);
and U1330 (N_1330,In_1179,In_1654);
and U1331 (N_1331,In_1020,In_920);
xnor U1332 (N_1332,In_6,In_686);
or U1333 (N_1333,In_447,In_483);
nand U1334 (N_1334,In_1862,In_1205);
xnor U1335 (N_1335,In_963,In_1638);
nand U1336 (N_1336,In_1786,In_644);
or U1337 (N_1337,In_1592,In_746);
nor U1338 (N_1338,In_1691,In_1136);
and U1339 (N_1339,In_281,In_235);
or U1340 (N_1340,In_1556,In_641);
or U1341 (N_1341,In_484,In_1167);
or U1342 (N_1342,In_1485,In_788);
and U1343 (N_1343,In_53,In_1164);
xor U1344 (N_1344,In_365,In_92);
or U1345 (N_1345,In_842,In_1142);
and U1346 (N_1346,In_1860,In_1231);
xor U1347 (N_1347,In_661,In_998);
and U1348 (N_1348,In_1994,In_1557);
and U1349 (N_1349,In_1639,In_1270);
nor U1350 (N_1350,In_1322,In_634);
xor U1351 (N_1351,In_423,In_148);
nor U1352 (N_1352,In_1165,In_46);
xor U1353 (N_1353,In_981,In_909);
nor U1354 (N_1354,In_264,In_1028);
nor U1355 (N_1355,In_1175,In_388);
nand U1356 (N_1356,In_208,In_1888);
or U1357 (N_1357,In_773,In_1585);
xor U1358 (N_1358,In_1310,In_1447);
nor U1359 (N_1359,In_1431,In_163);
nor U1360 (N_1360,In_1925,In_281);
or U1361 (N_1361,In_216,In_1904);
nand U1362 (N_1362,In_642,In_1228);
nand U1363 (N_1363,In_762,In_1869);
nor U1364 (N_1364,In_240,In_960);
xor U1365 (N_1365,In_1932,In_962);
or U1366 (N_1366,In_1698,In_1834);
xor U1367 (N_1367,In_1337,In_1576);
or U1368 (N_1368,In_1338,In_1295);
nand U1369 (N_1369,In_1578,In_884);
xor U1370 (N_1370,In_440,In_1906);
xor U1371 (N_1371,In_396,In_341);
nand U1372 (N_1372,In_1300,In_1259);
or U1373 (N_1373,In_665,In_327);
or U1374 (N_1374,In_702,In_1554);
nor U1375 (N_1375,In_692,In_482);
nand U1376 (N_1376,In_700,In_1872);
and U1377 (N_1377,In_115,In_1709);
nand U1378 (N_1378,In_207,In_1354);
xor U1379 (N_1379,In_512,In_1684);
xnor U1380 (N_1380,In_539,In_1131);
xnor U1381 (N_1381,In_256,In_1840);
nor U1382 (N_1382,In_790,In_1689);
and U1383 (N_1383,In_1606,In_212);
xor U1384 (N_1384,In_1636,In_692);
and U1385 (N_1385,In_123,In_1615);
nor U1386 (N_1386,In_786,In_1421);
nor U1387 (N_1387,In_1659,In_1531);
or U1388 (N_1388,In_1943,In_1335);
or U1389 (N_1389,In_308,In_260);
or U1390 (N_1390,In_141,In_321);
nand U1391 (N_1391,In_109,In_699);
and U1392 (N_1392,In_1520,In_1736);
nor U1393 (N_1393,In_877,In_1691);
or U1394 (N_1394,In_1680,In_641);
nand U1395 (N_1395,In_437,In_336);
or U1396 (N_1396,In_1163,In_575);
or U1397 (N_1397,In_71,In_1046);
or U1398 (N_1398,In_220,In_1460);
and U1399 (N_1399,In_880,In_38);
nand U1400 (N_1400,In_1649,In_1879);
nand U1401 (N_1401,In_867,In_1933);
xnor U1402 (N_1402,In_350,In_1554);
nand U1403 (N_1403,In_1471,In_1640);
nand U1404 (N_1404,In_1476,In_1556);
nand U1405 (N_1405,In_17,In_1886);
xor U1406 (N_1406,In_1779,In_1434);
nand U1407 (N_1407,In_1829,In_296);
xor U1408 (N_1408,In_1966,In_370);
nand U1409 (N_1409,In_1383,In_854);
xor U1410 (N_1410,In_1806,In_969);
or U1411 (N_1411,In_1809,In_22);
and U1412 (N_1412,In_259,In_1216);
xnor U1413 (N_1413,In_685,In_1179);
xor U1414 (N_1414,In_117,In_1369);
nand U1415 (N_1415,In_1464,In_873);
xor U1416 (N_1416,In_287,In_838);
xnor U1417 (N_1417,In_1494,In_120);
nand U1418 (N_1418,In_1612,In_123);
and U1419 (N_1419,In_1618,In_1600);
and U1420 (N_1420,In_1624,In_1743);
nor U1421 (N_1421,In_100,In_1911);
xor U1422 (N_1422,In_1605,In_1192);
or U1423 (N_1423,In_1401,In_722);
and U1424 (N_1424,In_424,In_106);
or U1425 (N_1425,In_1504,In_203);
nor U1426 (N_1426,In_64,In_243);
or U1427 (N_1427,In_893,In_847);
and U1428 (N_1428,In_454,In_1542);
nor U1429 (N_1429,In_1950,In_1102);
xnor U1430 (N_1430,In_473,In_703);
and U1431 (N_1431,In_1605,In_630);
xor U1432 (N_1432,In_793,In_1505);
nand U1433 (N_1433,In_169,In_1836);
and U1434 (N_1434,In_1414,In_1111);
nand U1435 (N_1435,In_1903,In_963);
and U1436 (N_1436,In_645,In_1391);
xnor U1437 (N_1437,In_360,In_1618);
nand U1438 (N_1438,In_439,In_332);
or U1439 (N_1439,In_940,In_1564);
nand U1440 (N_1440,In_1289,In_1938);
xnor U1441 (N_1441,In_1165,In_539);
xnor U1442 (N_1442,In_746,In_123);
nor U1443 (N_1443,In_1986,In_177);
nand U1444 (N_1444,In_28,In_731);
nor U1445 (N_1445,In_1582,In_268);
nor U1446 (N_1446,In_509,In_1946);
nand U1447 (N_1447,In_1956,In_55);
nor U1448 (N_1448,In_1018,In_912);
and U1449 (N_1449,In_1671,In_1031);
xor U1450 (N_1450,In_539,In_235);
and U1451 (N_1451,In_988,In_843);
xor U1452 (N_1452,In_113,In_1277);
nand U1453 (N_1453,In_1609,In_409);
nand U1454 (N_1454,In_330,In_1228);
or U1455 (N_1455,In_1282,In_1749);
nand U1456 (N_1456,In_14,In_294);
nor U1457 (N_1457,In_1233,In_812);
or U1458 (N_1458,In_966,In_5);
nand U1459 (N_1459,In_41,In_1918);
and U1460 (N_1460,In_1098,In_1224);
and U1461 (N_1461,In_1087,In_498);
xnor U1462 (N_1462,In_147,In_1866);
xor U1463 (N_1463,In_1297,In_1387);
and U1464 (N_1464,In_1696,In_501);
xnor U1465 (N_1465,In_1229,In_798);
and U1466 (N_1466,In_629,In_246);
nor U1467 (N_1467,In_102,In_1767);
and U1468 (N_1468,In_1632,In_153);
nand U1469 (N_1469,In_1999,In_371);
xnor U1470 (N_1470,In_725,In_15);
nor U1471 (N_1471,In_569,In_1131);
nand U1472 (N_1472,In_470,In_1824);
xor U1473 (N_1473,In_1965,In_120);
xnor U1474 (N_1474,In_1208,In_474);
nor U1475 (N_1475,In_1880,In_1729);
nand U1476 (N_1476,In_1052,In_1705);
xor U1477 (N_1477,In_697,In_1571);
nor U1478 (N_1478,In_427,In_1330);
xor U1479 (N_1479,In_174,In_1621);
nor U1480 (N_1480,In_1797,In_1186);
nand U1481 (N_1481,In_1466,In_355);
nor U1482 (N_1482,In_1966,In_1770);
nor U1483 (N_1483,In_988,In_695);
xnor U1484 (N_1484,In_901,In_1857);
or U1485 (N_1485,In_865,In_664);
and U1486 (N_1486,In_1565,In_1052);
nor U1487 (N_1487,In_324,In_1756);
nor U1488 (N_1488,In_1704,In_971);
xor U1489 (N_1489,In_699,In_906);
or U1490 (N_1490,In_707,In_576);
nand U1491 (N_1491,In_814,In_932);
nand U1492 (N_1492,In_83,In_1951);
and U1493 (N_1493,In_440,In_7);
or U1494 (N_1494,In_417,In_108);
xor U1495 (N_1495,In_281,In_650);
nand U1496 (N_1496,In_1650,In_1799);
xnor U1497 (N_1497,In_1340,In_578);
nand U1498 (N_1498,In_1024,In_455);
and U1499 (N_1499,In_1790,In_874);
or U1500 (N_1500,In_246,In_1737);
nand U1501 (N_1501,In_902,In_132);
and U1502 (N_1502,In_440,In_865);
and U1503 (N_1503,In_1436,In_202);
nand U1504 (N_1504,In_702,In_307);
nand U1505 (N_1505,In_965,In_1443);
nor U1506 (N_1506,In_1114,In_264);
and U1507 (N_1507,In_869,In_1931);
nand U1508 (N_1508,In_1136,In_1314);
nand U1509 (N_1509,In_1145,In_977);
nor U1510 (N_1510,In_1043,In_20);
nor U1511 (N_1511,In_1289,In_1852);
xor U1512 (N_1512,In_78,In_1846);
nor U1513 (N_1513,In_1070,In_1104);
nor U1514 (N_1514,In_1827,In_307);
or U1515 (N_1515,In_1606,In_329);
and U1516 (N_1516,In_1914,In_396);
nand U1517 (N_1517,In_1974,In_1954);
nand U1518 (N_1518,In_946,In_342);
xor U1519 (N_1519,In_1176,In_681);
nor U1520 (N_1520,In_1682,In_1143);
xnor U1521 (N_1521,In_75,In_785);
or U1522 (N_1522,In_1568,In_173);
nand U1523 (N_1523,In_1249,In_1443);
nand U1524 (N_1524,In_466,In_1360);
and U1525 (N_1525,In_1618,In_585);
nor U1526 (N_1526,In_1782,In_56);
xnor U1527 (N_1527,In_906,In_1807);
nor U1528 (N_1528,In_1533,In_1667);
xor U1529 (N_1529,In_811,In_1171);
nand U1530 (N_1530,In_1652,In_403);
and U1531 (N_1531,In_113,In_960);
xnor U1532 (N_1532,In_609,In_1684);
nor U1533 (N_1533,In_24,In_93);
xor U1534 (N_1534,In_1512,In_1798);
or U1535 (N_1535,In_1004,In_1444);
and U1536 (N_1536,In_1381,In_713);
xnor U1537 (N_1537,In_1150,In_1874);
xor U1538 (N_1538,In_649,In_260);
and U1539 (N_1539,In_1394,In_1726);
nor U1540 (N_1540,In_989,In_1845);
xnor U1541 (N_1541,In_1997,In_1728);
or U1542 (N_1542,In_1510,In_1600);
or U1543 (N_1543,In_1440,In_1015);
nand U1544 (N_1544,In_229,In_1685);
and U1545 (N_1545,In_1027,In_1799);
nor U1546 (N_1546,In_286,In_1305);
and U1547 (N_1547,In_1198,In_1105);
nand U1548 (N_1548,In_1719,In_1177);
and U1549 (N_1549,In_1033,In_1114);
and U1550 (N_1550,In_1400,In_1672);
nand U1551 (N_1551,In_1402,In_151);
or U1552 (N_1552,In_1258,In_798);
or U1553 (N_1553,In_840,In_1276);
nand U1554 (N_1554,In_1183,In_1482);
or U1555 (N_1555,In_1450,In_570);
nand U1556 (N_1556,In_756,In_1714);
nor U1557 (N_1557,In_1744,In_1137);
and U1558 (N_1558,In_1182,In_725);
xor U1559 (N_1559,In_1682,In_1759);
nor U1560 (N_1560,In_893,In_1981);
xor U1561 (N_1561,In_652,In_1127);
or U1562 (N_1562,In_439,In_1662);
xnor U1563 (N_1563,In_519,In_980);
xnor U1564 (N_1564,In_146,In_1320);
xor U1565 (N_1565,In_788,In_656);
xnor U1566 (N_1566,In_280,In_1058);
nor U1567 (N_1567,In_929,In_811);
and U1568 (N_1568,In_887,In_676);
nor U1569 (N_1569,In_406,In_1709);
xnor U1570 (N_1570,In_1582,In_1299);
nand U1571 (N_1571,In_526,In_607);
xnor U1572 (N_1572,In_1597,In_1639);
and U1573 (N_1573,In_1603,In_59);
and U1574 (N_1574,In_309,In_412);
xor U1575 (N_1575,In_1287,In_1566);
or U1576 (N_1576,In_1804,In_869);
and U1577 (N_1577,In_7,In_1785);
or U1578 (N_1578,In_243,In_1947);
xor U1579 (N_1579,In_259,In_1638);
nand U1580 (N_1580,In_640,In_657);
nor U1581 (N_1581,In_1097,In_1886);
xor U1582 (N_1582,In_1084,In_626);
and U1583 (N_1583,In_843,In_1626);
nand U1584 (N_1584,In_1207,In_1572);
and U1585 (N_1585,In_1226,In_1884);
or U1586 (N_1586,In_648,In_1560);
nor U1587 (N_1587,In_564,In_916);
and U1588 (N_1588,In_1323,In_1115);
and U1589 (N_1589,In_115,In_629);
and U1590 (N_1590,In_517,In_1162);
or U1591 (N_1591,In_1922,In_1225);
and U1592 (N_1592,In_615,In_1099);
and U1593 (N_1593,In_1416,In_199);
nor U1594 (N_1594,In_1531,In_497);
xnor U1595 (N_1595,In_1722,In_673);
xor U1596 (N_1596,In_1133,In_564);
and U1597 (N_1597,In_1959,In_184);
xor U1598 (N_1598,In_1532,In_1136);
nor U1599 (N_1599,In_205,In_701);
xnor U1600 (N_1600,In_1476,In_24);
xnor U1601 (N_1601,In_179,In_1183);
xnor U1602 (N_1602,In_1698,In_35);
nor U1603 (N_1603,In_1341,In_1117);
and U1604 (N_1604,In_1481,In_1325);
nand U1605 (N_1605,In_542,In_975);
nor U1606 (N_1606,In_1193,In_356);
xor U1607 (N_1607,In_1062,In_1692);
xor U1608 (N_1608,In_1645,In_194);
xnor U1609 (N_1609,In_1332,In_1883);
nor U1610 (N_1610,In_473,In_1266);
or U1611 (N_1611,In_1999,In_915);
and U1612 (N_1612,In_364,In_53);
nor U1613 (N_1613,In_1464,In_220);
or U1614 (N_1614,In_291,In_1416);
nor U1615 (N_1615,In_332,In_1939);
or U1616 (N_1616,In_1369,In_1790);
and U1617 (N_1617,In_921,In_1021);
nor U1618 (N_1618,In_1567,In_1377);
or U1619 (N_1619,In_1478,In_499);
xor U1620 (N_1620,In_927,In_358);
nand U1621 (N_1621,In_179,In_737);
xnor U1622 (N_1622,In_1750,In_1112);
xor U1623 (N_1623,In_770,In_733);
nand U1624 (N_1624,In_1273,In_891);
xor U1625 (N_1625,In_388,In_597);
or U1626 (N_1626,In_264,In_137);
and U1627 (N_1627,In_784,In_316);
nand U1628 (N_1628,In_1566,In_1201);
nand U1629 (N_1629,In_504,In_1687);
nor U1630 (N_1630,In_1283,In_1125);
and U1631 (N_1631,In_189,In_1159);
nor U1632 (N_1632,In_476,In_878);
nor U1633 (N_1633,In_967,In_771);
nor U1634 (N_1634,In_1031,In_988);
xor U1635 (N_1635,In_1689,In_430);
xnor U1636 (N_1636,In_26,In_213);
and U1637 (N_1637,In_538,In_328);
nand U1638 (N_1638,In_174,In_1238);
xnor U1639 (N_1639,In_1228,In_1059);
nor U1640 (N_1640,In_718,In_332);
and U1641 (N_1641,In_544,In_695);
and U1642 (N_1642,In_1907,In_1696);
xnor U1643 (N_1643,In_1910,In_463);
nand U1644 (N_1644,In_1325,In_1676);
nor U1645 (N_1645,In_1662,In_723);
xnor U1646 (N_1646,In_477,In_1405);
nor U1647 (N_1647,In_700,In_201);
and U1648 (N_1648,In_584,In_1356);
xnor U1649 (N_1649,In_1252,In_280);
nor U1650 (N_1650,In_1514,In_1573);
nor U1651 (N_1651,In_1871,In_187);
nor U1652 (N_1652,In_1459,In_77);
nand U1653 (N_1653,In_655,In_512);
or U1654 (N_1654,In_1545,In_1496);
nor U1655 (N_1655,In_1845,In_1005);
nand U1656 (N_1656,In_734,In_656);
nand U1657 (N_1657,In_455,In_789);
or U1658 (N_1658,In_390,In_1844);
nand U1659 (N_1659,In_459,In_630);
nor U1660 (N_1660,In_1869,In_267);
xor U1661 (N_1661,In_1763,In_1422);
xor U1662 (N_1662,In_981,In_1005);
xnor U1663 (N_1663,In_351,In_1850);
nor U1664 (N_1664,In_1554,In_803);
nand U1665 (N_1665,In_1126,In_1491);
nand U1666 (N_1666,In_1286,In_1556);
or U1667 (N_1667,In_376,In_117);
or U1668 (N_1668,In_1034,In_1898);
nand U1669 (N_1669,In_287,In_995);
or U1670 (N_1670,In_1652,In_1301);
nor U1671 (N_1671,In_560,In_901);
xor U1672 (N_1672,In_374,In_1925);
xor U1673 (N_1673,In_988,In_1956);
or U1674 (N_1674,In_1588,In_832);
nor U1675 (N_1675,In_580,In_1725);
and U1676 (N_1676,In_1372,In_1141);
xnor U1677 (N_1677,In_1285,In_1754);
xnor U1678 (N_1678,In_687,In_640);
xor U1679 (N_1679,In_1683,In_1913);
or U1680 (N_1680,In_1929,In_1759);
or U1681 (N_1681,In_11,In_912);
nand U1682 (N_1682,In_1395,In_1380);
and U1683 (N_1683,In_1696,In_185);
xnor U1684 (N_1684,In_1424,In_1279);
xnor U1685 (N_1685,In_30,In_1921);
xnor U1686 (N_1686,In_88,In_547);
and U1687 (N_1687,In_780,In_282);
or U1688 (N_1688,In_1229,In_295);
nor U1689 (N_1689,In_764,In_143);
nor U1690 (N_1690,In_1102,In_51);
and U1691 (N_1691,In_771,In_21);
and U1692 (N_1692,In_891,In_1535);
nor U1693 (N_1693,In_1040,In_223);
xnor U1694 (N_1694,In_1389,In_1063);
and U1695 (N_1695,In_643,In_1704);
xor U1696 (N_1696,In_450,In_37);
and U1697 (N_1697,In_211,In_1850);
or U1698 (N_1698,In_1491,In_455);
or U1699 (N_1699,In_1132,In_481);
nand U1700 (N_1700,In_240,In_1641);
nor U1701 (N_1701,In_1685,In_1509);
nor U1702 (N_1702,In_1212,In_1392);
nor U1703 (N_1703,In_236,In_862);
or U1704 (N_1704,In_534,In_985);
and U1705 (N_1705,In_566,In_579);
and U1706 (N_1706,In_1385,In_1411);
or U1707 (N_1707,In_1402,In_1421);
and U1708 (N_1708,In_1144,In_164);
nand U1709 (N_1709,In_1929,In_1805);
nor U1710 (N_1710,In_22,In_1886);
nor U1711 (N_1711,In_1257,In_630);
or U1712 (N_1712,In_727,In_1735);
nor U1713 (N_1713,In_185,In_1687);
nand U1714 (N_1714,In_1856,In_689);
nor U1715 (N_1715,In_680,In_1210);
nor U1716 (N_1716,In_1136,In_70);
nand U1717 (N_1717,In_1878,In_702);
or U1718 (N_1718,In_832,In_104);
xnor U1719 (N_1719,In_717,In_1982);
or U1720 (N_1720,In_1675,In_1936);
and U1721 (N_1721,In_430,In_1788);
xor U1722 (N_1722,In_1491,In_850);
nor U1723 (N_1723,In_1875,In_1509);
xnor U1724 (N_1724,In_201,In_588);
nand U1725 (N_1725,In_759,In_1602);
xnor U1726 (N_1726,In_1307,In_1234);
and U1727 (N_1727,In_713,In_1991);
and U1728 (N_1728,In_565,In_1161);
xnor U1729 (N_1729,In_1328,In_716);
nand U1730 (N_1730,In_1218,In_1348);
or U1731 (N_1731,In_985,In_346);
and U1732 (N_1732,In_1014,In_1301);
nand U1733 (N_1733,In_105,In_420);
and U1734 (N_1734,In_1345,In_599);
xor U1735 (N_1735,In_672,In_293);
nor U1736 (N_1736,In_597,In_1982);
nor U1737 (N_1737,In_1548,In_549);
and U1738 (N_1738,In_845,In_1057);
nor U1739 (N_1739,In_1964,In_439);
xnor U1740 (N_1740,In_1092,In_438);
or U1741 (N_1741,In_1844,In_1597);
or U1742 (N_1742,In_87,In_196);
or U1743 (N_1743,In_212,In_739);
nor U1744 (N_1744,In_1617,In_1620);
xnor U1745 (N_1745,In_1880,In_1568);
nor U1746 (N_1746,In_580,In_59);
xnor U1747 (N_1747,In_192,In_1632);
xnor U1748 (N_1748,In_1440,In_1414);
and U1749 (N_1749,In_1283,In_1884);
nand U1750 (N_1750,In_991,In_1192);
and U1751 (N_1751,In_1718,In_1433);
nor U1752 (N_1752,In_235,In_1118);
xor U1753 (N_1753,In_290,In_1820);
nand U1754 (N_1754,In_472,In_896);
and U1755 (N_1755,In_42,In_302);
nand U1756 (N_1756,In_1025,In_851);
xor U1757 (N_1757,In_1936,In_1488);
xor U1758 (N_1758,In_1900,In_1899);
nand U1759 (N_1759,In_1240,In_857);
or U1760 (N_1760,In_1451,In_1005);
or U1761 (N_1761,In_128,In_1629);
nand U1762 (N_1762,In_604,In_1345);
nand U1763 (N_1763,In_1365,In_445);
or U1764 (N_1764,In_389,In_720);
and U1765 (N_1765,In_225,In_1701);
nor U1766 (N_1766,In_1035,In_1989);
or U1767 (N_1767,In_1199,In_271);
xnor U1768 (N_1768,In_742,In_90);
and U1769 (N_1769,In_1208,In_41);
nor U1770 (N_1770,In_425,In_1850);
or U1771 (N_1771,In_1851,In_1929);
and U1772 (N_1772,In_60,In_1776);
or U1773 (N_1773,In_783,In_1614);
and U1774 (N_1774,In_724,In_907);
and U1775 (N_1775,In_1417,In_728);
xor U1776 (N_1776,In_164,In_636);
nand U1777 (N_1777,In_641,In_1829);
or U1778 (N_1778,In_687,In_1106);
or U1779 (N_1779,In_1202,In_947);
nor U1780 (N_1780,In_1264,In_1770);
xor U1781 (N_1781,In_59,In_701);
or U1782 (N_1782,In_484,In_1903);
and U1783 (N_1783,In_553,In_1888);
nor U1784 (N_1784,In_1864,In_587);
or U1785 (N_1785,In_438,In_571);
or U1786 (N_1786,In_617,In_1301);
xnor U1787 (N_1787,In_78,In_387);
xor U1788 (N_1788,In_1760,In_925);
nor U1789 (N_1789,In_11,In_466);
nor U1790 (N_1790,In_1414,In_1966);
xor U1791 (N_1791,In_1529,In_646);
or U1792 (N_1792,In_1360,In_854);
xnor U1793 (N_1793,In_757,In_1455);
nand U1794 (N_1794,In_1552,In_1727);
nand U1795 (N_1795,In_514,In_96);
and U1796 (N_1796,In_1752,In_232);
nand U1797 (N_1797,In_1585,In_705);
nor U1798 (N_1798,In_937,In_1237);
nor U1799 (N_1799,In_1427,In_992);
and U1800 (N_1800,In_1988,In_1134);
nor U1801 (N_1801,In_308,In_98);
nor U1802 (N_1802,In_892,In_285);
and U1803 (N_1803,In_1258,In_907);
or U1804 (N_1804,In_1445,In_774);
xor U1805 (N_1805,In_1897,In_1695);
nand U1806 (N_1806,In_888,In_1634);
nor U1807 (N_1807,In_865,In_1002);
or U1808 (N_1808,In_1667,In_574);
and U1809 (N_1809,In_786,In_840);
nand U1810 (N_1810,In_708,In_1970);
nand U1811 (N_1811,In_300,In_1936);
nand U1812 (N_1812,In_595,In_1066);
nand U1813 (N_1813,In_1556,In_1953);
nand U1814 (N_1814,In_754,In_122);
nand U1815 (N_1815,In_1559,In_705);
xnor U1816 (N_1816,In_1126,In_1607);
and U1817 (N_1817,In_1095,In_575);
or U1818 (N_1818,In_253,In_1691);
or U1819 (N_1819,In_99,In_1972);
and U1820 (N_1820,In_1515,In_1182);
xnor U1821 (N_1821,In_14,In_1675);
nor U1822 (N_1822,In_221,In_1237);
nand U1823 (N_1823,In_1666,In_715);
xnor U1824 (N_1824,In_433,In_1520);
or U1825 (N_1825,In_617,In_598);
nand U1826 (N_1826,In_1994,In_408);
or U1827 (N_1827,In_1618,In_1263);
nor U1828 (N_1828,In_1773,In_158);
nor U1829 (N_1829,In_841,In_1518);
nor U1830 (N_1830,In_1477,In_1352);
nor U1831 (N_1831,In_1531,In_1239);
nor U1832 (N_1832,In_1313,In_1728);
or U1833 (N_1833,In_12,In_534);
nand U1834 (N_1834,In_245,In_1538);
nor U1835 (N_1835,In_1338,In_35);
xor U1836 (N_1836,In_1242,In_537);
nand U1837 (N_1837,In_1448,In_56);
xnor U1838 (N_1838,In_381,In_27);
or U1839 (N_1839,In_1503,In_1685);
nor U1840 (N_1840,In_610,In_7);
nand U1841 (N_1841,In_1444,In_15);
nand U1842 (N_1842,In_1846,In_1528);
nand U1843 (N_1843,In_224,In_1277);
nor U1844 (N_1844,In_1506,In_1625);
and U1845 (N_1845,In_660,In_777);
and U1846 (N_1846,In_969,In_1720);
nand U1847 (N_1847,In_1257,In_532);
xor U1848 (N_1848,In_1195,In_1804);
nand U1849 (N_1849,In_126,In_488);
nor U1850 (N_1850,In_1186,In_1535);
nor U1851 (N_1851,In_44,In_457);
nor U1852 (N_1852,In_453,In_1269);
or U1853 (N_1853,In_1684,In_1578);
nor U1854 (N_1854,In_1016,In_399);
nand U1855 (N_1855,In_463,In_90);
xnor U1856 (N_1856,In_1611,In_109);
and U1857 (N_1857,In_1489,In_177);
or U1858 (N_1858,In_593,In_1670);
nand U1859 (N_1859,In_447,In_306);
nor U1860 (N_1860,In_1123,In_1324);
and U1861 (N_1861,In_108,In_1724);
xor U1862 (N_1862,In_768,In_1669);
nor U1863 (N_1863,In_1643,In_262);
xor U1864 (N_1864,In_77,In_1608);
or U1865 (N_1865,In_533,In_897);
xnor U1866 (N_1866,In_1017,In_1255);
or U1867 (N_1867,In_739,In_1925);
or U1868 (N_1868,In_432,In_902);
nand U1869 (N_1869,In_96,In_117);
or U1870 (N_1870,In_1878,In_892);
nand U1871 (N_1871,In_209,In_511);
and U1872 (N_1872,In_1808,In_1130);
xor U1873 (N_1873,In_1219,In_1184);
xor U1874 (N_1874,In_147,In_1715);
nand U1875 (N_1875,In_1748,In_397);
nand U1876 (N_1876,In_729,In_350);
or U1877 (N_1877,In_1586,In_693);
xnor U1878 (N_1878,In_37,In_590);
nor U1879 (N_1879,In_1372,In_863);
and U1880 (N_1880,In_1682,In_1813);
and U1881 (N_1881,In_344,In_1355);
or U1882 (N_1882,In_1325,In_607);
and U1883 (N_1883,In_1717,In_864);
nor U1884 (N_1884,In_716,In_935);
or U1885 (N_1885,In_1170,In_239);
xnor U1886 (N_1886,In_1280,In_1987);
xnor U1887 (N_1887,In_529,In_1808);
xnor U1888 (N_1888,In_1630,In_138);
nor U1889 (N_1889,In_201,In_495);
xor U1890 (N_1890,In_1044,In_1038);
nor U1891 (N_1891,In_1074,In_846);
xor U1892 (N_1892,In_107,In_1813);
and U1893 (N_1893,In_963,In_950);
and U1894 (N_1894,In_590,In_1098);
nor U1895 (N_1895,In_1944,In_1628);
xor U1896 (N_1896,In_1952,In_1223);
nand U1897 (N_1897,In_739,In_247);
or U1898 (N_1898,In_767,In_1104);
or U1899 (N_1899,In_1878,In_866);
nand U1900 (N_1900,In_1797,In_210);
nor U1901 (N_1901,In_232,In_238);
xor U1902 (N_1902,In_1420,In_100);
xor U1903 (N_1903,In_371,In_1941);
xor U1904 (N_1904,In_396,In_1808);
or U1905 (N_1905,In_462,In_132);
nand U1906 (N_1906,In_1222,In_1004);
xor U1907 (N_1907,In_1855,In_566);
nor U1908 (N_1908,In_833,In_717);
or U1909 (N_1909,In_1640,In_102);
and U1910 (N_1910,In_1290,In_1893);
nor U1911 (N_1911,In_755,In_182);
nand U1912 (N_1912,In_579,In_71);
and U1913 (N_1913,In_1521,In_718);
nor U1914 (N_1914,In_532,In_1723);
nor U1915 (N_1915,In_170,In_1998);
or U1916 (N_1916,In_141,In_81);
and U1917 (N_1917,In_1306,In_1597);
nand U1918 (N_1918,In_980,In_1807);
and U1919 (N_1919,In_982,In_608);
or U1920 (N_1920,In_888,In_913);
nand U1921 (N_1921,In_1314,In_1688);
xor U1922 (N_1922,In_888,In_1296);
and U1923 (N_1923,In_1962,In_818);
and U1924 (N_1924,In_386,In_1356);
xor U1925 (N_1925,In_1779,In_1121);
nor U1926 (N_1926,In_1325,In_1659);
xor U1927 (N_1927,In_1477,In_459);
nand U1928 (N_1928,In_37,In_1861);
or U1929 (N_1929,In_1352,In_592);
or U1930 (N_1930,In_1436,In_585);
or U1931 (N_1931,In_1566,In_1029);
or U1932 (N_1932,In_587,In_720);
and U1933 (N_1933,In_634,In_1188);
xnor U1934 (N_1934,In_1446,In_991);
nand U1935 (N_1935,In_119,In_1582);
nor U1936 (N_1936,In_976,In_1878);
or U1937 (N_1937,In_1727,In_256);
and U1938 (N_1938,In_1210,In_740);
and U1939 (N_1939,In_1983,In_217);
nand U1940 (N_1940,In_1307,In_1219);
or U1941 (N_1941,In_198,In_1578);
or U1942 (N_1942,In_1373,In_1422);
nor U1943 (N_1943,In_699,In_1132);
nand U1944 (N_1944,In_381,In_803);
or U1945 (N_1945,In_1323,In_1760);
and U1946 (N_1946,In_1726,In_1694);
xnor U1947 (N_1947,In_1904,In_1835);
and U1948 (N_1948,In_1498,In_15);
nor U1949 (N_1949,In_1360,In_748);
nand U1950 (N_1950,In_1313,In_1724);
xor U1951 (N_1951,In_1801,In_1984);
or U1952 (N_1952,In_1602,In_503);
nor U1953 (N_1953,In_35,In_231);
xnor U1954 (N_1954,In_57,In_840);
and U1955 (N_1955,In_1754,In_142);
and U1956 (N_1956,In_750,In_990);
or U1957 (N_1957,In_1870,In_1149);
xor U1958 (N_1958,In_1358,In_1725);
xor U1959 (N_1959,In_1987,In_180);
or U1960 (N_1960,In_1300,In_705);
or U1961 (N_1961,In_1876,In_1699);
nand U1962 (N_1962,In_384,In_1385);
nor U1963 (N_1963,In_898,In_760);
or U1964 (N_1964,In_391,In_1380);
or U1965 (N_1965,In_56,In_425);
and U1966 (N_1966,In_881,In_1442);
nor U1967 (N_1967,In_1487,In_248);
nand U1968 (N_1968,In_1628,In_340);
nor U1969 (N_1969,In_358,In_1241);
or U1970 (N_1970,In_1858,In_1296);
xnor U1971 (N_1971,In_842,In_205);
or U1972 (N_1972,In_818,In_157);
and U1973 (N_1973,In_1872,In_72);
or U1974 (N_1974,In_1171,In_1461);
and U1975 (N_1975,In_676,In_1526);
or U1976 (N_1976,In_1085,In_557);
nand U1977 (N_1977,In_3,In_1309);
nand U1978 (N_1978,In_819,In_57);
or U1979 (N_1979,In_1276,In_688);
and U1980 (N_1980,In_511,In_1107);
nand U1981 (N_1981,In_1482,In_1940);
nor U1982 (N_1982,In_1432,In_594);
nand U1983 (N_1983,In_1637,In_61);
xnor U1984 (N_1984,In_1715,In_734);
and U1985 (N_1985,In_1268,In_1845);
xnor U1986 (N_1986,In_86,In_1717);
and U1987 (N_1987,In_844,In_1607);
nand U1988 (N_1988,In_1028,In_516);
nand U1989 (N_1989,In_1695,In_455);
xnor U1990 (N_1990,In_1436,In_253);
nand U1991 (N_1991,In_1143,In_1990);
nor U1992 (N_1992,In_176,In_1130);
nand U1993 (N_1993,In_135,In_461);
nand U1994 (N_1994,In_1722,In_903);
or U1995 (N_1995,In_774,In_786);
xor U1996 (N_1996,In_1658,In_1948);
or U1997 (N_1997,In_1883,In_1567);
xnor U1998 (N_1998,In_700,In_782);
nor U1999 (N_1999,In_120,In_744);
nor U2000 (N_2000,N_61,N_1677);
and U2001 (N_2001,N_320,N_1261);
or U2002 (N_2002,N_1336,N_108);
xor U2003 (N_2003,N_1078,N_945);
xor U2004 (N_2004,N_275,N_272);
xor U2005 (N_2005,N_1787,N_1612);
nand U2006 (N_2006,N_1583,N_680);
or U2007 (N_2007,N_404,N_631);
and U2008 (N_2008,N_1609,N_1752);
nand U2009 (N_2009,N_258,N_106);
nand U2010 (N_2010,N_1150,N_1320);
xor U2011 (N_2011,N_1448,N_1420);
nand U2012 (N_2012,N_880,N_749);
xor U2013 (N_2013,N_122,N_1152);
nand U2014 (N_2014,N_1718,N_652);
nand U2015 (N_2015,N_530,N_1873);
and U2016 (N_2016,N_1364,N_1053);
or U2017 (N_2017,N_1490,N_1531);
or U2018 (N_2018,N_858,N_341);
or U2019 (N_2019,N_1138,N_725);
and U2020 (N_2020,N_940,N_1686);
and U2021 (N_2021,N_297,N_1333);
nand U2022 (N_2022,N_1041,N_635);
nand U2023 (N_2023,N_1253,N_529);
or U2024 (N_2024,N_954,N_1622);
xnor U2025 (N_2025,N_626,N_1780);
and U2026 (N_2026,N_864,N_797);
xor U2027 (N_2027,N_51,N_38);
xnor U2028 (N_2028,N_946,N_209);
and U2029 (N_2029,N_89,N_751);
nor U2030 (N_2030,N_1832,N_1514);
xor U2031 (N_2031,N_952,N_351);
or U2032 (N_2032,N_1380,N_1550);
xnor U2033 (N_2033,N_1808,N_687);
xnor U2034 (N_2034,N_1694,N_554);
xor U2035 (N_2035,N_644,N_845);
nor U2036 (N_2036,N_1696,N_746);
nand U2037 (N_2037,N_897,N_1123);
nand U2038 (N_2038,N_1613,N_212);
xor U2039 (N_2039,N_763,N_1203);
nor U2040 (N_2040,N_1049,N_618);
or U2041 (N_2041,N_1973,N_1265);
xor U2042 (N_2042,N_427,N_345);
xor U2043 (N_2043,N_1209,N_706);
nand U2044 (N_2044,N_1199,N_677);
xnor U2045 (N_2045,N_570,N_233);
and U2046 (N_2046,N_816,N_1865);
and U2047 (N_2047,N_1207,N_1857);
nand U2048 (N_2048,N_185,N_686);
nor U2049 (N_2049,N_484,N_616);
nand U2050 (N_2050,N_1652,N_1982);
or U2051 (N_2051,N_1515,N_741);
and U2052 (N_2052,N_1024,N_457);
or U2053 (N_2053,N_1487,N_338);
nor U2054 (N_2054,N_1169,N_558);
and U2055 (N_2055,N_443,N_1318);
and U2056 (N_2056,N_1640,N_1581);
xor U2057 (N_2057,N_1313,N_101);
xnor U2058 (N_2058,N_638,N_916);
and U2059 (N_2059,N_1451,N_761);
xnor U2060 (N_2060,N_1486,N_1941);
nand U2061 (N_2061,N_748,N_593);
xor U2062 (N_2062,N_164,N_302);
or U2063 (N_2063,N_1006,N_1903);
xor U2064 (N_2064,N_1863,N_823);
xnor U2065 (N_2065,N_17,N_736);
nand U2066 (N_2066,N_1356,N_1065);
xnor U2067 (N_2067,N_1171,N_1758);
xor U2068 (N_2068,N_1491,N_182);
and U2069 (N_2069,N_1061,N_1653);
nand U2070 (N_2070,N_572,N_1312);
xnor U2071 (N_2071,N_1461,N_1234);
and U2072 (N_2072,N_1258,N_1047);
and U2073 (N_2073,N_177,N_456);
nor U2074 (N_2074,N_278,N_1620);
nor U2075 (N_2075,N_970,N_1966);
and U2076 (N_2076,N_416,N_105);
or U2077 (N_2077,N_1409,N_1690);
and U2078 (N_2078,N_1423,N_1700);
nor U2079 (N_2079,N_1135,N_1034);
nand U2080 (N_2080,N_1990,N_811);
nor U2081 (N_2081,N_1554,N_1596);
and U2082 (N_2082,N_240,N_587);
xor U2083 (N_2083,N_401,N_664);
xor U2084 (N_2084,N_412,N_246);
or U2085 (N_2085,N_778,N_1826);
and U2086 (N_2086,N_1714,N_118);
nor U2087 (N_2087,N_1732,N_1761);
xnor U2088 (N_2088,N_228,N_1455);
xor U2089 (N_2089,N_1886,N_807);
nor U2090 (N_2090,N_1977,N_1287);
and U2091 (N_2091,N_1562,N_21);
nor U2092 (N_2092,N_1616,N_80);
nand U2093 (N_2093,N_773,N_1372);
nor U2094 (N_2094,N_1975,N_975);
nor U2095 (N_2095,N_1880,N_1172);
or U2096 (N_2096,N_1225,N_181);
nor U2097 (N_2097,N_1089,N_1481);
and U2098 (N_2098,N_413,N_1958);
nand U2099 (N_2099,N_1854,N_465);
xor U2100 (N_2100,N_1995,N_1556);
and U2101 (N_2101,N_1688,N_1501);
nor U2102 (N_2102,N_1631,N_204);
nor U2103 (N_2103,N_1391,N_1444);
nor U2104 (N_2104,N_0,N_1497);
or U2105 (N_2105,N_1870,N_422);
xnor U2106 (N_2106,N_301,N_1908);
and U2107 (N_2107,N_1155,N_727);
nand U2108 (N_2108,N_1248,N_1553);
or U2109 (N_2109,N_681,N_740);
nand U2110 (N_2110,N_260,N_1148);
and U2111 (N_2111,N_943,N_265);
nand U2112 (N_2112,N_1103,N_987);
and U2113 (N_2113,N_914,N_528);
and U2114 (N_2114,N_909,N_1713);
or U2115 (N_2115,N_728,N_1485);
nand U2116 (N_2116,N_678,N_565);
or U2117 (N_2117,N_1028,N_1750);
nor U2118 (N_2118,N_73,N_641);
or U2119 (N_2119,N_1608,N_460);
nand U2120 (N_2120,N_817,N_684);
and U2121 (N_2121,N_152,N_403);
or U2122 (N_2122,N_1195,N_515);
nand U2123 (N_2123,N_1347,N_601);
nor U2124 (N_2124,N_753,N_303);
nand U2125 (N_2125,N_1883,N_1915);
nor U2126 (N_2126,N_316,N_1228);
xor U2127 (N_2127,N_1840,N_1140);
or U2128 (N_2128,N_871,N_1416);
and U2129 (N_2129,N_6,N_332);
nor U2130 (N_2130,N_397,N_1378);
nor U2131 (N_2131,N_668,N_1370);
nor U2132 (N_2132,N_1398,N_659);
and U2133 (N_2133,N_1793,N_1593);
and U2134 (N_2134,N_1795,N_1799);
nor U2135 (N_2135,N_1587,N_969);
and U2136 (N_2136,N_1285,N_1949);
nand U2137 (N_2137,N_576,N_1104);
nand U2138 (N_2138,N_1937,N_155);
nand U2139 (N_2139,N_1101,N_1365);
nor U2140 (N_2140,N_1801,N_291);
nand U2141 (N_2141,N_64,N_1874);
nor U2142 (N_2142,N_474,N_733);
nand U2143 (N_2143,N_1842,N_436);
nor U2144 (N_2144,N_1022,N_206);
or U2145 (N_2145,N_653,N_508);
or U2146 (N_2146,N_178,N_1704);
and U2147 (N_2147,N_1746,N_1429);
nand U2148 (N_2148,N_785,N_649);
nor U2149 (N_2149,N_906,N_1030);
nor U2150 (N_2150,N_1316,N_514);
or U2151 (N_2151,N_1816,N_165);
or U2152 (N_2152,N_539,N_267);
or U2153 (N_2153,N_776,N_768);
nor U2154 (N_2154,N_1934,N_1067);
nand U2155 (N_2155,N_924,N_1557);
and U2156 (N_2156,N_1695,N_1633);
xor U2157 (N_2157,N_1667,N_4);
or U2158 (N_2158,N_802,N_578);
and U2159 (N_2159,N_113,N_1701);
xnor U2160 (N_2160,N_1406,N_1341);
nand U2161 (N_2161,N_990,N_1130);
or U2162 (N_2162,N_1668,N_167);
nor U2163 (N_2163,N_1379,N_435);
xor U2164 (N_2164,N_1764,N_657);
nor U2165 (N_2165,N_1855,N_1465);
or U2166 (N_2166,N_882,N_20);
and U2167 (N_2167,N_1721,N_1479);
nand U2168 (N_2168,N_1603,N_1950);
nor U2169 (N_2169,N_1196,N_1930);
xnor U2170 (N_2170,N_546,N_1456);
nor U2171 (N_2171,N_1584,N_663);
and U2172 (N_2172,N_82,N_1050);
nor U2173 (N_2173,N_770,N_1247);
nor U2174 (N_2174,N_1821,N_899);
nand U2175 (N_2175,N_1352,N_643);
nand U2176 (N_2176,N_679,N_561);
nor U2177 (N_2177,N_843,N_1021);
and U2178 (N_2178,N_1885,N_1951);
nand U2179 (N_2179,N_1805,N_1440);
nor U2180 (N_2180,N_1913,N_1529);
nand U2181 (N_2181,N_1566,N_229);
xor U2182 (N_2182,N_1804,N_1160);
xnor U2183 (N_2183,N_1670,N_900);
xor U2184 (N_2184,N_588,N_792);
nor U2185 (N_2185,N_1197,N_1322);
or U2186 (N_2186,N_1411,N_1710);
or U2187 (N_2187,N_138,N_518);
or U2188 (N_2188,N_314,N_1162);
or U2189 (N_2189,N_462,N_676);
nand U2190 (N_2190,N_1769,N_1093);
xnor U2191 (N_2191,N_550,N_1654);
nor U2192 (N_2192,N_1831,N_1290);
nand U2193 (N_2193,N_1575,N_488);
or U2194 (N_2194,N_1955,N_731);
nand U2195 (N_2195,N_473,N_451);
or U2196 (N_2196,N_1943,N_857);
xor U2197 (N_2197,N_415,N_148);
or U2198 (N_2198,N_1940,N_1295);
or U2199 (N_2199,N_1095,N_150);
nand U2200 (N_2200,N_1314,N_238);
or U2201 (N_2201,N_796,N_724);
nor U2202 (N_2202,N_949,N_926);
xor U2203 (N_2203,N_139,N_1549);
xor U2204 (N_2204,N_974,N_655);
and U2205 (N_2205,N_1102,N_375);
or U2206 (N_2206,N_1920,N_950);
xor U2207 (N_2207,N_1263,N_852);
nor U2208 (N_2208,N_222,N_188);
nand U2209 (N_2209,N_1499,N_1430);
xor U2210 (N_2210,N_1800,N_7);
or U2211 (N_2211,N_1747,N_344);
nor U2212 (N_2212,N_932,N_1590);
xnor U2213 (N_2213,N_389,N_1504);
nor U2214 (N_2214,N_931,N_1985);
nand U2215 (N_2215,N_68,N_690);
and U2216 (N_2216,N_1432,N_169);
nand U2217 (N_2217,N_266,N_1108);
nor U2218 (N_2218,N_1327,N_868);
or U2219 (N_2219,N_685,N_692);
xor U2220 (N_2220,N_311,N_1144);
and U2221 (N_2221,N_1981,N_771);
nand U2222 (N_2222,N_1588,N_1221);
nor U2223 (N_2223,N_1755,N_312);
or U2224 (N_2224,N_219,N_1473);
nor U2225 (N_2225,N_35,N_1509);
and U2226 (N_2226,N_119,N_476);
xor U2227 (N_2227,N_968,N_1214);
nor U2228 (N_2228,N_1879,N_720);
or U2229 (N_2229,N_170,N_767);
xor U2230 (N_2230,N_1905,N_750);
or U2231 (N_2231,N_22,N_1707);
nor U2232 (N_2232,N_1303,N_556);
xnor U2233 (N_2233,N_998,N_431);
xnor U2234 (N_2234,N_321,N_1099);
or U2235 (N_2235,N_56,N_1989);
nor U2236 (N_2236,N_501,N_1979);
nand U2237 (N_2237,N_1368,N_62);
nor U2238 (N_2238,N_840,N_1582);
or U2239 (N_2239,N_1773,N_1116);
xor U2240 (N_2240,N_854,N_1824);
or U2241 (N_2241,N_1656,N_1785);
or U2242 (N_2242,N_396,N_1904);
nand U2243 (N_2243,N_475,N_511);
and U2244 (N_2244,N_114,N_470);
and U2245 (N_2245,N_1781,N_699);
and U2246 (N_2246,N_509,N_205);
xnor U2247 (N_2247,N_149,N_83);
nand U2248 (N_2248,N_673,N_1968);
or U2249 (N_2249,N_617,N_377);
nand U2250 (N_2250,N_887,N_1991);
or U2251 (N_2251,N_42,N_446);
nor U2252 (N_2252,N_839,N_1643);
xor U2253 (N_2253,N_589,N_1993);
nand U2254 (N_2254,N_382,N_818);
nor U2255 (N_2255,N_1618,N_1117);
nand U2256 (N_2256,N_762,N_646);
nand U2257 (N_2257,N_1147,N_18);
and U2258 (N_2258,N_606,N_157);
nor U2259 (N_2259,N_1016,N_1572);
nand U2260 (N_2260,N_1462,N_45);
nor U2261 (N_2261,N_888,N_942);
nand U2262 (N_2262,N_1346,N_1646);
nor U2263 (N_2263,N_1107,N_1179);
xnor U2264 (N_2264,N_656,N_379);
xor U2265 (N_2265,N_1009,N_1133);
or U2266 (N_2266,N_709,N_1544);
or U2267 (N_2267,N_112,N_49);
and U2268 (N_2268,N_939,N_335);
xnor U2269 (N_2269,N_893,N_1308);
or U2270 (N_2270,N_1076,N_1177);
nor U2271 (N_2271,N_885,N_695);
or U2272 (N_2272,N_1924,N_1180);
xor U2273 (N_2273,N_1534,N_211);
and U2274 (N_2274,N_637,N_1530);
nand U2275 (N_2275,N_813,N_1453);
and U2276 (N_2276,N_1390,N_964);
and U2277 (N_2277,N_286,N_203);
nor U2278 (N_2278,N_594,N_3);
and U2279 (N_2279,N_1742,N_1252);
nor U2280 (N_2280,N_1242,N_195);
nand U2281 (N_2281,N_339,N_450);
nand U2282 (N_2282,N_1959,N_1273);
nand U2283 (N_2283,N_604,N_697);
nor U2284 (N_2284,N_775,N_147);
nand U2285 (N_2285,N_28,N_1829);
or U2286 (N_2286,N_1889,N_1141);
nor U2287 (N_2287,N_1579,N_689);
and U2288 (N_2288,N_1007,N_1326);
or U2289 (N_2289,N_1565,N_803);
and U2290 (N_2290,N_1510,N_1837);
xor U2291 (N_2291,N_911,N_534);
nand U2292 (N_2292,N_10,N_870);
xor U2293 (N_2293,N_959,N_1362);
nor U2294 (N_2294,N_394,N_1709);
or U2295 (N_2295,N_348,N_1118);
nand U2296 (N_2296,N_1743,N_1283);
or U2297 (N_2297,N_1216,N_116);
nor U2298 (N_2298,N_57,N_1426);
xnor U2299 (N_2299,N_1494,N_1843);
and U2300 (N_2300,N_598,N_1460);
and U2301 (N_2301,N_1875,N_1158);
and U2302 (N_2302,N_1794,N_694);
nor U2303 (N_2303,N_737,N_295);
nor U2304 (N_2304,N_1269,N_757);
nor U2305 (N_2305,N_1489,N_1676);
and U2306 (N_2306,N_756,N_904);
or U2307 (N_2307,N_300,N_322);
and U2308 (N_2308,N_1678,N_624);
nand U2309 (N_2309,N_1300,N_1035);
or U2310 (N_2310,N_134,N_513);
xor U2311 (N_2311,N_1422,N_779);
xor U2312 (N_2312,N_683,N_1080);
nor U2313 (N_2313,N_698,N_464);
and U2314 (N_2314,N_1703,N_1948);
and U2315 (N_2315,N_25,N_1627);
nand U2316 (N_2316,N_1286,N_1726);
or U2317 (N_2317,N_1001,N_128);
or U2318 (N_2318,N_77,N_11);
nand U2319 (N_2319,N_459,N_151);
nor U2320 (N_2320,N_1914,N_252);
xor U2321 (N_2321,N_244,N_1149);
xnor U2322 (N_2322,N_308,N_1017);
or U2323 (N_2323,N_292,N_787);
nand U2324 (N_2324,N_104,N_581);
xnor U2325 (N_2325,N_1784,N_1208);
and U2326 (N_2326,N_878,N_995);
nand U2327 (N_2327,N_1458,N_1896);
and U2328 (N_2328,N_279,N_726);
and U2329 (N_2329,N_1010,N_91);
nor U2330 (N_2330,N_1852,N_547);
or U2331 (N_2331,N_1776,N_795);
xor U2332 (N_2332,N_230,N_494);
nand U2333 (N_2333,N_1740,N_1847);
nor U2334 (N_2334,N_1675,N_1019);
and U2335 (N_2335,N_1639,N_1689);
and U2336 (N_2336,N_1483,N_154);
and U2337 (N_2337,N_1881,N_1057);
nand U2338 (N_2338,N_358,N_1340);
or U2339 (N_2339,N_745,N_1046);
and U2340 (N_2340,N_1292,N_1299);
xor U2341 (N_2341,N_548,N_283);
or U2342 (N_2342,N_304,N_960);
nor U2343 (N_2343,N_1815,N_962);
or U2344 (N_2344,N_1085,N_1827);
and U2345 (N_2345,N_1421,N_1988);
or U2346 (N_2346,N_1777,N_1381);
nand U2347 (N_2347,N_1888,N_1573);
or U2348 (N_2348,N_250,N_1906);
or U2349 (N_2349,N_1018,N_1239);
nand U2350 (N_2350,N_349,N_837);
or U2351 (N_2351,N_721,N_1268);
xnor U2352 (N_2352,N_1176,N_1728);
or U2353 (N_2353,N_1927,N_562);
xnor U2354 (N_2354,N_1305,N_859);
or U2355 (N_2355,N_1246,N_1054);
xor U2356 (N_2356,N_342,N_1111);
xor U2357 (N_2357,N_856,N_111);
or U2358 (N_2358,N_1122,N_1790);
nand U2359 (N_2359,N_898,N_956);
and U2360 (N_2360,N_1428,N_1386);
xor U2361 (N_2361,N_193,N_1436);
and U2362 (N_2362,N_1938,N_1056);
and U2363 (N_2363,N_281,N_1806);
or U2364 (N_2364,N_1139,N_237);
or U2365 (N_2365,N_1792,N_1545);
xnor U2366 (N_2366,N_936,N_850);
nand U2367 (N_2367,N_1164,N_809);
nor U2368 (N_2368,N_1224,N_1611);
or U2369 (N_2369,N_1860,N_1998);
nand U2370 (N_2370,N_471,N_1662);
xor U2371 (N_2371,N_433,N_538);
nor U2372 (N_2372,N_732,N_1297);
nor U2373 (N_2373,N_1516,N_1439);
nand U2374 (N_2374,N_674,N_235);
or U2375 (N_2375,N_325,N_1231);
or U2376 (N_2376,N_1963,N_1630);
nor U2377 (N_2377,N_1134,N_980);
and U2378 (N_2378,N_261,N_1745);
or U2379 (N_2379,N_248,N_497);
or U2380 (N_2380,N_754,N_1227);
nor U2381 (N_2381,N_55,N_1353);
xor U2382 (N_2382,N_1474,N_5);
xnor U2383 (N_2383,N_1232,N_1052);
or U2384 (N_2384,N_132,N_1559);
xor U2385 (N_2385,N_1454,N_506);
and U2386 (N_2386,N_52,N_1254);
nand U2387 (N_2387,N_365,N_407);
xor U2388 (N_2388,N_944,N_174);
or U2389 (N_2389,N_522,N_908);
and U2390 (N_2390,N_1508,N_1931);
nand U2391 (N_2391,N_876,N_1578);
xnor U2392 (N_2392,N_352,N_1674);
or U2393 (N_2393,N_1918,N_1450);
or U2394 (N_2394,N_1725,N_827);
and U2395 (N_2395,N_747,N_1729);
xnor U2396 (N_2396,N_1337,N_1218);
or U2397 (N_2397,N_253,N_996);
nor U2398 (N_2398,N_1763,N_1110);
xor U2399 (N_2399,N_1532,N_227);
nand U2400 (N_2400,N_665,N_1217);
nand U2401 (N_2401,N_120,N_1418);
xnor U2402 (N_2402,N_1468,N_1962);
or U2403 (N_2403,N_1774,N_1038);
and U2404 (N_2404,N_1614,N_48);
or U2405 (N_2405,N_1833,N_1797);
or U2406 (N_2406,N_429,N_221);
xor U2407 (N_2407,N_1778,N_444);
and U2408 (N_2408,N_140,N_866);
nand U2409 (N_2409,N_202,N_715);
and U2410 (N_2410,N_391,N_780);
or U2411 (N_2411,N_1571,N_241);
or U2412 (N_2412,N_1071,N_1251);
and U2413 (N_2413,N_296,N_597);
xor U2414 (N_2414,N_1058,N_1335);
and U2415 (N_2415,N_359,N_1151);
nand U2416 (N_2416,N_121,N_270);
nand U2417 (N_2417,N_1705,N_144);
xor U2418 (N_2418,N_1157,N_516);
and U2419 (N_2419,N_85,N_824);
and U2420 (N_2420,N_918,N_1533);
nand U2421 (N_2421,N_1909,N_392);
nand U2422 (N_2422,N_1502,N_1240);
xnor U2423 (N_2423,N_808,N_482);
or U2424 (N_2424,N_1192,N_1215);
nor U2425 (N_2425,N_1262,N_2);
nor U2426 (N_2426,N_172,N_483);
and U2427 (N_2427,N_1560,N_621);
nand U2428 (N_2428,N_420,N_1127);
nor U2429 (N_2429,N_842,N_499);
or U2430 (N_2430,N_1015,N_1693);
nor U2431 (N_2431,N_1617,N_1441);
xnor U2432 (N_2432,N_198,N_434);
or U2433 (N_2433,N_682,N_1082);
xor U2434 (N_2434,N_1062,N_449);
and U2435 (N_2435,N_1043,N_722);
and U2436 (N_2436,N_1412,N_317);
nand U2437 (N_2437,N_1926,N_1623);
nand U2438 (N_2438,N_855,N_1033);
xnor U2439 (N_2439,N_1088,N_1189);
nor U2440 (N_2440,N_1399,N_63);
nand U2441 (N_2441,N_1791,N_29);
nand U2442 (N_2442,N_1967,N_981);
or U2443 (N_2443,N_388,N_977);
and U2444 (N_2444,N_374,N_1280);
nand U2445 (N_2445,N_947,N_90);
xnor U2446 (N_2446,N_1457,N_224);
xor U2447 (N_2447,N_1408,N_1233);
xor U2448 (N_2448,N_602,N_505);
and U2449 (N_2449,N_535,N_232);
and U2450 (N_2450,N_1570,N_1744);
or U2451 (N_2451,N_934,N_1367);
or U2452 (N_2452,N_26,N_347);
nand U2453 (N_2453,N_33,N_1528);
and U2454 (N_2454,N_729,N_1407);
or U2455 (N_2455,N_276,N_719);
and U2456 (N_2456,N_1669,N_1779);
xnor U2457 (N_2457,N_874,N_1276);
and U2458 (N_2458,N_1229,N_819);
nor U2459 (N_2459,N_1789,N_1449);
nor U2460 (N_2460,N_1345,N_1766);
or U2461 (N_2461,N_448,N_361);
xor U2462 (N_2462,N_1072,N_1912);
xor U2463 (N_2463,N_171,N_1012);
or U2464 (N_2464,N_1115,N_1063);
and U2465 (N_2465,N_1891,N_441);
nor U2466 (N_2466,N_72,N_1201);
or U2467 (N_2467,N_1471,N_1351);
and U2468 (N_2468,N_8,N_354);
xnor U2469 (N_2469,N_832,N_972);
or U2470 (N_2470,N_1723,N_1576);
nand U2471 (N_2471,N_636,N_1861);
xnor U2472 (N_2472,N_577,N_1619);
and U2473 (N_2473,N_247,N_1921);
xnor U2474 (N_2474,N_376,N_1438);
nor U2475 (N_2475,N_385,N_1892);
nor U2476 (N_2476,N_1986,N_1706);
or U2477 (N_2477,N_97,N_15);
xor U2478 (N_2478,N_1055,N_1166);
or U2479 (N_2479,N_524,N_1666);
xor U2480 (N_2480,N_894,N_1629);
nand U2481 (N_2481,N_1547,N_1819);
nand U2482 (N_2482,N_136,N_287);
nor U2483 (N_2483,N_411,N_329);
and U2484 (N_2484,N_527,N_552);
nand U2485 (N_2485,N_1329,N_666);
nand U2486 (N_2486,N_1237,N_1392);
and U2487 (N_2487,N_1142,N_891);
xnor U2488 (N_2488,N_1469,N_1332);
or U2489 (N_2489,N_555,N_47);
nand U2490 (N_2490,N_1786,N_1665);
or U2491 (N_2491,N_1136,N_330);
nor U2492 (N_2492,N_196,N_1760);
xor U2493 (N_2493,N_452,N_583);
nand U2494 (N_2494,N_1070,N_1328);
and U2495 (N_2495,N_1568,N_163);
and U2496 (N_2496,N_985,N_1548);
and U2497 (N_2497,N_966,N_408);
and U2498 (N_2498,N_1304,N_141);
xnor U2499 (N_2499,N_1281,N_1417);
nand U2500 (N_2500,N_1467,N_622);
nor U2501 (N_2501,N_1389,N_1671);
xnor U2502 (N_2502,N_540,N_353);
xnor U2503 (N_2503,N_1624,N_738);
nor U2504 (N_2504,N_1355,N_1156);
nand U2505 (N_2505,N_1194,N_1595);
and U2506 (N_2506,N_159,N_1733);
nor U2507 (N_2507,N_559,N_1898);
xnor U2508 (N_2508,N_220,N_472);
and U2509 (N_2509,N_274,N_1165);
and U2510 (N_2510,N_124,N_810);
xnor U2511 (N_2511,N_1060,N_1944);
xor U2512 (N_2512,N_1031,N_187);
and U2513 (N_2513,N_289,N_280);
nand U2514 (N_2514,N_925,N_469);
nor U2515 (N_2515,N_600,N_1443);
xor U2516 (N_2516,N_830,N_1026);
nor U2517 (N_2517,N_362,N_299);
or U2518 (N_2518,N_913,N_418);
or U2519 (N_2519,N_479,N_919);
and U2520 (N_2520,N_784,N_1419);
or U2521 (N_2521,N_127,N_1679);
nand U2522 (N_2522,N_50,N_541);
or U2523 (N_2523,N_553,N_477);
and U2524 (N_2524,N_1782,N_953);
xor U2525 (N_2525,N_1591,N_129);
and U2526 (N_2526,N_210,N_777);
nand U2527 (N_2527,N_1238,N_574);
and U2528 (N_2528,N_1084,N_523);
and U2529 (N_2529,N_901,N_542);
or U2530 (N_2530,N_1294,N_1296);
and U2531 (N_2531,N_826,N_759);
or U2532 (N_2532,N_189,N_648);
nor U2533 (N_2533,N_491,N_324);
or U2534 (N_2534,N_1317,N_633);
xnor U2535 (N_2535,N_126,N_1206);
and U2536 (N_2536,N_532,N_1410);
or U2537 (N_2537,N_1524,N_1834);
and U2538 (N_2538,N_1161,N_1922);
xnor U2539 (N_2539,N_41,N_1284);
or U2540 (N_2540,N_405,N_1692);
nand U2541 (N_2541,N_658,N_1330);
nor U2542 (N_2542,N_1759,N_958);
or U2543 (N_2543,N_251,N_1244);
or U2544 (N_2544,N_557,N_1);
nand U2545 (N_2545,N_1558,N_971);
or U2546 (N_2546,N_896,N_1882);
nand U2547 (N_2547,N_507,N_1818);
xnor U2548 (N_2548,N_145,N_226);
xnor U2549 (N_2549,N_1505,N_1650);
or U2550 (N_2550,N_892,N_1267);
or U2551 (N_2551,N_458,N_510);
nor U2552 (N_2552,N_994,N_92);
and U2553 (N_2553,N_1075,N_1182);
nor U2554 (N_2554,N_1844,N_1878);
nand U2555 (N_2555,N_1869,N_1310);
or U2556 (N_2556,N_1601,N_1987);
and U2557 (N_2557,N_1213,N_1363);
and U2558 (N_2558,N_1040,N_639);
xnor U2559 (N_2559,N_1334,N_259);
xor U2560 (N_2560,N_1599,N_1856);
or U2561 (N_2561,N_1388,N_1220);
nor U2562 (N_2562,N_66,N_1339);
nor U2563 (N_2563,N_30,N_135);
nand U2564 (N_2564,N_1625,N_879);
or U2565 (N_2565,N_1274,N_873);
and U2566 (N_2566,N_531,N_298);
or U2567 (N_2567,N_1170,N_1178);
nor U2568 (N_2568,N_1561,N_372);
and U2569 (N_2569,N_710,N_1044);
and U2570 (N_2570,N_1023,N_1087);
nor U2571 (N_2571,N_1574,N_438);
and U2572 (N_2572,N_828,N_927);
and U2573 (N_2573,N_1521,N_1086);
xnor U2574 (N_2574,N_1538,N_1475);
nor U2575 (N_2575,N_468,N_1042);
nand U2576 (N_2576,N_1434,N_1589);
nand U2577 (N_2577,N_1191,N_1907);
xnor U2578 (N_2578,N_769,N_58);
xor U2579 (N_2579,N_419,N_1037);
nand U2580 (N_2580,N_1452,N_1059);
nand U2581 (N_2581,N_608,N_343);
and U2582 (N_2582,N_445,N_1459);
or U2583 (N_2583,N_502,N_1064);
nand U2584 (N_2584,N_1543,N_1106);
nand U2585 (N_2585,N_318,N_1371);
nor U2586 (N_2586,N_1185,N_1872);
nor U2587 (N_2587,N_1004,N_336);
or U2588 (N_2588,N_973,N_1083);
or U2589 (N_2589,N_1902,N_1928);
and U2590 (N_2590,N_1143,N_1293);
and U2591 (N_2591,N_65,N_789);
or U2592 (N_2592,N_1702,N_1796);
and U2593 (N_2593,N_1342,N_798);
nand U2594 (N_2594,N_1184,N_1682);
nand U2595 (N_2595,N_951,N_1527);
nor U2596 (N_2596,N_923,N_103);
or U2597 (N_2597,N_1664,N_1916);
or U2598 (N_2598,N_43,N_1522);
nor U2599 (N_2599,N_800,N_1684);
nand U2600 (N_2600,N_922,N_1867);
and U2601 (N_2601,N_786,N_1121);
nor U2602 (N_2602,N_1025,N_67);
xnor U2603 (N_2603,N_603,N_1894);
and U2604 (N_2604,N_820,N_208);
and U2605 (N_2605,N_625,N_1946);
nand U2606 (N_2606,N_1048,N_999);
nor U2607 (N_2607,N_1659,N_1315);
xor U2608 (N_2608,N_1839,N_1211);
nor U2609 (N_2609,N_1960,N_173);
or U2610 (N_2610,N_1235,N_1772);
and U2611 (N_2611,N_869,N_585);
nor U2612 (N_2612,N_921,N_1204);
or U2613 (N_2613,N_390,N_623);
or U2614 (N_2614,N_1632,N_1849);
or U2615 (N_2615,N_44,N_1716);
nor U2616 (N_2616,N_1969,N_1131);
or U2617 (N_2617,N_566,N_406);
and U2618 (N_2618,N_838,N_199);
or U2619 (N_2619,N_1727,N_264);
or U2620 (N_2620,N_1154,N_315);
and U2621 (N_2621,N_1301,N_1175);
nor U2622 (N_2622,N_384,N_1255);
nand U2623 (N_2623,N_560,N_1202);
nand U2624 (N_2624,N_183,N_442);
nor U2625 (N_2625,N_1278,N_1788);
or U2626 (N_2626,N_1919,N_1626);
nor U2627 (N_2627,N_1100,N_1649);
or U2628 (N_2628,N_1431,N_935);
nor U2629 (N_2629,N_640,N_1715);
nor U2630 (N_2630,N_319,N_1739);
and U2631 (N_2631,N_1537,N_846);
nor U2632 (N_2632,N_825,N_1971);
nor U2633 (N_2633,N_525,N_386);
or U2634 (N_2634,N_883,N_1511);
nor U2635 (N_2635,N_223,N_1563);
nor U2636 (N_2636,N_739,N_1645);
nand U2637 (N_2637,N_421,N_1096);
or U2638 (N_2638,N_1442,N_907);
nand U2639 (N_2639,N_1496,N_1864);
nor U2640 (N_2640,N_752,N_1817);
and U2641 (N_2641,N_402,N_545);
or U2642 (N_2642,N_1598,N_1503);
and U2643 (N_2643,N_1536,N_1910);
nand U2644 (N_2644,N_94,N_1564);
xnor U2645 (N_2645,N_1153,N_671);
nor U2646 (N_2646,N_1606,N_713);
and U2647 (N_2647,N_1027,N_1953);
or U2648 (N_2648,N_277,N_1724);
xnor U2649 (N_2649,N_1145,N_1394);
nand U2650 (N_2650,N_1414,N_1383);
and U2651 (N_2651,N_1167,N_862);
xor U2652 (N_2652,N_255,N_1424);
or U2653 (N_2653,N_992,N_902);
xnor U2654 (N_2654,N_439,N_1972);
xnor U2655 (N_2655,N_1719,N_822);
nand U2656 (N_2656,N_544,N_1338);
nor U2657 (N_2657,N_478,N_1687);
nand U2658 (N_2658,N_1586,N_1357);
nor U2659 (N_2659,N_582,N_133);
nor U2660 (N_2660,N_53,N_131);
nor U2661 (N_2661,N_1635,N_591);
or U2662 (N_2662,N_480,N_1935);
xor U2663 (N_2663,N_1754,N_1551);
xor U2664 (N_2664,N_979,N_596);
xnor U2665 (N_2665,N_723,N_1552);
nor U2666 (N_2666,N_380,N_708);
nor U2667 (N_2667,N_1994,N_1036);
nor U2668 (N_2668,N_218,N_957);
xor U2669 (N_2669,N_1757,N_1081);
and U2670 (N_2670,N_1066,N_424);
nand U2671 (N_2671,N_123,N_920);
xnor U2672 (N_2672,N_1567,N_1212);
or U2673 (N_2673,N_31,N_569);
nand U2674 (N_2674,N_1348,N_481);
nand U2675 (N_2675,N_1344,N_791);
xnor U2676 (N_2676,N_262,N_1200);
nor U2677 (N_2677,N_1114,N_701);
nand U2678 (N_2678,N_1405,N_1325);
and U2679 (N_2679,N_517,N_1900);
nand U2680 (N_2680,N_948,N_1478);
nand U2681 (N_2681,N_1711,N_1003);
and U2682 (N_2682,N_1846,N_1722);
and U2683 (N_2683,N_99,N_12);
and U2684 (N_2684,N_1382,N_231);
nor U2685 (N_2685,N_1512,N_1681);
or U2686 (N_2686,N_551,N_1306);
nand U2687 (N_2687,N_1513,N_1163);
or U2688 (N_2688,N_242,N_146);
nand U2689 (N_2689,N_1811,N_1482);
nand U2690 (N_2690,N_1376,N_306);
xor U2691 (N_2691,N_245,N_863);
nor U2692 (N_2692,N_801,N_912);
nand U2693 (N_2693,N_1395,N_288);
nor U2694 (N_2694,N_370,N_1542);
nor U2695 (N_2695,N_537,N_584);
nand U2696 (N_2696,N_93,N_16);
or U2697 (N_2697,N_1866,N_609);
and U2698 (N_2698,N_414,N_485);
or U2699 (N_2699,N_1259,N_213);
xnor U2700 (N_2700,N_794,N_463);
or U2701 (N_2701,N_1600,N_24);
or U2702 (N_2702,N_1809,N_1477);
nor U2703 (N_2703,N_1446,N_630);
nor U2704 (N_2704,N_730,N_168);
or U2705 (N_2705,N_1205,N_703);
nand U2706 (N_2706,N_180,N_430);
or U2707 (N_2707,N_651,N_1029);
and U2708 (N_2708,N_607,N_410);
or U2709 (N_2709,N_1309,N_425);
nor U2710 (N_2710,N_1845,N_929);
xor U2711 (N_2711,N_1493,N_1952);
nor U2712 (N_2712,N_437,N_1518);
and U2713 (N_2713,N_1112,N_294);
nor U2714 (N_2714,N_440,N_978);
nand U2715 (N_2715,N_1400,N_563);
nor U2716 (N_2716,N_707,N_184);
nor U2717 (N_2717,N_1762,N_629);
xnor U2718 (N_2718,N_495,N_100);
nand U2719 (N_2719,N_117,N_1607);
or U2720 (N_2720,N_39,N_905);
or U2721 (N_2721,N_1655,N_27);
or U2722 (N_2722,N_1272,N_860);
nor U2723 (N_2723,N_1198,N_1848);
or U2724 (N_2724,N_1266,N_1427);
nand U2725 (N_2725,N_844,N_941);
nand U2726 (N_2726,N_976,N_1470);
or U2727 (N_2727,N_1230,N_1541);
xnor U2728 (N_2728,N_95,N_700);
and U2729 (N_2729,N_1174,N_54);
nand U2730 (N_2730,N_611,N_13);
or U2731 (N_2731,N_1901,N_961);
nor U2732 (N_2732,N_1014,N_835);
or U2733 (N_2733,N_78,N_1525);
nand U2734 (N_2734,N_877,N_269);
xor U2735 (N_2735,N_1375,N_1307);
and U2736 (N_2736,N_360,N_69);
xor U2737 (N_2737,N_1539,N_1663);
or U2738 (N_2738,N_490,N_744);
and U2739 (N_2739,N_162,N_102);
or U2740 (N_2740,N_1647,N_1923);
or U2741 (N_2741,N_1243,N_313);
nor U2742 (N_2742,N_71,N_930);
xnor U2743 (N_2743,N_84,N_239);
nand U2744 (N_2744,N_1193,N_1097);
xor U2745 (N_2745,N_1862,N_1413);
xnor U2746 (N_2746,N_1814,N_1466);
nor U2747 (N_2747,N_87,N_1642);
nor U2748 (N_2748,N_1094,N_735);
xor U2749 (N_2749,N_107,N_1125);
or U2750 (N_2750,N_1321,N_243);
nand U2751 (N_2751,N_409,N_1868);
nor U2752 (N_2752,N_526,N_1850);
nand U2753 (N_2753,N_1288,N_519);
nor U2754 (N_2754,N_688,N_1585);
nor U2755 (N_2755,N_821,N_357);
nand U2756 (N_2756,N_1871,N_307);
and U2757 (N_2757,N_466,N_496);
xor U2758 (N_2758,N_1222,N_938);
xnor U2759 (N_2759,N_1091,N_718);
or U2760 (N_2760,N_520,N_1594);
xnor U2761 (N_2761,N_849,N_1683);
nand U2762 (N_2762,N_1289,N_693);
or U2763 (N_2763,N_1343,N_1997);
and U2764 (N_2764,N_1996,N_1492);
and U2765 (N_2765,N_1708,N_257);
xor U2766 (N_2766,N_1964,N_772);
xnor U2767 (N_2767,N_1011,N_1090);
or U2768 (N_2768,N_428,N_642);
nor U2769 (N_2769,N_1767,N_86);
and U2770 (N_2770,N_667,N_273);
nand U2771 (N_2771,N_1187,N_1895);
nand U2772 (N_2772,N_1523,N_1393);
and U2773 (N_2773,N_19,N_75);
and U2774 (N_2774,N_256,N_467);
or U2775 (N_2775,N_310,N_1402);
nor U2776 (N_2776,N_334,N_1569);
xor U2777 (N_2777,N_848,N_1691);
or U2778 (N_2778,N_37,N_890);
and U2779 (N_2779,N_1929,N_217);
nand U2780 (N_2780,N_1605,N_1592);
or U2781 (N_2781,N_1925,N_1820);
and U2782 (N_2782,N_965,N_933);
and U2783 (N_2783,N_176,N_1970);
xnor U2784 (N_2784,N_620,N_1159);
nor U2785 (N_2785,N_1825,N_166);
nor U2786 (N_2786,N_161,N_1366);
nor U2787 (N_2787,N_861,N_783);
xnor U2788 (N_2788,N_691,N_1917);
or U2789 (N_2789,N_1226,N_1956);
and U2790 (N_2790,N_654,N_1932);
nand U2791 (N_2791,N_503,N_937);
or U2792 (N_2792,N_1555,N_1768);
nand U2793 (N_2793,N_1730,N_613);
nand U2794 (N_2794,N_1644,N_1685);
xnor U2795 (N_2795,N_1331,N_1798);
and U2796 (N_2796,N_647,N_645);
and U2797 (N_2797,N_1068,N_851);
nand U2798 (N_2798,N_130,N_1546);
nor U2799 (N_2799,N_285,N_1965);
or U2800 (N_2800,N_1506,N_790);
or U2801 (N_2801,N_1349,N_1323);
and U2802 (N_2802,N_669,N_1476);
nand U2803 (N_2803,N_500,N_1680);
and U2804 (N_2804,N_799,N_493);
nand U2805 (N_2805,N_60,N_1146);
nand U2806 (N_2806,N_1621,N_1697);
and U2807 (N_2807,N_580,N_1186);
xnor U2808 (N_2808,N_1802,N_387);
nand U2809 (N_2809,N_1373,N_831);
or U2810 (N_2810,N_1851,N_1260);
and U2811 (N_2811,N_1188,N_781);
nand U2812 (N_2812,N_928,N_1736);
and U2813 (N_2813,N_1437,N_1813);
nor U2814 (N_2814,N_615,N_1480);
and U2815 (N_2815,N_712,N_614);
nor U2816 (N_2816,N_1602,N_1500);
and U2817 (N_2817,N_1980,N_521);
xnor U2818 (N_2818,N_331,N_399);
xor U2819 (N_2819,N_1947,N_23);
nand U2820 (N_2820,N_201,N_1822);
xor U2821 (N_2821,N_564,N_1999);
nor U2822 (N_2822,N_454,N_1435);
and U2823 (N_2823,N_1129,N_271);
nor U2824 (N_2824,N_834,N_895);
nor U2825 (N_2825,N_1628,N_1126);
and U2826 (N_2826,N_774,N_716);
and U2827 (N_2827,N_1360,N_1319);
or U2828 (N_2828,N_1484,N_903);
or U2829 (N_2829,N_889,N_1615);
or U2830 (N_2830,N_1717,N_263);
and U2831 (N_2831,N_1828,N_1853);
nand U2832 (N_2832,N_1580,N_1673);
xor U2833 (N_2833,N_917,N_328);
and U2834 (N_2834,N_1810,N_634);
xor U2835 (N_2835,N_383,N_1361);
nor U2836 (N_2836,N_549,N_815);
nand U2837 (N_2837,N_1812,N_1387);
or U2838 (N_2838,N_1660,N_175);
nand U2839 (N_2839,N_1638,N_1507);
and U2840 (N_2840,N_1636,N_194);
and U2841 (N_2841,N_366,N_81);
or U2842 (N_2842,N_417,N_1369);
xnor U2843 (N_2843,N_1637,N_1753);
nor U2844 (N_2844,N_1957,N_190);
nand U2845 (N_2845,N_1173,N_1897);
nor U2846 (N_2846,N_512,N_1119);
and U2847 (N_2847,N_1098,N_586);
xnor U2848 (N_2848,N_337,N_1245);
and U2849 (N_2849,N_142,N_788);
or U2850 (N_2850,N_1137,N_284);
nor U2851 (N_2851,N_309,N_1275);
and U2852 (N_2852,N_1890,N_423);
nand U2853 (N_2853,N_755,N_875);
nand U2854 (N_2854,N_812,N_1311);
nor U2855 (N_2855,N_492,N_1190);
nor U2856 (N_2856,N_568,N_1113);
and U2857 (N_2857,N_290,N_1359);
and U2858 (N_2858,N_1933,N_216);
nand U2859 (N_2859,N_743,N_661);
or U2860 (N_2860,N_326,N_1672);
or U2861 (N_2861,N_234,N_872);
nor U2862 (N_2862,N_1658,N_179);
or U2863 (N_2863,N_847,N_1069);
nor U2864 (N_2864,N_504,N_1358);
or U2865 (N_2865,N_333,N_1651);
nor U2866 (N_2866,N_356,N_1945);
or U2867 (N_2867,N_110,N_191);
nor U2868 (N_2868,N_605,N_1291);
nor U2869 (N_2869,N_1830,N_760);
xnor U2870 (N_2870,N_346,N_447);
nand U2871 (N_2871,N_610,N_461);
and U2872 (N_2872,N_1132,N_1495);
and U2873 (N_2873,N_1302,N_453);
or U2874 (N_2874,N_186,N_1535);
xnor U2875 (N_2875,N_1020,N_592);
nor U2876 (N_2876,N_268,N_363);
nand U2877 (N_2877,N_498,N_395);
and U2878 (N_2878,N_1783,N_1124);
nor U2879 (N_2879,N_381,N_1270);
nor U2880 (N_2880,N_867,N_1488);
or U2881 (N_2881,N_1836,N_1298);
and U2882 (N_2882,N_1983,N_991);
or U2883 (N_2883,N_1384,N_400);
xor U2884 (N_2884,N_1771,N_734);
nand U2885 (N_2885,N_355,N_14);
or U2886 (N_2886,N_1936,N_886);
xor U2887 (N_2887,N_1464,N_46);
nand U2888 (N_2888,N_1000,N_1385);
or U2889 (N_2889,N_590,N_1401);
nand U2890 (N_2890,N_1974,N_109);
nand U2891 (N_2891,N_543,N_1741);
nor U2892 (N_2892,N_225,N_215);
and U2893 (N_2893,N_1942,N_1841);
nor U2894 (N_2894,N_836,N_1109);
nor U2895 (N_2895,N_1051,N_1073);
nor U2896 (N_2896,N_207,N_1893);
or U2897 (N_2897,N_1279,N_702);
nor U2898 (N_2898,N_236,N_1354);
or U2899 (N_2899,N_1498,N_717);
or U2900 (N_2900,N_1045,N_650);
nand U2901 (N_2901,N_1734,N_1403);
nand U2902 (N_2902,N_1039,N_1013);
and U2903 (N_2903,N_1008,N_340);
xor U2904 (N_2904,N_1210,N_1256);
xnor U2905 (N_2905,N_1241,N_884);
xor U2906 (N_2906,N_612,N_143);
or U2907 (N_2907,N_575,N_536);
or U2908 (N_2908,N_1415,N_74);
nand U2909 (N_2909,N_573,N_373);
or U2910 (N_2910,N_200,N_98);
nand U2911 (N_2911,N_711,N_369);
xnor U2912 (N_2912,N_364,N_853);
nand U2913 (N_2913,N_1641,N_595);
nand U2914 (N_2914,N_1463,N_96);
or U2915 (N_2915,N_249,N_628);
xnor U2916 (N_2916,N_983,N_988);
and U2917 (N_2917,N_765,N_1236);
and U2918 (N_2918,N_214,N_9);
and U2919 (N_2919,N_1404,N_1005);
nor U2920 (N_2920,N_1249,N_955);
and U2921 (N_2921,N_997,N_34);
or U2922 (N_2922,N_1992,N_1731);
nor U2923 (N_2923,N_829,N_1425);
xor U2924 (N_2924,N_158,N_660);
or U2925 (N_2925,N_1105,N_1520);
nand U2926 (N_2926,N_1604,N_986);
nand U2927 (N_2927,N_1374,N_1120);
and U2928 (N_2928,N_1002,N_76);
nand U2929 (N_2929,N_1899,N_742);
nand U2930 (N_2930,N_984,N_371);
and U2931 (N_2931,N_599,N_1835);
nor U2932 (N_2932,N_1074,N_323);
and U2933 (N_2933,N_782,N_1433);
and U2934 (N_2934,N_1445,N_1939);
nand U2935 (N_2935,N_160,N_32);
nor U2936 (N_2936,N_1250,N_137);
nand U2937 (N_2937,N_40,N_993);
and U2938 (N_2938,N_982,N_764);
nand U2939 (N_2939,N_378,N_1838);
nor U2940 (N_2940,N_293,N_125);
or U2941 (N_2941,N_814,N_1610);
xor U2942 (N_2942,N_1396,N_1264);
xor U2943 (N_2943,N_533,N_1954);
and U2944 (N_2944,N_805,N_486);
or U2945 (N_2945,N_1720,N_1756);
xnor U2946 (N_2946,N_1324,N_197);
nor U2947 (N_2947,N_1032,N_350);
nor U2948 (N_2948,N_1472,N_766);
nor U2949 (N_2949,N_579,N_619);
or U2950 (N_2950,N_153,N_1887);
nor U2951 (N_2951,N_1657,N_327);
and U2952 (N_2952,N_192,N_1257);
nand U2953 (N_2953,N_567,N_881);
and U2954 (N_2954,N_758,N_1884);
nand U2955 (N_2955,N_1961,N_627);
nor U2956 (N_2956,N_1984,N_1735);
xor U2957 (N_2957,N_865,N_1447);
or U2958 (N_2958,N_1976,N_70);
nor U2959 (N_2959,N_662,N_1397);
xor U2960 (N_2960,N_426,N_804);
and U2961 (N_2961,N_368,N_1738);
or U2962 (N_2962,N_1128,N_967);
nor U2963 (N_2963,N_1271,N_1748);
nand U2964 (N_2964,N_79,N_1219);
nor U2965 (N_2965,N_841,N_1350);
xor U2966 (N_2966,N_1092,N_910);
nand U2967 (N_2967,N_115,N_1765);
or U2968 (N_2968,N_1699,N_254);
and U2969 (N_2969,N_1577,N_672);
nor U2970 (N_2970,N_670,N_88);
nand U2971 (N_2971,N_1876,N_1540);
xor U2972 (N_2972,N_393,N_432);
nand U2973 (N_2973,N_1077,N_156);
nor U2974 (N_2974,N_487,N_1377);
or U2975 (N_2975,N_1737,N_1823);
nand U2976 (N_2976,N_675,N_1775);
nand U2977 (N_2977,N_1859,N_1223);
or U2978 (N_2978,N_704,N_963);
or U2979 (N_2979,N_989,N_806);
xor U2980 (N_2980,N_1648,N_1749);
xor U2981 (N_2981,N_489,N_915);
nor U2982 (N_2982,N_1751,N_1978);
or U2983 (N_2983,N_1517,N_1877);
nand U2984 (N_2984,N_1698,N_1282);
nor U2985 (N_2985,N_1858,N_793);
and U2986 (N_2986,N_398,N_632);
nand U2987 (N_2987,N_282,N_1181);
or U2988 (N_2988,N_36,N_1277);
or U2989 (N_2989,N_1183,N_1597);
and U2990 (N_2990,N_305,N_1168);
nor U2991 (N_2991,N_571,N_1807);
or U2992 (N_2992,N_696,N_1911);
nor U2993 (N_2993,N_367,N_714);
or U2994 (N_2994,N_59,N_1526);
and U2995 (N_2995,N_833,N_1661);
nor U2996 (N_2996,N_455,N_1634);
nand U2997 (N_2997,N_1770,N_705);
xor U2998 (N_2998,N_1519,N_1803);
nor U2999 (N_2999,N_1079,N_1712);
nor U3000 (N_3000,N_1955,N_380);
nand U3001 (N_3001,N_845,N_20);
or U3002 (N_3002,N_708,N_1485);
and U3003 (N_3003,N_1368,N_1998);
and U3004 (N_3004,N_1603,N_1857);
nand U3005 (N_3005,N_1282,N_1995);
and U3006 (N_3006,N_364,N_1210);
nor U3007 (N_3007,N_1769,N_1481);
or U3008 (N_3008,N_1915,N_106);
nor U3009 (N_3009,N_1676,N_370);
and U3010 (N_3010,N_586,N_180);
nor U3011 (N_3011,N_345,N_225);
nand U3012 (N_3012,N_303,N_500);
and U3013 (N_3013,N_516,N_617);
and U3014 (N_3014,N_1475,N_1421);
and U3015 (N_3015,N_1605,N_1617);
xor U3016 (N_3016,N_1773,N_375);
and U3017 (N_3017,N_1985,N_679);
or U3018 (N_3018,N_566,N_203);
nand U3019 (N_3019,N_125,N_405);
nor U3020 (N_3020,N_1965,N_386);
or U3021 (N_3021,N_502,N_159);
xor U3022 (N_3022,N_1447,N_1316);
nor U3023 (N_3023,N_813,N_240);
or U3024 (N_3024,N_1317,N_1807);
nand U3025 (N_3025,N_1401,N_1338);
and U3026 (N_3026,N_529,N_758);
or U3027 (N_3027,N_899,N_1429);
nor U3028 (N_3028,N_1391,N_1132);
xnor U3029 (N_3029,N_398,N_822);
nor U3030 (N_3030,N_418,N_1070);
nand U3031 (N_3031,N_466,N_174);
xnor U3032 (N_3032,N_1471,N_1282);
nand U3033 (N_3033,N_1294,N_37);
nand U3034 (N_3034,N_1212,N_165);
nor U3035 (N_3035,N_1479,N_1751);
nand U3036 (N_3036,N_1091,N_228);
nand U3037 (N_3037,N_1952,N_1405);
and U3038 (N_3038,N_662,N_823);
nand U3039 (N_3039,N_563,N_510);
or U3040 (N_3040,N_1408,N_1409);
nand U3041 (N_3041,N_1135,N_452);
and U3042 (N_3042,N_865,N_672);
nor U3043 (N_3043,N_601,N_367);
and U3044 (N_3044,N_1614,N_1651);
xnor U3045 (N_3045,N_873,N_16);
nor U3046 (N_3046,N_122,N_1708);
nand U3047 (N_3047,N_80,N_266);
xor U3048 (N_3048,N_1380,N_227);
or U3049 (N_3049,N_1627,N_932);
and U3050 (N_3050,N_766,N_1797);
and U3051 (N_3051,N_226,N_1206);
xnor U3052 (N_3052,N_1320,N_72);
nor U3053 (N_3053,N_1247,N_289);
and U3054 (N_3054,N_1535,N_1115);
nor U3055 (N_3055,N_1891,N_245);
nand U3056 (N_3056,N_243,N_333);
and U3057 (N_3057,N_263,N_1244);
nand U3058 (N_3058,N_1982,N_113);
xor U3059 (N_3059,N_1103,N_985);
nor U3060 (N_3060,N_254,N_410);
nor U3061 (N_3061,N_1367,N_1373);
or U3062 (N_3062,N_1778,N_1418);
nand U3063 (N_3063,N_972,N_1460);
xor U3064 (N_3064,N_42,N_1515);
nand U3065 (N_3065,N_773,N_1041);
nand U3066 (N_3066,N_1972,N_1076);
nand U3067 (N_3067,N_1951,N_529);
or U3068 (N_3068,N_1452,N_100);
nand U3069 (N_3069,N_1704,N_1045);
and U3070 (N_3070,N_722,N_788);
xor U3071 (N_3071,N_91,N_1445);
nand U3072 (N_3072,N_1128,N_1400);
xnor U3073 (N_3073,N_636,N_1652);
or U3074 (N_3074,N_821,N_199);
and U3075 (N_3075,N_1989,N_856);
or U3076 (N_3076,N_135,N_1926);
nand U3077 (N_3077,N_1762,N_1898);
or U3078 (N_3078,N_718,N_1843);
xor U3079 (N_3079,N_987,N_252);
xnor U3080 (N_3080,N_54,N_1673);
nand U3081 (N_3081,N_1510,N_1799);
xor U3082 (N_3082,N_1480,N_158);
or U3083 (N_3083,N_1891,N_1017);
and U3084 (N_3084,N_1137,N_1058);
xor U3085 (N_3085,N_1894,N_1887);
nor U3086 (N_3086,N_707,N_992);
nand U3087 (N_3087,N_1994,N_796);
and U3088 (N_3088,N_1571,N_509);
nor U3089 (N_3089,N_447,N_172);
nor U3090 (N_3090,N_812,N_1567);
xor U3091 (N_3091,N_1859,N_1136);
nand U3092 (N_3092,N_56,N_1791);
nor U3093 (N_3093,N_1313,N_1236);
xnor U3094 (N_3094,N_437,N_137);
nor U3095 (N_3095,N_1906,N_143);
nand U3096 (N_3096,N_558,N_551);
and U3097 (N_3097,N_1210,N_1243);
nor U3098 (N_3098,N_439,N_1661);
and U3099 (N_3099,N_1481,N_1777);
nor U3100 (N_3100,N_382,N_1295);
xor U3101 (N_3101,N_412,N_539);
and U3102 (N_3102,N_1081,N_1436);
nand U3103 (N_3103,N_72,N_1167);
and U3104 (N_3104,N_1486,N_453);
xnor U3105 (N_3105,N_61,N_713);
xor U3106 (N_3106,N_1330,N_297);
or U3107 (N_3107,N_487,N_1343);
and U3108 (N_3108,N_670,N_976);
nor U3109 (N_3109,N_148,N_1749);
xnor U3110 (N_3110,N_844,N_1287);
nand U3111 (N_3111,N_1715,N_1255);
or U3112 (N_3112,N_600,N_688);
or U3113 (N_3113,N_1048,N_809);
nor U3114 (N_3114,N_1479,N_539);
nand U3115 (N_3115,N_397,N_1562);
xor U3116 (N_3116,N_252,N_1871);
xor U3117 (N_3117,N_1178,N_1619);
nand U3118 (N_3118,N_1058,N_799);
and U3119 (N_3119,N_1392,N_1532);
and U3120 (N_3120,N_1257,N_1116);
or U3121 (N_3121,N_1450,N_1623);
xor U3122 (N_3122,N_1678,N_1538);
or U3123 (N_3123,N_677,N_1352);
nand U3124 (N_3124,N_142,N_335);
xor U3125 (N_3125,N_1697,N_348);
nand U3126 (N_3126,N_41,N_1966);
nand U3127 (N_3127,N_533,N_1584);
nor U3128 (N_3128,N_682,N_940);
nand U3129 (N_3129,N_1542,N_1443);
nor U3130 (N_3130,N_1786,N_1627);
and U3131 (N_3131,N_1869,N_385);
and U3132 (N_3132,N_1657,N_559);
nor U3133 (N_3133,N_811,N_1363);
nor U3134 (N_3134,N_919,N_545);
nor U3135 (N_3135,N_1122,N_95);
and U3136 (N_3136,N_404,N_224);
nand U3137 (N_3137,N_945,N_260);
xnor U3138 (N_3138,N_683,N_759);
and U3139 (N_3139,N_916,N_597);
and U3140 (N_3140,N_1562,N_506);
or U3141 (N_3141,N_1381,N_1086);
and U3142 (N_3142,N_1341,N_428);
or U3143 (N_3143,N_1007,N_181);
nor U3144 (N_3144,N_1360,N_1815);
nand U3145 (N_3145,N_1082,N_416);
and U3146 (N_3146,N_582,N_810);
or U3147 (N_3147,N_943,N_223);
nand U3148 (N_3148,N_1473,N_315);
or U3149 (N_3149,N_1691,N_1651);
and U3150 (N_3150,N_1929,N_490);
nand U3151 (N_3151,N_876,N_1490);
and U3152 (N_3152,N_110,N_218);
nand U3153 (N_3153,N_1305,N_302);
and U3154 (N_3154,N_1554,N_381);
and U3155 (N_3155,N_1229,N_1500);
xor U3156 (N_3156,N_1845,N_537);
nor U3157 (N_3157,N_1769,N_1243);
nand U3158 (N_3158,N_1285,N_202);
nor U3159 (N_3159,N_1376,N_398);
nand U3160 (N_3160,N_1857,N_599);
nor U3161 (N_3161,N_617,N_216);
or U3162 (N_3162,N_1543,N_1943);
nor U3163 (N_3163,N_293,N_1550);
and U3164 (N_3164,N_1486,N_1362);
and U3165 (N_3165,N_761,N_101);
nand U3166 (N_3166,N_660,N_1292);
and U3167 (N_3167,N_1231,N_294);
and U3168 (N_3168,N_1954,N_226);
or U3169 (N_3169,N_1040,N_1535);
xor U3170 (N_3170,N_941,N_456);
nand U3171 (N_3171,N_1470,N_158);
or U3172 (N_3172,N_183,N_911);
or U3173 (N_3173,N_1171,N_1785);
nor U3174 (N_3174,N_1093,N_1179);
or U3175 (N_3175,N_1160,N_1286);
xnor U3176 (N_3176,N_969,N_354);
nor U3177 (N_3177,N_1540,N_999);
and U3178 (N_3178,N_1803,N_1310);
nand U3179 (N_3179,N_648,N_1817);
or U3180 (N_3180,N_978,N_1565);
nor U3181 (N_3181,N_1434,N_773);
nand U3182 (N_3182,N_1829,N_58);
nor U3183 (N_3183,N_599,N_858);
or U3184 (N_3184,N_169,N_365);
xor U3185 (N_3185,N_1140,N_1166);
and U3186 (N_3186,N_1682,N_635);
nand U3187 (N_3187,N_1794,N_470);
and U3188 (N_3188,N_42,N_113);
or U3189 (N_3189,N_1698,N_572);
and U3190 (N_3190,N_284,N_1279);
and U3191 (N_3191,N_105,N_173);
or U3192 (N_3192,N_1211,N_442);
xor U3193 (N_3193,N_573,N_153);
xnor U3194 (N_3194,N_1467,N_768);
nand U3195 (N_3195,N_640,N_1762);
and U3196 (N_3196,N_452,N_1047);
and U3197 (N_3197,N_1626,N_782);
nor U3198 (N_3198,N_1816,N_625);
and U3199 (N_3199,N_682,N_1009);
or U3200 (N_3200,N_537,N_1167);
and U3201 (N_3201,N_1711,N_1244);
and U3202 (N_3202,N_939,N_1567);
and U3203 (N_3203,N_1611,N_512);
nand U3204 (N_3204,N_606,N_981);
xnor U3205 (N_3205,N_1019,N_1811);
nor U3206 (N_3206,N_164,N_461);
and U3207 (N_3207,N_447,N_72);
xnor U3208 (N_3208,N_1422,N_725);
xnor U3209 (N_3209,N_1253,N_1450);
nand U3210 (N_3210,N_750,N_1158);
or U3211 (N_3211,N_91,N_347);
xnor U3212 (N_3212,N_157,N_1926);
or U3213 (N_3213,N_578,N_1310);
or U3214 (N_3214,N_1059,N_34);
or U3215 (N_3215,N_1426,N_1554);
and U3216 (N_3216,N_256,N_511);
and U3217 (N_3217,N_1635,N_385);
nand U3218 (N_3218,N_1495,N_1949);
nor U3219 (N_3219,N_1159,N_123);
or U3220 (N_3220,N_548,N_95);
or U3221 (N_3221,N_208,N_275);
nand U3222 (N_3222,N_56,N_683);
nand U3223 (N_3223,N_555,N_1864);
and U3224 (N_3224,N_1875,N_1008);
or U3225 (N_3225,N_1889,N_408);
nor U3226 (N_3226,N_1586,N_932);
and U3227 (N_3227,N_1800,N_216);
and U3228 (N_3228,N_1973,N_813);
nand U3229 (N_3229,N_550,N_946);
nor U3230 (N_3230,N_1761,N_1517);
xor U3231 (N_3231,N_1449,N_1024);
and U3232 (N_3232,N_213,N_765);
and U3233 (N_3233,N_798,N_1229);
or U3234 (N_3234,N_1599,N_1197);
or U3235 (N_3235,N_1823,N_738);
or U3236 (N_3236,N_1117,N_885);
and U3237 (N_3237,N_947,N_153);
nand U3238 (N_3238,N_106,N_1684);
and U3239 (N_3239,N_1622,N_695);
xor U3240 (N_3240,N_835,N_1601);
and U3241 (N_3241,N_560,N_1163);
nand U3242 (N_3242,N_1733,N_309);
nor U3243 (N_3243,N_1427,N_926);
and U3244 (N_3244,N_1544,N_635);
nand U3245 (N_3245,N_1077,N_960);
xor U3246 (N_3246,N_534,N_628);
xor U3247 (N_3247,N_123,N_1592);
nand U3248 (N_3248,N_679,N_1424);
or U3249 (N_3249,N_1513,N_700);
nand U3250 (N_3250,N_731,N_1747);
nand U3251 (N_3251,N_1232,N_1966);
nand U3252 (N_3252,N_1266,N_950);
nand U3253 (N_3253,N_882,N_1556);
nor U3254 (N_3254,N_1477,N_1847);
nor U3255 (N_3255,N_1207,N_421);
nor U3256 (N_3256,N_897,N_850);
or U3257 (N_3257,N_954,N_315);
and U3258 (N_3258,N_778,N_202);
or U3259 (N_3259,N_578,N_1470);
and U3260 (N_3260,N_1730,N_523);
nor U3261 (N_3261,N_141,N_632);
xor U3262 (N_3262,N_223,N_1824);
or U3263 (N_3263,N_1571,N_760);
nand U3264 (N_3264,N_264,N_1969);
nor U3265 (N_3265,N_356,N_1916);
or U3266 (N_3266,N_1890,N_1569);
or U3267 (N_3267,N_185,N_842);
xor U3268 (N_3268,N_1486,N_1474);
nor U3269 (N_3269,N_479,N_957);
xor U3270 (N_3270,N_1774,N_138);
xor U3271 (N_3271,N_91,N_182);
xnor U3272 (N_3272,N_1397,N_1243);
xnor U3273 (N_3273,N_1335,N_1756);
nand U3274 (N_3274,N_865,N_37);
xnor U3275 (N_3275,N_1273,N_250);
xor U3276 (N_3276,N_1811,N_309);
xor U3277 (N_3277,N_875,N_1618);
nor U3278 (N_3278,N_698,N_1485);
nor U3279 (N_3279,N_1239,N_360);
and U3280 (N_3280,N_907,N_193);
xor U3281 (N_3281,N_1003,N_988);
and U3282 (N_3282,N_1109,N_1257);
nor U3283 (N_3283,N_576,N_1489);
and U3284 (N_3284,N_1417,N_671);
nand U3285 (N_3285,N_1301,N_589);
nor U3286 (N_3286,N_1392,N_1152);
or U3287 (N_3287,N_1377,N_1418);
and U3288 (N_3288,N_685,N_25);
and U3289 (N_3289,N_1124,N_110);
nor U3290 (N_3290,N_867,N_1500);
and U3291 (N_3291,N_716,N_1862);
and U3292 (N_3292,N_1024,N_439);
nand U3293 (N_3293,N_1772,N_1598);
xnor U3294 (N_3294,N_84,N_1870);
or U3295 (N_3295,N_1872,N_1066);
nor U3296 (N_3296,N_138,N_1591);
xnor U3297 (N_3297,N_977,N_1369);
xnor U3298 (N_3298,N_253,N_1795);
xnor U3299 (N_3299,N_1675,N_809);
and U3300 (N_3300,N_505,N_1965);
nor U3301 (N_3301,N_188,N_1120);
nand U3302 (N_3302,N_197,N_1564);
xnor U3303 (N_3303,N_975,N_1708);
and U3304 (N_3304,N_877,N_1891);
and U3305 (N_3305,N_1897,N_210);
nor U3306 (N_3306,N_807,N_1409);
nand U3307 (N_3307,N_1265,N_321);
nand U3308 (N_3308,N_1936,N_477);
nor U3309 (N_3309,N_1374,N_1199);
nor U3310 (N_3310,N_1116,N_1749);
nor U3311 (N_3311,N_979,N_1681);
nand U3312 (N_3312,N_452,N_1704);
nor U3313 (N_3313,N_103,N_450);
xnor U3314 (N_3314,N_1236,N_925);
or U3315 (N_3315,N_396,N_1673);
and U3316 (N_3316,N_605,N_1530);
or U3317 (N_3317,N_572,N_1546);
xnor U3318 (N_3318,N_1314,N_528);
nand U3319 (N_3319,N_841,N_802);
or U3320 (N_3320,N_1662,N_1834);
xnor U3321 (N_3321,N_1763,N_1346);
xor U3322 (N_3322,N_1718,N_1510);
or U3323 (N_3323,N_1852,N_84);
nor U3324 (N_3324,N_1519,N_1215);
nor U3325 (N_3325,N_621,N_502);
and U3326 (N_3326,N_1523,N_1705);
and U3327 (N_3327,N_1560,N_526);
nand U3328 (N_3328,N_705,N_1319);
nor U3329 (N_3329,N_124,N_809);
nor U3330 (N_3330,N_44,N_1109);
and U3331 (N_3331,N_629,N_1756);
and U3332 (N_3332,N_1,N_72);
nand U3333 (N_3333,N_1460,N_921);
xor U3334 (N_3334,N_1773,N_1039);
or U3335 (N_3335,N_1939,N_1129);
xnor U3336 (N_3336,N_1891,N_671);
or U3337 (N_3337,N_378,N_476);
or U3338 (N_3338,N_1309,N_1988);
xnor U3339 (N_3339,N_465,N_860);
nand U3340 (N_3340,N_1420,N_232);
or U3341 (N_3341,N_1354,N_78);
and U3342 (N_3342,N_942,N_1208);
and U3343 (N_3343,N_349,N_718);
nor U3344 (N_3344,N_131,N_1992);
or U3345 (N_3345,N_430,N_845);
nand U3346 (N_3346,N_174,N_1333);
nor U3347 (N_3347,N_248,N_603);
xnor U3348 (N_3348,N_1445,N_220);
xnor U3349 (N_3349,N_762,N_808);
or U3350 (N_3350,N_1873,N_1585);
xor U3351 (N_3351,N_1434,N_595);
and U3352 (N_3352,N_1322,N_420);
nor U3353 (N_3353,N_601,N_1837);
xnor U3354 (N_3354,N_86,N_344);
xor U3355 (N_3355,N_786,N_1453);
and U3356 (N_3356,N_234,N_1797);
or U3357 (N_3357,N_1255,N_1196);
and U3358 (N_3358,N_1835,N_1341);
xor U3359 (N_3359,N_1655,N_840);
or U3360 (N_3360,N_835,N_1652);
nor U3361 (N_3361,N_1002,N_51);
nand U3362 (N_3362,N_905,N_1908);
or U3363 (N_3363,N_1605,N_1885);
nand U3364 (N_3364,N_543,N_707);
nand U3365 (N_3365,N_251,N_34);
nor U3366 (N_3366,N_397,N_425);
nor U3367 (N_3367,N_1554,N_1088);
and U3368 (N_3368,N_1308,N_1350);
or U3369 (N_3369,N_1972,N_26);
and U3370 (N_3370,N_230,N_1734);
nor U3371 (N_3371,N_1275,N_937);
xnor U3372 (N_3372,N_1315,N_1509);
xnor U3373 (N_3373,N_1013,N_130);
xnor U3374 (N_3374,N_1760,N_1170);
nor U3375 (N_3375,N_1182,N_1713);
nand U3376 (N_3376,N_1681,N_897);
or U3377 (N_3377,N_1333,N_1216);
and U3378 (N_3378,N_1188,N_1418);
and U3379 (N_3379,N_1981,N_564);
nor U3380 (N_3380,N_1748,N_1825);
nand U3381 (N_3381,N_47,N_42);
and U3382 (N_3382,N_1109,N_1204);
nand U3383 (N_3383,N_1889,N_1355);
or U3384 (N_3384,N_515,N_1352);
and U3385 (N_3385,N_1768,N_950);
and U3386 (N_3386,N_712,N_459);
and U3387 (N_3387,N_539,N_375);
xor U3388 (N_3388,N_1055,N_1451);
or U3389 (N_3389,N_1997,N_43);
nand U3390 (N_3390,N_1806,N_696);
nor U3391 (N_3391,N_556,N_1074);
and U3392 (N_3392,N_1354,N_147);
nor U3393 (N_3393,N_1570,N_82);
or U3394 (N_3394,N_1252,N_56);
nor U3395 (N_3395,N_1990,N_195);
xnor U3396 (N_3396,N_25,N_1600);
or U3397 (N_3397,N_107,N_99);
nor U3398 (N_3398,N_1093,N_873);
nor U3399 (N_3399,N_153,N_1783);
xnor U3400 (N_3400,N_1888,N_222);
or U3401 (N_3401,N_110,N_1433);
and U3402 (N_3402,N_1511,N_793);
xnor U3403 (N_3403,N_362,N_1046);
nor U3404 (N_3404,N_1840,N_117);
nor U3405 (N_3405,N_1123,N_810);
xnor U3406 (N_3406,N_480,N_722);
nand U3407 (N_3407,N_117,N_580);
nor U3408 (N_3408,N_1556,N_420);
or U3409 (N_3409,N_1403,N_155);
or U3410 (N_3410,N_760,N_1449);
nand U3411 (N_3411,N_108,N_1604);
xnor U3412 (N_3412,N_1461,N_1905);
nor U3413 (N_3413,N_679,N_1606);
xor U3414 (N_3414,N_1023,N_559);
nand U3415 (N_3415,N_1231,N_306);
nand U3416 (N_3416,N_1312,N_265);
or U3417 (N_3417,N_210,N_171);
or U3418 (N_3418,N_1632,N_634);
xor U3419 (N_3419,N_1427,N_75);
and U3420 (N_3420,N_6,N_1402);
xor U3421 (N_3421,N_656,N_960);
nor U3422 (N_3422,N_1535,N_320);
or U3423 (N_3423,N_581,N_117);
xnor U3424 (N_3424,N_575,N_339);
and U3425 (N_3425,N_1280,N_1117);
nand U3426 (N_3426,N_340,N_1514);
nand U3427 (N_3427,N_633,N_1516);
and U3428 (N_3428,N_334,N_1724);
xor U3429 (N_3429,N_1052,N_1144);
or U3430 (N_3430,N_1545,N_1732);
xor U3431 (N_3431,N_361,N_1722);
and U3432 (N_3432,N_1653,N_1075);
nand U3433 (N_3433,N_1653,N_1511);
or U3434 (N_3434,N_1859,N_160);
and U3435 (N_3435,N_253,N_258);
xnor U3436 (N_3436,N_214,N_1369);
nor U3437 (N_3437,N_986,N_1377);
xnor U3438 (N_3438,N_926,N_1322);
nand U3439 (N_3439,N_265,N_1645);
and U3440 (N_3440,N_372,N_679);
xnor U3441 (N_3441,N_345,N_1012);
or U3442 (N_3442,N_1835,N_378);
and U3443 (N_3443,N_1216,N_95);
xnor U3444 (N_3444,N_670,N_1479);
nand U3445 (N_3445,N_730,N_1845);
and U3446 (N_3446,N_1013,N_915);
and U3447 (N_3447,N_1448,N_438);
nor U3448 (N_3448,N_444,N_492);
and U3449 (N_3449,N_790,N_92);
or U3450 (N_3450,N_210,N_377);
nor U3451 (N_3451,N_901,N_283);
or U3452 (N_3452,N_1890,N_1401);
xor U3453 (N_3453,N_86,N_1687);
nand U3454 (N_3454,N_444,N_1945);
and U3455 (N_3455,N_1661,N_1068);
xnor U3456 (N_3456,N_1144,N_365);
xor U3457 (N_3457,N_1788,N_69);
xor U3458 (N_3458,N_851,N_888);
xnor U3459 (N_3459,N_1563,N_1665);
nand U3460 (N_3460,N_208,N_1625);
and U3461 (N_3461,N_1316,N_1408);
nand U3462 (N_3462,N_656,N_800);
nor U3463 (N_3463,N_236,N_1868);
nand U3464 (N_3464,N_1545,N_366);
or U3465 (N_3465,N_77,N_1773);
and U3466 (N_3466,N_1409,N_1905);
nand U3467 (N_3467,N_1159,N_1293);
nand U3468 (N_3468,N_803,N_1192);
nor U3469 (N_3469,N_1122,N_150);
nor U3470 (N_3470,N_1945,N_1196);
or U3471 (N_3471,N_5,N_705);
and U3472 (N_3472,N_484,N_1213);
or U3473 (N_3473,N_1315,N_491);
nand U3474 (N_3474,N_1183,N_679);
and U3475 (N_3475,N_93,N_1414);
nor U3476 (N_3476,N_1557,N_1638);
and U3477 (N_3477,N_761,N_1570);
and U3478 (N_3478,N_1455,N_683);
xnor U3479 (N_3479,N_18,N_1505);
nand U3480 (N_3480,N_1374,N_105);
and U3481 (N_3481,N_1408,N_86);
and U3482 (N_3482,N_1039,N_7);
nand U3483 (N_3483,N_1703,N_1728);
and U3484 (N_3484,N_41,N_220);
or U3485 (N_3485,N_1021,N_1088);
xor U3486 (N_3486,N_1429,N_1777);
nand U3487 (N_3487,N_1687,N_1557);
nand U3488 (N_3488,N_453,N_583);
and U3489 (N_3489,N_1425,N_1189);
and U3490 (N_3490,N_1042,N_958);
and U3491 (N_3491,N_1370,N_769);
and U3492 (N_3492,N_1692,N_596);
nor U3493 (N_3493,N_1270,N_383);
or U3494 (N_3494,N_1085,N_1117);
xor U3495 (N_3495,N_1644,N_896);
xnor U3496 (N_3496,N_1046,N_1347);
xor U3497 (N_3497,N_1980,N_1861);
nor U3498 (N_3498,N_761,N_292);
or U3499 (N_3499,N_554,N_1372);
xor U3500 (N_3500,N_1071,N_1642);
xnor U3501 (N_3501,N_1156,N_1249);
or U3502 (N_3502,N_1910,N_878);
and U3503 (N_3503,N_420,N_1138);
nand U3504 (N_3504,N_578,N_237);
nand U3505 (N_3505,N_1128,N_639);
or U3506 (N_3506,N_1614,N_1818);
and U3507 (N_3507,N_1143,N_179);
xnor U3508 (N_3508,N_589,N_782);
and U3509 (N_3509,N_561,N_1219);
nor U3510 (N_3510,N_1644,N_1282);
nor U3511 (N_3511,N_1538,N_1800);
nand U3512 (N_3512,N_1462,N_1300);
or U3513 (N_3513,N_571,N_493);
nand U3514 (N_3514,N_1470,N_610);
or U3515 (N_3515,N_147,N_236);
xnor U3516 (N_3516,N_78,N_1457);
or U3517 (N_3517,N_1178,N_847);
xor U3518 (N_3518,N_1319,N_1429);
or U3519 (N_3519,N_859,N_55);
xor U3520 (N_3520,N_831,N_217);
nand U3521 (N_3521,N_15,N_1566);
nor U3522 (N_3522,N_395,N_1988);
or U3523 (N_3523,N_342,N_189);
nand U3524 (N_3524,N_208,N_418);
and U3525 (N_3525,N_551,N_1426);
or U3526 (N_3526,N_1375,N_1967);
xor U3527 (N_3527,N_238,N_851);
xor U3528 (N_3528,N_125,N_983);
nor U3529 (N_3529,N_128,N_581);
xor U3530 (N_3530,N_1145,N_88);
nor U3531 (N_3531,N_1691,N_526);
xnor U3532 (N_3532,N_155,N_1584);
nand U3533 (N_3533,N_1858,N_997);
xor U3534 (N_3534,N_929,N_305);
nor U3535 (N_3535,N_1478,N_1528);
nor U3536 (N_3536,N_565,N_1696);
nand U3537 (N_3537,N_1492,N_564);
and U3538 (N_3538,N_1082,N_98);
and U3539 (N_3539,N_139,N_278);
xor U3540 (N_3540,N_801,N_1559);
nand U3541 (N_3541,N_1385,N_1930);
xor U3542 (N_3542,N_165,N_1963);
or U3543 (N_3543,N_1853,N_315);
xnor U3544 (N_3544,N_1196,N_767);
or U3545 (N_3545,N_1520,N_758);
nor U3546 (N_3546,N_1273,N_754);
xor U3547 (N_3547,N_861,N_333);
or U3548 (N_3548,N_848,N_1175);
or U3549 (N_3549,N_1217,N_1699);
and U3550 (N_3550,N_548,N_1519);
or U3551 (N_3551,N_1469,N_1520);
and U3552 (N_3552,N_256,N_1508);
nand U3553 (N_3553,N_366,N_663);
or U3554 (N_3554,N_1702,N_312);
or U3555 (N_3555,N_1947,N_1427);
nor U3556 (N_3556,N_678,N_964);
and U3557 (N_3557,N_1039,N_1940);
and U3558 (N_3558,N_1546,N_536);
xor U3559 (N_3559,N_478,N_869);
or U3560 (N_3560,N_617,N_543);
nor U3561 (N_3561,N_137,N_364);
nand U3562 (N_3562,N_1875,N_492);
xnor U3563 (N_3563,N_605,N_1516);
xor U3564 (N_3564,N_779,N_1254);
nor U3565 (N_3565,N_1706,N_1668);
nand U3566 (N_3566,N_1567,N_1872);
nor U3567 (N_3567,N_1470,N_208);
and U3568 (N_3568,N_586,N_1930);
nand U3569 (N_3569,N_1176,N_40);
xor U3570 (N_3570,N_1987,N_594);
nor U3571 (N_3571,N_1748,N_707);
and U3572 (N_3572,N_1410,N_1342);
or U3573 (N_3573,N_1759,N_237);
and U3574 (N_3574,N_1692,N_831);
and U3575 (N_3575,N_739,N_1234);
xnor U3576 (N_3576,N_1036,N_823);
nand U3577 (N_3577,N_1440,N_37);
nand U3578 (N_3578,N_1399,N_1445);
and U3579 (N_3579,N_1150,N_866);
nand U3580 (N_3580,N_205,N_1237);
and U3581 (N_3581,N_1220,N_977);
or U3582 (N_3582,N_1300,N_928);
or U3583 (N_3583,N_1406,N_676);
and U3584 (N_3584,N_1172,N_596);
xnor U3585 (N_3585,N_1990,N_800);
xor U3586 (N_3586,N_1782,N_1559);
xor U3587 (N_3587,N_434,N_1316);
and U3588 (N_3588,N_485,N_1763);
xor U3589 (N_3589,N_912,N_1222);
nor U3590 (N_3590,N_284,N_1816);
xor U3591 (N_3591,N_1619,N_331);
nor U3592 (N_3592,N_1032,N_348);
and U3593 (N_3593,N_73,N_513);
nand U3594 (N_3594,N_1078,N_121);
and U3595 (N_3595,N_1959,N_35);
and U3596 (N_3596,N_403,N_1963);
nand U3597 (N_3597,N_1471,N_588);
nand U3598 (N_3598,N_1760,N_1137);
nor U3599 (N_3599,N_1102,N_1947);
nor U3600 (N_3600,N_797,N_1979);
or U3601 (N_3601,N_1037,N_1904);
nand U3602 (N_3602,N_1900,N_338);
xor U3603 (N_3603,N_329,N_1983);
and U3604 (N_3604,N_1188,N_583);
nand U3605 (N_3605,N_1542,N_1884);
xor U3606 (N_3606,N_751,N_477);
and U3607 (N_3607,N_251,N_1315);
nand U3608 (N_3608,N_174,N_779);
nand U3609 (N_3609,N_482,N_1477);
nor U3610 (N_3610,N_1812,N_976);
and U3611 (N_3611,N_1906,N_1866);
xor U3612 (N_3612,N_1458,N_44);
and U3613 (N_3613,N_1667,N_414);
nand U3614 (N_3614,N_1064,N_1672);
nor U3615 (N_3615,N_1980,N_1011);
and U3616 (N_3616,N_540,N_844);
nand U3617 (N_3617,N_1291,N_1093);
nor U3618 (N_3618,N_222,N_608);
nand U3619 (N_3619,N_1928,N_122);
nor U3620 (N_3620,N_15,N_950);
and U3621 (N_3621,N_276,N_296);
nor U3622 (N_3622,N_494,N_462);
or U3623 (N_3623,N_1429,N_1569);
xor U3624 (N_3624,N_957,N_1794);
and U3625 (N_3625,N_1047,N_1728);
and U3626 (N_3626,N_1756,N_1279);
nor U3627 (N_3627,N_1549,N_1807);
nand U3628 (N_3628,N_1526,N_1315);
nand U3629 (N_3629,N_46,N_15);
nor U3630 (N_3630,N_1225,N_273);
nor U3631 (N_3631,N_1807,N_218);
and U3632 (N_3632,N_1274,N_838);
nand U3633 (N_3633,N_869,N_1517);
and U3634 (N_3634,N_656,N_576);
nor U3635 (N_3635,N_1387,N_878);
or U3636 (N_3636,N_1294,N_424);
and U3637 (N_3637,N_513,N_1275);
nor U3638 (N_3638,N_1130,N_353);
and U3639 (N_3639,N_1245,N_974);
or U3640 (N_3640,N_1436,N_1846);
nand U3641 (N_3641,N_864,N_1459);
nor U3642 (N_3642,N_1235,N_1407);
nand U3643 (N_3643,N_668,N_1347);
and U3644 (N_3644,N_1491,N_1545);
xor U3645 (N_3645,N_1663,N_855);
xnor U3646 (N_3646,N_1089,N_252);
nand U3647 (N_3647,N_798,N_208);
nor U3648 (N_3648,N_1516,N_1448);
and U3649 (N_3649,N_517,N_1671);
nor U3650 (N_3650,N_762,N_1646);
and U3651 (N_3651,N_766,N_147);
nor U3652 (N_3652,N_726,N_1146);
xnor U3653 (N_3653,N_1830,N_1359);
nor U3654 (N_3654,N_1727,N_942);
and U3655 (N_3655,N_1429,N_978);
nand U3656 (N_3656,N_805,N_1565);
and U3657 (N_3657,N_1044,N_47);
or U3658 (N_3658,N_349,N_466);
nand U3659 (N_3659,N_416,N_527);
or U3660 (N_3660,N_279,N_752);
and U3661 (N_3661,N_1355,N_1508);
nor U3662 (N_3662,N_1473,N_1543);
or U3663 (N_3663,N_371,N_1412);
xnor U3664 (N_3664,N_1650,N_1400);
and U3665 (N_3665,N_1736,N_671);
and U3666 (N_3666,N_268,N_1644);
and U3667 (N_3667,N_606,N_1567);
or U3668 (N_3668,N_1074,N_769);
nor U3669 (N_3669,N_1535,N_1476);
nand U3670 (N_3670,N_698,N_1832);
nand U3671 (N_3671,N_377,N_1952);
nand U3672 (N_3672,N_1649,N_395);
nor U3673 (N_3673,N_471,N_1142);
and U3674 (N_3674,N_1264,N_814);
xor U3675 (N_3675,N_741,N_1563);
xor U3676 (N_3676,N_1284,N_567);
nor U3677 (N_3677,N_1755,N_883);
and U3678 (N_3678,N_487,N_444);
xor U3679 (N_3679,N_1770,N_1092);
or U3680 (N_3680,N_1115,N_1771);
or U3681 (N_3681,N_993,N_1102);
xnor U3682 (N_3682,N_170,N_1357);
nand U3683 (N_3683,N_371,N_44);
or U3684 (N_3684,N_1983,N_1249);
nor U3685 (N_3685,N_711,N_875);
nand U3686 (N_3686,N_510,N_386);
nand U3687 (N_3687,N_1864,N_1731);
xor U3688 (N_3688,N_396,N_338);
nand U3689 (N_3689,N_300,N_1538);
nor U3690 (N_3690,N_718,N_1137);
and U3691 (N_3691,N_1270,N_215);
xor U3692 (N_3692,N_1428,N_551);
nand U3693 (N_3693,N_128,N_1072);
or U3694 (N_3694,N_1900,N_1017);
nor U3695 (N_3695,N_1891,N_675);
nor U3696 (N_3696,N_272,N_567);
or U3697 (N_3697,N_1190,N_1695);
nand U3698 (N_3698,N_943,N_1937);
nand U3699 (N_3699,N_999,N_418);
and U3700 (N_3700,N_1877,N_1731);
and U3701 (N_3701,N_980,N_1628);
xnor U3702 (N_3702,N_191,N_881);
xor U3703 (N_3703,N_1087,N_272);
and U3704 (N_3704,N_1205,N_1695);
and U3705 (N_3705,N_261,N_835);
or U3706 (N_3706,N_776,N_1580);
nor U3707 (N_3707,N_1646,N_437);
nor U3708 (N_3708,N_1692,N_453);
or U3709 (N_3709,N_357,N_1285);
nor U3710 (N_3710,N_1577,N_990);
and U3711 (N_3711,N_1735,N_564);
xor U3712 (N_3712,N_1685,N_1626);
and U3713 (N_3713,N_1935,N_492);
nand U3714 (N_3714,N_653,N_417);
and U3715 (N_3715,N_37,N_1072);
nand U3716 (N_3716,N_972,N_1930);
or U3717 (N_3717,N_1148,N_315);
nor U3718 (N_3718,N_412,N_1005);
and U3719 (N_3719,N_1680,N_902);
and U3720 (N_3720,N_45,N_553);
or U3721 (N_3721,N_1964,N_1643);
and U3722 (N_3722,N_63,N_163);
and U3723 (N_3723,N_736,N_955);
or U3724 (N_3724,N_535,N_560);
nor U3725 (N_3725,N_1224,N_1336);
and U3726 (N_3726,N_1247,N_1028);
or U3727 (N_3727,N_1309,N_1052);
nand U3728 (N_3728,N_1995,N_1238);
xnor U3729 (N_3729,N_1061,N_1148);
and U3730 (N_3730,N_599,N_1882);
xnor U3731 (N_3731,N_552,N_509);
and U3732 (N_3732,N_977,N_1973);
or U3733 (N_3733,N_692,N_1501);
nor U3734 (N_3734,N_990,N_1822);
nor U3735 (N_3735,N_1987,N_312);
xor U3736 (N_3736,N_738,N_1877);
nand U3737 (N_3737,N_272,N_66);
nor U3738 (N_3738,N_828,N_767);
nor U3739 (N_3739,N_760,N_1509);
or U3740 (N_3740,N_1091,N_591);
xnor U3741 (N_3741,N_656,N_1724);
nand U3742 (N_3742,N_1049,N_742);
and U3743 (N_3743,N_314,N_554);
or U3744 (N_3744,N_29,N_372);
nand U3745 (N_3745,N_1806,N_117);
and U3746 (N_3746,N_1273,N_689);
xnor U3747 (N_3747,N_314,N_1081);
nor U3748 (N_3748,N_53,N_945);
or U3749 (N_3749,N_934,N_668);
nand U3750 (N_3750,N_572,N_927);
nand U3751 (N_3751,N_169,N_1377);
nand U3752 (N_3752,N_1244,N_1822);
and U3753 (N_3753,N_766,N_988);
and U3754 (N_3754,N_1017,N_1053);
and U3755 (N_3755,N_561,N_1322);
and U3756 (N_3756,N_985,N_632);
xor U3757 (N_3757,N_1271,N_634);
and U3758 (N_3758,N_166,N_307);
nor U3759 (N_3759,N_635,N_1586);
nor U3760 (N_3760,N_226,N_1354);
and U3761 (N_3761,N_194,N_1748);
nand U3762 (N_3762,N_48,N_523);
nor U3763 (N_3763,N_944,N_1536);
or U3764 (N_3764,N_211,N_1135);
or U3765 (N_3765,N_210,N_815);
xor U3766 (N_3766,N_962,N_767);
nand U3767 (N_3767,N_492,N_402);
nor U3768 (N_3768,N_895,N_1265);
xor U3769 (N_3769,N_1825,N_1938);
nor U3770 (N_3770,N_1844,N_768);
nand U3771 (N_3771,N_1630,N_151);
xor U3772 (N_3772,N_920,N_1016);
or U3773 (N_3773,N_290,N_1073);
xnor U3774 (N_3774,N_1498,N_328);
nor U3775 (N_3775,N_137,N_1032);
nor U3776 (N_3776,N_1672,N_509);
nor U3777 (N_3777,N_660,N_190);
nand U3778 (N_3778,N_573,N_1713);
nand U3779 (N_3779,N_65,N_652);
nor U3780 (N_3780,N_793,N_1678);
or U3781 (N_3781,N_555,N_1401);
and U3782 (N_3782,N_472,N_1750);
nand U3783 (N_3783,N_1818,N_1969);
and U3784 (N_3784,N_496,N_1362);
and U3785 (N_3785,N_1624,N_1831);
xnor U3786 (N_3786,N_750,N_275);
and U3787 (N_3787,N_77,N_1064);
nor U3788 (N_3788,N_538,N_333);
nand U3789 (N_3789,N_583,N_392);
or U3790 (N_3790,N_312,N_135);
nor U3791 (N_3791,N_910,N_358);
nand U3792 (N_3792,N_534,N_1998);
and U3793 (N_3793,N_804,N_1082);
xor U3794 (N_3794,N_284,N_1911);
nand U3795 (N_3795,N_1836,N_458);
or U3796 (N_3796,N_1779,N_1659);
and U3797 (N_3797,N_853,N_407);
and U3798 (N_3798,N_1782,N_1776);
nor U3799 (N_3799,N_385,N_1307);
nand U3800 (N_3800,N_1535,N_187);
xnor U3801 (N_3801,N_1473,N_1579);
nand U3802 (N_3802,N_458,N_1456);
nand U3803 (N_3803,N_984,N_1570);
and U3804 (N_3804,N_269,N_902);
nand U3805 (N_3805,N_871,N_868);
and U3806 (N_3806,N_190,N_153);
or U3807 (N_3807,N_1660,N_990);
or U3808 (N_3808,N_253,N_76);
xor U3809 (N_3809,N_727,N_868);
nand U3810 (N_3810,N_63,N_1027);
xor U3811 (N_3811,N_1741,N_225);
and U3812 (N_3812,N_1951,N_1200);
or U3813 (N_3813,N_1794,N_166);
or U3814 (N_3814,N_1185,N_219);
and U3815 (N_3815,N_1007,N_1984);
xor U3816 (N_3816,N_1900,N_1605);
nand U3817 (N_3817,N_1190,N_1348);
xnor U3818 (N_3818,N_124,N_366);
xor U3819 (N_3819,N_204,N_23);
nor U3820 (N_3820,N_1259,N_553);
nor U3821 (N_3821,N_238,N_1741);
nand U3822 (N_3822,N_1828,N_1192);
or U3823 (N_3823,N_1697,N_1036);
xnor U3824 (N_3824,N_1327,N_631);
nand U3825 (N_3825,N_581,N_526);
nor U3826 (N_3826,N_364,N_608);
xor U3827 (N_3827,N_1381,N_990);
and U3828 (N_3828,N_690,N_308);
and U3829 (N_3829,N_513,N_401);
xor U3830 (N_3830,N_4,N_15);
nand U3831 (N_3831,N_1249,N_1964);
and U3832 (N_3832,N_1415,N_506);
nand U3833 (N_3833,N_1130,N_1926);
xnor U3834 (N_3834,N_625,N_370);
nor U3835 (N_3835,N_1081,N_1114);
xnor U3836 (N_3836,N_1750,N_818);
nand U3837 (N_3837,N_1723,N_1388);
xor U3838 (N_3838,N_912,N_856);
nor U3839 (N_3839,N_1623,N_63);
xnor U3840 (N_3840,N_1775,N_55);
nor U3841 (N_3841,N_235,N_929);
nand U3842 (N_3842,N_274,N_1635);
nor U3843 (N_3843,N_421,N_610);
nand U3844 (N_3844,N_1296,N_257);
and U3845 (N_3845,N_1106,N_1272);
xnor U3846 (N_3846,N_632,N_286);
nor U3847 (N_3847,N_1456,N_1025);
and U3848 (N_3848,N_1196,N_685);
xnor U3849 (N_3849,N_1563,N_659);
xnor U3850 (N_3850,N_1053,N_721);
nand U3851 (N_3851,N_926,N_1760);
or U3852 (N_3852,N_661,N_136);
or U3853 (N_3853,N_1068,N_1089);
xnor U3854 (N_3854,N_732,N_1863);
nor U3855 (N_3855,N_794,N_766);
nor U3856 (N_3856,N_1549,N_262);
nand U3857 (N_3857,N_661,N_66);
or U3858 (N_3858,N_491,N_1771);
nand U3859 (N_3859,N_774,N_126);
and U3860 (N_3860,N_1385,N_1148);
xnor U3861 (N_3861,N_74,N_1106);
xnor U3862 (N_3862,N_417,N_253);
nand U3863 (N_3863,N_333,N_1199);
nand U3864 (N_3864,N_409,N_320);
xor U3865 (N_3865,N_1404,N_99);
nor U3866 (N_3866,N_153,N_1912);
or U3867 (N_3867,N_1976,N_1186);
xnor U3868 (N_3868,N_892,N_169);
or U3869 (N_3869,N_1084,N_1894);
and U3870 (N_3870,N_1158,N_1828);
nor U3871 (N_3871,N_574,N_1173);
and U3872 (N_3872,N_496,N_770);
nor U3873 (N_3873,N_1054,N_1175);
and U3874 (N_3874,N_1463,N_1612);
xnor U3875 (N_3875,N_787,N_926);
nand U3876 (N_3876,N_1609,N_1473);
nor U3877 (N_3877,N_1590,N_978);
nand U3878 (N_3878,N_1639,N_1531);
and U3879 (N_3879,N_550,N_172);
nor U3880 (N_3880,N_1135,N_1339);
and U3881 (N_3881,N_1221,N_1738);
or U3882 (N_3882,N_528,N_663);
and U3883 (N_3883,N_835,N_805);
and U3884 (N_3884,N_388,N_1667);
and U3885 (N_3885,N_1308,N_858);
xnor U3886 (N_3886,N_577,N_501);
xor U3887 (N_3887,N_140,N_726);
nand U3888 (N_3888,N_927,N_444);
and U3889 (N_3889,N_1767,N_1836);
nor U3890 (N_3890,N_1059,N_449);
nand U3891 (N_3891,N_1675,N_1113);
xor U3892 (N_3892,N_1870,N_725);
nor U3893 (N_3893,N_659,N_1930);
or U3894 (N_3894,N_1618,N_741);
and U3895 (N_3895,N_574,N_907);
and U3896 (N_3896,N_1864,N_44);
and U3897 (N_3897,N_1574,N_553);
or U3898 (N_3898,N_1187,N_1899);
nor U3899 (N_3899,N_186,N_727);
nand U3900 (N_3900,N_1351,N_941);
xor U3901 (N_3901,N_1491,N_610);
xor U3902 (N_3902,N_1194,N_1453);
and U3903 (N_3903,N_1409,N_1461);
nand U3904 (N_3904,N_194,N_642);
or U3905 (N_3905,N_591,N_193);
and U3906 (N_3906,N_1201,N_1168);
or U3907 (N_3907,N_796,N_1491);
nand U3908 (N_3908,N_1168,N_521);
or U3909 (N_3909,N_874,N_1074);
or U3910 (N_3910,N_1543,N_8);
nor U3911 (N_3911,N_1751,N_727);
nand U3912 (N_3912,N_309,N_1963);
and U3913 (N_3913,N_1797,N_1473);
xor U3914 (N_3914,N_1591,N_448);
nor U3915 (N_3915,N_916,N_1456);
nor U3916 (N_3916,N_487,N_1164);
nor U3917 (N_3917,N_228,N_1730);
and U3918 (N_3918,N_697,N_1981);
xor U3919 (N_3919,N_1128,N_1776);
nor U3920 (N_3920,N_908,N_1333);
nand U3921 (N_3921,N_99,N_785);
or U3922 (N_3922,N_756,N_1185);
nand U3923 (N_3923,N_1579,N_74);
nand U3924 (N_3924,N_1992,N_299);
nor U3925 (N_3925,N_1202,N_397);
nor U3926 (N_3926,N_364,N_1721);
nand U3927 (N_3927,N_1859,N_1918);
and U3928 (N_3928,N_1889,N_14);
or U3929 (N_3929,N_373,N_789);
xor U3930 (N_3930,N_1043,N_1955);
and U3931 (N_3931,N_1896,N_1858);
xnor U3932 (N_3932,N_947,N_371);
and U3933 (N_3933,N_507,N_1919);
nand U3934 (N_3934,N_1824,N_1156);
or U3935 (N_3935,N_1477,N_1865);
xnor U3936 (N_3936,N_28,N_650);
xor U3937 (N_3937,N_1267,N_920);
nor U3938 (N_3938,N_432,N_1013);
xor U3939 (N_3939,N_424,N_261);
and U3940 (N_3940,N_1218,N_1197);
nand U3941 (N_3941,N_1930,N_209);
and U3942 (N_3942,N_1169,N_1008);
or U3943 (N_3943,N_795,N_1628);
or U3944 (N_3944,N_899,N_799);
xor U3945 (N_3945,N_1309,N_213);
nor U3946 (N_3946,N_1549,N_1198);
nor U3947 (N_3947,N_395,N_1180);
nand U3948 (N_3948,N_459,N_988);
or U3949 (N_3949,N_786,N_1417);
nand U3950 (N_3950,N_893,N_1565);
nor U3951 (N_3951,N_743,N_1806);
nor U3952 (N_3952,N_1898,N_1744);
nand U3953 (N_3953,N_60,N_261);
nor U3954 (N_3954,N_730,N_1549);
xnor U3955 (N_3955,N_1430,N_1996);
or U3956 (N_3956,N_1283,N_1960);
xor U3957 (N_3957,N_347,N_455);
nor U3958 (N_3958,N_1367,N_1843);
or U3959 (N_3959,N_1846,N_1862);
nand U3960 (N_3960,N_365,N_1748);
nor U3961 (N_3961,N_1275,N_882);
nand U3962 (N_3962,N_1534,N_603);
nor U3963 (N_3963,N_973,N_395);
xor U3964 (N_3964,N_1513,N_95);
nor U3965 (N_3965,N_1324,N_1609);
and U3966 (N_3966,N_285,N_1011);
xnor U3967 (N_3967,N_228,N_1096);
xnor U3968 (N_3968,N_1115,N_829);
and U3969 (N_3969,N_276,N_755);
or U3970 (N_3970,N_1941,N_1819);
xor U3971 (N_3971,N_143,N_1010);
or U3972 (N_3972,N_182,N_1268);
nand U3973 (N_3973,N_1544,N_881);
xor U3974 (N_3974,N_63,N_1556);
nand U3975 (N_3975,N_1158,N_1825);
or U3976 (N_3976,N_137,N_1223);
or U3977 (N_3977,N_1566,N_895);
xor U3978 (N_3978,N_948,N_1597);
nor U3979 (N_3979,N_1009,N_684);
and U3980 (N_3980,N_1966,N_1717);
nand U3981 (N_3981,N_1802,N_1234);
nor U3982 (N_3982,N_1659,N_930);
and U3983 (N_3983,N_1221,N_773);
xnor U3984 (N_3984,N_220,N_262);
and U3985 (N_3985,N_1852,N_1622);
nand U3986 (N_3986,N_1970,N_896);
or U3987 (N_3987,N_526,N_1477);
nor U3988 (N_3988,N_1059,N_1141);
or U3989 (N_3989,N_242,N_1259);
and U3990 (N_3990,N_1,N_1172);
nor U3991 (N_3991,N_1969,N_1543);
nor U3992 (N_3992,N_1140,N_152);
and U3993 (N_3993,N_107,N_1950);
xor U3994 (N_3994,N_1207,N_1390);
and U3995 (N_3995,N_656,N_1721);
or U3996 (N_3996,N_1524,N_312);
nor U3997 (N_3997,N_1468,N_887);
nand U3998 (N_3998,N_661,N_1362);
nand U3999 (N_3999,N_884,N_761);
and U4000 (N_4000,N_2199,N_3929);
nand U4001 (N_4001,N_2900,N_2757);
nor U4002 (N_4002,N_2304,N_2941);
nand U4003 (N_4003,N_2783,N_2574);
or U4004 (N_4004,N_2214,N_3866);
xor U4005 (N_4005,N_3449,N_3419);
xor U4006 (N_4006,N_2732,N_2874);
xnor U4007 (N_4007,N_3757,N_3874);
nand U4008 (N_4008,N_2228,N_3243);
and U4009 (N_4009,N_3325,N_2688);
nor U4010 (N_4010,N_2906,N_2849);
nand U4011 (N_4011,N_3463,N_3340);
nand U4012 (N_4012,N_3105,N_2240);
and U4013 (N_4013,N_2314,N_3931);
nor U4014 (N_4014,N_2663,N_3746);
and U4015 (N_4015,N_2829,N_2353);
nand U4016 (N_4016,N_3308,N_3457);
or U4017 (N_4017,N_2258,N_3290);
and U4018 (N_4018,N_2601,N_2848);
nand U4019 (N_4019,N_3641,N_3298);
nand U4020 (N_4020,N_3318,N_3333);
and U4021 (N_4021,N_3351,N_2492);
nor U4022 (N_4022,N_3363,N_3612);
and U4023 (N_4023,N_2552,N_2876);
nand U4024 (N_4024,N_3770,N_2315);
and U4025 (N_4025,N_3125,N_3403);
nand U4026 (N_4026,N_3763,N_2218);
nand U4027 (N_4027,N_2969,N_2821);
and U4028 (N_4028,N_2348,N_2665);
and U4029 (N_4029,N_2740,N_2145);
xor U4030 (N_4030,N_2632,N_3209);
nand U4031 (N_4031,N_3203,N_2546);
xnor U4032 (N_4032,N_2253,N_3794);
nand U4033 (N_4033,N_3568,N_3621);
and U4034 (N_4034,N_3188,N_2907);
xor U4035 (N_4035,N_2466,N_3811);
or U4036 (N_4036,N_3386,N_3010);
xor U4037 (N_4037,N_2898,N_2998);
and U4038 (N_4038,N_2417,N_3312);
nand U4039 (N_4039,N_3836,N_3354);
and U4040 (N_4040,N_2249,N_2010);
or U4041 (N_4041,N_2624,N_2252);
xor U4042 (N_4042,N_3075,N_2071);
and U4043 (N_4043,N_3091,N_3572);
xor U4044 (N_4044,N_3905,N_2099);
nor U4045 (N_4045,N_3971,N_3862);
nand U4046 (N_4046,N_3803,N_3431);
or U4047 (N_4047,N_2768,N_2398);
and U4048 (N_4048,N_2566,N_3838);
and U4049 (N_4049,N_2681,N_3871);
xor U4050 (N_4050,N_3288,N_3565);
and U4051 (N_4051,N_2208,N_2489);
or U4052 (N_4052,N_2739,N_3466);
xnor U4053 (N_4053,N_2058,N_3402);
and U4054 (N_4054,N_2219,N_2483);
or U4055 (N_4055,N_3528,N_3181);
nor U4056 (N_4056,N_2879,N_3983);
or U4057 (N_4057,N_2441,N_2079);
nor U4058 (N_4058,N_3549,N_2808);
nor U4059 (N_4059,N_2003,N_3483);
and U4060 (N_4060,N_3408,N_2231);
nor U4061 (N_4061,N_2561,N_3527);
nor U4062 (N_4062,N_2582,N_3121);
nor U4063 (N_4063,N_3877,N_3100);
xor U4064 (N_4064,N_2536,N_3057);
and U4065 (N_4065,N_2237,N_2480);
and U4066 (N_4066,N_2702,N_3782);
nand U4067 (N_4067,N_3192,N_2434);
or U4068 (N_4068,N_3675,N_3124);
xor U4069 (N_4069,N_3644,N_2455);
nor U4070 (N_4070,N_2795,N_2523);
nor U4071 (N_4071,N_3586,N_2952);
xnor U4072 (N_4072,N_3035,N_3952);
xor U4073 (N_4073,N_3812,N_3567);
nor U4074 (N_4074,N_3126,N_2356);
nor U4075 (N_4075,N_2942,N_2564);
xnor U4076 (N_4076,N_2467,N_2392);
nand U4077 (N_4077,N_2400,N_3349);
nand U4078 (N_4078,N_2233,N_2696);
xnor U4079 (N_4079,N_2838,N_3821);
nor U4080 (N_4080,N_2097,N_2837);
xor U4081 (N_4081,N_2641,N_3392);
xor U4082 (N_4082,N_2504,N_2769);
nand U4083 (N_4083,N_2568,N_2770);
nor U4084 (N_4084,N_2149,N_2081);
nand U4085 (N_4085,N_2545,N_3835);
nand U4086 (N_4086,N_2654,N_3008);
and U4087 (N_4087,N_2708,N_3226);
or U4088 (N_4088,N_3063,N_2130);
xnor U4089 (N_4089,N_3603,N_2780);
or U4090 (N_4090,N_3191,N_2432);
nand U4091 (N_4091,N_3925,N_3446);
xor U4092 (N_4092,N_2805,N_2767);
xor U4093 (N_4093,N_3602,N_3269);
nor U4094 (N_4094,N_2476,N_3564);
nand U4095 (N_4095,N_2494,N_3264);
nand U4096 (N_4096,N_2815,N_3393);
or U4097 (N_4097,N_3005,N_2435);
and U4098 (N_4098,N_2468,N_2165);
nand U4099 (N_4099,N_3535,N_3516);
xor U4100 (N_4100,N_3487,N_3132);
nor U4101 (N_4101,N_3846,N_3982);
or U4102 (N_4102,N_3588,N_3222);
nand U4103 (N_4103,N_3816,N_3878);
and U4104 (N_4104,N_2322,N_2448);
and U4105 (N_4105,N_3941,N_2736);
nand U4106 (N_4106,N_2285,N_2419);
nor U4107 (N_4107,N_3872,N_2096);
nand U4108 (N_4108,N_2631,N_2349);
xor U4109 (N_4109,N_3016,N_2313);
and U4110 (N_4110,N_3414,N_2728);
nand U4111 (N_4111,N_3475,N_3169);
xor U4112 (N_4112,N_3083,N_3617);
and U4113 (N_4113,N_3252,N_2008);
nand U4114 (N_4114,N_2430,N_2486);
xor U4115 (N_4115,N_3973,N_2209);
nor U4116 (N_4116,N_2800,N_2890);
nor U4117 (N_4117,N_3949,N_3537);
or U4118 (N_4118,N_2645,N_3421);
or U4119 (N_4119,N_2875,N_3037);
and U4120 (N_4120,N_2423,N_3733);
or U4121 (N_4121,N_3765,N_3476);
or U4122 (N_4122,N_2029,N_2181);
xor U4123 (N_4123,N_3798,N_2060);
xnor U4124 (N_4124,N_3906,N_2382);
nand U4125 (N_4125,N_2431,N_2034);
nand U4126 (N_4126,N_2857,N_2778);
and U4127 (N_4127,N_2286,N_2014);
nand U4128 (N_4128,N_2028,N_2174);
and U4129 (N_4129,N_2092,N_2465);
and U4130 (N_4130,N_2968,N_2846);
nor U4131 (N_4131,N_3719,N_2691);
nand U4132 (N_4132,N_2731,N_3923);
nand U4133 (N_4133,N_2446,N_2451);
and U4134 (N_4134,N_2371,N_2618);
or U4135 (N_4135,N_3772,N_3730);
nor U4136 (N_4136,N_3976,N_3825);
xor U4137 (N_4137,N_3359,N_3186);
xnor U4138 (N_4138,N_3627,N_2672);
and U4139 (N_4139,N_2461,N_2810);
and U4140 (N_4140,N_3227,N_2152);
xnor U4141 (N_4141,N_3331,N_2548);
nand U4142 (N_4142,N_3093,N_2171);
xnor U4143 (N_4143,N_2513,N_3390);
and U4144 (N_4144,N_3512,N_2527);
xnor U4145 (N_4145,N_3703,N_3357);
or U4146 (N_4146,N_3728,N_3070);
and U4147 (N_4147,N_2229,N_3190);
xor U4148 (N_4148,N_3807,N_2213);
or U4149 (N_4149,N_3805,N_3143);
nor U4150 (N_4150,N_2236,N_2210);
xnor U4151 (N_4151,N_2606,N_3287);
nor U4152 (N_4152,N_2717,N_2429);
nand U4153 (N_4153,N_3102,N_2019);
nand U4154 (N_4154,N_2211,N_2311);
xor U4155 (N_4155,N_2343,N_2345);
nor U4156 (N_4156,N_2359,N_2200);
or U4157 (N_4157,N_2710,N_2299);
nand U4158 (N_4158,N_2526,N_3336);
or U4159 (N_4159,N_3296,N_2608);
nor U4160 (N_4160,N_2027,N_2949);
and U4161 (N_4161,N_3327,N_3120);
or U4162 (N_4162,N_2743,N_2799);
nor U4163 (N_4163,N_3944,N_2948);
nand U4164 (N_4164,N_3684,N_2976);
xnor U4165 (N_4165,N_2648,N_3754);
or U4166 (N_4166,N_2847,N_2581);
nand U4167 (N_4167,N_2617,N_3558);
xor U4168 (N_4168,N_2960,N_2551);
nand U4169 (N_4169,N_2659,N_3793);
nor U4170 (N_4170,N_2675,N_3271);
or U4171 (N_4171,N_3249,N_3946);
and U4172 (N_4172,N_2281,N_3040);
nor U4173 (N_4173,N_3999,N_3180);
nor U4174 (N_4174,N_2414,N_2133);
nor U4175 (N_4175,N_2943,N_3638);
and U4176 (N_4176,N_2365,N_2487);
or U4177 (N_4177,N_3470,N_3267);
or U4178 (N_4178,N_3094,N_2610);
nor U4179 (N_4179,N_2031,N_3751);
or U4180 (N_4180,N_2753,N_3021);
or U4181 (N_4181,N_3240,N_2062);
or U4182 (N_4182,N_2297,N_2341);
xor U4183 (N_4183,N_2926,N_2626);
xor U4184 (N_4184,N_2784,N_2988);
and U4185 (N_4185,N_3117,N_2711);
xnor U4186 (N_4186,N_3755,N_3097);
nand U4187 (N_4187,N_2336,N_2911);
or U4188 (N_4188,N_2093,N_3954);
xnor U4189 (N_4189,N_2819,N_3508);
nor U4190 (N_4190,N_2761,N_2666);
xnor U4191 (N_4191,N_2354,N_2168);
and U4192 (N_4192,N_3967,N_3593);
and U4193 (N_4193,N_2685,N_3458);
xnor U4194 (N_4194,N_3138,N_3001);
nor U4195 (N_4195,N_2647,N_2039);
nand U4196 (N_4196,N_3039,N_3088);
and U4197 (N_4197,N_3864,N_2589);
or U4198 (N_4198,N_3560,N_3590);
and U4199 (N_4199,N_3334,N_3686);
nand U4200 (N_4200,N_3050,N_2169);
xor U4201 (N_4201,N_3631,N_2161);
or U4202 (N_4202,N_2403,N_3277);
and U4203 (N_4203,N_3199,N_2310);
and U4204 (N_4204,N_2505,N_2057);
xnor U4205 (N_4205,N_2289,N_2089);
and U4206 (N_4206,N_2444,N_3827);
nand U4207 (N_4207,N_3320,N_3036);
and U4208 (N_4208,N_3337,N_2918);
xor U4209 (N_4209,N_2103,N_2139);
and U4210 (N_4210,N_2215,N_3101);
nand U4211 (N_4211,N_3865,N_2335);
nor U4212 (N_4212,N_3348,N_3116);
nor U4213 (N_4213,N_3231,N_3651);
nor U4214 (N_4214,N_3921,N_3955);
nor U4215 (N_4215,N_2381,N_2571);
or U4216 (N_4216,N_2801,N_2121);
and U4217 (N_4217,N_3734,N_2687);
xnor U4218 (N_4218,N_2883,N_3996);
nand U4219 (N_4219,N_3851,N_2806);
nand U4220 (N_4220,N_2995,N_3215);
or U4221 (N_4221,N_3934,N_2195);
nor U4222 (N_4222,N_3969,N_3407);
and U4223 (N_4223,N_2892,N_2189);
and U4224 (N_4224,N_3064,N_3785);
xor U4225 (N_4225,N_2756,N_3498);
xor U4226 (N_4226,N_3702,N_2501);
or U4227 (N_4227,N_3889,N_3007);
or U4228 (N_4228,N_2100,N_2774);
nor U4229 (N_4229,N_3701,N_3899);
and U4230 (N_4230,N_2964,N_2935);
nand U4231 (N_4231,N_3551,N_2790);
and U4232 (N_4232,N_3898,N_3342);
nand U4233 (N_4233,N_3669,N_2026);
nor U4234 (N_4234,N_3176,N_3854);
nor U4235 (N_4235,N_3646,N_3553);
and U4236 (N_4236,N_3784,N_2813);
nor U4237 (N_4237,N_2167,N_3375);
or U4238 (N_4238,N_3009,N_3778);
or U4239 (N_4239,N_2376,N_2378);
xor U4240 (N_4240,N_3900,N_2114);
and U4241 (N_4241,N_3709,N_2042);
xnor U4242 (N_4242,N_2980,N_3647);
nor U4243 (N_4243,N_2817,N_3740);
or U4244 (N_4244,N_2190,N_2138);
nor U4245 (N_4245,N_2458,N_2294);
nor U4246 (N_4246,N_2803,N_3429);
or U4247 (N_4247,N_3073,N_2814);
xnor U4248 (N_4248,N_2424,N_3219);
and U4249 (N_4249,N_2202,N_2540);
xnor U4250 (N_4250,N_2120,N_3026);
nand U4251 (N_4251,N_3748,N_3945);
nand U4252 (N_4252,N_2604,N_2970);
xnor U4253 (N_4253,N_2987,N_2366);
or U4254 (N_4254,N_2035,N_2503);
nand U4255 (N_4255,N_3066,N_2021);
nand U4256 (N_4256,N_2325,N_2490);
nand U4257 (N_4257,N_3828,N_2357);
nor U4258 (N_4258,N_2113,N_3013);
or U4259 (N_4259,N_2607,N_2957);
and U4260 (N_4260,N_3980,N_3486);
nor U4261 (N_4261,N_3912,N_3167);
nand U4262 (N_4262,N_3159,N_2677);
nand U4263 (N_4263,N_2276,N_3711);
xor U4264 (N_4264,N_2535,N_3426);
xor U4265 (N_4265,N_3817,N_3937);
nor U4266 (N_4266,N_2390,N_2183);
xor U4267 (N_4267,N_2098,N_2088);
and U4268 (N_4268,N_3149,N_2971);
nor U4269 (N_4269,N_3310,N_3441);
xor U4270 (N_4270,N_3940,N_3510);
xor U4271 (N_4271,N_3196,N_3129);
and U4272 (N_4272,N_3975,N_2940);
nand U4273 (N_4273,N_3067,N_3378);
and U4274 (N_4274,N_2506,N_2525);
nor U4275 (N_4275,N_2726,N_2575);
or U4276 (N_4276,N_2061,N_3781);
xor U4277 (N_4277,N_3515,N_2766);
nand U4278 (N_4278,N_2497,N_2257);
or U4279 (N_4279,N_2084,N_3089);
and U4280 (N_4280,N_3238,N_2409);
or U4281 (N_4281,N_3847,N_3096);
or U4282 (N_4282,N_2981,N_2407);
and U4283 (N_4283,N_3724,N_3165);
and U4284 (N_4284,N_3536,N_3494);
or U4285 (N_4285,N_3843,N_3056);
or U4286 (N_4286,N_2695,N_3761);
and U4287 (N_4287,N_3532,N_3801);
nor U4288 (N_4288,N_2318,N_2004);
and U4289 (N_4289,N_3248,N_2983);
xor U4290 (N_4290,N_3777,N_2232);
nor U4291 (N_4291,N_2339,N_3541);
nor U4292 (N_4292,N_3552,N_3894);
nand U4293 (N_4293,N_3883,N_3480);
or U4294 (N_4294,N_2226,N_3239);
and U4295 (N_4295,N_2333,N_2261);
xor U4296 (N_4296,N_2760,N_3721);
nand U4297 (N_4297,N_3493,N_3632);
xor U4298 (N_4298,N_2812,N_3563);
nand U4299 (N_4299,N_2191,N_3489);
and U4300 (N_4300,N_2298,N_3488);
xor U4301 (N_4301,N_3957,N_2786);
xnor U4302 (N_4302,N_2277,N_3984);
nor U4303 (N_4303,N_3373,N_3525);
xnor U4304 (N_4304,N_3398,N_2243);
nand U4305 (N_4305,N_2899,N_2765);
or U4306 (N_4306,N_3385,N_2745);
xor U4307 (N_4307,N_2238,N_3428);
and U4308 (N_4308,N_3682,N_3942);
nand U4309 (N_4309,N_3915,N_2671);
or U4310 (N_4310,N_3388,N_3867);
and U4311 (N_4311,N_3034,N_2205);
nand U4312 (N_4312,N_2723,N_2246);
and U4313 (N_4313,N_3585,N_2854);
nor U4314 (N_4314,N_3744,N_3274);
xor U4315 (N_4315,N_2629,N_2358);
and U4316 (N_4316,N_3909,N_2402);
xor U4317 (N_4317,N_2603,N_2499);
and U4318 (N_4318,N_3321,N_3306);
xor U4319 (N_4319,N_2676,N_3051);
nor U4320 (N_4320,N_2993,N_3170);
nor U4321 (N_4321,N_3459,N_2612);
and U4322 (N_4322,N_3662,N_2377);
or U4323 (N_4323,N_3689,N_2040);
or U4324 (N_4324,N_2683,N_3988);
and U4325 (N_4325,N_2108,N_3078);
nor U4326 (N_4326,N_2420,N_2462);
or U4327 (N_4327,N_3216,N_2894);
xnor U4328 (N_4328,N_3384,N_3762);
nand U4329 (N_4329,N_2101,N_3972);
nor U4330 (N_4330,N_3224,N_2186);
or U4331 (N_4331,N_2234,N_3346);
nor U4332 (N_4332,N_3233,N_2599);
nand U4333 (N_4333,N_3573,N_3241);
and U4334 (N_4334,N_3890,N_2712);
nor U4335 (N_4335,N_2919,N_2045);
nor U4336 (N_4336,N_2584,N_2156);
xnor U4337 (N_4337,N_2818,N_2495);
and U4338 (N_4338,N_2146,N_2771);
nand U4339 (N_4339,N_3752,N_2449);
nor U4340 (N_4340,N_3456,N_3053);
xor U4341 (N_4341,N_3658,N_3205);
nand U4342 (N_4342,N_3491,N_3687);
and U4343 (N_4343,N_3304,N_2839);
nand U4344 (N_4344,N_2331,N_3897);
and U4345 (N_4345,N_3725,N_3693);
xor U4346 (N_4346,N_2915,N_2944);
nand U4347 (N_4347,N_3256,N_3047);
or U4348 (N_4348,N_2720,N_3142);
nor U4349 (N_4349,N_2187,N_3046);
xor U4350 (N_4350,N_3685,N_3146);
nor U4351 (N_4351,N_2751,N_2716);
nor U4352 (N_4352,N_2807,N_3438);
nand U4353 (N_4353,N_2539,N_3671);
nand U4354 (N_4354,N_2721,N_3044);
nor U4355 (N_4355,N_2621,N_2284);
and U4356 (N_4356,N_2518,N_2220);
xor U4357 (N_4357,N_2934,N_3855);
xnor U4358 (N_4358,N_3936,N_3011);
and U4359 (N_4359,N_2317,N_2782);
nand U4360 (N_4360,N_2212,N_3722);
xnor U4361 (N_4361,N_3148,N_2532);
xor U4362 (N_4362,N_2493,N_3079);
nand U4363 (N_4363,N_3624,N_2630);
and U4364 (N_4364,N_3642,N_2472);
xnor U4365 (N_4365,N_3300,N_3172);
xor U4366 (N_4366,N_3648,N_2206);
and U4367 (N_4367,N_2701,N_2851);
xnor U4368 (N_4368,N_2878,N_2881);
nand U4369 (N_4369,N_3024,N_3857);
and U4370 (N_4370,N_2707,N_3995);
or U4371 (N_4371,N_3679,N_2254);
xnor U4372 (N_4372,N_3891,N_3324);
nor U4373 (N_4373,N_2557,N_3739);
or U4374 (N_4374,N_2924,N_2986);
nor U4375 (N_4375,N_3886,N_2290);
or U4376 (N_4376,N_3140,N_2880);
nor U4377 (N_4377,N_2864,N_2262);
or U4378 (N_4378,N_2787,N_2689);
xnor U4379 (N_4379,N_2148,N_2306);
nor U4380 (N_4380,N_2410,N_3981);
xnor U4381 (N_4381,N_2305,N_3295);
nand U4382 (N_4382,N_2464,N_2150);
or U4383 (N_4383,N_3453,N_2048);
xor U4384 (N_4384,N_2990,N_3913);
or U4385 (N_4385,N_3555,N_2646);
nor U4386 (N_4386,N_3501,N_3979);
and U4387 (N_4387,N_3796,N_2699);
and U4388 (N_4388,N_2360,N_3107);
nand U4389 (N_4389,N_3853,N_2170);
nand U4390 (N_4390,N_2153,N_3768);
nand U4391 (N_4391,N_2555,N_2514);
nand U4392 (N_4392,N_2653,N_3868);
xor U4393 (N_4393,N_3485,N_3253);
nor U4394 (N_4394,N_3547,N_3879);
and U4395 (N_4395,N_3903,N_2855);
or U4396 (N_4396,N_2074,N_3681);
nor U4397 (N_4397,N_2627,N_3966);
and U4398 (N_4398,N_2634,N_2729);
and U4399 (N_4399,N_3882,N_2868);
nand U4400 (N_4400,N_2327,N_2908);
or U4401 (N_4401,N_2843,N_3815);
or U4402 (N_4402,N_3175,N_2512);
nand U4403 (N_4403,N_3221,N_3279);
nand U4404 (N_4404,N_2590,N_2893);
xor U4405 (N_4405,N_3137,N_3633);
xnor U4406 (N_4406,N_3775,N_3577);
nand U4407 (N_4407,N_3086,N_2477);
xor U4408 (N_4408,N_3518,N_2182);
and U4409 (N_4409,N_3634,N_2580);
nor U4410 (N_4410,N_2914,N_3484);
nand U4411 (N_4411,N_3389,N_3861);
nand U4412 (N_4412,N_3896,N_2866);
or U4413 (N_4413,N_3834,N_2871);
and U4414 (N_4414,N_3738,N_2852);
nor U4415 (N_4415,N_2072,N_2930);
nor U4416 (N_4416,N_2264,N_2734);
nor U4417 (N_4417,N_2985,N_3786);
or U4418 (N_4418,N_2973,N_2355);
xor U4419 (N_4419,N_2560,N_2379);
and U4420 (N_4420,N_2639,N_3395);
nand U4421 (N_4421,N_2340,N_3023);
nand U4422 (N_4422,N_3451,N_2860);
xnor U4423 (N_4423,N_3065,N_3171);
nor U4424 (N_4424,N_2362,N_2324);
xnor U4425 (N_4425,N_3122,N_2554);
nor U4426 (N_4426,N_3103,N_3380);
nand U4427 (N_4427,N_3901,N_2772);
nor U4428 (N_4428,N_2083,N_2678);
nor U4429 (N_4429,N_2762,N_2334);
nor U4430 (N_4430,N_2517,N_3997);
nor U4431 (N_4431,N_3144,N_2509);
xnor U4432 (N_4432,N_2958,N_2776);
and U4433 (N_4433,N_3992,N_3523);
or U4434 (N_4434,N_2012,N_2999);
xor U4435 (N_4435,N_2954,N_3893);
and U4436 (N_4436,N_3606,N_2920);
or U4437 (N_4437,N_3691,N_3742);
nor U4438 (N_4438,N_3970,N_3596);
and U4439 (N_4439,N_2667,N_2201);
nor U4440 (N_4440,N_3374,N_2296);
xor U4441 (N_4441,N_3411,N_2917);
nand U4442 (N_4442,N_3038,N_3873);
and U4443 (N_4443,N_2259,N_3666);
nor U4444 (N_4444,N_2406,N_3059);
nor U4445 (N_4445,N_3926,N_3607);
or U4446 (N_4446,N_3652,N_3452);
nand U4447 (N_4447,N_3908,N_2794);
or U4448 (N_4448,N_2134,N_2887);
nand U4449 (N_4449,N_3764,N_3280);
and U4450 (N_4450,N_2194,N_2478);
nor U4451 (N_4451,N_3579,N_3561);
xnor U4452 (N_4452,N_3704,N_2937);
nor U4453 (N_4453,N_2690,N_3756);
and U4454 (N_4454,N_3481,N_3571);
nor U4455 (N_4455,N_3783,N_2823);
nor U4456 (N_4456,N_3301,N_3259);
nand U4457 (N_4457,N_2303,N_3433);
nand U4458 (N_4458,N_2265,N_2865);
xor U4459 (N_4459,N_3178,N_2882);
nor U4460 (N_4460,N_2530,N_2158);
or U4461 (N_4461,N_3533,N_3307);
and U4462 (N_4462,N_3566,N_3998);
nand U4463 (N_4463,N_2565,N_3660);
and U4464 (N_4464,N_3258,N_2292);
or U4465 (N_4465,N_3524,N_3580);
nand U4466 (N_4466,N_2077,N_2657);
xor U4467 (N_4467,N_3594,N_3870);
nor U4468 (N_4468,N_2078,N_3068);
and U4469 (N_4469,N_2802,N_2656);
xor U4470 (N_4470,N_2352,N_3123);
and U4471 (N_4471,N_2175,N_2779);
xnor U4472 (N_4472,N_2351,N_2923);
xnor U4473 (N_4473,N_2850,N_3472);
nor U4474 (N_4474,N_2673,N_3358);
nand U4475 (N_4475,N_2680,N_2567);
and U4476 (N_4476,N_3605,N_2323);
nand U4477 (N_4477,N_2602,N_3242);
nand U4478 (N_4478,N_3099,N_2046);
nor U4479 (N_4479,N_2405,N_3299);
or U4480 (N_4480,N_3663,N_2006);
nor U4481 (N_4481,N_3985,N_3158);
xnor U4482 (N_4482,N_3977,N_2962);
nand U4483 (N_4483,N_3718,N_2834);
or U4484 (N_4484,N_3362,N_3554);
and U4485 (N_4485,N_2550,N_3714);
nor U4486 (N_4486,N_3006,N_3031);
and U4487 (N_4487,N_2269,N_2144);
and U4488 (N_4488,N_2788,N_3650);
nand U4489 (N_4489,N_3578,N_3829);
nor U4490 (N_4490,N_3887,N_3478);
nor U4491 (N_4491,N_3792,N_3749);
xor U4492 (N_4492,N_3273,N_3708);
xnor U4493 (N_4493,N_3856,N_2235);
nand U4494 (N_4494,N_2136,N_3697);
or U4495 (N_4495,N_2651,N_2694);
nand U4496 (N_4496,N_3225,N_2020);
xnor U4497 (N_4497,N_2227,N_2620);
nor U4498 (N_4498,N_2388,N_2982);
nor U4499 (N_4499,N_3027,N_3381);
and U4500 (N_4500,N_2367,N_2469);
xnor U4501 (N_4501,N_3157,N_3960);
or U4502 (N_4502,N_3015,N_3692);
or U4503 (N_4503,N_3993,N_3517);
or U4504 (N_4504,N_2330,N_3636);
nand U4505 (N_4505,N_3228,N_3439);
nor U4506 (N_4506,N_3022,N_3417);
and U4507 (N_4507,N_3072,N_2660);
nor U4508 (N_4508,N_3257,N_2591);
nor U4509 (N_4509,N_2605,N_2638);
nand U4510 (N_4510,N_3645,N_3622);
nor U4511 (N_4511,N_3344,N_3427);
nor U4512 (N_4512,N_2118,N_3788);
and U4513 (N_4513,N_2615,N_3455);
xnor U4514 (N_4514,N_3292,N_2346);
xor U4515 (N_4515,N_3664,N_3824);
nand U4516 (N_4516,N_3640,N_2534);
or U4517 (N_4517,N_2070,N_2411);
nand U4518 (N_4518,N_3902,N_2902);
xor U4519 (N_4519,N_2308,N_2422);
nand U4520 (N_4520,N_3473,N_3061);
nor U4521 (N_4521,N_2576,N_3163);
xnor U4522 (N_4522,N_2283,N_3881);
xnor U4523 (N_4523,N_3526,N_2307);
nand U4524 (N_4524,N_2280,N_3497);
nor U4525 (N_4525,N_3201,N_3443);
or U4526 (N_4526,N_3294,N_3230);
and U4527 (N_4527,N_2950,N_2749);
nor U4528 (N_4528,N_3630,N_3653);
or U4529 (N_4529,N_3418,N_3109);
nor U4530 (N_4530,N_2203,N_2816);
xor U4531 (N_4531,N_3405,N_3799);
nand U4532 (N_4532,N_3479,N_2752);
nor U4533 (N_4533,N_3601,N_2225);
nand U4534 (N_4534,N_2025,N_3968);
or U4535 (N_4535,N_2835,N_2904);
xnor U4536 (N_4536,N_2085,N_2510);
or U4537 (N_4537,N_3436,N_2706);
nor U4538 (N_4538,N_2750,N_2049);
and U4539 (N_4539,N_2413,N_2041);
or U4540 (N_4540,N_3635,N_3111);
nor U4541 (N_4541,N_3154,N_2515);
nand U4542 (N_4542,N_2586,N_2447);
and U4543 (N_4543,N_3323,N_2396);
nor U4544 (N_4544,N_3506,N_2984);
nor U4545 (N_4545,N_2374,N_2282);
nor U4546 (N_4546,N_3041,N_2528);
xor U4547 (N_4547,N_3826,N_2633);
xnor U4548 (N_4548,N_3018,N_3235);
xnor U4549 (N_4549,N_3326,N_3852);
nor U4550 (N_4550,N_2609,N_2542);
and U4551 (N_4551,N_2427,N_3254);
or U4552 (N_4552,N_2128,N_3437);
xnor U4553 (N_4553,N_3302,N_3160);
nand U4554 (N_4554,N_2556,N_3707);
and U4555 (N_4555,N_2877,N_3546);
xor U4556 (N_4556,N_3260,N_3499);
xor U4557 (N_4557,N_3876,N_2438);
and U4558 (N_4558,N_3759,N_2824);
nor U4559 (N_4559,N_3611,N_3831);
xor U4560 (N_4560,N_2112,N_2674);
nor U4561 (N_4561,N_2623,N_3619);
nor U4562 (N_4562,N_2544,N_3677);
nand U4563 (N_4563,N_2502,N_2401);
nand U4564 (N_4564,N_2485,N_3087);
and U4565 (N_4565,N_3655,N_3335);
or U4566 (N_4566,N_3048,N_2279);
xor U4567 (N_4567,N_3058,N_3394);
nor U4568 (N_4568,N_2155,N_3773);
xor U4569 (N_4569,N_2827,N_3432);
or U4570 (N_4570,N_3818,N_3069);
nor U4571 (N_4571,N_2337,N_2520);
xor U4572 (N_4572,N_3315,N_2047);
xor U4573 (N_4573,N_2033,N_3710);
and U4574 (N_4574,N_3716,N_3706);
xor U4575 (N_4575,N_3195,N_3543);
nor U4576 (N_4576,N_2030,N_2122);
and U4577 (N_4577,N_3164,N_2470);
xor U4578 (N_4578,N_3017,N_3207);
and U4579 (N_4579,N_3174,N_2754);
and U4580 (N_4580,N_2329,N_3106);
nand U4581 (N_4581,N_3353,N_3557);
xnor U4582 (N_4582,N_3185,N_2809);
xor U4583 (N_4583,N_2730,N_3343);
and U4584 (N_4584,N_2260,N_3391);
nand U4585 (N_4585,N_2989,N_3162);
nand U4586 (N_4586,N_3776,N_3347);
or U4587 (N_4587,N_2798,N_3444);
nor U4588 (N_4588,N_3521,N_2137);
nand U4589 (N_4589,N_2131,N_2649);
nor U4590 (N_4590,N_2763,N_3133);
xor U4591 (N_4591,N_2173,N_2714);
and U4592 (N_4592,N_3293,N_3003);
xor U4593 (N_4593,N_2291,N_2350);
and U4594 (N_4594,N_2453,N_3377);
or U4595 (N_4595,N_3625,N_3434);
or U4596 (N_4596,N_3055,N_3435);
or U4597 (N_4597,N_3193,N_3943);
and U4598 (N_4598,N_2570,N_2972);
and U4599 (N_4599,N_3467,N_2107);
or U4600 (N_4600,N_2826,N_3939);
xnor U4601 (N_4601,N_3839,N_3014);
and U4602 (N_4602,N_3382,N_2945);
nor U4603 (N_4603,N_3720,N_2775);
nor U4604 (N_4604,N_3237,N_2698);
nand U4605 (N_4605,N_2833,N_3700);
xor U4606 (N_4606,N_2052,N_3544);
and U4607 (N_4607,N_3990,N_2428);
nand U4608 (N_4608,N_2825,N_3823);
xnor U4609 (N_4609,N_3540,N_3500);
nor U4610 (N_4610,N_3859,N_3265);
or U4611 (N_4611,N_3182,N_2090);
or U4612 (N_4612,N_2463,N_2738);
and U4613 (N_4613,N_3139,N_2844);
nand U4614 (N_4614,N_2744,N_2384);
xnor U4615 (N_4615,N_3229,N_2263);
nor U4616 (N_4616,N_2166,N_2703);
or U4617 (N_4617,N_2588,N_3469);
or U4618 (N_4618,N_3189,N_3153);
nor U4619 (N_4619,N_3311,N_3263);
or U4620 (N_4620,N_2578,N_3737);
and U4621 (N_4621,N_2404,N_3210);
or U4622 (N_4622,N_3964,N_2387);
nor U4623 (N_4623,N_3275,N_2066);
nand U4624 (N_4624,N_3670,N_3085);
nand U4625 (N_4625,N_2443,N_3401);
nor U4626 (N_4626,N_3614,N_2022);
nand U4627 (N_4627,N_2936,N_2642);
nand U4628 (N_4628,N_2018,N_3667);
nand U4629 (N_4629,N_3758,N_2722);
and U4630 (N_4630,N_2828,N_2386);
nand U4631 (N_4631,N_3545,N_2758);
nor U4632 (N_4632,N_3104,N_3074);
or U4633 (N_4633,N_2091,N_3609);
xnor U4634 (N_4634,N_3383,N_3317);
nor U4635 (N_4635,N_3356,N_2938);
nand U4636 (N_4636,N_3002,N_2178);
or U4637 (N_4637,N_3529,N_2248);
or U4638 (N_4638,N_3134,N_3052);
and U4639 (N_4639,N_2163,N_3368);
or U4640 (N_4640,N_2585,N_2270);
and U4641 (N_4641,N_3986,N_3110);
or U4642 (N_4642,N_3316,N_2247);
nor U4643 (N_4643,N_3213,N_2188);
nor U4644 (N_4644,N_3464,N_2038);
or U4645 (N_4645,N_2764,N_3810);
xnor U4646 (N_4646,N_2644,N_3584);
xnor U4647 (N_4647,N_3042,N_2399);
or U4648 (N_4648,N_3626,N_3155);
xnor U4649 (N_4649,N_2068,N_3396);
nand U4650 (N_4650,N_3156,N_2037);
or U4651 (N_4651,N_3699,N_3511);
nor U4652 (N_4652,N_2891,N_2380);
xnor U4653 (N_4653,N_3629,N_2370);
or U4654 (N_4654,N_3212,N_3789);
and U4655 (N_4655,N_2622,N_3920);
and U4656 (N_4656,N_3179,N_2636);
and U4657 (N_4657,N_3076,N_2094);
nor U4658 (N_4658,N_2713,N_2619);
and U4659 (N_4659,N_3800,N_2076);
xor U4660 (N_4660,N_2484,N_3795);
and U4661 (N_4661,N_2301,N_2637);
xnor U4662 (N_4662,N_3399,N_3956);
and U4663 (N_4663,N_2951,N_2885);
or U4664 (N_4664,N_2748,N_3330);
and U4665 (N_4665,N_2300,N_3276);
or U4666 (N_4666,N_2491,N_2416);
nand U4667 (N_4667,N_2412,N_2928);
nor U4668 (N_4668,N_2715,N_2785);
and U4669 (N_4669,N_2547,N_3286);
nand U4670 (N_4670,N_3589,N_3369);
and U4671 (N_4671,N_2147,N_2583);
nor U4672 (N_4672,N_3610,N_3329);
and U4673 (N_4673,N_2916,N_2302);
xor U4674 (N_4674,N_3404,N_2975);
and U4675 (N_4675,N_3291,N_3582);
and U4676 (N_4676,N_3657,N_3019);
nor U4677 (N_4677,N_3234,N_2488);
nand U4678 (N_4678,N_3628,N_2363);
xnor U4679 (N_4679,N_3837,N_2563);
xnor U4680 (N_4680,N_2858,N_3948);
xor U4681 (N_4681,N_3032,N_2217);
or U4682 (N_4682,N_2635,N_2884);
and U4683 (N_4683,N_3345,N_3145);
nand U4684 (N_4684,N_2383,N_2577);
or U4685 (N_4685,N_3885,N_3570);
nor U4686 (N_4686,N_2682,N_2473);
and U4687 (N_4687,N_3071,N_3084);
xnor U4688 (N_4688,N_3400,N_3750);
and U4689 (N_4689,N_3303,N_2255);
xnor U4690 (N_4690,N_3410,N_3649);
xnor U4691 (N_4691,N_2397,N_3514);
xnor U4692 (N_4692,N_3416,N_2065);
xor U4693 (N_4693,N_3673,N_3232);
or U4694 (N_4694,N_2896,N_3974);
and U4695 (N_4695,N_2000,N_2393);
xor U4696 (N_4696,N_2440,N_3360);
or U4697 (N_4697,N_2737,N_2496);
nand U4698 (N_4698,N_2511,N_2176);
nor U4699 (N_4699,N_2143,N_3771);
xnor U4700 (N_4700,N_3531,N_2643);
nand U4701 (N_4701,N_2870,N_2347);
xor U4702 (N_4702,N_3251,N_3842);
or U4703 (N_4703,N_2159,N_2997);
xor U4704 (N_4704,N_2319,N_2275);
nand U4705 (N_4705,N_3208,N_2433);
or U4706 (N_4706,N_2459,N_2316);
nand U4707 (N_4707,N_3062,N_3848);
or U4708 (N_4708,N_3575,N_3415);
nor U4709 (N_4709,N_3916,N_2956);
nand U4710 (N_4710,N_3367,N_3413);
and U4711 (N_4711,N_3448,N_2073);
nor U4712 (N_4712,N_3152,N_2978);
or U4713 (N_4713,N_3933,N_3371);
or U4714 (N_4714,N_2955,N_2996);
nand U4715 (N_4715,N_2811,N_3098);
and U4716 (N_4716,N_2344,N_3365);
nor U4717 (N_4717,N_2154,N_3112);
xnor U4718 (N_4718,N_3236,N_3895);
nand U4719 (N_4719,N_2007,N_2069);
and U4720 (N_4720,N_3747,N_2587);
nor U4721 (N_4721,N_3665,N_2011);
and U4722 (N_4722,N_2905,N_2594);
and U4723 (N_4723,N_2221,N_3198);
xnor U4724 (N_4724,N_2538,N_2789);
or U4725 (N_4725,N_2321,N_3696);
and U4726 (N_4726,N_2054,N_3849);
xor U4727 (N_4727,N_3583,N_2250);
nand U4728 (N_4728,N_2693,N_2700);
and U4729 (N_4729,N_3250,N_3128);
and U4730 (N_4730,N_2192,N_2475);
xnor U4731 (N_4731,N_3715,N_2436);
and U4732 (N_4732,N_2670,N_3987);
nand U4733 (N_4733,N_2727,N_3054);
xnor U4734 (N_4734,N_3732,N_2132);
and U4735 (N_4735,N_2460,N_3092);
xor U4736 (N_4736,N_2064,N_2579);
or U4737 (N_4737,N_3978,N_2652);
or U4738 (N_4738,N_3904,N_3766);
nand U4739 (N_4739,N_3505,N_2036);
or U4740 (N_4740,N_2929,N_2177);
and U4741 (N_4741,N_3919,N_2123);
and U4742 (N_4742,N_3832,N_2831);
nor U4743 (N_4743,N_3530,N_3869);
nand U4744 (N_4744,N_3844,N_2223);
nor U4745 (N_4745,N_3643,N_3246);
nor U4746 (N_4746,N_3550,N_3991);
nor U4747 (N_4747,N_3151,N_2537);
or U4748 (N_4748,N_3261,N_2272);
nor U4749 (N_4749,N_3830,N_2705);
nand U4750 (N_4750,N_2001,N_3477);
nand U4751 (N_4751,N_3595,N_3780);
xnor U4752 (N_4752,N_3519,N_2309);
and U4753 (N_4753,N_2519,N_3928);
nor U4754 (N_4754,N_3202,N_3745);
xnor U4755 (N_4755,N_3000,N_2516);
or U4756 (N_4756,N_2592,N_3366);
xnor U4757 (N_4757,N_3049,N_3712);
nand U4758 (N_4758,N_2452,N_2394);
nor U4759 (N_4759,N_2921,N_2055);
or U4760 (N_4760,N_3965,N_2553);
xor U4761 (N_4761,N_3615,N_3833);
xnor U4762 (N_4762,N_2044,N_2104);
xor U4763 (N_4763,N_3813,N_2611);
xor U4764 (N_4764,N_2836,N_2051);
and U4765 (N_4765,N_2364,N_3474);
or U4766 (N_4766,N_3113,N_3951);
nor U4767 (N_4767,N_3678,N_2288);
nand U4768 (N_4768,N_3726,N_3409);
nor U4769 (N_4769,N_2886,N_3688);
or U4770 (N_4770,N_3694,N_3961);
or U4771 (N_4771,N_2965,N_2593);
and U4772 (N_4772,N_2024,N_3502);
or U4773 (N_4773,N_2105,N_2043);
xnor U4774 (N_4774,N_3661,N_2245);
or U4775 (N_4775,N_3460,N_3496);
xnor U4776 (N_4776,N_3574,N_3108);
and U4777 (N_4777,N_3461,N_2127);
xor U4778 (N_4778,N_3423,N_2500);
xor U4779 (N_4779,N_2342,N_2445);
nand U4780 (N_4780,N_2224,N_3447);
or U4781 (N_4781,N_2862,N_2655);
and U4782 (N_4782,N_2421,N_2781);
nor U4783 (N_4783,N_3791,N_3339);
nand U4784 (N_4784,N_3214,N_2053);
or U4785 (N_4785,N_2023,N_2110);
or U4786 (N_4786,N_3278,N_3723);
and U4787 (N_4787,N_2471,N_3372);
nand U4788 (N_4788,N_2415,N_3513);
nor U4789 (N_4789,N_3147,N_3808);
or U4790 (N_4790,N_2293,N_3690);
xnor U4791 (N_4791,N_2598,N_2456);
and U4792 (N_4792,N_2425,N_2658);
nor U4793 (N_4793,N_3522,N_2017);
or U4794 (N_4794,N_3422,N_3082);
nand U4795 (N_4795,N_2804,N_2820);
xor U4796 (N_4796,N_3820,N_2692);
xor U4797 (N_4797,N_3262,N_2185);
nand U4798 (N_4798,N_3503,N_3200);
or U4799 (N_4799,N_3599,N_2755);
and U4800 (N_4800,N_3425,N_3774);
nor U4801 (N_4801,N_3025,N_2373);
nor U4802 (N_4802,N_3471,N_3504);
xnor U4803 (N_4803,N_3183,N_2160);
or U4804 (N_4804,N_3695,N_2129);
nand U4805 (N_4805,N_2869,N_2596);
or U4806 (N_4806,N_3284,N_2498);
or U4807 (N_4807,N_2541,N_2974);
or U4808 (N_4808,N_3841,N_3814);
nand U4809 (N_4809,N_2222,N_3548);
xnor U4810 (N_4810,N_2932,N_2830);
and U4811 (N_4811,N_3328,N_3012);
and U4812 (N_4812,N_3166,N_2966);
and U4813 (N_4813,N_3639,N_3173);
nor U4814 (N_4814,N_2842,N_2867);
and U4815 (N_4815,N_2684,N_2650);
nand U4816 (N_4816,N_3043,N_2719);
and U4817 (N_4817,N_3204,N_2977);
nor U4818 (N_4818,N_2709,N_3319);
nand U4819 (N_4819,N_3220,N_3150);
nand U4820 (N_4820,N_2992,N_3802);
nor U4821 (N_4821,N_2369,N_3892);
and U4822 (N_4822,N_2009,N_2109);
nand U4823 (N_4823,N_2903,N_3539);
xor U4824 (N_4824,N_2140,N_3613);
nand U4825 (N_4825,N_2450,N_2013);
xnor U4826 (N_4826,N_3285,N_2278);
xnor U4827 (N_4827,N_2529,N_3309);
or U4828 (N_4828,N_2735,N_2408);
and U4829 (N_4829,N_3114,N_2856);
or U4830 (N_4830,N_3135,N_2558);
xor U4831 (N_4831,N_3045,N_3907);
or U4832 (N_4832,N_2747,N_3953);
nor U4833 (N_4833,N_2933,N_2822);
or U4834 (N_4834,N_3760,N_2273);
nand U4835 (N_4835,N_2863,N_2668);
and U4836 (N_4836,N_3958,N_2946);
or U4837 (N_4837,N_2927,N_3445);
nand U4838 (N_4838,N_2686,N_2116);
and U4839 (N_4839,N_3412,N_2242);
nor U4840 (N_4840,N_3559,N_2063);
xnor U4841 (N_4841,N_2895,N_2015);
xor U4842 (N_4842,N_2172,N_2910);
and U4843 (N_4843,N_3591,N_2141);
nand U4844 (N_4844,N_3674,N_2797);
or U4845 (N_4845,N_2338,N_3194);
nand U4846 (N_4846,N_2628,N_2859);
nor U4847 (N_4847,N_2274,N_3332);
and U4848 (N_4848,N_3197,N_2840);
xnor U4849 (N_4849,N_2395,N_3809);
nor U4850 (N_4850,N_3562,N_2664);
and U4851 (N_4851,N_3060,N_3576);
nand U4852 (N_4852,N_3592,N_2115);
nand U4853 (N_4853,N_3930,N_3963);
and U4854 (N_4854,N_2111,N_3717);
and U4855 (N_4855,N_2853,N_2075);
xor U4856 (N_4856,N_3440,N_2239);
or U4857 (N_4857,N_3822,N_3659);
xnor U4858 (N_4858,N_2016,N_3338);
or U4859 (N_4859,N_3989,N_3136);
xor U4860 (N_4860,N_2482,N_2389);
and U4861 (N_4861,N_3604,N_3654);
nor U4862 (N_4862,N_2102,N_2616);
nor U4863 (N_4863,N_3255,N_2204);
nand U4864 (N_4864,N_3080,N_2931);
and U4865 (N_4865,N_2162,N_2332);
and U4866 (N_4866,N_2426,N_3797);
nor U4867 (N_4867,N_3268,N_2549);
or U4868 (N_4868,N_2180,N_3569);
or U4869 (N_4869,N_2474,N_2963);
and U4870 (N_4870,N_3206,N_3779);
and U4871 (N_4871,N_3211,N_2372);
nand U4872 (N_4872,N_2569,N_2361);
and U4873 (N_4873,N_2184,N_3938);
and U4874 (N_4874,N_3376,N_2559);
nand U4875 (N_4875,N_2508,N_2095);
nor U4876 (N_4876,N_3884,N_3705);
nor U4877 (N_4877,N_3141,N_2531);
and U4878 (N_4878,N_2454,N_2193);
xor U4879 (N_4879,N_2953,N_2697);
nand U4880 (N_4880,N_2595,N_2059);
or U4881 (N_4881,N_2267,N_3492);
nand U4882 (N_4882,N_2326,N_3616);
or U4883 (N_4883,N_2922,N_3911);
or U4884 (N_4884,N_3361,N_3731);
nand U4885 (N_4885,N_3168,N_3313);
xor U4886 (N_4886,N_3266,N_2872);
xnor U4887 (N_4887,N_3880,N_3130);
and U4888 (N_4888,N_3450,N_3270);
or U4889 (N_4889,N_3713,N_3656);
or U4890 (N_4890,N_3028,N_3127);
or U4891 (N_4891,N_2164,N_3729);
and U4892 (N_4892,N_3077,N_3581);
or U4893 (N_4893,N_3587,N_3397);
or U4894 (N_4894,N_3495,N_2117);
nor U4895 (N_4895,N_3534,N_2244);
or U4896 (N_4896,N_2522,N_3917);
xnor U4897 (N_4897,N_3352,N_2913);
nor U4898 (N_4898,N_3283,N_2437);
nor U4899 (N_4899,N_2256,N_3910);
or U4900 (N_4900,N_2391,N_2087);
xor U4901 (N_4901,N_3932,N_3556);
or U4902 (N_4902,N_3245,N_2533);
xnor U4903 (N_4903,N_2320,N_3118);
nand U4904 (N_4904,N_3538,N_2613);
nor U4905 (N_4905,N_2661,N_3507);
and U4906 (N_4906,N_3637,N_2742);
nand U4907 (N_4907,N_2439,N_2086);
or U4908 (N_4908,N_2442,N_2793);
xnor U4909 (N_4909,N_3950,N_3819);
nor U4910 (N_4910,N_2792,N_2562);
xor U4911 (N_4911,N_3468,N_3623);
xnor U4912 (N_4912,N_3947,N_2746);
xor U4913 (N_4913,N_2796,N_2991);
nor U4914 (N_4914,N_3406,N_3914);
nand U4915 (N_4915,N_3090,N_2901);
nand U4916 (N_4916,N_3608,N_3727);
nand U4917 (N_4917,N_2873,N_2005);
or U4918 (N_4918,N_3217,N_3281);
or U4919 (N_4919,N_2124,N_3804);
and U4920 (N_4920,N_2889,N_3787);
nand U4921 (N_4921,N_2230,N_3462);
xnor U4922 (N_4922,N_3858,N_2759);
or U4923 (N_4923,N_2733,N_3600);
and U4924 (N_4924,N_3769,N_2573);
and U4925 (N_4925,N_3420,N_3935);
xnor U4926 (N_4926,N_3322,N_2080);
or U4927 (N_4927,N_2524,N_3922);
nor U4928 (N_4928,N_3218,N_2507);
xor U4929 (N_4929,N_2418,N_3364);
or U4930 (N_4930,N_3030,N_3597);
or U4931 (N_4931,N_2597,N_3962);
nor U4932 (N_4932,N_2888,N_3115);
xnor U4933 (N_4933,N_2614,N_2979);
and U4934 (N_4934,N_2106,N_2135);
or U4935 (N_4935,N_2151,N_3465);
xnor U4936 (N_4936,N_3959,N_3297);
nor U4937 (N_4937,N_2067,N_3119);
nand U4938 (N_4938,N_3424,N_3282);
nand U4939 (N_4939,N_3355,N_2912);
nand U4940 (N_4940,N_3289,N_3620);
and U4941 (N_4941,N_3542,N_3598);
or U4942 (N_4942,N_3131,N_2521);
and U4943 (N_4943,N_2791,N_3033);
xnor U4944 (N_4944,N_3004,N_3875);
nor U4945 (N_4945,N_3314,N_2197);
or U4946 (N_4946,N_3618,N_2925);
nand U4947 (N_4947,N_3350,N_2375);
nand U4948 (N_4948,N_2268,N_2845);
nor U4949 (N_4949,N_3741,N_2741);
and U4950 (N_4950,N_2704,N_2679);
xor U4951 (N_4951,N_3379,N_3187);
nor U4952 (N_4952,N_2157,N_2959);
and U4953 (N_4953,N_2271,N_2385);
and U4954 (N_4954,N_2196,N_2125);
xor U4955 (N_4955,N_3430,N_2994);
or U4956 (N_4956,N_3020,N_3994);
nand U4957 (N_4957,N_3029,N_2050);
xnor U4958 (N_4958,N_3806,N_2207);
or U4959 (N_4959,N_2662,N_2002);
and U4960 (N_4960,N_2572,N_2216);
and U4961 (N_4961,N_3735,N_3863);
nand U4962 (N_4962,N_3184,N_3683);
nor U4963 (N_4963,N_3743,N_3305);
nor U4964 (N_4964,N_3509,N_3490);
nor U4965 (N_4965,N_2832,N_2724);
and U4966 (N_4966,N_3736,N_2457);
or U4967 (N_4967,N_3927,N_2481);
nor U4968 (N_4968,N_3672,N_2266);
xnor U4969 (N_4969,N_2947,N_3850);
xor U4970 (N_4970,N_2625,N_2082);
or U4971 (N_4971,N_3676,N_2897);
and U4972 (N_4972,N_2287,N_3845);
nand U4973 (N_4973,N_2841,N_2777);
nand U4974 (N_4974,N_3924,N_2126);
or U4975 (N_4975,N_2241,N_2669);
or U4976 (N_4976,N_3790,N_3387);
and U4977 (N_4977,N_2861,N_3095);
and U4978 (N_4978,N_3520,N_2179);
xor U4979 (N_4979,N_3247,N_3161);
nor U4980 (N_4980,N_2368,N_2718);
nand U4981 (N_4981,N_2251,N_3680);
nand U4982 (N_4982,N_2312,N_3244);
xnor U4983 (N_4983,N_2640,N_3081);
nand U4984 (N_4984,N_2119,N_2479);
xnor U4985 (N_4985,N_2056,N_3860);
and U4986 (N_4986,N_2198,N_3272);
or U4987 (N_4987,N_3341,N_3668);
or U4988 (N_4988,N_3918,N_2600);
or U4989 (N_4989,N_3698,N_3223);
xnor U4990 (N_4990,N_2328,N_2142);
xor U4991 (N_4991,N_3840,N_2725);
xnor U4992 (N_4992,N_2967,N_2909);
and U4993 (N_4993,N_2295,N_3767);
xor U4994 (N_4994,N_2961,N_3454);
nand U4995 (N_4995,N_3482,N_3442);
nor U4996 (N_4996,N_2032,N_3370);
and U4997 (N_4997,N_3177,N_2543);
nand U4998 (N_4998,N_3888,N_3753);
nand U4999 (N_4999,N_2939,N_2773);
xor U5000 (N_5000,N_3887,N_3518);
and U5001 (N_5001,N_2809,N_2871);
and U5002 (N_5002,N_2550,N_3218);
nor U5003 (N_5003,N_3706,N_2387);
or U5004 (N_5004,N_2734,N_2934);
and U5005 (N_5005,N_3899,N_2439);
and U5006 (N_5006,N_3106,N_2820);
nand U5007 (N_5007,N_2437,N_2035);
nor U5008 (N_5008,N_3635,N_2289);
nand U5009 (N_5009,N_3247,N_3099);
nor U5010 (N_5010,N_3663,N_2317);
nor U5011 (N_5011,N_2479,N_2153);
or U5012 (N_5012,N_3381,N_2231);
or U5013 (N_5013,N_2423,N_3788);
and U5014 (N_5014,N_2369,N_2472);
and U5015 (N_5015,N_3969,N_2759);
nand U5016 (N_5016,N_3188,N_2029);
and U5017 (N_5017,N_3964,N_3492);
xor U5018 (N_5018,N_2787,N_2471);
and U5019 (N_5019,N_2342,N_3224);
and U5020 (N_5020,N_2236,N_3515);
and U5021 (N_5021,N_3560,N_3382);
or U5022 (N_5022,N_2251,N_3501);
xnor U5023 (N_5023,N_3030,N_3854);
xnor U5024 (N_5024,N_3315,N_2468);
or U5025 (N_5025,N_3228,N_3443);
nor U5026 (N_5026,N_3468,N_3184);
and U5027 (N_5027,N_3001,N_3592);
or U5028 (N_5028,N_2118,N_3544);
nand U5029 (N_5029,N_2701,N_2322);
nand U5030 (N_5030,N_3167,N_2454);
xor U5031 (N_5031,N_3985,N_3897);
nand U5032 (N_5032,N_2113,N_2624);
or U5033 (N_5033,N_2030,N_2140);
xor U5034 (N_5034,N_2159,N_3373);
xor U5035 (N_5035,N_3157,N_3216);
and U5036 (N_5036,N_2595,N_3458);
or U5037 (N_5037,N_3652,N_3041);
nand U5038 (N_5038,N_2100,N_3460);
or U5039 (N_5039,N_2601,N_3491);
nand U5040 (N_5040,N_2033,N_3312);
xnor U5041 (N_5041,N_2570,N_2026);
nand U5042 (N_5042,N_2551,N_3270);
or U5043 (N_5043,N_3524,N_3239);
nand U5044 (N_5044,N_3934,N_3498);
and U5045 (N_5045,N_3498,N_3897);
and U5046 (N_5046,N_2493,N_3156);
nor U5047 (N_5047,N_3658,N_2962);
xnor U5048 (N_5048,N_2525,N_2899);
xor U5049 (N_5049,N_3221,N_2869);
or U5050 (N_5050,N_3766,N_3043);
and U5051 (N_5051,N_2503,N_3262);
or U5052 (N_5052,N_2586,N_3655);
nor U5053 (N_5053,N_2060,N_3316);
nor U5054 (N_5054,N_2112,N_3100);
nand U5055 (N_5055,N_2230,N_3152);
or U5056 (N_5056,N_3354,N_2891);
xor U5057 (N_5057,N_3347,N_3846);
or U5058 (N_5058,N_3662,N_2124);
nand U5059 (N_5059,N_2015,N_2612);
nand U5060 (N_5060,N_2703,N_3562);
or U5061 (N_5061,N_3438,N_3929);
nand U5062 (N_5062,N_3562,N_3487);
nor U5063 (N_5063,N_3941,N_3894);
xor U5064 (N_5064,N_2199,N_3228);
and U5065 (N_5065,N_2741,N_3409);
or U5066 (N_5066,N_3072,N_2103);
and U5067 (N_5067,N_3665,N_3362);
nor U5068 (N_5068,N_2182,N_2564);
nor U5069 (N_5069,N_2052,N_3157);
xor U5070 (N_5070,N_3399,N_2719);
xnor U5071 (N_5071,N_3679,N_3911);
xor U5072 (N_5072,N_2133,N_2124);
nand U5073 (N_5073,N_2233,N_3366);
xor U5074 (N_5074,N_3094,N_2418);
or U5075 (N_5075,N_2802,N_2507);
or U5076 (N_5076,N_2859,N_2007);
xnor U5077 (N_5077,N_2792,N_2787);
xnor U5078 (N_5078,N_3743,N_2295);
xor U5079 (N_5079,N_2794,N_2932);
nor U5080 (N_5080,N_2060,N_2207);
nor U5081 (N_5081,N_3334,N_2252);
or U5082 (N_5082,N_3161,N_2259);
nor U5083 (N_5083,N_2747,N_2865);
and U5084 (N_5084,N_2773,N_3912);
or U5085 (N_5085,N_3184,N_3337);
nor U5086 (N_5086,N_2116,N_2492);
xor U5087 (N_5087,N_2030,N_3854);
and U5088 (N_5088,N_3484,N_3222);
or U5089 (N_5089,N_2412,N_2179);
xnor U5090 (N_5090,N_2851,N_3211);
or U5091 (N_5091,N_3363,N_2130);
or U5092 (N_5092,N_2948,N_2302);
xnor U5093 (N_5093,N_2519,N_3002);
nor U5094 (N_5094,N_3535,N_3995);
and U5095 (N_5095,N_3714,N_3068);
nor U5096 (N_5096,N_3415,N_3296);
and U5097 (N_5097,N_3556,N_3543);
nand U5098 (N_5098,N_2187,N_2046);
and U5099 (N_5099,N_2093,N_3437);
and U5100 (N_5100,N_3600,N_3164);
and U5101 (N_5101,N_3331,N_3171);
and U5102 (N_5102,N_3547,N_3414);
nor U5103 (N_5103,N_2586,N_2565);
and U5104 (N_5104,N_2185,N_2735);
nor U5105 (N_5105,N_2772,N_2176);
nand U5106 (N_5106,N_2793,N_3234);
or U5107 (N_5107,N_3607,N_2408);
nor U5108 (N_5108,N_3461,N_2826);
or U5109 (N_5109,N_3436,N_2500);
nor U5110 (N_5110,N_3206,N_2145);
xor U5111 (N_5111,N_2176,N_2854);
xor U5112 (N_5112,N_3800,N_3455);
or U5113 (N_5113,N_3984,N_2847);
or U5114 (N_5114,N_3621,N_3464);
xor U5115 (N_5115,N_2068,N_3149);
or U5116 (N_5116,N_3136,N_3807);
nand U5117 (N_5117,N_3429,N_2703);
nor U5118 (N_5118,N_2545,N_2799);
xnor U5119 (N_5119,N_3050,N_3890);
or U5120 (N_5120,N_2172,N_2408);
nand U5121 (N_5121,N_3798,N_3377);
or U5122 (N_5122,N_3660,N_2953);
xor U5123 (N_5123,N_3037,N_3459);
nor U5124 (N_5124,N_2899,N_3502);
xor U5125 (N_5125,N_3110,N_2704);
and U5126 (N_5126,N_2371,N_3165);
nand U5127 (N_5127,N_2548,N_3695);
xor U5128 (N_5128,N_2020,N_2493);
xor U5129 (N_5129,N_3183,N_3628);
nand U5130 (N_5130,N_3593,N_2295);
xor U5131 (N_5131,N_2244,N_3981);
xor U5132 (N_5132,N_3424,N_3962);
xnor U5133 (N_5133,N_3026,N_3744);
nand U5134 (N_5134,N_2849,N_3751);
xor U5135 (N_5135,N_2543,N_3540);
xnor U5136 (N_5136,N_3641,N_3195);
nand U5137 (N_5137,N_2463,N_2314);
nand U5138 (N_5138,N_2852,N_2240);
or U5139 (N_5139,N_3569,N_3871);
and U5140 (N_5140,N_3087,N_3678);
xnor U5141 (N_5141,N_2903,N_3615);
or U5142 (N_5142,N_2259,N_3293);
nand U5143 (N_5143,N_2355,N_3871);
xor U5144 (N_5144,N_2807,N_3417);
nand U5145 (N_5145,N_3794,N_2023);
or U5146 (N_5146,N_2572,N_3463);
xor U5147 (N_5147,N_3873,N_3298);
xor U5148 (N_5148,N_2192,N_2969);
or U5149 (N_5149,N_3017,N_3498);
or U5150 (N_5150,N_2706,N_2531);
and U5151 (N_5151,N_2577,N_2366);
nand U5152 (N_5152,N_3480,N_3292);
and U5153 (N_5153,N_2077,N_3583);
xor U5154 (N_5154,N_3389,N_3919);
xor U5155 (N_5155,N_3193,N_3297);
or U5156 (N_5156,N_3827,N_2369);
nor U5157 (N_5157,N_2982,N_2889);
nand U5158 (N_5158,N_2402,N_3690);
or U5159 (N_5159,N_3436,N_2319);
xnor U5160 (N_5160,N_2471,N_2598);
xor U5161 (N_5161,N_3728,N_3811);
xnor U5162 (N_5162,N_3487,N_2952);
nand U5163 (N_5163,N_2978,N_2830);
or U5164 (N_5164,N_2116,N_2581);
xnor U5165 (N_5165,N_2225,N_2936);
nor U5166 (N_5166,N_3971,N_3548);
xnor U5167 (N_5167,N_2553,N_2668);
nand U5168 (N_5168,N_3227,N_2591);
nor U5169 (N_5169,N_2842,N_3487);
nand U5170 (N_5170,N_2877,N_3818);
nand U5171 (N_5171,N_2539,N_3818);
nor U5172 (N_5172,N_3523,N_2540);
and U5173 (N_5173,N_2755,N_2032);
and U5174 (N_5174,N_2407,N_3725);
nand U5175 (N_5175,N_2736,N_2207);
nand U5176 (N_5176,N_2930,N_3695);
and U5177 (N_5177,N_3137,N_3718);
nand U5178 (N_5178,N_2667,N_2878);
nor U5179 (N_5179,N_2421,N_2101);
and U5180 (N_5180,N_2011,N_3021);
and U5181 (N_5181,N_2361,N_3035);
nor U5182 (N_5182,N_2422,N_3147);
and U5183 (N_5183,N_2083,N_3629);
nand U5184 (N_5184,N_3631,N_2425);
and U5185 (N_5185,N_2105,N_2278);
nor U5186 (N_5186,N_2603,N_3508);
xnor U5187 (N_5187,N_3896,N_3405);
or U5188 (N_5188,N_3623,N_3072);
or U5189 (N_5189,N_3206,N_2144);
nand U5190 (N_5190,N_2220,N_3711);
xnor U5191 (N_5191,N_2467,N_2765);
nor U5192 (N_5192,N_3546,N_3517);
and U5193 (N_5193,N_3025,N_2179);
and U5194 (N_5194,N_2661,N_3522);
and U5195 (N_5195,N_2682,N_3662);
or U5196 (N_5196,N_3210,N_2836);
nor U5197 (N_5197,N_2755,N_2175);
nand U5198 (N_5198,N_3902,N_2922);
or U5199 (N_5199,N_3883,N_3553);
xnor U5200 (N_5200,N_3104,N_2833);
xor U5201 (N_5201,N_2227,N_3265);
nor U5202 (N_5202,N_2267,N_2184);
nand U5203 (N_5203,N_2109,N_3403);
and U5204 (N_5204,N_3211,N_2509);
xor U5205 (N_5205,N_2191,N_2555);
xor U5206 (N_5206,N_2804,N_2754);
nor U5207 (N_5207,N_3013,N_3435);
nor U5208 (N_5208,N_2031,N_3261);
or U5209 (N_5209,N_3098,N_3865);
or U5210 (N_5210,N_3617,N_2410);
and U5211 (N_5211,N_3535,N_3912);
nor U5212 (N_5212,N_2603,N_2064);
nor U5213 (N_5213,N_2698,N_2603);
nor U5214 (N_5214,N_2212,N_2817);
nand U5215 (N_5215,N_3881,N_3836);
nor U5216 (N_5216,N_2050,N_2780);
nand U5217 (N_5217,N_3421,N_2307);
and U5218 (N_5218,N_2027,N_2897);
or U5219 (N_5219,N_2848,N_3736);
and U5220 (N_5220,N_2202,N_3670);
or U5221 (N_5221,N_3184,N_2998);
or U5222 (N_5222,N_2876,N_3238);
or U5223 (N_5223,N_3932,N_3869);
and U5224 (N_5224,N_3407,N_3913);
nand U5225 (N_5225,N_3780,N_2992);
xor U5226 (N_5226,N_2235,N_2148);
xnor U5227 (N_5227,N_3045,N_2091);
or U5228 (N_5228,N_2592,N_3705);
xnor U5229 (N_5229,N_2708,N_3588);
nand U5230 (N_5230,N_3211,N_2673);
nor U5231 (N_5231,N_3840,N_2881);
nor U5232 (N_5232,N_3720,N_2002);
and U5233 (N_5233,N_2928,N_3615);
nor U5234 (N_5234,N_2638,N_3641);
xor U5235 (N_5235,N_3902,N_2464);
xor U5236 (N_5236,N_2435,N_2656);
and U5237 (N_5237,N_3393,N_3699);
xor U5238 (N_5238,N_2994,N_3760);
nor U5239 (N_5239,N_2716,N_3556);
xnor U5240 (N_5240,N_2626,N_3888);
nand U5241 (N_5241,N_3694,N_3890);
xnor U5242 (N_5242,N_2281,N_3628);
nand U5243 (N_5243,N_2562,N_2983);
and U5244 (N_5244,N_3623,N_3286);
nor U5245 (N_5245,N_3735,N_2029);
xor U5246 (N_5246,N_3521,N_3240);
nand U5247 (N_5247,N_3574,N_2704);
nor U5248 (N_5248,N_3887,N_3857);
xor U5249 (N_5249,N_3890,N_3983);
nor U5250 (N_5250,N_2615,N_2583);
nand U5251 (N_5251,N_2597,N_3611);
xnor U5252 (N_5252,N_3179,N_3819);
nor U5253 (N_5253,N_3308,N_3352);
or U5254 (N_5254,N_2466,N_3828);
nor U5255 (N_5255,N_2130,N_3554);
xor U5256 (N_5256,N_2220,N_2487);
or U5257 (N_5257,N_2761,N_2623);
xnor U5258 (N_5258,N_3819,N_3515);
nor U5259 (N_5259,N_3840,N_2960);
nor U5260 (N_5260,N_2978,N_3428);
nand U5261 (N_5261,N_2767,N_3985);
xor U5262 (N_5262,N_2906,N_2317);
nor U5263 (N_5263,N_3561,N_2926);
xnor U5264 (N_5264,N_3661,N_3382);
and U5265 (N_5265,N_2742,N_3195);
xor U5266 (N_5266,N_2556,N_2067);
or U5267 (N_5267,N_3562,N_3371);
or U5268 (N_5268,N_3209,N_2374);
nor U5269 (N_5269,N_2779,N_3767);
and U5270 (N_5270,N_2566,N_3099);
and U5271 (N_5271,N_2421,N_2471);
or U5272 (N_5272,N_3264,N_2148);
xor U5273 (N_5273,N_3559,N_2621);
nand U5274 (N_5274,N_3523,N_2541);
nor U5275 (N_5275,N_2975,N_3944);
and U5276 (N_5276,N_3995,N_2032);
nor U5277 (N_5277,N_2021,N_3340);
nand U5278 (N_5278,N_3101,N_2196);
xor U5279 (N_5279,N_3948,N_3844);
nor U5280 (N_5280,N_3835,N_3987);
nor U5281 (N_5281,N_3719,N_2322);
or U5282 (N_5282,N_3257,N_3738);
nand U5283 (N_5283,N_2644,N_3951);
or U5284 (N_5284,N_3618,N_2271);
xor U5285 (N_5285,N_3495,N_2955);
nor U5286 (N_5286,N_3877,N_2964);
xor U5287 (N_5287,N_2902,N_3303);
or U5288 (N_5288,N_3812,N_2396);
or U5289 (N_5289,N_2656,N_2898);
and U5290 (N_5290,N_2051,N_2492);
and U5291 (N_5291,N_2606,N_3481);
and U5292 (N_5292,N_3613,N_3715);
xor U5293 (N_5293,N_2131,N_3803);
xor U5294 (N_5294,N_2113,N_2536);
and U5295 (N_5295,N_3725,N_2454);
and U5296 (N_5296,N_2760,N_2543);
or U5297 (N_5297,N_2650,N_2539);
nand U5298 (N_5298,N_3090,N_3303);
or U5299 (N_5299,N_3099,N_3075);
xor U5300 (N_5300,N_2529,N_3283);
and U5301 (N_5301,N_3283,N_3860);
xnor U5302 (N_5302,N_2912,N_2895);
xor U5303 (N_5303,N_2801,N_2406);
nor U5304 (N_5304,N_2566,N_3915);
nand U5305 (N_5305,N_2797,N_2197);
xor U5306 (N_5306,N_2064,N_3124);
nand U5307 (N_5307,N_2080,N_2938);
nand U5308 (N_5308,N_3231,N_2380);
nand U5309 (N_5309,N_2515,N_2569);
or U5310 (N_5310,N_2552,N_2195);
or U5311 (N_5311,N_2106,N_3917);
xnor U5312 (N_5312,N_2574,N_2486);
nand U5313 (N_5313,N_3925,N_3891);
xnor U5314 (N_5314,N_2621,N_3035);
and U5315 (N_5315,N_3200,N_3259);
xnor U5316 (N_5316,N_2547,N_2935);
nor U5317 (N_5317,N_2054,N_3757);
nand U5318 (N_5318,N_3474,N_2633);
xnor U5319 (N_5319,N_3819,N_2831);
xor U5320 (N_5320,N_2462,N_2984);
nand U5321 (N_5321,N_3475,N_3045);
and U5322 (N_5322,N_2521,N_3351);
and U5323 (N_5323,N_2616,N_2066);
xor U5324 (N_5324,N_3542,N_2302);
or U5325 (N_5325,N_3555,N_3504);
nand U5326 (N_5326,N_3377,N_2816);
or U5327 (N_5327,N_3899,N_2788);
nor U5328 (N_5328,N_3761,N_2933);
and U5329 (N_5329,N_3690,N_2299);
xnor U5330 (N_5330,N_3351,N_2799);
and U5331 (N_5331,N_2702,N_2020);
and U5332 (N_5332,N_2706,N_3251);
xnor U5333 (N_5333,N_3958,N_2980);
or U5334 (N_5334,N_3939,N_2728);
or U5335 (N_5335,N_2733,N_2100);
and U5336 (N_5336,N_3334,N_3554);
xor U5337 (N_5337,N_3136,N_2135);
xnor U5338 (N_5338,N_2190,N_2099);
or U5339 (N_5339,N_2876,N_2877);
nor U5340 (N_5340,N_2928,N_3156);
xnor U5341 (N_5341,N_2047,N_2421);
nand U5342 (N_5342,N_2978,N_2226);
or U5343 (N_5343,N_2301,N_2794);
nor U5344 (N_5344,N_3973,N_3630);
nand U5345 (N_5345,N_3295,N_3903);
xor U5346 (N_5346,N_2216,N_2068);
nand U5347 (N_5347,N_3122,N_2876);
xnor U5348 (N_5348,N_2573,N_3832);
xor U5349 (N_5349,N_2249,N_2702);
xor U5350 (N_5350,N_3057,N_3638);
xor U5351 (N_5351,N_3525,N_3144);
xnor U5352 (N_5352,N_2903,N_2846);
xnor U5353 (N_5353,N_3507,N_3289);
or U5354 (N_5354,N_2735,N_2941);
or U5355 (N_5355,N_3697,N_2149);
nor U5356 (N_5356,N_3890,N_3042);
nand U5357 (N_5357,N_3310,N_3453);
xnor U5358 (N_5358,N_3626,N_3002);
or U5359 (N_5359,N_3074,N_2646);
nand U5360 (N_5360,N_3432,N_2126);
or U5361 (N_5361,N_2545,N_2007);
and U5362 (N_5362,N_2887,N_3541);
nand U5363 (N_5363,N_3879,N_2839);
nor U5364 (N_5364,N_2404,N_2501);
nor U5365 (N_5365,N_3762,N_2658);
nor U5366 (N_5366,N_3284,N_3100);
or U5367 (N_5367,N_3166,N_3513);
xor U5368 (N_5368,N_2931,N_2526);
xor U5369 (N_5369,N_3165,N_3241);
nand U5370 (N_5370,N_3933,N_2292);
xor U5371 (N_5371,N_3262,N_3790);
nand U5372 (N_5372,N_3725,N_2175);
or U5373 (N_5373,N_3697,N_3674);
xor U5374 (N_5374,N_2936,N_3617);
nor U5375 (N_5375,N_3415,N_2942);
nand U5376 (N_5376,N_2449,N_2931);
xnor U5377 (N_5377,N_2968,N_3633);
nor U5378 (N_5378,N_3605,N_3513);
or U5379 (N_5379,N_2407,N_3026);
and U5380 (N_5380,N_3054,N_2427);
nand U5381 (N_5381,N_3546,N_2450);
or U5382 (N_5382,N_2482,N_3770);
xnor U5383 (N_5383,N_2083,N_3426);
or U5384 (N_5384,N_2492,N_2771);
and U5385 (N_5385,N_2807,N_3364);
nor U5386 (N_5386,N_3057,N_2362);
or U5387 (N_5387,N_3883,N_3151);
and U5388 (N_5388,N_3749,N_3480);
nand U5389 (N_5389,N_3991,N_3966);
and U5390 (N_5390,N_3358,N_2287);
nor U5391 (N_5391,N_2881,N_3645);
or U5392 (N_5392,N_2554,N_3229);
nor U5393 (N_5393,N_3177,N_3858);
or U5394 (N_5394,N_3548,N_3704);
or U5395 (N_5395,N_2552,N_2422);
nand U5396 (N_5396,N_3079,N_2890);
xnor U5397 (N_5397,N_3631,N_3725);
and U5398 (N_5398,N_2852,N_2233);
nand U5399 (N_5399,N_2203,N_3729);
or U5400 (N_5400,N_2062,N_3446);
and U5401 (N_5401,N_2833,N_2280);
or U5402 (N_5402,N_3572,N_3311);
nand U5403 (N_5403,N_3490,N_2257);
nor U5404 (N_5404,N_3254,N_3302);
nor U5405 (N_5405,N_3659,N_2635);
and U5406 (N_5406,N_3880,N_2887);
and U5407 (N_5407,N_2000,N_3504);
or U5408 (N_5408,N_2995,N_2536);
nand U5409 (N_5409,N_3928,N_3835);
or U5410 (N_5410,N_3711,N_3257);
or U5411 (N_5411,N_3276,N_3159);
or U5412 (N_5412,N_3008,N_2320);
or U5413 (N_5413,N_3401,N_2450);
xnor U5414 (N_5414,N_3297,N_3102);
and U5415 (N_5415,N_3375,N_3522);
and U5416 (N_5416,N_3514,N_3146);
xor U5417 (N_5417,N_3136,N_2906);
nor U5418 (N_5418,N_3986,N_3048);
nand U5419 (N_5419,N_2875,N_3869);
or U5420 (N_5420,N_2422,N_2570);
nor U5421 (N_5421,N_2582,N_3111);
nor U5422 (N_5422,N_3521,N_2651);
and U5423 (N_5423,N_3927,N_2975);
nor U5424 (N_5424,N_2219,N_3643);
or U5425 (N_5425,N_2776,N_2426);
nor U5426 (N_5426,N_3447,N_2338);
or U5427 (N_5427,N_3712,N_2447);
xor U5428 (N_5428,N_2948,N_3143);
nor U5429 (N_5429,N_3888,N_2414);
nand U5430 (N_5430,N_2980,N_2533);
nand U5431 (N_5431,N_3062,N_3169);
nor U5432 (N_5432,N_3715,N_3060);
and U5433 (N_5433,N_3268,N_2974);
nor U5434 (N_5434,N_2191,N_2927);
or U5435 (N_5435,N_2716,N_3545);
nor U5436 (N_5436,N_2057,N_2325);
nor U5437 (N_5437,N_2792,N_2830);
and U5438 (N_5438,N_2181,N_3410);
nand U5439 (N_5439,N_3662,N_3866);
xor U5440 (N_5440,N_2461,N_2334);
nand U5441 (N_5441,N_3565,N_3739);
nor U5442 (N_5442,N_2016,N_2706);
nand U5443 (N_5443,N_3813,N_2756);
and U5444 (N_5444,N_2826,N_3022);
and U5445 (N_5445,N_3959,N_2013);
xor U5446 (N_5446,N_3859,N_2723);
or U5447 (N_5447,N_3424,N_2121);
nand U5448 (N_5448,N_2286,N_3434);
nand U5449 (N_5449,N_3419,N_2885);
nor U5450 (N_5450,N_2256,N_2269);
or U5451 (N_5451,N_2133,N_2114);
xnor U5452 (N_5452,N_2235,N_2545);
nand U5453 (N_5453,N_3972,N_3268);
and U5454 (N_5454,N_3533,N_3914);
nor U5455 (N_5455,N_2645,N_2166);
nand U5456 (N_5456,N_2175,N_3048);
nand U5457 (N_5457,N_2295,N_2065);
nor U5458 (N_5458,N_2138,N_2602);
and U5459 (N_5459,N_2531,N_3227);
nand U5460 (N_5460,N_3938,N_2643);
nor U5461 (N_5461,N_2453,N_2435);
xnor U5462 (N_5462,N_2277,N_3430);
nand U5463 (N_5463,N_3244,N_2400);
nor U5464 (N_5464,N_3417,N_3510);
nor U5465 (N_5465,N_3580,N_3709);
nor U5466 (N_5466,N_2779,N_3243);
nor U5467 (N_5467,N_2739,N_3665);
and U5468 (N_5468,N_3061,N_3949);
xnor U5469 (N_5469,N_2415,N_2890);
nor U5470 (N_5470,N_2120,N_2942);
xor U5471 (N_5471,N_2761,N_2269);
xnor U5472 (N_5472,N_3748,N_3479);
nor U5473 (N_5473,N_2051,N_3858);
xnor U5474 (N_5474,N_2636,N_2548);
and U5475 (N_5475,N_2597,N_2123);
xnor U5476 (N_5476,N_2889,N_3197);
xor U5477 (N_5477,N_3236,N_2916);
and U5478 (N_5478,N_3846,N_2628);
or U5479 (N_5479,N_2629,N_2572);
nor U5480 (N_5480,N_2112,N_3389);
xor U5481 (N_5481,N_2331,N_2143);
xor U5482 (N_5482,N_3953,N_2244);
xor U5483 (N_5483,N_2552,N_2699);
xor U5484 (N_5484,N_2250,N_3919);
nand U5485 (N_5485,N_3766,N_3516);
nand U5486 (N_5486,N_3374,N_3545);
xnor U5487 (N_5487,N_2635,N_2764);
nand U5488 (N_5488,N_2026,N_3968);
nand U5489 (N_5489,N_2554,N_2245);
and U5490 (N_5490,N_3156,N_3829);
nor U5491 (N_5491,N_3501,N_2648);
nand U5492 (N_5492,N_2075,N_2298);
xor U5493 (N_5493,N_3283,N_2265);
or U5494 (N_5494,N_2094,N_2859);
xor U5495 (N_5495,N_2548,N_2376);
and U5496 (N_5496,N_2459,N_3660);
nor U5497 (N_5497,N_2993,N_3152);
and U5498 (N_5498,N_3965,N_2747);
xor U5499 (N_5499,N_3157,N_2847);
or U5500 (N_5500,N_3337,N_2353);
xor U5501 (N_5501,N_2047,N_2564);
or U5502 (N_5502,N_3277,N_2807);
and U5503 (N_5503,N_3417,N_3095);
xor U5504 (N_5504,N_2490,N_3295);
nor U5505 (N_5505,N_2126,N_3540);
and U5506 (N_5506,N_3994,N_2770);
nand U5507 (N_5507,N_2048,N_3087);
or U5508 (N_5508,N_3570,N_2635);
xnor U5509 (N_5509,N_3408,N_2489);
xor U5510 (N_5510,N_2446,N_2019);
and U5511 (N_5511,N_3031,N_2048);
nor U5512 (N_5512,N_3769,N_3568);
xor U5513 (N_5513,N_3436,N_2328);
xnor U5514 (N_5514,N_3181,N_3160);
nand U5515 (N_5515,N_3092,N_2915);
nand U5516 (N_5516,N_2835,N_3541);
or U5517 (N_5517,N_3634,N_3014);
and U5518 (N_5518,N_2991,N_3947);
or U5519 (N_5519,N_2277,N_3461);
or U5520 (N_5520,N_3832,N_3220);
and U5521 (N_5521,N_2497,N_3205);
and U5522 (N_5522,N_2255,N_2871);
nor U5523 (N_5523,N_3201,N_3920);
xor U5524 (N_5524,N_3652,N_3396);
or U5525 (N_5525,N_2825,N_2769);
nor U5526 (N_5526,N_3116,N_3811);
nand U5527 (N_5527,N_3235,N_2467);
and U5528 (N_5528,N_2716,N_2326);
xnor U5529 (N_5529,N_2972,N_3960);
nor U5530 (N_5530,N_2237,N_3844);
or U5531 (N_5531,N_2664,N_3434);
or U5532 (N_5532,N_3893,N_2481);
or U5533 (N_5533,N_2635,N_3852);
xnor U5534 (N_5534,N_2090,N_3574);
nor U5535 (N_5535,N_3902,N_3363);
xnor U5536 (N_5536,N_2349,N_2850);
nor U5537 (N_5537,N_3572,N_3512);
xor U5538 (N_5538,N_3880,N_2002);
nand U5539 (N_5539,N_2497,N_3638);
and U5540 (N_5540,N_3265,N_2484);
and U5541 (N_5541,N_3260,N_2129);
nand U5542 (N_5542,N_3246,N_2382);
or U5543 (N_5543,N_2936,N_3698);
and U5544 (N_5544,N_3679,N_2803);
nand U5545 (N_5545,N_2607,N_2223);
xor U5546 (N_5546,N_3007,N_3201);
xor U5547 (N_5547,N_2024,N_3542);
xnor U5548 (N_5548,N_3811,N_2125);
and U5549 (N_5549,N_3170,N_2994);
xnor U5550 (N_5550,N_3447,N_3802);
and U5551 (N_5551,N_2714,N_3473);
or U5552 (N_5552,N_3616,N_3795);
or U5553 (N_5553,N_2210,N_3220);
and U5554 (N_5554,N_3344,N_2041);
xnor U5555 (N_5555,N_3461,N_2317);
nor U5556 (N_5556,N_3600,N_2153);
nor U5557 (N_5557,N_2053,N_2216);
nand U5558 (N_5558,N_3006,N_2736);
or U5559 (N_5559,N_2833,N_3106);
and U5560 (N_5560,N_3620,N_3907);
and U5561 (N_5561,N_2093,N_2353);
and U5562 (N_5562,N_3714,N_3967);
or U5563 (N_5563,N_3835,N_2029);
nand U5564 (N_5564,N_3564,N_3843);
nor U5565 (N_5565,N_2152,N_2194);
nand U5566 (N_5566,N_2677,N_2382);
and U5567 (N_5567,N_2372,N_2336);
nor U5568 (N_5568,N_2607,N_2457);
or U5569 (N_5569,N_2914,N_2534);
and U5570 (N_5570,N_3686,N_2410);
and U5571 (N_5571,N_3062,N_2384);
xor U5572 (N_5572,N_3426,N_2357);
nand U5573 (N_5573,N_3139,N_3051);
or U5574 (N_5574,N_2543,N_3357);
nor U5575 (N_5575,N_2303,N_2994);
or U5576 (N_5576,N_2920,N_3727);
or U5577 (N_5577,N_2560,N_3257);
or U5578 (N_5578,N_3343,N_3823);
nor U5579 (N_5579,N_3224,N_2688);
or U5580 (N_5580,N_2996,N_2121);
xnor U5581 (N_5581,N_2636,N_3566);
and U5582 (N_5582,N_2813,N_3165);
or U5583 (N_5583,N_2940,N_3859);
nor U5584 (N_5584,N_3429,N_2925);
nand U5585 (N_5585,N_3839,N_2828);
nand U5586 (N_5586,N_2870,N_2333);
nand U5587 (N_5587,N_2655,N_3547);
or U5588 (N_5588,N_3884,N_2465);
nand U5589 (N_5589,N_2236,N_2946);
or U5590 (N_5590,N_3283,N_2745);
and U5591 (N_5591,N_3868,N_3902);
nor U5592 (N_5592,N_3785,N_3082);
xor U5593 (N_5593,N_3979,N_2693);
or U5594 (N_5594,N_3970,N_2858);
xnor U5595 (N_5595,N_2777,N_2786);
and U5596 (N_5596,N_2167,N_3936);
xor U5597 (N_5597,N_3571,N_3769);
xnor U5598 (N_5598,N_2005,N_3424);
or U5599 (N_5599,N_2328,N_3504);
xnor U5600 (N_5600,N_2860,N_3900);
or U5601 (N_5601,N_3398,N_3904);
or U5602 (N_5602,N_3764,N_2926);
nor U5603 (N_5603,N_3845,N_2548);
nor U5604 (N_5604,N_3857,N_2368);
xnor U5605 (N_5605,N_2885,N_3488);
nand U5606 (N_5606,N_3288,N_2370);
or U5607 (N_5607,N_2275,N_3940);
nand U5608 (N_5608,N_2643,N_3627);
or U5609 (N_5609,N_2288,N_3048);
nor U5610 (N_5610,N_2790,N_2312);
xor U5611 (N_5611,N_3729,N_3159);
nor U5612 (N_5612,N_3566,N_3521);
nand U5613 (N_5613,N_2707,N_2440);
nand U5614 (N_5614,N_2735,N_2203);
nor U5615 (N_5615,N_3894,N_3920);
nor U5616 (N_5616,N_3486,N_3447);
xnor U5617 (N_5617,N_3716,N_3762);
nand U5618 (N_5618,N_3699,N_2519);
and U5619 (N_5619,N_2472,N_2202);
nor U5620 (N_5620,N_2052,N_2967);
and U5621 (N_5621,N_3792,N_2418);
xor U5622 (N_5622,N_3543,N_2848);
or U5623 (N_5623,N_2995,N_2297);
or U5624 (N_5624,N_3888,N_3835);
nand U5625 (N_5625,N_2894,N_2796);
and U5626 (N_5626,N_3017,N_2589);
and U5627 (N_5627,N_3616,N_3598);
nand U5628 (N_5628,N_3634,N_3464);
and U5629 (N_5629,N_2828,N_3371);
or U5630 (N_5630,N_3893,N_2122);
and U5631 (N_5631,N_3122,N_3286);
xnor U5632 (N_5632,N_3107,N_3241);
nor U5633 (N_5633,N_2760,N_3603);
xor U5634 (N_5634,N_2106,N_3783);
and U5635 (N_5635,N_3867,N_3064);
or U5636 (N_5636,N_2442,N_2183);
xor U5637 (N_5637,N_2668,N_3854);
nand U5638 (N_5638,N_2791,N_2640);
nand U5639 (N_5639,N_2215,N_2270);
or U5640 (N_5640,N_2962,N_2466);
nand U5641 (N_5641,N_2717,N_2951);
xnor U5642 (N_5642,N_3034,N_3987);
and U5643 (N_5643,N_3385,N_3573);
or U5644 (N_5644,N_2944,N_2922);
nand U5645 (N_5645,N_3320,N_3731);
and U5646 (N_5646,N_3907,N_2374);
or U5647 (N_5647,N_3894,N_3090);
xnor U5648 (N_5648,N_3770,N_3829);
xnor U5649 (N_5649,N_2931,N_3456);
and U5650 (N_5650,N_3016,N_3228);
xnor U5651 (N_5651,N_2945,N_3708);
nand U5652 (N_5652,N_3161,N_2047);
and U5653 (N_5653,N_3710,N_2994);
xnor U5654 (N_5654,N_2982,N_2855);
nor U5655 (N_5655,N_2446,N_3437);
nand U5656 (N_5656,N_2468,N_2701);
nand U5657 (N_5657,N_3860,N_3091);
xnor U5658 (N_5658,N_2445,N_2300);
and U5659 (N_5659,N_3223,N_2584);
xnor U5660 (N_5660,N_3408,N_3244);
nand U5661 (N_5661,N_3144,N_3893);
nor U5662 (N_5662,N_2906,N_2408);
nand U5663 (N_5663,N_2773,N_2985);
or U5664 (N_5664,N_3884,N_3820);
xor U5665 (N_5665,N_3462,N_2621);
xor U5666 (N_5666,N_3056,N_3069);
nand U5667 (N_5667,N_3778,N_3377);
xnor U5668 (N_5668,N_3485,N_2769);
nand U5669 (N_5669,N_3281,N_2369);
and U5670 (N_5670,N_2218,N_3378);
nor U5671 (N_5671,N_2190,N_2536);
xnor U5672 (N_5672,N_2988,N_2948);
nand U5673 (N_5673,N_2782,N_2233);
nand U5674 (N_5674,N_2289,N_3292);
xnor U5675 (N_5675,N_2399,N_3976);
nor U5676 (N_5676,N_3918,N_2058);
and U5677 (N_5677,N_3121,N_3932);
and U5678 (N_5678,N_2555,N_3083);
or U5679 (N_5679,N_3860,N_3046);
and U5680 (N_5680,N_2223,N_3038);
nor U5681 (N_5681,N_2238,N_2057);
xor U5682 (N_5682,N_2529,N_3311);
or U5683 (N_5683,N_3359,N_2538);
xor U5684 (N_5684,N_3531,N_2414);
or U5685 (N_5685,N_2799,N_2667);
xor U5686 (N_5686,N_3171,N_2857);
or U5687 (N_5687,N_2494,N_3978);
and U5688 (N_5688,N_2077,N_2694);
xnor U5689 (N_5689,N_2519,N_3759);
or U5690 (N_5690,N_3212,N_2850);
and U5691 (N_5691,N_2114,N_3066);
or U5692 (N_5692,N_3849,N_3993);
xnor U5693 (N_5693,N_2302,N_3681);
or U5694 (N_5694,N_2541,N_2824);
xor U5695 (N_5695,N_2980,N_3974);
and U5696 (N_5696,N_3182,N_2896);
or U5697 (N_5697,N_2493,N_2356);
nand U5698 (N_5698,N_3505,N_2414);
nor U5699 (N_5699,N_2933,N_2258);
xor U5700 (N_5700,N_2919,N_3731);
nand U5701 (N_5701,N_3355,N_2457);
nand U5702 (N_5702,N_2366,N_3962);
and U5703 (N_5703,N_2121,N_3207);
xor U5704 (N_5704,N_3750,N_2400);
nand U5705 (N_5705,N_2676,N_3263);
and U5706 (N_5706,N_3817,N_2507);
and U5707 (N_5707,N_3423,N_3046);
nand U5708 (N_5708,N_3648,N_3177);
nand U5709 (N_5709,N_2983,N_3345);
or U5710 (N_5710,N_3428,N_2383);
nor U5711 (N_5711,N_2600,N_2812);
or U5712 (N_5712,N_2437,N_2280);
xnor U5713 (N_5713,N_2064,N_3329);
xnor U5714 (N_5714,N_2829,N_3324);
or U5715 (N_5715,N_2728,N_2968);
nor U5716 (N_5716,N_2166,N_2735);
nor U5717 (N_5717,N_2904,N_3429);
xnor U5718 (N_5718,N_2531,N_2493);
nor U5719 (N_5719,N_2663,N_3417);
xor U5720 (N_5720,N_2344,N_3847);
or U5721 (N_5721,N_2915,N_2429);
nor U5722 (N_5722,N_2189,N_2264);
or U5723 (N_5723,N_2150,N_2479);
or U5724 (N_5724,N_2922,N_2897);
nor U5725 (N_5725,N_2000,N_3030);
nor U5726 (N_5726,N_3078,N_2474);
nor U5727 (N_5727,N_3409,N_2579);
nor U5728 (N_5728,N_2488,N_2128);
and U5729 (N_5729,N_3223,N_3020);
nor U5730 (N_5730,N_3300,N_2374);
nor U5731 (N_5731,N_2275,N_2001);
and U5732 (N_5732,N_2217,N_2456);
nand U5733 (N_5733,N_2595,N_3119);
xnor U5734 (N_5734,N_2630,N_3419);
and U5735 (N_5735,N_3633,N_2319);
nor U5736 (N_5736,N_3883,N_3541);
xnor U5737 (N_5737,N_2362,N_3457);
and U5738 (N_5738,N_2425,N_3394);
or U5739 (N_5739,N_3314,N_2408);
xnor U5740 (N_5740,N_2610,N_2887);
xor U5741 (N_5741,N_2011,N_2626);
and U5742 (N_5742,N_3360,N_3141);
nor U5743 (N_5743,N_3222,N_2687);
xor U5744 (N_5744,N_3939,N_3131);
and U5745 (N_5745,N_3714,N_2145);
nor U5746 (N_5746,N_3943,N_2386);
and U5747 (N_5747,N_3155,N_2446);
xnor U5748 (N_5748,N_2359,N_2642);
nand U5749 (N_5749,N_2799,N_2116);
nor U5750 (N_5750,N_2888,N_2229);
nor U5751 (N_5751,N_3162,N_3506);
xnor U5752 (N_5752,N_2376,N_3974);
xnor U5753 (N_5753,N_3064,N_2023);
nor U5754 (N_5754,N_3609,N_2553);
nand U5755 (N_5755,N_3203,N_2744);
and U5756 (N_5756,N_2434,N_2501);
nor U5757 (N_5757,N_2792,N_3206);
and U5758 (N_5758,N_3492,N_3285);
xor U5759 (N_5759,N_3283,N_2223);
nor U5760 (N_5760,N_3011,N_2619);
nor U5761 (N_5761,N_3037,N_3373);
and U5762 (N_5762,N_3744,N_3007);
or U5763 (N_5763,N_3484,N_3365);
xnor U5764 (N_5764,N_3191,N_2203);
nand U5765 (N_5765,N_3592,N_3732);
and U5766 (N_5766,N_3344,N_2750);
nor U5767 (N_5767,N_2419,N_2527);
nor U5768 (N_5768,N_2485,N_3571);
nor U5769 (N_5769,N_2201,N_3480);
nor U5770 (N_5770,N_2265,N_3043);
and U5771 (N_5771,N_3324,N_2196);
and U5772 (N_5772,N_2225,N_2738);
or U5773 (N_5773,N_3895,N_3559);
or U5774 (N_5774,N_2436,N_2284);
nand U5775 (N_5775,N_3595,N_2146);
or U5776 (N_5776,N_2709,N_3726);
xnor U5777 (N_5777,N_3911,N_2633);
xnor U5778 (N_5778,N_3564,N_2351);
xor U5779 (N_5779,N_2402,N_3054);
nand U5780 (N_5780,N_3219,N_3273);
and U5781 (N_5781,N_2758,N_3387);
xnor U5782 (N_5782,N_2068,N_3425);
and U5783 (N_5783,N_3652,N_3568);
or U5784 (N_5784,N_2673,N_3530);
xor U5785 (N_5785,N_3445,N_3901);
nand U5786 (N_5786,N_2673,N_2102);
xnor U5787 (N_5787,N_3830,N_3253);
xor U5788 (N_5788,N_3422,N_3343);
nor U5789 (N_5789,N_2872,N_3486);
xor U5790 (N_5790,N_3836,N_2958);
xor U5791 (N_5791,N_2329,N_2521);
nand U5792 (N_5792,N_2402,N_3276);
nand U5793 (N_5793,N_3179,N_2565);
and U5794 (N_5794,N_3627,N_3134);
xor U5795 (N_5795,N_3641,N_3313);
or U5796 (N_5796,N_2617,N_2457);
and U5797 (N_5797,N_3335,N_3081);
and U5798 (N_5798,N_2437,N_3887);
nor U5799 (N_5799,N_3160,N_3941);
xnor U5800 (N_5800,N_2961,N_2416);
or U5801 (N_5801,N_3985,N_3747);
xor U5802 (N_5802,N_2110,N_3297);
xor U5803 (N_5803,N_2920,N_3829);
nand U5804 (N_5804,N_2368,N_2215);
or U5805 (N_5805,N_2643,N_2633);
nand U5806 (N_5806,N_2911,N_2944);
xor U5807 (N_5807,N_2679,N_2726);
or U5808 (N_5808,N_2457,N_3234);
nor U5809 (N_5809,N_3547,N_2344);
xor U5810 (N_5810,N_2185,N_3095);
nand U5811 (N_5811,N_2830,N_3775);
and U5812 (N_5812,N_2917,N_3971);
nor U5813 (N_5813,N_2691,N_3886);
xor U5814 (N_5814,N_3228,N_2213);
nand U5815 (N_5815,N_2097,N_2926);
nand U5816 (N_5816,N_3641,N_3814);
or U5817 (N_5817,N_3161,N_2484);
nor U5818 (N_5818,N_3823,N_2292);
and U5819 (N_5819,N_2097,N_2095);
and U5820 (N_5820,N_2868,N_2497);
or U5821 (N_5821,N_2410,N_2829);
nand U5822 (N_5822,N_2488,N_3414);
or U5823 (N_5823,N_2246,N_2705);
or U5824 (N_5824,N_2034,N_2828);
nor U5825 (N_5825,N_3661,N_3999);
and U5826 (N_5826,N_3515,N_3769);
and U5827 (N_5827,N_2199,N_2458);
nand U5828 (N_5828,N_2884,N_3200);
and U5829 (N_5829,N_2014,N_3696);
nand U5830 (N_5830,N_3645,N_2369);
and U5831 (N_5831,N_2705,N_2649);
or U5832 (N_5832,N_2080,N_3007);
xor U5833 (N_5833,N_2605,N_3256);
nand U5834 (N_5834,N_3677,N_2148);
and U5835 (N_5835,N_2823,N_3464);
and U5836 (N_5836,N_3906,N_2811);
or U5837 (N_5837,N_3123,N_2675);
xor U5838 (N_5838,N_2083,N_2532);
nor U5839 (N_5839,N_2296,N_2135);
and U5840 (N_5840,N_3352,N_2337);
xnor U5841 (N_5841,N_3573,N_2203);
or U5842 (N_5842,N_3420,N_3059);
xnor U5843 (N_5843,N_2673,N_2122);
xor U5844 (N_5844,N_3853,N_3467);
nand U5845 (N_5845,N_3634,N_2392);
and U5846 (N_5846,N_3424,N_3669);
xnor U5847 (N_5847,N_2022,N_3025);
xnor U5848 (N_5848,N_3315,N_2060);
or U5849 (N_5849,N_3038,N_2235);
xor U5850 (N_5850,N_2715,N_3324);
nor U5851 (N_5851,N_3553,N_2797);
nand U5852 (N_5852,N_2071,N_2001);
and U5853 (N_5853,N_3454,N_2499);
nor U5854 (N_5854,N_2113,N_3304);
and U5855 (N_5855,N_3017,N_2501);
or U5856 (N_5856,N_2103,N_2819);
nand U5857 (N_5857,N_3870,N_2534);
nand U5858 (N_5858,N_3762,N_2476);
nor U5859 (N_5859,N_2171,N_3564);
and U5860 (N_5860,N_3041,N_2311);
or U5861 (N_5861,N_3593,N_3336);
xnor U5862 (N_5862,N_3424,N_2267);
and U5863 (N_5863,N_2195,N_2075);
nand U5864 (N_5864,N_3350,N_3530);
and U5865 (N_5865,N_3361,N_3974);
or U5866 (N_5866,N_2439,N_3999);
and U5867 (N_5867,N_2925,N_2087);
and U5868 (N_5868,N_3954,N_3121);
nand U5869 (N_5869,N_2794,N_3732);
xnor U5870 (N_5870,N_2475,N_2329);
nand U5871 (N_5871,N_2428,N_2917);
nor U5872 (N_5872,N_2311,N_3721);
xnor U5873 (N_5873,N_2051,N_2116);
nand U5874 (N_5874,N_3652,N_3424);
xnor U5875 (N_5875,N_2596,N_3807);
nor U5876 (N_5876,N_3467,N_3087);
xor U5877 (N_5877,N_2668,N_2640);
or U5878 (N_5878,N_2964,N_3112);
nand U5879 (N_5879,N_3488,N_2430);
nand U5880 (N_5880,N_2232,N_3010);
nor U5881 (N_5881,N_2672,N_2164);
or U5882 (N_5882,N_2360,N_2696);
xnor U5883 (N_5883,N_2349,N_3338);
xnor U5884 (N_5884,N_3838,N_2635);
or U5885 (N_5885,N_2851,N_2353);
or U5886 (N_5886,N_2857,N_3033);
and U5887 (N_5887,N_2479,N_3251);
nor U5888 (N_5888,N_3096,N_2844);
or U5889 (N_5889,N_2314,N_3938);
nor U5890 (N_5890,N_2631,N_3320);
or U5891 (N_5891,N_2762,N_3115);
nor U5892 (N_5892,N_2797,N_2433);
and U5893 (N_5893,N_2735,N_3154);
nor U5894 (N_5894,N_2462,N_2629);
nand U5895 (N_5895,N_2218,N_3739);
or U5896 (N_5896,N_2801,N_3565);
and U5897 (N_5897,N_3350,N_3492);
or U5898 (N_5898,N_2561,N_3244);
or U5899 (N_5899,N_2183,N_2661);
nand U5900 (N_5900,N_3797,N_3698);
xor U5901 (N_5901,N_2695,N_2040);
nand U5902 (N_5902,N_2516,N_2686);
or U5903 (N_5903,N_3529,N_2387);
xnor U5904 (N_5904,N_3420,N_3839);
nand U5905 (N_5905,N_2694,N_3203);
xnor U5906 (N_5906,N_3042,N_2694);
xor U5907 (N_5907,N_2254,N_3592);
xnor U5908 (N_5908,N_2982,N_3891);
or U5909 (N_5909,N_2919,N_3210);
and U5910 (N_5910,N_2362,N_3836);
nor U5911 (N_5911,N_2196,N_3234);
nor U5912 (N_5912,N_2654,N_2739);
nand U5913 (N_5913,N_3621,N_2988);
or U5914 (N_5914,N_2859,N_2052);
nand U5915 (N_5915,N_3221,N_2283);
nor U5916 (N_5916,N_2417,N_2097);
nand U5917 (N_5917,N_3378,N_2625);
nor U5918 (N_5918,N_3240,N_3456);
and U5919 (N_5919,N_2927,N_2419);
nor U5920 (N_5920,N_3743,N_2398);
nor U5921 (N_5921,N_2153,N_2894);
nand U5922 (N_5922,N_3306,N_2914);
or U5923 (N_5923,N_3527,N_2887);
xnor U5924 (N_5924,N_2950,N_2516);
nor U5925 (N_5925,N_3984,N_3847);
nor U5926 (N_5926,N_3423,N_3169);
nand U5927 (N_5927,N_2288,N_3099);
nand U5928 (N_5928,N_3618,N_2089);
xnor U5929 (N_5929,N_3955,N_2616);
nand U5930 (N_5930,N_2177,N_3536);
or U5931 (N_5931,N_3500,N_2465);
nand U5932 (N_5932,N_2738,N_2309);
nand U5933 (N_5933,N_2895,N_2472);
nor U5934 (N_5934,N_3119,N_3080);
nand U5935 (N_5935,N_3155,N_2892);
and U5936 (N_5936,N_3912,N_2057);
nor U5937 (N_5937,N_2443,N_2216);
or U5938 (N_5938,N_2859,N_2468);
nor U5939 (N_5939,N_3251,N_2653);
and U5940 (N_5940,N_3892,N_3583);
nor U5941 (N_5941,N_3985,N_2920);
nor U5942 (N_5942,N_3600,N_2805);
and U5943 (N_5943,N_2804,N_2776);
and U5944 (N_5944,N_2424,N_2088);
nor U5945 (N_5945,N_3289,N_2448);
xor U5946 (N_5946,N_3788,N_3977);
or U5947 (N_5947,N_2878,N_3470);
or U5948 (N_5948,N_2683,N_3979);
xor U5949 (N_5949,N_3437,N_3332);
nand U5950 (N_5950,N_3963,N_3547);
or U5951 (N_5951,N_2041,N_3109);
nand U5952 (N_5952,N_2146,N_3084);
xnor U5953 (N_5953,N_3336,N_3842);
xor U5954 (N_5954,N_2905,N_2741);
nor U5955 (N_5955,N_2841,N_3616);
xor U5956 (N_5956,N_2642,N_3341);
or U5957 (N_5957,N_2630,N_2256);
and U5958 (N_5958,N_3007,N_3855);
and U5959 (N_5959,N_2853,N_2847);
nand U5960 (N_5960,N_2146,N_2050);
nand U5961 (N_5961,N_3029,N_3040);
or U5962 (N_5962,N_2541,N_3031);
xor U5963 (N_5963,N_2354,N_2914);
or U5964 (N_5964,N_2960,N_2402);
or U5965 (N_5965,N_2777,N_2486);
nor U5966 (N_5966,N_3048,N_3761);
or U5967 (N_5967,N_2356,N_3765);
xor U5968 (N_5968,N_2762,N_2054);
nor U5969 (N_5969,N_3042,N_3537);
xnor U5970 (N_5970,N_3289,N_2770);
and U5971 (N_5971,N_2428,N_2517);
nand U5972 (N_5972,N_2577,N_2648);
nor U5973 (N_5973,N_3828,N_2907);
nor U5974 (N_5974,N_2883,N_2088);
nand U5975 (N_5975,N_2360,N_3903);
or U5976 (N_5976,N_2578,N_3483);
and U5977 (N_5977,N_3899,N_2343);
nand U5978 (N_5978,N_3062,N_2001);
nor U5979 (N_5979,N_2356,N_3835);
or U5980 (N_5980,N_2711,N_2658);
nor U5981 (N_5981,N_3898,N_2242);
nand U5982 (N_5982,N_2193,N_2892);
and U5983 (N_5983,N_3143,N_3218);
nand U5984 (N_5984,N_3742,N_2063);
nand U5985 (N_5985,N_2019,N_3682);
xor U5986 (N_5986,N_2029,N_3777);
nor U5987 (N_5987,N_2279,N_3204);
or U5988 (N_5988,N_3678,N_3601);
xnor U5989 (N_5989,N_3245,N_2603);
or U5990 (N_5990,N_2413,N_2484);
and U5991 (N_5991,N_3981,N_3390);
nor U5992 (N_5992,N_3403,N_3140);
xor U5993 (N_5993,N_2911,N_3862);
or U5994 (N_5994,N_3804,N_2118);
xor U5995 (N_5995,N_3601,N_3972);
nor U5996 (N_5996,N_3140,N_3087);
and U5997 (N_5997,N_2955,N_2489);
or U5998 (N_5998,N_3720,N_2726);
or U5999 (N_5999,N_2191,N_3733);
xor U6000 (N_6000,N_4635,N_5603);
nor U6001 (N_6001,N_4016,N_5760);
nor U6002 (N_6002,N_5389,N_4186);
nor U6003 (N_6003,N_5573,N_4642);
nor U6004 (N_6004,N_4444,N_5981);
or U6005 (N_6005,N_5771,N_4643);
nor U6006 (N_6006,N_5480,N_4871);
xnor U6007 (N_6007,N_4725,N_4651);
nor U6008 (N_6008,N_5535,N_4422);
and U6009 (N_6009,N_4092,N_5166);
xor U6010 (N_6010,N_5158,N_4692);
or U6011 (N_6011,N_5410,N_4714);
nand U6012 (N_6012,N_4116,N_5505);
nor U6013 (N_6013,N_5422,N_5338);
nor U6014 (N_6014,N_5330,N_5185);
and U6015 (N_6015,N_4438,N_5590);
or U6016 (N_6016,N_5634,N_5472);
or U6017 (N_6017,N_4595,N_4830);
nand U6018 (N_6018,N_4787,N_4345);
xor U6019 (N_6019,N_4475,N_4081);
and U6020 (N_6020,N_4377,N_4279);
nand U6021 (N_6021,N_5041,N_4814);
nor U6022 (N_6022,N_4559,N_4056);
and U6023 (N_6023,N_4812,N_4716);
nor U6024 (N_6024,N_5841,N_4650);
nor U6025 (N_6025,N_5206,N_5163);
nand U6026 (N_6026,N_5600,N_5794);
nor U6027 (N_6027,N_5486,N_5701);
and U6028 (N_6028,N_4862,N_4959);
nor U6029 (N_6029,N_4682,N_5539);
and U6030 (N_6030,N_5609,N_5605);
or U6031 (N_6031,N_4143,N_5591);
nor U6032 (N_6032,N_5332,N_5902);
or U6033 (N_6033,N_5075,N_5008);
nand U6034 (N_6034,N_4407,N_4515);
nor U6035 (N_6035,N_5866,N_5584);
xor U6036 (N_6036,N_5226,N_5451);
xnor U6037 (N_6037,N_4263,N_4035);
nor U6038 (N_6038,N_4903,N_4027);
nor U6039 (N_6039,N_4057,N_5615);
nor U6040 (N_6040,N_5563,N_4397);
nand U6041 (N_6041,N_4896,N_4046);
nand U6042 (N_6042,N_4901,N_4111);
or U6043 (N_6043,N_5840,N_5756);
or U6044 (N_6044,N_5720,N_4165);
nor U6045 (N_6045,N_4512,N_5191);
or U6046 (N_6046,N_5703,N_5299);
nor U6047 (N_6047,N_5298,N_5820);
and U6048 (N_6048,N_5278,N_5414);
xor U6049 (N_6049,N_5254,N_4014);
nand U6050 (N_6050,N_4877,N_4630);
nand U6051 (N_6051,N_4693,N_5672);
xnor U6052 (N_6052,N_5138,N_4724);
nor U6053 (N_6053,N_5575,N_5196);
nor U6054 (N_6054,N_4169,N_4596);
or U6055 (N_6055,N_5343,N_5025);
nand U6056 (N_6056,N_5581,N_4529);
and U6057 (N_6057,N_4209,N_4711);
nor U6058 (N_6058,N_5007,N_5117);
and U6059 (N_6059,N_5790,N_4536);
or U6060 (N_6060,N_5893,N_4460);
and U6061 (N_6061,N_5839,N_4742);
xnor U6062 (N_6062,N_4308,N_4599);
nor U6063 (N_6063,N_5776,N_4341);
nor U6064 (N_6064,N_5415,N_5355);
nand U6065 (N_6065,N_5905,N_4328);
xor U6066 (N_6066,N_5228,N_4404);
and U6067 (N_6067,N_4082,N_4819);
xnor U6068 (N_6068,N_4031,N_5870);
or U6069 (N_6069,N_5656,N_4605);
nand U6070 (N_6070,N_4508,N_4996);
and U6071 (N_6071,N_5678,N_4876);
xor U6072 (N_6072,N_4421,N_5888);
nand U6073 (N_6073,N_5459,N_5210);
xnor U6074 (N_6074,N_4948,N_5111);
nor U6075 (N_6075,N_5379,N_5684);
and U6076 (N_6076,N_4006,N_5346);
xor U6077 (N_6077,N_4244,N_5294);
and U6078 (N_6078,N_4592,N_4990);
xnor U6079 (N_6079,N_5808,N_5824);
xnor U6080 (N_6080,N_5154,N_4322);
nand U6081 (N_6081,N_5412,N_5621);
and U6082 (N_6082,N_5903,N_5778);
or U6083 (N_6083,N_5217,N_4267);
nand U6084 (N_6084,N_4201,N_5243);
nor U6085 (N_6085,N_5620,N_4933);
xnor U6086 (N_6086,N_5939,N_5324);
and U6087 (N_6087,N_5682,N_5960);
or U6088 (N_6088,N_5876,N_5917);
and U6089 (N_6089,N_4668,N_5209);
nor U6090 (N_6090,N_4618,N_4989);
nor U6091 (N_6091,N_5491,N_4585);
xor U6092 (N_6092,N_5132,N_5918);
or U6093 (N_6093,N_5317,N_4502);
xor U6094 (N_6094,N_5947,N_5441);
xor U6095 (N_6095,N_4604,N_4778);
or U6096 (N_6096,N_5393,N_5815);
xor U6097 (N_6097,N_4089,N_5050);
nand U6098 (N_6098,N_4146,N_4252);
or U6099 (N_6099,N_4417,N_4325);
nor U6100 (N_6100,N_5433,N_5851);
nand U6101 (N_6101,N_4196,N_5817);
or U6102 (N_6102,N_4575,N_5349);
and U6103 (N_6103,N_4550,N_4398);
or U6104 (N_6104,N_4256,N_4374);
xor U6105 (N_6105,N_5353,N_5589);
nand U6106 (N_6106,N_5855,N_4227);
and U6107 (N_6107,N_5366,N_5085);
xor U6108 (N_6108,N_5836,N_5262);
and U6109 (N_6109,N_4570,N_5896);
xor U6110 (N_6110,N_4102,N_5694);
or U6111 (N_6111,N_4270,N_5199);
xor U6112 (N_6112,N_5499,N_4940);
and U6113 (N_6113,N_5181,N_4734);
and U6114 (N_6114,N_4891,N_4327);
and U6115 (N_6115,N_5922,N_4358);
or U6116 (N_6116,N_4426,N_4739);
nand U6117 (N_6117,N_4334,N_5301);
and U6118 (N_6118,N_4266,N_5979);
nand U6119 (N_6119,N_4413,N_5235);
nand U6120 (N_6120,N_5675,N_4880);
xnor U6121 (N_6121,N_4750,N_4507);
nand U6122 (N_6122,N_5380,N_4354);
nor U6123 (N_6123,N_5160,N_5009);
or U6124 (N_6124,N_4674,N_5048);
nor U6125 (N_6125,N_4535,N_4801);
xor U6126 (N_6126,N_4130,N_4123);
xor U6127 (N_6127,N_4818,N_4956);
nand U6128 (N_6128,N_5592,N_4236);
or U6129 (N_6129,N_5359,N_4984);
and U6130 (N_6130,N_5222,N_4136);
or U6131 (N_6131,N_4820,N_4297);
xor U6132 (N_6132,N_4237,N_5173);
or U6133 (N_6133,N_5819,N_5131);
nand U6134 (N_6134,N_5976,N_5424);
nand U6135 (N_6135,N_4802,N_5237);
nor U6136 (N_6136,N_4840,N_4690);
nand U6137 (N_6137,N_5143,N_4086);
nand U6138 (N_6138,N_4681,N_5497);
or U6139 (N_6139,N_5426,N_5205);
nor U6140 (N_6140,N_5345,N_5973);
or U6141 (N_6141,N_5718,N_4122);
nand U6142 (N_6142,N_5921,N_5202);
nand U6143 (N_6143,N_4405,N_5333);
nand U6144 (N_6144,N_4489,N_4101);
xor U6145 (N_6145,N_4803,N_5289);
xor U6146 (N_6146,N_5425,N_5619);
nand U6147 (N_6147,N_4845,N_5101);
xnor U6148 (N_6148,N_5381,N_5329);
and U6149 (N_6149,N_4694,N_4753);
nand U6150 (N_6150,N_4850,N_4077);
nand U6151 (N_6151,N_4906,N_4902);
nand U6152 (N_6152,N_5115,N_5428);
xor U6153 (N_6153,N_4305,N_5314);
nor U6154 (N_6154,N_5987,N_5477);
and U6155 (N_6155,N_4021,N_4163);
nor U6156 (N_6156,N_5285,N_5977);
and U6157 (N_6157,N_5027,N_5204);
xnor U6158 (N_6158,N_4556,N_4010);
and U6159 (N_6159,N_4540,N_4718);
or U6160 (N_6160,N_5526,N_5315);
xnor U6161 (N_6161,N_5668,N_5496);
xor U6162 (N_6162,N_5372,N_5689);
or U6163 (N_6163,N_4825,N_4464);
nor U6164 (N_6164,N_5801,N_5698);
or U6165 (N_6165,N_5242,N_4406);
or U6166 (N_6166,N_4329,N_5128);
or U6167 (N_6167,N_5089,N_4827);
and U6168 (N_6168,N_5554,N_5997);
nor U6169 (N_6169,N_5475,N_5356);
xor U6170 (N_6170,N_4688,N_4770);
or U6171 (N_6171,N_5853,N_4409);
nand U6172 (N_6172,N_5508,N_5377);
nor U6173 (N_6173,N_5963,N_5564);
xnor U6174 (N_6174,N_5003,N_5560);
xor U6175 (N_6175,N_5558,N_5275);
and U6176 (N_6176,N_5923,N_4894);
nor U6177 (N_6177,N_5419,N_4865);
or U6178 (N_6178,N_4441,N_4211);
nor U6179 (N_6179,N_4918,N_5889);
nor U6180 (N_6180,N_4979,N_4844);
nor U6181 (N_6181,N_5019,N_5829);
or U6182 (N_6182,N_4808,N_5962);
nor U6183 (N_6183,N_5369,N_5982);
and U6184 (N_6184,N_4188,N_4577);
nor U6185 (N_6185,N_4713,N_5442);
xnor U6186 (N_6186,N_5537,N_4612);
or U6187 (N_6187,N_5017,N_5717);
nand U6188 (N_6188,N_5719,N_4966);
nand U6189 (N_6189,N_5928,N_4275);
nand U6190 (N_6190,N_5268,N_5129);
nand U6191 (N_6191,N_5586,N_4884);
nor U6192 (N_6192,N_5772,N_5791);
or U6193 (N_6193,N_5283,N_5704);
nor U6194 (N_6194,N_4623,N_4302);
and U6195 (N_6195,N_5710,N_5403);
xnor U6196 (N_6196,N_4205,N_4704);
nor U6197 (N_6197,N_4180,N_4134);
or U6198 (N_6198,N_5904,N_5837);
xnor U6199 (N_6199,N_4272,N_5318);
nand U6200 (N_6200,N_4166,N_5616);
nand U6201 (N_6201,N_5219,N_4469);
or U6202 (N_6202,N_4799,N_5953);
nand U6203 (N_6203,N_4942,N_4888);
nor U6204 (N_6204,N_5809,N_4910);
and U6205 (N_6205,N_4593,N_4574);
nor U6206 (N_6206,N_4034,N_4747);
nor U6207 (N_6207,N_4361,N_4572);
or U6208 (N_6208,N_4622,N_5002);
nand U6209 (N_6209,N_5144,N_5378);
xnor U6210 (N_6210,N_4359,N_5828);
nor U6211 (N_6211,N_5340,N_5806);
and U6212 (N_6212,N_5660,N_4615);
nand U6213 (N_6213,N_4456,N_4994);
and U6214 (N_6214,N_5421,N_4241);
nand U6215 (N_6215,N_4706,N_5465);
nand U6216 (N_6216,N_5911,N_5733);
and U6217 (N_6217,N_5773,N_4807);
and U6218 (N_6218,N_5201,N_4659);
and U6219 (N_6219,N_4107,N_4664);
nor U6220 (N_6220,N_5388,N_4881);
or U6221 (N_6221,N_5082,N_4197);
or U6222 (N_6222,N_4523,N_5524);
and U6223 (N_6223,N_4946,N_4821);
nand U6224 (N_6224,N_4366,N_5813);
xor U6225 (N_6225,N_5259,N_5325);
xor U6226 (N_6226,N_4393,N_5513);
or U6227 (N_6227,N_4069,N_5382);
xor U6228 (N_6228,N_4727,N_4192);
nor U6229 (N_6229,N_4983,N_4723);
and U6230 (N_6230,N_4033,N_4153);
nor U6231 (N_6231,N_4829,N_5220);
xor U6232 (N_6232,N_4219,N_5188);
nor U6233 (N_6233,N_4066,N_5140);
or U6234 (N_6234,N_4721,N_4480);
nor U6235 (N_6235,N_4178,N_4396);
and U6236 (N_6236,N_4986,N_4553);
nor U6237 (N_6237,N_5081,N_5725);
or U6238 (N_6238,N_5948,N_5737);
or U6239 (N_6239,N_5444,N_5625);
nand U6240 (N_6240,N_4949,N_5578);
and U6241 (N_6241,N_5941,N_4832);
xnor U6242 (N_6242,N_5547,N_5241);
or U6243 (N_6243,N_5331,N_5116);
and U6244 (N_6244,N_5282,N_4943);
xnor U6245 (N_6245,N_5845,N_4506);
or U6246 (N_6246,N_4890,N_4194);
and U6247 (N_6247,N_5297,N_4045);
or U6248 (N_6248,N_4947,N_4970);
nand U6249 (N_6249,N_4783,N_4478);
nor U6250 (N_6250,N_5098,N_4108);
xnor U6251 (N_6251,N_4125,N_5856);
or U6252 (N_6252,N_5023,N_5553);
or U6253 (N_6253,N_5295,N_5057);
xnor U6254 (N_6254,N_5792,N_4632);
nand U6255 (N_6255,N_5247,N_5397);
or U6256 (N_6256,N_4927,N_5469);
nor U6257 (N_6257,N_5804,N_4520);
nor U6258 (N_6258,N_5047,N_4126);
nor U6259 (N_6259,N_4453,N_5165);
nor U6260 (N_6260,N_5988,N_4371);
xnor U6261 (N_6261,N_4479,N_5755);
nand U6262 (N_6262,N_5125,N_5763);
or U6263 (N_6263,N_5336,N_5245);
or U6264 (N_6264,N_4145,N_5074);
nand U6265 (N_6265,N_4864,N_5476);
and U6266 (N_6266,N_4709,N_4598);
or U6267 (N_6267,N_4156,N_4543);
nor U6268 (N_6268,N_5443,N_4376);
xnor U6269 (N_6269,N_5745,N_4809);
nand U6270 (N_6270,N_5086,N_4299);
or U6271 (N_6271,N_4050,N_4395);
nand U6272 (N_6272,N_4260,N_4815);
xnor U6273 (N_6273,N_4149,N_5139);
nand U6274 (N_6274,N_5944,N_4055);
xor U6275 (N_6275,N_4430,N_4262);
nor U6276 (N_6276,N_4836,N_4869);
xor U6277 (N_6277,N_4761,N_4843);
and U6278 (N_6278,N_4254,N_4895);
nand U6279 (N_6279,N_4442,N_5203);
xor U6280 (N_6280,N_4174,N_4995);
nand U6281 (N_6281,N_5651,N_5416);
xor U6282 (N_6282,N_5900,N_5863);
and U6283 (N_6283,N_5118,N_5797);
or U6284 (N_6284,N_5954,N_5385);
or U6285 (N_6285,N_5934,N_5438);
nand U6286 (N_6286,N_4513,N_5598);
or U6287 (N_6287,N_4641,N_4958);
xor U6288 (N_6288,N_4760,N_4032);
nand U6289 (N_6289,N_5396,N_4477);
xor U6290 (N_6290,N_4017,N_4660);
nor U6291 (N_6291,N_5536,N_4658);
xnor U6292 (N_6292,N_5847,N_4849);
and U6293 (N_6293,N_5290,N_5775);
or U6294 (N_6294,N_4204,N_5207);
xnor U6295 (N_6295,N_4128,N_4976);
nor U6296 (N_6296,N_4346,N_4719);
or U6297 (N_6297,N_4104,N_4624);
and U6298 (N_6298,N_5213,N_5585);
or U6299 (N_6299,N_4235,N_5796);
or U6300 (N_6300,N_4217,N_5636);
xor U6301 (N_6301,N_5423,N_5088);
xor U6302 (N_6302,N_4924,N_4846);
nor U6303 (N_6303,N_5602,N_4603);
or U6304 (N_6304,N_5559,N_5826);
or U6305 (N_6305,N_5194,N_4562);
xor U6306 (N_6306,N_4425,N_5622);
and U6307 (N_6307,N_5402,N_5884);
xor U6308 (N_6308,N_4310,N_4011);
and U6309 (N_6309,N_4487,N_5112);
nor U6310 (N_6310,N_4208,N_4732);
xnor U6311 (N_6311,N_4062,N_5453);
xor U6312 (N_6312,N_5649,N_5195);
nor U6313 (N_6313,N_5153,N_5093);
and U6314 (N_6314,N_4786,N_5488);
and U6315 (N_6315,N_5696,N_5838);
nand U6316 (N_6316,N_5229,N_4158);
nor U6317 (N_6317,N_4151,N_4993);
xnor U6318 (N_6318,N_5662,N_5786);
nand U6319 (N_6319,N_4403,N_5507);
nand U6320 (N_6320,N_5061,N_5261);
or U6321 (N_6321,N_5528,N_5858);
and U6322 (N_6322,N_4661,N_5454);
and U6323 (N_6323,N_4448,N_4736);
xor U6324 (N_6324,N_5542,N_4457);
nand U6325 (N_6325,N_5990,N_4588);
xor U6326 (N_6326,N_4646,N_5707);
xor U6327 (N_6327,N_5814,N_4283);
nor U6328 (N_6328,N_5551,N_4019);
or U6329 (N_6329,N_5159,N_4352);
nor U6330 (N_6330,N_5624,N_5799);
nor U6331 (N_6331,N_5640,N_4521);
xor U6332 (N_6332,N_4909,N_4029);
and U6333 (N_6333,N_4255,N_5652);
xor U6334 (N_6334,N_5168,N_4955);
or U6335 (N_6335,N_5852,N_5705);
nand U6336 (N_6336,N_5404,N_5642);
or U6337 (N_6337,N_4051,N_4185);
nand U6338 (N_6338,N_4571,N_4701);
or U6339 (N_6339,N_5092,N_4351);
xnor U6340 (N_6340,N_4720,N_4773);
nor U6341 (N_6341,N_5506,N_5321);
nor U6342 (N_6342,N_4386,N_5945);
and U6343 (N_6343,N_5328,N_4885);
xnor U6344 (N_6344,N_5780,N_4078);
or U6345 (N_6345,N_5060,N_5341);
xnor U6346 (N_6346,N_4852,N_4538);
nand U6347 (N_6347,N_5835,N_4580);
or U6348 (N_6348,N_4446,N_5255);
xor U6349 (N_6349,N_4755,N_5972);
nor U6350 (N_6350,N_5272,N_5909);
and U6351 (N_6351,N_5253,N_4440);
xor U6352 (N_6352,N_5955,N_4497);
nand U6353 (N_6353,N_5610,N_4917);
xor U6354 (N_6354,N_5680,N_5842);
and U6355 (N_6355,N_4929,N_5064);
and U6356 (N_6356,N_5104,N_4915);
nor U6357 (N_6357,N_4613,N_4080);
nor U6358 (N_6358,N_5788,N_4199);
nor U6359 (N_6359,N_4537,N_4301);
xnor U6360 (N_6360,N_4870,N_5930);
or U6361 (N_6361,N_4647,N_5239);
and U6362 (N_6362,N_4952,N_4191);
xor U6363 (N_6363,N_5054,N_5394);
or U6364 (N_6364,N_4127,N_4516);
xor U6365 (N_6365,N_5293,N_5561);
nor U6366 (N_6366,N_4431,N_4911);
nand U6367 (N_6367,N_4700,N_5761);
and U6368 (N_6368,N_5467,N_4542);
and U6369 (N_6369,N_4337,N_4519);
nand U6370 (N_6370,N_4118,N_4726);
and U6371 (N_6371,N_4054,N_4938);
and U6372 (N_6372,N_4638,N_5846);
and U6373 (N_6373,N_4968,N_5546);
nand U6374 (N_6374,N_4002,N_4967);
nor U6375 (N_6375,N_5574,N_4218);
or U6376 (N_6376,N_5249,N_5510);
nand U6377 (N_6377,N_5647,N_4388);
nand U6378 (N_6378,N_5304,N_5460);
nand U6379 (N_6379,N_4466,N_4913);
xor U6380 (N_6380,N_5823,N_5471);
xor U6381 (N_6381,N_4435,N_4212);
nand U6382 (N_6382,N_5549,N_5933);
and U6383 (N_6383,N_4291,N_4290);
nand U6384 (N_6384,N_4347,N_5937);
nand U6385 (N_6385,N_4539,N_4161);
or U6386 (N_6386,N_5100,N_4552);
nand U6387 (N_6387,N_4565,N_4988);
nand U6388 (N_6388,N_5248,N_4072);
nand U6389 (N_6389,N_5746,N_5929);
nor U6390 (N_6390,N_5627,N_5368);
and U6391 (N_6391,N_4309,N_4120);
nor U6392 (N_6392,N_4370,N_5663);
nand U6393 (N_6393,N_4600,N_4495);
and U6394 (N_6394,N_5674,N_4349);
nand U6395 (N_6395,N_4148,N_4978);
and U6396 (N_6396,N_4733,N_4528);
xnor U6397 (N_6397,N_5515,N_5391);
nor U6398 (N_6398,N_4883,N_5335);
xnor U6399 (N_6399,N_4231,N_4318);
and U6400 (N_6400,N_5572,N_4561);
nor U6401 (N_6401,N_4173,N_4831);
or U6402 (N_6402,N_4800,N_5969);
and U6403 (N_6403,N_5910,N_5735);
or U6404 (N_6404,N_4298,N_5031);
nand U6405 (N_6405,N_4926,N_4498);
or U6406 (N_6406,N_4566,N_5039);
xnor U6407 (N_6407,N_4243,N_4418);
nand U6408 (N_6408,N_5940,N_5730);
and U6409 (N_6409,N_4616,N_4476);
and U6410 (N_6410,N_5212,N_5258);
or U6411 (N_6411,N_5044,N_5223);
nand U6412 (N_6412,N_4645,N_5468);
xor U6413 (N_6413,N_5466,N_4568);
nor U6414 (N_6414,N_5700,N_5095);
xor U6415 (N_6415,N_4306,N_5626);
or U6416 (N_6416,N_4419,N_5908);
xor U6417 (N_6417,N_5018,N_5162);
xor U6418 (N_6418,N_5174,N_4109);
nor U6419 (N_6419,N_5952,N_4115);
nor U6420 (N_6420,N_5011,N_4810);
xor U6421 (N_6421,N_5270,N_5042);
and U6422 (N_6422,N_4432,N_4222);
xnor U6423 (N_6423,N_4505,N_4655);
nand U6424 (N_6424,N_5190,N_5458);
and U6425 (N_6425,N_5606,N_5915);
nor U6426 (N_6426,N_5277,N_5765);
and U6427 (N_6427,N_5512,N_5897);
xnor U6428 (N_6428,N_5296,N_5291);
and U6429 (N_6429,N_4246,N_4532);
or U6430 (N_6430,N_4841,N_5284);
nand U6431 (N_6431,N_5037,N_4024);
nor U6432 (N_6432,N_5807,N_5474);
nor U6433 (N_6433,N_5552,N_4065);
or U6434 (N_6434,N_4698,N_4551);
or U6435 (N_6435,N_4554,N_5545);
and U6436 (N_6436,N_5313,N_4385);
nand U6437 (N_6437,N_5722,N_4920);
xor U6438 (N_6438,N_4482,N_4640);
and U6439 (N_6439,N_4847,N_5518);
or U6440 (N_6440,N_5287,N_4304);
and U6441 (N_6441,N_4751,N_4467);
nor U6442 (N_6442,N_5795,N_4048);
or U6443 (N_6443,N_4030,N_5036);
xor U6444 (N_6444,N_4788,N_4708);
or U6445 (N_6445,N_5156,N_5005);
nor U6446 (N_6446,N_4908,N_5176);
nand U6447 (N_6447,N_4767,N_5126);
nand U6448 (N_6448,N_4590,N_5151);
or U6449 (N_6449,N_4360,N_5169);
nor U6450 (N_6450,N_4637,N_5757);
nor U6451 (N_6451,N_4144,N_5580);
nor U6452 (N_6452,N_5601,N_5992);
nand U6453 (N_6453,N_4930,N_5072);
xnor U6454 (N_6454,N_4768,N_5577);
nor U6455 (N_6455,N_4336,N_5736);
xor U6456 (N_6456,N_4277,N_4867);
nor U6457 (N_6457,N_4179,N_5094);
nor U6458 (N_6458,N_5727,N_4982);
nor U6459 (N_6459,N_4473,N_4129);
xnor U6460 (N_6460,N_4558,N_5632);
and U6461 (N_6461,N_5067,N_4228);
nor U6462 (N_6462,N_4198,N_5251);
nand U6463 (N_6463,N_4685,N_5032);
nand U6464 (N_6464,N_4587,N_4905);
xor U6465 (N_6465,N_5456,N_4594);
nand U6466 (N_6466,N_5702,N_5854);
and U6467 (N_6467,N_5492,N_4375);
and U6468 (N_6468,N_5256,N_5489);
nand U6469 (N_6469,N_4206,N_4147);
xor U6470 (N_6470,N_4712,N_4447);
and U6471 (N_6471,N_5175,N_5996);
or U6472 (N_6472,N_4973,N_4702);
xor U6473 (N_6473,N_5076,N_5646);
and U6474 (N_6474,N_5091,N_4644);
nor U6475 (N_6475,N_5161,N_5655);
nand U6476 (N_6476,N_4601,N_4541);
nor U6477 (N_6477,N_4063,N_5568);
and U6478 (N_6478,N_4088,N_4213);
and U6479 (N_6479,N_4221,N_5527);
xor U6480 (N_6480,N_5302,N_5058);
xor U6481 (N_6481,N_5635,N_4951);
or U6482 (N_6482,N_5015,N_5102);
xor U6483 (N_6483,N_4344,N_5699);
or U6484 (N_6484,N_4463,N_5420);
nand U6485 (N_6485,N_5119,N_4268);
nand U6486 (N_6486,N_5617,N_5726);
xor U6487 (N_6487,N_5978,N_5522);
xor U6488 (N_6488,N_4229,N_4522);
nand U6489 (N_6489,N_5122,N_5351);
nand U6490 (N_6490,N_5312,N_4546);
xor U6491 (N_6491,N_5950,N_4854);
and U6492 (N_6492,N_4292,N_4707);
nor U6493 (N_6493,N_5110,N_4452);
and U6494 (N_6494,N_4686,N_5305);
xor U6495 (N_6495,N_5965,N_4474);
and U6496 (N_6496,N_5501,N_5999);
nand U6497 (N_6497,N_5395,N_4459);
nor U6498 (N_6498,N_5686,N_4744);
or U6499 (N_6499,N_4012,N_5271);
or U6500 (N_6500,N_5715,N_4210);
and U6501 (N_6501,N_4060,N_5099);
nand U6502 (N_6502,N_5413,N_5511);
nor U6503 (N_6503,N_4090,N_4526);
nor U6504 (N_6504,N_4677,N_5754);
nand U6505 (N_6505,N_4294,N_5500);
nand U6506 (N_6506,N_5350,N_4455);
or U6507 (N_6507,N_4313,N_5376);
nor U6508 (N_6508,N_4443,N_4004);
xnor U6509 (N_6509,N_5728,N_4839);
nor U6510 (N_6510,N_5244,N_4873);
or U6511 (N_6511,N_4975,N_4138);
nor U6512 (N_6512,N_5430,N_5857);
nand U6513 (N_6513,N_4059,N_5665);
xnor U6514 (N_6514,N_4838,N_5805);
or U6515 (N_6515,N_4916,N_5850);
nor U6516 (N_6516,N_5648,N_4162);
and U6517 (N_6517,N_5587,N_4317);
and U6518 (N_6518,N_5743,N_5943);
or U6519 (N_6519,N_5409,N_5749);
and U6520 (N_6520,N_5777,N_5078);
or U6521 (N_6521,N_4289,N_5768);
nand U6522 (N_6522,N_5729,N_4240);
and U6523 (N_6523,N_5004,N_5803);
and U6524 (N_6524,N_5432,N_4022);
and U6525 (N_6525,N_5406,N_4094);
nor U6526 (N_6526,N_5583,N_4312);
and U6527 (N_6527,N_5874,N_4648);
and U6528 (N_6528,N_4972,N_4073);
nor U6529 (N_6529,N_5265,N_4544);
and U6530 (N_6530,N_4039,N_5567);
nor U6531 (N_6531,N_5225,N_5310);
or U6532 (N_6532,N_5907,N_5257);
or U6533 (N_6533,N_5431,N_4548);
nand U6534 (N_6534,N_4740,N_4020);
xnor U6535 (N_6535,N_4549,N_4139);
and U6536 (N_6536,N_5899,N_4414);
xor U6537 (N_6537,N_5849,N_4472);
nor U6538 (N_6538,N_5991,N_5557);
and U6539 (N_6539,N_4866,N_5967);
xnor U6540 (N_6540,N_5555,N_4484);
nand U6541 (N_6541,N_4944,N_4099);
and U6542 (N_6542,N_4335,N_4250);
and U6543 (N_6543,N_4665,N_4627);
xor U6544 (N_6544,N_5614,N_4857);
and U6545 (N_6545,N_5766,N_5523);
nor U6546 (N_6546,N_5582,N_4584);
or U6547 (N_6547,N_5800,N_4932);
xnor U6548 (N_6548,N_4569,N_5429);
and U6549 (N_6549,N_5079,N_4038);
nand U6550 (N_6550,N_4367,N_5071);
nor U6551 (N_6551,N_5604,N_4671);
nor U6552 (N_6552,N_5063,N_4183);
xnor U6553 (N_6553,N_4037,N_4348);
xnor U6554 (N_6554,N_4207,N_5473);
xnor U6555 (N_6555,N_5436,N_4889);
or U6556 (N_6556,N_4602,N_5623);
or U6557 (N_6557,N_5886,N_5654);
or U6558 (N_6558,N_4379,N_5938);
xor U6559 (N_6559,N_4981,N_4053);
nor U6560 (N_6560,N_5157,N_4415);
or U6561 (N_6561,N_4070,N_5731);
xor U6562 (N_6562,N_5949,N_5383);
or U6563 (N_6563,N_4084,N_4461);
and U6564 (N_6564,N_5155,N_5688);
nor U6565 (N_6565,N_5446,N_5274);
and U6566 (N_6566,N_5810,N_5762);
and U6567 (N_6567,N_4273,N_5146);
or U6568 (N_6568,N_5418,N_4257);
nand U6569 (N_6569,N_4606,N_4853);
nand U6570 (N_6570,N_4321,N_4992);
nand U6571 (N_6571,N_5266,N_4775);
and U6572 (N_6572,N_4485,N_5679);
xnor U6573 (N_6573,N_5924,N_4922);
nor U6574 (N_6574,N_5925,N_4675);
nand U6575 (N_6575,N_5040,N_4796);
xnor U6576 (N_6576,N_4776,N_4779);
xnor U6577 (N_6577,N_5137,N_5869);
or U6578 (N_6578,N_4074,N_4465);
nand U6579 (N_6579,N_4434,N_4381);
and U6580 (N_6580,N_4833,N_4611);
and U6581 (N_6581,N_5873,N_4728);
xor U6582 (N_6582,N_4261,N_4380);
or U6583 (N_6583,N_5448,N_5994);
and U6584 (N_6584,N_4657,N_5599);
nor U6585 (N_6585,N_5034,N_5142);
or U6586 (N_6586,N_4745,N_4445);
xor U6587 (N_6587,N_4481,N_4914);
and U6588 (N_6588,N_4639,N_4330);
nor U6589 (N_6589,N_5434,N_4295);
xnor U6590 (N_6590,N_5562,N_5883);
nor U6591 (N_6591,N_5734,N_4886);
nor U6592 (N_6592,N_4560,N_4965);
and U6593 (N_6593,N_4666,N_5200);
nor U6594 (N_6594,N_4503,N_4912);
and U6595 (N_6595,N_5407,N_5234);
nand U6596 (N_6596,N_4402,N_5957);
and U6597 (N_6597,N_4047,N_5352);
nand U6598 (N_6598,N_5216,N_5327);
nand U6599 (N_6599,N_5611,N_4389);
or U6600 (N_6600,N_4238,N_5891);
xor U6601 (N_6601,N_4654,N_5744);
and U6602 (N_6602,N_5830,N_5970);
nand U6603 (N_6603,N_4964,N_5090);
nand U6604 (N_6604,N_4769,N_4284);
or U6605 (N_6605,N_4937,N_5543);
xor U6606 (N_6606,N_4242,N_4851);
or U6607 (N_6607,N_4628,N_5759);
or U6608 (N_6608,N_5073,N_5676);
or U6609 (N_6609,N_4365,N_4510);
or U6610 (N_6610,N_5260,N_5875);
nand U6611 (N_6611,N_5692,N_5540);
xnor U6612 (N_6612,N_4372,N_4898);
nand U6613 (N_6613,N_5052,N_4509);
xnor U6614 (N_6614,N_5457,N_4200);
and U6615 (N_6615,N_5716,N_4251);
xor U6616 (N_6616,N_4499,N_4771);
nor U6617 (N_6617,N_4710,N_5816);
and U6618 (N_6618,N_5774,N_4245);
or U6619 (N_6619,N_4303,N_4676);
and U6620 (N_6620,N_4874,N_4044);
nor U6621 (N_6621,N_4177,N_4202);
or U6622 (N_6622,N_4095,N_5106);
nor U6623 (N_6623,N_5322,N_4400);
and U6624 (N_6624,N_5427,N_5781);
nor U6625 (N_6625,N_5693,N_4100);
xnor U6626 (N_6626,N_5831,N_4091);
and U6627 (N_6627,N_4555,N_4794);
nand U6628 (N_6628,N_4855,N_4806);
nand U6629 (N_6629,N_5645,N_5495);
and U6630 (N_6630,N_4680,N_4184);
and U6631 (N_6631,N_5303,N_4835);
and U6632 (N_6632,N_4015,N_5721);
nand U6633 (N_6633,N_5514,N_4316);
or U6634 (N_6634,N_5033,N_5931);
nand U6635 (N_6635,N_5877,N_4564);
nor U6636 (N_6636,N_4667,N_4311);
and U6637 (N_6637,N_4597,N_5152);
nand U6638 (N_6638,N_5758,N_4493);
or U6639 (N_6639,N_5215,N_5279);
nand U6640 (N_6640,N_4411,N_5739);
nand U6641 (N_6641,N_5983,N_5114);
nor U6642 (N_6642,N_5316,N_4176);
and U6643 (N_6643,N_5516,N_4936);
and U6644 (N_6644,N_5103,N_5898);
or U6645 (N_6645,N_4619,N_5386);
nor U6646 (N_6646,N_5461,N_5238);
or U6647 (N_6647,N_5502,N_5865);
xnor U6648 (N_6648,N_4097,N_5643);
or U6649 (N_6649,N_5861,N_5753);
xnor U6650 (N_6650,N_5764,N_5769);
nor U6651 (N_6651,N_5644,N_4882);
or U6652 (N_6652,N_5267,N_4036);
nand U6653 (N_6653,N_5405,N_5087);
nand U6654 (N_6654,N_4225,N_4717);
or U6655 (N_6655,N_4861,N_5821);
nor U6656 (N_6656,N_4678,N_4043);
or U6657 (N_6657,N_4563,N_5971);
nand U6658 (N_6658,N_5530,N_4813);
nand U6659 (N_6659,N_5198,N_5276);
nand U6660 (N_6660,N_5183,N_5319);
nand U6661 (N_6661,N_4899,N_4083);
or U6662 (N_6662,N_5641,N_4868);
nand U6663 (N_6663,N_4315,N_5784);
xor U6664 (N_6664,N_5056,N_4265);
nor U6665 (N_6665,N_5844,N_4963);
nor U6666 (N_6666,N_4061,N_4672);
or U6667 (N_6667,N_5484,N_4042);
or U6668 (N_6668,N_5463,N_5411);
nor U6669 (N_6669,N_5208,N_5452);
nand U6670 (N_6670,N_4649,N_5450);
nor U6671 (N_6671,N_5741,N_4534);
nor U6672 (N_6672,N_4817,N_4610);
or U6673 (N_6673,N_4919,N_4804);
nand U6674 (N_6674,N_5077,N_5280);
nand U6675 (N_6675,N_4621,N_4383);
xnor U6676 (N_6676,N_5892,N_5051);
nor U6677 (N_6677,N_4987,N_5782);
or U6678 (N_6678,N_4233,N_4106);
xor U6679 (N_6679,N_4772,N_4663);
nor U6680 (N_6680,N_4777,N_5334);
nor U6681 (N_6681,N_4282,N_4096);
and U6682 (N_6682,N_4164,N_5767);
nor U6683 (N_6683,N_5607,N_4793);
or U6684 (N_6684,N_4695,N_4009);
xor U6685 (N_6685,N_4697,N_4985);
nor U6686 (N_6686,N_4288,N_4028);
nor U6687 (N_6687,N_5447,N_5013);
xor U6688 (N_6688,N_4626,N_5485);
nor U6689 (N_6689,N_4382,N_5785);
xnor U6690 (N_6690,N_5479,N_4098);
and U6691 (N_6691,N_4064,N_4399);
nand U6692 (N_6692,N_4754,N_4150);
or U6693 (N_6693,N_5121,N_4759);
xnor U6694 (N_6694,N_4579,N_4140);
or U6695 (N_6695,N_5916,N_5001);
and U6696 (N_6696,N_5588,N_5390);
xnor U6697 (N_6697,N_5361,N_4068);
or U6698 (N_6698,N_4945,N_5868);
and U6699 (N_6699,N_4433,N_5521);
and U6700 (N_6700,N_5440,N_4629);
nor U6701 (N_6701,N_4897,N_4141);
nand U6702 (N_6702,N_5661,N_4175);
nand U6703 (N_6703,N_4974,N_4124);
and U6704 (N_6704,N_4232,N_5548);
or U6705 (N_6705,N_5935,N_4743);
nor U6706 (N_6706,N_4878,N_4041);
and U6707 (N_6707,N_5860,N_5659);
nand U6708 (N_6708,N_5273,N_5124);
and U6709 (N_6709,N_4320,N_5920);
nor U6710 (N_6710,N_4226,N_5113);
or U6711 (N_6711,N_4075,N_5365);
nand U6712 (N_6712,N_5020,N_5439);
xnor U6713 (N_6713,N_5141,N_4323);
nand U6714 (N_6714,N_5811,N_5747);
nor U6715 (N_6715,N_5519,N_4860);
or U6716 (N_6716,N_5148,N_4998);
or U6717 (N_6717,N_5083,N_5348);
nand U6718 (N_6718,N_5569,N_5362);
or U6719 (N_6719,N_4586,N_5197);
and U6720 (N_6720,N_5650,N_5887);
nor U6721 (N_6721,N_4748,N_4953);
nor U6722 (N_6722,N_4687,N_4731);
nand U6723 (N_6723,N_5264,N_4428);
and U6724 (N_6724,N_4935,N_4900);
and U6725 (N_6725,N_5049,N_5170);
or U6726 (N_6726,N_5862,N_4000);
nand U6727 (N_6727,N_5398,N_5914);
or U6728 (N_6728,N_4458,N_4187);
xor U6729 (N_6729,N_5483,N_5673);
nor U6730 (N_6730,N_4684,N_5751);
or U6731 (N_6731,N_5793,N_4362);
nand U6732 (N_6732,N_5010,N_5685);
nor U6733 (N_6733,N_4557,N_4790);
nor U6734 (N_6734,N_4110,N_4669);
xor U6735 (N_6735,N_4314,N_4858);
xnor U6736 (N_6736,N_4013,N_5022);
xnor U6737 (N_6737,N_5657,N_4780);
nor U6738 (N_6738,N_4633,N_4738);
nand U6739 (N_6739,N_4762,N_4269);
nor U6740 (N_6740,N_4872,N_4276);
xor U6741 (N_6741,N_4333,N_4494);
and U6742 (N_6742,N_4005,N_5164);
and U6743 (N_6743,N_4339,N_5375);
nand U6744 (N_6744,N_5566,N_4296);
or U6745 (N_6745,N_4950,N_4224);
and U6746 (N_6746,N_5520,N_4856);
nand U6747 (N_6747,N_5053,N_5724);
xor U6748 (N_6748,N_5783,N_5363);
nand U6749 (N_6749,N_5339,N_4368);
and U6750 (N_6750,N_4203,N_5133);
and U6751 (N_6751,N_4931,N_5400);
xor U6752 (N_6752,N_5630,N_4791);
nor U6753 (N_6753,N_5637,N_5787);
nand U6754 (N_6754,N_5211,N_5240);
nor U6755 (N_6755,N_5127,N_5681);
and U6756 (N_6756,N_4631,N_5822);
and U6757 (N_6757,N_4923,N_4159);
nand U6758 (N_6758,N_4999,N_5026);
nor U6759 (N_6759,N_4410,N_5344);
and U6760 (N_6760,N_5825,N_5509);
and U6761 (N_6761,N_4567,N_4749);
and U6762 (N_6762,N_5478,N_4249);
xor U6763 (N_6763,N_4271,N_5135);
or U6764 (N_6764,N_5014,N_4131);
xnor U6765 (N_6765,N_5712,N_4170);
nand U6766 (N_6766,N_4501,N_5354);
nand U6767 (N_6767,N_4798,N_5872);
and U6768 (N_6768,N_5045,N_5711);
nor U6769 (N_6769,N_5186,N_5926);
xor U6770 (N_6770,N_4067,N_5738);
xor U6771 (N_6771,N_4142,N_5859);
nand U6772 (N_6772,N_5108,N_4756);
nor U6773 (N_6773,N_4752,N_5084);
nor U6774 (N_6774,N_5848,N_4449);
and U6775 (N_6775,N_5030,N_4157);
xnor U6776 (N_6776,N_4531,N_5227);
and U6777 (N_6777,N_4525,N_4785);
or U6778 (N_6778,N_5269,N_4980);
xnor U6779 (N_6779,N_5946,N_4892);
nor U6780 (N_6780,N_5919,N_5812);
nand U6781 (N_6781,N_4451,N_5292);
nand U6782 (N_6782,N_4133,N_5843);
xnor U6783 (N_6783,N_4326,N_5667);
xnor U6784 (N_6784,N_5669,N_4488);
and U6785 (N_6785,N_4578,N_5529);
nor U6786 (N_6786,N_5105,N_4781);
xor U6787 (N_6787,N_4357,N_4114);
xnor U6788 (N_6788,N_5964,N_5232);
xor U6789 (N_6789,N_4617,N_4997);
nand U6790 (N_6790,N_4837,N_5628);
or U6791 (N_6791,N_5740,N_4008);
nand U6792 (N_6792,N_4450,N_5597);
nor U6793 (N_6793,N_4216,N_5579);
xnor U6794 (N_6794,N_5541,N_5570);
nand U6795 (N_6795,N_4258,N_5323);
nand U6796 (N_6796,N_4656,N_5288);
nand U6797 (N_6797,N_5593,N_5966);
and U6798 (N_6798,N_5069,N_4722);
nand U6799 (N_6799,N_4533,N_5912);
and U6800 (N_6800,N_5867,N_5462);
nor U6801 (N_6801,N_5281,N_5337);
or U6802 (N_6802,N_5770,N_5035);
and U6803 (N_6803,N_4904,N_4957);
and U6804 (N_6804,N_4928,N_5070);
or U6805 (N_6805,N_5818,N_5802);
xor U6806 (N_6806,N_4547,N_5311);
nor U6807 (N_6807,N_5986,N_4369);
and U6808 (N_6808,N_4182,N_5493);
nor U6809 (N_6809,N_4076,N_5732);
nand U6810 (N_6810,N_5913,N_4135);
and U6811 (N_6811,N_4653,N_4939);
or U6812 (N_6812,N_4782,N_5538);
nor U6813 (N_6813,N_4132,N_5576);
nor U6814 (N_6814,N_4757,N_4103);
xor U6815 (N_6815,N_4319,N_4679);
xnor U6816 (N_6816,N_4278,N_4789);
nor U6817 (N_6817,N_4573,N_5167);
and U6818 (N_6818,N_4391,N_4378);
or U6819 (N_6819,N_5445,N_4340);
nand U6820 (N_6820,N_5218,N_5374);
nand U6821 (N_6821,N_5998,N_5534);
and U6822 (N_6822,N_5000,N_4961);
nand U6823 (N_6823,N_5596,N_5307);
or U6824 (N_6824,N_5172,N_5029);
and U6825 (N_6825,N_4193,N_5308);
xnor U6826 (N_6826,N_5134,N_5482);
and U6827 (N_6827,N_4764,N_4941);
and U6828 (N_6828,N_5961,N_5878);
nor U6829 (N_6829,N_5958,N_5408);
and U6830 (N_6830,N_5360,N_5370);
or U6831 (N_6831,N_4471,N_4591);
and U6832 (N_6832,N_4816,N_5565);
and U6833 (N_6833,N_4427,N_5690);
and U6834 (N_6834,N_4576,N_5021);
nor U6835 (N_6835,N_5595,N_4287);
or U6836 (N_6836,N_4423,N_4589);
nand U6837 (N_6837,N_4625,N_5136);
nor U6838 (N_6838,N_5742,N_5687);
nor U6839 (N_6839,N_4355,N_5068);
nor U6840 (N_6840,N_4364,N_4137);
xnor U6841 (N_6841,N_4960,N_5714);
nor U6842 (N_6842,N_4514,N_4040);
and U6843 (N_6843,N_5189,N_4454);
nand U6844 (N_6844,N_5490,N_4470);
nand U6845 (N_6845,N_5371,N_4087);
or U6846 (N_6846,N_5193,N_5179);
nand U6847 (N_6847,N_5097,N_5401);
xnor U6848 (N_6848,N_4735,N_5932);
or U6849 (N_6849,N_5956,N_4343);
nor U6850 (N_6850,N_5286,N_4112);
or U6851 (N_6851,N_4079,N_4160);
nand U6852 (N_6852,N_4483,N_4052);
and U6853 (N_6853,N_4848,N_5177);
nand U6854 (N_6854,N_5658,N_4608);
nor U6855 (N_6855,N_5633,N_5171);
nand U6856 (N_6856,N_5880,N_5779);
nor U6857 (N_6857,N_5145,N_5709);
nand U6858 (N_6858,N_4392,N_5192);
nor U6859 (N_6859,N_4620,N_5503);
or U6860 (N_6860,N_4121,N_4307);
or U6861 (N_6861,N_4703,N_5594);
and U6862 (N_6862,N_4581,N_5481);
and U6863 (N_6863,N_4614,N_5901);
nor U6864 (N_6864,N_4977,N_4828);
and U6865 (N_6865,N_5464,N_5358);
nand U6866 (N_6866,N_4758,N_4007);
xor U6867 (N_6867,N_5985,N_4167);
nor U6868 (N_6868,N_4834,N_5455);
xor U6869 (N_6869,N_4673,N_4530);
and U6870 (N_6870,N_4018,N_5187);
or U6871 (N_6871,N_4492,N_5666);
nand U6872 (N_6872,N_4239,N_4954);
xor U6873 (N_6873,N_4893,N_5890);
nand U6874 (N_6874,N_5178,N_4293);
or U6875 (N_6875,N_5387,N_5180);
and U6876 (N_6876,N_4518,N_5533);
or U6877 (N_6877,N_4285,N_4181);
nor U6878 (N_6878,N_5989,N_4429);
and U6879 (N_6879,N_5392,N_4394);
nor U6880 (N_6880,N_4741,N_5833);
and U6881 (N_6881,N_4795,N_5437);
and U6882 (N_6882,N_4281,N_5384);
nor U6883 (N_6883,N_5066,N_4527);
nor U6884 (N_6884,N_5494,N_5012);
and U6885 (N_6885,N_4172,N_4921);
and U6886 (N_6886,N_4171,N_5043);
xor U6887 (N_6887,N_5252,N_5065);
nor U6888 (N_6888,N_4264,N_4154);
and U6889 (N_6889,N_4805,N_4253);
xnor U6890 (N_6890,N_5080,N_4350);
and U6891 (N_6891,N_5697,N_5695);
or U6892 (N_6892,N_5130,N_5364);
and U6893 (N_6893,N_4412,N_4907);
xor U6894 (N_6894,N_5671,N_5881);
xnor U6895 (N_6895,N_4496,N_4784);
xnor U6896 (N_6896,N_5357,N_4691);
and U6897 (N_6897,N_4859,N_4729);
and U6898 (N_6898,N_5230,N_5653);
nor U6899 (N_6899,N_5182,N_4113);
nor U6900 (N_6900,N_5214,N_4155);
and U6901 (N_6901,N_5885,N_5250);
xnor U6902 (N_6902,N_5750,N_4437);
xnor U6903 (N_6903,N_5417,N_5367);
or U6904 (N_6904,N_4408,N_5618);
xnor U6905 (N_6905,N_5062,N_5968);
or U6906 (N_6906,N_5571,N_5531);
nor U6907 (N_6907,N_5895,N_4730);
and U6908 (N_6908,N_5055,N_4105);
nand U6909 (N_6909,N_4274,N_5236);
nor U6910 (N_6910,N_5498,N_5347);
nor U6911 (N_6911,N_4468,N_5798);
nor U6912 (N_6912,N_4234,N_4765);
xnor U6913 (N_6913,N_5487,N_4524);
xor U6914 (N_6914,N_4436,N_5995);
or U6915 (N_6915,N_4195,N_4058);
nand U6916 (N_6916,N_5016,N_5677);
xnor U6917 (N_6917,N_4026,N_5879);
nor U6918 (N_6918,N_5894,N_4634);
or U6919 (N_6919,N_4420,N_5871);
or U6920 (N_6920,N_5613,N_4331);
nand U6921 (N_6921,N_4500,N_5399);
xor U6922 (N_6922,N_4763,N_4670);
xor U6923 (N_6923,N_5974,N_5748);
xor U6924 (N_6924,N_5300,N_5670);
nand U6925 (N_6925,N_4607,N_4025);
nand U6926 (N_6926,N_5942,N_4934);
and U6927 (N_6927,N_4925,N_5149);
and U6928 (N_6928,N_4168,N_4390);
or U6929 (N_6929,N_4300,N_5470);
and U6930 (N_6930,N_4824,N_4223);
or U6931 (N_6931,N_5984,N_5525);
and U6932 (N_6932,N_4545,N_5608);
nor U6933 (N_6933,N_4683,N_5306);
xor U6934 (N_6934,N_5975,N_5246);
nor U6935 (N_6935,N_5006,N_5096);
and U6936 (N_6936,N_5263,N_4511);
or U6937 (N_6937,N_5723,N_4491);
or U6938 (N_6938,N_4662,N_4792);
or U6939 (N_6939,N_5683,N_5951);
and U6940 (N_6940,N_5834,N_5713);
or U6941 (N_6941,N_4699,N_4774);
xor U6942 (N_6942,N_5224,N_4811);
xnor U6943 (N_6943,N_5936,N_4746);
and U6944 (N_6944,N_4490,N_4842);
nor U6945 (N_6945,N_4363,N_5664);
nand U6946 (N_6946,N_4356,N_5028);
xor U6947 (N_6947,N_5221,N_5449);
nand U6948 (N_6948,N_4280,N_4879);
xor U6949 (N_6949,N_4119,N_4715);
nand U6950 (N_6950,N_4230,N_5927);
nor U6951 (N_6951,N_4373,N_5147);
and U6952 (N_6952,N_5046,N_5231);
or U6953 (N_6953,N_4766,N_5059);
or U6954 (N_6954,N_4705,N_5504);
xor U6955 (N_6955,N_5435,N_4286);
and U6956 (N_6956,N_5320,N_5993);
nor U6957 (N_6957,N_5550,N_4214);
and U6958 (N_6958,N_4609,N_4384);
or U6959 (N_6959,N_4737,N_5959);
nor U6960 (N_6960,N_4247,N_4582);
nand U6961 (N_6961,N_5109,N_5038);
xor U6962 (N_6962,N_5544,N_5120);
or U6963 (N_6963,N_4875,N_5150);
nand U6964 (N_6964,N_4248,N_5373);
and U6965 (N_6965,N_4863,N_4689);
nand U6966 (N_6966,N_4342,N_4887);
and U6967 (N_6967,N_4049,N_5638);
xor U6968 (N_6968,N_4117,N_4324);
or U6969 (N_6969,N_5789,N_4152);
xor U6970 (N_6970,N_4822,N_5532);
and U6971 (N_6971,N_4416,N_5691);
and U6972 (N_6972,N_4401,N_4462);
and U6973 (N_6973,N_5342,N_4424);
or U6974 (N_6974,N_5980,N_4636);
or U6975 (N_6975,N_5827,N_5639);
and U6976 (N_6976,N_5706,N_4517);
nor U6977 (N_6977,N_4439,N_5629);
nand U6978 (N_6978,N_5631,N_4220);
nor U6979 (N_6979,N_5708,N_4093);
nor U6980 (N_6980,N_4338,N_4189);
nand U6981 (N_6981,N_4387,N_4071);
nor U6982 (N_6982,N_5906,N_4486);
xor U6983 (N_6983,N_4696,N_4826);
or U6984 (N_6984,N_5107,N_4971);
nand U6985 (N_6985,N_5556,N_4332);
nor U6986 (N_6986,N_4023,N_5864);
and U6987 (N_6987,N_4991,N_4215);
nor U6988 (N_6988,N_4583,N_5233);
xnor U6989 (N_6989,N_4962,N_4003);
nor U6990 (N_6990,N_4797,N_5184);
nor U6991 (N_6991,N_4259,N_5123);
nor U6992 (N_6992,N_4085,N_5024);
and U6993 (N_6993,N_5326,N_4353);
and U6994 (N_6994,N_5309,N_4969);
nor U6995 (N_6995,N_5612,N_4001);
and U6996 (N_6996,N_4504,N_5882);
nor U6997 (N_6997,N_5752,N_4190);
and U6998 (N_6998,N_4823,N_5832);
xnor U6999 (N_6999,N_4652,N_5517);
or U7000 (N_7000,N_4160,N_4621);
or U7001 (N_7001,N_4543,N_4633);
nand U7002 (N_7002,N_4496,N_4857);
nor U7003 (N_7003,N_5336,N_5562);
nor U7004 (N_7004,N_5638,N_4636);
and U7005 (N_7005,N_4625,N_5874);
xnor U7006 (N_7006,N_4706,N_4605);
nor U7007 (N_7007,N_5767,N_4227);
nor U7008 (N_7008,N_5061,N_5632);
nor U7009 (N_7009,N_4676,N_4456);
nand U7010 (N_7010,N_4140,N_4630);
or U7011 (N_7011,N_4792,N_4086);
and U7012 (N_7012,N_4769,N_5466);
or U7013 (N_7013,N_4916,N_5110);
xnor U7014 (N_7014,N_4487,N_5433);
or U7015 (N_7015,N_4466,N_5014);
and U7016 (N_7016,N_4544,N_4623);
and U7017 (N_7017,N_5689,N_4069);
or U7018 (N_7018,N_4723,N_4456);
or U7019 (N_7019,N_4126,N_5249);
or U7020 (N_7020,N_4948,N_4472);
nand U7021 (N_7021,N_4995,N_4762);
xnor U7022 (N_7022,N_4116,N_5930);
or U7023 (N_7023,N_5660,N_5574);
xnor U7024 (N_7024,N_5521,N_5343);
and U7025 (N_7025,N_5279,N_5899);
nor U7026 (N_7026,N_4391,N_4699);
nand U7027 (N_7027,N_5299,N_5311);
nor U7028 (N_7028,N_5887,N_5624);
xnor U7029 (N_7029,N_4583,N_4329);
nor U7030 (N_7030,N_5233,N_5911);
and U7031 (N_7031,N_5978,N_4522);
xnor U7032 (N_7032,N_5731,N_5767);
nor U7033 (N_7033,N_5098,N_5008);
nor U7034 (N_7034,N_5621,N_5937);
and U7035 (N_7035,N_5533,N_4473);
or U7036 (N_7036,N_5891,N_5000);
nor U7037 (N_7037,N_5552,N_4054);
and U7038 (N_7038,N_5956,N_5722);
nor U7039 (N_7039,N_5923,N_4706);
xor U7040 (N_7040,N_5574,N_4423);
xnor U7041 (N_7041,N_4204,N_4942);
xor U7042 (N_7042,N_4501,N_5467);
nor U7043 (N_7043,N_5858,N_5637);
xor U7044 (N_7044,N_5441,N_5555);
and U7045 (N_7045,N_5344,N_4092);
nand U7046 (N_7046,N_4560,N_5177);
or U7047 (N_7047,N_5981,N_4028);
and U7048 (N_7048,N_4039,N_4801);
xnor U7049 (N_7049,N_4133,N_5158);
or U7050 (N_7050,N_4175,N_5927);
nand U7051 (N_7051,N_5818,N_4129);
and U7052 (N_7052,N_4367,N_4574);
xor U7053 (N_7053,N_5874,N_4808);
nand U7054 (N_7054,N_5756,N_5422);
or U7055 (N_7055,N_5001,N_5091);
nor U7056 (N_7056,N_5256,N_4496);
or U7057 (N_7057,N_5230,N_5957);
nand U7058 (N_7058,N_5344,N_5916);
nand U7059 (N_7059,N_4808,N_5860);
and U7060 (N_7060,N_4158,N_5284);
and U7061 (N_7061,N_4108,N_5008);
xnor U7062 (N_7062,N_5702,N_5489);
or U7063 (N_7063,N_5949,N_4436);
or U7064 (N_7064,N_5846,N_4293);
and U7065 (N_7065,N_5991,N_5608);
xor U7066 (N_7066,N_4378,N_5771);
and U7067 (N_7067,N_4211,N_4593);
xnor U7068 (N_7068,N_5801,N_4599);
nand U7069 (N_7069,N_4042,N_5659);
nand U7070 (N_7070,N_5885,N_5106);
nand U7071 (N_7071,N_4809,N_4538);
or U7072 (N_7072,N_5633,N_5865);
nand U7073 (N_7073,N_4140,N_4214);
nor U7074 (N_7074,N_5930,N_5774);
nor U7075 (N_7075,N_5776,N_5661);
nor U7076 (N_7076,N_4875,N_5519);
xnor U7077 (N_7077,N_4897,N_5002);
xor U7078 (N_7078,N_4402,N_4406);
nor U7079 (N_7079,N_4603,N_4902);
and U7080 (N_7080,N_5341,N_4706);
nor U7081 (N_7081,N_5039,N_4955);
and U7082 (N_7082,N_5846,N_5497);
xnor U7083 (N_7083,N_5325,N_4747);
or U7084 (N_7084,N_5199,N_4347);
nor U7085 (N_7085,N_5019,N_5967);
nand U7086 (N_7086,N_4231,N_5738);
nand U7087 (N_7087,N_4257,N_5696);
nand U7088 (N_7088,N_4151,N_5129);
nor U7089 (N_7089,N_4918,N_4410);
nor U7090 (N_7090,N_5512,N_4567);
xor U7091 (N_7091,N_5709,N_4709);
and U7092 (N_7092,N_5601,N_5010);
or U7093 (N_7093,N_4342,N_5734);
xnor U7094 (N_7094,N_4933,N_5046);
xor U7095 (N_7095,N_4837,N_5417);
nand U7096 (N_7096,N_5145,N_4630);
or U7097 (N_7097,N_4999,N_5554);
and U7098 (N_7098,N_4514,N_4861);
nand U7099 (N_7099,N_5554,N_4374);
and U7100 (N_7100,N_4057,N_5419);
xnor U7101 (N_7101,N_5657,N_5624);
xor U7102 (N_7102,N_5516,N_5667);
nand U7103 (N_7103,N_5770,N_4567);
nor U7104 (N_7104,N_5702,N_5987);
or U7105 (N_7105,N_5571,N_4983);
xor U7106 (N_7106,N_4646,N_4880);
nand U7107 (N_7107,N_4430,N_4220);
nor U7108 (N_7108,N_5277,N_5165);
or U7109 (N_7109,N_5923,N_5316);
xor U7110 (N_7110,N_5132,N_5292);
nor U7111 (N_7111,N_5780,N_4199);
or U7112 (N_7112,N_5319,N_5817);
and U7113 (N_7113,N_5179,N_4957);
xnor U7114 (N_7114,N_5145,N_4545);
and U7115 (N_7115,N_5124,N_4185);
and U7116 (N_7116,N_4397,N_4919);
nand U7117 (N_7117,N_5113,N_4953);
or U7118 (N_7118,N_5702,N_4373);
and U7119 (N_7119,N_4965,N_5479);
nor U7120 (N_7120,N_4704,N_4286);
xor U7121 (N_7121,N_5746,N_4283);
xor U7122 (N_7122,N_4133,N_4086);
nand U7123 (N_7123,N_4977,N_4167);
nor U7124 (N_7124,N_4724,N_5180);
nor U7125 (N_7125,N_5458,N_4014);
nor U7126 (N_7126,N_5412,N_4660);
nor U7127 (N_7127,N_4144,N_5565);
and U7128 (N_7128,N_4143,N_5422);
xor U7129 (N_7129,N_4848,N_5050);
nand U7130 (N_7130,N_5986,N_5061);
and U7131 (N_7131,N_4211,N_5809);
nand U7132 (N_7132,N_4827,N_4209);
xor U7133 (N_7133,N_5049,N_5893);
nor U7134 (N_7134,N_5538,N_5474);
or U7135 (N_7135,N_4393,N_5644);
nand U7136 (N_7136,N_4680,N_5626);
nor U7137 (N_7137,N_5850,N_5540);
xnor U7138 (N_7138,N_4606,N_5948);
and U7139 (N_7139,N_5395,N_4491);
nor U7140 (N_7140,N_4212,N_5260);
xor U7141 (N_7141,N_5578,N_5213);
nor U7142 (N_7142,N_5884,N_5600);
and U7143 (N_7143,N_4993,N_4788);
nand U7144 (N_7144,N_4822,N_4528);
or U7145 (N_7145,N_5645,N_5094);
nand U7146 (N_7146,N_5592,N_4054);
nand U7147 (N_7147,N_5392,N_4535);
and U7148 (N_7148,N_5731,N_4915);
xnor U7149 (N_7149,N_4690,N_4590);
or U7150 (N_7150,N_4369,N_4575);
xnor U7151 (N_7151,N_4715,N_5617);
nand U7152 (N_7152,N_4411,N_5504);
or U7153 (N_7153,N_4909,N_5120);
and U7154 (N_7154,N_4958,N_4311);
nand U7155 (N_7155,N_5165,N_5416);
or U7156 (N_7156,N_5048,N_5270);
and U7157 (N_7157,N_4913,N_5909);
nand U7158 (N_7158,N_5988,N_4928);
xor U7159 (N_7159,N_4769,N_5152);
and U7160 (N_7160,N_5713,N_5181);
xnor U7161 (N_7161,N_5845,N_5041);
nor U7162 (N_7162,N_5287,N_4721);
or U7163 (N_7163,N_5360,N_4280);
or U7164 (N_7164,N_5128,N_4696);
nand U7165 (N_7165,N_5080,N_5408);
nor U7166 (N_7166,N_5777,N_5126);
xnor U7167 (N_7167,N_4041,N_5599);
and U7168 (N_7168,N_5683,N_4032);
nor U7169 (N_7169,N_5329,N_5911);
nand U7170 (N_7170,N_5480,N_4185);
nand U7171 (N_7171,N_5344,N_5729);
or U7172 (N_7172,N_5825,N_4471);
and U7173 (N_7173,N_4997,N_5854);
xnor U7174 (N_7174,N_4975,N_5812);
xnor U7175 (N_7175,N_4337,N_5067);
or U7176 (N_7176,N_5233,N_4725);
nor U7177 (N_7177,N_5754,N_5093);
nor U7178 (N_7178,N_4540,N_4430);
nor U7179 (N_7179,N_4751,N_4405);
nor U7180 (N_7180,N_4331,N_4549);
nand U7181 (N_7181,N_5256,N_5924);
nor U7182 (N_7182,N_4069,N_4609);
nand U7183 (N_7183,N_4331,N_5721);
nor U7184 (N_7184,N_5659,N_4782);
nor U7185 (N_7185,N_4815,N_4641);
or U7186 (N_7186,N_5797,N_5814);
nor U7187 (N_7187,N_5983,N_5110);
xor U7188 (N_7188,N_4297,N_5653);
and U7189 (N_7189,N_4645,N_5434);
nor U7190 (N_7190,N_5404,N_4095);
and U7191 (N_7191,N_4692,N_4842);
or U7192 (N_7192,N_4704,N_4900);
or U7193 (N_7193,N_5303,N_4093);
nand U7194 (N_7194,N_4541,N_4472);
nand U7195 (N_7195,N_5797,N_4323);
nand U7196 (N_7196,N_4092,N_5180);
nand U7197 (N_7197,N_4490,N_5017);
nand U7198 (N_7198,N_5618,N_5071);
xor U7199 (N_7199,N_4564,N_4301);
or U7200 (N_7200,N_5615,N_4912);
nor U7201 (N_7201,N_4537,N_4487);
or U7202 (N_7202,N_4120,N_4194);
nand U7203 (N_7203,N_5259,N_5786);
nor U7204 (N_7204,N_5133,N_4197);
nand U7205 (N_7205,N_4065,N_5299);
nor U7206 (N_7206,N_5305,N_5308);
xnor U7207 (N_7207,N_4431,N_5348);
xor U7208 (N_7208,N_4058,N_4141);
and U7209 (N_7209,N_5173,N_5452);
or U7210 (N_7210,N_5436,N_5625);
and U7211 (N_7211,N_5215,N_4360);
or U7212 (N_7212,N_4695,N_4064);
nor U7213 (N_7213,N_5058,N_5711);
or U7214 (N_7214,N_5873,N_5808);
xnor U7215 (N_7215,N_5782,N_4973);
or U7216 (N_7216,N_5258,N_4190);
nand U7217 (N_7217,N_4987,N_5787);
xor U7218 (N_7218,N_5330,N_5712);
nor U7219 (N_7219,N_5644,N_4161);
and U7220 (N_7220,N_4021,N_5470);
or U7221 (N_7221,N_5397,N_4720);
and U7222 (N_7222,N_4095,N_4993);
nand U7223 (N_7223,N_5317,N_5246);
nor U7224 (N_7224,N_5378,N_4622);
xnor U7225 (N_7225,N_4431,N_5012);
or U7226 (N_7226,N_5148,N_5024);
nor U7227 (N_7227,N_5141,N_4665);
and U7228 (N_7228,N_4087,N_4193);
xnor U7229 (N_7229,N_4045,N_4870);
nor U7230 (N_7230,N_4240,N_5626);
nor U7231 (N_7231,N_4536,N_4595);
and U7232 (N_7232,N_5467,N_4255);
nand U7233 (N_7233,N_5635,N_5447);
xnor U7234 (N_7234,N_4667,N_5404);
xnor U7235 (N_7235,N_4416,N_5059);
or U7236 (N_7236,N_5758,N_4370);
or U7237 (N_7237,N_5987,N_4676);
nand U7238 (N_7238,N_4582,N_4050);
or U7239 (N_7239,N_5614,N_4616);
xor U7240 (N_7240,N_4521,N_5383);
or U7241 (N_7241,N_5050,N_5659);
or U7242 (N_7242,N_5694,N_4017);
and U7243 (N_7243,N_5863,N_5041);
xnor U7244 (N_7244,N_5136,N_5780);
xor U7245 (N_7245,N_4219,N_4945);
xor U7246 (N_7246,N_5256,N_5525);
and U7247 (N_7247,N_4114,N_5241);
or U7248 (N_7248,N_5471,N_4676);
nand U7249 (N_7249,N_5832,N_5256);
and U7250 (N_7250,N_4411,N_5127);
nand U7251 (N_7251,N_4265,N_5535);
nor U7252 (N_7252,N_5305,N_4249);
xor U7253 (N_7253,N_4409,N_4966);
xor U7254 (N_7254,N_5655,N_5578);
and U7255 (N_7255,N_5575,N_4930);
nor U7256 (N_7256,N_4633,N_5030);
xor U7257 (N_7257,N_5385,N_5373);
nand U7258 (N_7258,N_5095,N_4394);
xnor U7259 (N_7259,N_5465,N_4379);
and U7260 (N_7260,N_4461,N_4469);
nand U7261 (N_7261,N_5168,N_4555);
nor U7262 (N_7262,N_5575,N_5283);
nand U7263 (N_7263,N_4501,N_4159);
or U7264 (N_7264,N_5231,N_5144);
or U7265 (N_7265,N_4717,N_5578);
and U7266 (N_7266,N_4875,N_5402);
or U7267 (N_7267,N_4804,N_5194);
xor U7268 (N_7268,N_5655,N_5621);
or U7269 (N_7269,N_4942,N_5788);
and U7270 (N_7270,N_5877,N_4893);
and U7271 (N_7271,N_5277,N_4608);
or U7272 (N_7272,N_5248,N_5723);
and U7273 (N_7273,N_4416,N_5227);
and U7274 (N_7274,N_5081,N_4048);
nor U7275 (N_7275,N_5197,N_5427);
and U7276 (N_7276,N_4904,N_4761);
nor U7277 (N_7277,N_4045,N_4768);
xnor U7278 (N_7278,N_5421,N_4955);
and U7279 (N_7279,N_4169,N_4159);
or U7280 (N_7280,N_4575,N_5600);
and U7281 (N_7281,N_4501,N_5840);
nand U7282 (N_7282,N_4605,N_4041);
or U7283 (N_7283,N_4217,N_5633);
or U7284 (N_7284,N_5112,N_5392);
nor U7285 (N_7285,N_5550,N_5177);
nor U7286 (N_7286,N_5773,N_4919);
xnor U7287 (N_7287,N_4584,N_4080);
and U7288 (N_7288,N_4793,N_4884);
nand U7289 (N_7289,N_5302,N_4444);
or U7290 (N_7290,N_4325,N_5988);
xor U7291 (N_7291,N_4721,N_5935);
nor U7292 (N_7292,N_5920,N_4237);
and U7293 (N_7293,N_4253,N_5194);
and U7294 (N_7294,N_4827,N_5584);
nor U7295 (N_7295,N_5969,N_4695);
nand U7296 (N_7296,N_5316,N_5546);
xnor U7297 (N_7297,N_5278,N_5439);
xnor U7298 (N_7298,N_4442,N_5027);
or U7299 (N_7299,N_4160,N_5308);
nand U7300 (N_7300,N_4769,N_4398);
nand U7301 (N_7301,N_4054,N_5822);
and U7302 (N_7302,N_5777,N_5631);
or U7303 (N_7303,N_5567,N_4736);
and U7304 (N_7304,N_5546,N_5614);
and U7305 (N_7305,N_5720,N_4017);
nor U7306 (N_7306,N_4698,N_4610);
nor U7307 (N_7307,N_4393,N_4811);
and U7308 (N_7308,N_5242,N_4882);
nor U7309 (N_7309,N_5678,N_5215);
or U7310 (N_7310,N_5830,N_5398);
or U7311 (N_7311,N_4611,N_4711);
and U7312 (N_7312,N_5986,N_5645);
or U7313 (N_7313,N_4293,N_5667);
and U7314 (N_7314,N_4195,N_4461);
nand U7315 (N_7315,N_4747,N_4477);
nor U7316 (N_7316,N_4680,N_4856);
or U7317 (N_7317,N_4266,N_4255);
and U7318 (N_7318,N_4280,N_4983);
nand U7319 (N_7319,N_4986,N_5304);
or U7320 (N_7320,N_5583,N_4407);
or U7321 (N_7321,N_4665,N_4754);
xnor U7322 (N_7322,N_5814,N_5860);
or U7323 (N_7323,N_5944,N_4637);
and U7324 (N_7324,N_4416,N_5895);
and U7325 (N_7325,N_4785,N_5325);
and U7326 (N_7326,N_4638,N_4516);
nor U7327 (N_7327,N_4553,N_4537);
xor U7328 (N_7328,N_5805,N_5654);
nand U7329 (N_7329,N_5860,N_5545);
nand U7330 (N_7330,N_4142,N_5502);
and U7331 (N_7331,N_4694,N_5622);
or U7332 (N_7332,N_5614,N_4550);
nand U7333 (N_7333,N_5078,N_4716);
nand U7334 (N_7334,N_4992,N_5911);
nand U7335 (N_7335,N_4872,N_5705);
nand U7336 (N_7336,N_4937,N_4423);
and U7337 (N_7337,N_4977,N_5371);
nand U7338 (N_7338,N_4648,N_4760);
xnor U7339 (N_7339,N_4028,N_5713);
xor U7340 (N_7340,N_5965,N_5843);
nor U7341 (N_7341,N_5089,N_5018);
nand U7342 (N_7342,N_4229,N_4601);
nand U7343 (N_7343,N_4439,N_5319);
and U7344 (N_7344,N_5985,N_4470);
xnor U7345 (N_7345,N_4115,N_5633);
and U7346 (N_7346,N_5676,N_5412);
nand U7347 (N_7347,N_5484,N_4675);
nor U7348 (N_7348,N_4488,N_4644);
xnor U7349 (N_7349,N_5592,N_5877);
and U7350 (N_7350,N_5859,N_4663);
and U7351 (N_7351,N_4414,N_4921);
xor U7352 (N_7352,N_4529,N_4203);
or U7353 (N_7353,N_5205,N_5124);
and U7354 (N_7354,N_4978,N_5330);
nor U7355 (N_7355,N_4744,N_5092);
nor U7356 (N_7356,N_5722,N_5206);
nand U7357 (N_7357,N_5743,N_5127);
nand U7358 (N_7358,N_4657,N_4918);
xnor U7359 (N_7359,N_5304,N_4305);
nor U7360 (N_7360,N_5461,N_4030);
and U7361 (N_7361,N_4494,N_4717);
xor U7362 (N_7362,N_5561,N_4002);
or U7363 (N_7363,N_4120,N_4650);
or U7364 (N_7364,N_5154,N_4149);
xor U7365 (N_7365,N_5453,N_4512);
or U7366 (N_7366,N_5698,N_4337);
nand U7367 (N_7367,N_4810,N_5416);
and U7368 (N_7368,N_5585,N_5182);
nor U7369 (N_7369,N_4983,N_5151);
and U7370 (N_7370,N_4195,N_4525);
xor U7371 (N_7371,N_4720,N_5163);
nand U7372 (N_7372,N_4489,N_5653);
and U7373 (N_7373,N_5673,N_5127);
nor U7374 (N_7374,N_5061,N_4695);
nor U7375 (N_7375,N_4820,N_5311);
nor U7376 (N_7376,N_4635,N_4243);
nand U7377 (N_7377,N_5831,N_5084);
or U7378 (N_7378,N_5162,N_5108);
and U7379 (N_7379,N_5909,N_4188);
or U7380 (N_7380,N_4176,N_5587);
xor U7381 (N_7381,N_5483,N_4173);
or U7382 (N_7382,N_5072,N_5294);
nor U7383 (N_7383,N_4795,N_5829);
or U7384 (N_7384,N_5178,N_4204);
xnor U7385 (N_7385,N_5076,N_5655);
and U7386 (N_7386,N_4217,N_4293);
and U7387 (N_7387,N_4880,N_5098);
nand U7388 (N_7388,N_5751,N_4574);
and U7389 (N_7389,N_4026,N_4998);
and U7390 (N_7390,N_4592,N_5380);
and U7391 (N_7391,N_4150,N_4788);
nor U7392 (N_7392,N_4929,N_5019);
and U7393 (N_7393,N_4759,N_5118);
and U7394 (N_7394,N_5677,N_5722);
xnor U7395 (N_7395,N_5368,N_5478);
nor U7396 (N_7396,N_5668,N_5359);
nor U7397 (N_7397,N_5796,N_4611);
nand U7398 (N_7398,N_4113,N_5410);
and U7399 (N_7399,N_4999,N_5334);
and U7400 (N_7400,N_4281,N_5731);
and U7401 (N_7401,N_4593,N_5032);
and U7402 (N_7402,N_5611,N_5196);
and U7403 (N_7403,N_4715,N_4381);
or U7404 (N_7404,N_4582,N_4070);
xor U7405 (N_7405,N_5561,N_5478);
nor U7406 (N_7406,N_4757,N_4811);
or U7407 (N_7407,N_4921,N_5576);
and U7408 (N_7408,N_5774,N_4536);
nor U7409 (N_7409,N_5440,N_4314);
or U7410 (N_7410,N_4032,N_4192);
or U7411 (N_7411,N_4698,N_4281);
xnor U7412 (N_7412,N_4864,N_4935);
or U7413 (N_7413,N_5413,N_5156);
xor U7414 (N_7414,N_5275,N_5515);
and U7415 (N_7415,N_5708,N_4468);
xor U7416 (N_7416,N_5172,N_5144);
nand U7417 (N_7417,N_4078,N_4285);
and U7418 (N_7418,N_5251,N_4521);
nor U7419 (N_7419,N_4813,N_4931);
xor U7420 (N_7420,N_4413,N_5503);
or U7421 (N_7421,N_5234,N_4915);
nand U7422 (N_7422,N_4194,N_4487);
xnor U7423 (N_7423,N_4657,N_4385);
or U7424 (N_7424,N_4866,N_4401);
nand U7425 (N_7425,N_5091,N_5158);
and U7426 (N_7426,N_4037,N_5864);
xor U7427 (N_7427,N_4419,N_4621);
nand U7428 (N_7428,N_4643,N_5297);
nor U7429 (N_7429,N_4721,N_5658);
or U7430 (N_7430,N_4526,N_4428);
nor U7431 (N_7431,N_5506,N_5029);
nand U7432 (N_7432,N_5383,N_5044);
or U7433 (N_7433,N_4301,N_5039);
nand U7434 (N_7434,N_4156,N_4830);
or U7435 (N_7435,N_4794,N_4435);
or U7436 (N_7436,N_4579,N_5324);
and U7437 (N_7437,N_4650,N_4994);
nand U7438 (N_7438,N_4182,N_4672);
xor U7439 (N_7439,N_4902,N_4006);
and U7440 (N_7440,N_4590,N_4329);
and U7441 (N_7441,N_4219,N_5513);
nand U7442 (N_7442,N_4477,N_4416);
xnor U7443 (N_7443,N_4831,N_4948);
and U7444 (N_7444,N_5423,N_5575);
xnor U7445 (N_7445,N_4662,N_5186);
and U7446 (N_7446,N_5887,N_5275);
or U7447 (N_7447,N_5525,N_5135);
nand U7448 (N_7448,N_5669,N_5889);
xor U7449 (N_7449,N_4713,N_5683);
nand U7450 (N_7450,N_5909,N_4874);
and U7451 (N_7451,N_4683,N_5427);
nor U7452 (N_7452,N_4168,N_4056);
nand U7453 (N_7453,N_4872,N_5151);
and U7454 (N_7454,N_5888,N_4562);
xnor U7455 (N_7455,N_5805,N_5407);
xnor U7456 (N_7456,N_5737,N_5960);
nand U7457 (N_7457,N_5092,N_5208);
and U7458 (N_7458,N_4056,N_4719);
and U7459 (N_7459,N_5590,N_5819);
or U7460 (N_7460,N_4975,N_4430);
nand U7461 (N_7461,N_4692,N_4753);
xnor U7462 (N_7462,N_4639,N_5928);
or U7463 (N_7463,N_4679,N_4275);
nand U7464 (N_7464,N_4847,N_5244);
xnor U7465 (N_7465,N_4688,N_4975);
xnor U7466 (N_7466,N_4672,N_5422);
or U7467 (N_7467,N_5065,N_4028);
nand U7468 (N_7468,N_5860,N_5799);
xnor U7469 (N_7469,N_5947,N_5279);
xor U7470 (N_7470,N_4413,N_5094);
xor U7471 (N_7471,N_5012,N_4666);
nand U7472 (N_7472,N_5563,N_5463);
or U7473 (N_7473,N_5732,N_4982);
nor U7474 (N_7474,N_4243,N_5284);
nor U7475 (N_7475,N_4752,N_5755);
xor U7476 (N_7476,N_5502,N_4411);
nor U7477 (N_7477,N_5865,N_4013);
or U7478 (N_7478,N_4174,N_4760);
nand U7479 (N_7479,N_4446,N_5078);
or U7480 (N_7480,N_4993,N_4470);
xnor U7481 (N_7481,N_4491,N_5512);
and U7482 (N_7482,N_4179,N_4227);
nor U7483 (N_7483,N_5686,N_5918);
nand U7484 (N_7484,N_4234,N_5275);
nand U7485 (N_7485,N_5654,N_5771);
or U7486 (N_7486,N_5785,N_5302);
or U7487 (N_7487,N_5280,N_4277);
and U7488 (N_7488,N_5654,N_5385);
or U7489 (N_7489,N_4222,N_4015);
nand U7490 (N_7490,N_4534,N_5650);
xnor U7491 (N_7491,N_4295,N_4893);
and U7492 (N_7492,N_4006,N_5436);
xnor U7493 (N_7493,N_4408,N_5183);
nor U7494 (N_7494,N_5164,N_5550);
and U7495 (N_7495,N_4970,N_4646);
or U7496 (N_7496,N_4825,N_4651);
nor U7497 (N_7497,N_4858,N_4604);
nand U7498 (N_7498,N_5653,N_5416);
or U7499 (N_7499,N_5926,N_5860);
and U7500 (N_7500,N_4592,N_5985);
and U7501 (N_7501,N_4352,N_4161);
and U7502 (N_7502,N_5666,N_5477);
or U7503 (N_7503,N_5216,N_4074);
and U7504 (N_7504,N_4319,N_5028);
and U7505 (N_7505,N_4306,N_5685);
xnor U7506 (N_7506,N_5601,N_4884);
and U7507 (N_7507,N_5389,N_5816);
and U7508 (N_7508,N_4625,N_5562);
xor U7509 (N_7509,N_5498,N_5126);
or U7510 (N_7510,N_4683,N_4548);
nor U7511 (N_7511,N_5242,N_4026);
xnor U7512 (N_7512,N_5328,N_4803);
nor U7513 (N_7513,N_5165,N_5438);
or U7514 (N_7514,N_5664,N_5858);
or U7515 (N_7515,N_4907,N_4245);
and U7516 (N_7516,N_5640,N_5201);
xnor U7517 (N_7517,N_4929,N_5322);
xnor U7518 (N_7518,N_4543,N_4389);
and U7519 (N_7519,N_5740,N_4343);
and U7520 (N_7520,N_5992,N_4853);
or U7521 (N_7521,N_5564,N_5125);
and U7522 (N_7522,N_4655,N_4562);
xor U7523 (N_7523,N_4100,N_5049);
or U7524 (N_7524,N_5701,N_4566);
nor U7525 (N_7525,N_4523,N_5413);
xor U7526 (N_7526,N_4278,N_5378);
nand U7527 (N_7527,N_4742,N_4305);
nor U7528 (N_7528,N_5167,N_4635);
and U7529 (N_7529,N_4293,N_4052);
nor U7530 (N_7530,N_4533,N_4406);
or U7531 (N_7531,N_5519,N_4174);
or U7532 (N_7532,N_4217,N_5403);
xor U7533 (N_7533,N_5310,N_4663);
xor U7534 (N_7534,N_4853,N_5467);
xor U7535 (N_7535,N_4327,N_5911);
nor U7536 (N_7536,N_5722,N_5272);
nor U7537 (N_7537,N_4604,N_4370);
or U7538 (N_7538,N_5946,N_5854);
xor U7539 (N_7539,N_5531,N_4664);
xnor U7540 (N_7540,N_5331,N_5198);
or U7541 (N_7541,N_5269,N_5945);
nor U7542 (N_7542,N_5684,N_4160);
and U7543 (N_7543,N_4113,N_4555);
nor U7544 (N_7544,N_4710,N_4232);
nor U7545 (N_7545,N_5432,N_4332);
nand U7546 (N_7546,N_5005,N_4613);
or U7547 (N_7547,N_4078,N_5613);
nand U7548 (N_7548,N_4398,N_4334);
or U7549 (N_7549,N_5065,N_4126);
xor U7550 (N_7550,N_4014,N_5707);
or U7551 (N_7551,N_4649,N_4250);
or U7552 (N_7552,N_4960,N_4836);
and U7553 (N_7553,N_5997,N_4845);
xor U7554 (N_7554,N_5335,N_4336);
or U7555 (N_7555,N_5788,N_5044);
or U7556 (N_7556,N_4347,N_5470);
nand U7557 (N_7557,N_5179,N_5415);
xor U7558 (N_7558,N_4565,N_4729);
and U7559 (N_7559,N_5496,N_4849);
nand U7560 (N_7560,N_5806,N_5239);
or U7561 (N_7561,N_5846,N_5078);
xnor U7562 (N_7562,N_5481,N_5466);
and U7563 (N_7563,N_4028,N_5690);
and U7564 (N_7564,N_4465,N_5435);
xnor U7565 (N_7565,N_4750,N_4252);
nand U7566 (N_7566,N_4060,N_4945);
xor U7567 (N_7567,N_4166,N_4721);
and U7568 (N_7568,N_4352,N_5771);
nand U7569 (N_7569,N_4557,N_4627);
xor U7570 (N_7570,N_4894,N_5722);
and U7571 (N_7571,N_5257,N_4081);
and U7572 (N_7572,N_4390,N_4914);
or U7573 (N_7573,N_5193,N_5612);
nor U7574 (N_7574,N_5884,N_5151);
or U7575 (N_7575,N_4518,N_5457);
and U7576 (N_7576,N_4139,N_5584);
nand U7577 (N_7577,N_5256,N_5646);
nor U7578 (N_7578,N_5585,N_4820);
nor U7579 (N_7579,N_5088,N_5071);
or U7580 (N_7580,N_4043,N_4105);
and U7581 (N_7581,N_5210,N_4341);
and U7582 (N_7582,N_4606,N_4538);
xor U7583 (N_7583,N_5391,N_5436);
or U7584 (N_7584,N_5772,N_5774);
nand U7585 (N_7585,N_4674,N_5343);
nor U7586 (N_7586,N_5214,N_4070);
or U7587 (N_7587,N_4291,N_4414);
and U7588 (N_7588,N_5856,N_4620);
nand U7589 (N_7589,N_4825,N_4729);
nor U7590 (N_7590,N_4358,N_4662);
xnor U7591 (N_7591,N_5084,N_5111);
and U7592 (N_7592,N_5708,N_4325);
and U7593 (N_7593,N_4600,N_4338);
nor U7594 (N_7594,N_5862,N_4479);
or U7595 (N_7595,N_5922,N_5916);
and U7596 (N_7596,N_5121,N_5409);
nor U7597 (N_7597,N_5242,N_4140);
and U7598 (N_7598,N_5682,N_5578);
and U7599 (N_7599,N_5446,N_4308);
xnor U7600 (N_7600,N_4286,N_5115);
nor U7601 (N_7601,N_5861,N_5310);
and U7602 (N_7602,N_5561,N_4354);
nand U7603 (N_7603,N_4053,N_5265);
xnor U7604 (N_7604,N_4516,N_5277);
or U7605 (N_7605,N_4925,N_4118);
nand U7606 (N_7606,N_5882,N_5104);
or U7607 (N_7607,N_4394,N_5821);
xor U7608 (N_7608,N_5945,N_4601);
or U7609 (N_7609,N_4319,N_5388);
xnor U7610 (N_7610,N_4085,N_5732);
and U7611 (N_7611,N_5696,N_4566);
or U7612 (N_7612,N_4020,N_4693);
and U7613 (N_7613,N_5117,N_5914);
nor U7614 (N_7614,N_5916,N_4851);
nand U7615 (N_7615,N_5262,N_5794);
xnor U7616 (N_7616,N_5363,N_4100);
nand U7617 (N_7617,N_4946,N_5268);
nand U7618 (N_7618,N_5287,N_4541);
nand U7619 (N_7619,N_4530,N_5188);
nand U7620 (N_7620,N_4516,N_5451);
nand U7621 (N_7621,N_4429,N_5514);
or U7622 (N_7622,N_4185,N_4876);
nor U7623 (N_7623,N_4040,N_5002);
and U7624 (N_7624,N_5016,N_4308);
nor U7625 (N_7625,N_5490,N_5596);
nand U7626 (N_7626,N_5385,N_5280);
nand U7627 (N_7627,N_5876,N_4572);
nor U7628 (N_7628,N_4472,N_5395);
or U7629 (N_7629,N_5073,N_5098);
nor U7630 (N_7630,N_5115,N_4703);
or U7631 (N_7631,N_4908,N_5592);
and U7632 (N_7632,N_5693,N_5117);
or U7633 (N_7633,N_5998,N_4193);
or U7634 (N_7634,N_4284,N_4007);
nand U7635 (N_7635,N_5777,N_4856);
and U7636 (N_7636,N_4581,N_5207);
or U7637 (N_7637,N_4442,N_4777);
nor U7638 (N_7638,N_4009,N_4357);
nand U7639 (N_7639,N_4455,N_4888);
xor U7640 (N_7640,N_4046,N_4736);
and U7641 (N_7641,N_5709,N_4626);
xnor U7642 (N_7642,N_5345,N_4611);
nand U7643 (N_7643,N_5110,N_5241);
nor U7644 (N_7644,N_5375,N_5585);
nand U7645 (N_7645,N_4778,N_4501);
nor U7646 (N_7646,N_4363,N_5707);
or U7647 (N_7647,N_5733,N_4906);
xnor U7648 (N_7648,N_5328,N_5636);
and U7649 (N_7649,N_5831,N_4847);
nor U7650 (N_7650,N_4480,N_4874);
nor U7651 (N_7651,N_5114,N_4591);
nor U7652 (N_7652,N_5240,N_5916);
and U7653 (N_7653,N_4805,N_4671);
nand U7654 (N_7654,N_4174,N_5839);
or U7655 (N_7655,N_4195,N_4886);
nor U7656 (N_7656,N_5166,N_4492);
and U7657 (N_7657,N_4406,N_5889);
nor U7658 (N_7658,N_5822,N_5235);
and U7659 (N_7659,N_4536,N_4408);
nor U7660 (N_7660,N_5513,N_4172);
nor U7661 (N_7661,N_5462,N_5808);
xor U7662 (N_7662,N_5757,N_4227);
or U7663 (N_7663,N_5216,N_5053);
xnor U7664 (N_7664,N_4869,N_5654);
xnor U7665 (N_7665,N_5783,N_4509);
xor U7666 (N_7666,N_5649,N_5431);
xor U7667 (N_7667,N_4590,N_5484);
and U7668 (N_7668,N_5951,N_4521);
nor U7669 (N_7669,N_5759,N_5879);
nor U7670 (N_7670,N_4362,N_5113);
or U7671 (N_7671,N_5047,N_4222);
and U7672 (N_7672,N_4559,N_4450);
and U7673 (N_7673,N_5209,N_4787);
and U7674 (N_7674,N_4416,N_4580);
xnor U7675 (N_7675,N_5528,N_4479);
or U7676 (N_7676,N_5649,N_4512);
nand U7677 (N_7677,N_5755,N_5844);
nand U7678 (N_7678,N_5486,N_4505);
nor U7679 (N_7679,N_4617,N_5324);
or U7680 (N_7680,N_5312,N_4806);
xor U7681 (N_7681,N_4133,N_4082);
nor U7682 (N_7682,N_4139,N_5988);
xnor U7683 (N_7683,N_5851,N_5736);
nor U7684 (N_7684,N_5642,N_4713);
xnor U7685 (N_7685,N_5694,N_5012);
and U7686 (N_7686,N_5032,N_4384);
nand U7687 (N_7687,N_4961,N_5520);
nand U7688 (N_7688,N_4840,N_4218);
or U7689 (N_7689,N_5159,N_4064);
xnor U7690 (N_7690,N_4999,N_4274);
nor U7691 (N_7691,N_4255,N_5348);
nand U7692 (N_7692,N_4709,N_5355);
and U7693 (N_7693,N_4287,N_5745);
nand U7694 (N_7694,N_4762,N_5806);
xor U7695 (N_7695,N_5217,N_4598);
or U7696 (N_7696,N_5828,N_4266);
or U7697 (N_7697,N_5453,N_4950);
and U7698 (N_7698,N_4722,N_5671);
xor U7699 (N_7699,N_4787,N_5271);
or U7700 (N_7700,N_5189,N_4215);
xnor U7701 (N_7701,N_5219,N_4340);
and U7702 (N_7702,N_4434,N_4424);
nor U7703 (N_7703,N_5211,N_4701);
xor U7704 (N_7704,N_4571,N_4039);
nand U7705 (N_7705,N_5246,N_4917);
and U7706 (N_7706,N_4574,N_5955);
xnor U7707 (N_7707,N_4618,N_5302);
nor U7708 (N_7708,N_5346,N_4213);
nand U7709 (N_7709,N_5689,N_5972);
or U7710 (N_7710,N_5646,N_4775);
nor U7711 (N_7711,N_5710,N_5016);
nand U7712 (N_7712,N_4888,N_4714);
or U7713 (N_7713,N_4412,N_5843);
nand U7714 (N_7714,N_4533,N_4117);
xnor U7715 (N_7715,N_5634,N_5690);
and U7716 (N_7716,N_4110,N_5367);
nand U7717 (N_7717,N_4832,N_5182);
or U7718 (N_7718,N_4202,N_4365);
nor U7719 (N_7719,N_5582,N_4154);
nor U7720 (N_7720,N_4192,N_4525);
xnor U7721 (N_7721,N_4427,N_4217);
xor U7722 (N_7722,N_5203,N_5314);
nor U7723 (N_7723,N_4842,N_4998);
nor U7724 (N_7724,N_5301,N_5669);
or U7725 (N_7725,N_4559,N_4391);
nor U7726 (N_7726,N_4456,N_4523);
nor U7727 (N_7727,N_5567,N_4871);
or U7728 (N_7728,N_4911,N_4298);
and U7729 (N_7729,N_5778,N_4838);
nor U7730 (N_7730,N_5231,N_5618);
nor U7731 (N_7731,N_5285,N_4413);
nand U7732 (N_7732,N_5604,N_5751);
or U7733 (N_7733,N_4945,N_5764);
xor U7734 (N_7734,N_4970,N_4114);
nor U7735 (N_7735,N_5987,N_5904);
or U7736 (N_7736,N_4153,N_4137);
or U7737 (N_7737,N_4244,N_5711);
nor U7738 (N_7738,N_5384,N_5032);
or U7739 (N_7739,N_5690,N_5458);
xor U7740 (N_7740,N_5697,N_4023);
or U7741 (N_7741,N_4799,N_4897);
and U7742 (N_7742,N_5773,N_4550);
and U7743 (N_7743,N_4575,N_4165);
and U7744 (N_7744,N_5646,N_5142);
or U7745 (N_7745,N_5654,N_5932);
and U7746 (N_7746,N_4658,N_5195);
nand U7747 (N_7747,N_5405,N_4337);
or U7748 (N_7748,N_4477,N_4489);
nor U7749 (N_7749,N_4395,N_5804);
nand U7750 (N_7750,N_5717,N_5518);
xnor U7751 (N_7751,N_4582,N_4897);
nand U7752 (N_7752,N_5260,N_5045);
xnor U7753 (N_7753,N_4146,N_4768);
nand U7754 (N_7754,N_5712,N_4531);
nand U7755 (N_7755,N_4739,N_4250);
nor U7756 (N_7756,N_5162,N_5886);
nand U7757 (N_7757,N_4953,N_4800);
xor U7758 (N_7758,N_5325,N_4461);
nor U7759 (N_7759,N_5887,N_4140);
nor U7760 (N_7760,N_5587,N_5241);
nor U7761 (N_7761,N_5287,N_5717);
or U7762 (N_7762,N_5388,N_5365);
and U7763 (N_7763,N_4878,N_4322);
nor U7764 (N_7764,N_4769,N_4385);
nand U7765 (N_7765,N_5141,N_4109);
xnor U7766 (N_7766,N_5947,N_4043);
or U7767 (N_7767,N_5601,N_5551);
xor U7768 (N_7768,N_4265,N_4402);
or U7769 (N_7769,N_4985,N_5155);
xnor U7770 (N_7770,N_4781,N_4700);
or U7771 (N_7771,N_4286,N_4048);
xor U7772 (N_7772,N_4023,N_4518);
and U7773 (N_7773,N_5360,N_4890);
and U7774 (N_7774,N_5904,N_4380);
and U7775 (N_7775,N_5755,N_5156);
nor U7776 (N_7776,N_5589,N_4002);
xor U7777 (N_7777,N_5577,N_5960);
xor U7778 (N_7778,N_5371,N_5614);
nor U7779 (N_7779,N_5655,N_5707);
nor U7780 (N_7780,N_4593,N_5368);
nand U7781 (N_7781,N_4539,N_5242);
nand U7782 (N_7782,N_4066,N_5376);
nor U7783 (N_7783,N_4501,N_4635);
xor U7784 (N_7784,N_4054,N_4680);
nand U7785 (N_7785,N_5488,N_4548);
or U7786 (N_7786,N_5212,N_5625);
and U7787 (N_7787,N_5191,N_4862);
nand U7788 (N_7788,N_4336,N_5040);
and U7789 (N_7789,N_5355,N_4561);
and U7790 (N_7790,N_5945,N_5657);
and U7791 (N_7791,N_4466,N_4341);
or U7792 (N_7792,N_4522,N_5352);
xor U7793 (N_7793,N_5280,N_4973);
or U7794 (N_7794,N_5513,N_5363);
xor U7795 (N_7795,N_4733,N_4399);
nor U7796 (N_7796,N_4695,N_4667);
and U7797 (N_7797,N_4118,N_5797);
xnor U7798 (N_7798,N_5489,N_4069);
nor U7799 (N_7799,N_4288,N_4603);
nand U7800 (N_7800,N_4197,N_5142);
and U7801 (N_7801,N_5518,N_4360);
nor U7802 (N_7802,N_4376,N_4459);
or U7803 (N_7803,N_4285,N_4652);
nand U7804 (N_7804,N_4859,N_4760);
nand U7805 (N_7805,N_4306,N_5420);
and U7806 (N_7806,N_4066,N_4418);
nor U7807 (N_7807,N_4471,N_4722);
xor U7808 (N_7808,N_5646,N_5271);
and U7809 (N_7809,N_4015,N_5643);
xor U7810 (N_7810,N_5509,N_5566);
or U7811 (N_7811,N_5482,N_4361);
nand U7812 (N_7812,N_5010,N_4963);
nand U7813 (N_7813,N_5678,N_4977);
and U7814 (N_7814,N_4633,N_4713);
and U7815 (N_7815,N_5263,N_5422);
nor U7816 (N_7816,N_4646,N_5708);
nor U7817 (N_7817,N_5567,N_4495);
or U7818 (N_7818,N_5036,N_4135);
nand U7819 (N_7819,N_4502,N_5580);
xor U7820 (N_7820,N_5983,N_5840);
nor U7821 (N_7821,N_4352,N_5595);
xor U7822 (N_7822,N_5044,N_4123);
nor U7823 (N_7823,N_4905,N_4833);
nor U7824 (N_7824,N_4090,N_4646);
nand U7825 (N_7825,N_4920,N_4721);
and U7826 (N_7826,N_4334,N_5899);
nand U7827 (N_7827,N_4021,N_4653);
nor U7828 (N_7828,N_5855,N_4821);
or U7829 (N_7829,N_4870,N_5434);
and U7830 (N_7830,N_4445,N_4118);
and U7831 (N_7831,N_4444,N_5748);
nand U7832 (N_7832,N_5598,N_5129);
or U7833 (N_7833,N_5685,N_4848);
and U7834 (N_7834,N_5413,N_5919);
and U7835 (N_7835,N_5320,N_5599);
xor U7836 (N_7836,N_4889,N_4273);
nor U7837 (N_7837,N_4443,N_4714);
and U7838 (N_7838,N_4616,N_4447);
nor U7839 (N_7839,N_5326,N_5271);
or U7840 (N_7840,N_5521,N_5880);
xnor U7841 (N_7841,N_4684,N_4157);
nor U7842 (N_7842,N_5922,N_5343);
and U7843 (N_7843,N_5050,N_4645);
nand U7844 (N_7844,N_5619,N_4457);
or U7845 (N_7845,N_4204,N_5298);
or U7846 (N_7846,N_5627,N_4461);
and U7847 (N_7847,N_4428,N_4619);
and U7848 (N_7848,N_5283,N_4948);
nor U7849 (N_7849,N_5877,N_4984);
xor U7850 (N_7850,N_5111,N_5471);
and U7851 (N_7851,N_5683,N_5750);
nor U7852 (N_7852,N_5533,N_5982);
nor U7853 (N_7853,N_4286,N_4202);
xnor U7854 (N_7854,N_5410,N_5503);
or U7855 (N_7855,N_4017,N_4335);
and U7856 (N_7856,N_4541,N_4129);
or U7857 (N_7857,N_4321,N_5784);
or U7858 (N_7858,N_5086,N_4981);
and U7859 (N_7859,N_4014,N_5887);
and U7860 (N_7860,N_4525,N_4537);
or U7861 (N_7861,N_4836,N_5065);
nand U7862 (N_7862,N_5366,N_4632);
xnor U7863 (N_7863,N_5582,N_4086);
nand U7864 (N_7864,N_5164,N_4449);
nand U7865 (N_7865,N_4302,N_5539);
nand U7866 (N_7866,N_5563,N_4528);
nor U7867 (N_7867,N_5541,N_5143);
nand U7868 (N_7868,N_4402,N_4565);
nand U7869 (N_7869,N_5996,N_4445);
and U7870 (N_7870,N_5724,N_4706);
nand U7871 (N_7871,N_5058,N_5189);
or U7872 (N_7872,N_5185,N_5458);
and U7873 (N_7873,N_5926,N_4134);
nor U7874 (N_7874,N_4318,N_5205);
nor U7875 (N_7875,N_4358,N_5383);
nor U7876 (N_7876,N_5979,N_4578);
xor U7877 (N_7877,N_4591,N_5685);
xor U7878 (N_7878,N_5878,N_5552);
and U7879 (N_7879,N_4777,N_4375);
nor U7880 (N_7880,N_4052,N_5946);
xnor U7881 (N_7881,N_4623,N_5474);
nand U7882 (N_7882,N_5157,N_4746);
nor U7883 (N_7883,N_5547,N_5814);
nor U7884 (N_7884,N_4384,N_4699);
nor U7885 (N_7885,N_5732,N_5009);
or U7886 (N_7886,N_5034,N_5992);
and U7887 (N_7887,N_5281,N_4224);
or U7888 (N_7888,N_5805,N_4709);
xor U7889 (N_7889,N_4177,N_4173);
nor U7890 (N_7890,N_5424,N_5876);
nor U7891 (N_7891,N_5146,N_4306);
or U7892 (N_7892,N_5241,N_4608);
nor U7893 (N_7893,N_4242,N_4412);
or U7894 (N_7894,N_5867,N_5185);
nor U7895 (N_7895,N_5505,N_4853);
nand U7896 (N_7896,N_5304,N_4960);
and U7897 (N_7897,N_5193,N_4499);
nand U7898 (N_7898,N_5759,N_5034);
or U7899 (N_7899,N_5908,N_4202);
or U7900 (N_7900,N_5383,N_5226);
nor U7901 (N_7901,N_4240,N_5383);
and U7902 (N_7902,N_5087,N_4191);
xnor U7903 (N_7903,N_4487,N_5795);
or U7904 (N_7904,N_5427,N_5454);
and U7905 (N_7905,N_4306,N_5319);
and U7906 (N_7906,N_5194,N_4070);
nand U7907 (N_7907,N_5364,N_5846);
xnor U7908 (N_7908,N_4830,N_5750);
nor U7909 (N_7909,N_4887,N_5067);
and U7910 (N_7910,N_4113,N_4756);
xnor U7911 (N_7911,N_5675,N_5753);
and U7912 (N_7912,N_5338,N_5285);
nor U7913 (N_7913,N_5637,N_5653);
or U7914 (N_7914,N_5193,N_5706);
nand U7915 (N_7915,N_4176,N_4813);
or U7916 (N_7916,N_5985,N_4362);
xnor U7917 (N_7917,N_5847,N_5934);
and U7918 (N_7918,N_4654,N_5414);
xnor U7919 (N_7919,N_4678,N_4644);
and U7920 (N_7920,N_4154,N_4888);
nor U7921 (N_7921,N_5830,N_4385);
xnor U7922 (N_7922,N_5242,N_5889);
or U7923 (N_7923,N_4523,N_5050);
nor U7924 (N_7924,N_5622,N_5395);
nor U7925 (N_7925,N_5588,N_5353);
xor U7926 (N_7926,N_5409,N_4136);
and U7927 (N_7927,N_5121,N_5231);
and U7928 (N_7928,N_4755,N_5376);
or U7929 (N_7929,N_4133,N_4247);
xor U7930 (N_7930,N_5063,N_4601);
xor U7931 (N_7931,N_4844,N_5758);
or U7932 (N_7932,N_5008,N_4842);
or U7933 (N_7933,N_4404,N_5344);
xor U7934 (N_7934,N_5675,N_5886);
nor U7935 (N_7935,N_5964,N_5982);
xnor U7936 (N_7936,N_5728,N_5304);
nand U7937 (N_7937,N_4073,N_4605);
xor U7938 (N_7938,N_4649,N_5988);
and U7939 (N_7939,N_4161,N_5578);
or U7940 (N_7940,N_5220,N_5991);
nor U7941 (N_7941,N_5987,N_4788);
nand U7942 (N_7942,N_4161,N_4240);
or U7943 (N_7943,N_5621,N_4310);
and U7944 (N_7944,N_5118,N_5123);
nand U7945 (N_7945,N_5280,N_4838);
or U7946 (N_7946,N_4979,N_5102);
nand U7947 (N_7947,N_4350,N_4058);
xnor U7948 (N_7948,N_5553,N_4635);
xnor U7949 (N_7949,N_4997,N_5721);
xor U7950 (N_7950,N_4558,N_5245);
or U7951 (N_7951,N_5078,N_4156);
or U7952 (N_7952,N_5730,N_5717);
nand U7953 (N_7953,N_4037,N_5972);
xor U7954 (N_7954,N_5411,N_5269);
or U7955 (N_7955,N_5790,N_5489);
nand U7956 (N_7956,N_5123,N_4780);
or U7957 (N_7957,N_5084,N_4694);
nand U7958 (N_7958,N_4490,N_4037);
or U7959 (N_7959,N_5594,N_5116);
and U7960 (N_7960,N_4709,N_5229);
nor U7961 (N_7961,N_4138,N_5644);
xnor U7962 (N_7962,N_5372,N_5080);
nand U7963 (N_7963,N_4168,N_5740);
or U7964 (N_7964,N_5519,N_5919);
and U7965 (N_7965,N_5392,N_5380);
nand U7966 (N_7966,N_5026,N_5225);
and U7967 (N_7967,N_4716,N_4492);
xnor U7968 (N_7968,N_4149,N_4290);
nand U7969 (N_7969,N_5992,N_5813);
nor U7970 (N_7970,N_5530,N_5888);
nor U7971 (N_7971,N_5876,N_5079);
nand U7972 (N_7972,N_4074,N_4501);
xnor U7973 (N_7973,N_4997,N_4426);
nor U7974 (N_7974,N_4904,N_4812);
xnor U7975 (N_7975,N_5421,N_5459);
and U7976 (N_7976,N_5152,N_5913);
xnor U7977 (N_7977,N_4343,N_5284);
and U7978 (N_7978,N_5393,N_4833);
nand U7979 (N_7979,N_4427,N_4073);
nor U7980 (N_7980,N_4820,N_4694);
and U7981 (N_7981,N_5795,N_4324);
nor U7982 (N_7982,N_4865,N_5110);
and U7983 (N_7983,N_5415,N_5387);
xnor U7984 (N_7984,N_5037,N_4659);
nor U7985 (N_7985,N_5637,N_5497);
xnor U7986 (N_7986,N_5172,N_5353);
or U7987 (N_7987,N_4590,N_4077);
or U7988 (N_7988,N_5362,N_4725);
nor U7989 (N_7989,N_5532,N_5104);
nand U7990 (N_7990,N_4264,N_5087);
or U7991 (N_7991,N_4818,N_5076);
xor U7992 (N_7992,N_5523,N_5251);
and U7993 (N_7993,N_5909,N_5247);
or U7994 (N_7994,N_4630,N_5093);
nor U7995 (N_7995,N_4356,N_5185);
and U7996 (N_7996,N_4660,N_5400);
nand U7997 (N_7997,N_4556,N_4148);
and U7998 (N_7998,N_4438,N_5876);
nand U7999 (N_7999,N_5514,N_5799);
nand U8000 (N_8000,N_7119,N_7592);
xnor U8001 (N_8001,N_6721,N_7266);
xnor U8002 (N_8002,N_6112,N_6533);
xnor U8003 (N_8003,N_6894,N_7216);
and U8004 (N_8004,N_6620,N_6786);
or U8005 (N_8005,N_7547,N_6541);
and U8006 (N_8006,N_7263,N_6836);
and U8007 (N_8007,N_6065,N_7910);
nor U8008 (N_8008,N_7027,N_7505);
nand U8009 (N_8009,N_6148,N_7156);
xnor U8010 (N_8010,N_6986,N_6519);
and U8011 (N_8011,N_7474,N_7179);
or U8012 (N_8012,N_6653,N_6466);
or U8013 (N_8013,N_7256,N_7258);
nand U8014 (N_8014,N_7674,N_7337);
xnor U8015 (N_8015,N_7432,N_7627);
nor U8016 (N_8016,N_7064,N_6480);
xnor U8017 (N_8017,N_7799,N_6957);
nor U8018 (N_8018,N_7545,N_6874);
nor U8019 (N_8019,N_6759,N_6204);
nor U8020 (N_8020,N_6387,N_7737);
xor U8021 (N_8021,N_6326,N_7588);
and U8022 (N_8022,N_6464,N_7334);
xnor U8023 (N_8023,N_7480,N_6214);
nor U8024 (N_8024,N_6779,N_6009);
and U8025 (N_8025,N_6956,N_6699);
nand U8026 (N_8026,N_6722,N_7819);
and U8027 (N_8027,N_7289,N_7053);
nor U8028 (N_8028,N_7300,N_7276);
or U8029 (N_8029,N_6709,N_6975);
or U8030 (N_8030,N_6943,N_7026);
and U8031 (N_8031,N_6820,N_7690);
and U8032 (N_8032,N_6461,N_6013);
and U8033 (N_8033,N_6069,N_7742);
nor U8034 (N_8034,N_7921,N_7257);
nor U8035 (N_8035,N_6598,N_6673);
nor U8036 (N_8036,N_7233,N_6187);
xnor U8037 (N_8037,N_7596,N_7293);
nand U8038 (N_8038,N_7701,N_6597);
or U8039 (N_8039,N_6645,N_7851);
or U8040 (N_8040,N_6737,N_6573);
and U8041 (N_8041,N_7291,N_7111);
and U8042 (N_8042,N_6727,N_6752);
xnor U8043 (N_8043,N_7907,N_7242);
and U8044 (N_8044,N_6562,N_6024);
or U8045 (N_8045,N_7063,N_7144);
xnor U8046 (N_8046,N_6321,N_7874);
and U8047 (N_8047,N_7767,N_6510);
nor U8048 (N_8048,N_6071,N_7172);
and U8049 (N_8049,N_6932,N_7735);
xor U8050 (N_8050,N_6879,N_6367);
nor U8051 (N_8051,N_7302,N_7724);
nand U8052 (N_8052,N_7857,N_6363);
nor U8053 (N_8053,N_6710,N_6790);
nor U8054 (N_8054,N_6294,N_6390);
and U8055 (N_8055,N_6073,N_7615);
or U8056 (N_8056,N_7294,N_7285);
and U8057 (N_8057,N_7830,N_6170);
nor U8058 (N_8058,N_6217,N_7990);
or U8059 (N_8059,N_6724,N_7653);
nand U8060 (N_8060,N_7782,N_6923);
nand U8061 (N_8061,N_6302,N_6010);
nand U8062 (N_8062,N_7981,N_7239);
xor U8063 (N_8063,N_7850,N_7862);
nor U8064 (N_8064,N_7549,N_6555);
nor U8065 (N_8065,N_7992,N_6140);
or U8066 (N_8066,N_6646,N_7071);
nand U8067 (N_8067,N_6816,N_7790);
or U8068 (N_8068,N_7430,N_7139);
nor U8069 (N_8069,N_6889,N_6843);
and U8070 (N_8070,N_7447,N_6216);
or U8071 (N_8071,N_7221,N_6354);
or U8072 (N_8072,N_6096,N_6058);
or U8073 (N_8073,N_7572,N_6019);
nor U8074 (N_8074,N_7884,N_7475);
or U8075 (N_8075,N_7299,N_7691);
xor U8076 (N_8076,N_7553,N_6772);
and U8077 (N_8077,N_6409,N_6091);
or U8078 (N_8078,N_6236,N_7120);
and U8079 (N_8079,N_7563,N_7567);
nand U8080 (N_8080,N_6094,N_6512);
nand U8081 (N_8081,N_6803,N_6522);
xor U8082 (N_8082,N_6574,N_7684);
nand U8083 (N_8083,N_7133,N_6421);
nor U8084 (N_8084,N_6213,N_7388);
nand U8085 (N_8085,N_6507,N_7312);
xor U8086 (N_8086,N_6600,N_7037);
nor U8087 (N_8087,N_6650,N_7279);
nor U8088 (N_8088,N_6061,N_7951);
or U8089 (N_8089,N_6121,N_6928);
and U8090 (N_8090,N_6591,N_6250);
xnor U8091 (N_8091,N_6442,N_7772);
xnor U8092 (N_8092,N_6278,N_7821);
nand U8093 (N_8093,N_6672,N_7496);
xnor U8094 (N_8094,N_7664,N_7775);
or U8095 (N_8095,N_7915,N_7384);
nand U8096 (N_8096,N_6137,N_7917);
nand U8097 (N_8097,N_6356,N_6883);
and U8098 (N_8098,N_6007,N_6253);
xor U8099 (N_8099,N_6114,N_6521);
nand U8100 (N_8100,N_7832,N_6345);
nand U8101 (N_8101,N_6775,N_6164);
xor U8102 (N_8102,N_7296,N_6540);
or U8103 (N_8103,N_6552,N_7713);
xor U8104 (N_8104,N_7804,N_6229);
and U8105 (N_8105,N_6748,N_7741);
xor U8106 (N_8106,N_6664,N_7333);
nand U8107 (N_8107,N_6324,N_6062);
nor U8108 (N_8108,N_6415,N_6159);
nand U8109 (N_8109,N_6681,N_7278);
nand U8110 (N_8110,N_6038,N_7065);
xor U8111 (N_8111,N_6304,N_7918);
nor U8112 (N_8112,N_7226,N_6477);
or U8113 (N_8113,N_6210,N_6362);
nor U8114 (N_8114,N_7222,N_7478);
or U8115 (N_8115,N_7513,N_6628);
and U8116 (N_8116,N_7632,N_7240);
xnor U8117 (N_8117,N_7671,N_6122);
or U8118 (N_8118,N_6799,N_7409);
nor U8119 (N_8119,N_7277,N_6386);
xor U8120 (N_8120,N_6968,N_6878);
nand U8121 (N_8121,N_7620,N_7765);
nor U8122 (N_8122,N_7326,N_6113);
or U8123 (N_8123,N_6614,N_6997);
or U8124 (N_8124,N_7571,N_7194);
or U8125 (N_8125,N_7131,N_6766);
xor U8126 (N_8126,N_7368,N_7739);
nand U8127 (N_8127,N_6316,N_7815);
xnor U8128 (N_8128,N_6310,N_6087);
xor U8129 (N_8129,N_6086,N_7077);
nor U8130 (N_8130,N_7249,N_6987);
nor U8131 (N_8131,N_7831,N_7055);
nor U8132 (N_8132,N_6385,N_7605);
nand U8133 (N_8133,N_7559,N_6166);
and U8134 (N_8134,N_6098,N_6792);
and U8135 (N_8135,N_6182,N_6670);
nand U8136 (N_8136,N_6129,N_6428);
xnor U8137 (N_8137,N_6378,N_6693);
or U8138 (N_8138,N_7116,N_6740);
and U8139 (N_8139,N_7982,N_6747);
or U8140 (N_8140,N_7953,N_6408);
xor U8141 (N_8141,N_6289,N_6831);
nand U8142 (N_8142,N_6089,N_6534);
nand U8143 (N_8143,N_7604,N_7134);
xor U8144 (N_8144,N_7047,N_6818);
or U8145 (N_8145,N_6863,N_6714);
xnor U8146 (N_8146,N_7526,N_7039);
nor U8147 (N_8147,N_7262,N_6280);
xnor U8148 (N_8148,N_6085,N_7636);
and U8149 (N_8149,N_6821,N_7577);
nand U8150 (N_8150,N_6485,N_7007);
nand U8151 (N_8151,N_7871,N_7978);
or U8152 (N_8152,N_6660,N_6003);
nand U8153 (N_8153,N_6504,N_6845);
and U8154 (N_8154,N_7361,N_7033);
xnor U8155 (N_8155,N_6041,N_6736);
xnor U8156 (N_8156,N_7730,N_7527);
and U8157 (N_8157,N_6801,N_7718);
nor U8158 (N_8158,N_6963,N_6617);
nand U8159 (N_8159,N_7667,N_7562);
nand U8160 (N_8160,N_7543,N_7974);
nor U8161 (N_8161,N_7237,N_7014);
nor U8162 (N_8162,N_7297,N_7695);
nor U8163 (N_8163,N_6804,N_6638);
or U8164 (N_8164,N_6719,N_6373);
nand U8165 (N_8165,N_7341,N_6847);
nand U8166 (N_8166,N_7252,N_6626);
or U8167 (N_8167,N_7646,N_7301);
and U8168 (N_8168,N_6494,N_7976);
nand U8169 (N_8169,N_7098,N_6520);
and U8170 (N_8170,N_7750,N_6870);
and U8171 (N_8171,N_7676,N_7687);
or U8172 (N_8172,N_7281,N_7184);
or U8173 (N_8173,N_7440,N_6749);
nand U8174 (N_8174,N_6579,N_6208);
and U8175 (N_8175,N_6469,N_6509);
and U8176 (N_8176,N_7408,N_7740);
and U8177 (N_8177,N_6109,N_6364);
and U8178 (N_8178,N_6704,N_6479);
nand U8179 (N_8179,N_6959,N_7497);
or U8180 (N_8180,N_7316,N_7158);
xnor U8181 (N_8181,N_7348,N_6970);
xnor U8182 (N_8182,N_7454,N_7437);
or U8183 (N_8183,N_7896,N_6791);
and U8184 (N_8184,N_6965,N_7255);
and U8185 (N_8185,N_6658,N_6769);
xor U8186 (N_8186,N_6679,N_6891);
xor U8187 (N_8187,N_7020,N_6738);
and U8188 (N_8188,N_7486,N_6331);
nor U8189 (N_8189,N_6339,N_7413);
xnor U8190 (N_8190,N_6794,N_6875);
or U8191 (N_8191,N_6106,N_7492);
xor U8192 (N_8192,N_6616,N_7731);
nor U8193 (N_8193,N_7253,N_6904);
nand U8194 (N_8194,N_6536,N_6424);
or U8195 (N_8195,N_6941,N_6695);
nand U8196 (N_8196,N_7135,N_7309);
xnor U8197 (N_8197,N_6404,N_7891);
or U8198 (N_8198,N_7833,N_7234);
and U8199 (N_8199,N_7322,N_6841);
or U8200 (N_8200,N_6989,N_7401);
or U8201 (N_8201,N_6272,N_6773);
and U8202 (N_8202,N_7814,N_6950);
nor U8203 (N_8203,N_6342,N_7160);
nor U8204 (N_8204,N_7888,N_6497);
nand U8205 (N_8205,N_7186,N_6276);
nand U8206 (N_8206,N_7611,N_7254);
nor U8207 (N_8207,N_7762,N_6335);
nor U8208 (N_8208,N_7363,N_6160);
nor U8209 (N_8209,N_6046,N_6806);
or U8210 (N_8210,N_7504,N_6982);
nand U8211 (N_8211,N_6256,N_6438);
and U8212 (N_8212,N_6221,N_7939);
nor U8213 (N_8213,N_7345,N_6005);
and U8214 (N_8214,N_6636,N_7783);
or U8215 (N_8215,N_6822,N_7425);
or U8216 (N_8216,N_6960,N_7268);
nand U8217 (N_8217,N_7335,N_6074);
xnor U8218 (N_8218,N_7968,N_6212);
xor U8219 (N_8219,N_7867,N_6683);
nand U8220 (N_8220,N_7847,N_7107);
xnor U8221 (N_8221,N_6267,N_6102);
nor U8222 (N_8222,N_7964,N_6254);
or U8223 (N_8223,N_7493,N_6535);
or U8224 (N_8224,N_6030,N_7054);
nor U8225 (N_8225,N_7954,N_6998);
nand U8226 (N_8226,N_6687,N_6674);
and U8227 (N_8227,N_6243,N_7359);
xor U8228 (N_8228,N_7072,N_6531);
xor U8229 (N_8229,N_6633,N_6036);
or U8230 (N_8230,N_6143,N_6783);
xnor U8231 (N_8231,N_6976,N_6282);
xnor U8232 (N_8232,N_6690,N_7641);
and U8233 (N_8233,N_6774,N_7423);
and U8234 (N_8234,N_7928,N_7069);
or U8235 (N_8235,N_7558,N_7381);
xnor U8236 (N_8236,N_6039,N_6973);
and U8237 (N_8237,N_6835,N_6516);
nand U8238 (N_8238,N_7882,N_7744);
or U8239 (N_8239,N_7931,N_6527);
nor U8240 (N_8240,N_7150,N_7868);
nor U8241 (N_8241,N_6120,N_7379);
or U8242 (N_8242,N_6517,N_6014);
or U8243 (N_8243,N_7115,N_6225);
or U8244 (N_8244,N_7930,N_6530);
or U8245 (N_8245,N_7052,N_6201);
and U8246 (N_8246,N_6788,N_7051);
and U8247 (N_8247,N_7102,N_7913);
or U8248 (N_8248,N_7777,N_7248);
nor U8249 (N_8249,N_6340,N_7709);
and U8250 (N_8250,N_6903,N_6427);
xor U8251 (N_8251,N_7898,N_7550);
nand U8252 (N_8252,N_6206,N_6172);
nand U8253 (N_8253,N_6183,N_7365);
xor U8254 (N_8254,N_6978,N_6162);
nand U8255 (N_8255,N_7328,N_6716);
xor U8256 (N_8256,N_7999,N_7199);
xnor U8257 (N_8257,N_6457,N_7344);
nand U8258 (N_8258,N_7477,N_6796);
nand U8259 (N_8259,N_6352,N_6819);
xnor U8260 (N_8260,N_7755,N_7729);
xnor U8261 (N_8261,N_6966,N_6499);
or U8262 (N_8262,N_7843,N_7142);
nand U8263 (N_8263,N_7987,N_7897);
nor U8264 (N_8264,N_6899,N_7370);
nand U8265 (N_8265,N_7151,N_6228);
nor U8266 (N_8266,N_7532,N_7637);
nand U8267 (N_8267,N_6478,N_6238);
and U8268 (N_8268,N_6505,N_7779);
nand U8269 (N_8269,N_7374,N_7812);
or U8270 (N_8270,N_7873,N_7795);
nand U8271 (N_8271,N_6262,N_6511);
xor U8272 (N_8272,N_6103,N_7323);
or U8273 (N_8273,N_7452,N_7540);
and U8274 (N_8274,N_6190,N_6887);
and U8275 (N_8275,N_6888,N_6919);
xor U8276 (N_8276,N_6460,N_6248);
nor U8277 (N_8277,N_7267,N_7236);
nor U8278 (N_8278,N_6800,N_6470);
or U8279 (N_8279,N_6615,N_7668);
nor U8280 (N_8280,N_7419,N_6564);
nor U8281 (N_8281,N_7171,N_7786);
xnor U8282 (N_8282,N_7863,N_7619);
nor U8283 (N_8283,N_6667,N_7778);
nor U8284 (N_8284,N_7209,N_7560);
nor U8285 (N_8285,N_6920,N_6380);
nor U8286 (N_8286,N_7925,N_6045);
and U8287 (N_8287,N_7745,N_6732);
nand U8288 (N_8288,N_7187,N_6741);
nand U8289 (N_8289,N_7317,N_7659);
or U8290 (N_8290,N_6589,N_6153);
xor U8291 (N_8291,N_6059,N_6951);
or U8292 (N_8292,N_6846,N_7938);
nand U8293 (N_8293,N_7483,N_7084);
or U8294 (N_8294,N_7869,N_6168);
or U8295 (N_8295,N_6524,N_6654);
xnor U8296 (N_8296,N_7114,N_7177);
nor U8297 (N_8297,N_6083,N_7679);
xnor U8298 (N_8298,N_7717,N_6451);
nor U8299 (N_8299,N_6441,N_6034);
and U8300 (N_8300,N_7660,N_7518);
nand U8301 (N_8301,N_6866,N_6247);
nand U8302 (N_8302,N_6056,N_7399);
and U8303 (N_8303,N_6506,N_7723);
nor U8304 (N_8304,N_7298,N_7510);
xor U8305 (N_8305,N_7716,N_7751);
nor U8306 (N_8306,N_6157,N_6076);
xor U8307 (N_8307,N_6163,N_7612);
or U8308 (N_8308,N_6420,N_7600);
or U8309 (N_8309,N_7929,N_6082);
nor U8310 (N_8310,N_6500,N_6662);
nand U8311 (N_8311,N_6015,N_6360);
nor U8312 (N_8312,N_6131,N_6832);
and U8313 (N_8313,N_7826,N_6611);
and U8314 (N_8314,N_7811,N_6604);
and U8315 (N_8315,N_7446,N_6697);
nor U8316 (N_8316,N_6227,N_6255);
nand U8317 (N_8317,N_6343,N_6379);
or U8318 (N_8318,N_6659,N_6447);
nand U8319 (N_8319,N_7960,N_7075);
or U8320 (N_8320,N_6576,N_7651);
xnor U8321 (N_8321,N_6651,N_6720);
and U8322 (N_8322,N_7643,N_6991);
xnor U8323 (N_8323,N_7083,N_6105);
or U8324 (N_8324,N_7235,N_7470);
or U8325 (N_8325,N_6433,N_7173);
nor U8326 (N_8326,N_7318,N_7774);
nand U8327 (N_8327,N_6055,N_6876);
xor U8328 (N_8328,N_6329,N_6900);
xor U8329 (N_8329,N_7011,N_6572);
or U8330 (N_8330,N_7642,N_6554);
or U8331 (N_8331,N_7906,N_6145);
and U8332 (N_8332,N_6458,N_7193);
xor U8333 (N_8333,N_6934,N_7472);
and U8334 (N_8334,N_6666,N_6043);
xnor U8335 (N_8335,N_6307,N_6117);
or U8336 (N_8336,N_6242,N_7336);
and U8337 (N_8337,N_7692,N_6301);
nand U8338 (N_8338,N_7168,N_7457);
or U8339 (N_8339,N_6205,N_7564);
xor U8340 (N_8340,N_7698,N_7424);
nand U8341 (N_8341,N_7061,N_6188);
and U8342 (N_8342,N_7155,N_7165);
nand U8343 (N_8343,N_6268,N_6209);
and U8344 (N_8344,N_6361,N_6634);
xor U8345 (N_8345,N_6156,N_6292);
or U8346 (N_8346,N_6703,N_6798);
and U8347 (N_8347,N_6669,N_7580);
or U8348 (N_8348,N_6068,N_7308);
xor U8349 (N_8349,N_7245,N_6141);
xor U8350 (N_8350,N_7124,N_7319);
nor U8351 (N_8351,N_7962,N_6501);
or U8352 (N_8352,N_7770,N_7176);
nor U8353 (N_8353,N_6244,N_7259);
xnor U8354 (N_8354,N_7228,N_7128);
xnor U8355 (N_8355,N_7736,N_6186);
or U8356 (N_8356,N_6211,N_7759);
and U8357 (N_8357,N_7449,N_6635);
and U8358 (N_8358,N_6912,N_6948);
nor U8359 (N_8359,N_7190,N_6868);
and U8360 (N_8360,N_6592,N_7840);
nor U8361 (N_8361,N_6486,N_6807);
nand U8362 (N_8362,N_6852,N_7028);
and U8363 (N_8363,N_7509,N_6627);
or U8364 (N_8364,N_7196,N_7043);
and U8365 (N_8365,N_7488,N_6622);
nand U8366 (N_8366,N_6528,N_6334);
and U8367 (N_8367,N_6685,N_7796);
or U8368 (N_8368,N_7614,N_7104);
xnor U8369 (N_8369,N_7665,N_7994);
nand U8370 (N_8370,N_6861,N_6290);
nor U8371 (N_8371,N_6696,N_6853);
nand U8372 (N_8372,N_7748,N_6151);
nand U8373 (N_8373,N_7973,N_7244);
and U8374 (N_8374,N_6601,N_7773);
and U8375 (N_8375,N_7024,N_7110);
nor U8376 (N_8376,N_7310,N_6608);
nor U8377 (N_8377,N_6291,N_6218);
and U8378 (N_8378,N_6179,N_7066);
nand U8379 (N_8379,N_7824,N_7481);
and U8380 (N_8380,N_6771,N_7108);
nand U8381 (N_8381,N_7441,N_6134);
nor U8382 (N_8382,N_7342,N_6181);
or U8383 (N_8383,N_7204,N_6896);
or U8384 (N_8384,N_7945,N_7476);
or U8385 (N_8385,N_6715,N_7264);
xnor U8386 (N_8386,N_7284,N_6728);
nand U8387 (N_8387,N_7434,N_6758);
nor U8388 (N_8388,N_6610,N_6926);
and U8389 (N_8389,N_6127,N_7975);
or U8390 (N_8390,N_7520,N_7576);
and U8391 (N_8391,N_6877,N_6124);
or U8392 (N_8392,N_6901,N_7188);
and U8393 (N_8393,N_7315,N_7680);
or U8394 (N_8394,N_6805,N_7455);
or U8395 (N_8395,N_6178,N_7087);
nor U8396 (N_8396,N_6906,N_7644);
and U8397 (N_8397,N_6964,N_7860);
nor U8398 (N_8398,N_6219,N_6746);
or U8399 (N_8399,N_7426,N_7835);
and U8400 (N_8400,N_7113,N_7827);
and U8401 (N_8401,N_7369,N_6049);
nor U8402 (N_8402,N_6882,N_6547);
and U8403 (N_8403,N_6436,N_6862);
nand U8404 (N_8404,N_7595,N_6128);
or U8405 (N_8405,N_7586,N_6471);
xnor U8406 (N_8406,N_7211,N_7057);
nor U8407 (N_8407,N_6979,N_7273);
and U8408 (N_8408,N_6871,N_6080);
or U8409 (N_8409,N_6180,N_7088);
or U8410 (N_8410,N_6169,N_6284);
xor U8411 (N_8411,N_7937,N_7602);
nand U8412 (N_8412,N_6817,N_7501);
nor U8413 (N_8413,N_6177,N_6135);
or U8414 (N_8414,N_7170,N_6851);
or U8415 (N_8415,N_6051,N_7531);
and U8416 (N_8416,N_6780,N_6189);
nor U8417 (N_8417,N_7996,N_6375);
nand U8418 (N_8418,N_6556,N_6526);
or U8419 (N_8419,N_6915,N_7629);
nor U8420 (N_8420,N_7569,N_6174);
nand U8421 (N_8421,N_7593,N_7608);
nor U8422 (N_8422,N_7045,N_7371);
xor U8423 (N_8423,N_7582,N_7375);
or U8424 (N_8424,N_7948,N_6435);
or U8425 (N_8425,N_6338,N_6084);
nand U8426 (N_8426,N_6833,N_7247);
nand U8427 (N_8427,N_6663,N_7157);
nand U8428 (N_8428,N_7422,N_7788);
and U8429 (N_8429,N_7373,N_6226);
xor U8430 (N_8430,N_6252,N_7224);
and U8431 (N_8431,N_6930,N_6040);
nand U8432 (N_8432,N_6612,N_7645);
nand U8433 (N_8433,N_6365,N_7597);
and U8434 (N_8434,N_6668,N_7140);
nand U8435 (N_8435,N_7838,N_7215);
nor U8436 (N_8436,N_7557,N_6023);
nand U8437 (N_8437,N_6462,N_7947);
nand U8438 (N_8438,N_7949,N_7647);
and U8439 (N_8439,N_6585,N_6347);
or U8440 (N_8440,N_6406,N_7428);
and U8441 (N_8441,N_6762,N_7243);
nor U8442 (N_8442,N_6575,N_6398);
xor U8443 (N_8443,N_6389,N_7924);
or U8444 (N_8444,N_7521,N_7306);
and U8445 (N_8445,N_7901,N_7433);
xor U8446 (N_8446,N_7585,N_6999);
and U8447 (N_8447,N_7519,N_7095);
nand U8448 (N_8448,N_7019,N_7436);
or U8449 (N_8449,N_7227,N_7936);
nor U8450 (N_8450,N_6656,N_6197);
or U8451 (N_8451,N_6465,N_7205);
and U8452 (N_8452,N_6273,N_6220);
nand U8453 (N_8453,N_7881,N_6152);
and U8454 (N_8454,N_6088,N_6767);
nand U8455 (N_8455,N_7386,N_7538);
nor U8456 (N_8456,N_7448,N_6760);
xor U8457 (N_8457,N_6570,N_7502);
and U8458 (N_8458,N_6557,N_6643);
and U8459 (N_8459,N_6823,N_7908);
xor U8460 (N_8460,N_6070,N_6605);
xor U8461 (N_8461,N_7984,N_7411);
and U8462 (N_8462,N_6311,N_7080);
or U8463 (N_8463,N_6132,N_6974);
nand U8464 (N_8464,N_7303,N_7806);
or U8465 (N_8465,N_6810,N_6498);
or U8466 (N_8466,N_6980,N_7435);
nor U8467 (N_8467,N_6949,N_7272);
nor U8468 (N_8468,N_7438,N_7805);
or U8469 (N_8469,N_6450,N_7185);
xnor U8470 (N_8470,N_7031,N_6239);
nor U8471 (N_8471,N_6448,N_6850);
or U8472 (N_8472,N_6495,N_7621);
and U8473 (N_8473,N_6582,N_7892);
nor U8474 (N_8474,N_7442,N_6586);
nor U8475 (N_8475,N_7813,N_7633);
nor U8476 (N_8476,N_7378,N_7453);
xor U8477 (N_8477,N_7630,N_7919);
xnor U8478 (N_8478,N_7872,N_6463);
nor U8479 (N_8479,N_7121,N_6092);
nor U8480 (N_8480,N_7997,N_6453);
xor U8481 (N_8481,N_6518,N_6558);
nand U8482 (N_8482,N_6158,N_6677);
nand U8483 (N_8483,N_7606,N_7752);
nand U8484 (N_8484,N_7710,N_7885);
xor U8485 (N_8485,N_6537,N_6118);
or U8486 (N_8486,N_7040,N_6684);
xnor U8487 (N_8487,N_7030,N_7327);
or U8488 (N_8488,N_6355,N_7785);
nand U8489 (N_8489,N_7986,N_7985);
nand U8490 (N_8490,N_7420,N_7587);
or U8491 (N_8491,N_6285,N_7566);
and U8492 (N_8492,N_7094,N_6348);
or U8493 (N_8493,N_6892,N_6496);
nor U8494 (N_8494,N_6545,N_6940);
nand U8495 (N_8495,N_7246,N_6542);
nor U8496 (N_8496,N_6712,N_7856);
nand U8497 (N_8497,N_6288,N_7141);
nand U8498 (N_8498,N_7610,N_7803);
or U8499 (N_8499,N_6490,N_6726);
nor U8500 (N_8500,N_6327,N_7229);
or U8501 (N_8501,N_7079,N_7666);
and U8502 (N_8502,N_6825,N_7387);
nor U8503 (N_8503,N_7561,N_7360);
and U8504 (N_8504,N_6430,N_7678);
or U8505 (N_8505,N_6493,N_6349);
and U8506 (N_8506,N_6731,N_7238);
nor U8507 (N_8507,N_7093,N_7212);
xor U8508 (N_8508,N_7340,N_6815);
nor U8509 (N_8509,N_7015,N_6370);
nor U8510 (N_8510,N_7200,N_7952);
nand U8511 (N_8511,N_7893,N_6245);
and U8512 (N_8512,N_6655,N_6006);
nor U8513 (N_8513,N_7078,N_6060);
nand U8514 (N_8514,N_6649,N_7681);
nand U8515 (N_8515,N_7980,N_7714);
xor U8516 (N_8516,N_6565,N_6864);
or U8517 (N_8517,N_6057,N_7904);
xor U8518 (N_8518,N_6613,N_7397);
nor U8519 (N_8519,N_6184,N_7848);
and U8520 (N_8520,N_7902,N_6175);
nand U8521 (N_8521,N_6011,N_7738);
xnor U8522 (N_8522,N_6962,N_7353);
xor U8523 (N_8523,N_6346,N_6539);
or U8524 (N_8524,N_7594,N_7351);
nor U8525 (N_8525,N_7797,N_7313);
nand U8526 (N_8526,N_6251,N_7943);
xor U8527 (N_8527,N_6199,N_7161);
or U8528 (N_8528,N_6277,N_7844);
or U8529 (N_8529,N_7617,N_7966);
and U8530 (N_8530,N_6571,N_6914);
xor U8531 (N_8531,N_7265,N_7495);
and U8532 (N_8532,N_7946,N_6032);
or U8533 (N_8533,N_7705,N_7164);
xnor U8534 (N_8534,N_6761,N_6328);
xor U8535 (N_8535,N_7972,N_7802);
xor U8536 (N_8536,N_6437,N_6624);
xnor U8537 (N_8537,N_7903,N_7129);
xor U8538 (N_8538,N_7590,N_6795);
nor U8539 (N_8539,N_7458,N_7622);
and U8540 (N_8540,N_7682,N_7760);
nand U8541 (N_8541,N_7537,N_6640);
nand U8542 (N_8542,N_6482,N_7696);
or U8543 (N_8543,N_7147,N_7749);
and U8544 (N_8544,N_6739,N_6925);
and U8545 (N_8545,N_7321,N_7971);
or U8546 (N_8546,N_6203,N_7747);
and U8547 (N_8547,N_7781,N_6647);
or U8548 (N_8548,N_6755,N_6858);
and U8549 (N_8549,N_7096,N_6675);
xnor U8550 (N_8550,N_7183,N_6033);
xor U8551 (N_8551,N_6336,N_7914);
xnor U8552 (N_8552,N_6322,N_7439);
and U8553 (N_8553,N_7117,N_7603);
or U8554 (N_8554,N_6566,N_6793);
nor U8555 (N_8555,N_7089,N_6723);
xor U8556 (N_8556,N_7726,N_7524);
nand U8557 (N_8557,N_6785,N_7876);
and U8558 (N_8558,N_6192,N_6394);
nor U8559 (N_8559,N_6742,N_6027);
and U8560 (N_8560,N_7837,N_6350);
nand U8561 (N_8561,N_6492,N_7877);
nor U8562 (N_8562,N_7712,N_6265);
nor U8563 (N_8563,N_6827,N_7648);
nand U8564 (N_8564,N_7287,N_6167);
or U8565 (N_8565,N_6577,N_6366);
and U8566 (N_8566,N_7103,N_7013);
or U8567 (N_8567,N_7589,N_6413);
nand U8568 (N_8568,N_7574,N_6995);
xnor U8569 (N_8569,N_7656,N_7555);
nand U8570 (N_8570,N_6898,N_7100);
xor U8571 (N_8571,N_7638,N_6020);
and U8572 (N_8572,N_7022,N_6559);
nand U8573 (N_8573,N_7029,N_7685);
and U8574 (N_8574,N_7325,N_6993);
nor U8575 (N_8575,N_6440,N_7444);
and U8576 (N_8576,N_6602,N_7776);
nand U8577 (N_8577,N_6484,N_6459);
nor U8578 (N_8578,N_7372,N_7208);
and U8579 (N_8579,N_6581,N_7652);
xnor U8580 (N_8580,N_7626,N_6468);
and U8581 (N_8581,N_7499,N_7197);
or U8582 (N_8582,N_6977,N_7230);
nand U8583 (N_8583,N_6176,N_6909);
or U8584 (N_8584,N_6308,N_6235);
and U8585 (N_8585,N_6917,N_6411);
or U8586 (N_8586,N_6309,N_6905);
or U8587 (N_8587,N_7828,N_7035);
nand U8588 (N_8588,N_7127,N_6115);
nor U8589 (N_8589,N_6711,N_7346);
nor U8590 (N_8590,N_7009,N_7533);
and U8591 (N_8591,N_6671,N_6947);
or U8592 (N_8592,N_7416,N_6475);
or U8593 (N_8593,N_7377,N_7355);
nor U8594 (N_8594,N_7733,N_7182);
or U8595 (N_8595,N_7471,N_7658);
and U8596 (N_8596,N_7757,N_6258);
nand U8597 (N_8597,N_7699,N_7989);
nand U8598 (N_8598,N_7864,N_6754);
xor U8599 (N_8599,N_6018,N_7922);
and U8600 (N_8600,N_6745,N_6708);
or U8601 (N_8601,N_6026,N_7214);
and U8602 (N_8602,N_7280,N_7283);
and U8603 (N_8603,N_6954,N_6416);
and U8604 (N_8604,N_7097,N_7271);
nor U8605 (N_8605,N_6502,N_6777);
and U8606 (N_8606,N_7583,N_6047);
nand U8607 (N_8607,N_6474,N_7106);
nand U8608 (N_8608,N_7356,N_7305);
or U8609 (N_8609,N_7941,N_7132);
nand U8610 (N_8610,N_6553,N_6231);
nand U8611 (N_8611,N_6418,N_6865);
nor U8612 (N_8612,N_7191,N_7203);
and U8613 (N_8613,N_6452,N_7787);
and U8614 (N_8614,N_7957,N_6397);
nand U8615 (N_8615,N_6908,N_6686);
or U8616 (N_8616,N_7702,N_6808);
nor U8617 (N_8617,N_6717,N_6637);
and U8618 (N_8618,N_6130,N_7414);
or U8619 (N_8619,N_6630,N_7081);
nand U8620 (N_8620,N_6374,N_7818);
and U8621 (N_8621,N_7807,N_6372);
nor U8622 (N_8622,N_6593,N_6263);
nor U8623 (N_8623,N_7711,N_6606);
nor U8624 (N_8624,N_7112,N_7822);
and U8625 (N_8625,N_7390,N_7181);
nand U8626 (N_8626,N_7940,N_7578);
xor U8627 (N_8627,N_6300,N_6369);
xor U8628 (N_8628,N_7508,N_7418);
nor U8629 (N_8629,N_7466,N_6902);
nor U8630 (N_8630,N_6002,N_7661);
nand U8631 (N_8631,N_6224,N_6546);
nor U8632 (N_8632,N_6139,N_7955);
nor U8633 (N_8633,N_7820,N_7693);
xnor U8634 (N_8634,N_6313,N_6296);
nand U8635 (N_8635,N_7662,N_6916);
and U8636 (N_8636,N_6391,N_6395);
nand U8637 (N_8637,N_6149,N_7138);
and U8638 (N_8638,N_6042,N_6481);
nand U8639 (N_8639,N_7146,N_7484);
or U8640 (N_8640,N_6569,N_6107);
nand U8641 (N_8641,N_7573,N_7849);
and U8642 (N_8642,N_6955,N_7366);
xor U8643 (N_8643,N_7825,N_7099);
nand U8644 (N_8644,N_7883,N_6483);
nor U8645 (N_8645,N_7082,N_6691);
nor U8646 (N_8646,N_7395,N_6330);
nand U8647 (N_8647,N_7003,N_6171);
nand U8648 (N_8648,N_6101,N_7808);
nand U8649 (N_8649,N_7076,N_6337);
and U8650 (N_8650,N_7991,N_6138);
and U8651 (N_8651,N_6532,N_6682);
or U8652 (N_8652,N_6580,N_6890);
and U8653 (N_8653,N_6994,N_7655);
nand U8654 (N_8654,N_6426,N_6417);
and U8655 (N_8655,N_6078,N_7367);
and U8656 (N_8656,N_7500,N_7528);
nand U8657 (N_8657,N_7012,N_6560);
nor U8658 (N_8658,N_7101,N_6401);
nor U8659 (N_8659,N_7514,N_6588);
nand U8660 (N_8660,N_7330,N_7609);
nor U8661 (N_8661,N_7581,N_6665);
xor U8662 (N_8662,N_6232,N_7565);
xor U8663 (N_8663,N_7923,N_7932);
nor U8664 (N_8664,N_6445,N_6393);
and U8665 (N_8665,N_7570,N_7899);
and U8666 (N_8666,N_6824,N_7137);
and U8667 (N_8667,N_6368,N_7122);
nor U8668 (N_8668,N_7362,N_6578);
nor U8669 (N_8669,N_6623,N_6990);
and U8670 (N_8670,N_6233,N_6155);
nand U8671 (N_8671,N_6895,N_7311);
or U8672 (N_8672,N_7412,N_7634);
or U8673 (N_8673,N_6194,N_6097);
nor U8674 (N_8674,N_7926,N_6881);
or U8675 (N_8675,N_6809,N_7331);
nor U8676 (N_8676,N_6467,N_7163);
or U8677 (N_8677,N_6312,N_7169);
and U8678 (N_8678,N_6142,N_7201);
nand U8679 (N_8679,N_7546,N_6029);
or U8680 (N_8680,N_6472,N_6066);
and U8681 (N_8681,N_7464,N_7631);
nor U8682 (N_8682,N_6414,N_7886);
xor U8683 (N_8683,N_7261,N_6111);
or U8684 (N_8684,N_6599,N_7324);
and U8685 (N_8685,N_6028,N_7092);
xnor U8686 (N_8686,N_7041,N_7220);
nor U8687 (N_8687,N_7544,N_7623);
nand U8688 (N_8688,N_7556,N_6644);
xnor U8689 (N_8689,N_6885,N_7548);
and U8690 (N_8690,N_6680,N_7942);
xor U8691 (N_8691,N_7450,N_6104);
nand U8692 (N_8692,N_7153,N_7858);
or U8693 (N_8693,N_6849,N_6688);
and U8694 (N_8694,N_7618,N_7639);
and U8695 (N_8695,N_7148,N_7697);
and U8696 (N_8696,N_6319,N_7460);
or U8697 (N_8697,N_6434,N_7451);
nand U8698 (N_8698,N_6207,N_7469);
and U8699 (N_8699,N_6778,N_7584);
xor U8700 (N_8700,N_7601,N_6607);
and U8701 (N_8701,N_7771,N_7516);
or U8702 (N_8702,N_6333,N_6828);
xor U8703 (N_8703,N_7491,N_7649);
xnor U8704 (N_8704,N_7743,N_6757);
xnor U8705 (N_8705,N_7398,N_6587);
and U8706 (N_8706,N_7912,N_7789);
xor U8707 (N_8707,N_6269,N_6857);
or U8708 (N_8708,N_6392,N_7406);
nor U8709 (N_8709,N_6842,N_7541);
and U8710 (N_8710,N_6971,N_6544);
nand U8711 (N_8711,N_6402,N_7959);
and U8712 (N_8712,N_7178,N_7956);
xnor U8713 (N_8713,N_7988,N_6025);
and U8714 (N_8714,N_7854,N_7599);
xnor U8715 (N_8715,N_7794,N_7274);
nand U8716 (N_8716,N_7720,N_7894);
xor U8717 (N_8717,N_7784,N_7607);
nand U8718 (N_8718,N_6240,N_6297);
nand U8719 (N_8719,N_7686,N_7551);
and U8720 (N_8720,N_6054,N_6455);
nand U8721 (N_8721,N_7405,N_7152);
or U8722 (N_8722,N_7706,N_6834);
or U8723 (N_8723,N_6859,N_7657);
and U8724 (N_8724,N_6924,N_7338);
or U8725 (N_8725,N_6515,N_7909);
or U8726 (N_8726,N_7675,N_6893);
nor U8727 (N_8727,N_6230,N_6323);
nor U8728 (N_8728,N_6306,N_6811);
nand U8729 (N_8729,N_7189,N_7517);
nand U8730 (N_8730,N_6927,N_7482);
or U8731 (N_8731,N_7880,N_6765);
or U8732 (N_8732,N_7260,N_6867);
xor U8733 (N_8733,N_7479,N_6734);
and U8734 (N_8734,N_7431,N_6261);
nor U8735 (N_8735,N_7207,N_6992);
nor U8736 (N_8736,N_7768,N_6946);
xnor U8737 (N_8737,N_6733,N_6972);
and U8738 (N_8738,N_6753,N_7391);
and U8739 (N_8739,N_6812,N_6953);
nand U8740 (N_8740,N_6529,N_7703);
and U8741 (N_8741,N_7766,N_6750);
or U8742 (N_8742,N_7126,N_6844);
xnor U8743 (N_8743,N_7722,N_6405);
or U8744 (N_8744,N_6826,N_6202);
nor U8745 (N_8745,N_7044,N_7801);
and U8746 (N_8746,N_7754,N_6359);
nand U8747 (N_8747,N_7732,N_6099);
xnor U8748 (N_8748,N_7654,N_6781);
and U8749 (N_8749,N_6707,N_6423);
xor U8750 (N_8750,N_6657,N_6584);
or U8751 (N_8751,N_6594,N_7143);
nor U8752 (N_8752,N_7979,N_7983);
or U8753 (N_8753,N_7753,N_7523);
and U8754 (N_8754,N_6488,N_6425);
and U8755 (N_8755,N_7878,N_6136);
and U8756 (N_8756,N_7792,N_6266);
nand U8757 (N_8757,N_6713,N_7049);
nor U8758 (N_8758,N_7445,N_7250);
and U8759 (N_8759,N_7352,N_7769);
nor U8760 (N_8760,N_7963,N_7403);
and U8761 (N_8761,N_7700,N_6035);
xor U8762 (N_8762,N_7853,N_7023);
nand U8763 (N_8763,N_7046,N_7154);
and U8764 (N_8764,N_7525,N_6476);
xor U8765 (N_8765,N_7993,N_6004);
nor U8766 (N_8766,N_6377,N_6249);
and U8767 (N_8767,N_6281,N_7383);
nor U8768 (N_8768,N_7846,N_7536);
nor U8769 (N_8769,N_6000,N_6921);
nand U8770 (N_8770,N_7694,N_6705);
nor U8771 (N_8771,N_6314,N_7034);
nand U8772 (N_8772,N_7887,N_7123);
or U8773 (N_8773,N_6489,N_6325);
and U8774 (N_8774,N_6017,N_7715);
xnor U8775 (N_8775,N_6195,N_6320);
and U8776 (N_8776,N_7487,N_6787);
xnor U8777 (N_8777,N_7042,N_7382);
xnor U8778 (N_8778,N_6133,N_6403);
xor U8779 (N_8779,N_7392,N_6855);
and U8780 (N_8780,N_6837,N_6603);
and U8781 (N_8781,N_6351,N_6317);
or U8782 (N_8782,N_7307,N_6439);
or U8783 (N_8783,N_6913,N_7074);
and U8784 (N_8784,N_7231,N_6075);
or U8785 (N_8785,N_6274,N_7018);
or U8786 (N_8786,N_7364,N_6886);
nor U8787 (N_8787,N_6422,N_6944);
xnor U8788 (N_8788,N_7206,N_6275);
xor U8789 (N_8789,N_7320,N_7977);
nor U8790 (N_8790,N_6725,N_7167);
nor U8791 (N_8791,N_7817,N_7210);
and U8792 (N_8792,N_6095,N_6631);
xor U8793 (N_8793,N_7162,N_7764);
and U8794 (N_8794,N_6371,N_7354);
nand U8795 (N_8795,N_6632,N_7396);
nand U8796 (N_8796,N_6967,N_6031);
nand U8797 (N_8797,N_6072,N_6341);
and U8798 (N_8798,N_7628,N_6456);
and U8799 (N_8799,N_7270,N_7761);
nand U8800 (N_8800,N_6193,N_7728);
nor U8801 (N_8801,N_6446,N_7841);
and U8802 (N_8802,N_6315,N_7879);
nor U8803 (N_8803,N_6081,N_6568);
and U8804 (N_8804,N_7008,N_7032);
and U8805 (N_8805,N_6550,N_6618);
or U8806 (N_8806,N_7515,N_6126);
nor U8807 (N_8807,N_7829,N_7816);
xor U8808 (N_8808,N_6751,N_6173);
xnor U8809 (N_8809,N_6399,N_6768);
or U8810 (N_8810,N_7062,N_6625);
xnor U8811 (N_8811,N_6939,N_7295);
nand U8812 (N_8812,N_7145,N_7404);
nor U8813 (N_8813,N_7852,N_6508);
xor U8814 (N_8814,N_6797,N_7934);
nor U8815 (N_8815,N_6802,N_6410);
and U8816 (N_8816,N_7670,N_7663);
and U8817 (N_8817,N_7021,N_6743);
and U8818 (N_8818,N_6305,N_7579);
or U8819 (N_8819,N_7719,N_7068);
or U8820 (N_8820,N_7625,N_6763);
and U8821 (N_8821,N_6384,N_7889);
nor U8822 (N_8822,N_7005,N_6264);
nor U8823 (N_8823,N_7180,N_7995);
and U8824 (N_8824,N_7218,N_6595);
nand U8825 (N_8825,N_6161,N_7050);
nor U8826 (N_8826,N_6165,N_6619);
nor U8827 (N_8827,N_6983,N_6567);
nand U8828 (N_8828,N_7329,N_6702);
nand U8829 (N_8829,N_6952,N_6454);
nand U8830 (N_8830,N_7010,N_6770);
xor U8831 (N_8831,N_6147,N_7689);
xnor U8832 (N_8832,N_7861,N_6191);
nor U8833 (N_8833,N_6357,N_6388);
nand U8834 (N_8834,N_7554,N_7870);
xor U8835 (N_8835,N_7056,N_7223);
and U8836 (N_8836,N_6150,N_6048);
nand U8837 (N_8837,N_7085,N_6872);
or U8838 (N_8838,N_7534,N_7834);
nand U8839 (N_8839,N_6590,N_6933);
xnor U8840 (N_8840,N_6583,N_7933);
xor U8841 (N_8841,N_6814,N_6503);
nor U8842 (N_8842,N_6694,N_7410);
or U8843 (N_8843,N_7006,N_6279);
or U8844 (N_8844,N_7017,N_7927);
or U8845 (N_8845,N_6922,N_7810);
nor U8846 (N_8846,N_7159,N_7839);
nand U8847 (N_8847,N_6856,N_7842);
nand U8848 (N_8848,N_7568,N_6829);
and U8849 (N_8849,N_6116,N_6839);
or U8850 (N_8850,N_6223,N_7195);
nand U8851 (N_8851,N_6196,N_7463);
or U8852 (N_8852,N_7911,N_7269);
nor U8853 (N_8853,N_7086,N_7961);
xnor U8854 (N_8854,N_6303,N_7746);
and U8855 (N_8855,N_7688,N_7467);
and U8856 (N_8856,N_7542,N_7462);
xnor U8857 (N_8857,N_6108,N_7241);
nor U8858 (N_8858,N_7865,N_6596);
or U8859 (N_8859,N_6958,N_6257);
or U8860 (N_8860,N_6563,N_7485);
and U8861 (N_8861,N_7530,N_6260);
nand U8862 (N_8862,N_7225,N_6396);
nand U8863 (N_8863,N_7512,N_6287);
or U8864 (N_8864,N_7202,N_7905);
nand U8865 (N_8865,N_6756,N_6077);
nor U8866 (N_8866,N_6044,N_7791);
and U8867 (N_8867,N_6419,N_7415);
and U8868 (N_8868,N_6945,N_6938);
nand U8869 (N_8869,N_6840,N_7036);
and U8870 (N_8870,N_7343,N_6241);
nor U8871 (N_8871,N_7166,N_6052);
nor U8872 (N_8872,N_7780,N_7136);
nand U8873 (N_8873,N_6286,N_6525);
or U8874 (N_8874,N_6910,N_7038);
nand U8875 (N_8875,N_7358,N_7393);
nand U8876 (N_8876,N_7800,N_7060);
xor U8877 (N_8877,N_7809,N_7456);
and U8878 (N_8878,N_6735,N_7616);
nor U8879 (N_8879,N_6090,N_6332);
nand U8880 (N_8880,N_6869,N_6609);
nor U8881 (N_8881,N_7461,N_7130);
or U8882 (N_8882,N_6293,N_7339);
or U8883 (N_8883,N_6271,N_6549);
and U8884 (N_8884,N_7473,N_6237);
and U8885 (N_8885,N_6784,N_6848);
and U8886 (N_8886,N_6432,N_7443);
xnor U8887 (N_8887,N_6146,N_6678);
nor U8888 (N_8888,N_7672,N_7059);
nand U8889 (N_8889,N_6523,N_6123);
xnor U8890 (N_8890,N_7635,N_6298);
nor U8891 (N_8891,N_6931,N_7763);
xnor U8892 (N_8892,N_7067,N_7823);
or U8893 (N_8893,N_7494,N_6730);
and U8894 (N_8894,N_6001,N_7349);
xnor U8895 (N_8895,N_6860,N_7669);
or U8896 (N_8896,N_7350,N_6144);
nor U8897 (N_8897,N_7468,N_7859);
xnor U8898 (N_8898,N_7969,N_7895);
xnor U8899 (N_8899,N_6429,N_7091);
nand U8900 (N_8900,N_6200,N_7109);
xor U8901 (N_8901,N_6789,N_7522);
xnor U8902 (N_8902,N_6079,N_6937);
nor U8903 (N_8903,N_6701,N_7198);
and U8904 (N_8904,N_7855,N_6813);
nor U8905 (N_8905,N_6400,N_7304);
and U8906 (N_8906,N_7707,N_6344);
or U8907 (N_8907,N_6961,N_7357);
nand U8908 (N_8908,N_6854,N_7174);
nor U8909 (N_8909,N_7465,N_6873);
nand U8910 (N_8910,N_7890,N_7798);
nor U8911 (N_8911,N_7640,N_7380);
nand U8912 (N_8912,N_6376,N_7677);
nand U8913 (N_8913,N_6154,N_7552);
or U8914 (N_8914,N_7944,N_7070);
nand U8915 (N_8915,N_7282,N_7002);
and U8916 (N_8916,N_6443,N_7965);
nand U8917 (N_8917,N_6358,N_6639);
and U8918 (N_8918,N_6067,N_6985);
xor U8919 (N_8919,N_6063,N_7935);
xnor U8920 (N_8920,N_6407,N_7004);
nand U8921 (N_8921,N_7175,N_6185);
nor U8922 (N_8922,N_6918,N_7118);
and U8923 (N_8923,N_7970,N_6911);
xor U8924 (N_8924,N_6100,N_6295);
nor U8925 (N_8925,N_6830,N_6353);
and U8926 (N_8926,N_7683,N_6383);
or U8927 (N_8927,N_6299,N_7090);
or U8928 (N_8928,N_7347,N_6996);
and U8929 (N_8929,N_6676,N_6050);
and U8930 (N_8930,N_7535,N_6884);
nand U8931 (N_8931,N_7489,N_7613);
nor U8932 (N_8932,N_6641,N_7598);
nor U8933 (N_8933,N_7125,N_6487);
or U8934 (N_8934,N_7385,N_6969);
or U8935 (N_8935,N_7967,N_6012);
nor U8936 (N_8936,N_7286,N_7048);
or U8937 (N_8937,N_6981,N_6431);
and U8938 (N_8938,N_7402,N_7498);
nand U8939 (N_8939,N_7490,N_6412);
or U8940 (N_8940,N_6648,N_6110);
or U8941 (N_8941,N_7251,N_6259);
or U8942 (N_8942,N_7950,N_6064);
nor U8943 (N_8943,N_6119,N_6548);
nor U8944 (N_8944,N_7332,N_6444);
nand U8945 (N_8945,N_6543,N_7793);
and U8946 (N_8946,N_7758,N_7407);
nor U8947 (N_8947,N_6198,N_7288);
nand U8948 (N_8948,N_6642,N_6318);
xor U8949 (N_8949,N_6729,N_7073);
and U8950 (N_8950,N_6698,N_7756);
or U8951 (N_8951,N_7427,N_7916);
and U8952 (N_8952,N_7275,N_6222);
or U8953 (N_8953,N_7650,N_7000);
nand U8954 (N_8954,N_6125,N_7900);
and U8955 (N_8955,N_7591,N_6053);
nor U8956 (N_8956,N_6907,N_7866);
or U8957 (N_8957,N_7727,N_6661);
and U8958 (N_8958,N_6692,N_6929);
nand U8959 (N_8959,N_6234,N_6776);
or U8960 (N_8960,N_7624,N_6382);
nand U8961 (N_8961,N_7836,N_6629);
nor U8962 (N_8962,N_7213,N_7292);
nand U8963 (N_8963,N_7920,N_7459);
and U8964 (N_8964,N_7025,N_7058);
and U8965 (N_8965,N_7429,N_6283);
nand U8966 (N_8966,N_7232,N_6270);
nor U8967 (N_8967,N_6449,N_6689);
nand U8968 (N_8968,N_7219,N_6215);
nand U8969 (N_8969,N_7673,N_7389);
nand U8970 (N_8970,N_7958,N_6942);
xnor U8971 (N_8971,N_6935,N_7734);
nor U8972 (N_8972,N_7721,N_7503);
nor U8973 (N_8973,N_6381,N_6491);
nand U8974 (N_8974,N_6764,N_7217);
and U8975 (N_8975,N_7149,N_6021);
and U8976 (N_8976,N_7001,N_6700);
and U8977 (N_8977,N_7290,N_6473);
nor U8978 (N_8978,N_6897,N_6022);
nor U8979 (N_8979,N_7016,N_6037);
xor U8980 (N_8980,N_7314,N_6551);
xnor U8981 (N_8981,N_7725,N_7575);
nor U8982 (N_8982,N_6621,N_6782);
nand U8983 (N_8983,N_7539,N_7417);
nor U8984 (N_8984,N_6744,N_6016);
and U8985 (N_8985,N_7394,N_7507);
nand U8986 (N_8986,N_7192,N_6513);
nand U8987 (N_8987,N_6538,N_6838);
and U8988 (N_8988,N_7529,N_6514);
nor U8989 (N_8989,N_6936,N_7506);
or U8990 (N_8990,N_6706,N_7421);
nor U8991 (N_8991,N_7708,N_7400);
or U8992 (N_8992,N_7376,N_7845);
and U8993 (N_8993,N_7105,N_6984);
xor U8994 (N_8994,N_6718,N_7704);
nor U8995 (N_8995,N_6093,N_7998);
and U8996 (N_8996,N_6880,N_7511);
and U8997 (N_8997,N_6652,N_6008);
nor U8998 (N_8998,N_6561,N_7875);
and U8999 (N_8999,N_6246,N_6988);
nor U9000 (N_9000,N_6678,N_6123);
nand U9001 (N_9001,N_6346,N_6028);
and U9002 (N_9002,N_6673,N_6607);
or U9003 (N_9003,N_7605,N_6802);
xor U9004 (N_9004,N_6948,N_6090);
xnor U9005 (N_9005,N_6386,N_7232);
nor U9006 (N_9006,N_7092,N_7626);
nand U9007 (N_9007,N_6544,N_6443);
nand U9008 (N_9008,N_6948,N_6038);
xor U9009 (N_9009,N_6883,N_6730);
or U9010 (N_9010,N_7125,N_7857);
nor U9011 (N_9011,N_7046,N_6410);
nor U9012 (N_9012,N_6322,N_7209);
and U9013 (N_9013,N_7268,N_6933);
nand U9014 (N_9014,N_7532,N_7554);
xor U9015 (N_9015,N_6110,N_7378);
nand U9016 (N_9016,N_6153,N_7089);
xnor U9017 (N_9017,N_7691,N_7348);
or U9018 (N_9018,N_7231,N_6780);
or U9019 (N_9019,N_6315,N_7292);
and U9020 (N_9020,N_6106,N_7140);
or U9021 (N_9021,N_6708,N_7765);
xnor U9022 (N_9022,N_7520,N_6418);
and U9023 (N_9023,N_7029,N_6122);
nor U9024 (N_9024,N_6063,N_6622);
and U9025 (N_9025,N_6250,N_6182);
xnor U9026 (N_9026,N_7139,N_6505);
or U9027 (N_9027,N_7990,N_7288);
nor U9028 (N_9028,N_6809,N_6045);
and U9029 (N_9029,N_6389,N_7334);
xnor U9030 (N_9030,N_7509,N_7283);
nor U9031 (N_9031,N_6341,N_6464);
or U9032 (N_9032,N_6954,N_6651);
nand U9033 (N_9033,N_6839,N_6340);
xnor U9034 (N_9034,N_7556,N_6295);
or U9035 (N_9035,N_7015,N_7283);
and U9036 (N_9036,N_6703,N_6781);
or U9037 (N_9037,N_7301,N_6840);
and U9038 (N_9038,N_6378,N_6861);
or U9039 (N_9039,N_7531,N_6972);
xor U9040 (N_9040,N_6501,N_6618);
and U9041 (N_9041,N_7804,N_7148);
nor U9042 (N_9042,N_7583,N_7175);
nor U9043 (N_9043,N_6801,N_6768);
and U9044 (N_9044,N_7420,N_7839);
nor U9045 (N_9045,N_6680,N_7955);
and U9046 (N_9046,N_6258,N_6697);
xnor U9047 (N_9047,N_6038,N_7275);
nor U9048 (N_9048,N_7192,N_7126);
nor U9049 (N_9049,N_7627,N_6705);
xor U9050 (N_9050,N_7590,N_7682);
or U9051 (N_9051,N_6753,N_7816);
and U9052 (N_9052,N_7840,N_7329);
nor U9053 (N_9053,N_6458,N_6017);
or U9054 (N_9054,N_7624,N_6431);
or U9055 (N_9055,N_6358,N_7608);
xnor U9056 (N_9056,N_7668,N_7140);
or U9057 (N_9057,N_7796,N_7497);
nand U9058 (N_9058,N_7922,N_7951);
xor U9059 (N_9059,N_6972,N_7771);
nand U9060 (N_9060,N_7879,N_7144);
or U9061 (N_9061,N_7027,N_6389);
or U9062 (N_9062,N_6669,N_6101);
or U9063 (N_9063,N_7602,N_6127);
nand U9064 (N_9064,N_6808,N_6205);
nand U9065 (N_9065,N_7242,N_7493);
nor U9066 (N_9066,N_7949,N_6370);
and U9067 (N_9067,N_7767,N_7408);
xor U9068 (N_9068,N_6462,N_6689);
nand U9069 (N_9069,N_7219,N_6737);
nand U9070 (N_9070,N_7298,N_6735);
xor U9071 (N_9071,N_6542,N_7871);
or U9072 (N_9072,N_7421,N_7720);
nand U9073 (N_9073,N_7949,N_6537);
or U9074 (N_9074,N_7624,N_7851);
or U9075 (N_9075,N_7936,N_7288);
nor U9076 (N_9076,N_6928,N_7284);
or U9077 (N_9077,N_7997,N_6801);
nor U9078 (N_9078,N_7054,N_6454);
nand U9079 (N_9079,N_6951,N_6780);
nand U9080 (N_9080,N_6466,N_6876);
nand U9081 (N_9081,N_7966,N_6425);
or U9082 (N_9082,N_6758,N_6078);
nor U9083 (N_9083,N_7203,N_6365);
or U9084 (N_9084,N_6924,N_6179);
nand U9085 (N_9085,N_6356,N_7420);
and U9086 (N_9086,N_7636,N_7829);
xor U9087 (N_9087,N_7840,N_6658);
xnor U9088 (N_9088,N_6007,N_7074);
or U9089 (N_9089,N_6149,N_7540);
or U9090 (N_9090,N_7717,N_7112);
xnor U9091 (N_9091,N_7177,N_6638);
or U9092 (N_9092,N_6111,N_7791);
xor U9093 (N_9093,N_6540,N_7441);
and U9094 (N_9094,N_6347,N_6471);
xor U9095 (N_9095,N_7771,N_6349);
and U9096 (N_9096,N_7237,N_7436);
nand U9097 (N_9097,N_6221,N_7126);
or U9098 (N_9098,N_7624,N_7888);
nand U9099 (N_9099,N_6313,N_7372);
and U9100 (N_9100,N_6733,N_7781);
nand U9101 (N_9101,N_7463,N_7376);
nand U9102 (N_9102,N_6493,N_6922);
and U9103 (N_9103,N_6024,N_6786);
nor U9104 (N_9104,N_7053,N_6497);
nor U9105 (N_9105,N_7544,N_7999);
and U9106 (N_9106,N_6498,N_6476);
and U9107 (N_9107,N_7193,N_7685);
or U9108 (N_9108,N_6182,N_6775);
xnor U9109 (N_9109,N_7425,N_7075);
nor U9110 (N_9110,N_6822,N_7720);
xnor U9111 (N_9111,N_7923,N_6367);
and U9112 (N_9112,N_7964,N_7164);
nand U9113 (N_9113,N_7366,N_6537);
and U9114 (N_9114,N_6262,N_6692);
or U9115 (N_9115,N_6927,N_7574);
nand U9116 (N_9116,N_7016,N_7705);
and U9117 (N_9117,N_7926,N_7233);
nor U9118 (N_9118,N_6365,N_6661);
nand U9119 (N_9119,N_7625,N_7620);
xor U9120 (N_9120,N_6914,N_6401);
xnor U9121 (N_9121,N_7141,N_7740);
nand U9122 (N_9122,N_6808,N_7946);
nand U9123 (N_9123,N_7028,N_7812);
and U9124 (N_9124,N_6092,N_6118);
and U9125 (N_9125,N_7883,N_7208);
nand U9126 (N_9126,N_7548,N_6137);
xnor U9127 (N_9127,N_7706,N_7970);
nand U9128 (N_9128,N_6672,N_6927);
xnor U9129 (N_9129,N_6257,N_6494);
xnor U9130 (N_9130,N_7799,N_7750);
nor U9131 (N_9131,N_7569,N_6504);
or U9132 (N_9132,N_7805,N_7982);
xor U9133 (N_9133,N_6924,N_7953);
nor U9134 (N_9134,N_7782,N_6085);
or U9135 (N_9135,N_6383,N_7473);
or U9136 (N_9136,N_7008,N_7696);
nand U9137 (N_9137,N_6906,N_6896);
xor U9138 (N_9138,N_6251,N_6739);
xnor U9139 (N_9139,N_6716,N_6213);
nand U9140 (N_9140,N_7365,N_7597);
and U9141 (N_9141,N_7000,N_6488);
nand U9142 (N_9142,N_7596,N_7951);
xor U9143 (N_9143,N_6305,N_7653);
or U9144 (N_9144,N_7303,N_7314);
xnor U9145 (N_9145,N_7441,N_7189);
and U9146 (N_9146,N_7598,N_7895);
nor U9147 (N_9147,N_7943,N_7939);
or U9148 (N_9148,N_7982,N_7257);
nor U9149 (N_9149,N_6550,N_7649);
or U9150 (N_9150,N_7275,N_7134);
xnor U9151 (N_9151,N_7723,N_6483);
or U9152 (N_9152,N_7064,N_7480);
xnor U9153 (N_9153,N_7318,N_6768);
nor U9154 (N_9154,N_7743,N_6383);
nor U9155 (N_9155,N_7424,N_6539);
xnor U9156 (N_9156,N_6949,N_6701);
xor U9157 (N_9157,N_6805,N_7025);
nor U9158 (N_9158,N_6304,N_6146);
xor U9159 (N_9159,N_6763,N_7699);
and U9160 (N_9160,N_7355,N_6187);
nand U9161 (N_9161,N_6021,N_6671);
nor U9162 (N_9162,N_7643,N_6729);
nor U9163 (N_9163,N_7954,N_7352);
xor U9164 (N_9164,N_6165,N_6403);
nor U9165 (N_9165,N_6963,N_6335);
and U9166 (N_9166,N_7888,N_7082);
or U9167 (N_9167,N_6859,N_6487);
and U9168 (N_9168,N_6906,N_7838);
nor U9169 (N_9169,N_7870,N_7590);
and U9170 (N_9170,N_7549,N_6619);
xnor U9171 (N_9171,N_6305,N_7742);
xnor U9172 (N_9172,N_6015,N_7063);
and U9173 (N_9173,N_7241,N_6626);
or U9174 (N_9174,N_7812,N_7105);
nand U9175 (N_9175,N_7609,N_7146);
or U9176 (N_9176,N_6027,N_6156);
and U9177 (N_9177,N_7542,N_6558);
xor U9178 (N_9178,N_7160,N_7538);
nand U9179 (N_9179,N_6237,N_6305);
and U9180 (N_9180,N_6880,N_7038);
nand U9181 (N_9181,N_6902,N_6821);
nand U9182 (N_9182,N_6344,N_7672);
and U9183 (N_9183,N_6500,N_6810);
nand U9184 (N_9184,N_7286,N_7496);
or U9185 (N_9185,N_6962,N_7651);
or U9186 (N_9186,N_6704,N_7411);
nor U9187 (N_9187,N_6199,N_6809);
nor U9188 (N_9188,N_7460,N_7001);
nand U9189 (N_9189,N_6662,N_7931);
xnor U9190 (N_9190,N_7324,N_7659);
nand U9191 (N_9191,N_7881,N_6221);
nor U9192 (N_9192,N_6167,N_7593);
nand U9193 (N_9193,N_7049,N_6574);
nor U9194 (N_9194,N_7447,N_6970);
or U9195 (N_9195,N_7617,N_6532);
or U9196 (N_9196,N_7137,N_6089);
or U9197 (N_9197,N_7133,N_7048);
nor U9198 (N_9198,N_6725,N_6039);
nand U9199 (N_9199,N_7701,N_6648);
nand U9200 (N_9200,N_6778,N_7361);
xor U9201 (N_9201,N_6523,N_6652);
nand U9202 (N_9202,N_7935,N_7229);
nor U9203 (N_9203,N_6515,N_6730);
or U9204 (N_9204,N_7269,N_7406);
nor U9205 (N_9205,N_6151,N_7472);
nor U9206 (N_9206,N_7276,N_7446);
and U9207 (N_9207,N_7632,N_6693);
nand U9208 (N_9208,N_7462,N_7534);
or U9209 (N_9209,N_7921,N_7458);
nand U9210 (N_9210,N_6345,N_7056);
nand U9211 (N_9211,N_6079,N_7751);
nor U9212 (N_9212,N_7784,N_6194);
xor U9213 (N_9213,N_6820,N_7738);
nand U9214 (N_9214,N_7908,N_7678);
nor U9215 (N_9215,N_6291,N_6485);
xor U9216 (N_9216,N_6801,N_6134);
or U9217 (N_9217,N_6932,N_7088);
nor U9218 (N_9218,N_7927,N_7867);
nor U9219 (N_9219,N_6661,N_6300);
or U9220 (N_9220,N_6790,N_7953);
nand U9221 (N_9221,N_6457,N_6966);
nor U9222 (N_9222,N_7138,N_6535);
and U9223 (N_9223,N_6393,N_7253);
nor U9224 (N_9224,N_7478,N_7932);
or U9225 (N_9225,N_7219,N_7202);
xor U9226 (N_9226,N_6536,N_7293);
and U9227 (N_9227,N_7117,N_7466);
nand U9228 (N_9228,N_7896,N_6101);
xor U9229 (N_9229,N_6864,N_7099);
xnor U9230 (N_9230,N_7284,N_6432);
or U9231 (N_9231,N_7170,N_6727);
nor U9232 (N_9232,N_6202,N_6512);
nand U9233 (N_9233,N_7294,N_6514);
xnor U9234 (N_9234,N_6115,N_7826);
nand U9235 (N_9235,N_6151,N_6713);
nand U9236 (N_9236,N_7739,N_6080);
nand U9237 (N_9237,N_7196,N_6223);
or U9238 (N_9238,N_6585,N_7091);
nand U9239 (N_9239,N_6955,N_7835);
and U9240 (N_9240,N_7226,N_6384);
or U9241 (N_9241,N_7146,N_7475);
xnor U9242 (N_9242,N_7288,N_7499);
and U9243 (N_9243,N_6454,N_7342);
or U9244 (N_9244,N_7440,N_6764);
or U9245 (N_9245,N_7432,N_6494);
nand U9246 (N_9246,N_6007,N_6869);
nand U9247 (N_9247,N_7309,N_6623);
nor U9248 (N_9248,N_6407,N_7807);
nor U9249 (N_9249,N_7777,N_6496);
nor U9250 (N_9250,N_7707,N_6475);
and U9251 (N_9251,N_7689,N_6853);
xor U9252 (N_9252,N_6195,N_6722);
nand U9253 (N_9253,N_6319,N_7047);
nand U9254 (N_9254,N_6599,N_6637);
nor U9255 (N_9255,N_6529,N_7944);
and U9256 (N_9256,N_6295,N_7200);
nor U9257 (N_9257,N_7111,N_6051);
and U9258 (N_9258,N_6879,N_7190);
nand U9259 (N_9259,N_6870,N_7564);
or U9260 (N_9260,N_6812,N_7949);
nor U9261 (N_9261,N_6352,N_7076);
nand U9262 (N_9262,N_7608,N_7374);
and U9263 (N_9263,N_6230,N_7042);
and U9264 (N_9264,N_6210,N_6031);
and U9265 (N_9265,N_7686,N_7546);
or U9266 (N_9266,N_6042,N_7271);
and U9267 (N_9267,N_6584,N_7327);
or U9268 (N_9268,N_7834,N_6507);
nand U9269 (N_9269,N_6366,N_7219);
or U9270 (N_9270,N_6555,N_7295);
nand U9271 (N_9271,N_6108,N_7245);
and U9272 (N_9272,N_6923,N_6092);
and U9273 (N_9273,N_6322,N_7053);
nand U9274 (N_9274,N_7694,N_7490);
xnor U9275 (N_9275,N_6816,N_6701);
or U9276 (N_9276,N_7362,N_7058);
nand U9277 (N_9277,N_7917,N_7196);
and U9278 (N_9278,N_6586,N_6829);
or U9279 (N_9279,N_7822,N_7256);
nor U9280 (N_9280,N_6611,N_7446);
nor U9281 (N_9281,N_6595,N_6930);
nand U9282 (N_9282,N_6786,N_7017);
nor U9283 (N_9283,N_6730,N_7546);
nand U9284 (N_9284,N_6198,N_6809);
nand U9285 (N_9285,N_6737,N_7362);
xor U9286 (N_9286,N_7146,N_6242);
or U9287 (N_9287,N_6940,N_7810);
and U9288 (N_9288,N_6720,N_7225);
nor U9289 (N_9289,N_7903,N_7396);
xor U9290 (N_9290,N_7429,N_6625);
nand U9291 (N_9291,N_7954,N_7820);
or U9292 (N_9292,N_7554,N_6933);
nand U9293 (N_9293,N_6655,N_7765);
and U9294 (N_9294,N_7222,N_7263);
nor U9295 (N_9295,N_6091,N_7284);
xor U9296 (N_9296,N_6964,N_7212);
xnor U9297 (N_9297,N_6245,N_6017);
nand U9298 (N_9298,N_6237,N_7303);
nor U9299 (N_9299,N_7204,N_7670);
nor U9300 (N_9300,N_7527,N_7536);
and U9301 (N_9301,N_7094,N_7723);
or U9302 (N_9302,N_7518,N_6106);
and U9303 (N_9303,N_6918,N_6907);
or U9304 (N_9304,N_7581,N_6039);
nand U9305 (N_9305,N_6770,N_6475);
nand U9306 (N_9306,N_6434,N_7925);
or U9307 (N_9307,N_7853,N_6007);
nor U9308 (N_9308,N_6333,N_7952);
or U9309 (N_9309,N_6813,N_7487);
and U9310 (N_9310,N_6603,N_7587);
and U9311 (N_9311,N_7336,N_6478);
nand U9312 (N_9312,N_6560,N_6983);
nor U9313 (N_9313,N_6040,N_6569);
and U9314 (N_9314,N_6976,N_6386);
and U9315 (N_9315,N_7347,N_7675);
nand U9316 (N_9316,N_6512,N_7804);
nor U9317 (N_9317,N_6598,N_6963);
and U9318 (N_9318,N_6634,N_6880);
nor U9319 (N_9319,N_7216,N_7546);
nor U9320 (N_9320,N_6824,N_7980);
xor U9321 (N_9321,N_7693,N_7138);
or U9322 (N_9322,N_6069,N_6347);
xor U9323 (N_9323,N_6219,N_6054);
nor U9324 (N_9324,N_6706,N_7631);
xnor U9325 (N_9325,N_6137,N_6260);
nand U9326 (N_9326,N_7270,N_6670);
xor U9327 (N_9327,N_7857,N_7556);
xnor U9328 (N_9328,N_6308,N_6909);
nand U9329 (N_9329,N_7604,N_7427);
and U9330 (N_9330,N_6285,N_7889);
nor U9331 (N_9331,N_7399,N_7183);
xor U9332 (N_9332,N_7291,N_6790);
nand U9333 (N_9333,N_7270,N_6928);
nand U9334 (N_9334,N_7560,N_6870);
or U9335 (N_9335,N_6755,N_7667);
nand U9336 (N_9336,N_6110,N_7869);
or U9337 (N_9337,N_6524,N_7588);
nor U9338 (N_9338,N_7564,N_7837);
xnor U9339 (N_9339,N_7504,N_6535);
nand U9340 (N_9340,N_6448,N_6345);
xnor U9341 (N_9341,N_7671,N_6698);
nand U9342 (N_9342,N_6164,N_6417);
nand U9343 (N_9343,N_7595,N_7502);
nand U9344 (N_9344,N_6976,N_6139);
nand U9345 (N_9345,N_6478,N_6397);
xor U9346 (N_9346,N_7972,N_6821);
and U9347 (N_9347,N_7471,N_7720);
or U9348 (N_9348,N_6060,N_6229);
or U9349 (N_9349,N_7245,N_6437);
and U9350 (N_9350,N_7672,N_6532);
xnor U9351 (N_9351,N_6046,N_7046);
nor U9352 (N_9352,N_7855,N_7839);
or U9353 (N_9353,N_6370,N_7632);
xor U9354 (N_9354,N_6985,N_7369);
and U9355 (N_9355,N_6958,N_6741);
nand U9356 (N_9356,N_7459,N_7881);
nor U9357 (N_9357,N_6896,N_6226);
and U9358 (N_9358,N_6051,N_7947);
xor U9359 (N_9359,N_6829,N_6154);
nand U9360 (N_9360,N_6166,N_7982);
or U9361 (N_9361,N_6775,N_6250);
and U9362 (N_9362,N_7954,N_6213);
and U9363 (N_9363,N_7263,N_6378);
or U9364 (N_9364,N_7549,N_7626);
nand U9365 (N_9365,N_7377,N_7695);
nand U9366 (N_9366,N_7385,N_6131);
or U9367 (N_9367,N_7335,N_7296);
nand U9368 (N_9368,N_7616,N_7358);
xnor U9369 (N_9369,N_7827,N_6302);
nor U9370 (N_9370,N_6045,N_6991);
xnor U9371 (N_9371,N_7140,N_7000);
and U9372 (N_9372,N_7857,N_6934);
nand U9373 (N_9373,N_6964,N_7449);
and U9374 (N_9374,N_6254,N_6690);
or U9375 (N_9375,N_6450,N_7373);
xor U9376 (N_9376,N_7437,N_7791);
and U9377 (N_9377,N_7171,N_6830);
and U9378 (N_9378,N_6596,N_7465);
xor U9379 (N_9379,N_7334,N_7650);
nor U9380 (N_9380,N_6702,N_7521);
nor U9381 (N_9381,N_7155,N_6380);
nor U9382 (N_9382,N_6073,N_6335);
nand U9383 (N_9383,N_6996,N_7581);
and U9384 (N_9384,N_6685,N_6968);
nor U9385 (N_9385,N_6487,N_6706);
nor U9386 (N_9386,N_7647,N_7864);
or U9387 (N_9387,N_7839,N_7482);
or U9388 (N_9388,N_6289,N_7849);
nor U9389 (N_9389,N_6793,N_7475);
xnor U9390 (N_9390,N_6434,N_7337);
xnor U9391 (N_9391,N_6041,N_6781);
and U9392 (N_9392,N_6119,N_7933);
or U9393 (N_9393,N_7678,N_7708);
and U9394 (N_9394,N_7449,N_6031);
nand U9395 (N_9395,N_6751,N_6838);
and U9396 (N_9396,N_7367,N_7998);
nor U9397 (N_9397,N_7183,N_7921);
nand U9398 (N_9398,N_7665,N_6325);
or U9399 (N_9399,N_7954,N_6143);
or U9400 (N_9400,N_7813,N_7012);
nor U9401 (N_9401,N_7024,N_6420);
or U9402 (N_9402,N_7804,N_7046);
nor U9403 (N_9403,N_7583,N_7239);
nor U9404 (N_9404,N_6802,N_6002);
or U9405 (N_9405,N_7216,N_7263);
nand U9406 (N_9406,N_7049,N_7051);
or U9407 (N_9407,N_7396,N_6229);
nand U9408 (N_9408,N_7085,N_7704);
and U9409 (N_9409,N_6039,N_6189);
nor U9410 (N_9410,N_7678,N_7059);
and U9411 (N_9411,N_7958,N_6194);
and U9412 (N_9412,N_6869,N_6264);
nor U9413 (N_9413,N_6408,N_7764);
or U9414 (N_9414,N_6987,N_6922);
nor U9415 (N_9415,N_7344,N_6925);
nor U9416 (N_9416,N_6909,N_7572);
nor U9417 (N_9417,N_6043,N_6987);
or U9418 (N_9418,N_6293,N_7904);
or U9419 (N_9419,N_6656,N_7797);
nor U9420 (N_9420,N_6987,N_6437);
xor U9421 (N_9421,N_7382,N_7898);
nand U9422 (N_9422,N_7267,N_6454);
or U9423 (N_9423,N_7260,N_6179);
xor U9424 (N_9424,N_6912,N_6169);
xor U9425 (N_9425,N_7792,N_6756);
nand U9426 (N_9426,N_6921,N_7629);
xor U9427 (N_9427,N_6994,N_7882);
or U9428 (N_9428,N_7364,N_6222);
and U9429 (N_9429,N_7696,N_7158);
xor U9430 (N_9430,N_7740,N_6568);
nor U9431 (N_9431,N_7230,N_6048);
or U9432 (N_9432,N_6660,N_7789);
and U9433 (N_9433,N_7489,N_7560);
or U9434 (N_9434,N_7306,N_6915);
or U9435 (N_9435,N_7059,N_7756);
nand U9436 (N_9436,N_7478,N_7560);
nand U9437 (N_9437,N_7370,N_6424);
and U9438 (N_9438,N_6952,N_6534);
xor U9439 (N_9439,N_7546,N_7489);
and U9440 (N_9440,N_6163,N_7944);
xor U9441 (N_9441,N_7405,N_6216);
or U9442 (N_9442,N_7214,N_6398);
or U9443 (N_9443,N_7428,N_6282);
nand U9444 (N_9444,N_6314,N_6384);
nor U9445 (N_9445,N_6225,N_7759);
nand U9446 (N_9446,N_7047,N_7871);
xnor U9447 (N_9447,N_7738,N_7727);
nand U9448 (N_9448,N_6631,N_6609);
nand U9449 (N_9449,N_7445,N_6707);
nor U9450 (N_9450,N_6345,N_7265);
nor U9451 (N_9451,N_7367,N_6404);
and U9452 (N_9452,N_7264,N_6370);
and U9453 (N_9453,N_7129,N_7285);
nor U9454 (N_9454,N_7227,N_7595);
nor U9455 (N_9455,N_6727,N_7986);
nor U9456 (N_9456,N_7924,N_6362);
and U9457 (N_9457,N_6661,N_6554);
nor U9458 (N_9458,N_7433,N_6719);
nand U9459 (N_9459,N_7702,N_6151);
nand U9460 (N_9460,N_6889,N_6104);
xnor U9461 (N_9461,N_6862,N_7153);
or U9462 (N_9462,N_7588,N_7581);
and U9463 (N_9463,N_6662,N_6826);
nand U9464 (N_9464,N_7465,N_7875);
xnor U9465 (N_9465,N_6193,N_7142);
and U9466 (N_9466,N_7194,N_6640);
nor U9467 (N_9467,N_7955,N_7190);
nor U9468 (N_9468,N_7935,N_7995);
nor U9469 (N_9469,N_6163,N_7374);
or U9470 (N_9470,N_7975,N_6370);
nand U9471 (N_9471,N_7188,N_6298);
nor U9472 (N_9472,N_7915,N_6758);
xor U9473 (N_9473,N_6402,N_7953);
or U9474 (N_9474,N_7261,N_6460);
or U9475 (N_9475,N_6792,N_7776);
nor U9476 (N_9476,N_7721,N_7282);
and U9477 (N_9477,N_7661,N_7543);
nor U9478 (N_9478,N_7265,N_6339);
xor U9479 (N_9479,N_6991,N_7306);
nor U9480 (N_9480,N_6435,N_6104);
or U9481 (N_9481,N_7767,N_7003);
xnor U9482 (N_9482,N_7417,N_6747);
nand U9483 (N_9483,N_6977,N_7341);
or U9484 (N_9484,N_7052,N_7081);
and U9485 (N_9485,N_7210,N_6707);
xnor U9486 (N_9486,N_6930,N_6172);
xnor U9487 (N_9487,N_7434,N_6115);
and U9488 (N_9488,N_7520,N_6248);
nand U9489 (N_9489,N_7509,N_6211);
and U9490 (N_9490,N_6623,N_7781);
and U9491 (N_9491,N_6700,N_6663);
or U9492 (N_9492,N_6244,N_6175);
and U9493 (N_9493,N_6674,N_6547);
xnor U9494 (N_9494,N_6715,N_6926);
nand U9495 (N_9495,N_6864,N_6518);
and U9496 (N_9496,N_6971,N_6752);
or U9497 (N_9497,N_6474,N_6546);
or U9498 (N_9498,N_6392,N_7847);
nand U9499 (N_9499,N_7555,N_6546);
nand U9500 (N_9500,N_7986,N_6867);
nor U9501 (N_9501,N_6990,N_6540);
xor U9502 (N_9502,N_6866,N_6230);
and U9503 (N_9503,N_6991,N_7799);
and U9504 (N_9504,N_6109,N_6860);
nand U9505 (N_9505,N_7241,N_6445);
nand U9506 (N_9506,N_7586,N_6380);
nor U9507 (N_9507,N_6090,N_7770);
nand U9508 (N_9508,N_7546,N_7932);
or U9509 (N_9509,N_7938,N_6278);
nor U9510 (N_9510,N_7509,N_7108);
nand U9511 (N_9511,N_7724,N_6245);
nor U9512 (N_9512,N_6450,N_7122);
and U9513 (N_9513,N_6430,N_7798);
or U9514 (N_9514,N_7145,N_7352);
and U9515 (N_9515,N_7463,N_7658);
and U9516 (N_9516,N_6255,N_7171);
xnor U9517 (N_9517,N_6610,N_6641);
nor U9518 (N_9518,N_7783,N_7071);
nand U9519 (N_9519,N_6040,N_6122);
xor U9520 (N_9520,N_7498,N_7054);
xnor U9521 (N_9521,N_6946,N_6741);
or U9522 (N_9522,N_6058,N_7333);
nand U9523 (N_9523,N_6205,N_7452);
or U9524 (N_9524,N_7356,N_6415);
and U9525 (N_9525,N_7791,N_7870);
nor U9526 (N_9526,N_7983,N_6367);
or U9527 (N_9527,N_7775,N_7215);
xnor U9528 (N_9528,N_6618,N_7731);
and U9529 (N_9529,N_7483,N_7843);
nand U9530 (N_9530,N_7725,N_6052);
or U9531 (N_9531,N_6627,N_7230);
nor U9532 (N_9532,N_7698,N_6027);
xnor U9533 (N_9533,N_7742,N_7203);
nand U9534 (N_9534,N_7281,N_7985);
nor U9535 (N_9535,N_7909,N_7127);
nand U9536 (N_9536,N_6850,N_7847);
xnor U9537 (N_9537,N_6533,N_6282);
and U9538 (N_9538,N_6252,N_6936);
or U9539 (N_9539,N_7182,N_6464);
and U9540 (N_9540,N_6184,N_6689);
or U9541 (N_9541,N_7130,N_7100);
or U9542 (N_9542,N_7142,N_7334);
nor U9543 (N_9543,N_7734,N_6563);
nor U9544 (N_9544,N_7925,N_7086);
xor U9545 (N_9545,N_7758,N_7980);
and U9546 (N_9546,N_6207,N_7546);
or U9547 (N_9547,N_6282,N_6314);
nand U9548 (N_9548,N_6167,N_7769);
xnor U9549 (N_9549,N_6933,N_6924);
xor U9550 (N_9550,N_6004,N_7517);
nor U9551 (N_9551,N_7406,N_6315);
and U9552 (N_9552,N_7852,N_7795);
or U9553 (N_9553,N_6428,N_6547);
xnor U9554 (N_9554,N_6490,N_6570);
nor U9555 (N_9555,N_7096,N_7188);
nor U9556 (N_9556,N_6290,N_6977);
nor U9557 (N_9557,N_6875,N_7247);
nand U9558 (N_9558,N_6824,N_7122);
xor U9559 (N_9559,N_7423,N_7453);
nand U9560 (N_9560,N_7535,N_6447);
and U9561 (N_9561,N_6614,N_7034);
nor U9562 (N_9562,N_6613,N_7972);
nor U9563 (N_9563,N_7660,N_7991);
and U9564 (N_9564,N_6587,N_6852);
xnor U9565 (N_9565,N_6328,N_7099);
xnor U9566 (N_9566,N_7918,N_7839);
xnor U9567 (N_9567,N_6781,N_7925);
nand U9568 (N_9568,N_6525,N_7531);
nand U9569 (N_9569,N_7111,N_7574);
nor U9570 (N_9570,N_6092,N_7744);
and U9571 (N_9571,N_7551,N_7926);
or U9572 (N_9572,N_7594,N_7390);
or U9573 (N_9573,N_6921,N_7452);
nand U9574 (N_9574,N_7780,N_7989);
and U9575 (N_9575,N_6418,N_6663);
or U9576 (N_9576,N_7548,N_6986);
nand U9577 (N_9577,N_7362,N_7272);
xnor U9578 (N_9578,N_7524,N_7143);
nand U9579 (N_9579,N_7433,N_7997);
and U9580 (N_9580,N_7623,N_7752);
nand U9581 (N_9581,N_7703,N_7392);
xnor U9582 (N_9582,N_6326,N_7658);
nand U9583 (N_9583,N_7978,N_7063);
and U9584 (N_9584,N_6075,N_6531);
nand U9585 (N_9585,N_6204,N_7268);
xnor U9586 (N_9586,N_6544,N_6236);
nor U9587 (N_9587,N_6116,N_6052);
or U9588 (N_9588,N_7869,N_7735);
xnor U9589 (N_9589,N_6027,N_6461);
xnor U9590 (N_9590,N_6026,N_6382);
nand U9591 (N_9591,N_7567,N_6248);
xor U9592 (N_9592,N_6247,N_7013);
and U9593 (N_9593,N_7159,N_6857);
xor U9594 (N_9594,N_7975,N_7277);
xor U9595 (N_9595,N_7689,N_6788);
nor U9596 (N_9596,N_6008,N_7681);
nor U9597 (N_9597,N_7959,N_6169);
and U9598 (N_9598,N_7267,N_7050);
xnor U9599 (N_9599,N_6940,N_6120);
nand U9600 (N_9600,N_6436,N_6461);
xnor U9601 (N_9601,N_7654,N_7881);
nand U9602 (N_9602,N_7109,N_7415);
xnor U9603 (N_9603,N_7498,N_6299);
and U9604 (N_9604,N_7766,N_7364);
or U9605 (N_9605,N_6297,N_7595);
and U9606 (N_9606,N_7365,N_6085);
nor U9607 (N_9607,N_6689,N_7043);
and U9608 (N_9608,N_6476,N_7787);
or U9609 (N_9609,N_7560,N_6377);
nor U9610 (N_9610,N_6894,N_7740);
nor U9611 (N_9611,N_7537,N_7079);
xnor U9612 (N_9612,N_6547,N_6949);
nand U9613 (N_9613,N_7356,N_6479);
xor U9614 (N_9614,N_7790,N_6050);
and U9615 (N_9615,N_6001,N_6109);
nand U9616 (N_9616,N_7265,N_7155);
or U9617 (N_9617,N_7855,N_7717);
nand U9618 (N_9618,N_7322,N_7994);
or U9619 (N_9619,N_6305,N_7409);
and U9620 (N_9620,N_7578,N_7444);
and U9621 (N_9621,N_6781,N_6652);
or U9622 (N_9622,N_6345,N_7209);
nor U9623 (N_9623,N_6904,N_7026);
nand U9624 (N_9624,N_6752,N_6459);
nor U9625 (N_9625,N_7875,N_6717);
xnor U9626 (N_9626,N_7135,N_7046);
nand U9627 (N_9627,N_6311,N_6573);
nand U9628 (N_9628,N_7859,N_7752);
and U9629 (N_9629,N_7824,N_6905);
or U9630 (N_9630,N_7472,N_7790);
nand U9631 (N_9631,N_6461,N_6371);
nand U9632 (N_9632,N_7645,N_7351);
and U9633 (N_9633,N_6220,N_6717);
xor U9634 (N_9634,N_7567,N_7549);
or U9635 (N_9635,N_7559,N_7406);
and U9636 (N_9636,N_6107,N_6633);
xor U9637 (N_9637,N_6715,N_6674);
and U9638 (N_9638,N_7446,N_7889);
or U9639 (N_9639,N_7131,N_7119);
or U9640 (N_9640,N_7461,N_6912);
or U9641 (N_9641,N_6356,N_7888);
xnor U9642 (N_9642,N_7868,N_6622);
nor U9643 (N_9643,N_6699,N_7383);
nand U9644 (N_9644,N_6356,N_6109);
nand U9645 (N_9645,N_7087,N_6623);
or U9646 (N_9646,N_6756,N_6326);
nand U9647 (N_9647,N_6776,N_7814);
nand U9648 (N_9648,N_7783,N_6943);
nor U9649 (N_9649,N_6209,N_6982);
xnor U9650 (N_9650,N_6782,N_7322);
xnor U9651 (N_9651,N_7683,N_6803);
or U9652 (N_9652,N_7842,N_7643);
or U9653 (N_9653,N_7043,N_7283);
and U9654 (N_9654,N_6912,N_6662);
nor U9655 (N_9655,N_6334,N_7045);
nand U9656 (N_9656,N_7632,N_6618);
nand U9657 (N_9657,N_7614,N_7879);
xor U9658 (N_9658,N_7191,N_6042);
nand U9659 (N_9659,N_7867,N_6612);
or U9660 (N_9660,N_6038,N_7555);
and U9661 (N_9661,N_6045,N_6214);
and U9662 (N_9662,N_7670,N_7232);
xor U9663 (N_9663,N_6547,N_6277);
and U9664 (N_9664,N_6832,N_6921);
nor U9665 (N_9665,N_6765,N_6278);
xor U9666 (N_9666,N_7822,N_6905);
nor U9667 (N_9667,N_7603,N_6992);
xor U9668 (N_9668,N_6208,N_6816);
nor U9669 (N_9669,N_7121,N_7739);
and U9670 (N_9670,N_7550,N_6262);
nand U9671 (N_9671,N_7075,N_7700);
nor U9672 (N_9672,N_7282,N_6072);
nand U9673 (N_9673,N_6046,N_6329);
and U9674 (N_9674,N_6301,N_6958);
and U9675 (N_9675,N_7482,N_7914);
and U9676 (N_9676,N_6151,N_7020);
xor U9677 (N_9677,N_7976,N_6400);
or U9678 (N_9678,N_6698,N_6957);
and U9679 (N_9679,N_6410,N_6272);
nor U9680 (N_9680,N_6161,N_7342);
nor U9681 (N_9681,N_6314,N_7811);
nand U9682 (N_9682,N_6112,N_6577);
nand U9683 (N_9683,N_7231,N_6498);
nor U9684 (N_9684,N_7792,N_6642);
and U9685 (N_9685,N_6734,N_7309);
xnor U9686 (N_9686,N_7607,N_6044);
or U9687 (N_9687,N_6005,N_7574);
or U9688 (N_9688,N_7949,N_6895);
nand U9689 (N_9689,N_6897,N_6606);
xor U9690 (N_9690,N_6779,N_7680);
or U9691 (N_9691,N_7081,N_7960);
nor U9692 (N_9692,N_7350,N_6259);
nand U9693 (N_9693,N_7452,N_6022);
nor U9694 (N_9694,N_6240,N_6996);
nand U9695 (N_9695,N_7723,N_7334);
nand U9696 (N_9696,N_7629,N_6883);
or U9697 (N_9697,N_6310,N_7797);
or U9698 (N_9698,N_7885,N_6727);
and U9699 (N_9699,N_7915,N_6618);
nor U9700 (N_9700,N_6456,N_7438);
and U9701 (N_9701,N_6093,N_6095);
and U9702 (N_9702,N_7611,N_7589);
nand U9703 (N_9703,N_7504,N_6592);
or U9704 (N_9704,N_6476,N_7034);
nor U9705 (N_9705,N_7806,N_7845);
nand U9706 (N_9706,N_7226,N_7979);
nor U9707 (N_9707,N_7410,N_7248);
nand U9708 (N_9708,N_6466,N_6587);
and U9709 (N_9709,N_6465,N_7195);
and U9710 (N_9710,N_7165,N_6145);
nand U9711 (N_9711,N_6395,N_7029);
or U9712 (N_9712,N_6521,N_7877);
nor U9713 (N_9713,N_6623,N_7232);
nand U9714 (N_9714,N_6195,N_6219);
and U9715 (N_9715,N_7748,N_6147);
or U9716 (N_9716,N_7243,N_7202);
xnor U9717 (N_9717,N_6636,N_7212);
nor U9718 (N_9718,N_7434,N_6162);
and U9719 (N_9719,N_7087,N_7703);
nor U9720 (N_9720,N_7275,N_6418);
nor U9721 (N_9721,N_7343,N_7850);
and U9722 (N_9722,N_7957,N_7770);
xnor U9723 (N_9723,N_7663,N_6408);
nand U9724 (N_9724,N_7632,N_6721);
nor U9725 (N_9725,N_6906,N_6050);
nand U9726 (N_9726,N_7849,N_7199);
or U9727 (N_9727,N_7066,N_6200);
or U9728 (N_9728,N_6909,N_6237);
nand U9729 (N_9729,N_6795,N_6943);
xor U9730 (N_9730,N_6083,N_7366);
xnor U9731 (N_9731,N_6219,N_7813);
xor U9732 (N_9732,N_6757,N_6906);
xnor U9733 (N_9733,N_7123,N_6804);
or U9734 (N_9734,N_7075,N_7952);
xor U9735 (N_9735,N_6545,N_7141);
nand U9736 (N_9736,N_7019,N_6422);
or U9737 (N_9737,N_7620,N_6573);
nor U9738 (N_9738,N_6351,N_7195);
nor U9739 (N_9739,N_6743,N_7111);
and U9740 (N_9740,N_7408,N_7611);
nand U9741 (N_9741,N_7412,N_6839);
or U9742 (N_9742,N_7675,N_7924);
xor U9743 (N_9743,N_7383,N_6239);
nand U9744 (N_9744,N_6399,N_7476);
and U9745 (N_9745,N_7116,N_6908);
or U9746 (N_9746,N_6391,N_7561);
and U9747 (N_9747,N_6208,N_7978);
xor U9748 (N_9748,N_6601,N_7449);
and U9749 (N_9749,N_7398,N_6380);
xor U9750 (N_9750,N_7599,N_7197);
xor U9751 (N_9751,N_6510,N_7402);
or U9752 (N_9752,N_6963,N_7169);
or U9753 (N_9753,N_6473,N_6039);
or U9754 (N_9754,N_6841,N_6826);
xnor U9755 (N_9755,N_6967,N_7497);
xnor U9756 (N_9756,N_7833,N_7396);
or U9757 (N_9757,N_7812,N_6927);
xor U9758 (N_9758,N_6912,N_7120);
xor U9759 (N_9759,N_6195,N_6965);
and U9760 (N_9760,N_6090,N_6254);
nor U9761 (N_9761,N_6246,N_7379);
nor U9762 (N_9762,N_7366,N_7449);
nor U9763 (N_9763,N_7405,N_7685);
and U9764 (N_9764,N_6009,N_6192);
xnor U9765 (N_9765,N_7582,N_7636);
and U9766 (N_9766,N_7863,N_6220);
or U9767 (N_9767,N_6607,N_7079);
xor U9768 (N_9768,N_6437,N_6366);
nand U9769 (N_9769,N_7599,N_6115);
or U9770 (N_9770,N_6751,N_7107);
and U9771 (N_9771,N_7937,N_7846);
or U9772 (N_9772,N_7280,N_7359);
and U9773 (N_9773,N_6284,N_7884);
or U9774 (N_9774,N_6194,N_6976);
or U9775 (N_9775,N_7688,N_6630);
and U9776 (N_9776,N_7753,N_7095);
or U9777 (N_9777,N_6556,N_7312);
and U9778 (N_9778,N_7062,N_7717);
xor U9779 (N_9779,N_6166,N_6409);
xor U9780 (N_9780,N_6890,N_6876);
xnor U9781 (N_9781,N_6521,N_6944);
xnor U9782 (N_9782,N_6431,N_7833);
and U9783 (N_9783,N_7249,N_6267);
nor U9784 (N_9784,N_7861,N_7248);
and U9785 (N_9785,N_6582,N_7553);
or U9786 (N_9786,N_7891,N_7291);
nor U9787 (N_9787,N_6906,N_6036);
nand U9788 (N_9788,N_6665,N_6690);
or U9789 (N_9789,N_6288,N_6357);
nor U9790 (N_9790,N_7782,N_6176);
xnor U9791 (N_9791,N_6964,N_6591);
and U9792 (N_9792,N_7708,N_7870);
nor U9793 (N_9793,N_6553,N_7729);
nor U9794 (N_9794,N_7189,N_6373);
and U9795 (N_9795,N_7429,N_7929);
xnor U9796 (N_9796,N_6195,N_6598);
xnor U9797 (N_9797,N_6985,N_6681);
nand U9798 (N_9798,N_7715,N_7196);
nor U9799 (N_9799,N_6313,N_6481);
xor U9800 (N_9800,N_7841,N_6160);
and U9801 (N_9801,N_7945,N_7439);
xor U9802 (N_9802,N_7220,N_7490);
nand U9803 (N_9803,N_6693,N_6396);
and U9804 (N_9804,N_7800,N_7302);
nand U9805 (N_9805,N_6018,N_6141);
or U9806 (N_9806,N_7487,N_7985);
nor U9807 (N_9807,N_6016,N_7943);
nor U9808 (N_9808,N_7206,N_7058);
nor U9809 (N_9809,N_7516,N_6833);
or U9810 (N_9810,N_7757,N_6417);
nand U9811 (N_9811,N_7311,N_7853);
and U9812 (N_9812,N_6132,N_6256);
nand U9813 (N_9813,N_7786,N_6022);
or U9814 (N_9814,N_7789,N_6014);
nand U9815 (N_9815,N_7440,N_6333);
nor U9816 (N_9816,N_7347,N_6810);
or U9817 (N_9817,N_6473,N_6612);
nand U9818 (N_9818,N_7536,N_7707);
nand U9819 (N_9819,N_6254,N_6329);
nor U9820 (N_9820,N_6502,N_6509);
or U9821 (N_9821,N_7284,N_7925);
or U9822 (N_9822,N_6542,N_6484);
nand U9823 (N_9823,N_7091,N_6818);
or U9824 (N_9824,N_6107,N_7748);
and U9825 (N_9825,N_6565,N_7500);
and U9826 (N_9826,N_7648,N_6504);
and U9827 (N_9827,N_6202,N_7250);
xor U9828 (N_9828,N_7743,N_7399);
and U9829 (N_9829,N_7704,N_7148);
and U9830 (N_9830,N_6027,N_6892);
nand U9831 (N_9831,N_7786,N_6794);
xnor U9832 (N_9832,N_7147,N_6285);
xnor U9833 (N_9833,N_6915,N_6363);
and U9834 (N_9834,N_6867,N_6651);
or U9835 (N_9835,N_7696,N_7380);
nand U9836 (N_9836,N_7663,N_6131);
or U9837 (N_9837,N_7357,N_7410);
xnor U9838 (N_9838,N_6182,N_7945);
or U9839 (N_9839,N_7649,N_7591);
or U9840 (N_9840,N_6914,N_7444);
and U9841 (N_9841,N_6122,N_6338);
or U9842 (N_9842,N_7753,N_6588);
nor U9843 (N_9843,N_7033,N_7596);
or U9844 (N_9844,N_7092,N_7048);
nand U9845 (N_9845,N_7764,N_6609);
xnor U9846 (N_9846,N_7409,N_7327);
or U9847 (N_9847,N_7220,N_6996);
and U9848 (N_9848,N_6055,N_7856);
nand U9849 (N_9849,N_7620,N_6559);
xnor U9850 (N_9850,N_6277,N_7684);
or U9851 (N_9851,N_7489,N_7014);
xor U9852 (N_9852,N_7484,N_6795);
xor U9853 (N_9853,N_6018,N_7299);
nor U9854 (N_9854,N_7683,N_7736);
nor U9855 (N_9855,N_6346,N_6353);
and U9856 (N_9856,N_7543,N_7787);
nand U9857 (N_9857,N_6411,N_7746);
xor U9858 (N_9858,N_7996,N_7838);
or U9859 (N_9859,N_6625,N_7788);
or U9860 (N_9860,N_6148,N_6653);
nand U9861 (N_9861,N_7647,N_7760);
nand U9862 (N_9862,N_7504,N_6041);
and U9863 (N_9863,N_6440,N_7870);
and U9864 (N_9864,N_7008,N_7739);
and U9865 (N_9865,N_7642,N_6753);
or U9866 (N_9866,N_7636,N_7674);
xor U9867 (N_9867,N_7090,N_7585);
nor U9868 (N_9868,N_7291,N_7921);
xnor U9869 (N_9869,N_6347,N_7999);
xor U9870 (N_9870,N_6518,N_6005);
or U9871 (N_9871,N_6002,N_6644);
nand U9872 (N_9872,N_7536,N_6091);
xor U9873 (N_9873,N_6422,N_7412);
xnor U9874 (N_9874,N_7342,N_7398);
and U9875 (N_9875,N_6043,N_6313);
nor U9876 (N_9876,N_6745,N_7016);
or U9877 (N_9877,N_7784,N_6384);
nand U9878 (N_9878,N_7376,N_7356);
nand U9879 (N_9879,N_6968,N_7307);
nand U9880 (N_9880,N_6156,N_6024);
xnor U9881 (N_9881,N_7755,N_6102);
xor U9882 (N_9882,N_7805,N_7617);
xnor U9883 (N_9883,N_6920,N_6260);
and U9884 (N_9884,N_6580,N_6230);
and U9885 (N_9885,N_7138,N_6654);
and U9886 (N_9886,N_7504,N_7596);
nand U9887 (N_9887,N_7045,N_7663);
nand U9888 (N_9888,N_7156,N_7696);
nor U9889 (N_9889,N_7401,N_6268);
xor U9890 (N_9890,N_7205,N_6323);
nand U9891 (N_9891,N_6309,N_6403);
and U9892 (N_9892,N_6847,N_7071);
and U9893 (N_9893,N_6549,N_6166);
xnor U9894 (N_9894,N_6116,N_6337);
nand U9895 (N_9895,N_7754,N_7407);
xor U9896 (N_9896,N_6206,N_6490);
and U9897 (N_9897,N_6528,N_7649);
xor U9898 (N_9898,N_6784,N_7899);
xnor U9899 (N_9899,N_7068,N_6790);
or U9900 (N_9900,N_7609,N_6315);
and U9901 (N_9901,N_6470,N_7709);
nor U9902 (N_9902,N_6657,N_6193);
nor U9903 (N_9903,N_7992,N_7197);
nor U9904 (N_9904,N_7425,N_6220);
or U9905 (N_9905,N_7607,N_6802);
xnor U9906 (N_9906,N_6128,N_7369);
nor U9907 (N_9907,N_6002,N_7905);
nand U9908 (N_9908,N_7685,N_7663);
xor U9909 (N_9909,N_6268,N_7398);
or U9910 (N_9910,N_7847,N_6308);
or U9911 (N_9911,N_6203,N_6255);
xnor U9912 (N_9912,N_7527,N_6603);
nand U9913 (N_9913,N_6886,N_6876);
nor U9914 (N_9914,N_7675,N_7251);
or U9915 (N_9915,N_7546,N_7471);
or U9916 (N_9916,N_6293,N_6650);
and U9917 (N_9917,N_6209,N_7993);
xnor U9918 (N_9918,N_6525,N_7928);
or U9919 (N_9919,N_7655,N_7934);
and U9920 (N_9920,N_6188,N_7726);
or U9921 (N_9921,N_7640,N_7944);
xor U9922 (N_9922,N_6082,N_6828);
nor U9923 (N_9923,N_6716,N_6378);
or U9924 (N_9924,N_7192,N_6340);
and U9925 (N_9925,N_7769,N_7499);
nor U9926 (N_9926,N_7505,N_6864);
xor U9927 (N_9927,N_6589,N_6356);
nand U9928 (N_9928,N_6259,N_7947);
nand U9929 (N_9929,N_7837,N_6110);
or U9930 (N_9930,N_7763,N_7623);
nor U9931 (N_9931,N_7315,N_6230);
nand U9932 (N_9932,N_6875,N_6001);
nor U9933 (N_9933,N_7774,N_7491);
nor U9934 (N_9934,N_7154,N_7505);
nor U9935 (N_9935,N_7682,N_7990);
or U9936 (N_9936,N_7914,N_6878);
xnor U9937 (N_9937,N_6575,N_7248);
xnor U9938 (N_9938,N_6010,N_6283);
xnor U9939 (N_9939,N_7275,N_7128);
nand U9940 (N_9940,N_7780,N_7851);
and U9941 (N_9941,N_7523,N_7649);
nor U9942 (N_9942,N_6268,N_7403);
and U9943 (N_9943,N_6314,N_6378);
xnor U9944 (N_9944,N_6704,N_6833);
or U9945 (N_9945,N_7931,N_7767);
xnor U9946 (N_9946,N_6728,N_6654);
and U9947 (N_9947,N_6132,N_6241);
and U9948 (N_9948,N_7514,N_6263);
nand U9949 (N_9949,N_6997,N_6315);
or U9950 (N_9950,N_7191,N_7946);
or U9951 (N_9951,N_7571,N_7989);
nand U9952 (N_9952,N_7481,N_7376);
or U9953 (N_9953,N_7977,N_6250);
nor U9954 (N_9954,N_6438,N_6564);
nand U9955 (N_9955,N_7641,N_6998);
nor U9956 (N_9956,N_7161,N_7910);
xnor U9957 (N_9957,N_6779,N_6008);
nor U9958 (N_9958,N_6505,N_6878);
nor U9959 (N_9959,N_7634,N_6641);
xor U9960 (N_9960,N_6383,N_6481);
nor U9961 (N_9961,N_6780,N_7275);
and U9962 (N_9962,N_7773,N_7994);
xor U9963 (N_9963,N_7661,N_6582);
xor U9964 (N_9964,N_6875,N_6650);
nor U9965 (N_9965,N_7175,N_7780);
xnor U9966 (N_9966,N_7154,N_7098);
or U9967 (N_9967,N_7635,N_7238);
xor U9968 (N_9968,N_6466,N_7917);
nand U9969 (N_9969,N_6406,N_7695);
nor U9970 (N_9970,N_7825,N_7437);
and U9971 (N_9971,N_6166,N_6851);
or U9972 (N_9972,N_7715,N_6490);
nand U9973 (N_9973,N_6308,N_7172);
and U9974 (N_9974,N_7884,N_7914);
nand U9975 (N_9975,N_6275,N_7469);
nor U9976 (N_9976,N_6010,N_7204);
nor U9977 (N_9977,N_6518,N_6880);
xor U9978 (N_9978,N_6309,N_7353);
and U9979 (N_9979,N_6676,N_6925);
nand U9980 (N_9980,N_6250,N_7457);
and U9981 (N_9981,N_7664,N_6896);
and U9982 (N_9982,N_7740,N_6974);
and U9983 (N_9983,N_7559,N_6168);
or U9984 (N_9984,N_6864,N_7104);
nand U9985 (N_9985,N_6602,N_6981);
and U9986 (N_9986,N_7676,N_7885);
nor U9987 (N_9987,N_6895,N_7771);
nor U9988 (N_9988,N_7002,N_6045);
nand U9989 (N_9989,N_7209,N_7191);
nor U9990 (N_9990,N_6535,N_6067);
and U9991 (N_9991,N_6715,N_7518);
nand U9992 (N_9992,N_7812,N_7018);
nand U9993 (N_9993,N_7301,N_6020);
xor U9994 (N_9994,N_6148,N_6547);
and U9995 (N_9995,N_7616,N_7181);
nand U9996 (N_9996,N_6912,N_6188);
xor U9997 (N_9997,N_6755,N_6776);
or U9998 (N_9998,N_7011,N_7376);
and U9999 (N_9999,N_6191,N_6046);
nor U10000 (N_10000,N_9227,N_9317);
nand U10001 (N_10001,N_9395,N_9532);
xnor U10002 (N_10002,N_8544,N_9255);
nand U10003 (N_10003,N_9727,N_8634);
nand U10004 (N_10004,N_8513,N_9959);
or U10005 (N_10005,N_8049,N_8398);
and U10006 (N_10006,N_8459,N_9072);
or U10007 (N_10007,N_8461,N_8880);
xor U10008 (N_10008,N_9294,N_9987);
xor U10009 (N_10009,N_8023,N_9304);
or U10010 (N_10010,N_8234,N_8556);
nand U10011 (N_10011,N_9437,N_9512);
xor U10012 (N_10012,N_8682,N_9180);
nand U10013 (N_10013,N_8550,N_8265);
or U10014 (N_10014,N_8577,N_9209);
nand U10015 (N_10015,N_8034,N_8699);
and U10016 (N_10016,N_9846,N_8570);
nor U10017 (N_10017,N_9129,N_9262);
or U10018 (N_10018,N_8965,N_9176);
nor U10019 (N_10019,N_8167,N_9174);
and U10020 (N_10020,N_9049,N_8002);
and U10021 (N_10021,N_8610,N_8165);
nand U10022 (N_10022,N_8404,N_9808);
nor U10023 (N_10023,N_9700,N_8527);
nor U10024 (N_10024,N_9245,N_8428);
nand U10025 (N_10025,N_9800,N_8869);
nand U10026 (N_10026,N_9004,N_9517);
nor U10027 (N_10027,N_9472,N_8684);
or U10028 (N_10028,N_8803,N_9545);
or U10029 (N_10029,N_8594,N_8901);
nand U10030 (N_10030,N_8957,N_8316);
nor U10031 (N_10031,N_9177,N_9113);
and U10032 (N_10032,N_8296,N_9336);
xnor U10033 (N_10033,N_9888,N_9300);
or U10034 (N_10034,N_8505,N_8017);
nor U10035 (N_10035,N_9046,N_9155);
nor U10036 (N_10036,N_9675,N_9875);
or U10037 (N_10037,N_9196,N_9951);
nand U10038 (N_10038,N_9983,N_9471);
nor U10039 (N_10039,N_8648,N_8623);
nand U10040 (N_10040,N_9058,N_8253);
or U10041 (N_10041,N_8319,N_8693);
xnor U10042 (N_10042,N_9642,N_9765);
nor U10043 (N_10043,N_8419,N_9082);
xnor U10044 (N_10044,N_8379,N_9956);
xnor U10045 (N_10045,N_9565,N_9443);
nand U10046 (N_10046,N_9486,N_9130);
nand U10047 (N_10047,N_9663,N_9370);
xor U10048 (N_10048,N_8827,N_8816);
nor U10049 (N_10049,N_9450,N_8559);
xnor U10050 (N_10050,N_8009,N_9065);
and U10051 (N_10051,N_9272,N_8406);
xor U10052 (N_10052,N_8552,N_8192);
or U10053 (N_10053,N_9056,N_9104);
or U10054 (N_10054,N_8276,N_9275);
nand U10055 (N_10055,N_8738,N_8408);
xnor U10056 (N_10056,N_8251,N_9407);
nor U10057 (N_10057,N_8670,N_8173);
and U10058 (N_10058,N_9077,N_9710);
nor U10059 (N_10059,N_8657,N_9935);
and U10060 (N_10060,N_8858,N_8347);
xnor U10061 (N_10061,N_8627,N_8717);
nor U10062 (N_10062,N_9198,N_9857);
nor U10063 (N_10063,N_9789,N_9842);
or U10064 (N_10064,N_8388,N_8365);
nand U10065 (N_10065,N_9869,N_8808);
xor U10066 (N_10066,N_8776,N_9687);
or U10067 (N_10067,N_8946,N_9362);
or U10068 (N_10068,N_9702,N_9210);
or U10069 (N_10069,N_8155,N_9464);
nand U10070 (N_10070,N_8035,N_8641);
nand U10071 (N_10071,N_8212,N_9341);
nor U10072 (N_10072,N_8895,N_8663);
or U10073 (N_10073,N_8958,N_8130);
nor U10074 (N_10074,N_8284,N_9240);
nor U10075 (N_10075,N_9896,N_9440);
xor U10076 (N_10076,N_8604,N_9215);
or U10077 (N_10077,N_8575,N_8087);
nand U10078 (N_10078,N_8063,N_8557);
and U10079 (N_10079,N_9225,N_8665);
nand U10080 (N_10080,N_9723,N_9587);
nand U10081 (N_10081,N_8525,N_8994);
xnor U10082 (N_10082,N_9513,N_9006);
nor U10083 (N_10083,N_9099,N_8332);
xnor U10084 (N_10084,N_9405,N_8982);
xnor U10085 (N_10085,N_8156,N_8233);
xnor U10086 (N_10086,N_8184,N_9848);
or U10087 (N_10087,N_9055,N_9193);
and U10088 (N_10088,N_9022,N_9994);
or U10089 (N_10089,N_9812,N_8083);
nor U10090 (N_10090,N_8990,N_9992);
and U10091 (N_10091,N_8888,N_9826);
and U10092 (N_10092,N_8567,N_9281);
xnor U10093 (N_10093,N_9829,N_9349);
xnor U10094 (N_10094,N_8462,N_9166);
and U10095 (N_10095,N_9673,N_8216);
and U10096 (N_10096,N_8908,N_9076);
or U10097 (N_10097,N_8686,N_9365);
xnor U10098 (N_10098,N_8135,N_8182);
and U10099 (N_10099,N_9684,N_9277);
and U10100 (N_10100,N_8169,N_9618);
nand U10101 (N_10101,N_9485,N_8681);
nor U10102 (N_10102,N_9912,N_8317);
nand U10103 (N_10103,N_8064,N_9679);
or U10104 (N_10104,N_8407,N_9915);
nand U10105 (N_10105,N_8042,N_9916);
and U10106 (N_10106,N_9861,N_9446);
nor U10107 (N_10107,N_8781,N_8578);
xnor U10108 (N_10108,N_9524,N_8057);
nor U10109 (N_10109,N_8259,N_8497);
nand U10110 (N_10110,N_9051,N_8336);
nor U10111 (N_10111,N_8915,N_9882);
nor U10112 (N_10112,N_9345,N_8724);
xor U10113 (N_10113,N_9045,N_9368);
nand U10114 (N_10114,N_8041,N_8626);
xnor U10115 (N_10115,N_9731,N_8645);
xnor U10116 (N_10116,N_9386,N_9630);
xnor U10117 (N_10117,N_8861,N_9698);
or U10118 (N_10118,N_8873,N_9161);
nor U10119 (N_10119,N_8044,N_9397);
nor U10120 (N_10120,N_9910,N_9554);
nand U10121 (N_10121,N_8831,N_9489);
xor U10122 (N_10122,N_8405,N_9263);
xnor U10123 (N_10123,N_8524,N_9760);
nor U10124 (N_10124,N_9584,N_8380);
xnor U10125 (N_10125,N_8555,N_8582);
and U10126 (N_10126,N_8005,N_9353);
and U10127 (N_10127,N_9518,N_8792);
and U10128 (N_10128,N_9794,N_9749);
or U10129 (N_10129,N_8980,N_8095);
and U10130 (N_10130,N_9550,N_8467);
or U10131 (N_10131,N_9572,N_8472);
xor U10132 (N_10132,N_8817,N_9886);
xor U10133 (N_10133,N_8385,N_8387);
or U10134 (N_10134,N_8774,N_9776);
and U10135 (N_10135,N_8585,N_8186);
or U10136 (N_10136,N_8521,N_9465);
and U10137 (N_10137,N_8073,N_8753);
or U10138 (N_10138,N_8903,N_9028);
nand U10139 (N_10139,N_8254,N_8833);
nand U10140 (N_10140,N_8938,N_8615);
and U10141 (N_10141,N_8490,N_8089);
or U10142 (N_10142,N_8386,N_8307);
nand U10143 (N_10143,N_9175,N_8722);
and U10144 (N_10144,N_9574,N_9746);
nand U10145 (N_10145,N_9964,N_9396);
nor U10146 (N_10146,N_8484,N_8327);
and U10147 (N_10147,N_9707,N_8881);
nor U10148 (N_10148,N_8787,N_8200);
nand U10149 (N_10149,N_8230,N_9639);
nor U10150 (N_10150,N_8756,N_8399);
xor U10151 (N_10151,N_8761,N_8890);
nand U10152 (N_10152,N_9629,N_8789);
nor U10153 (N_10153,N_8146,N_8763);
nand U10154 (N_10154,N_8417,N_9784);
or U10155 (N_10155,N_8059,N_9701);
or U10156 (N_10156,N_8003,N_9930);
or U10157 (N_10157,N_8204,N_8168);
nand U10158 (N_10158,N_9936,N_8710);
nand U10159 (N_10159,N_8126,N_8261);
nor U10160 (N_10160,N_9297,N_9555);
or U10161 (N_10161,N_8409,N_9751);
xnor U10162 (N_10162,N_8811,N_8099);
xnor U10163 (N_10163,N_9753,N_8275);
nand U10164 (N_10164,N_8109,N_9873);
nor U10165 (N_10165,N_8152,N_9863);
xnor U10166 (N_10166,N_8967,N_9266);
and U10167 (N_10167,N_9925,N_9868);
nor U10168 (N_10168,N_8164,N_8536);
nor U10169 (N_10169,N_9635,N_9773);
nand U10170 (N_10170,N_8326,N_8048);
or U10171 (N_10171,N_9285,N_8143);
xnor U10172 (N_10172,N_8759,N_9820);
and U10173 (N_10173,N_8197,N_8075);
nand U10174 (N_10174,N_8569,N_9391);
xor U10175 (N_10175,N_8036,N_8481);
or U10176 (N_10176,N_8766,N_8289);
nand U10177 (N_10177,N_9995,N_9590);
or U10178 (N_10178,N_8157,N_9414);
xnor U10179 (N_10179,N_9109,N_8802);
nor U10180 (N_10180,N_8826,N_8416);
and U10181 (N_10181,N_8286,N_9854);
or U10182 (N_10182,N_8836,N_8180);
xor U10183 (N_10183,N_9614,N_9913);
or U10184 (N_10184,N_8742,N_8032);
or U10185 (N_10185,N_8824,N_9503);
xor U10186 (N_10186,N_8560,N_9007);
and U10187 (N_10187,N_9020,N_9411);
or U10188 (N_10188,N_9534,N_9095);
and U10189 (N_10189,N_9354,N_9436);
xnor U10190 (N_10190,N_9268,N_9348);
or U10191 (N_10191,N_9378,N_9972);
xor U10192 (N_10192,N_9254,N_9595);
or U10193 (N_10193,N_8899,N_9408);
nand U10194 (N_10194,N_8225,N_9261);
nor U10195 (N_10195,N_8444,N_8972);
nand U10196 (N_10196,N_8315,N_9508);
or U10197 (N_10197,N_9952,N_8907);
xnor U10198 (N_10198,N_8176,N_8856);
or U10199 (N_10199,N_9783,N_9351);
nor U10200 (N_10200,N_9325,N_9217);
nor U10201 (N_10201,N_8008,N_9205);
nor U10202 (N_10202,N_8943,N_9732);
xor U10203 (N_10203,N_9769,N_8728);
or U10204 (N_10204,N_9228,N_8221);
nor U10205 (N_10205,N_8170,N_9091);
nor U10206 (N_10206,N_9954,N_9066);
and U10207 (N_10207,N_8345,N_8629);
or U10208 (N_10208,N_9074,N_9081);
and U10209 (N_10209,N_9119,N_8934);
nor U10210 (N_10210,N_9187,N_9745);
xor U10211 (N_10211,N_8374,N_8847);
or U10212 (N_10212,N_8716,N_9548);
nand U10213 (N_10213,N_9521,N_9226);
nand U10214 (N_10214,N_9706,N_9649);
nand U10215 (N_10215,N_8208,N_9990);
or U10216 (N_10216,N_8272,N_8866);
xor U10217 (N_10217,N_8605,N_9329);
and U10218 (N_10218,N_8391,N_8183);
nor U10219 (N_10219,N_9164,N_8624);
nor U10220 (N_10220,N_9087,N_9722);
and U10221 (N_10221,N_9571,N_8614);
xor U10222 (N_10222,N_8607,N_9797);
nand U10223 (N_10223,N_8479,N_9945);
xnor U10224 (N_10224,N_9360,N_8707);
nand U10225 (N_10225,N_8851,N_9017);
and U10226 (N_10226,N_9064,N_8447);
xor U10227 (N_10227,N_9905,N_9840);
and U10228 (N_10228,N_8203,N_8020);
nor U10229 (N_10229,N_8672,N_8715);
xnor U10230 (N_10230,N_8141,N_8726);
nand U10231 (N_10231,N_9016,N_8542);
or U10232 (N_10232,N_9439,N_9755);
nor U10233 (N_10233,N_9207,N_9515);
nor U10234 (N_10234,N_9836,N_9549);
and U10235 (N_10235,N_8050,N_9880);
and U10236 (N_10236,N_8733,N_8441);
nand U10237 (N_10237,N_8979,N_9984);
or U10238 (N_10238,N_9757,N_9214);
xnor U10239 (N_10239,N_9425,N_8342);
or U10240 (N_10240,N_8543,N_9451);
nor U10241 (N_10241,N_8477,N_9703);
or U10242 (N_10242,N_8778,N_9246);
xnor U10243 (N_10243,N_9509,N_9578);
nor U10244 (N_10244,N_8389,N_8288);
or U10245 (N_10245,N_9721,N_8346);
xnor U10246 (N_10246,N_9139,N_9522);
xnor U10247 (N_10247,N_9822,N_9202);
xor U10248 (N_10248,N_8928,N_8632);
xnor U10249 (N_10249,N_9303,N_8951);
and U10250 (N_10250,N_8683,N_8767);
nor U10251 (N_10251,N_9674,N_9319);
and U10252 (N_10252,N_8991,N_8538);
xor U10253 (N_10253,N_8078,N_9677);
nor U10254 (N_10254,N_9821,N_8440);
and U10255 (N_10255,N_8819,N_8503);
and U10256 (N_10256,N_8066,N_8223);
nand U10257 (N_10257,N_8674,N_9815);
and U10258 (N_10258,N_9010,N_9566);
xnor U10259 (N_10259,N_8476,N_9434);
nand U10260 (N_10260,N_8874,N_9320);
nand U10261 (N_10261,N_9942,N_8860);
nand U10262 (N_10262,N_9827,N_8217);
or U10263 (N_10263,N_8077,N_9352);
nor U10264 (N_10264,N_9709,N_8986);
nor U10265 (N_10265,N_8478,N_8936);
or U10266 (N_10266,N_8252,N_8944);
nor U10267 (N_10267,N_8457,N_8362);
and U10268 (N_10268,N_9188,N_8740);
and U10269 (N_10269,N_8518,N_9791);
or U10270 (N_10270,N_9200,N_9874);
nand U10271 (N_10271,N_8033,N_8746);
and U10272 (N_10272,N_8120,N_9393);
nor U10273 (N_10273,N_9357,N_9544);
nand U10274 (N_10274,N_9775,N_9400);
xor U10275 (N_10275,N_8611,N_9490);
or U10276 (N_10276,N_9605,N_9381);
nor U10277 (N_10277,N_8372,N_8381);
or U10278 (N_10278,N_9904,N_8533);
or U10279 (N_10279,N_8650,N_9787);
xnor U10280 (N_10280,N_8893,N_8311);
nand U10281 (N_10281,N_9009,N_8804);
nand U10282 (N_10282,N_8973,N_8865);
nor U10283 (N_10283,N_8985,N_8673);
and U10284 (N_10284,N_8660,N_9218);
xnor U10285 (N_10285,N_8675,N_9906);
or U10286 (N_10286,N_9718,N_8801);
nand U10287 (N_10287,N_8098,N_9314);
or U10288 (N_10288,N_9488,N_8134);
and U10289 (N_10289,N_8121,N_9617);
nor U10290 (N_10290,N_8705,N_8592);
or U10291 (N_10291,N_9585,N_8268);
nor U10292 (N_10292,N_8909,N_9053);
xnor U10293 (N_10293,N_9292,N_8815);
nand U10294 (N_10294,N_8963,N_9308);
or U10295 (N_10295,N_9948,N_8661);
nor U10296 (N_10296,N_8247,N_8771);
nand U10297 (N_10297,N_8514,N_8413);
nand U10298 (N_10298,N_9851,N_9478);
and U10299 (N_10299,N_9390,N_9531);
or U10300 (N_10300,N_8599,N_8045);
xnor U10301 (N_10301,N_9785,N_8402);
and U10302 (N_10302,N_8834,N_8721);
nand U10303 (N_10303,N_9422,N_8085);
xnor U10304 (N_10304,N_9733,N_9852);
nand U10305 (N_10305,N_9219,N_9047);
xor U10306 (N_10306,N_9713,N_9170);
xnor U10307 (N_10307,N_9415,N_9057);
or U10308 (N_10308,N_9132,N_8297);
or U10309 (N_10309,N_8016,N_9979);
nor U10310 (N_10310,N_8264,N_8517);
xnor U10311 (N_10311,N_8698,N_8941);
nand U10312 (N_10312,N_9855,N_9213);
nor U10313 (N_10313,N_8090,N_9309);
and U10314 (N_10314,N_8433,N_9274);
or U10315 (N_10315,N_9146,N_9641);
xnor U10316 (N_10316,N_9593,N_8425);
or U10317 (N_10317,N_8117,N_8174);
nor U10318 (N_10318,N_8487,N_9279);
nand U10319 (N_10319,N_8222,N_9890);
or U10320 (N_10320,N_8158,N_9944);
xor U10321 (N_10321,N_9011,N_9652);
nand U10322 (N_10322,N_8148,N_9473);
or U10323 (N_10323,N_8432,N_8199);
nand U10324 (N_10324,N_9982,N_8287);
and U10325 (N_10325,N_9969,N_8012);
or U10326 (N_10326,N_8747,N_9729);
or U10327 (N_10327,N_8153,N_8981);
nand U10328 (N_10328,N_9030,N_8921);
nand U10329 (N_10329,N_8734,N_8482);
nand U10330 (N_10330,N_8652,N_9256);
nor U10331 (N_10331,N_9416,N_8248);
nand U10332 (N_10332,N_8812,N_9817);
nor U10333 (N_10333,N_8474,N_8056);
nor U10334 (N_10334,N_9691,N_8102);
or U10335 (N_10335,N_8519,N_8953);
or U10336 (N_10336,N_9567,N_9239);
xor U10337 (N_10337,N_9569,N_9887);
xnor U10338 (N_10338,N_9301,N_9250);
and U10339 (N_10339,N_8788,N_8685);
nor U10340 (N_10340,N_9922,N_8328);
xnor U10341 (N_10341,N_9625,N_9101);
and U10342 (N_10342,N_9530,N_8279);
nor U10343 (N_10343,N_9697,N_8468);
xor U10344 (N_10344,N_9159,N_8886);
xnor U10345 (N_10345,N_9670,N_9844);
xnor U10346 (N_10346,N_9603,N_9212);
nand U10347 (N_10347,N_8917,N_9803);
xnor U10348 (N_10348,N_9665,N_9404);
xnor U10349 (N_10349,N_9133,N_8838);
nor U10350 (N_10350,N_8736,N_9655);
nand U10351 (N_10351,N_9172,N_8922);
nand U10352 (N_10352,N_9909,N_8298);
nor U10353 (N_10353,N_8832,N_8855);
nand U10354 (N_10354,N_8828,N_9334);
or U10355 (N_10355,N_9445,N_9034);
or U10356 (N_10356,N_8446,N_8600);
or U10357 (N_10357,N_9893,N_9481);
xnor U10358 (N_10358,N_9282,N_8281);
or U10359 (N_10359,N_8696,N_9197);
and U10360 (N_10360,N_9038,N_9553);
and U10361 (N_10361,N_8343,N_8976);
nor U10362 (N_10362,N_9654,N_9778);
and U10363 (N_10363,N_9908,N_9993);
nor U10364 (N_10364,N_8800,N_8000);
xnor U10365 (N_10365,N_9100,N_9249);
nand U10366 (N_10366,N_9154,N_8794);
nor U10367 (N_10367,N_8541,N_8160);
and U10368 (N_10368,N_8266,N_9127);
and U10369 (N_10369,N_8280,N_8823);
nand U10370 (N_10370,N_8350,N_9376);
nand U10371 (N_10371,N_8798,N_9612);
or U10372 (N_10372,N_9955,N_9189);
or U10373 (N_10373,N_8231,N_9331);
and U10374 (N_10374,N_8451,N_9001);
xor U10375 (N_10375,N_9824,N_8238);
nand U10376 (N_10376,N_9728,N_9623);
nor U10377 (N_10377,N_8480,N_8612);
or U10378 (N_10378,N_8574,N_9105);
nor U10379 (N_10379,N_8608,N_9454);
nor U10380 (N_10380,N_8105,N_8878);
or U10381 (N_10381,N_8974,N_8240);
xor U10382 (N_10382,N_8654,N_9788);
and U10383 (N_10383,N_8357,N_9809);
nor U10384 (N_10384,N_9298,N_9157);
nand U10385 (N_10385,N_9616,N_9343);
nor U10386 (N_10386,N_8344,N_8129);
nor U10387 (N_10387,N_9377,N_8891);
nand U10388 (N_10388,N_9192,N_9040);
or U10389 (N_10389,N_8978,N_9421);
nand U10390 (N_10390,N_9997,N_8845);
nor U10391 (N_10391,N_9431,N_9068);
nor U10392 (N_10392,N_8712,N_9651);
and U10393 (N_10393,N_9734,N_9234);
nand U10394 (N_10394,N_8260,N_8697);
nand U10395 (N_10395,N_8587,N_9685);
or U10396 (N_10396,N_8473,N_8151);
nand U10397 (N_10397,N_8637,N_8303);
and U10398 (N_10398,N_8027,N_8580);
or U10399 (N_10399,N_9793,N_9790);
and U10400 (N_10400,N_9845,N_9284);
xnor U10401 (N_10401,N_9506,N_8583);
xor U10402 (N_10402,N_9183,N_8925);
and U10403 (N_10403,N_8030,N_8784);
and U10404 (N_10404,N_9000,N_8571);
nand U10405 (N_10405,N_9712,N_9537);
nor U10406 (N_10406,N_9427,N_8383);
nor U10407 (N_10407,N_8520,N_8884);
nor U10408 (N_10408,N_8492,N_9122);
or U10409 (N_10409,N_8731,N_8422);
xor U10410 (N_10410,N_8494,N_8862);
or U10411 (N_10411,N_8299,N_9278);
and U10412 (N_10412,N_9097,N_9088);
nor U10413 (N_10413,N_8366,N_8876);
nand U10414 (N_10414,N_8945,N_9950);
or U10415 (N_10415,N_9579,N_8360);
nand U10416 (N_10416,N_9135,N_9355);
or U10417 (N_10417,N_8708,N_8015);
or U10418 (N_10418,N_8772,N_8456);
xnor U10419 (N_10419,N_9551,N_9560);
or U10420 (N_10420,N_9676,N_9143);
or U10421 (N_10421,N_8331,N_9867);
nor U10422 (N_10422,N_9694,N_8115);
xor U10423 (N_10423,N_9632,N_8218);
and U10424 (N_10424,N_9070,N_8159);
nand U10425 (N_10425,N_8338,N_9025);
and U10426 (N_10426,N_9069,N_9762);
or U10427 (N_10427,N_9795,N_9973);
nand U10428 (N_10428,N_8037,N_9932);
nand U10429 (N_10429,N_8655,N_9504);
nor U10430 (N_10430,N_9469,N_9123);
and U10431 (N_10431,N_8664,N_8822);
nand U10432 (N_10432,N_9126,N_9374);
xor U10433 (N_10433,N_8438,N_9704);
xor U10434 (N_10434,N_9418,N_9475);
and U10435 (N_10435,N_9409,N_8370);
xnor U10436 (N_10436,N_9160,N_8700);
xnor U10437 (N_10437,N_9849,N_8224);
nand U10438 (N_10438,N_9724,N_9441);
nor U10439 (N_10439,N_8061,N_9716);
nand U10440 (N_10440,N_9291,N_8396);
xor U10441 (N_10441,N_8595,N_8760);
nor U10442 (N_10442,N_9985,N_8894);
and U10443 (N_10443,N_8445,N_9224);
and U10444 (N_10444,N_8162,N_9540);
or U10445 (N_10445,N_9211,N_8701);
and U10446 (N_10446,N_8131,N_8962);
xor U10447 (N_10447,N_8410,N_9967);
and U10448 (N_10448,N_9535,N_8961);
or U10449 (N_10449,N_9356,N_9860);
nor U10450 (N_10450,N_9247,N_9599);
nor U10451 (N_10451,N_9696,N_8508);
or U10452 (N_10452,N_8026,N_8201);
and U10453 (N_10453,N_9466,N_8163);
nor U10454 (N_10454,N_8219,N_9897);
xor U10455 (N_10455,N_8852,N_9523);
xnor U10456 (N_10456,N_8426,N_9991);
xnor U10457 (N_10457,N_9067,N_9657);
nand U10458 (N_10458,N_9961,N_9027);
xor U10459 (N_10459,N_9774,N_8080);
xnor U10460 (N_10460,N_9310,N_8584);
nor U10461 (N_10461,N_8730,N_8597);
nor U10462 (N_10462,N_9433,N_8321);
xor U10463 (N_10463,N_9621,N_9739);
or U10464 (N_10464,N_9387,N_8547);
or U10465 (N_10465,N_9686,N_9152);
and U10466 (N_10466,N_9919,N_9546);
nor U10467 (N_10467,N_9777,N_8935);
xnor U10468 (N_10468,N_9204,N_9692);
or U10469 (N_10469,N_9717,N_9257);
or U10470 (N_10470,N_9244,N_9735);
nor U10471 (N_10471,N_9662,N_9726);
and U10472 (N_10472,N_9496,N_8304);
xnor U10473 (N_10473,N_9048,N_9558);
nor U10474 (N_10474,N_8313,N_8640);
nor U10475 (N_10475,N_8437,N_8609);
or U10476 (N_10476,N_8244,N_9165);
or U10477 (N_10477,N_8821,N_9720);
nor U10478 (N_10478,N_9302,N_9561);
nand U10479 (N_10479,N_9792,N_8485);
nor U10480 (N_10480,N_8081,N_8564);
nor U10481 (N_10481,N_9804,N_9666);
and U10482 (N_10482,N_9032,N_8933);
xor U10483 (N_10483,N_9669,N_9287);
or U10484 (N_10484,N_9940,N_9738);
nor U10485 (N_10485,N_9359,N_8807);
and U10486 (N_10486,N_8455,N_8308);
or U10487 (N_10487,N_8662,N_9493);
xnor U10488 (N_10488,N_9516,N_8052);
nand U10489 (N_10489,N_8070,N_9158);
nor U10490 (N_10490,N_9410,N_9491);
and U10491 (N_10491,N_9121,N_8142);
nand U10492 (N_10492,N_8322,N_8601);
nand U10493 (N_10493,N_8237,N_9598);
nor U10494 (N_10494,N_9190,N_8507);
xnor U10495 (N_10495,N_8711,N_9380);
nand U10496 (N_10496,N_9767,N_9645);
and U10497 (N_10497,N_9367,N_8805);
nor U10498 (N_10498,N_9575,N_9273);
and U10499 (N_10499,N_9231,N_8889);
nand U10500 (N_10500,N_9646,N_9019);
xor U10501 (N_10501,N_9941,N_8735);
nand U10502 (N_10502,N_8628,N_8046);
or U10503 (N_10503,N_9145,N_9452);
nor U10504 (N_10504,N_8116,N_8523);
or U10505 (N_10505,N_8373,N_8750);
nor U10506 (N_10506,N_9693,N_9970);
xor U10507 (N_10507,N_9858,N_8795);
nor U10508 (N_10508,N_9276,N_9801);
nand U10509 (N_10509,N_9962,N_9741);
or U10510 (N_10510,N_9021,N_9293);
and U10511 (N_10511,N_9759,N_9748);
nand U10512 (N_10512,N_8329,N_9251);
xnor U10513 (N_10513,N_8335,N_8988);
nor U10514 (N_10514,N_9609,N_9447);
or U10515 (N_10515,N_8679,N_9080);
xnor U10516 (N_10516,N_8214,N_9606);
or U10517 (N_10517,N_9457,N_8242);
nor U10518 (N_10518,N_8576,N_8436);
or U10519 (N_10519,N_9570,N_9862);
xnor U10520 (N_10520,N_9502,N_8097);
nand U10521 (N_10521,N_8897,N_9182);
and U10522 (N_10522,N_9823,N_8561);
xnor U10523 (N_10523,N_8442,N_9881);
nand U10524 (N_10524,N_9108,N_8414);
nor U10525 (N_10525,N_9667,N_9853);
or U10526 (N_10526,N_9086,N_8205);
or U10527 (N_10527,N_8213,N_9449);
or U10528 (N_10528,N_8086,N_9914);
or U10529 (N_10529,N_8590,N_8659);
or U10530 (N_10530,N_9333,N_9151);
and U10531 (N_10531,N_9819,N_9772);
nor U10532 (N_10532,N_8745,N_8400);
nand U10533 (N_10533,N_8937,N_8695);
nand U10534 (N_10534,N_9843,N_8188);
or U10535 (N_10535,N_8429,N_8314);
or U10536 (N_10536,N_9798,N_8902);
nand U10537 (N_10537,N_8359,N_8718);
nor U10538 (N_10538,N_9664,N_9085);
and U10539 (N_10539,N_8123,N_9871);
xnor U10540 (N_10540,N_9974,N_9744);
or U10541 (N_10541,N_8616,N_8051);
or U10542 (N_10542,N_8094,N_9607);
or U10543 (N_10543,N_9658,N_9953);
xnor U10544 (N_10544,N_9090,N_8687);
nor U10545 (N_10545,N_8295,N_8024);
nor U10546 (N_10546,N_9063,N_9986);
xnor U10547 (N_10547,N_8274,N_8995);
nor U10548 (N_10548,N_8668,N_8535);
or U10549 (N_10549,N_8598,N_8806);
and U10550 (N_10550,N_8458,N_8647);
nor U10551 (N_10551,N_8107,N_8103);
xor U10552 (N_10552,N_9814,N_9557);
nor U10553 (N_10553,N_9156,N_8954);
xnor U10554 (N_10554,N_8565,N_9168);
or U10555 (N_10555,N_9660,N_9459);
nand U10556 (N_10556,N_9668,N_9901);
or U10557 (N_10557,N_9125,N_8150);
nand U10558 (N_10558,N_9847,N_9315);
xnor U10559 (N_10559,N_8491,N_9903);
nor U10560 (N_10560,N_8434,N_8431);
or U10561 (N_10561,N_8622,N_9740);
nand U10562 (N_10562,N_9178,N_8189);
nand U10563 (N_10563,N_9999,N_9003);
nor U10564 (N_10564,N_9036,N_9562);
or U10565 (N_10565,N_9615,N_9511);
nor U10566 (N_10566,N_8149,N_9628);
nor U10567 (N_10567,N_8942,N_8125);
nand U10568 (N_10568,N_9895,N_9911);
xor U10569 (N_10569,N_9044,N_9269);
xor U10570 (N_10570,N_8777,N_8950);
and U10571 (N_10571,N_8101,N_8093);
nor U10572 (N_10572,N_9347,N_9556);
or U10573 (N_10573,N_9520,N_9059);
xor U10574 (N_10574,N_9384,N_8703);
or U10575 (N_10575,N_8337,N_8154);
and U10576 (N_10576,N_8486,N_9949);
xnor U10577 (N_10577,N_9201,N_8190);
nor U10578 (N_10578,N_9206,N_9461);
or U10579 (N_10579,N_9098,N_8285);
or U10580 (N_10580,N_8356,N_8723);
xnor U10581 (N_10581,N_9631,N_8144);
xnor U10582 (N_10582,N_9456,N_8110);
xor U10583 (N_10583,N_9763,N_8423);
xor U10584 (N_10584,N_9866,N_8923);
or U10585 (N_10585,N_8341,N_9839);
and U10586 (N_10586,N_8349,N_9600);
and U10587 (N_10587,N_9543,N_9467);
or U10588 (N_10588,N_8235,N_9476);
or U10589 (N_10589,N_8074,N_9375);
or U10590 (N_10590,N_9026,N_9596);
nor U10591 (N_10591,N_9417,N_8330);
and U10592 (N_10592,N_8725,N_8546);
and U10593 (N_10593,N_9379,N_8940);
or U10594 (N_10594,N_8868,N_8864);
and U10595 (N_10595,N_9564,N_9114);
or U10596 (N_10596,N_9462,N_9243);
or U10597 (N_10597,N_8835,N_9388);
or U10598 (N_10598,N_8470,N_9781);
nand U10599 (N_10599,N_9805,N_8108);
nand U10600 (N_10600,N_8351,N_8566);
nand U10601 (N_10601,N_8185,N_8239);
and U10602 (N_10602,N_8226,N_8796);
xnor U10603 (N_10603,N_8452,N_8512);
nor U10604 (N_10604,N_9761,N_9818);
and U10605 (N_10605,N_8006,N_8172);
xnor U10606 (N_10606,N_9877,N_8989);
xnor U10607 (N_10607,N_8646,N_9771);
nor U10608 (N_10608,N_8970,N_8920);
and U10609 (N_10609,N_8857,N_9093);
and U10610 (N_10610,N_9002,N_8175);
and U10611 (N_10611,N_8011,N_9296);
and U10612 (N_10612,N_8975,N_8568);
nand U10613 (N_10613,N_8502,N_8987);
and U10614 (N_10614,N_9383,N_9307);
or U10615 (N_10615,N_9638,N_8053);
nand U10616 (N_10616,N_8291,N_9611);
and U10617 (N_10617,N_9444,N_8691);
or U10618 (N_10618,N_8054,N_9902);
or U10619 (N_10619,N_8114,N_8515);
xnor U10620 (N_10620,N_8939,N_9719);
or U10621 (N_10621,N_8229,N_9957);
xnor U10622 (N_10622,N_8912,N_9078);
and U10623 (N_10623,N_8591,N_8136);
xor U10624 (N_10624,N_8191,N_9998);
and U10625 (N_10625,N_8018,N_8392);
or U10626 (N_10626,N_8992,N_8773);
xnor U10627 (N_10627,N_9601,N_9094);
or U10628 (N_10628,N_9743,N_8882);
or U10629 (N_10629,N_8060,N_8088);
nor U10630 (N_10630,N_9656,N_8139);
xnor U10631 (N_10631,N_9042,N_8306);
xnor U10632 (N_10632,N_8900,N_8178);
nor U10633 (N_10633,N_9037,N_9392);
xnor U10634 (N_10634,N_9938,N_9659);
nor U10635 (N_10635,N_8118,N_8764);
nor U10636 (N_10636,N_8949,N_8522);
or U10637 (N_10637,N_8464,N_9112);
and U10638 (N_10638,N_8501,N_8215);
xor U10639 (N_10639,N_8892,N_9920);
xor U10640 (N_10640,N_9463,N_9876);
nand U10641 (N_10641,N_8765,N_9423);
nor U10642 (N_10642,N_8510,N_8013);
nand U10643 (N_10643,N_9260,N_9171);
nand U10644 (N_10644,N_9385,N_8529);
or U10645 (N_10645,N_8531,N_8952);
xnor U10646 (N_10646,N_8739,N_9364);
or U10647 (N_10647,N_8076,N_8460);
or U10648 (N_10648,N_9084,N_9526);
nand U10649 (N_10649,N_8166,N_9191);
nor U10650 (N_10650,N_8082,N_9937);
and U10651 (N_10651,N_8509,N_8530);
and U10652 (N_10652,N_8273,N_8558);
or U10653 (N_10653,N_9043,N_9754);
or U10654 (N_10654,N_9661,N_9012);
xor U10655 (N_10655,N_9831,N_8755);
nor U10656 (N_10656,N_9029,N_9313);
or U10657 (N_10657,N_8825,N_8688);
and U10658 (N_10658,N_8004,N_8068);
and U10659 (N_10659,N_9806,N_8228);
xor U10660 (N_10660,N_8551,N_9889);
nand U10661 (N_10661,N_9162,N_8334);
nor U10662 (N_10662,N_8333,N_9323);
xor U10663 (N_10663,N_9927,N_9406);
nor U10664 (N_10664,N_9453,N_9235);
nand U10665 (N_10665,N_9148,N_9619);
nor U10666 (N_10666,N_9637,N_9163);
nand U10667 (N_10667,N_8927,N_9715);
and U10668 (N_10668,N_9116,N_8929);
xor U10669 (N_10669,N_8282,N_9730);
nor U10670 (N_10670,N_9033,N_8029);
and U10671 (N_10671,N_9883,N_9528);
and U10672 (N_10672,N_8256,N_9136);
or U10673 (N_10673,N_9435,N_8667);
or U10674 (N_10674,N_8883,N_9372);
nand U10675 (N_10675,N_9539,N_8368);
nand U10676 (N_10676,N_9832,N_8642);
nand U10677 (N_10677,N_8187,N_8727);
nor U10678 (N_10678,N_9144,N_8177);
xnor U10679 (N_10679,N_8534,N_9120);
nand U10680 (N_10680,N_8206,N_8849);
or U10681 (N_10681,N_9725,N_9203);
nand U10682 (N_10682,N_8926,N_9173);
xor U10683 (N_10683,N_8999,N_8161);
or U10684 (N_10684,N_8966,N_8814);
xor U10685 (N_10685,N_9358,N_9926);
xor U10686 (N_10686,N_8618,N_8636);
nor U10687 (N_10687,N_8780,N_8403);
and U10688 (N_10688,N_8500,N_9604);
or U10689 (N_10689,N_9229,N_8209);
nor U10690 (N_10690,N_9194,N_8475);
nand U10691 (N_10691,N_9758,N_9402);
nand U10692 (N_10692,N_8047,N_8853);
nand U10693 (N_10693,N_8964,N_8848);
or U10694 (N_10694,N_9884,N_9865);
xnor U10695 (N_10695,N_8713,N_9420);
and U10696 (N_10696,N_8867,N_8841);
nor U10697 (N_10697,N_9939,N_8573);
xor U10698 (N_10698,N_8785,N_9633);
and U10699 (N_10699,N_8799,N_9432);
or U10700 (N_10700,N_9828,N_9216);
and U10701 (N_10701,N_8309,N_9138);
xor U10702 (N_10702,N_8412,N_9005);
and U10703 (N_10703,N_8621,N_9779);
nor U10704 (N_10704,N_8448,N_8863);
nor U10705 (N_10705,N_8352,N_9737);
or U10706 (N_10706,N_9330,N_9394);
nand U10707 (N_10707,N_9267,N_8656);
or U10708 (N_10708,N_9613,N_8471);
and U10709 (N_10709,N_8496,N_9265);
nor U10710 (N_10710,N_8689,N_8232);
nand U10711 (N_10711,N_8732,N_8589);
nand U10712 (N_10712,N_8540,N_8258);
or U10713 (N_10713,N_9573,N_8752);
xnor U10714 (N_10714,N_9366,N_9960);
nor U10715 (N_10715,N_8133,N_8055);
nand U10716 (N_10716,N_9978,N_8719);
or U10717 (N_10717,N_9591,N_8751);
or U10718 (N_10718,N_8720,N_9841);
and U10719 (N_10719,N_8124,N_9023);
or U10720 (N_10720,N_8666,N_9766);
or U10721 (N_10721,N_8324,N_9460);
nand U10722 (N_10722,N_9241,N_8353);
xnor U10723 (N_10723,N_9141,N_9859);
and U10724 (N_10724,N_8430,N_9280);
nand U10725 (N_10725,N_8022,N_9186);
xnor U10726 (N_10726,N_8007,N_9653);
nor U10727 (N_10727,N_9167,N_9369);
or U10728 (N_10728,N_8021,N_8931);
xor U10729 (N_10729,N_9499,N_9311);
and U10730 (N_10730,N_8579,N_9928);
nor U10731 (N_10731,N_8246,N_8677);
or U10732 (N_10732,N_9533,N_8602);
and U10733 (N_10733,N_8181,N_9339);
xor U10734 (N_10734,N_8278,N_9864);
and U10735 (N_10735,N_9492,N_8692);
or U10736 (N_10736,N_9102,N_9946);
nor U10737 (N_10737,N_9327,N_8411);
or U10738 (N_10738,N_9131,N_9626);
nand U10739 (N_10739,N_9468,N_9594);
nand U10740 (N_10740,N_8709,N_8643);
xnor U10741 (N_10741,N_9419,N_9885);
nor U10742 (N_10742,N_8019,N_8270);
nand U10743 (N_10743,N_9054,N_9110);
or U10744 (N_10744,N_9350,N_8786);
or U10745 (N_10745,N_8528,N_8549);
and U10746 (N_10746,N_9830,N_8450);
xnor U10747 (N_10747,N_9872,N_9577);
and U10748 (N_10748,N_8348,N_9305);
and U10749 (N_10749,N_8010,N_9096);
nand U10750 (N_10750,N_9248,N_9923);
xnor U10751 (N_10751,N_8318,N_9742);
nand U10752 (N_10752,N_8914,N_8993);
nand U10753 (N_10753,N_8421,N_9340);
nand U10754 (N_10754,N_8554,N_8932);
or U10755 (N_10755,N_8871,N_8948);
nor U10756 (N_10756,N_8390,N_9971);
and U10757 (N_10757,N_8395,N_8495);
or U10758 (N_10758,N_8638,N_8202);
xnor U10759 (N_10759,N_9035,N_8769);
nor U10760 (N_10760,N_8748,N_8122);
xor U10761 (N_10761,N_8910,N_8111);
nor U10762 (N_10762,N_9966,N_9232);
and U10763 (N_10763,N_9083,N_9286);
nor U10764 (N_10764,N_9650,N_9181);
or U10765 (N_10765,N_8147,N_8250);
and U10766 (N_10766,N_9780,N_9290);
nand U10767 (N_10767,N_8096,N_8269);
nand U10768 (N_10768,N_9681,N_9062);
xnor U10769 (N_10769,N_9586,N_8998);
xor U10770 (N_10770,N_8112,N_8617);
nand U10771 (N_10771,N_9222,N_9321);
nand U10772 (N_10772,N_9796,N_9115);
or U10773 (N_10773,N_8757,N_9929);
or U10774 (N_10774,N_8690,N_8371);
and U10775 (N_10775,N_8499,N_9835);
and U10776 (N_10776,N_9947,N_9238);
or U10777 (N_10777,N_9147,N_9917);
and U10778 (N_10778,N_8393,N_8511);
nor U10779 (N_10779,N_8820,N_8516);
nand U10780 (N_10780,N_8581,N_9501);
nand U10781 (N_10781,N_9223,N_8984);
xor U10782 (N_10782,N_9878,N_8758);
nand U10783 (N_10783,N_9306,N_9965);
or U10784 (N_10784,N_9592,N_8493);
and U10785 (N_10785,N_8960,N_8671);
and U10786 (N_10786,N_9918,N_9879);
nor U10787 (N_10787,N_9438,N_9071);
nand U10788 (N_10788,N_8603,N_9061);
nor U10789 (N_10789,N_8294,N_8846);
nand U10790 (N_10790,N_9117,N_8069);
nand U10791 (N_10791,N_8924,N_8572);
or U10792 (N_10792,N_8791,N_8427);
nor U10793 (N_10793,N_8394,N_8263);
xnor U10794 (N_10794,N_9620,N_8651);
nor U10795 (N_10795,N_8211,N_8454);
xor U10796 (N_10796,N_9199,N_9474);
nor U10797 (N_10797,N_9898,N_9338);
nand U10798 (N_10798,N_8301,N_8714);
or U10799 (N_10799,N_9140,N_9542);
nor U10800 (N_10800,N_8539,N_9015);
and U10801 (N_10801,N_8469,N_8593);
and U10802 (N_10802,N_8844,N_8596);
xor U10803 (N_10803,N_9756,N_9221);
or U10804 (N_10804,N_9089,N_9559);
nor U10805 (N_10805,N_9931,N_9149);
nand U10806 (N_10806,N_9708,N_9429);
and U10807 (N_10807,N_9128,N_8100);
nand U10808 (N_10808,N_8977,N_8062);
or U10809 (N_10809,N_8694,N_8678);
nand U10810 (N_10810,N_8375,N_9690);
nand U10811 (N_10811,N_8439,N_9563);
nand U10812 (N_10812,N_9363,N_8898);
or U10813 (N_10813,N_9714,N_8905);
nor U10814 (N_10814,N_9484,N_8323);
nor U10815 (N_10815,N_9608,N_9870);
or U10816 (N_10816,N_8255,N_8067);
nor U10817 (N_10817,N_9318,N_9024);
nand U10818 (N_10818,N_8267,N_9252);
and U10819 (N_10819,N_8630,N_8290);
xor U10820 (N_10820,N_9283,N_8532);
and U10821 (N_10821,N_8906,N_8783);
nand U10822 (N_10822,N_9008,N_8236);
and U10823 (N_10823,N_8782,N_8872);
nor U10824 (N_10824,N_9344,N_8810);
nand U10825 (N_10825,N_9271,N_8877);
nand U10826 (N_10826,N_8930,N_9118);
nand U10827 (N_10827,N_8850,N_8283);
nor U10828 (N_10828,N_9894,N_8220);
nand U10829 (N_10829,N_9671,N_8367);
or U10830 (N_10830,N_9736,N_8377);
xnor U10831 (N_10831,N_9541,N_8384);
xnor U10832 (N_10832,N_9695,N_8382);
nor U10833 (N_10833,N_8588,N_9934);
xnor U10834 (N_10834,N_8424,N_9495);
or U10835 (N_10835,N_9482,N_9589);
xnor U10836 (N_10836,N_9134,N_9031);
or U10837 (N_10837,N_9426,N_9892);
or U10838 (N_10838,N_9018,N_9634);
nand U10839 (N_10839,N_8132,N_9153);
and U10840 (N_10840,N_8744,N_8839);
nand U10841 (N_10841,N_8702,N_8737);
or U10842 (N_10842,N_8065,N_9813);
xnor U10843 (N_10843,N_9424,N_9647);
nand U10844 (N_10844,N_9052,N_8031);
or U10845 (N_10845,N_8194,N_9747);
nor U10846 (N_10846,N_9361,N_9602);
nor U10847 (N_10847,N_9624,N_8001);
and U10848 (N_10848,N_9519,N_9289);
nor U10849 (N_10849,N_9013,N_9636);
xor U10850 (N_10850,N_8210,N_8829);
or U10851 (N_10851,N_9833,N_9258);
nor U10852 (N_10852,N_8562,N_9299);
or U10853 (N_10853,N_8378,N_8840);
nor U10854 (N_10854,N_9907,N_8706);
nor U10855 (N_10855,N_9092,N_8271);
xor U10856 (N_10856,N_8241,N_9498);
and U10857 (N_10857,N_9312,N_8918);
and U10858 (N_10858,N_8644,N_9041);
xor U10859 (N_10859,N_9403,N_9678);
or U10860 (N_10860,N_9111,N_9799);
nor U10861 (N_10861,N_9943,N_9470);
xnor U10862 (N_10862,N_8453,N_9382);
nand U10863 (N_10863,N_8489,N_9371);
xor U10864 (N_10864,N_9184,N_8790);
xnor U10865 (N_10865,N_9583,N_9672);
or U10866 (N_10866,N_8537,N_9597);
or U10867 (N_10867,N_8179,N_8361);
or U10868 (N_10868,N_9220,N_8959);
nor U10869 (N_10869,N_9014,N_8916);
nor U10870 (N_10870,N_9680,N_9689);
nor U10871 (N_10871,N_8207,N_9398);
xnor U10872 (N_10872,N_8354,N_8859);
or U10873 (N_10873,N_8729,N_8553);
and U10874 (N_10874,N_9924,N_9428);
xor U10875 (N_10875,N_9968,N_8364);
xnor U10876 (N_10876,N_8653,N_9039);
xor U10877 (N_10877,N_9075,N_9253);
or U10878 (N_10878,N_9242,N_8243);
nor U10879 (N_10879,N_8257,N_8443);
xor U10880 (N_10880,N_9295,N_8340);
and U10881 (N_10881,N_9770,N_8754);
or U10882 (N_10882,N_9479,N_8137);
and U10883 (N_10883,N_8127,N_9169);
nand U10884 (N_10884,N_9683,N_8983);
nand U10885 (N_10885,N_8669,N_8904);
nor U10886 (N_10886,N_9975,N_9568);
and U10887 (N_10887,N_9455,N_8358);
and U10888 (N_10888,N_9480,N_9552);
nand U10889 (N_10889,N_8997,N_9208);
xor U10890 (N_10890,N_8092,N_8770);
nor U10891 (N_10891,N_8138,N_8606);
nor U10892 (N_10892,N_8227,N_9547);
nor U10893 (N_10893,N_8956,N_9580);
xnor U10894 (N_10894,N_9230,N_9510);
and U10895 (N_10895,N_9536,N_8631);
nand U10896 (N_10896,N_9764,N_8586);
and U10897 (N_10897,N_8506,N_9588);
or U10898 (N_10898,N_8913,N_8830);
and U10899 (N_10899,N_9786,N_8854);
nand U10900 (N_10900,N_9103,N_9494);
nand U10901 (N_10901,N_8809,N_9958);
nor U10902 (N_10902,N_9399,N_9483);
xor U10903 (N_10903,N_8145,N_9529);
nor U10904 (N_10904,N_9837,N_9079);
and U10905 (N_10905,N_8466,N_8465);
nor U10906 (N_10906,N_9648,N_9810);
and U10907 (N_10907,N_9507,N_8058);
nor U10908 (N_10908,N_8040,N_8749);
or U10909 (N_10909,N_8435,N_8043);
or U10910 (N_10910,N_9442,N_8488);
or U10911 (N_10911,N_8071,N_9150);
or U10912 (N_10912,N_9581,N_9989);
and U10913 (N_10913,N_9899,N_8870);
xnor U10914 (N_10914,N_8969,N_8545);
xor U10915 (N_10915,N_8277,N_9921);
or U10916 (N_10916,N_9328,N_8768);
and U10917 (N_10917,N_9448,N_8420);
and U10918 (N_10918,N_8140,N_8039);
xor U10919 (N_10919,N_9963,N_8797);
nand U10920 (N_10920,N_9525,N_8312);
or U10921 (N_10921,N_9270,N_9816);
xor U10922 (N_10922,N_8305,N_8463);
nand U10923 (N_10923,N_9500,N_9838);
xnor U10924 (N_10924,N_9811,N_9981);
nor U10925 (N_10925,N_9233,N_8842);
and U10926 (N_10926,N_8919,N_9622);
nor U10927 (N_10927,N_9412,N_8620);
and U10928 (N_10928,N_8837,N_8875);
xnor U10929 (N_10929,N_9891,N_9124);
nor U10930 (N_10930,N_8198,N_9335);
xnor U10931 (N_10931,N_8563,N_8704);
nand U10932 (N_10932,N_9807,N_8548);
xnor U10933 (N_10933,N_8639,N_9976);
nor U10934 (N_10934,N_8038,N_8196);
nor U10935 (N_10935,N_9389,N_8818);
xnor U10936 (N_10936,N_8193,N_8292);
nor U10937 (N_10937,N_8996,N_8635);
or U10938 (N_10938,N_9316,N_9373);
xnor U10939 (N_10939,N_8128,N_8397);
xnor U10940 (N_10940,N_9142,N_9834);
xnor U10941 (N_10941,N_8762,N_8028);
xor U10942 (N_10942,N_9514,N_9752);
nor U10943 (N_10943,N_9996,N_9538);
nand U10944 (N_10944,N_8119,N_9802);
and U10945 (N_10945,N_8293,N_8025);
or U10946 (N_10946,N_8415,N_9643);
nand U10947 (N_10947,N_8449,N_8320);
or U10948 (N_10948,N_8955,N_8879);
or U10949 (N_10949,N_8310,N_8526);
xnor U10950 (N_10950,N_8363,N_8775);
or U10951 (N_10951,N_8014,N_9900);
nor U10952 (N_10952,N_9711,N_8483);
xnor U10953 (N_10953,N_8676,N_9750);
xnor U10954 (N_10954,N_9259,N_9137);
and U10955 (N_10955,N_9050,N_9627);
xnor U10956 (N_10956,N_8619,N_9768);
xnor U10957 (N_10957,N_9106,N_9324);
and U10958 (N_10958,N_9705,N_8741);
or U10959 (N_10959,N_8911,N_9073);
or U10960 (N_10960,N_8649,N_9782);
xnor U10961 (N_10961,N_8084,N_8401);
xnor U10962 (N_10962,N_9688,N_8625);
nand U10963 (N_10963,N_9582,N_8813);
or U10964 (N_10964,N_8896,N_9640);
nand U10965 (N_10965,N_8680,N_9497);
and U10966 (N_10966,N_8633,N_9060);
nand U10967 (N_10967,N_9337,N_8106);
and U10968 (N_10968,N_9195,N_8195);
and U10969 (N_10969,N_9342,N_9401);
and U10970 (N_10970,N_8079,N_8971);
or U10971 (N_10971,N_8262,N_9610);
nand U10972 (N_10972,N_9477,N_9825);
nand U10973 (N_10973,N_9185,N_8504);
nor U10974 (N_10974,N_9322,N_9236);
nand U10975 (N_10975,N_8245,N_8355);
or U10976 (N_10976,N_9332,N_8843);
xor U10977 (N_10977,N_8072,N_8743);
xnor U10978 (N_10978,N_9933,N_9346);
nor U10979 (N_10979,N_8091,N_8887);
or U10980 (N_10980,N_8793,N_9980);
and U10981 (N_10981,N_9264,N_8947);
or U10982 (N_10982,N_8418,N_8249);
nand U10983 (N_10983,N_9179,N_8498);
xor U10984 (N_10984,N_8376,N_8113);
nor U10985 (N_10985,N_8302,N_8300);
or U10986 (N_10986,N_9430,N_9487);
and U10987 (N_10987,N_9107,N_8968);
or U10988 (N_10988,N_9237,N_9576);
and U10989 (N_10989,N_8613,N_8885);
and U10990 (N_10990,N_8339,N_9505);
and U10991 (N_10991,N_9682,N_9288);
xnor U10992 (N_10992,N_9699,N_8369);
nand U10993 (N_10993,N_9988,N_8325);
nor U10994 (N_10994,N_9458,N_8171);
nand U10995 (N_10995,N_9413,N_8658);
nand U10996 (N_10996,N_8104,N_9850);
and U10997 (N_10997,N_9326,N_9527);
and U10998 (N_10998,N_9644,N_9977);
nand U10999 (N_10999,N_9856,N_8779);
xor U11000 (N_11000,N_9524,N_8323);
nor U11001 (N_11001,N_9961,N_8384);
or U11002 (N_11002,N_8715,N_8218);
or U11003 (N_11003,N_8441,N_9668);
and U11004 (N_11004,N_9665,N_9640);
nand U11005 (N_11005,N_9790,N_8672);
or U11006 (N_11006,N_9082,N_8301);
xnor U11007 (N_11007,N_9524,N_9032);
and U11008 (N_11008,N_9101,N_8049);
nor U11009 (N_11009,N_9251,N_9551);
nor U11010 (N_11010,N_8965,N_8354);
nor U11011 (N_11011,N_9230,N_9602);
and U11012 (N_11012,N_9742,N_8691);
nor U11013 (N_11013,N_8647,N_9658);
xnor U11014 (N_11014,N_8530,N_9737);
nand U11015 (N_11015,N_8526,N_9549);
nand U11016 (N_11016,N_9402,N_8891);
and U11017 (N_11017,N_9534,N_9527);
nand U11018 (N_11018,N_8857,N_8376);
or U11019 (N_11019,N_9456,N_9155);
nor U11020 (N_11020,N_8411,N_9349);
nand U11021 (N_11021,N_8307,N_8339);
or U11022 (N_11022,N_9619,N_9929);
nand U11023 (N_11023,N_9030,N_8531);
xor U11024 (N_11024,N_9420,N_8192);
xnor U11025 (N_11025,N_8014,N_9044);
or U11026 (N_11026,N_8955,N_9814);
xnor U11027 (N_11027,N_9103,N_9891);
nor U11028 (N_11028,N_8999,N_8948);
and U11029 (N_11029,N_9477,N_9773);
nand U11030 (N_11030,N_8987,N_8738);
nand U11031 (N_11031,N_8331,N_9027);
and U11032 (N_11032,N_9949,N_9315);
and U11033 (N_11033,N_8490,N_8678);
or U11034 (N_11034,N_9666,N_9286);
and U11035 (N_11035,N_9875,N_9523);
nor U11036 (N_11036,N_8536,N_9193);
and U11037 (N_11037,N_8322,N_8903);
or U11038 (N_11038,N_8892,N_8759);
or U11039 (N_11039,N_8478,N_9302);
nand U11040 (N_11040,N_8507,N_8935);
nor U11041 (N_11041,N_9271,N_8314);
or U11042 (N_11042,N_8548,N_9630);
nand U11043 (N_11043,N_9823,N_9394);
nor U11044 (N_11044,N_8748,N_8531);
nand U11045 (N_11045,N_9454,N_8869);
and U11046 (N_11046,N_9086,N_8304);
xor U11047 (N_11047,N_8532,N_9922);
and U11048 (N_11048,N_8202,N_9765);
nand U11049 (N_11049,N_9999,N_8728);
and U11050 (N_11050,N_9445,N_8539);
nor U11051 (N_11051,N_8537,N_9715);
nor U11052 (N_11052,N_9719,N_9885);
nor U11053 (N_11053,N_8555,N_9705);
nor U11054 (N_11054,N_8596,N_8616);
or U11055 (N_11055,N_8035,N_8675);
or U11056 (N_11056,N_9956,N_8337);
and U11057 (N_11057,N_9326,N_9748);
or U11058 (N_11058,N_8221,N_9129);
nor U11059 (N_11059,N_8556,N_8954);
nand U11060 (N_11060,N_9791,N_8153);
or U11061 (N_11061,N_8909,N_9398);
or U11062 (N_11062,N_9668,N_9146);
and U11063 (N_11063,N_9932,N_8171);
nor U11064 (N_11064,N_9582,N_9394);
nand U11065 (N_11065,N_9949,N_8374);
xnor U11066 (N_11066,N_8293,N_8469);
or U11067 (N_11067,N_8984,N_9243);
and U11068 (N_11068,N_9346,N_8800);
and U11069 (N_11069,N_9979,N_8929);
xor U11070 (N_11070,N_8032,N_8167);
and U11071 (N_11071,N_8193,N_9625);
and U11072 (N_11072,N_8193,N_9673);
and U11073 (N_11073,N_8676,N_9724);
nand U11074 (N_11074,N_9059,N_8240);
xor U11075 (N_11075,N_8960,N_9633);
nor U11076 (N_11076,N_9097,N_8566);
nand U11077 (N_11077,N_8479,N_8143);
xnor U11078 (N_11078,N_9059,N_9992);
nor U11079 (N_11079,N_8764,N_8620);
xor U11080 (N_11080,N_8041,N_9250);
and U11081 (N_11081,N_8563,N_9912);
nor U11082 (N_11082,N_8734,N_8826);
xnor U11083 (N_11083,N_8422,N_9865);
xor U11084 (N_11084,N_9512,N_9920);
xnor U11085 (N_11085,N_9438,N_8969);
nor U11086 (N_11086,N_8067,N_9842);
xor U11087 (N_11087,N_9252,N_8668);
nand U11088 (N_11088,N_9428,N_9346);
and U11089 (N_11089,N_8066,N_8092);
xnor U11090 (N_11090,N_8745,N_8750);
nor U11091 (N_11091,N_9354,N_8010);
nand U11092 (N_11092,N_9709,N_8164);
and U11093 (N_11093,N_8603,N_8278);
or U11094 (N_11094,N_9942,N_8166);
and U11095 (N_11095,N_8607,N_8520);
nor U11096 (N_11096,N_9556,N_9990);
xor U11097 (N_11097,N_8827,N_9500);
or U11098 (N_11098,N_9389,N_8737);
or U11099 (N_11099,N_9097,N_8276);
nor U11100 (N_11100,N_8669,N_8413);
nor U11101 (N_11101,N_8322,N_8910);
and U11102 (N_11102,N_8766,N_9659);
nand U11103 (N_11103,N_9260,N_9265);
nor U11104 (N_11104,N_8876,N_9371);
and U11105 (N_11105,N_8866,N_9162);
xnor U11106 (N_11106,N_8470,N_9897);
xnor U11107 (N_11107,N_9124,N_8007);
nand U11108 (N_11108,N_8124,N_8415);
or U11109 (N_11109,N_8370,N_8498);
or U11110 (N_11110,N_9343,N_9734);
nand U11111 (N_11111,N_9853,N_8232);
nor U11112 (N_11112,N_8521,N_8888);
xor U11113 (N_11113,N_8486,N_8543);
nor U11114 (N_11114,N_8444,N_9430);
nand U11115 (N_11115,N_8576,N_9461);
or U11116 (N_11116,N_8401,N_8089);
nand U11117 (N_11117,N_8316,N_8327);
nor U11118 (N_11118,N_9994,N_9299);
or U11119 (N_11119,N_8303,N_8236);
nor U11120 (N_11120,N_8036,N_9866);
xor U11121 (N_11121,N_8549,N_9914);
or U11122 (N_11122,N_8168,N_9642);
xor U11123 (N_11123,N_9795,N_9419);
nand U11124 (N_11124,N_8992,N_8107);
or U11125 (N_11125,N_8138,N_9443);
xnor U11126 (N_11126,N_9465,N_8865);
nand U11127 (N_11127,N_8817,N_9487);
xor U11128 (N_11128,N_9323,N_9539);
and U11129 (N_11129,N_8899,N_9948);
or U11130 (N_11130,N_8056,N_8178);
or U11131 (N_11131,N_9230,N_8487);
and U11132 (N_11132,N_9349,N_8816);
xor U11133 (N_11133,N_8180,N_9019);
xor U11134 (N_11134,N_9546,N_9420);
or U11135 (N_11135,N_8751,N_8873);
or U11136 (N_11136,N_9826,N_8828);
or U11137 (N_11137,N_9270,N_8552);
and U11138 (N_11138,N_8601,N_9479);
nand U11139 (N_11139,N_8652,N_9742);
and U11140 (N_11140,N_9169,N_8736);
xor U11141 (N_11141,N_9783,N_9473);
or U11142 (N_11142,N_9506,N_9872);
and U11143 (N_11143,N_9719,N_8856);
nand U11144 (N_11144,N_8895,N_8331);
nand U11145 (N_11145,N_8897,N_8415);
nand U11146 (N_11146,N_9630,N_9265);
or U11147 (N_11147,N_9428,N_9676);
nand U11148 (N_11148,N_8661,N_8252);
nor U11149 (N_11149,N_8655,N_8653);
xnor U11150 (N_11150,N_8434,N_8072);
nand U11151 (N_11151,N_8162,N_9781);
or U11152 (N_11152,N_9591,N_9924);
xnor U11153 (N_11153,N_9158,N_8613);
nand U11154 (N_11154,N_8343,N_9410);
and U11155 (N_11155,N_8072,N_9031);
and U11156 (N_11156,N_9171,N_8209);
nand U11157 (N_11157,N_8748,N_9181);
or U11158 (N_11158,N_9894,N_9789);
and U11159 (N_11159,N_8282,N_9154);
or U11160 (N_11160,N_8824,N_9540);
xor U11161 (N_11161,N_8359,N_8276);
nand U11162 (N_11162,N_9786,N_9760);
nor U11163 (N_11163,N_8915,N_9213);
xnor U11164 (N_11164,N_9727,N_9170);
and U11165 (N_11165,N_9763,N_9277);
xnor U11166 (N_11166,N_8395,N_9638);
nor U11167 (N_11167,N_9459,N_9114);
or U11168 (N_11168,N_8728,N_8820);
and U11169 (N_11169,N_9598,N_8117);
and U11170 (N_11170,N_9079,N_9157);
nand U11171 (N_11171,N_8204,N_8237);
nand U11172 (N_11172,N_8084,N_9978);
xnor U11173 (N_11173,N_8512,N_9261);
xor U11174 (N_11174,N_9919,N_8334);
nand U11175 (N_11175,N_9099,N_9161);
nor U11176 (N_11176,N_8068,N_8610);
or U11177 (N_11177,N_9312,N_9349);
nand U11178 (N_11178,N_9705,N_8359);
xor U11179 (N_11179,N_9825,N_8716);
nor U11180 (N_11180,N_8111,N_9848);
nor U11181 (N_11181,N_9787,N_8713);
nand U11182 (N_11182,N_8060,N_9062);
or U11183 (N_11183,N_9468,N_8309);
xnor U11184 (N_11184,N_9626,N_9973);
xor U11185 (N_11185,N_9440,N_8543);
xnor U11186 (N_11186,N_9682,N_9635);
nor U11187 (N_11187,N_8843,N_9290);
xnor U11188 (N_11188,N_9636,N_9914);
nand U11189 (N_11189,N_9536,N_8495);
and U11190 (N_11190,N_9415,N_8271);
xor U11191 (N_11191,N_8360,N_8293);
and U11192 (N_11192,N_9090,N_8189);
or U11193 (N_11193,N_9473,N_8424);
and U11194 (N_11194,N_9068,N_9823);
or U11195 (N_11195,N_8899,N_9228);
or U11196 (N_11196,N_9509,N_9283);
nand U11197 (N_11197,N_8077,N_8857);
and U11198 (N_11198,N_8300,N_9046);
and U11199 (N_11199,N_9978,N_8506);
and U11200 (N_11200,N_8932,N_9901);
xor U11201 (N_11201,N_9557,N_9749);
or U11202 (N_11202,N_8673,N_8503);
and U11203 (N_11203,N_9204,N_9473);
and U11204 (N_11204,N_8644,N_9516);
xnor U11205 (N_11205,N_8278,N_9449);
or U11206 (N_11206,N_8130,N_8979);
nor U11207 (N_11207,N_9379,N_9155);
nor U11208 (N_11208,N_8401,N_8026);
or U11209 (N_11209,N_8302,N_9745);
nand U11210 (N_11210,N_9315,N_8866);
nor U11211 (N_11211,N_8325,N_9468);
and U11212 (N_11212,N_9591,N_9521);
xnor U11213 (N_11213,N_9568,N_8992);
xnor U11214 (N_11214,N_9310,N_9991);
nor U11215 (N_11215,N_8537,N_9519);
and U11216 (N_11216,N_8192,N_8786);
xor U11217 (N_11217,N_8638,N_9517);
nor U11218 (N_11218,N_8129,N_8876);
nor U11219 (N_11219,N_8200,N_8352);
nand U11220 (N_11220,N_9572,N_8561);
xor U11221 (N_11221,N_9269,N_9860);
nor U11222 (N_11222,N_8312,N_8462);
nand U11223 (N_11223,N_8343,N_9671);
nor U11224 (N_11224,N_8891,N_9758);
xor U11225 (N_11225,N_8056,N_8947);
nand U11226 (N_11226,N_8618,N_8972);
and U11227 (N_11227,N_8850,N_8224);
or U11228 (N_11228,N_8588,N_8355);
nand U11229 (N_11229,N_8592,N_8422);
and U11230 (N_11230,N_9431,N_9416);
or U11231 (N_11231,N_9038,N_9844);
nor U11232 (N_11232,N_9923,N_8212);
nor U11233 (N_11233,N_8588,N_9455);
nor U11234 (N_11234,N_8758,N_9611);
and U11235 (N_11235,N_9538,N_9219);
nand U11236 (N_11236,N_9070,N_8062);
xnor U11237 (N_11237,N_9415,N_9293);
or U11238 (N_11238,N_9889,N_8854);
nor U11239 (N_11239,N_9966,N_8686);
nand U11240 (N_11240,N_9231,N_8852);
nand U11241 (N_11241,N_8356,N_8759);
or U11242 (N_11242,N_8415,N_8833);
nor U11243 (N_11243,N_8704,N_8992);
nor U11244 (N_11244,N_9635,N_9487);
or U11245 (N_11245,N_9530,N_8443);
and U11246 (N_11246,N_8006,N_9342);
nand U11247 (N_11247,N_9091,N_8328);
and U11248 (N_11248,N_8713,N_9048);
nand U11249 (N_11249,N_8573,N_9508);
nor U11250 (N_11250,N_9952,N_8297);
nand U11251 (N_11251,N_8557,N_9539);
nand U11252 (N_11252,N_9880,N_8702);
or U11253 (N_11253,N_8622,N_9553);
and U11254 (N_11254,N_8962,N_9280);
and U11255 (N_11255,N_9148,N_8201);
nor U11256 (N_11256,N_8969,N_9611);
nor U11257 (N_11257,N_8670,N_9305);
nand U11258 (N_11258,N_8340,N_9469);
xnor U11259 (N_11259,N_9672,N_9190);
and U11260 (N_11260,N_9424,N_8757);
or U11261 (N_11261,N_8709,N_9670);
or U11262 (N_11262,N_9558,N_9685);
xnor U11263 (N_11263,N_8986,N_9013);
and U11264 (N_11264,N_9056,N_8314);
and U11265 (N_11265,N_9571,N_8822);
nand U11266 (N_11266,N_9709,N_9773);
and U11267 (N_11267,N_8335,N_8392);
xnor U11268 (N_11268,N_9200,N_9187);
nor U11269 (N_11269,N_8719,N_8652);
or U11270 (N_11270,N_8261,N_8800);
and U11271 (N_11271,N_8191,N_8472);
xnor U11272 (N_11272,N_9731,N_8170);
xnor U11273 (N_11273,N_8669,N_8841);
or U11274 (N_11274,N_8937,N_9250);
or U11275 (N_11275,N_9505,N_9419);
and U11276 (N_11276,N_9543,N_8080);
xnor U11277 (N_11277,N_8212,N_8733);
nor U11278 (N_11278,N_9992,N_9021);
xnor U11279 (N_11279,N_9294,N_9875);
nor U11280 (N_11280,N_9942,N_8434);
xor U11281 (N_11281,N_9630,N_8685);
xor U11282 (N_11282,N_8816,N_9684);
nor U11283 (N_11283,N_8932,N_9905);
nand U11284 (N_11284,N_9226,N_8047);
nor U11285 (N_11285,N_8979,N_9507);
nor U11286 (N_11286,N_9182,N_8155);
nor U11287 (N_11287,N_9705,N_8140);
nor U11288 (N_11288,N_9758,N_8453);
xnor U11289 (N_11289,N_9339,N_8911);
nand U11290 (N_11290,N_9614,N_9502);
and U11291 (N_11291,N_8288,N_9315);
xor U11292 (N_11292,N_9843,N_8218);
nand U11293 (N_11293,N_8591,N_8398);
and U11294 (N_11294,N_9408,N_8105);
or U11295 (N_11295,N_9727,N_8388);
xor U11296 (N_11296,N_9188,N_9925);
nor U11297 (N_11297,N_9110,N_8459);
nor U11298 (N_11298,N_9792,N_9110);
nor U11299 (N_11299,N_8144,N_9969);
nand U11300 (N_11300,N_8988,N_8200);
nor U11301 (N_11301,N_9488,N_9071);
or U11302 (N_11302,N_9705,N_8774);
or U11303 (N_11303,N_8392,N_9544);
or U11304 (N_11304,N_9580,N_9649);
and U11305 (N_11305,N_9337,N_8102);
and U11306 (N_11306,N_9415,N_8513);
nand U11307 (N_11307,N_9716,N_8809);
and U11308 (N_11308,N_9204,N_8388);
nand U11309 (N_11309,N_8608,N_8023);
nand U11310 (N_11310,N_9066,N_9712);
nand U11311 (N_11311,N_8088,N_8739);
nand U11312 (N_11312,N_8735,N_9700);
nor U11313 (N_11313,N_9997,N_8990);
nor U11314 (N_11314,N_8040,N_9471);
or U11315 (N_11315,N_9411,N_8047);
or U11316 (N_11316,N_9206,N_9880);
nand U11317 (N_11317,N_8950,N_9574);
xnor U11318 (N_11318,N_9736,N_9602);
and U11319 (N_11319,N_9804,N_9501);
nor U11320 (N_11320,N_9235,N_9098);
and U11321 (N_11321,N_8504,N_9236);
xnor U11322 (N_11322,N_8782,N_9609);
and U11323 (N_11323,N_8824,N_9119);
xor U11324 (N_11324,N_8719,N_8351);
nand U11325 (N_11325,N_9762,N_8776);
xor U11326 (N_11326,N_9093,N_9124);
or U11327 (N_11327,N_8207,N_8606);
or U11328 (N_11328,N_8842,N_8959);
or U11329 (N_11329,N_9242,N_9778);
xor U11330 (N_11330,N_8301,N_9456);
nand U11331 (N_11331,N_8833,N_8708);
xor U11332 (N_11332,N_8406,N_9896);
or U11333 (N_11333,N_9230,N_9150);
or U11334 (N_11334,N_9150,N_9428);
xnor U11335 (N_11335,N_8663,N_9951);
nand U11336 (N_11336,N_9130,N_8897);
xor U11337 (N_11337,N_8424,N_9188);
xor U11338 (N_11338,N_8524,N_9884);
nand U11339 (N_11339,N_8649,N_9844);
nand U11340 (N_11340,N_9463,N_8411);
and U11341 (N_11341,N_9789,N_9455);
xor U11342 (N_11342,N_9123,N_9461);
xnor U11343 (N_11343,N_9784,N_8600);
nor U11344 (N_11344,N_9599,N_8265);
and U11345 (N_11345,N_8416,N_8532);
and U11346 (N_11346,N_8715,N_9073);
nand U11347 (N_11347,N_9545,N_8225);
and U11348 (N_11348,N_8968,N_9705);
or U11349 (N_11349,N_8329,N_9953);
and U11350 (N_11350,N_8332,N_9775);
nand U11351 (N_11351,N_9972,N_8985);
nand U11352 (N_11352,N_8922,N_9690);
nor U11353 (N_11353,N_8700,N_8643);
nand U11354 (N_11354,N_8691,N_9641);
xor U11355 (N_11355,N_8414,N_9996);
nor U11356 (N_11356,N_8273,N_9805);
or U11357 (N_11357,N_9883,N_8956);
nand U11358 (N_11358,N_8117,N_8508);
nand U11359 (N_11359,N_8936,N_8120);
nor U11360 (N_11360,N_8970,N_8063);
and U11361 (N_11361,N_9780,N_8910);
nand U11362 (N_11362,N_9575,N_9580);
or U11363 (N_11363,N_8012,N_9281);
nor U11364 (N_11364,N_9169,N_8597);
nand U11365 (N_11365,N_8993,N_8327);
or U11366 (N_11366,N_9338,N_9658);
and U11367 (N_11367,N_8573,N_8234);
xor U11368 (N_11368,N_9353,N_9025);
nand U11369 (N_11369,N_8150,N_8883);
nand U11370 (N_11370,N_8877,N_9233);
nand U11371 (N_11371,N_8649,N_8305);
xnor U11372 (N_11372,N_8806,N_8218);
or U11373 (N_11373,N_8400,N_9041);
or U11374 (N_11374,N_8737,N_8470);
and U11375 (N_11375,N_9181,N_9778);
nand U11376 (N_11376,N_8712,N_8943);
or U11377 (N_11377,N_9897,N_9727);
nor U11378 (N_11378,N_9959,N_9061);
or U11379 (N_11379,N_9658,N_8616);
nand U11380 (N_11380,N_9638,N_9229);
and U11381 (N_11381,N_9714,N_9801);
or U11382 (N_11382,N_9066,N_9210);
and U11383 (N_11383,N_9474,N_8686);
or U11384 (N_11384,N_9968,N_8652);
or U11385 (N_11385,N_9164,N_8136);
nand U11386 (N_11386,N_8265,N_8873);
or U11387 (N_11387,N_8616,N_9592);
or U11388 (N_11388,N_9545,N_9932);
nand U11389 (N_11389,N_8275,N_9928);
xor U11390 (N_11390,N_8527,N_9354);
nand U11391 (N_11391,N_8803,N_8907);
xnor U11392 (N_11392,N_8007,N_8967);
nand U11393 (N_11393,N_8952,N_8091);
nor U11394 (N_11394,N_8990,N_8552);
or U11395 (N_11395,N_9841,N_8388);
and U11396 (N_11396,N_9796,N_9274);
nand U11397 (N_11397,N_9672,N_8265);
nor U11398 (N_11398,N_9728,N_9220);
xor U11399 (N_11399,N_9863,N_9237);
nand U11400 (N_11400,N_9776,N_9722);
nand U11401 (N_11401,N_9335,N_9944);
nand U11402 (N_11402,N_8942,N_8853);
or U11403 (N_11403,N_8952,N_8310);
or U11404 (N_11404,N_9028,N_9001);
nand U11405 (N_11405,N_9618,N_9197);
nor U11406 (N_11406,N_8293,N_9362);
and U11407 (N_11407,N_9325,N_8035);
xor U11408 (N_11408,N_9346,N_9074);
xnor U11409 (N_11409,N_9815,N_9675);
xnor U11410 (N_11410,N_9293,N_9857);
nor U11411 (N_11411,N_9632,N_8976);
or U11412 (N_11412,N_8171,N_9634);
nand U11413 (N_11413,N_8172,N_9872);
and U11414 (N_11414,N_8603,N_8126);
nand U11415 (N_11415,N_9731,N_8367);
or U11416 (N_11416,N_9031,N_8625);
and U11417 (N_11417,N_9814,N_8244);
or U11418 (N_11418,N_8041,N_8069);
and U11419 (N_11419,N_8478,N_8845);
nor U11420 (N_11420,N_9173,N_9956);
and U11421 (N_11421,N_9637,N_9688);
and U11422 (N_11422,N_9682,N_8038);
and U11423 (N_11423,N_8189,N_8416);
xor U11424 (N_11424,N_9243,N_8951);
nand U11425 (N_11425,N_8491,N_9828);
and U11426 (N_11426,N_9399,N_9585);
nor U11427 (N_11427,N_8419,N_8847);
or U11428 (N_11428,N_9197,N_8272);
xnor U11429 (N_11429,N_8559,N_8305);
xor U11430 (N_11430,N_8354,N_9538);
xor U11431 (N_11431,N_8416,N_8482);
xnor U11432 (N_11432,N_8783,N_9954);
nor U11433 (N_11433,N_9798,N_9692);
nor U11434 (N_11434,N_9500,N_9642);
nand U11435 (N_11435,N_8069,N_8632);
and U11436 (N_11436,N_9769,N_9914);
xor U11437 (N_11437,N_8026,N_9570);
and U11438 (N_11438,N_9898,N_9073);
and U11439 (N_11439,N_8694,N_8386);
nor U11440 (N_11440,N_8857,N_8306);
or U11441 (N_11441,N_8859,N_9568);
or U11442 (N_11442,N_8713,N_9235);
xnor U11443 (N_11443,N_9974,N_8472);
nor U11444 (N_11444,N_9950,N_8644);
or U11445 (N_11445,N_9231,N_9315);
and U11446 (N_11446,N_9330,N_8928);
xnor U11447 (N_11447,N_8891,N_8703);
xnor U11448 (N_11448,N_8630,N_9966);
or U11449 (N_11449,N_8791,N_8491);
xnor U11450 (N_11450,N_9537,N_8281);
nor U11451 (N_11451,N_9432,N_8922);
or U11452 (N_11452,N_9060,N_8805);
and U11453 (N_11453,N_9564,N_8547);
xnor U11454 (N_11454,N_8001,N_8188);
and U11455 (N_11455,N_8387,N_8340);
or U11456 (N_11456,N_8423,N_9107);
nand U11457 (N_11457,N_8499,N_8879);
nor U11458 (N_11458,N_9527,N_8558);
xnor U11459 (N_11459,N_8867,N_9755);
xor U11460 (N_11460,N_8553,N_8415);
and U11461 (N_11461,N_8832,N_8241);
and U11462 (N_11462,N_9781,N_9448);
nand U11463 (N_11463,N_8905,N_8222);
xor U11464 (N_11464,N_8832,N_9742);
nand U11465 (N_11465,N_8478,N_8831);
and U11466 (N_11466,N_8382,N_8835);
or U11467 (N_11467,N_8159,N_9919);
nand U11468 (N_11468,N_8924,N_8132);
or U11469 (N_11469,N_9785,N_8058);
nand U11470 (N_11470,N_8762,N_9075);
nand U11471 (N_11471,N_8303,N_8480);
nand U11472 (N_11472,N_9612,N_8424);
and U11473 (N_11473,N_8372,N_9978);
nor U11474 (N_11474,N_8360,N_9274);
xor U11475 (N_11475,N_8924,N_9558);
xor U11476 (N_11476,N_8903,N_8941);
xnor U11477 (N_11477,N_8804,N_9236);
xor U11478 (N_11478,N_9009,N_8273);
nor U11479 (N_11479,N_8926,N_9094);
xor U11480 (N_11480,N_9135,N_8542);
xor U11481 (N_11481,N_9963,N_9357);
nor U11482 (N_11482,N_8772,N_8518);
nand U11483 (N_11483,N_9910,N_8140);
and U11484 (N_11484,N_9937,N_9282);
xor U11485 (N_11485,N_8848,N_8803);
nor U11486 (N_11486,N_8981,N_8003);
nor U11487 (N_11487,N_8742,N_8768);
and U11488 (N_11488,N_9484,N_9379);
xor U11489 (N_11489,N_8937,N_9247);
xor U11490 (N_11490,N_8357,N_9649);
and U11491 (N_11491,N_8198,N_9318);
and U11492 (N_11492,N_9893,N_9075);
xnor U11493 (N_11493,N_8250,N_9376);
xor U11494 (N_11494,N_9555,N_9812);
and U11495 (N_11495,N_8893,N_9521);
and U11496 (N_11496,N_8098,N_8935);
nand U11497 (N_11497,N_9849,N_9071);
or U11498 (N_11498,N_9678,N_9260);
nor U11499 (N_11499,N_8033,N_9924);
nand U11500 (N_11500,N_9607,N_9725);
nor U11501 (N_11501,N_9497,N_9515);
and U11502 (N_11502,N_8091,N_8561);
or U11503 (N_11503,N_9527,N_8938);
nand U11504 (N_11504,N_8867,N_8495);
xor U11505 (N_11505,N_8977,N_8111);
nor U11506 (N_11506,N_8557,N_9122);
nor U11507 (N_11507,N_8621,N_8316);
or U11508 (N_11508,N_8376,N_8566);
xor U11509 (N_11509,N_9759,N_9679);
nor U11510 (N_11510,N_9217,N_8844);
nand U11511 (N_11511,N_8131,N_9758);
and U11512 (N_11512,N_8405,N_9600);
xnor U11513 (N_11513,N_8914,N_8097);
and U11514 (N_11514,N_9317,N_8589);
xor U11515 (N_11515,N_8666,N_8465);
xnor U11516 (N_11516,N_8927,N_9925);
and U11517 (N_11517,N_8939,N_9236);
or U11518 (N_11518,N_9197,N_8317);
nand U11519 (N_11519,N_9919,N_8121);
xor U11520 (N_11520,N_8685,N_9698);
nor U11521 (N_11521,N_9233,N_8723);
and U11522 (N_11522,N_9759,N_8088);
nor U11523 (N_11523,N_8526,N_9384);
or U11524 (N_11524,N_9357,N_8471);
nand U11525 (N_11525,N_9381,N_9514);
or U11526 (N_11526,N_9040,N_8118);
nand U11527 (N_11527,N_9159,N_8687);
and U11528 (N_11528,N_8750,N_9378);
xor U11529 (N_11529,N_8855,N_8993);
nand U11530 (N_11530,N_9932,N_9333);
and U11531 (N_11531,N_9759,N_9793);
nor U11532 (N_11532,N_9600,N_8493);
and U11533 (N_11533,N_8008,N_9277);
xor U11534 (N_11534,N_8174,N_9378);
or U11535 (N_11535,N_8461,N_8800);
nor U11536 (N_11536,N_9692,N_9130);
or U11537 (N_11537,N_9555,N_8896);
or U11538 (N_11538,N_8926,N_8731);
nor U11539 (N_11539,N_8654,N_9599);
nor U11540 (N_11540,N_9079,N_9260);
and U11541 (N_11541,N_9097,N_9214);
nand U11542 (N_11542,N_8499,N_9981);
nor U11543 (N_11543,N_9135,N_9281);
nand U11544 (N_11544,N_9480,N_9257);
nor U11545 (N_11545,N_9424,N_8489);
xnor U11546 (N_11546,N_8893,N_8106);
or U11547 (N_11547,N_9272,N_9501);
nand U11548 (N_11548,N_8543,N_8295);
and U11549 (N_11549,N_8877,N_9591);
or U11550 (N_11550,N_9784,N_9660);
nor U11551 (N_11551,N_8703,N_9808);
xnor U11552 (N_11552,N_8503,N_8559);
xor U11553 (N_11553,N_9636,N_9601);
nand U11554 (N_11554,N_8252,N_8289);
xor U11555 (N_11555,N_8373,N_9374);
nor U11556 (N_11556,N_9995,N_9839);
xnor U11557 (N_11557,N_8932,N_9208);
and U11558 (N_11558,N_8822,N_8284);
or U11559 (N_11559,N_9201,N_8432);
xnor U11560 (N_11560,N_9082,N_8613);
xor U11561 (N_11561,N_8804,N_8192);
nand U11562 (N_11562,N_9357,N_8829);
and U11563 (N_11563,N_8737,N_9348);
nor U11564 (N_11564,N_8224,N_8707);
or U11565 (N_11565,N_8759,N_9144);
nand U11566 (N_11566,N_8050,N_9685);
nor U11567 (N_11567,N_8475,N_8517);
nand U11568 (N_11568,N_8591,N_8046);
nor U11569 (N_11569,N_8234,N_9200);
or U11570 (N_11570,N_8867,N_8993);
and U11571 (N_11571,N_8843,N_9145);
xnor U11572 (N_11572,N_8033,N_9441);
and U11573 (N_11573,N_8229,N_9082);
nor U11574 (N_11574,N_9045,N_9770);
nand U11575 (N_11575,N_9591,N_8257);
xnor U11576 (N_11576,N_8729,N_8270);
and U11577 (N_11577,N_9896,N_9071);
and U11578 (N_11578,N_8599,N_8273);
nor U11579 (N_11579,N_8871,N_9355);
nor U11580 (N_11580,N_9675,N_8900);
nor U11581 (N_11581,N_9926,N_8845);
xor U11582 (N_11582,N_9405,N_9181);
nand U11583 (N_11583,N_9287,N_8839);
and U11584 (N_11584,N_8400,N_9819);
xor U11585 (N_11585,N_9687,N_9109);
nor U11586 (N_11586,N_9253,N_8346);
xnor U11587 (N_11587,N_9252,N_8989);
and U11588 (N_11588,N_9676,N_8458);
xor U11589 (N_11589,N_8277,N_8654);
xor U11590 (N_11590,N_9514,N_9560);
nor U11591 (N_11591,N_9059,N_9649);
xor U11592 (N_11592,N_8547,N_9083);
nor U11593 (N_11593,N_9082,N_8342);
xor U11594 (N_11594,N_9780,N_9658);
and U11595 (N_11595,N_8943,N_8972);
nand U11596 (N_11596,N_8636,N_9453);
nor U11597 (N_11597,N_9768,N_9263);
nand U11598 (N_11598,N_9346,N_8267);
nor U11599 (N_11599,N_9894,N_9955);
and U11600 (N_11600,N_9474,N_9047);
nor U11601 (N_11601,N_8660,N_8452);
xnor U11602 (N_11602,N_8717,N_8632);
nand U11603 (N_11603,N_8960,N_8181);
nand U11604 (N_11604,N_8071,N_9077);
xor U11605 (N_11605,N_9732,N_8877);
or U11606 (N_11606,N_8294,N_8908);
nand U11607 (N_11607,N_8011,N_9397);
and U11608 (N_11608,N_8327,N_9342);
nand U11609 (N_11609,N_9207,N_8396);
xnor U11610 (N_11610,N_9595,N_8640);
xnor U11611 (N_11611,N_9025,N_8774);
nand U11612 (N_11612,N_8104,N_8479);
xnor U11613 (N_11613,N_9831,N_9460);
nand U11614 (N_11614,N_9459,N_9396);
nand U11615 (N_11615,N_8303,N_8800);
xor U11616 (N_11616,N_9675,N_8805);
nand U11617 (N_11617,N_8286,N_8690);
nand U11618 (N_11618,N_9203,N_8697);
xor U11619 (N_11619,N_9078,N_9404);
or U11620 (N_11620,N_8012,N_8825);
nand U11621 (N_11621,N_9708,N_8427);
xor U11622 (N_11622,N_8958,N_9385);
nor U11623 (N_11623,N_9009,N_8291);
nand U11624 (N_11624,N_9230,N_8272);
xnor U11625 (N_11625,N_8492,N_9014);
nor U11626 (N_11626,N_9956,N_9158);
nand U11627 (N_11627,N_8386,N_8558);
or U11628 (N_11628,N_8480,N_9793);
xor U11629 (N_11629,N_9474,N_8969);
xor U11630 (N_11630,N_8505,N_9277);
and U11631 (N_11631,N_9802,N_9437);
nor U11632 (N_11632,N_8288,N_8890);
nand U11633 (N_11633,N_9640,N_8823);
or U11634 (N_11634,N_9489,N_8174);
or U11635 (N_11635,N_8497,N_9777);
and U11636 (N_11636,N_9682,N_9334);
nand U11637 (N_11637,N_9321,N_9313);
xor U11638 (N_11638,N_8151,N_9721);
xor U11639 (N_11639,N_8379,N_8811);
or U11640 (N_11640,N_8825,N_9665);
and U11641 (N_11641,N_8067,N_8170);
nor U11642 (N_11642,N_9647,N_9482);
nand U11643 (N_11643,N_9821,N_9317);
or U11644 (N_11644,N_8730,N_8367);
nand U11645 (N_11645,N_9961,N_8853);
nand U11646 (N_11646,N_9226,N_8948);
xnor U11647 (N_11647,N_9962,N_9826);
nand U11648 (N_11648,N_8962,N_9224);
nor U11649 (N_11649,N_8238,N_8092);
and U11650 (N_11650,N_9807,N_9936);
or U11651 (N_11651,N_8684,N_8007);
xor U11652 (N_11652,N_9457,N_8412);
xor U11653 (N_11653,N_8996,N_8165);
xor U11654 (N_11654,N_8171,N_8044);
xor U11655 (N_11655,N_9371,N_9897);
nand U11656 (N_11656,N_8689,N_8908);
or U11657 (N_11657,N_8920,N_8659);
xnor U11658 (N_11658,N_8050,N_9442);
xor U11659 (N_11659,N_9022,N_8920);
or U11660 (N_11660,N_9061,N_8505);
and U11661 (N_11661,N_8011,N_9000);
or U11662 (N_11662,N_9995,N_8346);
or U11663 (N_11663,N_8331,N_9115);
or U11664 (N_11664,N_8243,N_8477);
nand U11665 (N_11665,N_8647,N_9985);
nand U11666 (N_11666,N_8308,N_8583);
and U11667 (N_11667,N_8727,N_9325);
xnor U11668 (N_11668,N_8286,N_8994);
nor U11669 (N_11669,N_8179,N_8053);
and U11670 (N_11670,N_8251,N_8277);
nor U11671 (N_11671,N_9474,N_8218);
nor U11672 (N_11672,N_9288,N_9247);
nand U11673 (N_11673,N_8644,N_8185);
xnor U11674 (N_11674,N_8834,N_8174);
or U11675 (N_11675,N_9694,N_9828);
xor U11676 (N_11676,N_9492,N_8520);
nand U11677 (N_11677,N_8537,N_9580);
nand U11678 (N_11678,N_8706,N_9579);
and U11679 (N_11679,N_8932,N_9512);
nor U11680 (N_11680,N_8478,N_9468);
nand U11681 (N_11681,N_8690,N_8438);
and U11682 (N_11682,N_8407,N_8962);
xor U11683 (N_11683,N_8310,N_8260);
xor U11684 (N_11684,N_9627,N_8053);
xnor U11685 (N_11685,N_8607,N_9748);
xnor U11686 (N_11686,N_9629,N_8169);
nor U11687 (N_11687,N_9061,N_8617);
xnor U11688 (N_11688,N_9984,N_8888);
xnor U11689 (N_11689,N_8724,N_8428);
xnor U11690 (N_11690,N_8097,N_8860);
xnor U11691 (N_11691,N_9786,N_8487);
and U11692 (N_11692,N_9329,N_9518);
or U11693 (N_11693,N_8012,N_9658);
and U11694 (N_11694,N_8004,N_8256);
nor U11695 (N_11695,N_8351,N_9438);
nand U11696 (N_11696,N_9428,N_8759);
nand U11697 (N_11697,N_9925,N_9596);
and U11698 (N_11698,N_8674,N_9295);
nor U11699 (N_11699,N_8144,N_8621);
or U11700 (N_11700,N_9917,N_8591);
and U11701 (N_11701,N_9861,N_9400);
and U11702 (N_11702,N_8971,N_9242);
or U11703 (N_11703,N_9403,N_9047);
nand U11704 (N_11704,N_8443,N_9748);
xor U11705 (N_11705,N_9842,N_9644);
and U11706 (N_11706,N_8774,N_9124);
or U11707 (N_11707,N_9446,N_9967);
or U11708 (N_11708,N_9826,N_9681);
nor U11709 (N_11709,N_9302,N_9287);
nand U11710 (N_11710,N_8271,N_8052);
or U11711 (N_11711,N_8919,N_9851);
xor U11712 (N_11712,N_8398,N_9514);
nor U11713 (N_11713,N_8958,N_9273);
or U11714 (N_11714,N_9329,N_9407);
nand U11715 (N_11715,N_8390,N_9958);
nand U11716 (N_11716,N_8803,N_9776);
or U11717 (N_11717,N_8918,N_9464);
or U11718 (N_11718,N_8073,N_8400);
xor U11719 (N_11719,N_9447,N_8951);
xor U11720 (N_11720,N_8608,N_8857);
nor U11721 (N_11721,N_8040,N_8485);
or U11722 (N_11722,N_8005,N_9005);
nor U11723 (N_11723,N_8828,N_8076);
xnor U11724 (N_11724,N_9178,N_8396);
nor U11725 (N_11725,N_9415,N_9628);
nand U11726 (N_11726,N_9289,N_8592);
or U11727 (N_11727,N_9414,N_8140);
xor U11728 (N_11728,N_8651,N_9553);
or U11729 (N_11729,N_8329,N_9220);
and U11730 (N_11730,N_8488,N_9062);
xor U11731 (N_11731,N_9764,N_8672);
nor U11732 (N_11732,N_8979,N_9882);
and U11733 (N_11733,N_8823,N_8381);
or U11734 (N_11734,N_8672,N_8985);
nand U11735 (N_11735,N_8677,N_9876);
or U11736 (N_11736,N_8721,N_9422);
nor U11737 (N_11737,N_9411,N_8588);
nand U11738 (N_11738,N_8189,N_8670);
and U11739 (N_11739,N_9656,N_8432);
or U11740 (N_11740,N_8554,N_9680);
or U11741 (N_11741,N_9035,N_9869);
xor U11742 (N_11742,N_8766,N_9035);
xor U11743 (N_11743,N_8771,N_9887);
or U11744 (N_11744,N_9664,N_8203);
nor U11745 (N_11745,N_9341,N_8695);
nor U11746 (N_11746,N_9744,N_9230);
nor U11747 (N_11747,N_8735,N_9807);
or U11748 (N_11748,N_9879,N_8478);
nor U11749 (N_11749,N_8977,N_9629);
or U11750 (N_11750,N_8091,N_8306);
nor U11751 (N_11751,N_9509,N_8496);
or U11752 (N_11752,N_8308,N_9531);
or U11753 (N_11753,N_8627,N_8839);
xnor U11754 (N_11754,N_9323,N_8699);
or U11755 (N_11755,N_8493,N_9402);
or U11756 (N_11756,N_8638,N_8908);
or U11757 (N_11757,N_8102,N_8549);
xor U11758 (N_11758,N_9680,N_9402);
or U11759 (N_11759,N_9163,N_8981);
nand U11760 (N_11760,N_9123,N_8885);
or U11761 (N_11761,N_9160,N_9110);
and U11762 (N_11762,N_8038,N_8678);
or U11763 (N_11763,N_8263,N_8127);
and U11764 (N_11764,N_9949,N_8405);
nand U11765 (N_11765,N_9250,N_8064);
xor U11766 (N_11766,N_9536,N_8881);
or U11767 (N_11767,N_8910,N_8760);
nor U11768 (N_11768,N_8102,N_8985);
nor U11769 (N_11769,N_9480,N_8747);
and U11770 (N_11770,N_9664,N_8274);
nand U11771 (N_11771,N_9182,N_8821);
xor U11772 (N_11772,N_9011,N_8933);
nand U11773 (N_11773,N_8615,N_9934);
nand U11774 (N_11774,N_9070,N_8673);
or U11775 (N_11775,N_8855,N_9793);
nand U11776 (N_11776,N_9728,N_8366);
xnor U11777 (N_11777,N_9256,N_8720);
nand U11778 (N_11778,N_8728,N_8325);
xnor U11779 (N_11779,N_9767,N_9775);
or U11780 (N_11780,N_8084,N_9757);
and U11781 (N_11781,N_9172,N_9971);
and U11782 (N_11782,N_8051,N_8235);
or U11783 (N_11783,N_9253,N_8034);
or U11784 (N_11784,N_9666,N_9430);
and U11785 (N_11785,N_8125,N_9629);
or U11786 (N_11786,N_9699,N_8308);
nand U11787 (N_11787,N_9552,N_8847);
or U11788 (N_11788,N_9882,N_9754);
and U11789 (N_11789,N_8762,N_9168);
or U11790 (N_11790,N_9404,N_8040);
nand U11791 (N_11791,N_8004,N_8153);
nand U11792 (N_11792,N_9175,N_9595);
nor U11793 (N_11793,N_8246,N_9488);
nor U11794 (N_11794,N_9951,N_9703);
and U11795 (N_11795,N_8689,N_8255);
or U11796 (N_11796,N_8088,N_8989);
and U11797 (N_11797,N_8764,N_8544);
xor U11798 (N_11798,N_8985,N_8000);
nand U11799 (N_11799,N_8397,N_9436);
and U11800 (N_11800,N_8933,N_8385);
or U11801 (N_11801,N_9257,N_9050);
nand U11802 (N_11802,N_8699,N_8247);
nor U11803 (N_11803,N_9071,N_8050);
nand U11804 (N_11804,N_8240,N_8297);
and U11805 (N_11805,N_9801,N_8571);
xor U11806 (N_11806,N_8839,N_9295);
xnor U11807 (N_11807,N_9876,N_8214);
xnor U11808 (N_11808,N_9295,N_8348);
and U11809 (N_11809,N_9524,N_9561);
nor U11810 (N_11810,N_9771,N_9598);
and U11811 (N_11811,N_9575,N_8324);
nand U11812 (N_11812,N_9049,N_9280);
or U11813 (N_11813,N_8433,N_9201);
nor U11814 (N_11814,N_9773,N_9981);
nor U11815 (N_11815,N_8444,N_8881);
nand U11816 (N_11816,N_9741,N_8193);
nand U11817 (N_11817,N_9532,N_9634);
nand U11818 (N_11818,N_8295,N_9757);
nand U11819 (N_11819,N_8724,N_9201);
or U11820 (N_11820,N_8043,N_8327);
nor U11821 (N_11821,N_9476,N_8690);
nor U11822 (N_11822,N_9860,N_9718);
or U11823 (N_11823,N_9948,N_8869);
nand U11824 (N_11824,N_8468,N_9734);
nand U11825 (N_11825,N_8123,N_8794);
or U11826 (N_11826,N_9489,N_8561);
and U11827 (N_11827,N_8426,N_8031);
nor U11828 (N_11828,N_9812,N_9462);
nand U11829 (N_11829,N_9489,N_9658);
nor U11830 (N_11830,N_9964,N_9685);
nand U11831 (N_11831,N_8032,N_8295);
or U11832 (N_11832,N_9537,N_8151);
nand U11833 (N_11833,N_8075,N_8631);
and U11834 (N_11834,N_8262,N_9704);
and U11835 (N_11835,N_9197,N_9059);
nand U11836 (N_11836,N_9332,N_9256);
xor U11837 (N_11837,N_8214,N_8263);
nor U11838 (N_11838,N_9134,N_9051);
nand U11839 (N_11839,N_9462,N_8604);
xnor U11840 (N_11840,N_8747,N_9172);
nand U11841 (N_11841,N_8919,N_8246);
nor U11842 (N_11842,N_8609,N_9164);
or U11843 (N_11843,N_8111,N_9564);
nand U11844 (N_11844,N_8764,N_9754);
nor U11845 (N_11845,N_9305,N_9998);
xor U11846 (N_11846,N_8330,N_8348);
xor U11847 (N_11847,N_9567,N_8141);
nor U11848 (N_11848,N_8194,N_9680);
or U11849 (N_11849,N_9454,N_9963);
and U11850 (N_11850,N_8797,N_8699);
nand U11851 (N_11851,N_8734,N_9076);
or U11852 (N_11852,N_9612,N_8643);
and U11853 (N_11853,N_8908,N_8038);
nand U11854 (N_11854,N_8757,N_8948);
or U11855 (N_11855,N_9638,N_8309);
or U11856 (N_11856,N_9236,N_8491);
xnor U11857 (N_11857,N_9268,N_9484);
and U11858 (N_11858,N_8811,N_9629);
or U11859 (N_11859,N_8986,N_8049);
and U11860 (N_11860,N_9137,N_8916);
or U11861 (N_11861,N_9027,N_8268);
and U11862 (N_11862,N_9231,N_9332);
and U11863 (N_11863,N_9321,N_9931);
nand U11864 (N_11864,N_9801,N_8501);
nor U11865 (N_11865,N_8852,N_9442);
xor U11866 (N_11866,N_8293,N_9233);
nand U11867 (N_11867,N_9469,N_9231);
nand U11868 (N_11868,N_9124,N_9725);
nor U11869 (N_11869,N_9229,N_9680);
nand U11870 (N_11870,N_9759,N_8652);
nand U11871 (N_11871,N_8867,N_8186);
nand U11872 (N_11872,N_9577,N_9131);
xor U11873 (N_11873,N_8439,N_9619);
or U11874 (N_11874,N_8753,N_8736);
or U11875 (N_11875,N_8913,N_8371);
or U11876 (N_11876,N_8878,N_9136);
nor U11877 (N_11877,N_9091,N_8182);
xor U11878 (N_11878,N_8556,N_9645);
nand U11879 (N_11879,N_8746,N_9279);
xor U11880 (N_11880,N_9955,N_8001);
and U11881 (N_11881,N_9728,N_8846);
xnor U11882 (N_11882,N_9805,N_9415);
and U11883 (N_11883,N_9856,N_9895);
or U11884 (N_11884,N_8673,N_8358);
xor U11885 (N_11885,N_8425,N_8363);
xor U11886 (N_11886,N_9955,N_9571);
nor U11887 (N_11887,N_8071,N_9387);
and U11888 (N_11888,N_9413,N_9100);
and U11889 (N_11889,N_8004,N_9354);
nand U11890 (N_11890,N_8944,N_9067);
and U11891 (N_11891,N_9637,N_9912);
nor U11892 (N_11892,N_9510,N_9813);
xor U11893 (N_11893,N_8517,N_9258);
or U11894 (N_11894,N_8822,N_9032);
nand U11895 (N_11895,N_9396,N_9742);
or U11896 (N_11896,N_9362,N_8119);
or U11897 (N_11897,N_9273,N_8083);
or U11898 (N_11898,N_8150,N_9953);
nand U11899 (N_11899,N_9834,N_9556);
or U11900 (N_11900,N_8737,N_9166);
and U11901 (N_11901,N_9817,N_9978);
or U11902 (N_11902,N_9285,N_9818);
or U11903 (N_11903,N_8760,N_8804);
nor U11904 (N_11904,N_9419,N_8147);
nand U11905 (N_11905,N_9206,N_9148);
nor U11906 (N_11906,N_8124,N_8667);
and U11907 (N_11907,N_9196,N_8398);
nor U11908 (N_11908,N_8147,N_8061);
nor U11909 (N_11909,N_9596,N_9305);
or U11910 (N_11910,N_9639,N_8024);
or U11911 (N_11911,N_9672,N_9665);
and U11912 (N_11912,N_9801,N_8318);
nand U11913 (N_11913,N_8515,N_9420);
and U11914 (N_11914,N_9546,N_9364);
xnor U11915 (N_11915,N_8364,N_9725);
and U11916 (N_11916,N_8039,N_8574);
and U11917 (N_11917,N_9276,N_8583);
and U11918 (N_11918,N_9600,N_9599);
nor U11919 (N_11919,N_9764,N_8471);
and U11920 (N_11920,N_8072,N_9818);
nor U11921 (N_11921,N_8332,N_9451);
nand U11922 (N_11922,N_9073,N_9146);
or U11923 (N_11923,N_9467,N_9406);
and U11924 (N_11924,N_9547,N_8767);
or U11925 (N_11925,N_9328,N_9025);
and U11926 (N_11926,N_9637,N_9021);
nor U11927 (N_11927,N_9681,N_8487);
xnor U11928 (N_11928,N_8323,N_8865);
and U11929 (N_11929,N_9192,N_8370);
xnor U11930 (N_11930,N_9559,N_8033);
or U11931 (N_11931,N_8592,N_9858);
nor U11932 (N_11932,N_9260,N_8949);
nor U11933 (N_11933,N_9092,N_8044);
nand U11934 (N_11934,N_8623,N_9177);
xnor U11935 (N_11935,N_8698,N_9725);
xor U11936 (N_11936,N_9377,N_9034);
xnor U11937 (N_11937,N_9288,N_8326);
and U11938 (N_11938,N_9116,N_9371);
nor U11939 (N_11939,N_8265,N_9747);
and U11940 (N_11940,N_8044,N_8866);
and U11941 (N_11941,N_8244,N_9579);
or U11942 (N_11942,N_8092,N_8125);
nor U11943 (N_11943,N_9129,N_9507);
xor U11944 (N_11944,N_9569,N_8221);
xnor U11945 (N_11945,N_8944,N_8616);
xnor U11946 (N_11946,N_8746,N_9230);
nand U11947 (N_11947,N_8841,N_8562);
and U11948 (N_11948,N_8756,N_9772);
xnor U11949 (N_11949,N_9657,N_9945);
or U11950 (N_11950,N_8218,N_8051);
xnor U11951 (N_11951,N_8952,N_9306);
and U11952 (N_11952,N_8775,N_8971);
and U11953 (N_11953,N_8635,N_8328);
nor U11954 (N_11954,N_9881,N_8408);
or U11955 (N_11955,N_8185,N_8051);
or U11956 (N_11956,N_8434,N_9070);
xor U11957 (N_11957,N_8576,N_8880);
nand U11958 (N_11958,N_9783,N_9782);
nand U11959 (N_11959,N_9760,N_9318);
nand U11960 (N_11960,N_8282,N_9468);
or U11961 (N_11961,N_9035,N_8999);
or U11962 (N_11962,N_9281,N_8130);
nor U11963 (N_11963,N_8659,N_8213);
nor U11964 (N_11964,N_8271,N_9827);
and U11965 (N_11965,N_9889,N_8676);
nor U11966 (N_11966,N_9134,N_9823);
nor U11967 (N_11967,N_8445,N_8958);
and U11968 (N_11968,N_9035,N_9036);
nand U11969 (N_11969,N_8587,N_8634);
xnor U11970 (N_11970,N_9360,N_9770);
nor U11971 (N_11971,N_8445,N_9925);
nand U11972 (N_11972,N_9699,N_8886);
nand U11973 (N_11973,N_9037,N_9223);
xnor U11974 (N_11974,N_8998,N_9279);
or U11975 (N_11975,N_8091,N_9073);
nor U11976 (N_11976,N_8269,N_8932);
nand U11977 (N_11977,N_8714,N_8300);
nand U11978 (N_11978,N_8911,N_9714);
xnor U11979 (N_11979,N_9380,N_9799);
nand U11980 (N_11980,N_9085,N_9026);
nand U11981 (N_11981,N_9200,N_8560);
and U11982 (N_11982,N_8493,N_8723);
xnor U11983 (N_11983,N_9250,N_8526);
and U11984 (N_11984,N_9622,N_8392);
and U11985 (N_11985,N_8344,N_8756);
and U11986 (N_11986,N_9848,N_9376);
nand U11987 (N_11987,N_9226,N_8856);
xnor U11988 (N_11988,N_8302,N_9402);
xnor U11989 (N_11989,N_8481,N_8424);
nand U11990 (N_11990,N_8473,N_8214);
nor U11991 (N_11991,N_8496,N_9334);
xor U11992 (N_11992,N_8388,N_9570);
nor U11993 (N_11993,N_8607,N_9589);
or U11994 (N_11994,N_9317,N_8385);
nand U11995 (N_11995,N_8957,N_9135);
and U11996 (N_11996,N_9925,N_8544);
nand U11997 (N_11997,N_9480,N_9998);
or U11998 (N_11998,N_9390,N_9088);
or U11999 (N_11999,N_9733,N_8497);
or U12000 (N_12000,N_10166,N_10141);
nor U12001 (N_12001,N_10011,N_10394);
and U12002 (N_12002,N_11055,N_10750);
and U12003 (N_12003,N_11825,N_10013);
xnor U12004 (N_12004,N_10960,N_11320);
nand U12005 (N_12005,N_11927,N_11839);
xor U12006 (N_12006,N_11246,N_10824);
nand U12007 (N_12007,N_11326,N_10036);
nand U12008 (N_12008,N_11422,N_10583);
xnor U12009 (N_12009,N_10457,N_11955);
nand U12010 (N_12010,N_11756,N_11216);
nor U12011 (N_12011,N_11318,N_10804);
or U12012 (N_12012,N_10536,N_10444);
and U12013 (N_12013,N_11574,N_10061);
xor U12014 (N_12014,N_10834,N_11810);
nor U12015 (N_12015,N_10529,N_11153);
nand U12016 (N_12016,N_10606,N_10274);
xor U12017 (N_12017,N_11190,N_11709);
and U12018 (N_12018,N_11462,N_11308);
xor U12019 (N_12019,N_11464,N_11553);
xor U12020 (N_12020,N_10706,N_11288);
or U12021 (N_12021,N_10389,N_11355);
nand U12022 (N_12022,N_11097,N_10110);
and U12023 (N_12023,N_11297,N_10962);
nor U12024 (N_12024,N_11032,N_10652);
xor U12025 (N_12025,N_10910,N_10755);
nand U12026 (N_12026,N_11831,N_10589);
nand U12027 (N_12027,N_11440,N_11775);
and U12028 (N_12028,N_10168,N_10470);
nand U12029 (N_12029,N_11439,N_11542);
and U12030 (N_12030,N_11799,N_10841);
nor U12031 (N_12031,N_10702,N_11105);
or U12032 (N_12032,N_10932,N_11127);
or U12033 (N_12033,N_11473,N_11581);
or U12034 (N_12034,N_10655,N_10335);
nand U12035 (N_12035,N_10758,N_11836);
and U12036 (N_12036,N_10759,N_11585);
xor U12037 (N_12037,N_11084,N_10486);
nand U12038 (N_12038,N_10762,N_10008);
and U12039 (N_12039,N_10934,N_10359);
xor U12040 (N_12040,N_10403,N_10154);
xnor U12041 (N_12041,N_10845,N_11205);
nor U12042 (N_12042,N_11466,N_10975);
or U12043 (N_12043,N_10734,N_10575);
or U12044 (N_12044,N_11313,N_11513);
nand U12045 (N_12045,N_11787,N_11652);
nor U12046 (N_12046,N_11527,N_10404);
and U12047 (N_12047,N_11414,N_10580);
or U12048 (N_12048,N_11434,N_11941);
nand U12049 (N_12049,N_10891,N_10030);
nand U12050 (N_12050,N_10653,N_10305);
nand U12051 (N_12051,N_10139,N_10007);
nor U12052 (N_12052,N_10095,N_10948);
nor U12053 (N_12053,N_11432,N_11938);
nor U12054 (N_12054,N_11474,N_10693);
nand U12055 (N_12055,N_11532,N_11807);
nand U12056 (N_12056,N_11199,N_10374);
xor U12057 (N_12057,N_10566,N_10542);
xor U12058 (N_12058,N_10793,N_10924);
nand U12059 (N_12059,N_11011,N_10640);
nand U12060 (N_12060,N_10654,N_10667);
xnor U12061 (N_12061,N_11536,N_11183);
nor U12062 (N_12062,N_10393,N_10809);
or U12063 (N_12063,N_11106,N_10108);
or U12064 (N_12064,N_10093,N_11041);
or U12065 (N_12065,N_10228,N_11817);
nor U12066 (N_12066,N_10282,N_11167);
nand U12067 (N_12067,N_11904,N_11385);
nand U12068 (N_12068,N_11537,N_11811);
and U12069 (N_12069,N_10626,N_11509);
nor U12070 (N_12070,N_10921,N_11266);
xnor U12071 (N_12071,N_10749,N_11400);
nor U12072 (N_12072,N_11263,N_10101);
nand U12073 (N_12073,N_11600,N_11991);
and U12074 (N_12074,N_11114,N_10747);
nor U12075 (N_12075,N_11983,N_11144);
and U12076 (N_12076,N_11822,N_10897);
and U12077 (N_12077,N_10195,N_10516);
nand U12078 (N_12078,N_10153,N_10767);
nand U12079 (N_12079,N_10491,N_11323);
nand U12080 (N_12080,N_10796,N_10662);
and U12081 (N_12081,N_11777,N_11576);
nand U12082 (N_12082,N_10300,N_10303);
nand U12083 (N_12083,N_11354,N_10576);
and U12084 (N_12084,N_10885,N_10386);
xor U12085 (N_12085,N_11182,N_11245);
and U12086 (N_12086,N_10893,N_10694);
nor U12087 (N_12087,N_10387,N_11281);
xor U12088 (N_12088,N_11240,N_10106);
xnor U12089 (N_12089,N_11875,N_10937);
xnor U12090 (N_12090,N_10976,N_11175);
and U12091 (N_12091,N_10596,N_11830);
and U12092 (N_12092,N_11868,N_11025);
xor U12093 (N_12093,N_10760,N_11088);
or U12094 (N_12094,N_11430,N_10043);
and U12095 (N_12095,N_11671,N_11007);
xor U12096 (N_12096,N_10239,N_11197);
or U12097 (N_12097,N_11699,N_10617);
nor U12098 (N_12098,N_10521,N_10838);
xnor U12099 (N_12099,N_10026,N_10420);
or U12100 (N_12100,N_11647,N_11277);
nor U12101 (N_12101,N_10898,N_10116);
xnor U12102 (N_12102,N_11715,N_10120);
nand U12103 (N_12103,N_10573,N_11573);
nand U12104 (N_12104,N_10276,N_10244);
nor U12105 (N_12105,N_11828,N_10006);
nor U12106 (N_12106,N_11203,N_11776);
or U12107 (N_12107,N_11195,N_10735);
nand U12108 (N_12108,N_10454,N_11934);
xor U12109 (N_12109,N_11207,N_10205);
and U12110 (N_12110,N_10237,N_10740);
and U12111 (N_12111,N_10671,N_11670);
and U12112 (N_12112,N_11117,N_10524);
xor U12113 (N_12113,N_11595,N_11568);
or U12114 (N_12114,N_10051,N_10741);
nor U12115 (N_12115,N_10969,N_10314);
nand U12116 (N_12116,N_10811,N_11802);
nand U12117 (N_12117,N_11497,N_10795);
nor U12118 (N_12118,N_11310,N_10788);
xnor U12119 (N_12119,N_10649,N_10187);
xor U12120 (N_12120,N_11408,N_10049);
xnor U12121 (N_12121,N_10900,N_11342);
nor U12122 (N_12122,N_10451,N_10504);
nand U12123 (N_12123,N_11001,N_10604);
and U12124 (N_12124,N_11601,N_11036);
and U12125 (N_12125,N_11303,N_11349);
xnor U12126 (N_12126,N_11230,N_10500);
nand U12127 (N_12127,N_10967,N_10324);
nand U12128 (N_12128,N_10193,N_11689);
nand U12129 (N_12129,N_10854,N_11402);
nor U12130 (N_12130,N_11919,N_10831);
nor U12131 (N_12131,N_11760,N_10047);
xnor U12132 (N_12132,N_11631,N_11389);
and U12133 (N_12133,N_10226,N_10764);
and U12134 (N_12134,N_11696,N_11999);
and U12135 (N_12135,N_10126,N_11970);
nand U12136 (N_12136,N_11341,N_10395);
nor U12137 (N_12137,N_11994,N_11339);
or U12138 (N_12138,N_11618,N_10002);
nor U12139 (N_12139,N_11470,N_11102);
nor U12140 (N_12140,N_11192,N_11833);
xor U12141 (N_12141,N_10643,N_10115);
and U12142 (N_12142,N_11805,N_11617);
xor U12143 (N_12143,N_11383,N_10460);
nor U12144 (N_12144,N_11605,N_10235);
nor U12145 (N_12145,N_10316,N_10497);
nand U12146 (N_12146,N_10243,N_10015);
nor U12147 (N_12147,N_11120,N_11265);
xnor U12148 (N_12148,N_10466,N_10376);
and U12149 (N_12149,N_11923,N_11176);
and U12150 (N_12150,N_11596,N_10288);
nand U12151 (N_12151,N_11003,N_10123);
nand U12152 (N_12152,N_11899,N_10950);
nor U12153 (N_12153,N_11249,N_10603);
nor U12154 (N_12154,N_11543,N_11364);
or U12155 (N_12155,N_11482,N_11993);
and U12156 (N_12156,N_11194,N_11594);
nor U12157 (N_12157,N_11356,N_11572);
nor U12158 (N_12158,N_10790,N_10806);
or U12159 (N_12159,N_10940,N_10328);
nand U12160 (N_12160,N_11334,N_11714);
nand U12161 (N_12161,N_10301,N_10971);
nand U12162 (N_12162,N_10505,N_10582);
nand U12163 (N_12163,N_10961,N_11332);
and U12164 (N_12164,N_11759,N_10634);
nand U12165 (N_12165,N_10939,N_10369);
nor U12166 (N_12166,N_10904,N_10765);
xnor U12167 (N_12167,N_11163,N_10778);
xnor U12168 (N_12168,N_10943,N_10579);
nand U12169 (N_12169,N_11673,N_11258);
and U12170 (N_12170,N_11020,N_11599);
xor U12171 (N_12171,N_10996,N_11271);
xor U12172 (N_12172,N_10528,N_11902);
nand U12173 (N_12173,N_11534,N_11159);
xnor U12174 (N_12174,N_10771,N_10068);
nor U12175 (N_12175,N_11896,N_11416);
and U12176 (N_12176,N_10103,N_10434);
or U12177 (N_12177,N_11152,N_11417);
nand U12178 (N_12178,N_11038,N_11446);
nand U12179 (N_12179,N_11523,N_11247);
or U12180 (N_12180,N_11401,N_11141);
xor U12181 (N_12181,N_10357,N_10842);
or U12182 (N_12182,N_11680,N_11161);
and U12183 (N_12183,N_10232,N_11888);
nand U12184 (N_12184,N_10724,N_11920);
nor U12185 (N_12185,N_11312,N_11498);
xnor U12186 (N_12186,N_11067,N_10159);
xor U12187 (N_12187,N_10056,N_11837);
or U12188 (N_12188,N_10787,N_10089);
xnor U12189 (N_12189,N_10614,N_10913);
nand U12190 (N_12190,N_11877,N_10259);
and U12191 (N_12191,N_11338,N_11615);
and U12192 (N_12192,N_10517,N_10443);
or U12193 (N_12193,N_11373,N_11587);
nor U12194 (N_12194,N_11008,N_11283);
xor U12195 (N_12195,N_11517,N_11979);
nand U12196 (N_12196,N_11257,N_10400);
nand U12197 (N_12197,N_10630,N_10099);
xor U12198 (N_12198,N_10507,N_11094);
nand U12199 (N_12199,N_10745,N_11031);
and U12200 (N_12200,N_10894,N_11765);
and U12201 (N_12201,N_11487,N_10202);
or U12202 (N_12202,N_11704,N_11525);
or U12203 (N_12203,N_10287,N_10465);
xnor U12204 (N_12204,N_10025,N_11835);
or U12205 (N_12205,N_11891,N_10856);
or U12206 (N_12206,N_10931,N_10463);
xnor U12207 (N_12207,N_10121,N_11445);
and U12208 (N_12208,N_10769,N_10612);
nor U12209 (N_12209,N_10479,N_10508);
nand U12210 (N_12210,N_11869,N_10742);
and U12211 (N_12211,N_11851,N_10902);
and U12212 (N_12212,N_10797,N_10585);
nand U12213 (N_12213,N_10746,N_11588);
nand U12214 (N_12214,N_10339,N_11597);
xor U12215 (N_12215,N_10514,N_10416);
xnor U12216 (N_12216,N_11479,N_11713);
and U12217 (N_12217,N_10544,N_10726);
xnor U12218 (N_12218,N_11329,N_11638);
or U12219 (N_12219,N_10737,N_11989);
nor U12220 (N_12220,N_10307,N_10494);
or U12221 (N_12221,N_10225,N_10851);
or U12222 (N_12222,N_11060,N_11206);
nor U12223 (N_12223,N_10993,N_11812);
and U12224 (N_12224,N_11790,N_10447);
xnor U12225 (N_12225,N_11004,N_11437);
or U12226 (N_12226,N_10016,N_10175);
nor U12227 (N_12227,N_11550,N_11253);
xnor U12228 (N_12228,N_10965,N_11508);
nand U12229 (N_12229,N_10938,N_10496);
nand U12230 (N_12230,N_11900,N_11380);
xor U12231 (N_12231,N_11040,N_11413);
nor U12232 (N_12232,N_10846,N_11959);
nand U12233 (N_12233,N_11580,N_11629);
nand U12234 (N_12234,N_10130,N_11619);
nand U12235 (N_12235,N_10651,N_10406);
nand U12236 (N_12236,N_10538,N_10555);
and U12237 (N_12237,N_11026,N_11926);
nand U12238 (N_12238,N_10919,N_10128);
and U12239 (N_12239,N_11614,N_11411);
nand U12240 (N_12240,N_11065,N_11975);
and U12241 (N_12241,N_11908,N_10313);
xnor U12242 (N_12242,N_10293,N_10147);
xnor U12243 (N_12243,N_10333,N_10431);
nand U12244 (N_12244,N_11823,N_10722);
or U12245 (N_12245,N_10928,N_10010);
and U12246 (N_12246,N_10032,N_11488);
nand U12247 (N_12247,N_11085,N_10060);
nor U12248 (N_12248,N_11820,N_11870);
or U12249 (N_12249,N_10438,N_11274);
or U12250 (N_12250,N_10058,N_11819);
nand U12251 (N_12251,N_11030,N_10363);
nor U12252 (N_12252,N_11808,N_11235);
xnor U12253 (N_12253,N_11366,N_11078);
or U12254 (N_12254,N_11645,N_10432);
and U12255 (N_12255,N_11973,N_10294);
nand U12256 (N_12256,N_11186,N_10714);
xor U12257 (N_12257,N_10292,N_10349);
nor U12258 (N_12258,N_10268,N_10847);
nor U12259 (N_12259,N_10968,N_11307);
xor U12260 (N_12260,N_10623,N_11495);
and U12261 (N_12261,N_11452,N_10245);
and U12262 (N_12262,N_11984,N_10484);
and U12263 (N_12263,N_10161,N_10481);
xnor U12264 (N_12264,N_10345,N_11855);
xor U12265 (N_12265,N_10568,N_10889);
xor U12266 (N_12266,N_10914,N_10413);
xor U12267 (N_12267,N_11276,N_10468);
xnor U12268 (N_12268,N_10241,N_10152);
xor U12269 (N_12269,N_10028,N_10029);
nor U12270 (N_12270,N_10005,N_10658);
or U12271 (N_12271,N_11000,N_11363);
or U12272 (N_12272,N_11490,N_10590);
nor U12273 (N_12273,N_10880,N_11173);
and U12274 (N_12274,N_10318,N_11267);
xor U12275 (N_12275,N_10285,N_10201);
or U12276 (N_12276,N_11539,N_11353);
nor U12277 (N_12277,N_10077,N_11949);
nand U12278 (N_12278,N_11304,N_10577);
xor U12279 (N_12279,N_11145,N_11123);
and U12280 (N_12280,N_11384,N_11890);
nor U12281 (N_12281,N_11922,N_11579);
nor U12282 (N_12282,N_10901,N_10743);
xor U12283 (N_12283,N_10183,N_10180);
or U12284 (N_12284,N_10203,N_11796);
or U12285 (N_12285,N_10422,N_10559);
and U12286 (N_12286,N_11268,N_10926);
nor U12287 (N_12287,N_11282,N_10320);
and U12288 (N_12288,N_11551,N_11138);
and U12289 (N_12289,N_11419,N_11940);
xnor U12290 (N_12290,N_11119,N_10732);
xnor U12291 (N_12291,N_10124,N_11672);
or U12292 (N_12292,N_11345,N_11763);
or U12293 (N_12293,N_11767,N_10679);
and U12294 (N_12294,N_11842,N_10753);
xnor U12295 (N_12295,N_10189,N_10805);
nor U12296 (N_12296,N_11412,N_10137);
xnor U12297 (N_12297,N_11590,N_11985);
xor U12298 (N_12298,N_11129,N_11586);
and U12299 (N_12299,N_10877,N_11511);
or U12300 (N_12300,N_11604,N_11967);
nor U12301 (N_12301,N_10208,N_11721);
and U12302 (N_12302,N_10905,N_11952);
or U12303 (N_12303,N_10263,N_10781);
xor U12304 (N_12304,N_11476,N_10022);
or U12305 (N_12305,N_11570,N_10859);
nand U12306 (N_12306,N_10867,N_10079);
or U12307 (N_12307,N_11730,N_10808);
or U12308 (N_12308,N_11174,N_10362);
or U12309 (N_12309,N_10234,N_10227);
xnor U12310 (N_12310,N_11861,N_11644);
nor U12311 (N_12311,N_11557,N_10719);
or U12312 (N_12312,N_11793,N_10262);
or U12313 (N_12313,N_10117,N_10267);
or U12314 (N_12314,N_10858,N_11727);
nand U12315 (N_12315,N_10511,N_10534);
xnor U12316 (N_12316,N_11058,N_11204);
or U12317 (N_12317,N_11901,N_11944);
nor U12318 (N_12318,N_11359,N_11347);
xnor U12319 (N_12319,N_10372,N_11331);
nand U12320 (N_12320,N_10250,N_10249);
nand U12321 (N_12321,N_11724,N_11181);
xor U12322 (N_12322,N_11782,N_10170);
and U12323 (N_12323,N_11212,N_11228);
or U12324 (N_12324,N_10629,N_11740);
xor U12325 (N_12325,N_11781,N_11471);
or U12326 (N_12326,N_10866,N_10642);
nor U12327 (N_12327,N_11660,N_11154);
and U12328 (N_12328,N_11054,N_10140);
nand U12329 (N_12329,N_10081,N_10983);
and U12330 (N_12330,N_11280,N_10260);
nand U12331 (N_12331,N_10855,N_10247);
nand U12332 (N_12332,N_11410,N_11530);
xor U12333 (N_12333,N_11602,N_11243);
or U12334 (N_12334,N_10622,N_10423);
nand U12335 (N_12335,N_10472,N_10306);
nand U12336 (N_12336,N_11333,N_10001);
and U12337 (N_12337,N_10739,N_10777);
or U12338 (N_12338,N_10186,N_10090);
or U12339 (N_12339,N_10863,N_11438);
xnor U12340 (N_12340,N_11700,N_11388);
xor U12341 (N_12341,N_10815,N_10144);
xor U12342 (N_12342,N_11939,N_11749);
nor U12343 (N_12343,N_10836,N_10609);
nor U12344 (N_12344,N_11424,N_10238);
nand U12345 (N_12345,N_11758,N_11296);
nor U12346 (N_12346,N_11079,N_10399);
xor U12347 (N_12347,N_11703,N_10696);
nand U12348 (N_12348,N_11361,N_11914);
nand U12349 (N_12349,N_11104,N_10476);
nor U12350 (N_12350,N_10122,N_11878);
nand U12351 (N_12351,N_11957,N_10150);
nor U12352 (N_12352,N_10543,N_10532);
nor U12353 (N_12353,N_11061,N_10118);
or U12354 (N_12354,N_10903,N_10502);
xor U12355 (N_12355,N_11905,N_10289);
nand U12356 (N_12356,N_11491,N_11012);
nand U12357 (N_12357,N_11744,N_10136);
xnor U12358 (N_12358,N_11829,N_11290);
and U12359 (N_12359,N_10786,N_11126);
and U12360 (N_12360,N_11502,N_11451);
xor U12361 (N_12361,N_11856,N_11221);
and U12362 (N_12362,N_10888,N_10673);
nor U12363 (N_12363,N_11695,N_10218);
and U12364 (N_12364,N_10455,N_11978);
xnor U12365 (N_12365,N_10733,N_11177);
or U12366 (N_12366,N_10211,N_10572);
nand U12367 (N_12367,N_10074,N_10995);
and U12368 (N_12368,N_10265,N_10003);
or U12369 (N_12369,N_10474,N_11386);
nor U12370 (N_12370,N_11073,N_11954);
xnor U12371 (N_12371,N_10094,N_11664);
and U12372 (N_12372,N_11217,N_10627);
and U12373 (N_12373,N_11809,N_11208);
nor U12374 (N_12374,N_10207,N_11883);
and U12375 (N_12375,N_11658,N_10471);
xnor U12376 (N_12376,N_10200,N_10309);
nand U12377 (N_12377,N_11946,N_11650);
or U12378 (N_12378,N_11780,N_10537);
nor U12379 (N_12379,N_11365,N_11494);
or U12380 (N_12380,N_11379,N_10927);
or U12381 (N_12381,N_11876,N_11128);
nor U12382 (N_12382,N_10224,N_10744);
nor U12383 (N_12383,N_11444,N_11679);
nor U12384 (N_12384,N_11591,N_10196);
or U12385 (N_12385,N_10701,N_11107);
xor U12386 (N_12386,N_10246,N_10280);
nand U12387 (N_12387,N_10584,N_11395);
nor U12388 (N_12388,N_11251,N_11771);
and U12389 (N_12389,N_10433,N_10929);
nand U12390 (N_12390,N_11571,N_11215);
and U12391 (N_12391,N_10972,N_10730);
nor U12392 (N_12392,N_11248,N_10176);
nand U12393 (N_12393,N_10252,N_10379);
nand U12394 (N_12394,N_11858,N_10217);
xnor U12395 (N_12395,N_11827,N_10270);
nor U12396 (N_12396,N_10297,N_11643);
nand U12397 (N_12397,N_10984,N_10639);
or U12398 (N_12398,N_11512,N_11610);
nor U12399 (N_12399,N_10558,N_11209);
and U12400 (N_12400,N_11783,N_11314);
and U12401 (N_12401,N_10601,N_11840);
nand U12402 (N_12402,N_10849,N_11706);
and U12403 (N_12403,N_11879,N_10105);
nand U12404 (N_12404,N_11800,N_10873);
and U12405 (N_12405,N_10564,N_11506);
nor U12406 (N_12406,N_10182,N_10830);
nand U12407 (N_12407,N_11168,N_10633);
xnor U12408 (N_12408,N_10650,N_11640);
and U12409 (N_12409,N_10419,N_10160);
and U12410 (N_12410,N_10553,N_10367);
xnor U12411 (N_12411,N_10213,N_10146);
nand U12412 (N_12412,N_11428,N_10353);
xor U12413 (N_12413,N_11351,N_11301);
or U12414 (N_12414,N_11447,N_10704);
and U12415 (N_12415,N_11484,N_10409);
and U12416 (N_12416,N_11567,N_10779);
nand U12417 (N_12417,N_10813,N_10381);
and U12418 (N_12418,N_10659,N_10084);
nor U12419 (N_12419,N_11801,N_11300);
xnor U12420 (N_12420,N_10024,N_11261);
and U12421 (N_12421,N_11387,N_11130);
or U12422 (N_12422,N_10608,N_11225);
and U12423 (N_12423,N_11016,N_11298);
nand U12424 (N_12424,N_11892,N_10665);
or U12425 (N_12425,N_10113,N_10329);
nor U12426 (N_12426,N_10242,N_10989);
nor U12427 (N_12427,N_10518,N_10034);
nand U12428 (N_12428,N_10019,N_10944);
nand U12429 (N_12429,N_10802,N_10946);
nor U12430 (N_12430,N_11913,N_11232);
nand U12431 (N_12431,N_10982,N_10377);
and U12432 (N_12432,N_11947,N_11371);
or U12433 (N_12433,N_11370,N_11755);
or U12434 (N_12434,N_10776,N_10539);
or U12435 (N_12435,N_11798,N_11327);
or U12436 (N_12436,N_10883,N_10269);
and U12437 (N_12437,N_10865,N_10214);
and U12438 (N_12438,N_10695,N_10828);
nor U12439 (N_12439,N_10046,N_11467);
and U12440 (N_12440,N_10461,N_10258);
or U12441 (N_12441,N_10050,N_10446);
or U12442 (N_12442,N_10857,N_10216);
xor U12443 (N_12443,N_11394,N_10499);
xnor U12444 (N_12444,N_11937,N_11986);
and U12445 (N_12445,N_10647,N_11753);
xor U12446 (N_12446,N_10040,N_11961);
nor U12447 (N_12447,N_10772,N_10418);
or U12448 (N_12448,N_10261,N_11035);
nand U12449 (N_12449,N_11843,N_11171);
or U12450 (N_12450,N_11239,N_11918);
nand U12451 (N_12451,N_11712,N_10009);
or U12452 (N_12452,N_10998,N_10916);
and U12453 (N_12453,N_10325,N_10266);
nand U12454 (N_12454,N_11360,N_11734);
nand U12455 (N_12455,N_10941,N_11874);
nand U12456 (N_12456,N_11815,N_10763);
or U12457 (N_12457,N_11732,N_11113);
nand U12458 (N_12458,N_11684,N_10281);
or U12459 (N_12459,N_10680,N_10979);
xor U12460 (N_12460,N_11133,N_11165);
nor U12461 (N_12461,N_11146,N_10057);
or U12462 (N_12462,N_10563,N_10812);
nand U12463 (N_12463,N_10296,N_10512);
and U12464 (N_12464,N_10490,N_10892);
xnor U12465 (N_12465,N_11273,N_10371);
or U12466 (N_12466,N_10284,N_11982);
nor U12467 (N_12467,N_11059,N_10337);
xor U12468 (N_12468,N_10908,N_11050);
xnor U12469 (N_12469,N_10964,N_10798);
xor U12470 (N_12470,N_11864,N_10799);
or U12471 (N_12471,N_10545,N_10299);
and U12472 (N_12472,N_11972,N_10692);
nor U12473 (N_12473,N_11448,N_10663);
or U12474 (N_12474,N_10700,N_11854);
or U12475 (N_12475,N_10233,N_10358);
and U12476 (N_12476,N_11997,N_11393);
or U12477 (N_12477,N_10062,N_11136);
and U12478 (N_12478,N_11784,N_11045);
or U12479 (N_12479,N_11449,N_10560);
and U12480 (N_12480,N_10954,N_10052);
and U12481 (N_12481,N_10145,N_11917);
nand U12482 (N_12482,N_10114,N_10063);
or U12483 (N_12483,N_10638,N_11907);
xnor U12484 (N_12484,N_11708,N_11089);
nor U12485 (N_12485,N_11654,N_11531);
or U12486 (N_12486,N_10999,N_11358);
nor U12487 (N_12487,N_10493,N_11222);
and U12488 (N_12488,N_11124,N_11633);
and U12489 (N_12489,N_10458,N_10185);
and U12490 (N_12490,N_11569,N_10044);
nand U12491 (N_12491,N_10330,N_10864);
nor U12492 (N_12492,N_11951,N_11659);
nor U12493 (N_12493,N_11010,N_10597);
nand U12494 (N_12494,N_11931,N_10223);
and U12495 (N_12495,N_11023,N_10986);
nor U12496 (N_12496,N_10111,N_10748);
nor U12497 (N_12497,N_11849,N_11233);
and U12498 (N_12498,N_11048,N_10801);
nand U12499 (N_12499,N_11287,N_11289);
and U12500 (N_12500,N_10957,N_11226);
nand U12501 (N_12501,N_11071,N_11237);
nand U12502 (N_12502,N_10323,N_11223);
nand U12503 (N_12503,N_10669,N_11733);
or U12504 (N_12504,N_11125,N_10509);
or U12505 (N_12505,N_11948,N_10531);
or U12506 (N_12506,N_11608,N_10738);
or U12507 (N_12507,N_10442,N_10076);
nand U12508 (N_12508,N_10341,N_11200);
xnor U12509 (N_12509,N_11850,N_11737);
nor U12510 (N_12510,N_10038,N_11785);
and U12511 (N_12511,N_11321,N_10412);
and U12512 (N_12512,N_10023,N_10054);
nor U12513 (N_12513,N_10818,N_10966);
nand U12514 (N_12514,N_11166,N_11916);
xnor U12515 (N_12515,N_11966,N_11871);
nand U12516 (N_12516,N_10985,N_10519);
xnor U12517 (N_12517,N_11987,N_11122);
nor U12518 (N_12518,N_10448,N_10810);
or U12519 (N_12519,N_10833,N_11435);
nand U12520 (N_12520,N_11806,N_10478);
nand U12521 (N_12521,N_10310,N_10955);
and U12522 (N_12522,N_10319,N_11076);
and U12523 (N_12523,N_10370,N_10075);
xor U12524 (N_12524,N_10085,N_11172);
xnor U12525 (N_12525,N_10197,N_11803);
nor U12526 (N_12526,N_11528,N_11074);
nand U12527 (N_12527,N_10298,N_11158);
nand U12528 (N_12528,N_10549,N_11728);
nor U12529 (N_12529,N_10548,N_11179);
and U12530 (N_12530,N_11773,N_10872);
or U12531 (N_12531,N_10721,N_11657);
or U12532 (N_12532,N_11853,N_10206);
xnor U12533 (N_12533,N_11865,N_10194);
and U12534 (N_12534,N_10783,N_11091);
nand U12535 (N_12535,N_10578,N_10988);
or U12536 (N_12536,N_11971,N_11838);
and U12537 (N_12537,N_10495,N_11562);
xnor U12538 (N_12538,N_10906,N_10012);
nor U12539 (N_12539,N_11661,N_10248);
and U12540 (N_12540,N_11147,N_11472);
and U12541 (N_12541,N_10594,N_10177);
xnor U12542 (N_12542,N_10621,N_10624);
nor U12543 (N_12543,N_11552,N_11108);
xnor U12544 (N_12544,N_10648,N_11156);
or U12545 (N_12545,N_11750,N_11033);
and U12546 (N_12546,N_11747,N_10593);
and U12547 (N_12547,N_11286,N_11889);
nand U12548 (N_12548,N_11407,N_10396);
or U12549 (N_12549,N_11887,N_11431);
nand U12550 (N_12550,N_11824,N_11350);
or U12551 (N_12551,N_10611,N_10498);
xor U12552 (N_12552,N_10800,N_10978);
or U12553 (N_12553,N_11852,N_10148);
xor U12554 (N_12554,N_10078,N_10354);
nand U12555 (N_12555,N_10343,N_11752);
xnor U12556 (N_12556,N_10426,N_11911);
nor U12557 (N_12557,N_11507,N_11293);
nor U12558 (N_12558,N_10322,N_11455);
and U12559 (N_12559,N_11037,N_11459);
or U12560 (N_12560,N_11157,N_11468);
and U12561 (N_12561,N_11231,N_10550);
nor U12562 (N_12562,N_11390,N_10882);
and U12563 (N_12563,N_11762,N_11169);
or U12564 (N_12564,N_11667,N_10618);
nand U12565 (N_12565,N_11519,N_10109);
xnor U12566 (N_12566,N_10896,N_11882);
nor U12567 (N_12567,N_11284,N_11362);
nand U12568 (N_12568,N_10708,N_11992);
or U12569 (N_12569,N_10766,N_10190);
nand U12570 (N_12570,N_10156,N_11062);
xor U12571 (N_12571,N_11019,N_10429);
nor U12572 (N_12572,N_10331,N_10042);
and U12573 (N_12573,N_11066,N_11518);
nand U12574 (N_12574,N_11956,N_11403);
and U12575 (N_12575,N_10685,N_10164);
xnor U12576 (N_12576,N_10876,N_10761);
nand U12577 (N_12577,N_10482,N_10464);
xnor U12578 (N_12578,N_10340,N_10088);
nand U12579 (N_12579,N_11229,N_10321);
nand U12580 (N_12580,N_11639,N_10586);
and U12581 (N_12581,N_10821,N_10713);
or U12582 (N_12582,N_11315,N_10636);
or U12583 (N_12583,N_10871,N_10411);
or U12584 (N_12584,N_10129,N_11786);
or U12585 (N_12585,N_10449,N_11690);
xor U12586 (N_12586,N_11906,N_11463);
or U12587 (N_12587,N_11184,N_11555);
and U12588 (N_12588,N_11945,N_11486);
nand U12589 (N_12589,N_10687,N_10033);
xor U12590 (N_12590,N_11118,N_10427);
nand U12591 (N_12591,N_11409,N_10417);
and U12592 (N_12592,N_11185,N_11969);
xor U12593 (N_12593,N_10192,N_10501);
and U12594 (N_12594,N_11541,N_11735);
xor U12595 (N_12595,N_10541,N_11404);
nor U12596 (N_12596,N_11558,N_11028);
nand U12597 (N_12597,N_10414,N_11272);
and U12598 (N_12598,N_11236,N_10890);
nor U12599 (N_12599,N_10171,N_11457);
nor U12600 (N_12600,N_11632,N_10958);
or U12601 (N_12601,N_11324,N_10264);
and U12602 (N_12602,N_10041,N_11592);
nor U12603 (N_12603,N_11547,N_11529);
and U12604 (N_12604,N_10131,N_10415);
nor U12605 (N_12605,N_10881,N_10151);
nor U12606 (N_12606,N_11540,N_11860);
nor U12607 (N_12607,N_10690,N_10086);
or U12608 (N_12608,N_10149,N_10535);
nor U12609 (N_12609,N_10717,N_10348);
and U12610 (N_12610,N_11627,N_11336);
nor U12611 (N_12611,N_11425,N_10547);
and U12612 (N_12612,N_11244,N_10308);
or U12613 (N_12613,N_10785,N_11291);
xnor U12614 (N_12614,N_11881,N_10467);
and U12615 (N_12615,N_10645,N_10675);
nor U12616 (N_12616,N_10616,N_10725);
and U12617 (N_12617,N_10691,N_11160);
and U12618 (N_12618,N_10729,N_10751);
or U12619 (N_12619,N_10631,N_10561);
or U12620 (N_12620,N_10104,N_10435);
nor U12621 (N_12621,N_11278,N_11501);
xnor U12622 (N_12622,N_11505,N_10020);
or U12623 (N_12623,N_11420,N_10424);
nand U12624 (N_12624,N_10731,N_10342);
or U12625 (N_12625,N_10421,N_10364);
xnor U12626 (N_12626,N_11250,N_11674);
and U12627 (N_12627,N_11503,N_10789);
nand U12628 (N_12628,N_11087,N_10257);
xnor U12629 (N_12629,N_11396,N_11554);
xnor U12630 (N_12630,N_10922,N_11788);
or U12631 (N_12631,N_10332,N_11832);
and U12632 (N_12632,N_10157,N_11990);
xnor U12633 (N_12633,N_10398,N_11720);
or U12634 (N_12634,N_10951,N_10625);
nor U12635 (N_12635,N_10768,N_10097);
nand U12636 (N_12636,N_11426,N_10683);
or U12637 (N_12637,N_11722,N_11685);
nor U12638 (N_12638,N_11710,N_11668);
and U12639 (N_12639,N_10551,N_10070);
xnor U12640 (N_12640,N_11962,N_11317);
and U12641 (N_12641,N_11017,N_10489);
nor U12642 (N_12642,N_10254,N_10304);
and U12643 (N_12643,N_10657,N_10181);
nand U12644 (N_12644,N_10826,N_10162);
or U12645 (N_12645,N_11813,N_11357);
nor U12646 (N_12646,N_11450,N_11898);
nand U12647 (N_12647,N_11863,N_11259);
or U12648 (N_12648,N_10782,N_10615);
nor U12649 (N_12649,N_11862,N_10716);
nor U12650 (N_12650,N_10574,N_10119);
or U12651 (N_12651,N_11584,N_10632);
xnor U12652 (N_12652,N_11611,N_10952);
xor U12653 (N_12653,N_11791,N_10473);
or U12654 (N_12654,N_10368,N_10271);
xnor U12655 (N_12655,N_10219,N_10803);
xnor U12656 (N_12656,N_11306,N_11841);
and U12657 (N_12657,N_10992,N_11729);
xnor U12658 (N_12658,N_10071,N_10327);
nor U12659 (N_12659,N_11148,N_11151);
or U12660 (N_12660,N_11804,N_10728);
and U12661 (N_12661,N_11150,N_10822);
xor U12662 (N_12662,N_11335,N_10911);
nand U12663 (N_12663,N_11707,N_10311);
or U12664 (N_12664,N_10956,N_10945);
nand U12665 (N_12665,N_10503,N_10697);
nand U12666 (N_12666,N_11859,N_11305);
or U12667 (N_12667,N_11039,N_11378);
nand U12668 (N_12668,N_10091,N_11092);
xor U12669 (N_12669,N_10172,N_11816);
or U12670 (N_12670,N_11454,N_10492);
nand U12671 (N_12671,N_11834,N_10820);
or U12672 (N_12672,N_10456,N_11220);
and U12673 (N_12673,N_10366,N_11285);
and U12674 (N_12674,N_11260,N_10198);
xor U12675 (N_12675,N_10380,N_10953);
xor U12676 (N_12676,N_11063,N_11337);
and U12677 (N_12677,N_10912,N_10723);
xor U12678 (N_12678,N_11262,N_10819);
nor U12679 (N_12679,N_10727,N_10977);
or U12680 (N_12680,N_11693,N_10522);
nor U12681 (N_12681,N_11702,N_11149);
nor U12682 (N_12682,N_10487,N_10598);
nor U12683 (N_12683,N_11953,N_11625);
or U12684 (N_12684,N_10688,N_10334);
xor U12685 (N_12685,N_11343,N_11292);
xor U12686 (N_12686,N_11264,N_11504);
nand U12687 (N_12687,N_10143,N_10336);
nor U12688 (N_12688,N_10844,N_11924);
nor U12689 (N_12689,N_11316,N_11399);
nor U12690 (N_12690,N_11493,N_10592);
nand U12691 (N_12691,N_11719,N_10437);
or U12692 (N_12692,N_10083,N_11049);
xor U12693 (N_12693,N_10791,N_10231);
xor U12694 (N_12694,N_10096,N_10981);
nor U12695 (N_12695,N_10527,N_11034);
xnor U12696 (N_12696,N_11723,N_10391);
nand U12697 (N_12697,N_10251,N_10588);
and U12698 (N_12698,N_11626,N_10158);
nand U12699 (N_12699,N_10523,N_11081);
or U12700 (N_12700,N_11681,N_10600);
nand U12701 (N_12701,N_11461,N_10868);
nor U12702 (N_12702,N_11027,N_10107);
xnor U12703 (N_12703,N_11489,N_10506);
and U12704 (N_12704,N_10664,N_11392);
or U12705 (N_12705,N_10917,N_11052);
nand U12706 (N_12706,N_11238,N_11029);
nand U12707 (N_12707,N_10477,N_10641);
or U12708 (N_12708,N_11738,N_11739);
or U12709 (N_12709,N_10283,N_11477);
nor U12710 (N_12710,N_11469,N_11692);
nor U12711 (N_12711,N_11193,N_11072);
or U12712 (N_12712,N_10255,N_10567);
xnor U12713 (N_12713,N_11772,N_10861);
nand U12714 (N_12714,N_11928,N_11884);
and U12715 (N_12715,N_10970,N_11090);
and U12716 (N_12716,N_11742,N_11566);
or U12717 (N_12717,N_11648,N_10125);
or U12718 (N_12718,N_10445,N_10138);
xnor U12719 (N_12719,N_11224,N_10619);
nor U12720 (N_12720,N_10720,N_11642);
nand U12721 (N_12721,N_11082,N_11634);
xor U12722 (N_12722,N_10613,N_11270);
xnor U12723 (N_12723,N_10605,N_10709);
xor U12724 (N_12724,N_11134,N_10378);
or U12725 (N_12725,N_11548,N_11613);
and U12726 (N_12726,N_10887,N_11694);
or U12727 (N_12727,N_11051,N_11930);
or U12728 (N_12728,N_11698,N_10347);
nor U12729 (N_12729,N_11545,N_11111);
nand U12730 (N_12730,N_10530,N_11521);
xor U12731 (N_12731,N_11697,N_10707);
and U12732 (N_12732,N_10899,N_11427);
and U12733 (N_12733,N_10817,N_11603);
nor U12734 (N_12734,N_11748,N_11418);
nor U12735 (N_12735,N_10382,N_11083);
or U12736 (N_12736,N_11656,N_11340);
and U12737 (N_12737,N_11188,N_11976);
nand U12738 (N_12738,N_11751,N_10816);
and U12739 (N_12739,N_10014,N_11499);
nor U12740 (N_12740,N_11348,N_11736);
and U12741 (N_12741,N_11524,N_10385);
and U12742 (N_12742,N_11936,N_11381);
nor U12743 (N_12743,N_10850,N_11612);
xor U12744 (N_12744,N_10407,N_10973);
nand U12745 (N_12745,N_10210,N_11018);
nor U12746 (N_12746,N_11683,N_11406);
nor U12747 (N_12747,N_11295,N_10515);
xnor U12748 (N_12748,N_10488,N_11846);
nor U12749 (N_12749,N_10222,N_11682);
nor U12750 (N_12750,N_11560,N_10770);
or U12751 (N_12751,N_11121,N_10661);
nor U12752 (N_12752,N_10930,N_11582);
or U12753 (N_12753,N_11779,N_10754);
or U12754 (N_12754,N_10048,N_10773);
nand U12755 (N_12755,N_11429,N_10021);
or U12756 (N_12756,N_10188,N_10475);
and U12757 (N_12757,N_11180,N_11279);
nor U12758 (N_12758,N_11139,N_11669);
nand U12759 (N_12759,N_11637,N_11974);
nand U12760 (N_12760,N_10169,N_11095);
or U12761 (N_12761,N_10942,N_10569);
nand U12762 (N_12762,N_11778,N_11935);
nor U12763 (N_12763,N_11311,N_10829);
nand U12764 (N_12764,N_11635,N_10272);
xnor U12765 (N_12765,N_11024,N_10780);
nand U12766 (N_12766,N_10869,N_10055);
nor U12767 (N_12767,N_11598,N_10587);
and U12768 (N_12768,N_10452,N_10037);
nand U12769 (N_12769,N_10546,N_11086);
nor U12770 (N_12770,N_10756,N_11367);
or U12771 (N_12771,N_11510,N_10286);
nor U12772 (N_12772,N_11021,N_11620);
xnor U12773 (N_12773,N_11483,N_11958);
and U12774 (N_12774,N_11302,N_11630);
nand U12775 (N_12775,N_10644,N_11005);
and U12776 (N_12776,N_10552,N_11241);
or U12777 (N_12777,N_10165,N_10557);
nor U12778 (N_12778,N_11319,N_10825);
xor U12779 (N_12779,N_10059,N_10684);
or U12780 (N_12780,N_11857,N_11275);
or U12781 (N_12781,N_10874,N_11549);
and U12782 (N_12782,N_10990,N_11140);
or U12783 (N_12783,N_10835,N_10935);
and U12784 (N_12784,N_10229,N_10752);
xor U12785 (N_12785,N_11607,N_10256);
and U12786 (N_12786,N_10591,N_10092);
xor U12787 (N_12787,N_11538,N_11110);
nand U12788 (N_12788,N_10959,N_10221);
nand U12789 (N_12789,N_11903,N_10000);
nand U12790 (N_12790,N_10936,N_11565);
nor U12791 (N_12791,N_10073,N_11770);
and U12792 (N_12792,N_11500,N_10923);
and U12793 (N_12793,N_10290,N_10875);
nor U12794 (N_12794,N_10994,N_11142);
nand U12795 (N_12795,N_10862,N_11925);
nor U12796 (N_12796,N_11254,N_11794);
and U12797 (N_12797,N_11202,N_11405);
or U12798 (N_12798,N_11252,N_10277);
and U12799 (N_12799,N_10390,N_11046);
nor U12800 (N_12800,N_11933,N_10067);
and U12801 (N_12801,N_11950,N_11578);
and U12802 (N_12802,N_11821,N_10167);
or U12803 (N_12803,N_11352,N_11655);
xor U12804 (N_12804,N_11042,N_10672);
and U12805 (N_12805,N_11745,N_11746);
xor U12806 (N_12806,N_10163,N_11628);
xnor U12807 (N_12807,N_11577,N_10142);
and U12808 (N_12808,N_11792,N_11492);
nor U12809 (N_12809,N_11564,N_11069);
xor U12810 (N_12810,N_10082,N_11867);
or U12811 (N_12811,N_10453,N_10253);
and U12812 (N_12812,N_11609,N_11070);
or U12813 (N_12813,N_10599,N_11044);
nand U12814 (N_12814,N_11616,N_11932);
nand U12815 (N_12815,N_10275,N_10656);
nand U12816 (N_12816,N_11170,N_10610);
nor U12817 (N_12817,N_10689,N_11397);
xor U12818 (N_12818,N_11795,N_11546);
or U12819 (N_12819,N_11897,N_11143);
or U12820 (N_12820,N_10430,N_11761);
or U12821 (N_12821,N_11330,N_11769);
xor U12822 (N_12822,N_11109,N_10918);
xor U12823 (N_12823,N_10439,N_11057);
and U12824 (N_12824,N_10401,N_10031);
or U12825 (N_12825,N_11006,N_11132);
xnor U12826 (N_12826,N_10017,N_11663);
nand U12827 (N_12827,N_11242,N_10794);
nor U12828 (N_12828,N_11442,N_11711);
or U12829 (N_12829,N_11187,N_10155);
nand U12830 (N_12830,N_11196,N_11651);
xnor U12831 (N_12831,N_11299,N_10326);
xnor U12832 (N_12832,N_11137,N_10637);
or U12833 (N_12833,N_11575,N_10064);
nor U12834 (N_12834,N_10666,N_11213);
nand U12835 (N_12835,N_10204,N_10027);
xnor U12836 (N_12836,N_10035,N_11556);
xnor U12837 (N_12837,N_11915,N_10628);
xnor U12838 (N_12838,N_10397,N_11101);
xnor U12839 (N_12839,N_11687,N_11995);
nor U12840 (N_12840,N_11514,N_11662);
nor U12841 (N_12841,N_10581,N_11929);
and U12842 (N_12842,N_10191,N_11624);
or U12843 (N_12843,N_10199,N_10273);
or U12844 (N_12844,N_10678,N_11014);
or U12845 (N_12845,N_11743,N_11872);
and U12846 (N_12846,N_11369,N_10408);
nand U12847 (N_12847,N_10909,N_10510);
nand U12848 (N_12848,N_11981,N_11112);
nor U12849 (N_12849,N_10556,N_11725);
and U12850 (N_12850,N_10562,N_10839);
nand U12851 (N_12851,N_11328,N_11064);
nand U12852 (N_12852,N_10686,N_11666);
xnor U12853 (N_12853,N_10315,N_10646);
and U12854 (N_12854,N_10045,N_11013);
nand U12855 (N_12855,N_11015,N_11096);
and U12856 (N_12856,N_11844,N_10295);
nand U12857 (N_12857,N_10571,N_10388);
nor U12858 (N_12858,N_10784,N_10072);
xor U12859 (N_12859,N_10963,N_11421);
and U12860 (N_12860,N_10698,N_11135);
xnor U12861 (N_12861,N_11098,N_11056);
or U12862 (N_12862,N_11678,N_10526);
xnor U12863 (N_12863,N_10792,N_10436);
xnor U12864 (N_12864,N_11115,N_11218);
or U12865 (N_12865,N_10383,N_11910);
nor U12866 (N_12866,N_11481,N_11155);
nand U12867 (N_12867,N_10485,N_11346);
nand U12868 (N_12868,N_10827,N_11227);
nand U12869 (N_12869,N_11515,N_10668);
and U12870 (N_12870,N_11255,N_10483);
or U12871 (N_12871,N_11583,N_10710);
xor U12872 (N_12872,N_11022,N_10907);
xor U12873 (N_12873,N_11377,N_10705);
nor U12874 (N_12874,N_10209,N_11496);
nand U12875 (N_12875,N_11533,N_10607);
and U12876 (N_12876,N_11433,N_10127);
xnor U12877 (N_12877,N_11641,N_11921);
nor U12878 (N_12878,N_10069,N_11943);
or U12879 (N_12879,N_10291,N_11726);
nor U12880 (N_12880,N_11009,N_10405);
or U12881 (N_12881,N_10620,N_11960);
or U12882 (N_12882,N_11053,N_11099);
or U12883 (N_12883,N_10715,N_11234);
nor U12884 (N_12884,N_10525,N_11436);
xnor U12885 (N_12885,N_10459,N_11741);
nand U12886 (N_12886,N_11526,N_11043);
xor U12887 (N_12887,N_10682,N_10848);
nor U12888 (N_12888,N_11475,N_10302);
and U12889 (N_12889,N_11372,N_11423);
and U12890 (N_12890,N_10718,N_10133);
xnor U12891 (N_12891,N_11646,N_10565);
and U12892 (N_12892,N_10886,N_11942);
and U12893 (N_12893,N_11522,N_10814);
and U12894 (N_12894,N_10392,N_10450);
xnor U12895 (N_12895,N_11873,N_11676);
nand U12896 (N_12896,N_11563,N_10018);
nor U12897 (N_12897,N_10278,N_11382);
nor U12898 (N_12898,N_11325,N_11458);
nand U12899 (N_12899,N_11465,N_10373);
or U12900 (N_12900,N_11621,N_10980);
nor U12901 (N_12901,N_10915,N_11768);
xor U12902 (N_12902,N_11415,N_11814);
and U12903 (N_12903,N_10215,N_11988);
or U12904 (N_12904,N_11589,N_10832);
and U12905 (N_12905,N_11456,N_10212);
nand U12906 (N_12906,N_10823,N_11980);
nand U12907 (N_12907,N_10540,N_11516);
xnor U12908 (N_12908,N_11131,N_10711);
nand U12909 (N_12909,N_11309,N_11201);
nor U12910 (N_12910,N_11485,N_11191);
nor U12911 (N_12911,N_10660,N_10098);
nor U12912 (N_12912,N_11398,N_10997);
xor U12913 (N_12913,N_11677,N_10513);
and U12914 (N_12914,N_10920,N_11701);
or U12915 (N_12915,N_10775,N_11688);
nor U12916 (N_12916,N_11374,N_11893);
and U12917 (N_12917,N_10184,N_10004);
or U12918 (N_12918,N_10135,N_11885);
or U12919 (N_12919,N_11544,N_11080);
nor U12920 (N_12920,N_10879,N_11077);
xnor U12921 (N_12921,N_10134,N_10220);
xnor U12922 (N_12922,N_11757,N_11716);
nor U12923 (N_12923,N_10533,N_11103);
and U12924 (N_12924,N_10317,N_10087);
or U12925 (N_12925,N_10355,N_10895);
nor U12926 (N_12926,N_11210,N_11964);
xor U12927 (N_12927,N_11774,N_11848);
or U12928 (N_12928,N_11269,N_11623);
xor U12929 (N_12929,N_10344,N_10974);
or U12930 (N_12930,N_11895,N_10852);
and U12931 (N_12931,N_10102,N_10840);
and U12932 (N_12932,N_11375,N_10554);
xnor U12933 (N_12933,N_11606,N_11211);
xnor U12934 (N_12934,N_10469,N_10338);
and U12935 (N_12935,N_11559,N_11162);
xnor U12936 (N_12936,N_11535,N_11754);
and U12937 (N_12937,N_11731,N_10681);
nand U12938 (N_12938,N_10279,N_11453);
nand U12939 (N_12939,N_10949,N_11189);
nand U12940 (N_12940,N_10361,N_10428);
xor U12941 (N_12941,N_10402,N_11636);
or U12942 (N_12942,N_11068,N_10179);
xnor U12943 (N_12943,N_11912,N_11047);
nor U12944 (N_12944,N_10100,N_11797);
nor U12945 (N_12945,N_10480,N_10925);
and U12946 (N_12946,N_11789,N_10774);
or U12947 (N_12947,N_10375,N_11909);
and U12948 (N_12948,N_11665,N_11691);
or U12949 (N_12949,N_11460,N_11965);
nor U12950 (N_12950,N_11116,N_10843);
and U12951 (N_12951,N_11368,N_11705);
or U12952 (N_12952,N_11478,N_11322);
xnor U12953 (N_12953,N_11391,N_11214);
nor U12954 (N_12954,N_10703,N_11977);
and U12955 (N_12955,N_11764,N_11880);
nand U12956 (N_12956,N_11593,N_11443);
nand U12957 (N_12957,N_11178,N_11845);
xor U12958 (N_12958,N_10441,N_11561);
xor U12959 (N_12959,N_10853,N_11653);
xor U12960 (N_12960,N_11075,N_11886);
nor U12961 (N_12961,N_10240,N_10352);
or U12962 (N_12962,N_10635,N_10236);
or U12963 (N_12963,N_10570,N_11376);
xor U12964 (N_12964,N_11441,N_10039);
nor U12965 (N_12965,N_10173,N_10462);
and U12966 (N_12966,N_11686,N_10807);
nand U12967 (N_12967,N_11766,N_11826);
and U12968 (N_12968,N_11718,N_11622);
and U12969 (N_12969,N_10837,N_10736);
xor U12970 (N_12970,N_10440,N_10520);
xnor U12971 (N_12971,N_11294,N_11649);
xnor U12972 (N_12972,N_10699,N_11344);
or U12973 (N_12973,N_11100,N_10132);
or U12974 (N_12974,N_11198,N_10356);
and U12975 (N_12975,N_10112,N_10670);
xnor U12976 (N_12976,N_10065,N_10066);
and U12977 (N_12977,N_10991,N_10987);
nor U12978 (N_12978,N_10350,N_11996);
nor U12979 (N_12979,N_11675,N_10595);
xnor U12980 (N_12980,N_10878,N_10365);
nand U12981 (N_12981,N_10312,N_11480);
nor U12982 (N_12982,N_11256,N_10080);
nor U12983 (N_12983,N_11093,N_10230);
nand U12984 (N_12984,N_11968,N_11818);
xnor U12985 (N_12985,N_10602,N_11998);
or U12986 (N_12986,N_10351,N_11219);
and U12987 (N_12987,N_11894,N_10178);
xor U12988 (N_12988,N_11164,N_10384);
or U12989 (N_12989,N_11847,N_10174);
xnor U12990 (N_12990,N_10712,N_10674);
nor U12991 (N_12991,N_10346,N_11520);
nand U12992 (N_12992,N_10860,N_11002);
xnor U12993 (N_12993,N_10870,N_10757);
and U12994 (N_12994,N_10360,N_10425);
and U12995 (N_12995,N_10053,N_11963);
or U12996 (N_12996,N_10884,N_10410);
and U12997 (N_12997,N_10933,N_10677);
and U12998 (N_12998,N_10676,N_10947);
xor U12999 (N_12999,N_11717,N_11866);
nand U13000 (N_13000,N_10240,N_10236);
and U13001 (N_13001,N_10252,N_11332);
or U13002 (N_13002,N_10510,N_10262);
or U13003 (N_13003,N_11839,N_11858);
nand U13004 (N_13004,N_10963,N_11288);
or U13005 (N_13005,N_11890,N_10222);
and U13006 (N_13006,N_11474,N_11871);
or U13007 (N_13007,N_11564,N_11072);
and U13008 (N_13008,N_11076,N_10494);
xor U13009 (N_13009,N_11497,N_11668);
nor U13010 (N_13010,N_11377,N_11490);
xor U13011 (N_13011,N_11932,N_10261);
and U13012 (N_13012,N_10766,N_10511);
nand U13013 (N_13013,N_11374,N_11081);
xnor U13014 (N_13014,N_11380,N_10134);
nand U13015 (N_13015,N_10518,N_11083);
and U13016 (N_13016,N_11832,N_11049);
nand U13017 (N_13017,N_11241,N_11011);
or U13018 (N_13018,N_11740,N_10500);
xor U13019 (N_13019,N_11534,N_10678);
or U13020 (N_13020,N_10046,N_11335);
nand U13021 (N_13021,N_11129,N_11955);
nand U13022 (N_13022,N_10134,N_11547);
xor U13023 (N_13023,N_11859,N_10485);
and U13024 (N_13024,N_10399,N_10630);
nand U13025 (N_13025,N_11684,N_10442);
xor U13026 (N_13026,N_10825,N_11485);
or U13027 (N_13027,N_11521,N_10055);
and U13028 (N_13028,N_10814,N_11447);
nand U13029 (N_13029,N_11711,N_11418);
xor U13030 (N_13030,N_11190,N_10899);
nand U13031 (N_13031,N_10441,N_10555);
or U13032 (N_13032,N_11034,N_11558);
or U13033 (N_13033,N_11037,N_10595);
and U13034 (N_13034,N_10794,N_10608);
xor U13035 (N_13035,N_11457,N_10701);
xor U13036 (N_13036,N_11594,N_10541);
nand U13037 (N_13037,N_11066,N_11661);
or U13038 (N_13038,N_10817,N_11260);
xor U13039 (N_13039,N_10062,N_10194);
nor U13040 (N_13040,N_11401,N_11469);
xor U13041 (N_13041,N_10470,N_10933);
and U13042 (N_13042,N_10504,N_11609);
and U13043 (N_13043,N_10554,N_11049);
xnor U13044 (N_13044,N_11728,N_10854);
xnor U13045 (N_13045,N_10898,N_10589);
nand U13046 (N_13046,N_10783,N_10578);
and U13047 (N_13047,N_11318,N_10795);
nand U13048 (N_13048,N_10483,N_10388);
or U13049 (N_13049,N_10749,N_11906);
nor U13050 (N_13050,N_11441,N_10024);
xor U13051 (N_13051,N_11385,N_10065);
nor U13052 (N_13052,N_11922,N_11306);
or U13053 (N_13053,N_10654,N_10752);
and U13054 (N_13054,N_11409,N_11896);
nor U13055 (N_13055,N_10699,N_10185);
xnor U13056 (N_13056,N_10122,N_11359);
and U13057 (N_13057,N_10512,N_11191);
nand U13058 (N_13058,N_11579,N_11921);
nor U13059 (N_13059,N_10543,N_11206);
and U13060 (N_13060,N_11771,N_10410);
or U13061 (N_13061,N_10607,N_10117);
or U13062 (N_13062,N_10936,N_11733);
and U13063 (N_13063,N_10847,N_10033);
and U13064 (N_13064,N_10713,N_10861);
or U13065 (N_13065,N_11938,N_11514);
nor U13066 (N_13066,N_10505,N_10023);
and U13067 (N_13067,N_11555,N_11875);
or U13068 (N_13068,N_10315,N_10016);
and U13069 (N_13069,N_11766,N_11509);
nor U13070 (N_13070,N_11495,N_10522);
or U13071 (N_13071,N_10451,N_10911);
nand U13072 (N_13072,N_10011,N_11222);
and U13073 (N_13073,N_11434,N_11931);
or U13074 (N_13074,N_11699,N_10575);
or U13075 (N_13075,N_11184,N_10384);
or U13076 (N_13076,N_11156,N_10464);
nand U13077 (N_13077,N_11796,N_10689);
nor U13078 (N_13078,N_11399,N_10578);
nand U13079 (N_13079,N_10076,N_10346);
and U13080 (N_13080,N_10100,N_11386);
and U13081 (N_13081,N_11364,N_10355);
and U13082 (N_13082,N_11242,N_11330);
xor U13083 (N_13083,N_11519,N_11405);
nor U13084 (N_13084,N_10038,N_11150);
and U13085 (N_13085,N_10191,N_10912);
xor U13086 (N_13086,N_10752,N_11924);
xnor U13087 (N_13087,N_10975,N_10932);
nor U13088 (N_13088,N_11325,N_10860);
nor U13089 (N_13089,N_11717,N_11874);
or U13090 (N_13090,N_11056,N_10106);
and U13091 (N_13091,N_11649,N_11704);
nor U13092 (N_13092,N_10285,N_11002);
xnor U13093 (N_13093,N_10353,N_10730);
xor U13094 (N_13094,N_10137,N_10568);
and U13095 (N_13095,N_10061,N_10506);
nand U13096 (N_13096,N_11471,N_10867);
xnor U13097 (N_13097,N_10043,N_10377);
nand U13098 (N_13098,N_10814,N_10273);
nor U13099 (N_13099,N_11808,N_11798);
nand U13100 (N_13100,N_11069,N_11375);
nor U13101 (N_13101,N_11127,N_11392);
xor U13102 (N_13102,N_11596,N_10974);
nor U13103 (N_13103,N_11857,N_11237);
and U13104 (N_13104,N_10578,N_11313);
and U13105 (N_13105,N_10011,N_11192);
xnor U13106 (N_13106,N_11400,N_10545);
or U13107 (N_13107,N_11370,N_11268);
nand U13108 (N_13108,N_10000,N_11176);
or U13109 (N_13109,N_11278,N_11687);
or U13110 (N_13110,N_10284,N_10456);
xnor U13111 (N_13111,N_11105,N_10910);
nor U13112 (N_13112,N_11910,N_11849);
xnor U13113 (N_13113,N_11532,N_11483);
or U13114 (N_13114,N_10441,N_11689);
nor U13115 (N_13115,N_11608,N_10142);
and U13116 (N_13116,N_10925,N_11838);
xnor U13117 (N_13117,N_11955,N_10036);
or U13118 (N_13118,N_10595,N_11268);
and U13119 (N_13119,N_10143,N_10569);
or U13120 (N_13120,N_11930,N_11420);
or U13121 (N_13121,N_11941,N_10565);
or U13122 (N_13122,N_11424,N_10922);
xnor U13123 (N_13123,N_10580,N_11416);
xnor U13124 (N_13124,N_11246,N_10650);
nand U13125 (N_13125,N_10372,N_11888);
nand U13126 (N_13126,N_11402,N_10186);
nand U13127 (N_13127,N_10197,N_11341);
and U13128 (N_13128,N_11960,N_10698);
nand U13129 (N_13129,N_11078,N_10991);
xnor U13130 (N_13130,N_10017,N_10231);
xor U13131 (N_13131,N_11727,N_11777);
xor U13132 (N_13132,N_10165,N_11610);
xor U13133 (N_13133,N_10080,N_11613);
or U13134 (N_13134,N_11993,N_10756);
xor U13135 (N_13135,N_11754,N_10904);
nor U13136 (N_13136,N_10238,N_10637);
nor U13137 (N_13137,N_11980,N_10535);
xnor U13138 (N_13138,N_10212,N_10858);
nand U13139 (N_13139,N_10540,N_10572);
xor U13140 (N_13140,N_11494,N_10654);
xnor U13141 (N_13141,N_11173,N_11123);
nor U13142 (N_13142,N_11554,N_10439);
nand U13143 (N_13143,N_10952,N_10004);
xor U13144 (N_13144,N_11011,N_10243);
nor U13145 (N_13145,N_11361,N_10132);
xor U13146 (N_13146,N_11494,N_10697);
nor U13147 (N_13147,N_11999,N_11039);
nand U13148 (N_13148,N_11133,N_10178);
nor U13149 (N_13149,N_10778,N_10102);
nor U13150 (N_13150,N_10898,N_10120);
xor U13151 (N_13151,N_11294,N_10496);
nand U13152 (N_13152,N_10761,N_10637);
nor U13153 (N_13153,N_10818,N_11200);
or U13154 (N_13154,N_11466,N_10589);
and U13155 (N_13155,N_11853,N_11672);
xor U13156 (N_13156,N_10435,N_11125);
nand U13157 (N_13157,N_10684,N_10981);
nor U13158 (N_13158,N_10534,N_11485);
or U13159 (N_13159,N_11415,N_10845);
nor U13160 (N_13160,N_10718,N_11581);
or U13161 (N_13161,N_11325,N_11528);
nor U13162 (N_13162,N_11814,N_11225);
nand U13163 (N_13163,N_10678,N_11302);
and U13164 (N_13164,N_11242,N_11854);
or U13165 (N_13165,N_11045,N_10502);
nand U13166 (N_13166,N_10791,N_11289);
or U13167 (N_13167,N_10050,N_11592);
nand U13168 (N_13168,N_10267,N_11325);
nand U13169 (N_13169,N_10921,N_10875);
xor U13170 (N_13170,N_11863,N_11113);
nand U13171 (N_13171,N_11649,N_10242);
and U13172 (N_13172,N_11472,N_10145);
nand U13173 (N_13173,N_11644,N_10498);
nor U13174 (N_13174,N_10369,N_11844);
nor U13175 (N_13175,N_11464,N_10759);
or U13176 (N_13176,N_11166,N_11341);
nand U13177 (N_13177,N_10300,N_11034);
nand U13178 (N_13178,N_11967,N_11633);
and U13179 (N_13179,N_10985,N_11090);
nand U13180 (N_13180,N_11305,N_10988);
and U13181 (N_13181,N_10292,N_11033);
nor U13182 (N_13182,N_11872,N_11135);
nand U13183 (N_13183,N_11573,N_10350);
and U13184 (N_13184,N_11969,N_10411);
xnor U13185 (N_13185,N_10857,N_11708);
or U13186 (N_13186,N_11743,N_10783);
nand U13187 (N_13187,N_11192,N_11262);
nor U13188 (N_13188,N_10727,N_10880);
and U13189 (N_13189,N_11544,N_10662);
and U13190 (N_13190,N_11051,N_10495);
and U13191 (N_13191,N_10839,N_11133);
nand U13192 (N_13192,N_11235,N_11885);
nor U13193 (N_13193,N_10175,N_10829);
or U13194 (N_13194,N_11007,N_11248);
and U13195 (N_13195,N_10022,N_11374);
and U13196 (N_13196,N_10620,N_11402);
nor U13197 (N_13197,N_11312,N_11524);
xnor U13198 (N_13198,N_10818,N_11579);
and U13199 (N_13199,N_11234,N_11202);
xnor U13200 (N_13200,N_11211,N_11993);
nand U13201 (N_13201,N_10182,N_10138);
xnor U13202 (N_13202,N_10475,N_11211);
nor U13203 (N_13203,N_11187,N_11815);
and U13204 (N_13204,N_11155,N_11607);
nor U13205 (N_13205,N_10380,N_10701);
or U13206 (N_13206,N_11398,N_10362);
and U13207 (N_13207,N_10633,N_10725);
xnor U13208 (N_13208,N_11407,N_10912);
xor U13209 (N_13209,N_10014,N_11204);
or U13210 (N_13210,N_11578,N_11140);
nor U13211 (N_13211,N_11965,N_11059);
or U13212 (N_13212,N_10689,N_10731);
and U13213 (N_13213,N_10439,N_11361);
nor U13214 (N_13214,N_11596,N_10654);
xnor U13215 (N_13215,N_11566,N_10757);
nor U13216 (N_13216,N_10792,N_10090);
or U13217 (N_13217,N_10281,N_10770);
and U13218 (N_13218,N_10818,N_10837);
xnor U13219 (N_13219,N_10720,N_10325);
and U13220 (N_13220,N_10937,N_11386);
or U13221 (N_13221,N_11574,N_11341);
nor U13222 (N_13222,N_10247,N_11835);
or U13223 (N_13223,N_11071,N_10533);
nand U13224 (N_13224,N_10591,N_10049);
nor U13225 (N_13225,N_11016,N_10148);
or U13226 (N_13226,N_10769,N_11565);
and U13227 (N_13227,N_10456,N_10401);
and U13228 (N_13228,N_11630,N_10467);
xnor U13229 (N_13229,N_10808,N_11892);
or U13230 (N_13230,N_11421,N_10929);
nand U13231 (N_13231,N_11842,N_10322);
or U13232 (N_13232,N_11528,N_11894);
and U13233 (N_13233,N_10460,N_10698);
xor U13234 (N_13234,N_11924,N_10465);
and U13235 (N_13235,N_10651,N_10065);
nand U13236 (N_13236,N_10966,N_10435);
or U13237 (N_13237,N_10783,N_10545);
nor U13238 (N_13238,N_10194,N_10650);
and U13239 (N_13239,N_10099,N_11373);
or U13240 (N_13240,N_10880,N_10152);
nor U13241 (N_13241,N_11647,N_10052);
xor U13242 (N_13242,N_11269,N_11823);
or U13243 (N_13243,N_10959,N_11706);
xor U13244 (N_13244,N_11110,N_11537);
or U13245 (N_13245,N_10676,N_10967);
nand U13246 (N_13246,N_10584,N_11587);
nand U13247 (N_13247,N_10828,N_10725);
xor U13248 (N_13248,N_10562,N_10224);
or U13249 (N_13249,N_11230,N_10054);
xor U13250 (N_13250,N_11801,N_10727);
nand U13251 (N_13251,N_11258,N_10882);
nor U13252 (N_13252,N_11526,N_11444);
xor U13253 (N_13253,N_10223,N_10518);
nor U13254 (N_13254,N_11098,N_11886);
nor U13255 (N_13255,N_10183,N_11397);
and U13256 (N_13256,N_10132,N_11989);
and U13257 (N_13257,N_10694,N_11793);
nand U13258 (N_13258,N_10245,N_10552);
xnor U13259 (N_13259,N_10012,N_11619);
and U13260 (N_13260,N_10054,N_10172);
nand U13261 (N_13261,N_11266,N_11943);
nand U13262 (N_13262,N_11741,N_10409);
xor U13263 (N_13263,N_10410,N_11658);
and U13264 (N_13264,N_10239,N_11647);
and U13265 (N_13265,N_10831,N_11395);
or U13266 (N_13266,N_10593,N_10821);
nor U13267 (N_13267,N_11878,N_10339);
or U13268 (N_13268,N_11316,N_10626);
nor U13269 (N_13269,N_11498,N_10878);
or U13270 (N_13270,N_11628,N_10546);
nor U13271 (N_13271,N_10975,N_10859);
and U13272 (N_13272,N_10376,N_11464);
and U13273 (N_13273,N_11181,N_10294);
nand U13274 (N_13274,N_11279,N_11634);
and U13275 (N_13275,N_10040,N_10401);
nor U13276 (N_13276,N_10185,N_10332);
xor U13277 (N_13277,N_10869,N_10529);
and U13278 (N_13278,N_11895,N_10015);
xor U13279 (N_13279,N_11247,N_11091);
and U13280 (N_13280,N_10211,N_11923);
and U13281 (N_13281,N_11119,N_11044);
nand U13282 (N_13282,N_10864,N_11055);
or U13283 (N_13283,N_10756,N_11114);
nor U13284 (N_13284,N_10076,N_10407);
xnor U13285 (N_13285,N_11856,N_11990);
or U13286 (N_13286,N_10935,N_10694);
or U13287 (N_13287,N_11536,N_10413);
and U13288 (N_13288,N_10444,N_11979);
nor U13289 (N_13289,N_11817,N_11250);
or U13290 (N_13290,N_10624,N_10583);
xnor U13291 (N_13291,N_10885,N_10297);
or U13292 (N_13292,N_11850,N_10427);
nor U13293 (N_13293,N_10063,N_10868);
or U13294 (N_13294,N_11161,N_10440);
xnor U13295 (N_13295,N_11605,N_10020);
nor U13296 (N_13296,N_11804,N_10587);
nor U13297 (N_13297,N_10821,N_11009);
nor U13298 (N_13298,N_10092,N_11109);
nor U13299 (N_13299,N_10388,N_10675);
xor U13300 (N_13300,N_10097,N_11087);
and U13301 (N_13301,N_11670,N_10967);
or U13302 (N_13302,N_11141,N_11417);
nand U13303 (N_13303,N_11981,N_10603);
nand U13304 (N_13304,N_10378,N_11609);
xnor U13305 (N_13305,N_10470,N_11738);
nor U13306 (N_13306,N_10437,N_11381);
xor U13307 (N_13307,N_11180,N_11447);
nor U13308 (N_13308,N_10508,N_11271);
xnor U13309 (N_13309,N_10860,N_10902);
and U13310 (N_13310,N_11358,N_11222);
xnor U13311 (N_13311,N_11567,N_10525);
nor U13312 (N_13312,N_11346,N_10137);
or U13313 (N_13313,N_11954,N_10239);
and U13314 (N_13314,N_11721,N_11346);
and U13315 (N_13315,N_11340,N_10078);
and U13316 (N_13316,N_11832,N_10173);
nor U13317 (N_13317,N_10583,N_11522);
or U13318 (N_13318,N_10838,N_11715);
nor U13319 (N_13319,N_10104,N_10998);
and U13320 (N_13320,N_11040,N_10498);
or U13321 (N_13321,N_11865,N_11688);
xnor U13322 (N_13322,N_10617,N_11352);
or U13323 (N_13323,N_11464,N_10076);
or U13324 (N_13324,N_11173,N_11375);
or U13325 (N_13325,N_11667,N_10382);
nor U13326 (N_13326,N_10979,N_11072);
xor U13327 (N_13327,N_10581,N_10842);
xor U13328 (N_13328,N_11181,N_10863);
and U13329 (N_13329,N_11634,N_10544);
or U13330 (N_13330,N_10127,N_10507);
xor U13331 (N_13331,N_10526,N_11615);
nand U13332 (N_13332,N_11221,N_11665);
nand U13333 (N_13333,N_11851,N_10151);
xnor U13334 (N_13334,N_10564,N_10650);
or U13335 (N_13335,N_10576,N_11939);
nand U13336 (N_13336,N_11376,N_11938);
nand U13337 (N_13337,N_11495,N_10034);
nor U13338 (N_13338,N_10909,N_11911);
or U13339 (N_13339,N_11005,N_11522);
nand U13340 (N_13340,N_10705,N_10326);
nand U13341 (N_13341,N_10516,N_11643);
or U13342 (N_13342,N_10909,N_10910);
and U13343 (N_13343,N_10681,N_11842);
xor U13344 (N_13344,N_10559,N_11240);
nor U13345 (N_13345,N_10228,N_11277);
nand U13346 (N_13346,N_10461,N_10513);
nand U13347 (N_13347,N_11047,N_10531);
or U13348 (N_13348,N_11645,N_11371);
xnor U13349 (N_13349,N_10034,N_11757);
nor U13350 (N_13350,N_11251,N_10002);
or U13351 (N_13351,N_10628,N_11322);
xor U13352 (N_13352,N_11514,N_10499);
nor U13353 (N_13353,N_10702,N_10238);
nor U13354 (N_13354,N_10865,N_11791);
nor U13355 (N_13355,N_11463,N_11277);
or U13356 (N_13356,N_11596,N_10909);
xnor U13357 (N_13357,N_10310,N_11562);
xor U13358 (N_13358,N_10524,N_11042);
or U13359 (N_13359,N_10156,N_10382);
or U13360 (N_13360,N_11533,N_10718);
nand U13361 (N_13361,N_10679,N_10544);
or U13362 (N_13362,N_11296,N_10101);
nor U13363 (N_13363,N_10350,N_10731);
and U13364 (N_13364,N_10200,N_11199);
and U13365 (N_13365,N_10522,N_11457);
and U13366 (N_13366,N_11995,N_10050);
and U13367 (N_13367,N_11072,N_11885);
xnor U13368 (N_13368,N_11672,N_10220);
and U13369 (N_13369,N_10117,N_10332);
and U13370 (N_13370,N_11489,N_10855);
and U13371 (N_13371,N_10251,N_10542);
nand U13372 (N_13372,N_11242,N_11687);
or U13373 (N_13373,N_11888,N_10331);
or U13374 (N_13374,N_11778,N_11739);
nand U13375 (N_13375,N_10031,N_11228);
nand U13376 (N_13376,N_10134,N_11272);
and U13377 (N_13377,N_10073,N_11538);
nor U13378 (N_13378,N_11030,N_11074);
nor U13379 (N_13379,N_11914,N_10969);
xnor U13380 (N_13380,N_11577,N_10867);
or U13381 (N_13381,N_11812,N_10546);
and U13382 (N_13382,N_10422,N_10101);
nand U13383 (N_13383,N_10555,N_11090);
nor U13384 (N_13384,N_11899,N_10769);
xor U13385 (N_13385,N_11253,N_11380);
nand U13386 (N_13386,N_10628,N_10108);
xnor U13387 (N_13387,N_11483,N_11460);
nor U13388 (N_13388,N_11177,N_10310);
and U13389 (N_13389,N_10515,N_11375);
or U13390 (N_13390,N_10704,N_10171);
nor U13391 (N_13391,N_10931,N_10173);
and U13392 (N_13392,N_11106,N_11205);
or U13393 (N_13393,N_11539,N_11012);
xor U13394 (N_13394,N_11385,N_10298);
or U13395 (N_13395,N_10643,N_10766);
or U13396 (N_13396,N_11065,N_11431);
nor U13397 (N_13397,N_10515,N_10902);
or U13398 (N_13398,N_10666,N_10781);
nand U13399 (N_13399,N_11264,N_10355);
nor U13400 (N_13400,N_11879,N_11137);
nor U13401 (N_13401,N_10399,N_11435);
and U13402 (N_13402,N_11444,N_11883);
and U13403 (N_13403,N_10553,N_11853);
nand U13404 (N_13404,N_10340,N_11188);
nand U13405 (N_13405,N_11337,N_10765);
or U13406 (N_13406,N_11766,N_10876);
xnor U13407 (N_13407,N_11875,N_10114);
and U13408 (N_13408,N_10484,N_11606);
or U13409 (N_13409,N_11783,N_10069);
or U13410 (N_13410,N_10974,N_10504);
nand U13411 (N_13411,N_10847,N_11825);
nand U13412 (N_13412,N_11421,N_10060);
nor U13413 (N_13413,N_10831,N_10154);
nand U13414 (N_13414,N_11081,N_11891);
nand U13415 (N_13415,N_11522,N_10362);
nor U13416 (N_13416,N_10440,N_10756);
or U13417 (N_13417,N_10676,N_10487);
and U13418 (N_13418,N_11525,N_11185);
or U13419 (N_13419,N_11465,N_11565);
nor U13420 (N_13420,N_11350,N_10537);
nor U13421 (N_13421,N_11549,N_11110);
or U13422 (N_13422,N_11653,N_11453);
and U13423 (N_13423,N_10304,N_11926);
or U13424 (N_13424,N_10605,N_11602);
xor U13425 (N_13425,N_10309,N_11227);
nor U13426 (N_13426,N_11738,N_10065);
nor U13427 (N_13427,N_11520,N_11930);
nor U13428 (N_13428,N_10867,N_11624);
or U13429 (N_13429,N_10806,N_11645);
nand U13430 (N_13430,N_10913,N_11363);
and U13431 (N_13431,N_11443,N_11880);
xnor U13432 (N_13432,N_10169,N_10139);
or U13433 (N_13433,N_10644,N_11833);
and U13434 (N_13434,N_10868,N_10366);
xnor U13435 (N_13435,N_10961,N_11262);
nand U13436 (N_13436,N_10938,N_11625);
and U13437 (N_13437,N_11557,N_11106);
or U13438 (N_13438,N_11311,N_10234);
xor U13439 (N_13439,N_11096,N_11317);
nor U13440 (N_13440,N_11482,N_11546);
nand U13441 (N_13441,N_11764,N_11438);
nor U13442 (N_13442,N_11659,N_10288);
nor U13443 (N_13443,N_10112,N_11890);
and U13444 (N_13444,N_10178,N_10338);
or U13445 (N_13445,N_11724,N_10401);
or U13446 (N_13446,N_11193,N_10908);
nand U13447 (N_13447,N_10896,N_10837);
or U13448 (N_13448,N_11725,N_10513);
nand U13449 (N_13449,N_10734,N_10350);
or U13450 (N_13450,N_10093,N_11720);
xnor U13451 (N_13451,N_11065,N_11399);
xnor U13452 (N_13452,N_11887,N_11819);
or U13453 (N_13453,N_11072,N_10718);
nor U13454 (N_13454,N_11876,N_11510);
nand U13455 (N_13455,N_11170,N_10856);
nor U13456 (N_13456,N_11698,N_11627);
and U13457 (N_13457,N_10147,N_11035);
and U13458 (N_13458,N_11119,N_10608);
nor U13459 (N_13459,N_11445,N_10525);
nor U13460 (N_13460,N_11799,N_10363);
or U13461 (N_13461,N_11373,N_11244);
xor U13462 (N_13462,N_10331,N_10639);
nor U13463 (N_13463,N_11936,N_10555);
and U13464 (N_13464,N_10672,N_11797);
nor U13465 (N_13465,N_11411,N_11107);
and U13466 (N_13466,N_11648,N_10614);
nor U13467 (N_13467,N_10590,N_10487);
nor U13468 (N_13468,N_11731,N_10861);
xnor U13469 (N_13469,N_10306,N_10242);
and U13470 (N_13470,N_10661,N_10484);
nor U13471 (N_13471,N_11756,N_10561);
xnor U13472 (N_13472,N_10367,N_10156);
xor U13473 (N_13473,N_11918,N_10876);
nand U13474 (N_13474,N_11718,N_11944);
nand U13475 (N_13475,N_11895,N_10228);
nor U13476 (N_13476,N_11069,N_11135);
and U13477 (N_13477,N_11388,N_11027);
xor U13478 (N_13478,N_11966,N_11530);
and U13479 (N_13479,N_10275,N_11312);
or U13480 (N_13480,N_10501,N_10813);
nor U13481 (N_13481,N_10244,N_10987);
and U13482 (N_13482,N_10360,N_11209);
nand U13483 (N_13483,N_10161,N_11906);
and U13484 (N_13484,N_11669,N_10990);
nand U13485 (N_13485,N_10872,N_10683);
nand U13486 (N_13486,N_11522,N_10913);
and U13487 (N_13487,N_11132,N_11452);
nand U13488 (N_13488,N_10722,N_10246);
or U13489 (N_13489,N_11623,N_10099);
xnor U13490 (N_13490,N_10116,N_11746);
nor U13491 (N_13491,N_10177,N_11273);
and U13492 (N_13492,N_10901,N_11210);
nor U13493 (N_13493,N_11610,N_10301);
nor U13494 (N_13494,N_11820,N_11792);
nand U13495 (N_13495,N_11222,N_10195);
xnor U13496 (N_13496,N_11835,N_11317);
xor U13497 (N_13497,N_10830,N_11019);
or U13498 (N_13498,N_10247,N_10764);
nand U13499 (N_13499,N_10731,N_10137);
nor U13500 (N_13500,N_10458,N_11632);
or U13501 (N_13501,N_11013,N_10552);
nand U13502 (N_13502,N_11011,N_10029);
xnor U13503 (N_13503,N_11177,N_10615);
xnor U13504 (N_13504,N_11119,N_10965);
and U13505 (N_13505,N_11670,N_11801);
or U13506 (N_13506,N_11303,N_10235);
nor U13507 (N_13507,N_10852,N_10303);
nand U13508 (N_13508,N_10182,N_10859);
or U13509 (N_13509,N_10801,N_11647);
or U13510 (N_13510,N_10393,N_11969);
nand U13511 (N_13511,N_11083,N_11703);
and U13512 (N_13512,N_11955,N_10261);
nor U13513 (N_13513,N_10575,N_10061);
and U13514 (N_13514,N_11101,N_10839);
or U13515 (N_13515,N_11812,N_11169);
xnor U13516 (N_13516,N_11228,N_10017);
and U13517 (N_13517,N_11696,N_10498);
or U13518 (N_13518,N_10310,N_11227);
and U13519 (N_13519,N_10571,N_11656);
nand U13520 (N_13520,N_10597,N_11425);
or U13521 (N_13521,N_11469,N_10117);
nand U13522 (N_13522,N_11626,N_11287);
and U13523 (N_13523,N_10574,N_10823);
or U13524 (N_13524,N_11266,N_10081);
nor U13525 (N_13525,N_10804,N_11789);
and U13526 (N_13526,N_11075,N_11870);
and U13527 (N_13527,N_10000,N_10064);
nand U13528 (N_13528,N_10817,N_11573);
xnor U13529 (N_13529,N_11493,N_10603);
nand U13530 (N_13530,N_10702,N_10980);
and U13531 (N_13531,N_11738,N_11844);
nor U13532 (N_13532,N_10237,N_10760);
nor U13533 (N_13533,N_10346,N_10410);
or U13534 (N_13534,N_11637,N_10050);
nor U13535 (N_13535,N_11099,N_11694);
nor U13536 (N_13536,N_11561,N_11878);
nor U13537 (N_13537,N_11539,N_10158);
nand U13538 (N_13538,N_11196,N_10708);
nor U13539 (N_13539,N_11534,N_10567);
or U13540 (N_13540,N_11553,N_10782);
and U13541 (N_13541,N_11908,N_10889);
or U13542 (N_13542,N_11800,N_10063);
or U13543 (N_13543,N_10023,N_11674);
nor U13544 (N_13544,N_11659,N_10621);
nand U13545 (N_13545,N_11945,N_11627);
and U13546 (N_13546,N_11902,N_10307);
nor U13547 (N_13547,N_10380,N_11019);
xor U13548 (N_13548,N_10768,N_10638);
nor U13549 (N_13549,N_10102,N_11722);
nand U13550 (N_13550,N_11845,N_11141);
nand U13551 (N_13551,N_10858,N_11967);
and U13552 (N_13552,N_11784,N_10444);
or U13553 (N_13553,N_10916,N_11790);
xnor U13554 (N_13554,N_10749,N_11703);
xnor U13555 (N_13555,N_11904,N_10163);
nor U13556 (N_13556,N_11991,N_10761);
or U13557 (N_13557,N_10914,N_10342);
xnor U13558 (N_13558,N_11638,N_10928);
or U13559 (N_13559,N_10957,N_10943);
nor U13560 (N_13560,N_10996,N_10798);
nor U13561 (N_13561,N_11579,N_11893);
nand U13562 (N_13562,N_11901,N_10038);
nor U13563 (N_13563,N_11029,N_10199);
nand U13564 (N_13564,N_11161,N_11047);
and U13565 (N_13565,N_11241,N_11638);
nor U13566 (N_13566,N_11399,N_11427);
nand U13567 (N_13567,N_10889,N_11807);
xor U13568 (N_13568,N_10877,N_11959);
or U13569 (N_13569,N_11439,N_10647);
or U13570 (N_13570,N_10834,N_11624);
xnor U13571 (N_13571,N_11434,N_11525);
and U13572 (N_13572,N_11573,N_10811);
and U13573 (N_13573,N_11130,N_10889);
or U13574 (N_13574,N_11835,N_11450);
or U13575 (N_13575,N_11174,N_10739);
nand U13576 (N_13576,N_10979,N_11762);
or U13577 (N_13577,N_10233,N_11724);
or U13578 (N_13578,N_11510,N_10846);
and U13579 (N_13579,N_10944,N_11283);
and U13580 (N_13580,N_11488,N_11771);
xor U13581 (N_13581,N_10237,N_10040);
and U13582 (N_13582,N_11106,N_10868);
or U13583 (N_13583,N_10644,N_10783);
nor U13584 (N_13584,N_11785,N_11082);
nor U13585 (N_13585,N_11801,N_10691);
nor U13586 (N_13586,N_10629,N_11395);
xor U13587 (N_13587,N_10208,N_10316);
xnor U13588 (N_13588,N_10939,N_11525);
or U13589 (N_13589,N_10499,N_11760);
xor U13590 (N_13590,N_11118,N_10133);
and U13591 (N_13591,N_11307,N_11733);
nand U13592 (N_13592,N_10545,N_11598);
and U13593 (N_13593,N_10382,N_11500);
or U13594 (N_13594,N_11519,N_10271);
and U13595 (N_13595,N_11074,N_10206);
and U13596 (N_13596,N_11687,N_10598);
xor U13597 (N_13597,N_11625,N_11902);
or U13598 (N_13598,N_11901,N_10601);
or U13599 (N_13599,N_10905,N_11336);
or U13600 (N_13600,N_11068,N_10743);
and U13601 (N_13601,N_10914,N_11078);
xnor U13602 (N_13602,N_10902,N_10286);
nand U13603 (N_13603,N_10592,N_10817);
and U13604 (N_13604,N_10171,N_10709);
xnor U13605 (N_13605,N_11642,N_10644);
xnor U13606 (N_13606,N_11772,N_11988);
xnor U13607 (N_13607,N_10727,N_11555);
nand U13608 (N_13608,N_10289,N_10220);
and U13609 (N_13609,N_10365,N_10440);
nor U13610 (N_13610,N_10019,N_10195);
nand U13611 (N_13611,N_11544,N_11333);
or U13612 (N_13612,N_11934,N_10919);
nand U13613 (N_13613,N_10039,N_11711);
nor U13614 (N_13614,N_11667,N_11381);
xnor U13615 (N_13615,N_10170,N_10468);
nor U13616 (N_13616,N_11685,N_11996);
nor U13617 (N_13617,N_10026,N_10642);
or U13618 (N_13618,N_11115,N_11879);
or U13619 (N_13619,N_11993,N_10188);
nand U13620 (N_13620,N_11382,N_11101);
nor U13621 (N_13621,N_10965,N_11863);
nor U13622 (N_13622,N_10249,N_10349);
and U13623 (N_13623,N_10705,N_10683);
or U13624 (N_13624,N_11802,N_11038);
nor U13625 (N_13625,N_11418,N_11929);
or U13626 (N_13626,N_10282,N_10346);
nor U13627 (N_13627,N_10672,N_10653);
nand U13628 (N_13628,N_10443,N_10785);
nand U13629 (N_13629,N_11387,N_11845);
nand U13630 (N_13630,N_11529,N_10157);
or U13631 (N_13631,N_11157,N_10907);
nand U13632 (N_13632,N_10896,N_11863);
xor U13633 (N_13633,N_11922,N_11006);
xnor U13634 (N_13634,N_11423,N_10639);
or U13635 (N_13635,N_11783,N_11340);
xor U13636 (N_13636,N_11756,N_10263);
xor U13637 (N_13637,N_10987,N_10349);
or U13638 (N_13638,N_10755,N_10908);
and U13639 (N_13639,N_10536,N_10217);
xor U13640 (N_13640,N_11707,N_10204);
nand U13641 (N_13641,N_11386,N_10502);
nor U13642 (N_13642,N_11286,N_11102);
xor U13643 (N_13643,N_11586,N_10835);
xnor U13644 (N_13644,N_10620,N_10011);
or U13645 (N_13645,N_10788,N_10902);
and U13646 (N_13646,N_10242,N_10548);
xnor U13647 (N_13647,N_10865,N_11947);
nand U13648 (N_13648,N_11374,N_11971);
or U13649 (N_13649,N_11241,N_11442);
xnor U13650 (N_13650,N_11554,N_10233);
nor U13651 (N_13651,N_10223,N_11539);
nor U13652 (N_13652,N_10266,N_11638);
nand U13653 (N_13653,N_11080,N_10522);
nor U13654 (N_13654,N_11207,N_11995);
nand U13655 (N_13655,N_11618,N_10830);
xnor U13656 (N_13656,N_10841,N_11620);
xnor U13657 (N_13657,N_10553,N_11704);
and U13658 (N_13658,N_10262,N_11696);
nor U13659 (N_13659,N_11037,N_10822);
nor U13660 (N_13660,N_10043,N_11915);
xnor U13661 (N_13661,N_10061,N_11918);
nor U13662 (N_13662,N_10654,N_11887);
nand U13663 (N_13663,N_10068,N_10257);
nor U13664 (N_13664,N_10021,N_10042);
or U13665 (N_13665,N_10400,N_11092);
or U13666 (N_13666,N_11190,N_10071);
or U13667 (N_13667,N_10255,N_11878);
and U13668 (N_13668,N_10892,N_11958);
nor U13669 (N_13669,N_11744,N_11526);
and U13670 (N_13670,N_10554,N_10006);
nor U13671 (N_13671,N_11570,N_11189);
xor U13672 (N_13672,N_10702,N_11265);
nor U13673 (N_13673,N_10306,N_11440);
xor U13674 (N_13674,N_10441,N_10023);
xor U13675 (N_13675,N_10057,N_11323);
or U13676 (N_13676,N_10850,N_11912);
nor U13677 (N_13677,N_10922,N_10089);
and U13678 (N_13678,N_11094,N_11373);
or U13679 (N_13679,N_11137,N_11423);
or U13680 (N_13680,N_11266,N_11336);
nand U13681 (N_13681,N_11299,N_11166);
xnor U13682 (N_13682,N_11943,N_11848);
nor U13683 (N_13683,N_11615,N_11470);
nand U13684 (N_13684,N_10486,N_11286);
and U13685 (N_13685,N_10224,N_11733);
and U13686 (N_13686,N_11058,N_11217);
xnor U13687 (N_13687,N_11518,N_11437);
or U13688 (N_13688,N_11329,N_11555);
xnor U13689 (N_13689,N_10929,N_11661);
nor U13690 (N_13690,N_11951,N_11849);
nand U13691 (N_13691,N_11641,N_10732);
xor U13692 (N_13692,N_11285,N_10288);
nand U13693 (N_13693,N_10798,N_11332);
nand U13694 (N_13694,N_10993,N_11956);
xor U13695 (N_13695,N_11504,N_11867);
and U13696 (N_13696,N_10709,N_10799);
or U13697 (N_13697,N_10905,N_10477);
and U13698 (N_13698,N_10659,N_11954);
xnor U13699 (N_13699,N_10442,N_10203);
nand U13700 (N_13700,N_11801,N_10359);
nor U13701 (N_13701,N_10115,N_11802);
nor U13702 (N_13702,N_10162,N_10879);
and U13703 (N_13703,N_11409,N_10433);
nand U13704 (N_13704,N_11966,N_10895);
and U13705 (N_13705,N_11184,N_10962);
xnor U13706 (N_13706,N_10781,N_11083);
xor U13707 (N_13707,N_10330,N_10962);
xnor U13708 (N_13708,N_10289,N_11133);
or U13709 (N_13709,N_11295,N_10446);
or U13710 (N_13710,N_11023,N_10248);
nand U13711 (N_13711,N_10473,N_10884);
nor U13712 (N_13712,N_11975,N_10239);
nand U13713 (N_13713,N_10069,N_11076);
nand U13714 (N_13714,N_10884,N_11569);
xnor U13715 (N_13715,N_10700,N_11110);
nor U13716 (N_13716,N_11902,N_10591);
xnor U13717 (N_13717,N_10801,N_10861);
xnor U13718 (N_13718,N_10371,N_10947);
nand U13719 (N_13719,N_10943,N_10418);
and U13720 (N_13720,N_11231,N_10766);
xnor U13721 (N_13721,N_10678,N_10188);
or U13722 (N_13722,N_11726,N_10958);
and U13723 (N_13723,N_10147,N_11324);
and U13724 (N_13724,N_10724,N_10695);
xor U13725 (N_13725,N_11261,N_10723);
nand U13726 (N_13726,N_11267,N_11632);
or U13727 (N_13727,N_10299,N_11207);
and U13728 (N_13728,N_11627,N_11944);
nand U13729 (N_13729,N_11084,N_11729);
or U13730 (N_13730,N_11011,N_11342);
or U13731 (N_13731,N_10499,N_10236);
xor U13732 (N_13732,N_11981,N_11975);
and U13733 (N_13733,N_11011,N_10187);
xor U13734 (N_13734,N_11966,N_10781);
nand U13735 (N_13735,N_11945,N_10210);
xnor U13736 (N_13736,N_10155,N_11827);
xor U13737 (N_13737,N_11565,N_11144);
nor U13738 (N_13738,N_10750,N_11967);
and U13739 (N_13739,N_11563,N_11911);
or U13740 (N_13740,N_11249,N_10615);
and U13741 (N_13741,N_11515,N_10037);
nand U13742 (N_13742,N_11259,N_10262);
nand U13743 (N_13743,N_10641,N_11479);
nand U13744 (N_13744,N_10476,N_10553);
nand U13745 (N_13745,N_10173,N_10177);
xor U13746 (N_13746,N_11235,N_10796);
and U13747 (N_13747,N_10190,N_10316);
nor U13748 (N_13748,N_11677,N_11165);
or U13749 (N_13749,N_11311,N_11167);
and U13750 (N_13750,N_11125,N_11640);
and U13751 (N_13751,N_10821,N_11441);
xnor U13752 (N_13752,N_10388,N_10833);
or U13753 (N_13753,N_11724,N_10574);
xnor U13754 (N_13754,N_11609,N_10123);
xor U13755 (N_13755,N_11188,N_10999);
and U13756 (N_13756,N_10519,N_10136);
and U13757 (N_13757,N_11264,N_10047);
xor U13758 (N_13758,N_11185,N_11803);
xnor U13759 (N_13759,N_11968,N_10769);
xnor U13760 (N_13760,N_10224,N_10655);
and U13761 (N_13761,N_10309,N_11650);
and U13762 (N_13762,N_10327,N_10406);
and U13763 (N_13763,N_11652,N_11569);
xor U13764 (N_13764,N_11648,N_10242);
or U13765 (N_13765,N_11361,N_10274);
or U13766 (N_13766,N_10015,N_11871);
or U13767 (N_13767,N_11263,N_10636);
xor U13768 (N_13768,N_11211,N_11406);
xnor U13769 (N_13769,N_10863,N_11012);
or U13770 (N_13770,N_10916,N_10143);
xor U13771 (N_13771,N_11201,N_10713);
nand U13772 (N_13772,N_11383,N_11526);
and U13773 (N_13773,N_10773,N_10690);
and U13774 (N_13774,N_11981,N_11784);
nor U13775 (N_13775,N_10454,N_10408);
and U13776 (N_13776,N_11076,N_11804);
xnor U13777 (N_13777,N_11421,N_11493);
or U13778 (N_13778,N_10273,N_11359);
xnor U13779 (N_13779,N_11021,N_11596);
xnor U13780 (N_13780,N_11247,N_11906);
xnor U13781 (N_13781,N_10783,N_10892);
and U13782 (N_13782,N_11821,N_11692);
nand U13783 (N_13783,N_11252,N_10436);
nor U13784 (N_13784,N_10090,N_10801);
xor U13785 (N_13785,N_11397,N_10458);
nand U13786 (N_13786,N_10200,N_10724);
nor U13787 (N_13787,N_11810,N_10301);
nand U13788 (N_13788,N_10036,N_10701);
or U13789 (N_13789,N_10286,N_11124);
and U13790 (N_13790,N_11932,N_10136);
and U13791 (N_13791,N_11054,N_10053);
xor U13792 (N_13792,N_10058,N_10577);
nor U13793 (N_13793,N_10771,N_10215);
nand U13794 (N_13794,N_11979,N_11254);
nor U13795 (N_13795,N_11757,N_10128);
nand U13796 (N_13796,N_11413,N_10527);
xor U13797 (N_13797,N_11226,N_11667);
nand U13798 (N_13798,N_11540,N_11747);
nand U13799 (N_13799,N_10986,N_10418);
nor U13800 (N_13800,N_10469,N_11130);
nor U13801 (N_13801,N_11867,N_10642);
and U13802 (N_13802,N_11568,N_11737);
xor U13803 (N_13803,N_10272,N_11123);
nand U13804 (N_13804,N_10003,N_11262);
nand U13805 (N_13805,N_11355,N_10873);
nor U13806 (N_13806,N_11906,N_11748);
or U13807 (N_13807,N_11673,N_11337);
xnor U13808 (N_13808,N_10693,N_10957);
nand U13809 (N_13809,N_10018,N_10508);
nand U13810 (N_13810,N_11264,N_11430);
nor U13811 (N_13811,N_11085,N_10526);
nor U13812 (N_13812,N_10637,N_10885);
nor U13813 (N_13813,N_11493,N_10392);
nor U13814 (N_13814,N_11560,N_10031);
nand U13815 (N_13815,N_11359,N_10477);
xor U13816 (N_13816,N_11991,N_10681);
or U13817 (N_13817,N_11672,N_11704);
nor U13818 (N_13818,N_10204,N_11401);
or U13819 (N_13819,N_11398,N_10097);
and U13820 (N_13820,N_11855,N_11783);
or U13821 (N_13821,N_10646,N_10598);
nand U13822 (N_13822,N_11981,N_11002);
xor U13823 (N_13823,N_10097,N_10274);
and U13824 (N_13824,N_10390,N_10363);
or U13825 (N_13825,N_11456,N_11192);
or U13826 (N_13826,N_10471,N_11479);
and U13827 (N_13827,N_10780,N_10733);
nand U13828 (N_13828,N_11639,N_11573);
nand U13829 (N_13829,N_10442,N_11342);
nor U13830 (N_13830,N_10188,N_11979);
nor U13831 (N_13831,N_10778,N_11939);
xnor U13832 (N_13832,N_11156,N_11759);
nand U13833 (N_13833,N_10249,N_10133);
nand U13834 (N_13834,N_11165,N_11422);
nor U13835 (N_13835,N_10016,N_10226);
nand U13836 (N_13836,N_11357,N_10153);
nor U13837 (N_13837,N_11165,N_11102);
and U13838 (N_13838,N_10408,N_10481);
xor U13839 (N_13839,N_11132,N_10747);
nand U13840 (N_13840,N_11201,N_11092);
and U13841 (N_13841,N_11977,N_11930);
xor U13842 (N_13842,N_11062,N_10840);
nor U13843 (N_13843,N_10655,N_10942);
or U13844 (N_13844,N_10100,N_10963);
xnor U13845 (N_13845,N_10279,N_11914);
or U13846 (N_13846,N_10661,N_11733);
nand U13847 (N_13847,N_11022,N_11246);
and U13848 (N_13848,N_10158,N_11724);
or U13849 (N_13849,N_10863,N_10148);
nand U13850 (N_13850,N_10790,N_11559);
or U13851 (N_13851,N_11316,N_11188);
nand U13852 (N_13852,N_10881,N_10559);
nor U13853 (N_13853,N_10935,N_10398);
nor U13854 (N_13854,N_11867,N_11208);
xnor U13855 (N_13855,N_10969,N_10423);
nor U13856 (N_13856,N_11230,N_11084);
or U13857 (N_13857,N_10924,N_11363);
xnor U13858 (N_13858,N_11621,N_10482);
xnor U13859 (N_13859,N_10546,N_10181);
nor U13860 (N_13860,N_10193,N_10385);
xor U13861 (N_13861,N_11607,N_11927);
nor U13862 (N_13862,N_11875,N_10128);
nor U13863 (N_13863,N_11286,N_11460);
or U13864 (N_13864,N_10749,N_10534);
xnor U13865 (N_13865,N_10713,N_10607);
xnor U13866 (N_13866,N_11882,N_11277);
nand U13867 (N_13867,N_11222,N_11286);
xor U13868 (N_13868,N_11779,N_10003);
nand U13869 (N_13869,N_11547,N_10783);
nand U13870 (N_13870,N_10139,N_10155);
and U13871 (N_13871,N_11608,N_11816);
and U13872 (N_13872,N_10210,N_11422);
and U13873 (N_13873,N_10811,N_10535);
and U13874 (N_13874,N_11702,N_10939);
nor U13875 (N_13875,N_11626,N_10431);
nor U13876 (N_13876,N_11816,N_10971);
nand U13877 (N_13877,N_11484,N_11584);
nand U13878 (N_13878,N_10450,N_10367);
nand U13879 (N_13879,N_10587,N_10630);
and U13880 (N_13880,N_10633,N_10265);
nand U13881 (N_13881,N_11634,N_10248);
nor U13882 (N_13882,N_11269,N_10363);
and U13883 (N_13883,N_10988,N_10950);
or U13884 (N_13884,N_10843,N_10152);
nor U13885 (N_13885,N_11115,N_10252);
xnor U13886 (N_13886,N_11619,N_10260);
nor U13887 (N_13887,N_11725,N_11920);
nor U13888 (N_13888,N_10064,N_11072);
nand U13889 (N_13889,N_10848,N_10910);
nor U13890 (N_13890,N_11723,N_10207);
nand U13891 (N_13891,N_10838,N_11722);
nor U13892 (N_13892,N_11766,N_11977);
and U13893 (N_13893,N_11949,N_10143);
xor U13894 (N_13894,N_11866,N_11013);
nand U13895 (N_13895,N_10113,N_10391);
nand U13896 (N_13896,N_11856,N_11138);
xor U13897 (N_13897,N_11717,N_10473);
nor U13898 (N_13898,N_11863,N_11269);
or U13899 (N_13899,N_10708,N_11903);
xor U13900 (N_13900,N_10804,N_11131);
nand U13901 (N_13901,N_10840,N_10876);
nand U13902 (N_13902,N_11605,N_11692);
and U13903 (N_13903,N_11896,N_10431);
nand U13904 (N_13904,N_10101,N_11896);
xnor U13905 (N_13905,N_10258,N_11616);
or U13906 (N_13906,N_11993,N_10045);
or U13907 (N_13907,N_10775,N_11432);
or U13908 (N_13908,N_10576,N_10971);
or U13909 (N_13909,N_11487,N_11007);
nor U13910 (N_13910,N_10843,N_10925);
xnor U13911 (N_13911,N_10377,N_10557);
nand U13912 (N_13912,N_11675,N_10268);
nor U13913 (N_13913,N_11518,N_11651);
and U13914 (N_13914,N_11191,N_10717);
and U13915 (N_13915,N_11040,N_11161);
xnor U13916 (N_13916,N_10588,N_11827);
nand U13917 (N_13917,N_10361,N_11561);
nor U13918 (N_13918,N_10613,N_10549);
xor U13919 (N_13919,N_10593,N_10412);
and U13920 (N_13920,N_11202,N_11056);
nand U13921 (N_13921,N_10980,N_10900);
or U13922 (N_13922,N_11915,N_10865);
or U13923 (N_13923,N_10229,N_11764);
nand U13924 (N_13924,N_10696,N_11865);
xor U13925 (N_13925,N_10399,N_11990);
and U13926 (N_13926,N_11156,N_10509);
and U13927 (N_13927,N_10936,N_11411);
or U13928 (N_13928,N_11438,N_10037);
nand U13929 (N_13929,N_10454,N_10782);
xor U13930 (N_13930,N_10781,N_10428);
nor U13931 (N_13931,N_11325,N_11288);
or U13932 (N_13932,N_11858,N_10527);
or U13933 (N_13933,N_11244,N_11170);
and U13934 (N_13934,N_11477,N_11863);
or U13935 (N_13935,N_10669,N_11864);
or U13936 (N_13936,N_10035,N_10962);
and U13937 (N_13937,N_10348,N_11478);
nand U13938 (N_13938,N_10198,N_11302);
xor U13939 (N_13939,N_10224,N_11795);
or U13940 (N_13940,N_11251,N_11033);
and U13941 (N_13941,N_11855,N_10939);
nand U13942 (N_13942,N_10319,N_10591);
xor U13943 (N_13943,N_10338,N_10478);
or U13944 (N_13944,N_11142,N_11516);
nand U13945 (N_13945,N_10159,N_10959);
xor U13946 (N_13946,N_11609,N_10940);
or U13947 (N_13947,N_11175,N_11246);
or U13948 (N_13948,N_11960,N_11637);
or U13949 (N_13949,N_11894,N_10070);
nor U13950 (N_13950,N_11677,N_10376);
or U13951 (N_13951,N_10287,N_10587);
nor U13952 (N_13952,N_11668,N_11384);
xnor U13953 (N_13953,N_11993,N_11041);
nand U13954 (N_13954,N_11533,N_10374);
nand U13955 (N_13955,N_10112,N_11484);
nor U13956 (N_13956,N_10454,N_11749);
and U13957 (N_13957,N_11312,N_11010);
or U13958 (N_13958,N_10350,N_10169);
or U13959 (N_13959,N_11216,N_11419);
nor U13960 (N_13960,N_10386,N_10354);
or U13961 (N_13961,N_10148,N_11159);
nor U13962 (N_13962,N_11616,N_10604);
or U13963 (N_13963,N_11899,N_10631);
nand U13964 (N_13964,N_10798,N_10705);
nand U13965 (N_13965,N_10782,N_10858);
nor U13966 (N_13966,N_11923,N_11059);
or U13967 (N_13967,N_10099,N_10766);
nand U13968 (N_13968,N_11952,N_10645);
nor U13969 (N_13969,N_10979,N_10208);
xor U13970 (N_13970,N_10500,N_10527);
nand U13971 (N_13971,N_10726,N_11644);
and U13972 (N_13972,N_11815,N_10761);
and U13973 (N_13973,N_10115,N_10875);
and U13974 (N_13974,N_11160,N_10782);
or U13975 (N_13975,N_11046,N_10607);
or U13976 (N_13976,N_11901,N_10094);
or U13977 (N_13977,N_10051,N_10590);
nand U13978 (N_13978,N_11411,N_11369);
or U13979 (N_13979,N_11884,N_11637);
xnor U13980 (N_13980,N_11189,N_11707);
nand U13981 (N_13981,N_10830,N_10606);
or U13982 (N_13982,N_10560,N_10123);
and U13983 (N_13983,N_10441,N_11811);
nor U13984 (N_13984,N_11340,N_11888);
xor U13985 (N_13985,N_10759,N_11234);
nor U13986 (N_13986,N_11614,N_10545);
nand U13987 (N_13987,N_11547,N_11436);
nor U13988 (N_13988,N_10020,N_10607);
xor U13989 (N_13989,N_11097,N_11244);
nor U13990 (N_13990,N_10660,N_10685);
and U13991 (N_13991,N_11900,N_11117);
and U13992 (N_13992,N_10018,N_10778);
nor U13993 (N_13993,N_11783,N_10190);
nor U13994 (N_13994,N_11802,N_11622);
xor U13995 (N_13995,N_11585,N_10898);
xnor U13996 (N_13996,N_11528,N_11596);
xnor U13997 (N_13997,N_10676,N_10873);
or U13998 (N_13998,N_10925,N_10162);
nor U13999 (N_13999,N_10285,N_11493);
nor U14000 (N_14000,N_13842,N_12240);
and U14001 (N_14001,N_13172,N_13581);
nor U14002 (N_14002,N_13052,N_13532);
or U14003 (N_14003,N_12319,N_12654);
nand U14004 (N_14004,N_13942,N_13112);
nand U14005 (N_14005,N_12115,N_12710);
or U14006 (N_14006,N_12127,N_12216);
and U14007 (N_14007,N_13086,N_13839);
xor U14008 (N_14008,N_12904,N_13654);
xor U14009 (N_14009,N_12510,N_12041);
or U14010 (N_14010,N_12967,N_13117);
nor U14011 (N_14011,N_13108,N_12593);
nand U14012 (N_14012,N_12984,N_12065);
nor U14013 (N_14013,N_13412,N_12946);
nand U14014 (N_14014,N_12006,N_13167);
nand U14015 (N_14015,N_12440,N_13500);
nor U14016 (N_14016,N_12947,N_12188);
xor U14017 (N_14017,N_12378,N_13012);
or U14018 (N_14018,N_12540,N_12467);
and U14019 (N_14019,N_12524,N_13717);
or U14020 (N_14020,N_12345,N_12857);
nor U14021 (N_14021,N_12701,N_13480);
nor U14022 (N_14022,N_13189,N_12886);
and U14023 (N_14023,N_13276,N_12563);
xnor U14024 (N_14024,N_13763,N_12075);
and U14025 (N_14025,N_13390,N_12082);
xnor U14026 (N_14026,N_13036,N_12343);
xnor U14027 (N_14027,N_13026,N_13337);
and U14028 (N_14028,N_13280,N_13099);
nor U14029 (N_14029,N_12841,N_13999);
xnor U14030 (N_14030,N_12254,N_13622);
xnor U14031 (N_14031,N_13956,N_13905);
nand U14032 (N_14032,N_12097,N_12965);
and U14033 (N_14033,N_12085,N_13491);
or U14034 (N_14034,N_13241,N_13268);
nand U14035 (N_14035,N_13639,N_13409);
or U14036 (N_14036,N_12511,N_12724);
or U14037 (N_14037,N_12474,N_13510);
and U14038 (N_14038,N_13650,N_13104);
nor U14039 (N_14039,N_13297,N_13512);
or U14040 (N_14040,N_12777,N_13073);
nor U14041 (N_14041,N_12641,N_13661);
nand U14042 (N_14042,N_13809,N_13105);
and U14043 (N_14043,N_12611,N_13525);
nand U14044 (N_14044,N_13695,N_12410);
and U14045 (N_14045,N_12809,N_13102);
and U14046 (N_14046,N_13439,N_12741);
or U14047 (N_14047,N_12294,N_12035);
and U14048 (N_14048,N_12738,N_13185);
nand U14049 (N_14049,N_13752,N_12719);
nor U14050 (N_14050,N_12036,N_12770);
nand U14051 (N_14051,N_13747,N_13699);
xor U14052 (N_14052,N_12288,N_13203);
xor U14053 (N_14053,N_13386,N_13147);
xor U14054 (N_14054,N_12346,N_13827);
xor U14055 (N_14055,N_12480,N_13056);
or U14056 (N_14056,N_13642,N_13188);
or U14057 (N_14057,N_13298,N_13119);
or U14058 (N_14058,N_12399,N_13255);
and U14059 (N_14059,N_13804,N_13240);
nand U14060 (N_14060,N_12373,N_13085);
nor U14061 (N_14061,N_13092,N_13933);
nand U14062 (N_14062,N_13126,N_12726);
and U14063 (N_14063,N_12771,N_13230);
and U14064 (N_14064,N_13600,N_12183);
nor U14065 (N_14065,N_13380,N_13209);
xor U14066 (N_14066,N_13150,N_12455);
and U14067 (N_14067,N_12964,N_13447);
or U14068 (N_14068,N_13305,N_13611);
nand U14069 (N_14069,N_13045,N_12772);
xnor U14070 (N_14070,N_13178,N_12019);
nor U14071 (N_14071,N_12321,N_13693);
and U14072 (N_14072,N_13708,N_12312);
or U14073 (N_14073,N_12368,N_13775);
nor U14074 (N_14074,N_13862,N_12223);
or U14075 (N_14075,N_12181,N_13617);
or U14076 (N_14076,N_12887,N_13633);
nand U14077 (N_14077,N_12761,N_13379);
xor U14078 (N_14078,N_12478,N_13474);
xnor U14079 (N_14079,N_12443,N_12674);
or U14080 (N_14080,N_12987,N_13811);
and U14081 (N_14081,N_13536,N_13858);
xnor U14082 (N_14082,N_12490,N_12644);
nor U14083 (N_14083,N_13646,N_13992);
nor U14084 (N_14084,N_13553,N_13274);
xor U14085 (N_14085,N_12049,N_13151);
nand U14086 (N_14086,N_13488,N_12898);
xnor U14087 (N_14087,N_13433,N_12918);
xnor U14088 (N_14088,N_13455,N_12460);
xor U14089 (N_14089,N_12270,N_13829);
and U14090 (N_14090,N_12465,N_12083);
and U14091 (N_14091,N_13743,N_12689);
nor U14092 (N_14092,N_12406,N_13967);
or U14093 (N_14093,N_13397,N_13417);
xor U14094 (N_14094,N_13391,N_12598);
nand U14095 (N_14095,N_12118,N_13795);
nand U14096 (N_14096,N_13173,N_13736);
xnor U14097 (N_14097,N_12371,N_12140);
and U14098 (N_14098,N_12512,N_13023);
nand U14099 (N_14099,N_12204,N_12028);
nand U14100 (N_14100,N_13060,N_13954);
and U14101 (N_14101,N_12193,N_13413);
nand U14102 (N_14102,N_13183,N_12434);
xnor U14103 (N_14103,N_13937,N_12499);
xor U14104 (N_14104,N_13801,N_12381);
xor U14105 (N_14105,N_12506,N_13777);
nor U14106 (N_14106,N_12925,N_13363);
nor U14107 (N_14107,N_12583,N_13050);
or U14108 (N_14108,N_12736,N_12929);
or U14109 (N_14109,N_13979,N_13278);
nor U14110 (N_14110,N_12757,N_13601);
nand U14111 (N_14111,N_13849,N_13725);
and U14112 (N_14112,N_13113,N_13761);
nand U14113 (N_14113,N_12937,N_13078);
nand U14114 (N_14114,N_12386,N_12235);
and U14115 (N_14115,N_12200,N_12859);
nand U14116 (N_14116,N_13746,N_12832);
nor U14117 (N_14117,N_12128,N_13182);
xnor U14118 (N_14118,N_12180,N_12136);
nor U14119 (N_14119,N_13103,N_13984);
and U14120 (N_14120,N_12673,N_12495);
nand U14121 (N_14121,N_12392,N_13832);
nand U14122 (N_14122,N_13095,N_12520);
nand U14123 (N_14123,N_12034,N_13121);
and U14124 (N_14124,N_13475,N_12778);
nor U14125 (N_14125,N_12069,N_13507);
or U14126 (N_14126,N_12975,N_12768);
and U14127 (N_14127,N_13263,N_13015);
or U14128 (N_14128,N_13533,N_12628);
nand U14129 (N_14129,N_12620,N_13081);
nand U14130 (N_14130,N_13591,N_13783);
and U14131 (N_14131,N_12500,N_12135);
or U14132 (N_14132,N_12941,N_13909);
and U14133 (N_14133,N_13790,N_13406);
xor U14134 (N_14134,N_13576,N_13587);
nor U14135 (N_14135,N_12693,N_13681);
nand U14136 (N_14136,N_12040,N_12309);
or U14137 (N_14137,N_13088,N_12218);
and U14138 (N_14138,N_12954,N_13816);
or U14139 (N_14139,N_12414,N_12201);
nor U14140 (N_14140,N_13302,N_12942);
xnor U14141 (N_14141,N_12126,N_12527);
or U14142 (N_14142,N_13155,N_13245);
nand U14143 (N_14143,N_12195,N_12285);
nor U14144 (N_14144,N_13978,N_12403);
or U14145 (N_14145,N_12023,N_12291);
xor U14146 (N_14146,N_13653,N_12978);
or U14147 (N_14147,N_12293,N_12372);
or U14148 (N_14148,N_13649,N_13850);
or U14149 (N_14149,N_12461,N_12005);
nor U14150 (N_14150,N_13722,N_12472);
nand U14151 (N_14151,N_12518,N_12086);
xor U14152 (N_14152,N_12427,N_13669);
or U14153 (N_14153,N_12990,N_13010);
nand U14154 (N_14154,N_12882,N_12281);
and U14155 (N_14155,N_13888,N_12554);
xor U14156 (N_14156,N_12526,N_12928);
and U14157 (N_14157,N_13058,N_12073);
or U14158 (N_14158,N_12926,N_12544);
xor U14159 (N_14159,N_13421,N_13028);
and U14160 (N_14160,N_12170,N_12477);
nor U14161 (N_14161,N_13213,N_12376);
xor U14162 (N_14162,N_13200,N_12679);
or U14163 (N_14163,N_12426,N_13382);
and U14164 (N_14164,N_12418,N_13748);
nand U14165 (N_14165,N_12740,N_13079);
nor U14166 (N_14166,N_13547,N_12144);
xnor U14167 (N_14167,N_12446,N_13062);
xor U14168 (N_14168,N_13089,N_13440);
nor U14169 (N_14169,N_13392,N_12709);
and U14170 (N_14170,N_13469,N_12564);
nor U14171 (N_14171,N_12432,N_12915);
nor U14172 (N_14172,N_13146,N_13574);
or U14173 (N_14173,N_12924,N_13176);
nor U14174 (N_14174,N_12971,N_13335);
xor U14175 (N_14175,N_13877,N_13466);
nor U14176 (N_14176,N_13282,N_12380);
or U14177 (N_14177,N_12631,N_12447);
xor U14178 (N_14178,N_12154,N_12962);
nor U14179 (N_14179,N_12442,N_13358);
or U14180 (N_14180,N_12423,N_13934);
and U14181 (N_14181,N_12542,N_13890);
and U14182 (N_14182,N_13915,N_13950);
nand U14183 (N_14183,N_13420,N_13524);
xnor U14184 (N_14184,N_12879,N_12058);
xnor U14185 (N_14185,N_12529,N_13714);
nand U14186 (N_14186,N_12634,N_12791);
nor U14187 (N_14187,N_12858,N_13879);
or U14188 (N_14188,N_12063,N_13446);
or U14189 (N_14189,N_12237,N_12643);
or U14190 (N_14190,N_12732,N_12341);
xor U14191 (N_14191,N_13604,N_13061);
and U14192 (N_14192,N_12746,N_12627);
nor U14193 (N_14193,N_13840,N_12064);
xnor U14194 (N_14194,N_13891,N_12923);
nor U14195 (N_14195,N_12864,N_12896);
xor U14196 (N_14196,N_12800,N_13552);
nor U14197 (N_14197,N_13368,N_13364);
nand U14198 (N_14198,N_13257,N_12002);
xor U14199 (N_14199,N_12823,N_13628);
xor U14200 (N_14200,N_13039,N_13407);
nand U14201 (N_14201,N_13575,N_13786);
xnor U14202 (N_14202,N_13424,N_12256);
or U14203 (N_14203,N_12754,N_12448);
xor U14204 (N_14204,N_12286,N_13142);
or U14205 (N_14205,N_12586,N_13830);
xor U14206 (N_14206,N_13442,N_13157);
nor U14207 (N_14207,N_13757,N_13353);
and U14208 (N_14208,N_13265,N_12642);
nand U14209 (N_14209,N_13139,N_13878);
nand U14210 (N_14210,N_12919,N_12071);
nand U14211 (N_14211,N_13797,N_13366);
or U14212 (N_14212,N_12534,N_12578);
xor U14213 (N_14213,N_13679,N_13375);
nor U14214 (N_14214,N_13031,N_13145);
or U14215 (N_14215,N_12671,N_13111);
nand U14216 (N_14216,N_12050,N_12938);
nand U14217 (N_14217,N_13917,N_12483);
and U14218 (N_14218,N_13460,N_12438);
nor U14219 (N_14219,N_13875,N_13149);
nor U14220 (N_14220,N_13707,N_13501);
nor U14221 (N_14221,N_12007,N_12272);
xnor U14222 (N_14222,N_12959,N_13378);
nand U14223 (N_14223,N_13426,N_13626);
and U14224 (N_14224,N_12375,N_12197);
nand U14225 (N_14225,N_12481,N_12314);
xor U14226 (N_14226,N_13516,N_13819);
and U14227 (N_14227,N_12782,N_12001);
nor U14228 (N_14228,N_12025,N_13499);
or U14229 (N_14229,N_12769,N_13206);
nor U14230 (N_14230,N_13994,N_13896);
or U14231 (N_14231,N_13311,N_13349);
or U14232 (N_14232,N_13310,N_12377);
xor U14233 (N_14233,N_13494,N_13193);
or U14234 (N_14234,N_12514,N_12352);
or U14235 (N_14235,N_13238,N_12382);
nand U14236 (N_14236,N_12979,N_12908);
or U14237 (N_14237,N_12102,N_13037);
xnor U14238 (N_14238,N_13360,N_12704);
and U14239 (N_14239,N_13481,N_12817);
or U14240 (N_14240,N_13027,N_13168);
xnor U14241 (N_14241,N_12484,N_12226);
nand U14242 (N_14242,N_13486,N_12548);
and U14243 (N_14243,N_13670,N_13067);
xor U14244 (N_14244,N_12988,N_13548);
or U14245 (N_14245,N_13005,N_13207);
or U14246 (N_14246,N_12525,N_12420);
nor U14247 (N_14247,N_12556,N_12715);
nand U14248 (N_14248,N_12119,N_13696);
and U14249 (N_14249,N_12501,N_13734);
or U14250 (N_14250,N_12716,N_13541);
xnor U14251 (N_14251,N_12825,N_13244);
nor U14252 (N_14252,N_13662,N_12277);
nor U14253 (N_14253,N_12466,N_12998);
and U14254 (N_14254,N_12282,N_13874);
or U14255 (N_14255,N_12523,N_12072);
xnor U14256 (N_14256,N_13952,N_13509);
nor U14257 (N_14257,N_12977,N_13610);
nand U14258 (N_14258,N_12950,N_12462);
xor U14259 (N_14259,N_13980,N_13222);
or U14260 (N_14260,N_13082,N_12935);
nand U14261 (N_14261,N_13721,N_12911);
xor U14262 (N_14262,N_12310,N_13171);
or U14263 (N_14263,N_13973,N_13640);
xor U14264 (N_14264,N_13431,N_12151);
nand U14265 (N_14265,N_12703,N_13443);
nor U14266 (N_14266,N_12271,N_12122);
or U14267 (N_14267,N_12883,N_12081);
nand U14268 (N_14268,N_12493,N_13289);
and U14269 (N_14269,N_13822,N_13330);
nand U14270 (N_14270,N_12785,N_12878);
or U14271 (N_14271,N_13573,N_13846);
and U14272 (N_14272,N_12225,N_13427);
nor U14273 (N_14273,N_13419,N_13718);
and U14274 (N_14274,N_12812,N_12795);
or U14275 (N_14275,N_12055,N_12516);
nor U14276 (N_14276,N_13434,N_13051);
and U14277 (N_14277,N_12194,N_12905);
nand U14278 (N_14278,N_13982,N_13715);
nand U14279 (N_14279,N_13961,N_12565);
and U14280 (N_14280,N_12498,N_13165);
nor U14281 (N_14281,N_12186,N_12596);
xnor U14282 (N_14282,N_12632,N_12212);
and U14283 (N_14283,N_13348,N_13989);
xor U14284 (N_14284,N_13986,N_12155);
or U14285 (N_14285,N_12960,N_13011);
nor U14286 (N_14286,N_13926,N_13549);
nand U14287 (N_14287,N_12362,N_12318);
nor U14288 (N_14288,N_13866,N_12305);
or U14289 (N_14289,N_13234,N_12617);
xor U14290 (N_14290,N_12874,N_13071);
nor U14291 (N_14291,N_13910,N_13258);
nand U14292 (N_14292,N_13338,N_13690);
xor U14293 (N_14293,N_13281,N_13000);
and U14294 (N_14294,N_13665,N_13457);
xnor U14295 (N_14295,N_12968,N_12259);
nand U14296 (N_14296,N_12255,N_12422);
or U14297 (N_14297,N_12624,N_13958);
nand U14298 (N_14298,N_13400,N_12684);
xnor U14299 (N_14299,N_13678,N_12742);
xor U14300 (N_14300,N_13588,N_12835);
nand U14301 (N_14301,N_12297,N_13347);
or U14302 (N_14302,N_12330,N_13847);
and U14303 (N_14303,N_13564,N_12391);
xor U14304 (N_14304,N_13876,N_12022);
xor U14305 (N_14305,N_13396,N_12012);
xnor U14306 (N_14306,N_13658,N_12158);
xor U14307 (N_14307,N_13381,N_13100);
nor U14308 (N_14308,N_13769,N_13365);
and U14309 (N_14309,N_13566,N_12338);
and U14310 (N_14310,N_12798,N_13064);
nand U14311 (N_14311,N_12553,N_12672);
xnor U14312 (N_14312,N_12405,N_13737);
nor U14313 (N_14313,N_13318,N_12149);
and U14314 (N_14314,N_13966,N_12325);
or U14315 (N_14315,N_13550,N_12452);
nor U14316 (N_14316,N_13852,N_12413);
nand U14317 (N_14317,N_12326,N_12080);
or U14318 (N_14318,N_13492,N_13158);
or U14319 (N_14319,N_13329,N_13461);
xnor U14320 (N_14320,N_13343,N_12751);
xnor U14321 (N_14321,N_13114,N_13503);
nor U14322 (N_14322,N_12045,N_13941);
or U14323 (N_14323,N_12897,N_13191);
nor U14324 (N_14324,N_12360,N_12209);
nor U14325 (N_14325,N_12892,N_13186);
nor U14326 (N_14326,N_12171,N_13024);
nor U14327 (N_14327,N_12630,N_12052);
xor U14328 (N_14328,N_13354,N_13767);
xnor U14329 (N_14329,N_13868,N_13927);
nor U14330 (N_14330,N_13881,N_13456);
nor U14331 (N_14331,N_12206,N_12513);
xor U14332 (N_14332,N_13136,N_13243);
nand U14333 (N_14333,N_13159,N_12130);
and U14334 (N_14334,N_12993,N_13672);
or U14335 (N_14335,N_13865,N_13470);
and U14336 (N_14336,N_12192,N_12875);
nand U14337 (N_14337,N_13416,N_12914);
xnor U14338 (N_14338,N_12311,N_13843);
or U14339 (N_14339,N_13402,N_13798);
and U14340 (N_14340,N_12011,N_12856);
nand U14341 (N_14341,N_13166,N_12284);
nor U14342 (N_14342,N_12349,N_12232);
xnor U14343 (N_14343,N_13700,N_12304);
nand U14344 (N_14344,N_13569,N_12436);
or U14345 (N_14345,N_12390,N_13704);
nor U14346 (N_14346,N_12789,N_12334);
or U14347 (N_14347,N_12503,N_13703);
nor U14348 (N_14348,N_12801,N_13740);
nor U14349 (N_14349,N_13997,N_13387);
or U14350 (N_14350,N_13657,N_12449);
xor U14351 (N_14351,N_13556,N_13428);
or U14352 (N_14352,N_13049,N_13249);
nand U14353 (N_14353,N_13070,N_13815);
or U14354 (N_14354,N_13648,N_12845);
xor U14355 (N_14355,N_13647,N_12657);
or U14356 (N_14356,N_12107,N_12737);
nor U14357 (N_14357,N_13560,N_12894);
nand U14358 (N_14358,N_13643,N_13351);
nor U14359 (N_14359,N_12120,N_13083);
or U14360 (N_14360,N_12532,N_13948);
nand U14361 (N_14361,N_12515,N_12780);
or U14362 (N_14362,N_12502,N_12307);
nand U14363 (N_14363,N_13451,N_13749);
nand U14364 (N_14364,N_12273,N_13283);
or U14365 (N_14365,N_12039,N_12916);
nor U14366 (N_14366,N_13559,N_12543);
nand U14367 (N_14367,N_12541,N_13259);
and U14368 (N_14368,N_13730,N_13663);
and U14369 (N_14369,N_12331,N_12669);
nand U14370 (N_14370,N_13291,N_12214);
and U14371 (N_14371,N_12221,N_12091);
and U14372 (N_14372,N_12488,N_12054);
nor U14373 (N_14373,N_12880,N_12504);
nand U14374 (N_14374,N_13945,N_12779);
nand U14375 (N_14375,N_13220,N_13030);
nor U14376 (N_14376,N_13435,N_12702);
xnor U14377 (N_14377,N_12607,N_12820);
or U14378 (N_14378,N_13701,N_12354);
nor U14379 (N_14379,N_13898,N_13618);
xnor U14380 (N_14380,N_12755,N_13912);
or U14381 (N_14381,N_12339,N_13562);
or U14382 (N_14382,N_13163,N_12230);
nor U14383 (N_14383,N_12622,N_13996);
and U14384 (N_14384,N_13543,N_12748);
and U14385 (N_14385,N_12681,N_12995);
or U14386 (N_14386,N_13233,N_12656);
and U14387 (N_14387,N_12215,N_13963);
xnor U14388 (N_14388,N_12698,N_12165);
nor U14389 (N_14389,N_13317,N_13346);
nor U14390 (N_14390,N_13399,N_12393);
or U14391 (N_14391,N_13022,N_12639);
and U14392 (N_14392,N_13921,N_13627);
xnor U14393 (N_14393,N_13528,N_12729);
nor U14394 (N_14394,N_12295,N_12930);
nor U14395 (N_14395,N_13886,N_12148);
nand U14396 (N_14396,N_12290,N_13659);
xor U14397 (N_14397,N_13441,N_12412);
and U14398 (N_14398,N_12601,N_13579);
xor U14399 (N_14399,N_12246,N_13892);
nor U14400 (N_14400,N_12976,N_13334);
nand U14401 (N_14401,N_12138,N_12792);
xor U14402 (N_14402,N_12750,N_13928);
nor U14403 (N_14403,N_13674,N_12863);
and U14404 (N_14404,N_12603,N_13870);
or U14405 (N_14405,N_13393,N_12332);
nor U14406 (N_14406,N_13116,N_12621);
xor U14407 (N_14407,N_13629,N_12098);
and U14408 (N_14408,N_13632,N_12991);
nand U14409 (N_14409,N_13059,N_12612);
nor U14410 (N_14410,N_13813,N_12227);
and U14411 (N_14411,N_13991,N_12558);
nand U14412 (N_14412,N_13808,N_13975);
xnor U14413 (N_14413,N_13765,N_12353);
or U14414 (N_14414,N_13517,N_13256);
and U14415 (N_14415,N_12067,N_13152);
nand U14416 (N_14416,N_13773,N_13925);
or U14417 (N_14417,N_13977,N_13586);
or U14418 (N_14418,N_12152,N_13987);
and U14419 (N_14419,N_13389,N_12927);
nand U14420 (N_14420,N_12912,N_13493);
nor U14421 (N_14421,N_13606,N_13333);
and U14422 (N_14422,N_12999,N_12059);
nor U14423 (N_14423,N_12431,N_12647);
and U14424 (N_14424,N_13615,N_12308);
nor U14425 (N_14425,N_13459,N_13593);
xor U14426 (N_14426,N_13356,N_12257);
or U14427 (N_14427,N_12057,N_12853);
and U14428 (N_14428,N_13504,N_12891);
nand U14429 (N_14429,N_12335,N_12666);
nor U14430 (N_14430,N_12722,N_13831);
nor U14431 (N_14431,N_12804,N_12574);
and U14432 (N_14432,N_13527,N_12106);
or U14433 (N_14433,N_12134,N_12616);
xnor U14434 (N_14434,N_12132,N_12619);
xor U14435 (N_14435,N_12653,N_12569);
xnor U14436 (N_14436,N_13160,N_13571);
and U14437 (N_14437,N_12871,N_12096);
nand U14438 (N_14438,N_13228,N_13855);
or U14439 (N_14439,N_12608,N_13901);
nor U14440 (N_14440,N_12184,N_12579);
nor U14441 (N_14441,N_12383,N_12707);
xor U14442 (N_14442,N_13132,N_13101);
xor U14443 (N_14443,N_13612,N_12571);
and U14444 (N_14444,N_13357,N_12557);
xor U14445 (N_14445,N_12117,N_13034);
and U14446 (N_14446,N_13841,N_13713);
or U14447 (N_14447,N_13140,N_12141);
and U14448 (N_14448,N_12670,N_12017);
nand U14449 (N_14449,N_12150,N_13780);
and U14450 (N_14450,N_13472,N_12773);
or U14451 (N_14451,N_13482,N_12159);
nor U14452 (N_14452,N_13902,N_13692);
xor U14453 (N_14453,N_12267,N_12580);
and U14454 (N_14454,N_12783,N_12730);
nor U14455 (N_14455,N_13807,N_12944);
xor U14456 (N_14456,N_13208,N_12907);
nor U14457 (N_14457,N_13211,N_12568);
and U14458 (N_14458,N_12744,N_12087);
nor U14459 (N_14459,N_12996,N_12328);
or U14460 (N_14460,N_13520,N_13107);
nor U14461 (N_14461,N_13995,N_12796);
or U14462 (N_14462,N_13403,N_13570);
or U14463 (N_14463,N_12459,N_12476);
or U14464 (N_14464,N_12862,N_13754);
xnor U14465 (N_14465,N_13742,N_13479);
nand U14466 (N_14466,N_12760,N_13511);
and U14467 (N_14467,N_12992,N_12357);
or U14468 (N_14468,N_13820,N_12695);
xor U14469 (N_14469,N_13723,N_12348);
xnor U14470 (N_14470,N_12044,N_13667);
nand U14471 (N_14471,N_12298,N_12686);
nor U14472 (N_14472,N_13959,N_12970);
xnor U14473 (N_14473,N_12655,N_13306);
xor U14474 (N_14474,N_13044,N_12487);
nand U14475 (N_14475,N_13949,N_12873);
and U14476 (N_14476,N_12444,N_12337);
and U14477 (N_14477,N_13733,N_12419);
nor U14478 (N_14478,N_13294,N_12890);
nand U14479 (N_14479,N_13731,N_13080);
nor U14480 (N_14480,N_12169,N_12109);
and U14481 (N_14481,N_13554,N_12112);
and U14482 (N_14482,N_12092,N_12070);
or U14483 (N_14483,N_12660,N_13792);
nor U14484 (N_14484,N_12408,N_12932);
nand U14485 (N_14485,N_12893,N_13194);
or U14486 (N_14486,N_12191,N_13201);
xnor U14487 (N_14487,N_13181,N_13017);
and U14488 (N_14488,N_13998,N_13624);
nand U14489 (N_14489,N_13018,N_13432);
nand U14490 (N_14490,N_12706,N_12471);
or U14491 (N_14491,N_13753,N_13857);
nand U14492 (N_14492,N_13098,N_12901);
nor U14493 (N_14493,N_13938,N_12302);
xnor U14494 (N_14494,N_12433,N_13066);
or U14495 (N_14495,N_12983,N_12803);
xor U14496 (N_14496,N_12179,N_12217);
nor U14497 (N_14497,N_12592,N_13584);
and U14498 (N_14498,N_13859,N_12060);
nand U14499 (N_14499,N_13613,N_12366);
xnor U14500 (N_14500,N_13502,N_12688);
or U14501 (N_14501,N_13248,N_13597);
nor U14502 (N_14502,N_12198,N_13534);
xor U14503 (N_14503,N_13833,N_13197);
nor U14504 (N_14504,N_13677,N_12156);
nor U14505 (N_14505,N_13008,N_13918);
nand U14506 (N_14506,N_12089,N_13214);
or U14507 (N_14507,N_12280,N_12238);
xor U14508 (N_14508,N_13908,N_12199);
nand U14509 (N_14509,N_13582,N_12489);
and U14510 (N_14510,N_12735,N_13621);
and U14511 (N_14511,N_13376,N_13710);
nand U14512 (N_14512,N_13776,N_13580);
nor U14513 (N_14513,N_12986,N_12807);
xor U14514 (N_14514,N_12416,N_12113);
nor U14515 (N_14515,N_12989,N_12486);
xor U14516 (N_14516,N_13838,N_12590);
or U14517 (N_14517,N_13602,N_13694);
and U14518 (N_14518,N_13932,N_13887);
xnor U14519 (N_14519,N_13539,N_13063);
nand U14520 (N_14520,N_12635,N_12178);
or U14521 (N_14521,N_12651,N_13720);
nor U14522 (N_14522,N_13477,N_12275);
and U14523 (N_14523,N_12105,N_13020);
or U14524 (N_14524,N_13545,N_13530);
xor U14525 (N_14525,N_12177,N_13706);
nand U14526 (N_14526,N_12680,N_13712);
nor U14527 (N_14527,N_12766,N_13322);
and U14528 (N_14528,N_13002,N_12143);
and U14529 (N_14529,N_12394,N_12561);
xnor U14530 (N_14530,N_13180,N_13096);
or U14531 (N_14531,N_12865,N_12682);
or U14532 (N_14532,N_12145,N_12242);
nor U14533 (N_14533,N_13895,N_13880);
or U14534 (N_14534,N_13930,N_13968);
and U14535 (N_14535,N_13762,N_12854);
nand U14536 (N_14536,N_13065,N_12129);
nor U14537 (N_14537,N_12969,N_13048);
and U14538 (N_14538,N_13906,N_13686);
or U14539 (N_14539,N_12450,N_13885);
nand U14540 (N_14540,N_12327,N_13490);
or U14541 (N_14541,N_12324,N_12015);
and U14542 (N_14542,N_12313,N_12668);
xor U14543 (N_14543,N_13785,N_13883);
nand U14544 (N_14544,N_13135,N_13485);
or U14545 (N_14545,N_13212,N_13009);
nor U14546 (N_14546,N_13914,N_12885);
nand U14547 (N_14547,N_12699,N_13423);
nand U14548 (N_14548,N_12231,N_13589);
or U14549 (N_14549,N_12837,N_13625);
and U14550 (N_14550,N_12125,N_12551);
and U14551 (N_14551,N_12016,N_12537);
and U14552 (N_14552,N_13242,N_13131);
nor U14553 (N_14553,N_13312,N_12224);
nand U14554 (N_14554,N_12815,N_13097);
nor U14555 (N_14555,N_12457,N_13907);
nand U14556 (N_14556,N_12676,N_12110);
xor U14557 (N_14557,N_13745,N_12061);
or U14558 (N_14558,N_12776,N_13137);
or U14559 (N_14559,N_12479,N_12265);
or U14560 (N_14560,N_13544,N_13250);
nand U14561 (N_14561,N_12861,N_13483);
nand U14562 (N_14562,N_13093,N_12734);
and U14563 (N_14563,N_13035,N_12278);
or U14564 (N_14564,N_13043,N_13755);
nor U14565 (N_14565,N_13319,N_12078);
xor U14566 (N_14566,N_13174,N_13266);
and U14567 (N_14567,N_13215,N_12831);
nand U14568 (N_14568,N_12855,N_13156);
nand U14569 (N_14569,N_13361,N_13538);
nand U14570 (N_14570,N_12222,N_13947);
xnor U14571 (N_14571,N_13372,N_12395);
or U14572 (N_14572,N_13960,N_13109);
nand U14573 (N_14573,N_12210,N_12981);
xnor U14574 (N_14574,N_12010,N_13519);
nor U14575 (N_14575,N_12340,N_13636);
xnor U14576 (N_14576,N_13771,N_13796);
xor U14577 (N_14577,N_12625,N_12765);
nand U14578 (N_14578,N_12301,N_13143);
and U14579 (N_14579,N_13592,N_13429);
and U14580 (N_14580,N_13025,N_12691);
or U14581 (N_14581,N_13448,N_13826);
or U14582 (N_14582,N_12220,N_13974);
or U14583 (N_14583,N_12767,N_13084);
nor U14584 (N_14584,N_13897,N_12665);
nand U14585 (N_14585,N_12629,N_12658);
and U14586 (N_14586,N_13635,N_12714);
nand U14587 (N_14587,N_13837,N_13729);
and U14588 (N_14588,N_13869,N_12095);
nor U14589 (N_14589,N_13936,N_12725);
or U14590 (N_14590,N_13410,N_12234);
or U14591 (N_14591,N_13969,N_13408);
nand U14592 (N_14592,N_13106,N_12902);
and U14593 (N_14593,N_13972,N_12638);
nand U14594 (N_14594,N_13922,N_12453);
xnor U14595 (N_14595,N_12424,N_12175);
xor U14596 (N_14596,N_12300,N_12961);
xnor U14597 (N_14597,N_12196,N_13835);
and U14598 (N_14598,N_12404,N_12781);
nand U14599 (N_14599,N_13284,N_12043);
and U14600 (N_14600,N_12866,N_12811);
nor U14601 (N_14601,N_13976,N_13515);
or U14602 (N_14602,N_12843,N_13342);
xor U14603 (N_14603,N_12369,N_12633);
xor U14604 (N_14604,N_12650,N_12547);
or U14605 (N_14605,N_13793,N_13221);
nor U14606 (N_14606,N_12496,N_13645);
nand U14607 (N_14607,N_12131,N_12100);
xnor U14608 (N_14608,N_12509,N_12367);
nor U14609 (N_14609,N_12591,N_12116);
xnor U14610 (N_14610,N_12636,N_13239);
nor U14611 (N_14611,N_12920,N_12764);
or U14612 (N_14612,N_12207,N_12808);
or U14613 (N_14613,N_12958,N_13444);
or U14614 (N_14614,N_12402,N_12762);
nand U14615 (N_14615,N_12881,N_13848);
nand U14616 (N_14616,N_12475,N_12219);
nor U14617 (N_14617,N_12167,N_13732);
nor U14618 (N_14618,N_13384,N_13697);
xor U14619 (N_14619,N_12208,N_12957);
or U14620 (N_14620,N_13300,N_12463);
nor U14621 (N_14621,N_12121,N_12187);
and U14622 (N_14622,N_13634,N_13789);
or U14623 (N_14623,N_13894,N_13814);
and U14624 (N_14624,N_13198,N_12094);
xor U14625 (N_14625,N_12101,N_13616);
or U14626 (N_14626,N_12365,N_13287);
xor U14627 (N_14627,N_13675,N_13664);
xnor U14628 (N_14628,N_12640,N_13964);
or U14629 (N_14629,N_13844,N_12336);
xor U14630 (N_14630,N_12355,N_12948);
xor U14631 (N_14631,N_13046,N_13235);
or U14632 (N_14632,N_12482,N_12844);
nand U14633 (N_14633,N_13970,N_13558);
xor U14634 (N_14634,N_12939,N_13683);
nor U14635 (N_14635,N_13385,N_13555);
or U14636 (N_14636,N_12084,N_13129);
or U14637 (N_14637,N_13301,N_13518);
xor U14638 (N_14638,N_13130,N_13449);
or U14639 (N_14639,N_12868,N_12245);
xor U14640 (N_14640,N_12415,N_12731);
or U14641 (N_14641,N_12163,N_13689);
and U14642 (N_14642,N_13595,N_13016);
xnor U14643 (N_14643,N_12895,N_12696);
nand U14644 (N_14644,N_12697,N_12774);
nand U14645 (N_14645,N_12229,N_13940);
or U14646 (N_14646,N_13314,N_12980);
nand U14647 (N_14647,N_12648,N_12824);
or U14648 (N_14648,N_12316,N_13118);
xnor U14649 (N_14649,N_13398,N_12536);
and U14650 (N_14650,N_13824,N_13040);
xnor U14651 (N_14651,N_13542,N_13341);
nand U14652 (N_14652,N_12053,N_12784);
xnor U14653 (N_14653,N_12153,N_12400);
or U14654 (N_14654,N_13175,N_12922);
and U14655 (N_14655,N_13271,N_13484);
and U14656 (N_14656,N_12840,N_12146);
and U14657 (N_14657,N_12519,N_13467);
nor U14658 (N_14658,N_13851,N_12468);
or U14659 (N_14659,N_12753,N_13900);
xor U14660 (N_14660,N_12610,N_13205);
xnor U14661 (N_14661,N_12533,N_12176);
and U14662 (N_14662,N_12262,N_13567);
nand U14663 (N_14663,N_12430,N_12609);
or U14664 (N_14664,N_12877,N_12705);
and U14665 (N_14665,N_12869,N_12168);
nor U14666 (N_14666,N_12264,N_12560);
or U14667 (N_14667,N_12026,N_12745);
and U14668 (N_14668,N_13120,N_13540);
or U14669 (N_14669,N_12306,N_13531);
xor U14670 (N_14670,N_13463,N_12550);
nor U14671 (N_14671,N_13609,N_13004);
nor U14672 (N_14672,N_12123,N_13828);
and U14673 (N_14673,N_12469,N_12910);
and U14674 (N_14674,N_12661,N_13817);
and U14675 (N_14675,N_13436,N_12921);
nand U14676 (N_14676,N_12029,N_13465);
nor U14677 (N_14677,N_13585,N_13939);
nand U14678 (N_14678,N_12582,N_12142);
and U14679 (N_14679,N_13247,N_13091);
nor U14680 (N_14680,N_12909,N_12775);
nor U14681 (N_14681,N_12963,N_12985);
xor U14682 (N_14682,N_12664,N_12847);
nor U14683 (N_14683,N_12172,N_13577);
nor U14684 (N_14684,N_12974,N_13110);
or U14685 (N_14685,N_12677,N_12396);
nor U14686 (N_14686,N_13074,N_12692);
xor U14687 (N_14687,N_13273,N_13007);
nand U14688 (N_14688,N_13369,N_13931);
nor U14689 (N_14689,N_12364,N_13450);
xor U14690 (N_14690,N_13315,N_12456);
and U14691 (N_14691,N_13452,N_12949);
xnor U14692 (N_14692,N_13328,N_12303);
and U14693 (N_14693,N_13856,N_13596);
or U14694 (N_14694,N_13430,N_12236);
nor U14695 (N_14695,N_13087,N_13962);
or U14696 (N_14696,N_12623,N_13578);
xnor U14697 (N_14697,N_13836,N_12822);
or U14698 (N_14698,N_13845,N_12752);
xnor U14699 (N_14699,N_13513,N_13702);
and U14700 (N_14700,N_13668,N_13161);
and U14701 (N_14701,N_13882,N_13935);
nand U14702 (N_14702,N_12850,N_13884);
nand U14703 (N_14703,N_12690,N_12385);
or U14704 (N_14704,N_12269,N_12899);
nor U14705 (N_14705,N_12934,N_12559);
nor U14706 (N_14706,N_12802,N_12613);
nand U14707 (N_14707,N_12389,N_12763);
xnor U14708 (N_14708,N_12827,N_13818);
or U14709 (N_14709,N_12521,N_13778);
and U14710 (N_14710,N_13903,N_12649);
or U14711 (N_14711,N_13688,N_13453);
or U14712 (N_14712,N_12077,N_13770);
xnor U14713 (N_14713,N_12458,N_12570);
or U14714 (N_14714,N_13943,N_12008);
xor U14715 (N_14715,N_12683,N_13304);
or U14716 (N_14716,N_13326,N_13041);
and U14717 (N_14717,N_12370,N_12814);
or U14718 (N_14718,N_13437,N_12538);
and U14719 (N_14719,N_12268,N_12955);
nor U14720 (N_14720,N_13812,N_12090);
and U14721 (N_14721,N_13682,N_12439);
nor U14722 (N_14722,N_12494,N_13216);
nand U14723 (N_14723,N_12718,N_13651);
and U14724 (N_14724,N_13124,N_12497);
and U14725 (N_14725,N_13316,N_13803);
xnor U14726 (N_14726,N_12576,N_12972);
xnor U14727 (N_14727,N_12816,N_13231);
nand U14728 (N_14728,N_12933,N_13299);
or U14729 (N_14729,N_13473,N_13638);
or U14730 (N_14730,N_13860,N_13068);
and U14731 (N_14731,N_13802,N_13227);
and U14732 (N_14732,N_12943,N_13327);
xor U14733 (N_14733,N_13759,N_13383);
nor U14734 (N_14734,N_13537,N_13929);
nand U14735 (N_14735,N_12031,N_13806);
and U14736 (N_14736,N_13766,N_13955);
or U14737 (N_14737,N_12913,N_12797);
or U14738 (N_14738,N_12344,N_12239);
nand U14739 (N_14739,N_12758,N_13951);
or U14740 (N_14740,N_12317,N_12530);
nor U14741 (N_14741,N_13295,N_12573);
xor U14742 (N_14742,N_13462,N_12906);
or U14743 (N_14743,N_12492,N_12485);
xor U14744 (N_14744,N_13458,N_12250);
xnor U14745 (N_14745,N_13454,N_12903);
nor U14746 (N_14746,N_12411,N_12021);
or U14747 (N_14747,N_12952,N_12261);
and U14748 (N_14748,N_12333,N_13047);
nor U14749 (N_14749,N_13340,N_12846);
xor U14750 (N_14750,N_12445,N_13506);
xor U14751 (N_14751,N_13388,N_13787);
and U14752 (N_14752,N_13735,N_13029);
or U14753 (N_14753,N_13190,N_13652);
nand U14754 (N_14754,N_12435,N_13144);
or U14755 (N_14755,N_12584,N_13122);
nor U14756 (N_14756,N_13889,N_13394);
xor U14757 (N_14757,N_13496,N_13277);
nand U14758 (N_14758,N_13415,N_13006);
or U14759 (N_14759,N_13303,N_13148);
nand U14760 (N_14760,N_13904,N_12663);
nor U14761 (N_14761,N_12830,N_12838);
or U14762 (N_14762,N_12243,N_12088);
or U14763 (N_14763,N_12421,N_13853);
or U14764 (N_14764,N_13744,N_12508);
nor U14765 (N_14765,N_13799,N_12276);
nor U14766 (N_14766,N_13345,N_13127);
nand U14767 (N_14767,N_13598,N_12618);
nand U14768 (N_14768,N_12329,N_12829);
and U14769 (N_14769,N_13224,N_12739);
nor U14770 (N_14770,N_13709,N_12545);
nor U14771 (N_14771,N_12552,N_13768);
or U14772 (N_14772,N_13953,N_13003);
or U14773 (N_14773,N_13605,N_13262);
and U14774 (N_14774,N_13698,N_13021);
nand U14775 (N_14775,N_12379,N_12567);
nand U14776 (N_14776,N_12093,N_12248);
nor U14777 (N_14777,N_12042,N_13631);
nand U14778 (N_14778,N_12205,N_12805);
nand U14779 (N_14779,N_13204,N_13267);
nand U14780 (N_14780,N_12384,N_12441);
and U14781 (N_14781,N_12388,N_12733);
xnor U14782 (N_14782,N_13614,N_13561);
and U14783 (N_14783,N_12018,N_12173);
or U14784 (N_14784,N_13362,N_12675);
and U14785 (N_14785,N_13072,N_13237);
xnor U14786 (N_14786,N_13981,N_12821);
or U14787 (N_14787,N_13873,N_12687);
and U14788 (N_14788,N_12566,N_12111);
nor U14789 (N_14789,N_13464,N_12605);
and U14790 (N_14790,N_13535,N_13660);
nor U14791 (N_14791,N_13210,N_12292);
nor U14792 (N_14792,N_13115,N_13162);
and U14793 (N_14793,N_12048,N_12247);
xnor U14794 (N_14794,N_12788,N_12531);
or U14795 (N_14795,N_13422,N_13321);
and U14796 (N_14796,N_13965,N_13522);
xnor U14797 (N_14797,N_12162,N_12678);
xor U14798 (N_14798,N_13308,N_12562);
nor U14799 (N_14799,N_13055,N_13603);
xnor U14800 (N_14800,N_13285,N_12595);
nand U14801 (N_14801,N_12409,N_13924);
and U14802 (N_14802,N_12876,N_13899);
nand U14803 (N_14803,N_12581,N_12727);
nor U14804 (N_14804,N_13069,N_12315);
nor U14805 (N_14805,N_13042,N_12464);
or U14806 (N_14806,N_13716,N_13134);
nor U14807 (N_14807,N_13350,N_12546);
nor U14808 (N_14808,N_13275,N_12507);
nor U14809 (N_14809,N_12549,N_12363);
xnor U14810 (N_14810,N_13246,N_12322);
nand U14811 (N_14811,N_13325,N_13772);
xnor U14812 (N_14812,N_13551,N_12046);
xor U14813 (N_14813,N_13054,N_12037);
nand U14814 (N_14814,N_13546,N_13196);
or U14815 (N_14815,N_13764,N_12720);
or U14816 (N_14816,N_12166,N_12397);
or U14817 (N_14817,N_12032,N_13154);
nor U14818 (N_14818,N_13871,N_13565);
and U14819 (N_14819,N_12834,N_12491);
nand U14820 (N_14820,N_12712,N_12244);
and U14821 (N_14821,N_13666,N_13983);
xnor U14822 (N_14822,N_13404,N_12842);
nand U14823 (N_14823,N_13478,N_12818);
nand U14824 (N_14824,N_12700,N_12066);
and U14825 (N_14825,N_12794,N_13332);
nand U14826 (N_14826,N_13727,N_12585);
nand U14827 (N_14827,N_13352,N_13563);
or U14828 (N_14828,N_13825,N_12274);
nor U14829 (N_14829,N_13791,N_13620);
xor U14830 (N_14830,N_12685,N_12251);
xor U14831 (N_14831,N_13864,N_12667);
or U14832 (N_14832,N_13607,N_12350);
xnor U14833 (N_14833,N_13254,N_12626);
or U14834 (N_14834,N_13760,N_13425);
or U14835 (N_14835,N_13758,N_13313);
nor U14836 (N_14836,N_13619,N_12147);
xnor U14837 (N_14837,N_13863,N_13684);
xor U14838 (N_14838,N_12361,N_12713);
nand U14839 (N_14839,N_12572,N_12139);
nand U14840 (N_14840,N_13252,N_12068);
nand U14841 (N_14841,N_12851,N_13377);
nand U14842 (N_14842,N_13990,N_13810);
and U14843 (N_14843,N_13782,N_13170);
and U14844 (N_14844,N_13557,N_13323);
nor U14845 (N_14845,N_12522,N_13053);
and U14846 (N_14846,N_12711,N_13685);
nand U14847 (N_14847,N_12074,N_12401);
nand U14848 (N_14848,N_13355,N_12104);
xnor U14849 (N_14849,N_13225,N_13033);
xor U14850 (N_14850,N_12872,N_13032);
nand U14851 (N_14851,N_12014,N_12828);
nand U14852 (N_14852,N_13339,N_13805);
nor U14853 (N_14853,N_13202,N_12202);
nand U14854 (N_14854,N_13946,N_12597);
xor U14855 (N_14855,N_13184,N_13495);
nand U14856 (N_14856,N_13445,N_12645);
nor U14857 (N_14857,N_13911,N_12606);
xnor U14858 (N_14858,N_13741,N_12099);
nand U14859 (N_14859,N_13823,N_13013);
xnor U14860 (N_14860,N_13800,N_13128);
and U14861 (N_14861,N_13153,N_12614);
xor U14862 (N_14862,N_13395,N_12033);
nor U14863 (N_14863,N_12615,N_12425);
or U14864 (N_14864,N_13498,N_13834);
and U14865 (N_14865,N_13738,N_12283);
xnor U14866 (N_14866,N_13309,N_13232);
or U14867 (N_14867,N_12819,N_12211);
nand U14868 (N_14868,N_12185,N_13487);
xor U14869 (N_14869,N_13526,N_13944);
xnor U14870 (N_14870,N_12994,N_12973);
and U14871 (N_14871,N_13141,N_13217);
nor U14872 (N_14872,N_13913,N_13821);
nor U14873 (N_14873,N_13599,N_12124);
nand U14874 (N_14874,N_13226,N_12299);
or U14875 (N_14875,N_13019,N_12253);
xnor U14876 (N_14876,N_13001,N_13336);
nor U14877 (N_14877,N_13367,N_13590);
nor U14878 (N_14878,N_12694,N_12662);
nor U14879 (N_14879,N_13296,N_12997);
or U14880 (N_14880,N_12038,N_13728);
and U14881 (N_14881,N_12289,N_13123);
nand U14882 (N_14882,N_13133,N_13192);
nor U14883 (N_14883,N_12852,N_13919);
and U14884 (N_14884,N_13784,N_13687);
or U14885 (N_14885,N_12799,N_13094);
nand U14886 (N_14886,N_13691,N_13292);
nand U14887 (N_14887,N_13656,N_13568);
or U14888 (N_14888,N_13438,N_13505);
nand U14889 (N_14889,N_12539,N_13414);
nor U14890 (N_14890,N_12867,N_13508);
and U14891 (N_14891,N_13750,N_12940);
nor U14892 (N_14892,N_13794,N_12917);
nand U14893 (N_14893,N_12717,N_12956);
nand U14894 (N_14894,N_12429,N_13971);
nor U14895 (N_14895,N_12323,N_12951);
or U14896 (N_14896,N_12786,N_13594);
and U14897 (N_14897,N_12160,N_12407);
nand U14898 (N_14898,N_13038,N_12594);
and U14899 (N_14899,N_13867,N_13370);
xor U14900 (N_14900,N_12428,N_12203);
nor U14901 (N_14901,N_12945,N_12263);
nor U14902 (N_14902,N_12437,N_12342);
nand U14903 (N_14903,N_12659,N_12721);
nand U14904 (N_14904,N_12953,N_13671);
and U14905 (N_14905,N_12287,N_12787);
nor U14906 (N_14906,N_13644,N_13290);
nand U14907 (N_14907,N_13489,N_13253);
nand U14908 (N_14908,N_13497,N_13705);
xor U14909 (N_14909,N_13985,N_12810);
or U14910 (N_14910,N_12505,N_12587);
nand U14911 (N_14911,N_12241,N_13359);
and U14912 (N_14912,N_13779,N_12759);
xor U14913 (N_14913,N_12884,N_12728);
and U14914 (N_14914,N_12588,N_13075);
nand U14915 (N_14915,N_13608,N_13471);
xnor U14916 (N_14916,N_12473,N_13077);
xnor U14917 (N_14917,N_13411,N_13169);
nor U14918 (N_14918,N_13655,N_12347);
xnor U14919 (N_14919,N_12793,N_12966);
nor U14920 (N_14920,N_13676,N_13572);
or U14921 (N_14921,N_13993,N_12079);
nor U14922 (N_14922,N_12826,N_12849);
and U14923 (N_14923,N_12133,N_13270);
nor U14924 (N_14924,N_13751,N_13893);
nand U14925 (N_14925,N_13711,N_13177);
nor U14926 (N_14926,N_13264,N_13774);
nand U14927 (N_14927,N_12213,N_13229);
nor U14928 (N_14928,N_13090,N_12189);
and U14929 (N_14929,N_13724,N_12839);
nor U14930 (N_14930,N_13331,N_13125);
and U14931 (N_14931,N_13623,N_13236);
nand U14932 (N_14932,N_12359,N_13218);
nand U14933 (N_14933,N_12454,N_13920);
nor U14934 (N_14934,N_12637,N_12260);
and U14935 (N_14935,N_13916,N_12599);
nor U14936 (N_14936,N_12047,N_12743);
and U14937 (N_14937,N_13476,N_13279);
xor U14938 (N_14938,N_13199,N_12108);
and U14939 (N_14939,N_13260,N_12000);
nand U14940 (N_14940,N_12747,N_13307);
and U14941 (N_14941,N_12451,N_13288);
or U14942 (N_14942,N_12320,N_13076);
xor U14943 (N_14943,N_13637,N_12790);
or U14944 (N_14944,N_12233,N_12279);
nand U14945 (N_14945,N_13057,N_12009);
nor U14946 (N_14946,N_13014,N_12398);
xor U14947 (N_14947,N_12888,N_12931);
nand U14948 (N_14948,N_13923,N_12003);
and U14949 (N_14949,N_12936,N_13523);
nor U14950 (N_14950,N_12013,N_12604);
xor U14951 (N_14951,N_13521,N_12027);
nor U14952 (N_14952,N_13739,N_12870);
xor U14953 (N_14953,N_13187,N_13418);
and U14954 (N_14954,N_12174,N_12103);
nand U14955 (N_14955,N_13630,N_13680);
nand U14956 (N_14956,N_13223,N_12575);
or U14957 (N_14957,N_12266,N_12836);
and U14958 (N_14958,N_12056,N_13861);
or U14959 (N_14959,N_12157,N_12600);
nor U14960 (N_14960,N_13373,N_13293);
nor U14961 (N_14961,N_13269,N_12024);
or U14962 (N_14962,N_13468,N_12517);
nand U14963 (N_14963,N_13514,N_12228);
xor U14964 (N_14964,N_12164,N_12577);
or U14965 (N_14965,N_12062,N_12356);
nand U14966 (N_14966,N_12161,N_13726);
or U14967 (N_14967,N_12351,N_12602);
nand U14968 (N_14968,N_12258,N_12051);
nand U14969 (N_14969,N_12982,N_12020);
nor U14970 (N_14970,N_13164,N_13138);
nand U14971 (N_14971,N_13251,N_13529);
and U14972 (N_14972,N_12723,N_13371);
or U14973 (N_14973,N_12889,N_13219);
and U14974 (N_14974,N_12417,N_12249);
or U14975 (N_14975,N_12806,N_13286);
nor U14976 (N_14976,N_13405,N_13583);
nor U14977 (N_14977,N_13788,N_12535);
and U14978 (N_14978,N_12756,N_13374);
and U14979 (N_14979,N_13320,N_13957);
nand U14980 (N_14980,N_12358,N_13401);
xnor U14981 (N_14981,N_12813,N_12374);
xor U14982 (N_14982,N_12708,N_12528);
nor U14983 (N_14983,N_13261,N_13195);
and U14984 (N_14984,N_13272,N_12646);
xnor U14985 (N_14985,N_12137,N_12004);
nor U14986 (N_14986,N_12589,N_13641);
nor U14987 (N_14987,N_12848,N_13324);
and U14988 (N_14988,N_13988,N_12296);
nor U14989 (N_14989,N_13872,N_12387);
xor U14990 (N_14990,N_12030,N_12555);
nor U14991 (N_14991,N_13719,N_12182);
nand U14992 (N_14992,N_12833,N_13344);
xnor U14993 (N_14993,N_13179,N_13854);
xnor U14994 (N_14994,N_13756,N_12190);
xnor U14995 (N_14995,N_13781,N_12252);
and U14996 (N_14996,N_12900,N_12749);
and U14997 (N_14997,N_13673,N_12860);
or U14998 (N_14998,N_12076,N_12470);
nor U14999 (N_14999,N_12652,N_12114);
and U15000 (N_15000,N_13679,N_12797);
and U15001 (N_15001,N_13530,N_12519);
xor U15002 (N_15002,N_12930,N_13244);
nand U15003 (N_15003,N_13442,N_12070);
or U15004 (N_15004,N_13406,N_13534);
and U15005 (N_15005,N_12473,N_13766);
and U15006 (N_15006,N_12327,N_12586);
and U15007 (N_15007,N_12117,N_13279);
xor U15008 (N_15008,N_13811,N_13139);
nor U15009 (N_15009,N_12037,N_13088);
nor U15010 (N_15010,N_12382,N_12609);
xor U15011 (N_15011,N_13349,N_12839);
and U15012 (N_15012,N_13980,N_12589);
nor U15013 (N_15013,N_12304,N_13562);
xnor U15014 (N_15014,N_13267,N_12532);
nor U15015 (N_15015,N_13364,N_12305);
xnor U15016 (N_15016,N_13955,N_12932);
or U15017 (N_15017,N_12921,N_13697);
or U15018 (N_15018,N_13679,N_12538);
xnor U15019 (N_15019,N_13112,N_13266);
nand U15020 (N_15020,N_12266,N_13735);
or U15021 (N_15021,N_12819,N_13031);
xnor U15022 (N_15022,N_13538,N_13369);
nand U15023 (N_15023,N_13342,N_13779);
and U15024 (N_15024,N_13534,N_13189);
and U15025 (N_15025,N_13229,N_12093);
or U15026 (N_15026,N_13576,N_12320);
xnor U15027 (N_15027,N_12274,N_13069);
nand U15028 (N_15028,N_13089,N_13228);
nor U15029 (N_15029,N_13133,N_12626);
xor U15030 (N_15030,N_12874,N_13325);
xor U15031 (N_15031,N_12618,N_12328);
or U15032 (N_15032,N_12806,N_12081);
and U15033 (N_15033,N_12523,N_12549);
or U15034 (N_15034,N_12939,N_12999);
and U15035 (N_15035,N_12539,N_13420);
nand U15036 (N_15036,N_12379,N_13795);
or U15037 (N_15037,N_12448,N_13401);
and U15038 (N_15038,N_13455,N_12856);
nor U15039 (N_15039,N_12289,N_13749);
xnor U15040 (N_15040,N_13151,N_13345);
or U15041 (N_15041,N_13953,N_12734);
nor U15042 (N_15042,N_13007,N_12433);
and U15043 (N_15043,N_12754,N_13845);
nor U15044 (N_15044,N_12694,N_13815);
xor U15045 (N_15045,N_13244,N_12772);
nor U15046 (N_15046,N_13725,N_12657);
or U15047 (N_15047,N_13612,N_13653);
nand U15048 (N_15048,N_12260,N_12417);
nor U15049 (N_15049,N_13166,N_12398);
xor U15050 (N_15050,N_13228,N_13350);
or U15051 (N_15051,N_13669,N_13996);
nand U15052 (N_15052,N_13628,N_13844);
or U15053 (N_15053,N_12270,N_13553);
xor U15054 (N_15054,N_12744,N_13221);
and U15055 (N_15055,N_12297,N_12634);
nand U15056 (N_15056,N_13278,N_13770);
and U15057 (N_15057,N_12511,N_13301);
xnor U15058 (N_15058,N_12520,N_12277);
nor U15059 (N_15059,N_12785,N_13778);
nor U15060 (N_15060,N_13356,N_12139);
or U15061 (N_15061,N_13273,N_13644);
nand U15062 (N_15062,N_13609,N_13551);
xnor U15063 (N_15063,N_13031,N_13728);
nand U15064 (N_15064,N_13375,N_13523);
nor U15065 (N_15065,N_12912,N_13072);
nor U15066 (N_15066,N_12471,N_12151);
or U15067 (N_15067,N_13068,N_13289);
and U15068 (N_15068,N_13316,N_13518);
and U15069 (N_15069,N_13863,N_12459);
nand U15070 (N_15070,N_12964,N_12719);
xor U15071 (N_15071,N_12473,N_12478);
and U15072 (N_15072,N_13794,N_12827);
nand U15073 (N_15073,N_13045,N_13179);
or U15074 (N_15074,N_13618,N_12227);
nor U15075 (N_15075,N_13917,N_13046);
nand U15076 (N_15076,N_13683,N_13081);
and U15077 (N_15077,N_13946,N_12745);
and U15078 (N_15078,N_12046,N_12632);
xor U15079 (N_15079,N_13500,N_12281);
and U15080 (N_15080,N_12809,N_12206);
nor U15081 (N_15081,N_13114,N_13244);
nor U15082 (N_15082,N_13815,N_12002);
nand U15083 (N_15083,N_13506,N_12819);
or U15084 (N_15084,N_13361,N_12045);
and U15085 (N_15085,N_13836,N_12488);
nor U15086 (N_15086,N_13730,N_13941);
or U15087 (N_15087,N_13582,N_13873);
and U15088 (N_15088,N_12718,N_12747);
xnor U15089 (N_15089,N_12280,N_13041);
and U15090 (N_15090,N_12092,N_13299);
xnor U15091 (N_15091,N_13683,N_13480);
nand U15092 (N_15092,N_12357,N_12682);
xor U15093 (N_15093,N_13013,N_13133);
or U15094 (N_15094,N_13302,N_13771);
nand U15095 (N_15095,N_13088,N_12458);
and U15096 (N_15096,N_12840,N_13633);
and U15097 (N_15097,N_12879,N_12000);
or U15098 (N_15098,N_13695,N_12164);
or U15099 (N_15099,N_12458,N_12055);
xor U15100 (N_15100,N_13670,N_13804);
or U15101 (N_15101,N_13160,N_13078);
and U15102 (N_15102,N_12181,N_12564);
nor U15103 (N_15103,N_12940,N_12377);
or U15104 (N_15104,N_13101,N_12490);
nor U15105 (N_15105,N_12276,N_13284);
nor U15106 (N_15106,N_12354,N_13880);
or U15107 (N_15107,N_12886,N_13393);
xnor U15108 (N_15108,N_12538,N_13561);
xor U15109 (N_15109,N_12908,N_13251);
and U15110 (N_15110,N_13894,N_13029);
or U15111 (N_15111,N_12057,N_12503);
and U15112 (N_15112,N_12539,N_13459);
nand U15113 (N_15113,N_12769,N_13392);
or U15114 (N_15114,N_13937,N_13662);
or U15115 (N_15115,N_13815,N_13779);
nand U15116 (N_15116,N_13224,N_13491);
or U15117 (N_15117,N_12928,N_12139);
or U15118 (N_15118,N_13653,N_12176);
nor U15119 (N_15119,N_12981,N_12216);
nor U15120 (N_15120,N_13198,N_13142);
nor U15121 (N_15121,N_12792,N_13380);
or U15122 (N_15122,N_12972,N_12277);
xnor U15123 (N_15123,N_13569,N_13752);
nand U15124 (N_15124,N_12470,N_13799);
and U15125 (N_15125,N_13332,N_12668);
nand U15126 (N_15126,N_13244,N_12730);
and U15127 (N_15127,N_13248,N_12610);
nand U15128 (N_15128,N_12769,N_12000);
xor U15129 (N_15129,N_13728,N_12951);
nand U15130 (N_15130,N_13092,N_13593);
or U15131 (N_15131,N_13345,N_13098);
nand U15132 (N_15132,N_12272,N_13182);
nand U15133 (N_15133,N_13937,N_13033);
xor U15134 (N_15134,N_13464,N_13486);
and U15135 (N_15135,N_12307,N_12141);
nand U15136 (N_15136,N_12458,N_13435);
xor U15137 (N_15137,N_13901,N_13297);
and U15138 (N_15138,N_13984,N_13194);
nor U15139 (N_15139,N_12700,N_12596);
and U15140 (N_15140,N_12871,N_13134);
nor U15141 (N_15141,N_12440,N_13102);
nand U15142 (N_15142,N_12975,N_13411);
and U15143 (N_15143,N_12587,N_13876);
xnor U15144 (N_15144,N_13704,N_13369);
nor U15145 (N_15145,N_13151,N_12609);
or U15146 (N_15146,N_13068,N_13980);
nand U15147 (N_15147,N_12767,N_13223);
xor U15148 (N_15148,N_13178,N_12823);
nand U15149 (N_15149,N_13654,N_13622);
and U15150 (N_15150,N_12185,N_13181);
or U15151 (N_15151,N_12407,N_12790);
nor U15152 (N_15152,N_12903,N_13254);
nand U15153 (N_15153,N_13264,N_13188);
xor U15154 (N_15154,N_12558,N_13262);
nand U15155 (N_15155,N_13754,N_13514);
xnor U15156 (N_15156,N_13244,N_13483);
xnor U15157 (N_15157,N_12895,N_12823);
and U15158 (N_15158,N_12800,N_12296);
xor U15159 (N_15159,N_12207,N_12625);
and U15160 (N_15160,N_12662,N_13371);
and U15161 (N_15161,N_12759,N_12750);
nor U15162 (N_15162,N_13333,N_13983);
nand U15163 (N_15163,N_13997,N_12551);
nand U15164 (N_15164,N_13104,N_12767);
nand U15165 (N_15165,N_12095,N_13239);
nor U15166 (N_15166,N_13427,N_13316);
nor U15167 (N_15167,N_13258,N_13853);
and U15168 (N_15168,N_13166,N_12773);
or U15169 (N_15169,N_13275,N_12563);
and U15170 (N_15170,N_12129,N_12342);
xor U15171 (N_15171,N_12803,N_12189);
or U15172 (N_15172,N_12525,N_12348);
or U15173 (N_15173,N_12114,N_12349);
nand U15174 (N_15174,N_13802,N_13360);
xor U15175 (N_15175,N_13359,N_13054);
and U15176 (N_15176,N_13046,N_13757);
nor U15177 (N_15177,N_13456,N_12455);
and U15178 (N_15178,N_13529,N_12542);
nand U15179 (N_15179,N_13915,N_13131);
or U15180 (N_15180,N_13687,N_13522);
nor U15181 (N_15181,N_12240,N_12186);
and U15182 (N_15182,N_12766,N_13882);
or U15183 (N_15183,N_12186,N_12657);
or U15184 (N_15184,N_13621,N_13584);
or U15185 (N_15185,N_12806,N_12327);
or U15186 (N_15186,N_13174,N_13742);
and U15187 (N_15187,N_13992,N_12312);
or U15188 (N_15188,N_13812,N_12954);
and U15189 (N_15189,N_12103,N_12047);
nor U15190 (N_15190,N_13689,N_12045);
nand U15191 (N_15191,N_12299,N_13306);
and U15192 (N_15192,N_12027,N_12599);
nand U15193 (N_15193,N_13383,N_13144);
xor U15194 (N_15194,N_12379,N_13635);
nor U15195 (N_15195,N_12370,N_12687);
xnor U15196 (N_15196,N_13966,N_13804);
and U15197 (N_15197,N_12854,N_13742);
nor U15198 (N_15198,N_13723,N_12460);
nor U15199 (N_15199,N_13191,N_13631);
nor U15200 (N_15200,N_12269,N_13433);
or U15201 (N_15201,N_12271,N_13735);
nand U15202 (N_15202,N_12287,N_12385);
nand U15203 (N_15203,N_13380,N_12938);
and U15204 (N_15204,N_13169,N_12807);
xor U15205 (N_15205,N_12148,N_13134);
and U15206 (N_15206,N_12473,N_12075);
or U15207 (N_15207,N_12304,N_13817);
nand U15208 (N_15208,N_13982,N_12450);
and U15209 (N_15209,N_13093,N_13588);
or U15210 (N_15210,N_13353,N_12439);
nand U15211 (N_15211,N_13631,N_12348);
nor U15212 (N_15212,N_12260,N_12257);
nand U15213 (N_15213,N_12148,N_13982);
nor U15214 (N_15214,N_13127,N_13772);
nand U15215 (N_15215,N_12996,N_13230);
and U15216 (N_15216,N_12336,N_13374);
and U15217 (N_15217,N_12465,N_13043);
or U15218 (N_15218,N_12804,N_13842);
or U15219 (N_15219,N_13460,N_12541);
nor U15220 (N_15220,N_12447,N_12309);
nand U15221 (N_15221,N_12404,N_12591);
or U15222 (N_15222,N_12755,N_12691);
nand U15223 (N_15223,N_13354,N_12769);
and U15224 (N_15224,N_12659,N_13680);
and U15225 (N_15225,N_12722,N_13574);
and U15226 (N_15226,N_12446,N_12273);
and U15227 (N_15227,N_12935,N_12042);
nand U15228 (N_15228,N_13678,N_12697);
and U15229 (N_15229,N_12181,N_12094);
and U15230 (N_15230,N_13310,N_12522);
and U15231 (N_15231,N_13816,N_13973);
nor U15232 (N_15232,N_13254,N_12037);
nand U15233 (N_15233,N_13731,N_13742);
nand U15234 (N_15234,N_13039,N_13339);
and U15235 (N_15235,N_13454,N_13635);
nor U15236 (N_15236,N_13239,N_13994);
nand U15237 (N_15237,N_12243,N_13674);
and U15238 (N_15238,N_12132,N_13874);
nor U15239 (N_15239,N_12187,N_12372);
nand U15240 (N_15240,N_12449,N_12328);
nor U15241 (N_15241,N_12723,N_13574);
and U15242 (N_15242,N_13552,N_12328);
nor U15243 (N_15243,N_13336,N_13523);
xnor U15244 (N_15244,N_13471,N_13169);
xor U15245 (N_15245,N_12612,N_12893);
nor U15246 (N_15246,N_12807,N_13602);
nand U15247 (N_15247,N_13172,N_12476);
nor U15248 (N_15248,N_13809,N_12352);
or U15249 (N_15249,N_12191,N_12729);
and U15250 (N_15250,N_13992,N_13236);
nor U15251 (N_15251,N_12870,N_13508);
and U15252 (N_15252,N_12548,N_12243);
nor U15253 (N_15253,N_12557,N_12981);
and U15254 (N_15254,N_13503,N_12195);
nand U15255 (N_15255,N_13696,N_13175);
nor U15256 (N_15256,N_12014,N_12515);
xor U15257 (N_15257,N_13125,N_13991);
xor U15258 (N_15258,N_12332,N_13456);
xor U15259 (N_15259,N_12351,N_13647);
and U15260 (N_15260,N_12158,N_12098);
xnor U15261 (N_15261,N_13081,N_13610);
xor U15262 (N_15262,N_13353,N_12514);
nand U15263 (N_15263,N_13362,N_12604);
xnor U15264 (N_15264,N_13175,N_13292);
xnor U15265 (N_15265,N_13014,N_13725);
and U15266 (N_15266,N_12046,N_13502);
nand U15267 (N_15267,N_12840,N_12642);
nand U15268 (N_15268,N_13144,N_13832);
or U15269 (N_15269,N_12856,N_12453);
nand U15270 (N_15270,N_13248,N_12784);
nor U15271 (N_15271,N_13256,N_12591);
or U15272 (N_15272,N_12414,N_12003);
or U15273 (N_15273,N_12983,N_13410);
nor U15274 (N_15274,N_12149,N_12303);
nand U15275 (N_15275,N_12544,N_13780);
xor U15276 (N_15276,N_13429,N_12033);
nand U15277 (N_15277,N_13554,N_13169);
xor U15278 (N_15278,N_13881,N_12888);
or U15279 (N_15279,N_13027,N_12391);
nor U15280 (N_15280,N_13899,N_12550);
nor U15281 (N_15281,N_13573,N_12691);
nor U15282 (N_15282,N_12367,N_13166);
nor U15283 (N_15283,N_13474,N_12653);
nor U15284 (N_15284,N_12200,N_13630);
and U15285 (N_15285,N_13102,N_13255);
nor U15286 (N_15286,N_13685,N_12522);
nand U15287 (N_15287,N_13256,N_12580);
or U15288 (N_15288,N_12535,N_13465);
nor U15289 (N_15289,N_12488,N_13147);
nand U15290 (N_15290,N_12329,N_12755);
nand U15291 (N_15291,N_12107,N_12284);
or U15292 (N_15292,N_13280,N_13901);
nor U15293 (N_15293,N_12086,N_13547);
nand U15294 (N_15294,N_12575,N_13134);
or U15295 (N_15295,N_13276,N_13642);
nor U15296 (N_15296,N_13928,N_12552);
nand U15297 (N_15297,N_12959,N_13504);
xnor U15298 (N_15298,N_12076,N_12621);
or U15299 (N_15299,N_12996,N_13175);
xnor U15300 (N_15300,N_12001,N_13894);
nand U15301 (N_15301,N_12139,N_12628);
or U15302 (N_15302,N_12979,N_12558);
nand U15303 (N_15303,N_13519,N_12743);
xor U15304 (N_15304,N_12286,N_13457);
or U15305 (N_15305,N_12402,N_13224);
and U15306 (N_15306,N_13931,N_13870);
nand U15307 (N_15307,N_12671,N_12947);
and U15308 (N_15308,N_13047,N_13091);
xnor U15309 (N_15309,N_13507,N_12045);
nor U15310 (N_15310,N_12079,N_13067);
nand U15311 (N_15311,N_13034,N_13710);
nor U15312 (N_15312,N_13936,N_13133);
nand U15313 (N_15313,N_13365,N_13416);
and U15314 (N_15314,N_13780,N_13125);
nor U15315 (N_15315,N_12277,N_12463);
or U15316 (N_15316,N_12460,N_13499);
nor U15317 (N_15317,N_12104,N_12492);
or U15318 (N_15318,N_13051,N_13812);
or U15319 (N_15319,N_13483,N_13054);
or U15320 (N_15320,N_12959,N_12903);
or U15321 (N_15321,N_12574,N_13047);
nand U15322 (N_15322,N_13022,N_12965);
xnor U15323 (N_15323,N_13866,N_12192);
xor U15324 (N_15324,N_12481,N_13832);
and U15325 (N_15325,N_13315,N_13131);
nor U15326 (N_15326,N_12051,N_13250);
nand U15327 (N_15327,N_12031,N_12034);
xnor U15328 (N_15328,N_13680,N_13407);
nor U15329 (N_15329,N_12137,N_12406);
and U15330 (N_15330,N_12555,N_12484);
xnor U15331 (N_15331,N_13584,N_12887);
nor U15332 (N_15332,N_13293,N_13191);
nor U15333 (N_15333,N_13118,N_13663);
or U15334 (N_15334,N_13723,N_13774);
nor U15335 (N_15335,N_12102,N_13381);
xor U15336 (N_15336,N_13245,N_12556);
and U15337 (N_15337,N_13767,N_12870);
or U15338 (N_15338,N_12284,N_12677);
and U15339 (N_15339,N_12052,N_13750);
xor U15340 (N_15340,N_13519,N_12642);
or U15341 (N_15341,N_12483,N_13059);
xnor U15342 (N_15342,N_13960,N_13828);
xnor U15343 (N_15343,N_13705,N_13319);
or U15344 (N_15344,N_12275,N_13410);
and U15345 (N_15345,N_13827,N_13453);
nand U15346 (N_15346,N_12589,N_12293);
and U15347 (N_15347,N_12870,N_13786);
and U15348 (N_15348,N_12459,N_13132);
nand U15349 (N_15349,N_12091,N_13001);
or U15350 (N_15350,N_13589,N_12026);
or U15351 (N_15351,N_12401,N_13688);
nor U15352 (N_15352,N_12352,N_12837);
or U15353 (N_15353,N_13441,N_12288);
nand U15354 (N_15354,N_13482,N_13968);
xnor U15355 (N_15355,N_13922,N_13690);
nor U15356 (N_15356,N_13689,N_13697);
xnor U15357 (N_15357,N_12691,N_12978);
nor U15358 (N_15358,N_12529,N_12246);
nand U15359 (N_15359,N_12514,N_12472);
xnor U15360 (N_15360,N_13027,N_13330);
or U15361 (N_15361,N_13261,N_13133);
and U15362 (N_15362,N_13377,N_12877);
nand U15363 (N_15363,N_13256,N_12705);
and U15364 (N_15364,N_13225,N_13860);
or U15365 (N_15365,N_12877,N_13551);
xor U15366 (N_15366,N_13709,N_12464);
or U15367 (N_15367,N_13387,N_13344);
or U15368 (N_15368,N_12992,N_12155);
nor U15369 (N_15369,N_12253,N_12357);
xnor U15370 (N_15370,N_13764,N_13063);
nand U15371 (N_15371,N_13709,N_13417);
nor U15372 (N_15372,N_13876,N_12311);
and U15373 (N_15373,N_13077,N_12162);
nor U15374 (N_15374,N_13884,N_12230);
nor U15375 (N_15375,N_12359,N_13572);
and U15376 (N_15376,N_12787,N_13446);
xnor U15377 (N_15377,N_13544,N_13869);
or U15378 (N_15378,N_12911,N_12645);
nand U15379 (N_15379,N_13857,N_13409);
nand U15380 (N_15380,N_12551,N_13079);
nand U15381 (N_15381,N_12506,N_12573);
or U15382 (N_15382,N_12291,N_13584);
nand U15383 (N_15383,N_12883,N_13019);
or U15384 (N_15384,N_13909,N_12614);
and U15385 (N_15385,N_13152,N_13873);
nor U15386 (N_15386,N_12420,N_12481);
xor U15387 (N_15387,N_12927,N_13701);
or U15388 (N_15388,N_13877,N_12502);
and U15389 (N_15389,N_12579,N_13677);
nand U15390 (N_15390,N_12035,N_13178);
or U15391 (N_15391,N_12702,N_12670);
nor U15392 (N_15392,N_13988,N_12188);
or U15393 (N_15393,N_13625,N_13563);
xnor U15394 (N_15394,N_12563,N_12921);
nor U15395 (N_15395,N_13073,N_12725);
xnor U15396 (N_15396,N_13128,N_12994);
and U15397 (N_15397,N_13340,N_13324);
and U15398 (N_15398,N_13597,N_13585);
nor U15399 (N_15399,N_13154,N_13126);
nor U15400 (N_15400,N_13076,N_12579);
nand U15401 (N_15401,N_12235,N_12332);
nand U15402 (N_15402,N_13167,N_12575);
or U15403 (N_15403,N_13273,N_12194);
and U15404 (N_15404,N_12639,N_12494);
nand U15405 (N_15405,N_13085,N_13552);
and U15406 (N_15406,N_12599,N_13922);
nor U15407 (N_15407,N_13121,N_13124);
or U15408 (N_15408,N_13720,N_13040);
or U15409 (N_15409,N_12195,N_12309);
xor U15410 (N_15410,N_12746,N_13216);
nand U15411 (N_15411,N_12947,N_12982);
nor U15412 (N_15412,N_12602,N_13834);
or U15413 (N_15413,N_13049,N_13519);
and U15414 (N_15414,N_12863,N_13182);
or U15415 (N_15415,N_12391,N_12803);
nand U15416 (N_15416,N_13744,N_13033);
nor U15417 (N_15417,N_12555,N_13930);
xnor U15418 (N_15418,N_13202,N_12592);
nor U15419 (N_15419,N_12420,N_12395);
xor U15420 (N_15420,N_13801,N_13263);
and U15421 (N_15421,N_13260,N_12292);
and U15422 (N_15422,N_13427,N_12813);
nor U15423 (N_15423,N_12218,N_13367);
and U15424 (N_15424,N_13582,N_13865);
xnor U15425 (N_15425,N_12708,N_12033);
nor U15426 (N_15426,N_13029,N_12672);
or U15427 (N_15427,N_13217,N_13013);
nor U15428 (N_15428,N_13987,N_12177);
or U15429 (N_15429,N_12732,N_13843);
nor U15430 (N_15430,N_12064,N_13316);
and U15431 (N_15431,N_12018,N_13650);
nor U15432 (N_15432,N_13020,N_13681);
or U15433 (N_15433,N_12546,N_12040);
and U15434 (N_15434,N_13986,N_12868);
nand U15435 (N_15435,N_13693,N_12150);
nor U15436 (N_15436,N_12109,N_13008);
xnor U15437 (N_15437,N_13740,N_12597);
and U15438 (N_15438,N_13380,N_12837);
nand U15439 (N_15439,N_12615,N_12252);
nand U15440 (N_15440,N_12955,N_13366);
and U15441 (N_15441,N_12539,N_13789);
nand U15442 (N_15442,N_12375,N_13908);
nor U15443 (N_15443,N_12996,N_12057);
and U15444 (N_15444,N_12010,N_12392);
or U15445 (N_15445,N_13283,N_13873);
nor U15446 (N_15446,N_13620,N_13538);
or U15447 (N_15447,N_12622,N_12952);
nand U15448 (N_15448,N_12753,N_12756);
nand U15449 (N_15449,N_13341,N_12863);
nand U15450 (N_15450,N_12759,N_12870);
nand U15451 (N_15451,N_12017,N_13559);
nand U15452 (N_15452,N_12883,N_12092);
or U15453 (N_15453,N_13464,N_13592);
nand U15454 (N_15454,N_12233,N_12120);
or U15455 (N_15455,N_12478,N_13723);
xor U15456 (N_15456,N_13744,N_13621);
xnor U15457 (N_15457,N_13321,N_12303);
nor U15458 (N_15458,N_12130,N_13743);
or U15459 (N_15459,N_13839,N_13650);
nand U15460 (N_15460,N_12479,N_12830);
nand U15461 (N_15461,N_12565,N_12518);
nor U15462 (N_15462,N_12067,N_12330);
and U15463 (N_15463,N_12601,N_12232);
and U15464 (N_15464,N_12270,N_13947);
nand U15465 (N_15465,N_13282,N_12983);
nor U15466 (N_15466,N_13148,N_12279);
or U15467 (N_15467,N_12086,N_13609);
nand U15468 (N_15468,N_12261,N_13103);
nand U15469 (N_15469,N_12476,N_12555);
or U15470 (N_15470,N_12266,N_12642);
or U15471 (N_15471,N_13293,N_12023);
nand U15472 (N_15472,N_13491,N_13843);
and U15473 (N_15473,N_13053,N_12666);
or U15474 (N_15474,N_12702,N_12682);
nand U15475 (N_15475,N_12173,N_13914);
or U15476 (N_15476,N_13668,N_13058);
or U15477 (N_15477,N_12580,N_12498);
xor U15478 (N_15478,N_12209,N_13247);
nor U15479 (N_15479,N_13056,N_13806);
and U15480 (N_15480,N_13508,N_12392);
nor U15481 (N_15481,N_13086,N_13677);
xor U15482 (N_15482,N_13264,N_13006);
and U15483 (N_15483,N_13716,N_13388);
and U15484 (N_15484,N_13564,N_12221);
nand U15485 (N_15485,N_12116,N_12816);
nand U15486 (N_15486,N_12929,N_13019);
and U15487 (N_15487,N_13340,N_13088);
nor U15488 (N_15488,N_13491,N_12160);
or U15489 (N_15489,N_12824,N_12993);
nor U15490 (N_15490,N_13646,N_12888);
and U15491 (N_15491,N_12951,N_13819);
or U15492 (N_15492,N_13140,N_12887);
or U15493 (N_15493,N_13035,N_12006);
nor U15494 (N_15494,N_13907,N_13040);
and U15495 (N_15495,N_12722,N_12103);
or U15496 (N_15496,N_13837,N_13312);
xnor U15497 (N_15497,N_13251,N_12429);
and U15498 (N_15498,N_13887,N_12566);
and U15499 (N_15499,N_13742,N_12005);
or U15500 (N_15500,N_13998,N_13198);
nor U15501 (N_15501,N_13921,N_13903);
xnor U15502 (N_15502,N_12878,N_12781);
nand U15503 (N_15503,N_12420,N_12323);
and U15504 (N_15504,N_13789,N_12518);
or U15505 (N_15505,N_13111,N_12795);
or U15506 (N_15506,N_13511,N_13547);
nand U15507 (N_15507,N_12821,N_12598);
and U15508 (N_15508,N_13741,N_13227);
nand U15509 (N_15509,N_13459,N_12924);
nor U15510 (N_15510,N_12217,N_13898);
and U15511 (N_15511,N_12812,N_13456);
xor U15512 (N_15512,N_13695,N_13639);
nand U15513 (N_15513,N_12983,N_13948);
nand U15514 (N_15514,N_12917,N_12784);
xnor U15515 (N_15515,N_13000,N_12017);
xor U15516 (N_15516,N_12473,N_12693);
and U15517 (N_15517,N_12970,N_13804);
xor U15518 (N_15518,N_13231,N_13724);
nand U15519 (N_15519,N_12187,N_12255);
nand U15520 (N_15520,N_12710,N_12066);
or U15521 (N_15521,N_13893,N_13212);
nand U15522 (N_15522,N_12147,N_12337);
or U15523 (N_15523,N_13355,N_12070);
xnor U15524 (N_15524,N_12835,N_13044);
xor U15525 (N_15525,N_13648,N_12244);
xnor U15526 (N_15526,N_13252,N_12036);
nor U15527 (N_15527,N_13214,N_13320);
nor U15528 (N_15528,N_13076,N_13046);
or U15529 (N_15529,N_12307,N_13996);
and U15530 (N_15530,N_13578,N_12008);
xor U15531 (N_15531,N_13886,N_12141);
and U15532 (N_15532,N_12843,N_12467);
or U15533 (N_15533,N_13369,N_13478);
xnor U15534 (N_15534,N_13286,N_13382);
or U15535 (N_15535,N_12626,N_12981);
xnor U15536 (N_15536,N_13409,N_13798);
and U15537 (N_15537,N_12689,N_12632);
and U15538 (N_15538,N_12216,N_13349);
and U15539 (N_15539,N_12651,N_12655);
and U15540 (N_15540,N_13335,N_13097);
and U15541 (N_15541,N_13207,N_13155);
xor U15542 (N_15542,N_13578,N_13907);
xor U15543 (N_15543,N_12922,N_12178);
and U15544 (N_15544,N_12144,N_12820);
or U15545 (N_15545,N_13982,N_12085);
nor U15546 (N_15546,N_13700,N_13835);
nand U15547 (N_15547,N_13823,N_12517);
or U15548 (N_15548,N_12758,N_12840);
and U15549 (N_15549,N_12519,N_12437);
xor U15550 (N_15550,N_12725,N_12987);
xnor U15551 (N_15551,N_13802,N_12729);
nor U15552 (N_15552,N_13807,N_12616);
or U15553 (N_15553,N_13839,N_13299);
and U15554 (N_15554,N_13903,N_13623);
xnor U15555 (N_15555,N_13124,N_13826);
and U15556 (N_15556,N_12883,N_12467);
or U15557 (N_15557,N_12407,N_13559);
nor U15558 (N_15558,N_12762,N_13318);
or U15559 (N_15559,N_12680,N_13397);
xnor U15560 (N_15560,N_13876,N_12594);
and U15561 (N_15561,N_13564,N_13395);
or U15562 (N_15562,N_13148,N_12450);
or U15563 (N_15563,N_13496,N_12924);
nor U15564 (N_15564,N_13586,N_12888);
nor U15565 (N_15565,N_13267,N_13450);
or U15566 (N_15566,N_12197,N_13101);
nand U15567 (N_15567,N_13578,N_13509);
or U15568 (N_15568,N_13115,N_12399);
or U15569 (N_15569,N_12578,N_13598);
nand U15570 (N_15570,N_12682,N_13512);
xor U15571 (N_15571,N_12586,N_12556);
nand U15572 (N_15572,N_12983,N_12804);
xnor U15573 (N_15573,N_13375,N_12921);
nand U15574 (N_15574,N_13178,N_12309);
nand U15575 (N_15575,N_12498,N_12988);
xor U15576 (N_15576,N_13278,N_12561);
nor U15577 (N_15577,N_13614,N_12781);
nor U15578 (N_15578,N_12583,N_12202);
and U15579 (N_15579,N_12803,N_13741);
or U15580 (N_15580,N_12330,N_12104);
nand U15581 (N_15581,N_12963,N_12283);
nor U15582 (N_15582,N_13534,N_13658);
or U15583 (N_15583,N_12323,N_13881);
and U15584 (N_15584,N_12775,N_13529);
and U15585 (N_15585,N_12304,N_13329);
nor U15586 (N_15586,N_12837,N_13794);
or U15587 (N_15587,N_13214,N_13671);
nand U15588 (N_15588,N_12017,N_12402);
xnor U15589 (N_15589,N_12160,N_13057);
or U15590 (N_15590,N_13552,N_12319);
and U15591 (N_15591,N_13812,N_12465);
nand U15592 (N_15592,N_13248,N_13288);
and U15593 (N_15593,N_13321,N_13641);
nand U15594 (N_15594,N_13526,N_13709);
nor U15595 (N_15595,N_13642,N_13522);
xnor U15596 (N_15596,N_12034,N_13197);
and U15597 (N_15597,N_12564,N_12593);
nor U15598 (N_15598,N_12431,N_13574);
or U15599 (N_15599,N_13214,N_13241);
xnor U15600 (N_15600,N_12671,N_13634);
or U15601 (N_15601,N_12916,N_12321);
xnor U15602 (N_15602,N_13961,N_12379);
and U15603 (N_15603,N_13218,N_12127);
and U15604 (N_15604,N_12416,N_12935);
xor U15605 (N_15605,N_12740,N_12491);
or U15606 (N_15606,N_13717,N_13738);
nor U15607 (N_15607,N_12273,N_13762);
nand U15608 (N_15608,N_12255,N_13909);
nor U15609 (N_15609,N_12058,N_12129);
xor U15610 (N_15610,N_13810,N_12199);
xor U15611 (N_15611,N_13451,N_12514);
xor U15612 (N_15612,N_13934,N_12084);
nor U15613 (N_15613,N_13988,N_12433);
and U15614 (N_15614,N_13197,N_13621);
or U15615 (N_15615,N_12719,N_12134);
nor U15616 (N_15616,N_12195,N_13472);
and U15617 (N_15617,N_12172,N_12464);
nor U15618 (N_15618,N_13606,N_12046);
and U15619 (N_15619,N_13719,N_12665);
and U15620 (N_15620,N_12771,N_13664);
or U15621 (N_15621,N_13967,N_13411);
or U15622 (N_15622,N_12850,N_13414);
nor U15623 (N_15623,N_13976,N_13656);
nor U15624 (N_15624,N_13633,N_13615);
nor U15625 (N_15625,N_12174,N_13445);
and U15626 (N_15626,N_12224,N_12778);
nor U15627 (N_15627,N_13144,N_13061);
nand U15628 (N_15628,N_13096,N_13839);
nor U15629 (N_15629,N_12276,N_12036);
nor U15630 (N_15630,N_12585,N_12229);
and U15631 (N_15631,N_12330,N_12232);
nor U15632 (N_15632,N_13802,N_13746);
or U15633 (N_15633,N_12358,N_13460);
and U15634 (N_15634,N_13417,N_12933);
nor U15635 (N_15635,N_12418,N_13146);
nand U15636 (N_15636,N_13057,N_13620);
or U15637 (N_15637,N_13870,N_13999);
nand U15638 (N_15638,N_12685,N_13085);
nand U15639 (N_15639,N_13151,N_12824);
nand U15640 (N_15640,N_13279,N_13728);
nor U15641 (N_15641,N_12444,N_13193);
xor U15642 (N_15642,N_12503,N_12400);
or U15643 (N_15643,N_13954,N_13887);
nand U15644 (N_15644,N_12259,N_13559);
xor U15645 (N_15645,N_13332,N_12104);
and U15646 (N_15646,N_13945,N_12051);
xor U15647 (N_15647,N_12713,N_12379);
nand U15648 (N_15648,N_12493,N_13989);
nand U15649 (N_15649,N_13858,N_12599);
xor U15650 (N_15650,N_13254,N_13285);
nand U15651 (N_15651,N_13192,N_13070);
and U15652 (N_15652,N_12155,N_12379);
xnor U15653 (N_15653,N_12621,N_13581);
nor U15654 (N_15654,N_13495,N_12899);
xnor U15655 (N_15655,N_12392,N_12296);
nand U15656 (N_15656,N_13248,N_13371);
nand U15657 (N_15657,N_13662,N_13657);
or U15658 (N_15658,N_12720,N_12300);
nor U15659 (N_15659,N_13387,N_13107);
xnor U15660 (N_15660,N_12402,N_12209);
xnor U15661 (N_15661,N_13044,N_12339);
or U15662 (N_15662,N_13510,N_13049);
and U15663 (N_15663,N_12690,N_12543);
nand U15664 (N_15664,N_13310,N_13280);
xnor U15665 (N_15665,N_12121,N_12985);
nand U15666 (N_15666,N_12078,N_12602);
nor U15667 (N_15667,N_12681,N_13707);
nor U15668 (N_15668,N_13242,N_13196);
or U15669 (N_15669,N_13075,N_13117);
and U15670 (N_15670,N_13486,N_12603);
nor U15671 (N_15671,N_12037,N_13371);
and U15672 (N_15672,N_13882,N_13330);
nand U15673 (N_15673,N_12788,N_12214);
nand U15674 (N_15674,N_13009,N_13765);
nand U15675 (N_15675,N_12165,N_12275);
and U15676 (N_15676,N_12560,N_12069);
nand U15677 (N_15677,N_12265,N_12186);
or U15678 (N_15678,N_13588,N_13552);
and U15679 (N_15679,N_12711,N_13178);
xnor U15680 (N_15680,N_13220,N_12791);
or U15681 (N_15681,N_13551,N_12832);
nand U15682 (N_15682,N_12031,N_12953);
xnor U15683 (N_15683,N_13634,N_12273);
nor U15684 (N_15684,N_13976,N_13947);
and U15685 (N_15685,N_12813,N_12741);
and U15686 (N_15686,N_12020,N_12281);
nor U15687 (N_15687,N_13282,N_12671);
and U15688 (N_15688,N_13954,N_13763);
and U15689 (N_15689,N_12026,N_13359);
xnor U15690 (N_15690,N_12964,N_13906);
or U15691 (N_15691,N_12635,N_12020);
or U15692 (N_15692,N_12644,N_12280);
nor U15693 (N_15693,N_13338,N_13296);
nor U15694 (N_15694,N_13549,N_12148);
and U15695 (N_15695,N_12326,N_13263);
xnor U15696 (N_15696,N_12413,N_13056);
or U15697 (N_15697,N_13274,N_12031);
nor U15698 (N_15698,N_13675,N_13862);
and U15699 (N_15699,N_12520,N_12061);
xor U15700 (N_15700,N_13775,N_13593);
xor U15701 (N_15701,N_12289,N_12055);
nand U15702 (N_15702,N_13440,N_12917);
and U15703 (N_15703,N_13980,N_12764);
nand U15704 (N_15704,N_12217,N_12583);
nor U15705 (N_15705,N_13707,N_13314);
nor U15706 (N_15706,N_13555,N_13019);
and U15707 (N_15707,N_12387,N_13045);
xnor U15708 (N_15708,N_12767,N_12427);
nor U15709 (N_15709,N_13425,N_12516);
xor U15710 (N_15710,N_13511,N_12017);
and U15711 (N_15711,N_13065,N_13129);
xnor U15712 (N_15712,N_12605,N_12850);
or U15713 (N_15713,N_13169,N_13458);
xnor U15714 (N_15714,N_13202,N_12268);
nor U15715 (N_15715,N_12751,N_13290);
nor U15716 (N_15716,N_12819,N_13729);
and U15717 (N_15717,N_13661,N_13360);
and U15718 (N_15718,N_12598,N_13316);
and U15719 (N_15719,N_13367,N_12139);
nor U15720 (N_15720,N_12743,N_12008);
and U15721 (N_15721,N_13165,N_13060);
or U15722 (N_15722,N_13468,N_13562);
xor U15723 (N_15723,N_13127,N_13001);
nor U15724 (N_15724,N_12877,N_12829);
and U15725 (N_15725,N_12830,N_12822);
or U15726 (N_15726,N_13663,N_12913);
or U15727 (N_15727,N_12421,N_12262);
and U15728 (N_15728,N_13914,N_12212);
nor U15729 (N_15729,N_13152,N_12018);
and U15730 (N_15730,N_12469,N_13218);
xnor U15731 (N_15731,N_13509,N_12548);
or U15732 (N_15732,N_12851,N_13822);
or U15733 (N_15733,N_12343,N_13562);
or U15734 (N_15734,N_13321,N_13991);
nor U15735 (N_15735,N_12747,N_13946);
and U15736 (N_15736,N_12035,N_13896);
and U15737 (N_15737,N_13402,N_12069);
nand U15738 (N_15738,N_13324,N_13558);
or U15739 (N_15739,N_12411,N_12680);
nand U15740 (N_15740,N_12883,N_12921);
xor U15741 (N_15741,N_12155,N_12169);
xor U15742 (N_15742,N_12574,N_13561);
or U15743 (N_15743,N_13057,N_12168);
nor U15744 (N_15744,N_13682,N_13925);
xor U15745 (N_15745,N_13789,N_12624);
nor U15746 (N_15746,N_13499,N_12154);
and U15747 (N_15747,N_12768,N_12604);
and U15748 (N_15748,N_12981,N_12463);
nand U15749 (N_15749,N_13503,N_12849);
or U15750 (N_15750,N_13884,N_13549);
or U15751 (N_15751,N_12939,N_13948);
or U15752 (N_15752,N_13604,N_13522);
and U15753 (N_15753,N_12473,N_13083);
and U15754 (N_15754,N_13701,N_13026);
nor U15755 (N_15755,N_12313,N_13611);
or U15756 (N_15756,N_12534,N_13422);
and U15757 (N_15757,N_13086,N_13403);
and U15758 (N_15758,N_13086,N_12407);
xnor U15759 (N_15759,N_13037,N_12117);
xor U15760 (N_15760,N_12426,N_12821);
xnor U15761 (N_15761,N_12351,N_12247);
nor U15762 (N_15762,N_12195,N_12198);
nand U15763 (N_15763,N_13984,N_13325);
and U15764 (N_15764,N_13923,N_12317);
nand U15765 (N_15765,N_12871,N_12209);
nor U15766 (N_15766,N_13995,N_12034);
xnor U15767 (N_15767,N_13239,N_13417);
nand U15768 (N_15768,N_13455,N_12020);
xnor U15769 (N_15769,N_12915,N_12651);
nand U15770 (N_15770,N_12444,N_12483);
or U15771 (N_15771,N_12771,N_13399);
and U15772 (N_15772,N_13297,N_13542);
xnor U15773 (N_15773,N_12295,N_12156);
nand U15774 (N_15774,N_13419,N_12968);
or U15775 (N_15775,N_12918,N_13977);
and U15776 (N_15776,N_13820,N_13052);
and U15777 (N_15777,N_13017,N_13400);
xnor U15778 (N_15778,N_13788,N_12243);
xnor U15779 (N_15779,N_12681,N_12219);
and U15780 (N_15780,N_12260,N_13539);
and U15781 (N_15781,N_12782,N_13740);
xnor U15782 (N_15782,N_13188,N_12134);
nand U15783 (N_15783,N_13250,N_13875);
nor U15784 (N_15784,N_12076,N_13738);
nor U15785 (N_15785,N_12082,N_13705);
xor U15786 (N_15786,N_13173,N_13412);
nor U15787 (N_15787,N_13129,N_13604);
xnor U15788 (N_15788,N_13066,N_12515);
or U15789 (N_15789,N_12361,N_12973);
or U15790 (N_15790,N_13679,N_13390);
and U15791 (N_15791,N_12189,N_13343);
and U15792 (N_15792,N_12498,N_13701);
xor U15793 (N_15793,N_12741,N_13988);
xor U15794 (N_15794,N_13010,N_12216);
and U15795 (N_15795,N_12057,N_12922);
or U15796 (N_15796,N_12100,N_12519);
and U15797 (N_15797,N_13262,N_13127);
and U15798 (N_15798,N_12305,N_12189);
or U15799 (N_15799,N_12866,N_13003);
nor U15800 (N_15800,N_12194,N_13216);
or U15801 (N_15801,N_13142,N_12004);
xnor U15802 (N_15802,N_13768,N_13557);
or U15803 (N_15803,N_13148,N_13464);
nor U15804 (N_15804,N_13861,N_13079);
or U15805 (N_15805,N_13326,N_13208);
or U15806 (N_15806,N_13091,N_12330);
nand U15807 (N_15807,N_12742,N_13413);
or U15808 (N_15808,N_12997,N_12463);
nand U15809 (N_15809,N_13380,N_12303);
or U15810 (N_15810,N_13798,N_13712);
nor U15811 (N_15811,N_12764,N_12761);
or U15812 (N_15812,N_12814,N_13660);
nor U15813 (N_15813,N_13361,N_13042);
and U15814 (N_15814,N_13219,N_13332);
and U15815 (N_15815,N_12440,N_13465);
xor U15816 (N_15816,N_13939,N_12434);
and U15817 (N_15817,N_12598,N_13062);
xnor U15818 (N_15818,N_12793,N_12061);
xnor U15819 (N_15819,N_12799,N_13528);
or U15820 (N_15820,N_13633,N_13354);
xnor U15821 (N_15821,N_12552,N_13542);
nor U15822 (N_15822,N_13406,N_13543);
xnor U15823 (N_15823,N_13485,N_12466);
and U15824 (N_15824,N_12150,N_13073);
and U15825 (N_15825,N_12568,N_12781);
xor U15826 (N_15826,N_13096,N_13092);
and U15827 (N_15827,N_13840,N_13048);
and U15828 (N_15828,N_12859,N_13625);
nand U15829 (N_15829,N_12558,N_13311);
nor U15830 (N_15830,N_13310,N_12574);
xnor U15831 (N_15831,N_13146,N_12736);
nand U15832 (N_15832,N_12558,N_12291);
and U15833 (N_15833,N_12931,N_13998);
or U15834 (N_15834,N_13910,N_13308);
xnor U15835 (N_15835,N_13820,N_12931);
xor U15836 (N_15836,N_12252,N_13903);
nor U15837 (N_15837,N_12190,N_12228);
and U15838 (N_15838,N_13677,N_13959);
and U15839 (N_15839,N_12890,N_13216);
nand U15840 (N_15840,N_12908,N_13262);
nor U15841 (N_15841,N_12076,N_13833);
xor U15842 (N_15842,N_12656,N_12555);
xnor U15843 (N_15843,N_13953,N_13973);
nand U15844 (N_15844,N_13255,N_13758);
and U15845 (N_15845,N_13638,N_12289);
nand U15846 (N_15846,N_12284,N_12315);
nor U15847 (N_15847,N_12957,N_12246);
nor U15848 (N_15848,N_13302,N_13142);
and U15849 (N_15849,N_12627,N_13006);
xor U15850 (N_15850,N_12077,N_13142);
and U15851 (N_15851,N_13615,N_12061);
xor U15852 (N_15852,N_12744,N_12565);
or U15853 (N_15853,N_13846,N_12302);
xnor U15854 (N_15854,N_12597,N_13426);
or U15855 (N_15855,N_12923,N_12636);
nand U15856 (N_15856,N_12657,N_12905);
and U15857 (N_15857,N_13182,N_13507);
nand U15858 (N_15858,N_12798,N_12082);
and U15859 (N_15859,N_12195,N_12437);
nand U15860 (N_15860,N_13431,N_13839);
nor U15861 (N_15861,N_13797,N_13652);
nor U15862 (N_15862,N_13124,N_13713);
xnor U15863 (N_15863,N_12791,N_12524);
or U15864 (N_15864,N_13942,N_13187);
xor U15865 (N_15865,N_13191,N_12583);
nor U15866 (N_15866,N_13238,N_12913);
nand U15867 (N_15867,N_13324,N_13796);
nor U15868 (N_15868,N_13184,N_13783);
nor U15869 (N_15869,N_13892,N_13116);
nor U15870 (N_15870,N_13830,N_13210);
or U15871 (N_15871,N_12106,N_12400);
nor U15872 (N_15872,N_13243,N_12259);
xnor U15873 (N_15873,N_13426,N_13806);
nor U15874 (N_15874,N_12493,N_12979);
xnor U15875 (N_15875,N_13233,N_13147);
or U15876 (N_15876,N_13279,N_13953);
and U15877 (N_15877,N_13232,N_13354);
nor U15878 (N_15878,N_12981,N_12488);
xnor U15879 (N_15879,N_12552,N_12085);
xor U15880 (N_15880,N_12298,N_12980);
nand U15881 (N_15881,N_12116,N_13131);
and U15882 (N_15882,N_13153,N_12163);
nand U15883 (N_15883,N_12328,N_13374);
nand U15884 (N_15884,N_13516,N_13082);
or U15885 (N_15885,N_13798,N_12050);
or U15886 (N_15886,N_12485,N_12376);
and U15887 (N_15887,N_12137,N_12352);
nor U15888 (N_15888,N_12837,N_13596);
nor U15889 (N_15889,N_13705,N_13059);
or U15890 (N_15890,N_12448,N_13532);
nor U15891 (N_15891,N_12176,N_13176);
nand U15892 (N_15892,N_13208,N_13495);
or U15893 (N_15893,N_12514,N_13285);
xnor U15894 (N_15894,N_13488,N_12606);
xnor U15895 (N_15895,N_12141,N_12234);
nor U15896 (N_15896,N_13324,N_12819);
nand U15897 (N_15897,N_13077,N_13196);
nor U15898 (N_15898,N_12254,N_12700);
xor U15899 (N_15899,N_12785,N_12288);
and U15900 (N_15900,N_13035,N_13361);
nor U15901 (N_15901,N_13081,N_12114);
nor U15902 (N_15902,N_12895,N_12730);
xnor U15903 (N_15903,N_12900,N_13665);
nor U15904 (N_15904,N_12451,N_12166);
and U15905 (N_15905,N_12441,N_12069);
xnor U15906 (N_15906,N_13488,N_13434);
nand U15907 (N_15907,N_12809,N_12707);
xnor U15908 (N_15908,N_12055,N_13207);
nor U15909 (N_15909,N_13049,N_13320);
nor U15910 (N_15910,N_12565,N_13410);
and U15911 (N_15911,N_13701,N_12228);
nor U15912 (N_15912,N_13003,N_12606);
xor U15913 (N_15913,N_12786,N_13076);
or U15914 (N_15914,N_13297,N_13675);
nand U15915 (N_15915,N_12217,N_12531);
nand U15916 (N_15916,N_12530,N_13414);
and U15917 (N_15917,N_12035,N_12029);
nor U15918 (N_15918,N_12997,N_12990);
and U15919 (N_15919,N_13855,N_13814);
or U15920 (N_15920,N_13361,N_12162);
nor U15921 (N_15921,N_13727,N_13149);
nand U15922 (N_15922,N_13633,N_12088);
or U15923 (N_15923,N_13072,N_13925);
and U15924 (N_15924,N_13187,N_12462);
or U15925 (N_15925,N_12794,N_12499);
or U15926 (N_15926,N_12220,N_13889);
nor U15927 (N_15927,N_13315,N_13388);
nand U15928 (N_15928,N_13528,N_12425);
or U15929 (N_15929,N_13429,N_13378);
nand U15930 (N_15930,N_13176,N_13730);
nor U15931 (N_15931,N_12879,N_12822);
or U15932 (N_15932,N_13533,N_12316);
nor U15933 (N_15933,N_12952,N_13320);
nand U15934 (N_15934,N_12438,N_13857);
xor U15935 (N_15935,N_12182,N_13053);
or U15936 (N_15936,N_12357,N_12197);
nand U15937 (N_15937,N_13673,N_13284);
xnor U15938 (N_15938,N_13195,N_12604);
and U15939 (N_15939,N_13814,N_13378);
and U15940 (N_15940,N_13551,N_12267);
nor U15941 (N_15941,N_13023,N_13496);
nand U15942 (N_15942,N_13377,N_13438);
and U15943 (N_15943,N_13695,N_13835);
nor U15944 (N_15944,N_13299,N_13916);
nor U15945 (N_15945,N_13964,N_12504);
and U15946 (N_15946,N_13984,N_13009);
xnor U15947 (N_15947,N_13682,N_12789);
nand U15948 (N_15948,N_12445,N_13285);
and U15949 (N_15949,N_12899,N_12199);
nor U15950 (N_15950,N_12236,N_12863);
xor U15951 (N_15951,N_12454,N_13114);
xor U15952 (N_15952,N_13458,N_12856);
and U15953 (N_15953,N_12380,N_12916);
or U15954 (N_15954,N_12901,N_13269);
nand U15955 (N_15955,N_13494,N_13339);
nand U15956 (N_15956,N_12667,N_13685);
nor U15957 (N_15957,N_12491,N_13934);
nor U15958 (N_15958,N_12329,N_13838);
xor U15959 (N_15959,N_12340,N_13772);
or U15960 (N_15960,N_12061,N_12203);
nor U15961 (N_15961,N_12674,N_12049);
nand U15962 (N_15962,N_12051,N_12478);
and U15963 (N_15963,N_12416,N_13129);
and U15964 (N_15964,N_13010,N_12127);
or U15965 (N_15965,N_12909,N_13939);
and U15966 (N_15966,N_12481,N_12641);
nor U15967 (N_15967,N_12215,N_12619);
nand U15968 (N_15968,N_12212,N_13729);
nand U15969 (N_15969,N_12592,N_12542);
or U15970 (N_15970,N_12682,N_12538);
nor U15971 (N_15971,N_13039,N_13701);
and U15972 (N_15972,N_12823,N_13118);
or U15973 (N_15973,N_12426,N_12081);
xor U15974 (N_15974,N_12732,N_12397);
nor U15975 (N_15975,N_13331,N_12448);
or U15976 (N_15976,N_12901,N_13016);
and U15977 (N_15977,N_12096,N_12410);
nand U15978 (N_15978,N_12929,N_12331);
and U15979 (N_15979,N_12623,N_13882);
xor U15980 (N_15980,N_12809,N_12390);
and U15981 (N_15981,N_12029,N_13311);
and U15982 (N_15982,N_13172,N_12384);
and U15983 (N_15983,N_13233,N_13422);
nor U15984 (N_15984,N_12851,N_13459);
xnor U15985 (N_15985,N_12808,N_13662);
nor U15986 (N_15986,N_13085,N_12446);
nand U15987 (N_15987,N_13840,N_12388);
and U15988 (N_15988,N_12515,N_13389);
or U15989 (N_15989,N_12388,N_13738);
nor U15990 (N_15990,N_12846,N_13836);
or U15991 (N_15991,N_13589,N_12840);
and U15992 (N_15992,N_13439,N_12850);
nand U15993 (N_15993,N_12648,N_12397);
nand U15994 (N_15994,N_12154,N_13318);
or U15995 (N_15995,N_12832,N_13675);
or U15996 (N_15996,N_12241,N_13117);
and U15997 (N_15997,N_12775,N_13681);
nor U15998 (N_15998,N_13264,N_12134);
xnor U15999 (N_15999,N_13209,N_13365);
xor U16000 (N_16000,N_14424,N_14796);
or U16001 (N_16001,N_14539,N_15952);
nand U16002 (N_16002,N_15075,N_14713);
or U16003 (N_16003,N_15712,N_14377);
xor U16004 (N_16004,N_15532,N_15426);
or U16005 (N_16005,N_14008,N_14920);
or U16006 (N_16006,N_15269,N_14064);
nor U16007 (N_16007,N_14396,N_14432);
and U16008 (N_16008,N_14697,N_15924);
or U16009 (N_16009,N_14642,N_14020);
xnor U16010 (N_16010,N_15962,N_15812);
nand U16011 (N_16011,N_15583,N_14669);
xnor U16012 (N_16012,N_15702,N_15987);
and U16013 (N_16013,N_14726,N_14462);
or U16014 (N_16014,N_15415,N_15997);
nor U16015 (N_16015,N_14223,N_15796);
and U16016 (N_16016,N_14908,N_15528);
nand U16017 (N_16017,N_15525,N_14698);
nor U16018 (N_16018,N_14655,N_15916);
nor U16019 (N_16019,N_14932,N_15259);
nor U16020 (N_16020,N_15792,N_14980);
nand U16021 (N_16021,N_15331,N_15040);
xnor U16022 (N_16022,N_14962,N_14944);
xnor U16023 (N_16023,N_14525,N_14488);
nor U16024 (N_16024,N_15939,N_15563);
nor U16025 (N_16025,N_14171,N_15582);
xnor U16026 (N_16026,N_15758,N_15300);
nand U16027 (N_16027,N_14004,N_14670);
and U16028 (N_16028,N_15615,N_14092);
nor U16029 (N_16029,N_14493,N_15188);
or U16030 (N_16030,N_14125,N_15743);
and U16031 (N_16031,N_14343,N_15646);
and U16032 (N_16032,N_15619,N_14138);
xnor U16033 (N_16033,N_15233,N_15690);
or U16034 (N_16034,N_14904,N_15840);
nand U16035 (N_16035,N_15598,N_15481);
xor U16036 (N_16036,N_15340,N_14659);
nor U16037 (N_16037,N_15904,N_15310);
nor U16038 (N_16038,N_15291,N_14498);
or U16039 (N_16039,N_14351,N_15096);
nand U16040 (N_16040,N_14985,N_14452);
xor U16041 (N_16041,N_14835,N_14853);
nand U16042 (N_16042,N_14286,N_14666);
and U16043 (N_16043,N_14943,N_14194);
xnor U16044 (N_16044,N_14584,N_15375);
xnor U16045 (N_16045,N_15492,N_14549);
nor U16046 (N_16046,N_14618,N_14088);
nand U16047 (N_16047,N_15860,N_14271);
or U16048 (N_16048,N_14316,N_15482);
nand U16049 (N_16049,N_15465,N_15639);
or U16050 (N_16050,N_14490,N_14024);
xnor U16051 (N_16051,N_15317,N_14550);
nand U16052 (N_16052,N_15377,N_15342);
or U16053 (N_16053,N_14656,N_15183);
and U16054 (N_16054,N_15795,N_14800);
or U16055 (N_16055,N_15202,N_15436);
or U16056 (N_16056,N_14945,N_15098);
xnor U16057 (N_16057,N_14581,N_15651);
or U16058 (N_16058,N_14610,N_15894);
and U16059 (N_16059,N_15210,N_15955);
nand U16060 (N_16060,N_15235,N_15884);
nor U16061 (N_16061,N_14863,N_15655);
nand U16062 (N_16062,N_14443,N_15130);
nand U16063 (N_16063,N_15455,N_15029);
nand U16064 (N_16064,N_14395,N_14535);
or U16065 (N_16065,N_14645,N_15006);
or U16066 (N_16066,N_15268,N_15156);
and U16067 (N_16067,N_14155,N_14891);
xor U16068 (N_16068,N_15921,N_14249);
xor U16069 (N_16069,N_14999,N_14942);
nor U16070 (N_16070,N_14455,N_15391);
or U16071 (N_16071,N_14928,N_14570);
and U16072 (N_16072,N_14430,N_14255);
nor U16073 (N_16073,N_14187,N_15135);
and U16074 (N_16074,N_14021,N_14977);
xor U16075 (N_16075,N_14912,N_14494);
xor U16076 (N_16076,N_14522,N_14289);
xnor U16077 (N_16077,N_15345,N_15679);
nand U16078 (N_16078,N_14317,N_14858);
and U16079 (N_16079,N_15585,N_14700);
nand U16080 (N_16080,N_15283,N_14299);
nor U16081 (N_16081,N_15402,N_15044);
or U16082 (N_16082,N_14056,N_15204);
and U16083 (N_16083,N_14936,N_14449);
nor U16084 (N_16084,N_14164,N_14716);
and U16085 (N_16085,N_15879,N_15062);
and U16086 (N_16086,N_14690,N_15666);
xnor U16087 (N_16087,N_15799,N_15922);
nand U16088 (N_16088,N_15733,N_14414);
nand U16089 (N_16089,N_15024,N_14173);
and U16090 (N_16090,N_15963,N_14308);
and U16091 (N_16091,N_15989,N_15330);
and U16092 (N_16092,N_15520,N_15947);
nand U16093 (N_16093,N_14120,N_14189);
and U16094 (N_16094,N_15530,N_14634);
or U16095 (N_16095,N_14394,N_14224);
or U16096 (N_16096,N_15087,N_14495);
nor U16097 (N_16097,N_15049,N_15635);
or U16098 (N_16098,N_15439,N_15643);
or U16099 (N_16099,N_14709,N_14210);
nand U16100 (N_16100,N_14941,N_15086);
nor U16101 (N_16101,N_15236,N_14680);
or U16102 (N_16102,N_15606,N_15027);
nor U16103 (N_16103,N_15322,N_15241);
xor U16104 (N_16104,N_14433,N_15009);
nand U16105 (N_16105,N_15373,N_15901);
and U16106 (N_16106,N_14112,N_15010);
or U16107 (N_16107,N_14346,N_14459);
or U16108 (N_16108,N_15416,N_15282);
nand U16109 (N_16109,N_14970,N_15853);
nor U16110 (N_16110,N_14244,N_15247);
nor U16111 (N_16111,N_15015,N_15621);
or U16112 (N_16112,N_15461,N_14415);
nand U16113 (N_16113,N_14053,N_15638);
and U16114 (N_16114,N_15554,N_15862);
nand U16115 (N_16115,N_14267,N_15320);
xor U16116 (N_16116,N_15943,N_14180);
and U16117 (N_16117,N_14751,N_15677);
and U16118 (N_16118,N_15699,N_14429);
or U16119 (N_16119,N_14009,N_15326);
xor U16120 (N_16120,N_14184,N_15155);
xnor U16121 (N_16121,N_15116,N_15034);
nor U16122 (N_16122,N_15097,N_15669);
or U16123 (N_16123,N_14016,N_15703);
xnor U16124 (N_16124,N_15008,N_14453);
xor U16125 (N_16125,N_15036,N_15389);
nand U16126 (N_16126,N_15052,N_14534);
nand U16127 (N_16127,N_15101,N_15307);
nor U16128 (N_16128,N_15208,N_14178);
xnor U16129 (N_16129,N_15986,N_15581);
nor U16130 (N_16130,N_14695,N_14901);
nor U16131 (N_16131,N_14843,N_15608);
nand U16132 (N_16132,N_15789,N_14597);
and U16133 (N_16133,N_14090,N_15216);
and U16134 (N_16134,N_14134,N_14815);
and U16135 (N_16135,N_14593,N_15452);
nor U16136 (N_16136,N_15944,N_15025);
nand U16137 (N_16137,N_15542,N_14717);
xnor U16138 (N_16138,N_15765,N_14849);
or U16139 (N_16139,N_14010,N_14371);
and U16140 (N_16140,N_14362,N_15493);
or U16141 (N_16141,N_14294,N_15467);
nor U16142 (N_16142,N_14756,N_14313);
and U16143 (N_16143,N_15763,N_14761);
nor U16144 (N_16144,N_15013,N_14935);
nand U16145 (N_16145,N_15736,N_14086);
nand U16146 (N_16146,N_15256,N_14297);
xor U16147 (N_16147,N_14794,N_15411);
and U16148 (N_16148,N_15772,N_14749);
nand U16149 (N_16149,N_15321,N_14589);
nand U16150 (N_16150,N_15141,N_14026);
nand U16151 (N_16151,N_14934,N_15961);
nor U16152 (N_16152,N_14334,N_15577);
xor U16153 (N_16153,N_14620,N_15738);
nand U16154 (N_16154,N_14003,N_14132);
or U16155 (N_16155,N_14614,N_14206);
xnor U16156 (N_16156,N_14917,N_14623);
and U16157 (N_16157,N_15475,N_15578);
nand U16158 (N_16158,N_15149,N_14781);
and U16159 (N_16159,N_14091,N_14662);
xnor U16160 (N_16160,N_15037,N_15797);
and U16161 (N_16161,N_14583,N_14520);
or U16162 (N_16162,N_15223,N_15565);
nor U16163 (N_16163,N_15447,N_14885);
xor U16164 (N_16164,N_14875,N_15787);
or U16165 (N_16165,N_15337,N_15936);
and U16166 (N_16166,N_15382,N_15502);
and U16167 (N_16167,N_15880,N_14261);
or U16168 (N_16168,N_14409,N_15238);
nand U16169 (N_16169,N_14532,N_14950);
nand U16170 (N_16170,N_15686,N_14473);
and U16171 (N_16171,N_15122,N_14119);
nand U16172 (N_16172,N_15773,N_14191);
nor U16173 (N_16173,N_15984,N_15403);
nand U16174 (N_16174,N_14504,N_14306);
nor U16175 (N_16175,N_14197,N_14454);
or U16176 (N_16176,N_14046,N_14959);
xor U16177 (N_16177,N_14325,N_15591);
nand U16178 (N_16178,N_14152,N_14921);
and U16179 (N_16179,N_14651,N_14693);
or U16180 (N_16180,N_14890,N_14233);
or U16181 (N_16181,N_14611,N_14207);
or U16182 (N_16182,N_15129,N_14186);
and U16183 (N_16183,N_14257,N_14675);
and U16184 (N_16184,N_14032,N_15151);
xor U16185 (N_16185,N_14211,N_14365);
nand U16186 (N_16186,N_14837,N_14661);
nor U16187 (N_16187,N_15140,N_15038);
and U16188 (N_16188,N_15804,N_14332);
or U16189 (N_16189,N_15000,N_15705);
xor U16190 (N_16190,N_14270,N_14410);
nand U16191 (N_16191,N_14804,N_14467);
xor U16192 (N_16192,N_15971,N_14688);
nand U16193 (N_16193,N_14169,N_14949);
nor U16194 (N_16194,N_14038,N_15991);
nor U16195 (N_16195,N_15350,N_14911);
and U16196 (N_16196,N_14353,N_15248);
nand U16197 (N_16197,N_14636,N_14340);
nor U16198 (N_16198,N_15304,N_15381);
and U16199 (N_16199,N_14701,N_15338);
nor U16200 (N_16200,N_15127,N_14657);
xor U16201 (N_16201,N_14141,N_15771);
or U16202 (N_16202,N_14392,N_15668);
nand U16203 (N_16203,N_15616,N_15275);
and U16204 (N_16204,N_14547,N_15464);
nor U16205 (N_16205,N_15001,N_14451);
nand U16206 (N_16206,N_14710,N_15510);
or U16207 (N_16207,N_14083,N_15665);
xor U16208 (N_16208,N_15294,N_15566);
nor U16209 (N_16209,N_15061,N_14914);
or U16210 (N_16210,N_15301,N_14412);
and U16211 (N_16211,N_15158,N_15995);
nand U16212 (N_16212,N_15656,N_14456);
nand U16213 (N_16213,N_15254,N_15480);
or U16214 (N_16214,N_14879,N_15169);
xor U16215 (N_16215,N_14407,N_15740);
xor U16216 (N_16216,N_14280,N_14314);
nand U16217 (N_16217,N_15245,N_14627);
and U16218 (N_16218,N_15746,N_15888);
and U16219 (N_16219,N_14007,N_14981);
nand U16220 (N_16220,N_15430,N_15752);
nor U16221 (N_16221,N_15325,N_15735);
nand U16222 (N_16222,N_14357,N_15385);
nor U16223 (N_16223,N_14384,N_14703);
nor U16224 (N_16224,N_15309,N_15339);
or U16225 (N_16225,N_15166,N_15045);
nor U16226 (N_16226,N_15640,N_14438);
nand U16227 (N_16227,N_14577,N_15343);
xnor U16228 (N_16228,N_14100,N_14747);
and U16229 (N_16229,N_14696,N_15368);
or U16230 (N_16230,N_15095,N_14876);
or U16231 (N_16231,N_14375,N_15867);
nand U16232 (N_16232,N_14420,N_14296);
xor U16233 (N_16233,N_15004,N_15653);
nand U16234 (N_16234,N_14199,N_14530);
nor U16235 (N_16235,N_14059,N_14093);
and U16236 (N_16236,N_15200,N_14587);
xor U16237 (N_16237,N_15648,N_14102);
nor U16238 (N_16238,N_14905,N_15196);
or U16239 (N_16239,N_15393,N_15568);
and U16240 (N_16240,N_14201,N_14531);
nor U16241 (N_16241,N_14312,N_14916);
nand U16242 (N_16242,N_15890,N_15866);
and U16243 (N_16243,N_14505,N_15246);
and U16244 (N_16244,N_14050,N_14826);
nor U16245 (N_16245,N_14877,N_14888);
nand U16246 (N_16246,N_15114,N_15965);
nor U16247 (N_16247,N_14082,N_15546);
xnor U16248 (N_16248,N_14964,N_15637);
nand U16249 (N_16249,N_15280,N_15413);
and U16250 (N_16250,N_15572,N_14315);
xnor U16251 (N_16251,N_14735,N_15126);
xnor U16252 (N_16252,N_14291,N_15976);
and U16253 (N_16253,N_15891,N_14813);
nand U16254 (N_16254,N_15460,N_15312);
nand U16255 (N_16255,N_14881,N_14247);
or U16256 (N_16256,N_14436,N_14418);
xnor U16257 (N_16257,N_14519,N_14963);
nand U16258 (N_16258,N_14730,N_15769);
nor U16259 (N_16259,N_15448,N_14033);
and U16260 (N_16260,N_15687,N_14886);
and U16261 (N_16261,N_14622,N_15975);
nor U16262 (N_16262,N_14209,N_15704);
or U16263 (N_16263,N_15897,N_14724);
and U16264 (N_16264,N_15993,N_15070);
nor U16265 (N_16265,N_14445,N_15555);
nand U16266 (N_16266,N_15323,N_14148);
and U16267 (N_16267,N_14967,N_15611);
nor U16268 (N_16268,N_15220,N_15770);
xor U16269 (N_16269,N_14071,N_15833);
or U16270 (N_16270,N_14218,N_15082);
nor U16271 (N_16271,N_15016,N_14660);
or U16272 (N_16272,N_15764,N_15443);
nand U16273 (N_16273,N_15721,N_14869);
xor U16274 (N_16274,N_14250,N_14857);
nor U16275 (N_16275,N_15819,N_14615);
nand U16276 (N_16276,N_14567,N_15173);
nand U16277 (N_16277,N_14476,N_15751);
nand U16278 (N_16278,N_14135,N_15861);
nor U16279 (N_16279,N_15685,N_15234);
nand U16280 (N_16280,N_14202,N_15556);
or U16281 (N_16281,N_14711,N_15816);
or U16282 (N_16282,N_14108,N_15881);
nand U16283 (N_16283,N_14416,N_15980);
nor U16284 (N_16284,N_14236,N_14447);
nand U16285 (N_16285,N_14245,N_15485);
or U16286 (N_16286,N_15949,N_14149);
and U16287 (N_16287,N_14075,N_14425);
and U16288 (N_16288,N_15755,N_15418);
nor U16289 (N_16289,N_14692,N_15967);
nor U16290 (N_16290,N_14281,N_14130);
nor U16291 (N_16291,N_15263,N_15698);
nand U16292 (N_16292,N_14159,N_14128);
or U16293 (N_16293,N_14385,N_14041);
or U16294 (N_16294,N_14689,N_15002);
or U16295 (N_16295,N_14907,N_14774);
nand U16296 (N_16296,N_14569,N_14952);
or U16297 (N_16297,N_15023,N_14256);
nor U16298 (N_16298,N_14227,N_15371);
nand U16299 (N_16299,N_15454,N_14328);
nor U16300 (N_16300,N_14933,N_14938);
nand U16301 (N_16301,N_14176,N_14491);
nand U16302 (N_16302,N_15194,N_15931);
and U16303 (N_16303,N_15588,N_14242);
nor U16304 (N_16304,N_14025,N_14744);
nand U16305 (N_16305,N_15815,N_15078);
and U16306 (N_16306,N_14573,N_14366);
nand U16307 (N_16307,N_15663,N_15620);
xor U16308 (N_16308,N_15868,N_14354);
and U16309 (N_16309,N_14789,N_15761);
or U16310 (N_16310,N_15741,N_14262);
or U16311 (N_16311,N_14345,N_14166);
nor U16312 (N_16312,N_15298,N_14376);
nand U16313 (N_16313,N_15693,N_14860);
nor U16314 (N_16314,N_14198,N_15882);
nand U16315 (N_16315,N_15131,N_14419);
or U16316 (N_16316,N_14402,N_14607);
xor U16317 (N_16317,N_14983,N_15473);
and U16318 (N_16318,N_14464,N_14553);
or U16319 (N_16319,N_14598,N_14926);
nor U16320 (N_16320,N_15344,N_14827);
nand U16321 (N_16321,N_14533,N_14542);
nand U16322 (N_16322,N_15192,N_14819);
and U16323 (N_16323,N_14892,N_14285);
and U16324 (N_16324,N_14027,N_15111);
and U16325 (N_16325,N_15242,N_15933);
and U16326 (N_16326,N_15725,N_14958);
nor U16327 (N_16327,N_15251,N_14554);
and U16328 (N_16328,N_14563,N_15011);
nand U16329 (N_16329,N_15274,N_14292);
nor U16330 (N_16330,N_15333,N_15435);
nor U16331 (N_16331,N_14327,N_15032);
or U16332 (N_16332,N_14105,N_14903);
xnor U16333 (N_16333,N_15273,N_14302);
xor U16334 (N_16334,N_15354,N_15970);
xnor U16335 (N_16335,N_14600,N_15123);
nor U16336 (N_16336,N_14763,N_15424);
and U16337 (N_16337,N_15186,N_14874);
and U16338 (N_16338,N_14682,N_14671);
xnor U16339 (N_16339,N_15187,N_15745);
xnor U16340 (N_16340,N_14040,N_15491);
nand U16341 (N_16341,N_15564,N_15946);
xor U16342 (N_16342,N_15077,N_15596);
nand U16343 (N_16343,N_15734,N_15658);
nor U16344 (N_16344,N_14168,N_14954);
nand U16345 (N_16345,N_14831,N_14864);
and U16346 (N_16346,N_15033,N_14946);
nor U16347 (N_16347,N_15361,N_15831);
nor U16348 (N_16348,N_15297,N_14183);
nor U16349 (N_16349,N_15171,N_15811);
nor U16350 (N_16350,N_15412,N_15278);
xnor U16351 (N_16351,N_15243,N_15453);
nor U16352 (N_16352,N_14558,N_15311);
and U16353 (N_16353,N_14324,N_14548);
xor U16354 (N_16354,N_15570,N_15896);
and U16355 (N_16355,N_15903,N_14431);
or U16356 (N_16356,N_14783,N_14764);
or U16357 (N_16357,N_14018,N_15524);
and U16358 (N_16358,N_14214,N_15213);
nand U16359 (N_16359,N_14736,N_14014);
and U16360 (N_16360,N_14626,N_14940);
nor U16361 (N_16361,N_14859,N_14768);
nand U16362 (N_16362,N_15364,N_14497);
xnor U16363 (N_16363,N_14140,N_15641);
nand U16364 (N_16364,N_15526,N_14413);
nand U16365 (N_16365,N_14617,N_14672);
or U16366 (N_16366,N_14582,N_15226);
nor U16367 (N_16367,N_14011,N_14708);
xnor U16368 (N_16368,N_14323,N_15346);
nand U16369 (N_16369,N_14422,N_14400);
xor U16370 (N_16370,N_14821,N_14537);
xnor U16371 (N_16371,N_14485,N_14792);
or U16372 (N_16372,N_15514,N_14188);
nor U16373 (N_16373,N_15406,N_15938);
or U16374 (N_16374,N_14643,N_15807);
or U16375 (N_16375,N_15372,N_15821);
or U16376 (N_16376,N_15429,N_15231);
nor U16377 (N_16377,N_15654,N_15817);
nand U16378 (N_16378,N_14992,N_15162);
xor U16379 (N_16379,N_15031,N_15912);
xnor U16380 (N_16380,N_15914,N_14157);
nand U16381 (N_16381,N_14028,N_14918);
xnor U16382 (N_16382,N_15607,N_15864);
and U16383 (N_16383,N_14117,N_14369);
and U16384 (N_16384,N_14975,N_14096);
or U16385 (N_16385,N_14062,N_14095);
and U16386 (N_16386,N_15966,N_15545);
xnor U16387 (N_16387,N_14068,N_15314);
or U16388 (N_16388,N_15915,N_14367);
and U16389 (N_16389,N_15329,N_15700);
nand U16390 (N_16390,N_14702,N_15762);
or U16391 (N_16391,N_14805,N_15165);
and U16392 (N_16392,N_15255,N_15053);
xnor U16393 (N_16393,N_14665,N_14674);
nand U16394 (N_16394,N_14103,N_14889);
and U16395 (N_16395,N_15749,N_15613);
nand U16396 (N_16396,N_14755,N_15422);
nand U16397 (N_16397,N_15295,N_14023);
and U16398 (N_16398,N_15253,N_14240);
xor U16399 (N_16399,N_14536,N_15875);
or U16400 (N_16400,N_14521,N_15468);
nor U16401 (N_16401,N_15674,N_14254);
xnor U16402 (N_16402,N_14374,N_14741);
nor U16403 (N_16403,N_14144,N_14825);
nor U16404 (N_16404,N_15533,N_15369);
nor U16405 (N_16405,N_15920,N_15522);
or U16406 (N_16406,N_14044,N_14591);
xor U16407 (N_16407,N_14580,N_14733);
xnor U16408 (N_16408,N_15985,N_14423);
xnor U16409 (N_16409,N_15800,N_15215);
or U16410 (N_16410,N_14398,N_15292);
and U16411 (N_16411,N_15190,N_15929);
and U16412 (N_16412,N_15272,N_14212);
nand U16413 (N_16413,N_14760,N_14871);
and U16414 (N_16414,N_14274,N_15137);
nand U16415 (N_16415,N_14668,N_14808);
or U16416 (N_16416,N_15713,N_15678);
or U16417 (N_16417,N_15232,N_14143);
and U16418 (N_16418,N_15571,N_15541);
nand U16419 (N_16419,N_14508,N_14237);
or U16420 (N_16420,N_14426,N_14571);
nor U16421 (N_16421,N_14506,N_15444);
and U16422 (N_16422,N_15604,N_14277);
xor U16423 (N_16423,N_15163,N_15394);
nor U16424 (N_16424,N_15209,N_14704);
and U16425 (N_16425,N_15100,N_15113);
and U16426 (N_16426,N_15205,N_15632);
nor U16427 (N_16427,N_14797,N_14965);
nand U16428 (N_16428,N_15125,N_15237);
or U16429 (N_16429,N_14080,N_14336);
nor U16430 (N_16430,N_15917,N_14200);
and U16431 (N_16431,N_15121,N_14727);
nor U16432 (N_16432,N_14370,N_15265);
xnor U16433 (N_16433,N_15872,N_15780);
nand U16434 (N_16434,N_15146,N_14646);
nor U16435 (N_16435,N_14639,N_15617);
nor U16436 (N_16436,N_15737,N_14195);
nor U16437 (N_16437,N_14116,N_15108);
xor U16438 (N_16438,N_14993,N_14440);
xor U16439 (N_16439,N_15661,N_15644);
or U16440 (N_16440,N_14382,N_14560);
or U16441 (N_16441,N_14818,N_15355);
nand U16442 (N_16442,N_15516,N_14264);
nand U16443 (N_16443,N_14087,N_15992);
and U16444 (N_16444,N_15334,N_15509);
nor U16445 (N_16445,N_15094,N_14812);
nor U16446 (N_16446,N_14074,N_15396);
xnor U16447 (N_16447,N_15018,N_14060);
nand U16448 (N_16448,N_15826,N_14439);
nor U16449 (N_16449,N_15488,N_15513);
and U16450 (N_16450,N_15064,N_14785);
and U16451 (N_16451,N_14552,N_15595);
nand U16452 (N_16452,N_15449,N_15701);
xor U16453 (N_16453,N_14851,N_14300);
nor U16454 (N_16454,N_15539,N_15281);
nor U16455 (N_16455,N_15080,N_15470);
and U16456 (N_16456,N_15562,N_15120);
nor U16457 (N_16457,N_15768,N_14241);
nand U16458 (N_16458,N_15074,N_15362);
and U16459 (N_16459,N_15534,N_14182);
nand U16460 (N_16460,N_15636,N_14192);
and U16461 (N_16461,N_15494,N_14017);
nand U16462 (N_16462,N_15197,N_15567);
or U16463 (N_16463,N_14216,N_14019);
or U16464 (N_16464,N_14585,N_15747);
xnor U16465 (N_16465,N_14349,N_15547);
xnor U16466 (N_16466,N_14121,N_14801);
xnor U16467 (N_16467,N_14106,N_14609);
or U16468 (N_16468,N_15090,N_15252);
and U16469 (N_16469,N_14486,N_14720);
or U16470 (N_16470,N_14356,N_15221);
nand U16471 (N_16471,N_14854,N_14790);
or U16472 (N_16472,N_15118,N_15561);
and U16473 (N_16473,N_14765,N_15089);
xor U16474 (N_16474,N_14404,N_14619);
and U16475 (N_16475,N_14273,N_14605);
or U16476 (N_16476,N_14097,N_15782);
and U16477 (N_16477,N_14731,N_14806);
xnor U16478 (N_16478,N_15791,N_14960);
or U16479 (N_16479,N_15843,N_14406);
or U16480 (N_16480,N_14780,N_15498);
xnor U16481 (N_16481,N_15594,N_14156);
nand U16482 (N_16482,N_15612,N_15136);
nor U16483 (N_16483,N_14867,N_14947);
or U16484 (N_16484,N_15774,N_15718);
or U16485 (N_16485,N_14559,N_15115);
or U16486 (N_16486,N_15172,N_15633);
xnor U16487 (N_16487,N_15844,N_14442);
nand U16488 (N_16488,N_14725,N_15557);
xor U16489 (N_16489,N_14978,N_15979);
or U16490 (N_16490,N_14740,N_15072);
nand U16491 (N_16491,N_15692,N_15388);
and U16492 (N_16492,N_14880,N_14971);
nand U16493 (N_16493,N_15353,N_15732);
nand U16494 (N_16494,N_14883,N_14239);
xnor U16495 (N_16495,N_15626,N_14759);
nand U16496 (N_16496,N_15580,N_15047);
nand U16497 (N_16497,N_15257,N_14070);
and U16498 (N_16498,N_14715,N_15964);
and U16499 (N_16499,N_14061,N_15073);
nor U16500 (N_16500,N_14109,N_14150);
or U16501 (N_16501,N_14047,N_14363);
nor U16502 (N_16502,N_15726,N_14172);
nor U16503 (N_16503,N_14072,N_15240);
and U16504 (N_16504,N_14984,N_14850);
nor U16505 (N_16505,N_15974,N_15174);
xor U16506 (N_16506,N_15676,N_15569);
nor U16507 (N_16507,N_15709,N_14364);
or U16508 (N_16508,N_15066,N_14006);
nor U16509 (N_16509,N_14997,N_15261);
xnor U16510 (N_16510,N_15214,N_14807);
nor U16511 (N_16511,N_15757,N_15442);
or U16512 (N_16512,N_15390,N_14865);
or U16513 (N_16513,N_14217,N_14810);
or U16514 (N_16514,N_14745,N_15825);
or U16515 (N_16515,N_15998,N_15012);
nor U16516 (N_16516,N_14750,N_15652);
nand U16517 (N_16517,N_15184,N_14101);
nand U16518 (N_16518,N_14786,N_15508);
nor U16519 (N_16519,N_15405,N_15065);
or U16520 (N_16520,N_15863,N_15722);
or U16521 (N_16521,N_14652,N_14397);
and U16522 (N_16522,N_15206,N_14145);
and U16523 (N_16523,N_14359,N_15303);
or U16524 (N_16524,N_15558,N_15328);
nand U16525 (N_16525,N_14995,N_15667);
xnor U16526 (N_16526,N_15942,N_15332);
nand U16527 (N_16527,N_14177,N_15048);
and U16528 (N_16528,N_15907,N_15289);
xor U16529 (N_16529,N_15370,N_15871);
nor U16530 (N_16530,N_14654,N_14146);
nor U16531 (N_16531,N_14649,N_15848);
xnor U16532 (N_16532,N_15968,N_15590);
nor U16533 (N_16533,N_15739,N_14284);
nand U16534 (N_16534,N_15505,N_15544);
and U16535 (N_16535,N_15822,N_15398);
nand U16536 (N_16536,N_15540,N_14778);
or U16537 (N_16537,N_14243,N_15483);
or U16538 (N_16538,N_15150,N_15729);
and U16539 (N_16539,N_14979,N_14136);
and U16540 (N_16540,N_15463,N_14896);
xor U16541 (N_16541,N_14321,N_15076);
nor U16542 (N_16542,N_15176,N_15927);
and U16543 (N_16543,N_14699,N_14906);
nand U16544 (N_16544,N_15978,N_15972);
and U16545 (N_16545,N_14753,N_14540);
nand U16546 (N_16546,N_14893,N_14151);
and U16547 (N_16547,N_14076,N_14077);
and U16548 (N_16548,N_14721,N_15079);
and U16549 (N_16549,N_15602,N_15576);
nor U16550 (N_16550,N_14085,N_14293);
xor U16551 (N_16551,N_14803,N_14546);
nand U16552 (N_16552,N_14722,N_15809);
and U16553 (N_16553,N_14909,N_14127);
and U16554 (N_16554,N_15645,N_14602);
nor U16555 (N_16555,N_14311,N_15610);
xor U16556 (N_16556,N_15711,N_14283);
nand U16557 (N_16557,N_15625,N_14002);
and U16558 (N_16558,N_14931,N_15551);
or U16559 (N_16559,N_14089,N_14079);
nand U16560 (N_16560,N_14973,N_14408);
xor U16561 (N_16561,N_14625,N_15021);
or U16562 (N_16562,N_14969,N_15911);
nor U16563 (N_16563,N_14196,N_15781);
nor U16564 (N_16564,N_14322,N_14518);
or U16565 (N_16565,N_14204,N_15306);
or U16566 (N_16566,N_15808,N_15177);
xor U16567 (N_16567,N_14603,N_15271);
or U16568 (N_16568,N_14956,N_15456);
or U16569 (N_16569,N_15478,N_15587);
or U16570 (N_16570,N_15543,N_15983);
xnor U16571 (N_16571,N_15586,N_15068);
xnor U16572 (N_16572,N_14922,N_14923);
xor U16573 (N_16573,N_14350,N_15858);
xor U16574 (N_16574,N_14167,N_15103);
and U16575 (N_16575,N_14222,N_14870);
or U16576 (N_16576,N_14809,N_15058);
or U16577 (N_16577,N_15417,N_14986);
or U16578 (N_16578,N_14746,N_14052);
or U16579 (N_16579,N_15662,N_15727);
xor U16580 (N_16580,N_14953,N_15940);
or U16581 (N_16581,N_15348,N_15553);
nor U16582 (N_16582,N_14094,N_15117);
xnor U16583 (N_16583,N_14544,N_14579);
nand U16584 (N_16584,N_15497,N_15603);
nand U16585 (N_16585,N_14872,N_14225);
or U16586 (N_16586,N_14595,N_15105);
and U16587 (N_16587,N_14644,N_15753);
and U16588 (N_16588,N_15874,N_14824);
nand U16589 (N_16589,N_15697,N_15358);
nand U16590 (N_16590,N_15446,N_15512);
nor U16591 (N_16591,N_14814,N_14976);
and U16592 (N_16592,N_14887,N_15837);
or U16593 (N_16593,N_14830,N_14787);
or U16594 (N_16594,N_15500,N_14129);
or U16595 (N_16595,N_15056,N_15973);
or U16596 (N_16596,N_14673,N_14691);
or U16597 (N_16597,N_14502,N_14613);
xor U16598 (N_16598,N_15401,N_14499);
or U16599 (N_16599,N_15287,N_15723);
xor U16600 (N_16600,N_14503,N_15093);
nand U16601 (N_16601,N_15106,N_15883);
and U16602 (N_16602,N_14458,N_14919);
xor U16603 (N_16603,N_14939,N_14137);
nand U16604 (N_16604,N_15028,N_15457);
xnor U16605 (N_16605,N_14538,N_14477);
or U16606 (N_16606,N_14590,N_14450);
nand U16607 (N_16607,N_15849,N_14310);
and U16608 (N_16608,N_15951,N_15324);
nor U16609 (N_16609,N_15918,N_15395);
nor U16610 (N_16610,N_14913,N_15445);
nand U16611 (N_16611,N_15574,N_15597);
or U16612 (N_16612,N_14510,N_15486);
nor U16613 (N_16613,N_15956,N_14466);
nor U16614 (N_16614,N_15820,N_15785);
nor U16615 (N_16615,N_15438,N_15296);
and U16616 (N_16616,N_15928,N_14866);
nor U16617 (N_16617,N_15351,N_15941);
nand U16618 (N_16618,N_15144,N_14057);
nand U16619 (N_16619,N_15496,N_14001);
xor U16620 (N_16620,N_14592,N_14215);
xnor U16621 (N_16621,N_15694,N_15504);
or U16622 (N_16622,N_15293,N_15990);
or U16623 (N_16623,N_14303,N_15499);
nor U16624 (N_16624,N_15472,N_14739);
and U16625 (N_16625,N_15451,N_14160);
nor U16626 (N_16626,N_15828,N_14035);
or U16627 (N_16627,N_15876,N_15039);
nor U16628 (N_16628,N_15357,N_15537);
xnor U16629 (N_16629,N_14457,N_15776);
or U16630 (N_16630,N_15748,N_14653);
nand U16631 (N_16631,N_15627,N_15051);
nor U16632 (N_16632,N_15392,N_14681);
nor U16633 (N_16633,N_14344,N_14898);
or U16634 (N_16634,N_14378,N_15802);
nor U16635 (N_16635,N_14203,N_15829);
nand U16636 (N_16636,N_14358,N_14482);
nand U16637 (N_16637,N_14122,N_14335);
xor U16638 (N_16638,N_15950,N_15160);
and U16639 (N_16639,N_15476,N_14463);
nand U16640 (N_16640,N_15327,N_15731);
xor U16641 (N_16641,N_14073,N_14728);
xnor U16642 (N_16642,N_14162,N_15207);
xor U16643 (N_16643,N_15414,N_14873);
nor U16644 (N_16644,N_14678,N_15352);
and U16645 (N_16645,N_14427,N_14234);
and U16646 (N_16646,N_15277,N_15649);
and U16647 (N_16647,N_14469,N_14799);
and U16648 (N_16648,N_14638,N_14776);
nor U16649 (N_16649,N_14005,N_15302);
xnor U16650 (N_16650,N_14930,N_15400);
xor U16651 (N_16651,N_15664,N_15179);
or U16652 (N_16652,N_14347,N_15847);
and U16653 (N_16653,N_14480,N_14758);
and U16654 (N_16654,N_15258,N_15262);
nor U16655 (N_16655,N_14561,N_14528);
and U16656 (N_16656,N_14268,N_14855);
or U16657 (N_16657,N_15279,N_15407);
nand U16658 (N_16658,N_14968,N_15592);
nor U16659 (N_16659,N_14051,N_15462);
nor U16660 (N_16660,N_15379,N_15818);
nand U16661 (N_16661,N_14118,N_15181);
nor U16662 (N_16662,N_14368,N_14686);
nand U16663 (N_16663,N_14629,N_14706);
xor U16664 (N_16664,N_15286,N_15495);
and U16665 (N_16665,N_15614,N_15359);
nor U16666 (N_16666,N_15360,N_14446);
nand U16667 (N_16667,N_14219,N_14238);
or U16668 (N_16668,N_15019,N_14478);
nor U16669 (N_16669,N_15284,N_14228);
nand U16670 (N_16670,N_14460,N_14389);
xnor U16671 (N_16671,N_14966,N_14738);
or U16672 (N_16672,N_14705,N_15766);
and U16673 (N_16673,N_14034,N_14572);
nor U16674 (N_16674,N_14793,N_15088);
nor U16675 (N_16675,N_14820,N_14428);
or U16676 (N_16676,N_14836,N_15810);
or U16677 (N_16677,N_14361,N_15191);
and U16678 (N_16678,N_14337,N_14779);
nand U16679 (N_16679,N_15431,N_15474);
xnor U16680 (N_16680,N_15798,N_15175);
and U16681 (N_16681,N_15366,N_15926);
and U16682 (N_16682,N_15707,N_15601);
nand U16683 (N_16683,N_15906,N_14258);
xor U16684 (N_16684,N_14621,N_14265);
nor U16685 (N_16685,N_15624,N_14526);
or U16686 (N_16686,N_14320,N_14948);
nand U16687 (N_16687,N_15827,N_15779);
nor U16688 (N_16688,N_14846,N_14276);
xor U16689 (N_16689,N_15374,N_15788);
xnor U16690 (N_16690,N_15022,N_14326);
or U16691 (N_16691,N_14957,N_14513);
or U16692 (N_16692,N_14142,N_15441);
xnor U16693 (N_16693,N_15043,N_15691);
nand U16694 (N_16694,N_14996,N_14165);
nor U16695 (N_16695,N_14496,N_15182);
or U16696 (N_16696,N_14848,N_15425);
or U16697 (N_16697,N_15318,N_14015);
xor U16698 (N_16698,N_15249,N_15132);
or U16699 (N_16699,N_14220,N_14329);
xnor U16700 (N_16700,N_14042,N_14514);
nand U16701 (N_16701,N_15969,N_15218);
or U16702 (N_16702,N_15609,N_15201);
and U16703 (N_16703,N_14676,N_15290);
nor U16704 (N_16704,N_15689,N_14110);
nor U16705 (N_16705,N_14816,N_14489);
nand U16706 (N_16706,N_14856,N_15152);
or U16707 (N_16707,N_14288,N_15519);
nand U16708 (N_16708,N_15466,N_15315);
nor U16709 (N_16709,N_15139,N_15489);
nand U16710 (N_16710,N_14829,N_14507);
or U16711 (N_16711,N_14301,N_14754);
and U16712 (N_16712,N_14269,N_14266);
nor U16713 (N_16713,N_15316,N_14900);
nor U16714 (N_16714,N_14757,N_15856);
and U16715 (N_16715,N_15628,N_14055);
nor U16716 (N_16716,N_15178,N_14380);
nand U16717 (N_16717,N_14628,N_14330);
and U16718 (N_16718,N_14541,N_14599);
and U16719 (N_16719,N_14568,N_14512);
and U16720 (N_16720,N_14817,N_15285);
nor U16721 (N_16721,N_14078,N_14037);
nand U16722 (N_16722,N_15250,N_14065);
nor U16723 (N_16723,N_14461,N_14260);
nand U16724 (N_16724,N_14500,N_14472);
and U16725 (N_16725,N_15046,N_14471);
nand U16726 (N_16726,N_15133,N_15518);
or U16727 (N_16727,N_15511,N_14048);
or U16728 (N_16728,N_14099,N_15267);
nor U16729 (N_16729,N_15437,N_15842);
xor U16730 (N_16730,N_14383,N_14773);
nor U16731 (N_16731,N_15003,N_14190);
nand U16732 (N_16732,N_14213,N_14937);
nor U16733 (N_16733,N_14511,N_14246);
nand U16734 (N_16734,N_14987,N_14714);
nand U16735 (N_16735,N_15937,N_15092);
xor U16736 (N_16736,N_14732,N_15007);
xor U16737 (N_16737,N_15909,N_15948);
xor U16738 (N_16738,N_15650,N_14766);
xnor U16739 (N_16739,N_14578,N_14338);
or U16740 (N_16740,N_14683,N_15119);
xor U16741 (N_16741,N_15552,N_15957);
nand U16742 (N_16742,N_15754,N_15893);
nor U16743 (N_16743,N_15905,N_15124);
nor U16744 (N_16744,N_14632,N_15630);
or U16745 (N_16745,N_15716,N_15264);
nand U16746 (N_16746,N_14576,N_15803);
or U16747 (N_16747,N_14333,N_14586);
nor U16748 (N_16748,N_14282,N_15908);
or U16749 (N_16749,N_15109,N_15423);
nand U16750 (N_16750,N_15579,N_14902);
and U16751 (N_16751,N_15988,N_14054);
nor U16752 (N_16752,N_14718,N_15982);
or U16753 (N_16753,N_15618,N_14861);
or U16754 (N_16754,N_15839,N_15672);
or U16755 (N_16755,N_14307,N_15854);
or U16756 (N_16756,N_14982,N_15421);
or U16757 (N_16757,N_15996,N_14951);
xor U16758 (N_16758,N_15067,N_14601);
xnor U16759 (N_16759,N_14878,N_14972);
nand U16760 (N_16760,N_15521,N_15783);
xor U16761 (N_16761,N_15313,N_14441);
or U16762 (N_16762,N_15887,N_15767);
nor U16763 (N_16763,N_14465,N_15673);
xnor U16764 (N_16764,N_15835,N_15877);
nor U16765 (N_16765,N_14915,N_15549);
nand U16766 (N_16766,N_14492,N_15189);
nand U16767 (N_16767,N_15069,N_15230);
or U16768 (N_16768,N_14604,N_14232);
and U16769 (N_16769,N_15660,N_15222);
xnor U16770 (N_16770,N_15684,N_14153);
xor U16771 (N_16771,N_15459,N_14650);
nand U16772 (N_16772,N_14483,N_15410);
and U16773 (N_16773,N_14253,N_15180);
xor U16774 (N_16774,N_15659,N_14403);
and U16775 (N_16775,N_15035,N_14381);
and U16776 (N_16776,N_14862,N_14379);
nor U16777 (N_16777,N_15902,N_14252);
and U16778 (N_16778,N_14475,N_15977);
or U16779 (N_16779,N_15865,N_15376);
or U16780 (N_16780,N_14339,N_14565);
or U16781 (N_16781,N_15365,N_15288);
xnor U16782 (N_16782,N_15550,N_15305);
or U16783 (N_16783,N_15091,N_14107);
nor U16784 (N_16784,N_14596,N_15775);
nand U16785 (N_16785,N_15958,N_15212);
nor U16786 (N_16786,N_14897,N_15164);
nor U16787 (N_16787,N_15538,N_14748);
and U16788 (N_16788,N_15529,N_14179);
nand U16789 (N_16789,N_14484,N_15527);
nor U16790 (N_16790,N_15104,N_15851);
or U16791 (N_16791,N_14840,N_15107);
nand U16792 (N_16792,N_14635,N_15380);
or U16793 (N_16793,N_14111,N_14631);
and U16794 (N_16794,N_15134,N_14386);
or U16795 (N_16795,N_14743,N_15154);
xnor U16796 (N_16796,N_14181,N_14098);
or U16797 (N_16797,N_14828,N_14842);
nor U16798 (N_16798,N_15110,N_15657);
nand U16799 (N_16799,N_14557,N_14719);
xnor U16800 (N_16800,N_14290,N_15229);
nor U16801 (N_16801,N_15469,N_14272);
xor U16802 (N_16802,N_14998,N_14594);
nand U16803 (N_16803,N_14788,N_14043);
and U16804 (N_16804,N_15934,N_14133);
or U16805 (N_16805,N_14575,N_15560);
and U16806 (N_16806,N_14248,N_15777);
and U16807 (N_16807,N_14388,N_15953);
xnor U16808 (N_16808,N_15145,N_15599);
or U16809 (N_16809,N_15517,N_14304);
or U16810 (N_16810,N_15959,N_14263);
nor U16811 (N_16811,N_15085,N_15490);
nand U16812 (N_16812,N_14988,N_15889);
nor U16813 (N_16813,N_14648,N_14417);
nor U16814 (N_16814,N_14278,N_14468);
xnor U16815 (N_16815,N_14752,N_15805);
nand U16816 (N_16816,N_15193,N_14566);
nor U16817 (N_16817,N_15299,N_14124);
xor U16818 (N_16818,N_14448,N_15081);
or U16819 (N_16819,N_14927,N_14067);
xor U16820 (N_16820,N_15605,N_14515);
nand U16821 (N_16821,N_14139,N_14606);
nand U16822 (N_16822,N_14193,N_14235);
nor U16823 (N_16823,N_14154,N_15167);
xor U16824 (N_16824,N_14355,N_14066);
nor U16825 (N_16825,N_14298,N_15244);
or U16826 (N_16826,N_15720,N_14393);
or U16827 (N_16827,N_15487,N_14045);
nor U16828 (N_16828,N_14113,N_14523);
xor U16829 (N_16829,N_15593,N_14318);
and U16830 (N_16830,N_14275,N_15270);
nor U16831 (N_16831,N_15041,N_14685);
nor U16832 (N_16832,N_15960,N_14527);
nand U16833 (N_16833,N_15143,N_14707);
nor U16834 (N_16834,N_14974,N_15913);
nor U16835 (N_16835,N_15784,N_14158);
nand U16836 (N_16836,N_14147,N_15634);
or U16837 (N_16837,N_15153,N_15760);
or U16838 (N_16838,N_15199,N_14161);
or U16839 (N_16839,N_15170,N_15147);
xor U16840 (N_16840,N_14163,N_14791);
nand U16841 (N_16841,N_14069,N_14822);
xor U16842 (N_16842,N_15935,N_14770);
and U16843 (N_16843,N_14838,N_14841);
xor U16844 (N_16844,N_14955,N_15719);
or U16845 (N_16845,N_14767,N_14723);
xnor U16846 (N_16846,N_15128,N_15515);
xor U16847 (N_16847,N_15841,N_15142);
nor U16848 (N_16848,N_14574,N_14663);
xor U16849 (N_16849,N_14664,N_15824);
nor U16850 (N_16850,N_14734,N_15696);
nand U16851 (N_16851,N_15857,N_14226);
and U16852 (N_16852,N_15336,N_15071);
nand U16853 (N_16853,N_14868,N_15794);
nor U16854 (N_16854,N_15112,N_15419);
nand U16855 (N_16855,N_14742,N_15440);
nor U16856 (N_16856,N_15715,N_15059);
xor U16857 (N_16857,N_14174,N_14616);
xnor U16858 (N_16858,N_14910,N_14802);
nor U16859 (N_16859,N_14221,N_14063);
nor U16860 (N_16860,N_15397,N_15363);
nand U16861 (N_16861,N_14319,N_14782);
nor U16862 (N_16862,N_14811,N_15778);
and U16863 (N_16863,N_14543,N_15932);
nand U16864 (N_16864,N_15548,N_15471);
nand U16865 (N_16865,N_15217,N_15793);
and U16866 (N_16866,N_15895,N_15600);
nand U16867 (N_16867,N_15161,N_15404);
xnor U16868 (N_16868,N_15790,N_14884);
xnor U16869 (N_16869,N_15910,N_14331);
nand U16870 (N_16870,N_14342,N_15629);
or U16871 (N_16871,N_15823,N_14229);
nor U16872 (N_16872,N_15349,N_14775);
xnor U16873 (N_16873,N_14555,N_14772);
nor U16874 (N_16874,N_14029,N_15870);
nand U16875 (N_16875,N_14401,N_15227);
or U16876 (N_16876,N_15647,N_15695);
and U16877 (N_16877,N_14641,N_15347);
nor U16878 (N_16878,N_14516,N_15060);
and U16879 (N_16879,N_15138,N_14712);
and U16880 (N_16880,N_15020,N_15892);
nand U16881 (N_16881,N_15814,N_15484);
nor U16882 (N_16882,N_14529,N_15930);
or U16883 (N_16883,N_14444,N_14039);
and U16884 (N_16884,N_15458,N_15945);
and U16885 (N_16885,N_14435,N_15083);
nand U16886 (N_16886,N_14123,N_14205);
or U16887 (N_16887,N_15584,N_15742);
nand U16888 (N_16888,N_15408,N_14899);
and U16889 (N_16889,N_14479,N_14114);
and U16890 (N_16890,N_15531,N_14013);
xnor U16891 (N_16891,N_14658,N_15450);
nand U16892 (N_16892,N_14434,N_14852);
or U16893 (N_16893,N_15503,N_14104);
nor U16894 (N_16894,N_15838,N_14588);
or U16895 (N_16895,N_15168,N_15846);
or U16896 (N_16896,N_14170,N_14630);
and U16897 (N_16897,N_15900,N_15623);
xnor U16898 (N_16898,N_14131,N_14437);
and U16899 (N_16899,N_15683,N_15219);
and U16900 (N_16900,N_15157,N_15919);
xor U16901 (N_16901,N_15055,N_15148);
or U16902 (N_16902,N_15852,N_15428);
and U16903 (N_16903,N_14115,N_15399);
nand U16904 (N_16904,N_15420,N_14030);
or U16905 (N_16905,N_14839,N_14470);
or U16906 (N_16906,N_15999,N_15432);
nor U16907 (N_16907,N_15159,N_15708);
xnor U16908 (N_16908,N_14175,N_15054);
xnor U16909 (N_16909,N_15981,N_15195);
xnor U16910 (N_16910,N_14989,N_14509);
and U16911 (N_16911,N_15225,N_15501);
or U16912 (N_16912,N_14295,N_15575);
nand U16913 (N_16913,N_14737,N_15224);
or U16914 (N_16914,N_15830,N_14231);
nand U16915 (N_16915,N_14000,N_15386);
nor U16916 (N_16916,N_14762,N_15756);
and U16917 (N_16917,N_14798,N_15266);
nor U16918 (N_16918,N_15675,N_14845);
xor U16919 (N_16919,N_15084,N_15536);
nand U16920 (N_16920,N_14305,N_15850);
or U16921 (N_16921,N_14405,N_15994);
nor U16922 (N_16922,N_14769,N_14279);
nor U16923 (N_16923,N_14287,N_15017);
and U16924 (N_16924,N_14832,N_15276);
nand U16925 (N_16925,N_15387,N_15260);
xor U16926 (N_16926,N_14784,N_14084);
xnor U16927 (N_16927,N_14729,N_14924);
xor U16928 (N_16928,N_15198,N_15706);
or U16929 (N_16929,N_14058,N_14694);
nor U16930 (N_16930,N_14031,N_14771);
xnor U16931 (N_16931,N_14309,N_14036);
xnor U16932 (N_16932,N_14991,N_15813);
or U16933 (N_16933,N_14524,N_15728);
nand U16934 (N_16934,N_14551,N_14081);
nor U16935 (N_16935,N_14259,N_15005);
xnor U16936 (N_16936,N_14777,N_15750);
and U16937 (N_16937,N_15642,N_15710);
nor U16938 (N_16938,N_15319,N_15523);
nand U16939 (N_16939,N_15507,N_15680);
nor U16940 (N_16940,N_14637,N_14894);
nand U16941 (N_16941,N_14390,N_15682);
xor U16942 (N_16942,N_15878,N_15859);
or U16943 (N_16943,N_14677,N_15714);
nor U16944 (N_16944,N_15211,N_14925);
and U16945 (N_16945,N_14961,N_14684);
xor U16946 (N_16946,N_15724,N_14994);
nand U16947 (N_16947,N_15954,N_15559);
nor U16948 (N_16948,N_14126,N_15427);
xnor U16949 (N_16949,N_14022,N_15308);
nor U16950 (N_16950,N_15786,N_15631);
xor U16951 (N_16951,N_15367,N_14372);
nor U16952 (N_16952,N_15688,N_14391);
and U16953 (N_16953,N_15923,N_15506);
or U16954 (N_16954,N_15681,N_15869);
nand U16955 (N_16955,N_15806,N_15384);
or U16956 (N_16956,N_14612,N_14387);
xor U16957 (N_16957,N_14564,N_14481);
or U16958 (N_16958,N_14847,N_15925);
and U16959 (N_16959,N_14421,N_14833);
and U16960 (N_16960,N_14049,N_14844);
or U16961 (N_16961,N_15014,N_15042);
nand U16962 (N_16962,N_15239,N_15099);
nand U16963 (N_16963,N_14633,N_14399);
and U16964 (N_16964,N_15717,N_15759);
or U16965 (N_16965,N_14474,N_15409);
and U16966 (N_16966,N_14895,N_15228);
and U16967 (N_16967,N_15203,N_14251);
or U16968 (N_16968,N_15356,N_15185);
xnor U16969 (N_16969,N_15886,N_15622);
nand U16970 (N_16970,N_14360,N_14517);
and U16971 (N_16971,N_14640,N_15801);
and U16972 (N_16972,N_15026,N_15589);
nor U16973 (N_16973,N_15573,N_14208);
xor U16974 (N_16974,N_14608,N_14667);
and U16975 (N_16975,N_14823,N_14556);
nor U16976 (N_16976,N_14545,N_15341);
xnor U16977 (N_16977,N_14185,N_14373);
or U16978 (N_16978,N_14012,N_15102);
nand U16979 (N_16979,N_15050,N_15479);
and U16980 (N_16980,N_15836,N_15744);
xor U16981 (N_16981,N_15063,N_14687);
nand U16982 (N_16982,N_14929,N_14348);
nor U16983 (N_16983,N_14795,N_15834);
nor U16984 (N_16984,N_14501,N_15535);
and U16985 (N_16985,N_15477,N_15845);
and U16986 (N_16986,N_14624,N_15057);
and U16987 (N_16987,N_15030,N_14487);
nand U16988 (N_16988,N_15855,N_14647);
and U16989 (N_16989,N_14834,N_15671);
and U16990 (N_16990,N_14411,N_14990);
and U16991 (N_16991,N_15899,N_15670);
nor U16992 (N_16992,N_14679,N_14230);
or U16993 (N_16993,N_15730,N_15885);
nor U16994 (N_16994,N_15433,N_15383);
and U16995 (N_16995,N_15434,N_15898);
or U16996 (N_16996,N_14341,N_15832);
nor U16997 (N_16997,N_14882,N_15378);
nand U16998 (N_16998,N_15873,N_15335);
nor U16999 (N_16999,N_14562,N_14352);
nand U17000 (N_17000,N_14478,N_15130);
nor U17001 (N_17001,N_15897,N_15424);
nand U17002 (N_17002,N_15900,N_14074);
nand U17003 (N_17003,N_14264,N_14612);
and U17004 (N_17004,N_15123,N_14143);
xnor U17005 (N_17005,N_14565,N_14796);
nor U17006 (N_17006,N_14860,N_14631);
xor U17007 (N_17007,N_15423,N_15652);
nor U17008 (N_17008,N_14304,N_14747);
xnor U17009 (N_17009,N_14071,N_14731);
nor U17010 (N_17010,N_14853,N_14552);
nor U17011 (N_17011,N_14042,N_15938);
xor U17012 (N_17012,N_15540,N_14503);
and U17013 (N_17013,N_15939,N_15417);
nor U17014 (N_17014,N_15255,N_14707);
and U17015 (N_17015,N_15380,N_15241);
or U17016 (N_17016,N_15499,N_14701);
and U17017 (N_17017,N_14466,N_15369);
nor U17018 (N_17018,N_15038,N_14572);
nor U17019 (N_17019,N_14445,N_15621);
or U17020 (N_17020,N_14326,N_15865);
nand U17021 (N_17021,N_14308,N_15415);
or U17022 (N_17022,N_15089,N_14289);
or U17023 (N_17023,N_15925,N_14721);
nor U17024 (N_17024,N_14089,N_15337);
xor U17025 (N_17025,N_14945,N_15160);
or U17026 (N_17026,N_14091,N_14808);
nand U17027 (N_17027,N_15811,N_14594);
and U17028 (N_17028,N_14795,N_14024);
and U17029 (N_17029,N_15367,N_14226);
nand U17030 (N_17030,N_15550,N_14534);
nand U17031 (N_17031,N_15638,N_14488);
nand U17032 (N_17032,N_14049,N_15080);
nor U17033 (N_17033,N_14199,N_14080);
xnor U17034 (N_17034,N_14165,N_14096);
and U17035 (N_17035,N_15783,N_14907);
nor U17036 (N_17036,N_14391,N_15296);
nand U17037 (N_17037,N_15762,N_15736);
and U17038 (N_17038,N_14720,N_14730);
xor U17039 (N_17039,N_14653,N_14374);
and U17040 (N_17040,N_15086,N_15628);
nor U17041 (N_17041,N_15406,N_14156);
and U17042 (N_17042,N_14011,N_15159);
xor U17043 (N_17043,N_14043,N_15579);
and U17044 (N_17044,N_14740,N_14282);
nand U17045 (N_17045,N_14124,N_15736);
or U17046 (N_17046,N_15677,N_14967);
and U17047 (N_17047,N_14721,N_15959);
nor U17048 (N_17048,N_14735,N_15645);
and U17049 (N_17049,N_15414,N_14564);
xor U17050 (N_17050,N_15085,N_15702);
and U17051 (N_17051,N_15687,N_15193);
nor U17052 (N_17052,N_14114,N_15858);
nand U17053 (N_17053,N_14563,N_14516);
nor U17054 (N_17054,N_15377,N_14594);
xor U17055 (N_17055,N_15217,N_14158);
or U17056 (N_17056,N_14147,N_15288);
nor U17057 (N_17057,N_14256,N_15649);
nor U17058 (N_17058,N_14712,N_14838);
nand U17059 (N_17059,N_14880,N_14380);
nor U17060 (N_17060,N_15309,N_15587);
and U17061 (N_17061,N_15619,N_15906);
and U17062 (N_17062,N_14363,N_14180);
or U17063 (N_17063,N_14016,N_15059);
or U17064 (N_17064,N_14641,N_15496);
nand U17065 (N_17065,N_14284,N_15064);
nand U17066 (N_17066,N_15933,N_14923);
or U17067 (N_17067,N_14444,N_15851);
and U17068 (N_17068,N_14001,N_14517);
xnor U17069 (N_17069,N_14803,N_14357);
nand U17070 (N_17070,N_14616,N_15139);
and U17071 (N_17071,N_14765,N_15732);
and U17072 (N_17072,N_15495,N_14938);
or U17073 (N_17073,N_15387,N_14506);
or U17074 (N_17074,N_15680,N_14213);
and U17075 (N_17075,N_15333,N_15445);
xnor U17076 (N_17076,N_14391,N_14642);
nand U17077 (N_17077,N_15605,N_14643);
nand U17078 (N_17078,N_14181,N_14581);
nand U17079 (N_17079,N_15637,N_15332);
xnor U17080 (N_17080,N_14455,N_15145);
xnor U17081 (N_17081,N_15408,N_15647);
xnor U17082 (N_17082,N_14315,N_15467);
and U17083 (N_17083,N_14723,N_15871);
or U17084 (N_17084,N_14786,N_15903);
and U17085 (N_17085,N_15868,N_15731);
xnor U17086 (N_17086,N_14445,N_14026);
xnor U17087 (N_17087,N_15235,N_14980);
nand U17088 (N_17088,N_15282,N_14030);
xnor U17089 (N_17089,N_14573,N_14805);
xor U17090 (N_17090,N_15965,N_15674);
or U17091 (N_17091,N_15847,N_14680);
nand U17092 (N_17092,N_14000,N_15927);
xor U17093 (N_17093,N_14097,N_14375);
nand U17094 (N_17094,N_15273,N_14909);
xor U17095 (N_17095,N_15749,N_14203);
nor U17096 (N_17096,N_14977,N_15207);
or U17097 (N_17097,N_15413,N_15766);
xnor U17098 (N_17098,N_14211,N_14835);
nand U17099 (N_17099,N_15893,N_15181);
xor U17100 (N_17100,N_14787,N_14695);
and U17101 (N_17101,N_15008,N_14316);
xor U17102 (N_17102,N_14101,N_14064);
or U17103 (N_17103,N_15698,N_15966);
xnor U17104 (N_17104,N_14834,N_15901);
nand U17105 (N_17105,N_15308,N_15980);
and U17106 (N_17106,N_14578,N_14742);
nand U17107 (N_17107,N_14499,N_15073);
nand U17108 (N_17108,N_15180,N_15573);
and U17109 (N_17109,N_14738,N_15505);
and U17110 (N_17110,N_15541,N_14857);
nor U17111 (N_17111,N_15584,N_14223);
nor U17112 (N_17112,N_15857,N_15820);
or U17113 (N_17113,N_15280,N_15318);
xor U17114 (N_17114,N_15695,N_15023);
nand U17115 (N_17115,N_15176,N_15980);
or U17116 (N_17116,N_15721,N_15520);
or U17117 (N_17117,N_15473,N_14683);
nand U17118 (N_17118,N_15747,N_15842);
nor U17119 (N_17119,N_14642,N_14847);
nand U17120 (N_17120,N_15004,N_15773);
xor U17121 (N_17121,N_15978,N_14628);
xor U17122 (N_17122,N_15931,N_15794);
xor U17123 (N_17123,N_15308,N_15824);
and U17124 (N_17124,N_15810,N_14407);
nand U17125 (N_17125,N_15244,N_14543);
xor U17126 (N_17126,N_15306,N_15549);
and U17127 (N_17127,N_14106,N_15058);
or U17128 (N_17128,N_15342,N_14300);
nor U17129 (N_17129,N_15077,N_14339);
xnor U17130 (N_17130,N_15070,N_15457);
nor U17131 (N_17131,N_15033,N_14152);
nand U17132 (N_17132,N_15509,N_15301);
nand U17133 (N_17133,N_15994,N_15307);
xnor U17134 (N_17134,N_14929,N_15767);
nand U17135 (N_17135,N_15236,N_14467);
xor U17136 (N_17136,N_14375,N_14043);
and U17137 (N_17137,N_14011,N_15745);
or U17138 (N_17138,N_14754,N_15461);
and U17139 (N_17139,N_14015,N_15119);
or U17140 (N_17140,N_15066,N_14597);
or U17141 (N_17141,N_15746,N_15902);
and U17142 (N_17142,N_14090,N_15706);
or U17143 (N_17143,N_15340,N_15091);
xor U17144 (N_17144,N_15096,N_14418);
nand U17145 (N_17145,N_14630,N_15605);
nor U17146 (N_17146,N_15942,N_14485);
nor U17147 (N_17147,N_15286,N_15684);
nand U17148 (N_17148,N_15794,N_15855);
nand U17149 (N_17149,N_14958,N_14382);
nand U17150 (N_17150,N_14064,N_15816);
nor U17151 (N_17151,N_15257,N_15213);
and U17152 (N_17152,N_15482,N_14186);
nand U17153 (N_17153,N_14329,N_14641);
nand U17154 (N_17154,N_14488,N_14811);
xnor U17155 (N_17155,N_15906,N_15806);
nor U17156 (N_17156,N_15171,N_15038);
and U17157 (N_17157,N_15166,N_15712);
nand U17158 (N_17158,N_15769,N_14421);
or U17159 (N_17159,N_14096,N_15261);
and U17160 (N_17160,N_15682,N_14848);
or U17161 (N_17161,N_15679,N_15932);
or U17162 (N_17162,N_14992,N_15213);
and U17163 (N_17163,N_14849,N_14646);
nor U17164 (N_17164,N_15377,N_15649);
nand U17165 (N_17165,N_15950,N_15108);
and U17166 (N_17166,N_14665,N_15301);
or U17167 (N_17167,N_14985,N_14486);
nor U17168 (N_17168,N_14956,N_14354);
and U17169 (N_17169,N_14049,N_15529);
nand U17170 (N_17170,N_15980,N_14173);
or U17171 (N_17171,N_15067,N_15417);
or U17172 (N_17172,N_15937,N_14147);
nand U17173 (N_17173,N_14244,N_15390);
or U17174 (N_17174,N_14712,N_14539);
and U17175 (N_17175,N_14211,N_15259);
nor U17176 (N_17176,N_14812,N_15122);
nand U17177 (N_17177,N_15318,N_15879);
or U17178 (N_17178,N_15282,N_14233);
or U17179 (N_17179,N_15331,N_14106);
nor U17180 (N_17180,N_14965,N_14541);
xor U17181 (N_17181,N_15246,N_14620);
nand U17182 (N_17182,N_14406,N_15144);
nor U17183 (N_17183,N_14514,N_15272);
nor U17184 (N_17184,N_15648,N_15174);
and U17185 (N_17185,N_15750,N_14720);
or U17186 (N_17186,N_15214,N_15782);
nor U17187 (N_17187,N_15432,N_15033);
nand U17188 (N_17188,N_14682,N_14582);
xnor U17189 (N_17189,N_15898,N_15062);
nand U17190 (N_17190,N_14427,N_15755);
nor U17191 (N_17191,N_14333,N_14788);
and U17192 (N_17192,N_15152,N_15081);
or U17193 (N_17193,N_14558,N_15094);
nand U17194 (N_17194,N_14171,N_15859);
or U17195 (N_17195,N_14330,N_14032);
nor U17196 (N_17196,N_14067,N_14569);
nor U17197 (N_17197,N_15476,N_14645);
or U17198 (N_17198,N_15282,N_15360);
and U17199 (N_17199,N_14224,N_15810);
and U17200 (N_17200,N_14725,N_14039);
xnor U17201 (N_17201,N_15449,N_14377);
xor U17202 (N_17202,N_15510,N_15243);
nor U17203 (N_17203,N_14351,N_14985);
nor U17204 (N_17204,N_15508,N_14956);
nor U17205 (N_17205,N_15572,N_14025);
or U17206 (N_17206,N_15856,N_14666);
nand U17207 (N_17207,N_15130,N_14725);
or U17208 (N_17208,N_15407,N_14429);
nand U17209 (N_17209,N_15387,N_15143);
nor U17210 (N_17210,N_14407,N_15681);
and U17211 (N_17211,N_14811,N_15307);
nand U17212 (N_17212,N_15566,N_15192);
nor U17213 (N_17213,N_14002,N_15431);
or U17214 (N_17214,N_15634,N_15932);
nor U17215 (N_17215,N_15452,N_14650);
and U17216 (N_17216,N_14278,N_14589);
xor U17217 (N_17217,N_15132,N_14384);
nand U17218 (N_17218,N_15059,N_15267);
nand U17219 (N_17219,N_15565,N_14927);
or U17220 (N_17220,N_15133,N_14128);
xor U17221 (N_17221,N_14856,N_14158);
xnor U17222 (N_17222,N_15857,N_14815);
xor U17223 (N_17223,N_14970,N_14060);
and U17224 (N_17224,N_15755,N_14402);
nand U17225 (N_17225,N_15032,N_15451);
and U17226 (N_17226,N_14330,N_14590);
or U17227 (N_17227,N_14196,N_15539);
or U17228 (N_17228,N_15713,N_14240);
or U17229 (N_17229,N_15379,N_14468);
or U17230 (N_17230,N_15558,N_15952);
nor U17231 (N_17231,N_14107,N_15480);
and U17232 (N_17232,N_15030,N_15143);
nand U17233 (N_17233,N_15112,N_14702);
nor U17234 (N_17234,N_15179,N_15741);
or U17235 (N_17235,N_14486,N_14635);
and U17236 (N_17236,N_15444,N_14372);
or U17237 (N_17237,N_14868,N_15326);
xnor U17238 (N_17238,N_14179,N_15909);
xor U17239 (N_17239,N_14325,N_15151);
nand U17240 (N_17240,N_15106,N_15847);
xnor U17241 (N_17241,N_14343,N_14113);
and U17242 (N_17242,N_15641,N_15761);
or U17243 (N_17243,N_14726,N_14991);
nand U17244 (N_17244,N_14213,N_15445);
or U17245 (N_17245,N_14594,N_14328);
or U17246 (N_17246,N_15040,N_14098);
xnor U17247 (N_17247,N_15384,N_14527);
nor U17248 (N_17248,N_15342,N_14615);
xor U17249 (N_17249,N_14808,N_14277);
xor U17250 (N_17250,N_14163,N_14323);
xor U17251 (N_17251,N_15577,N_14886);
nand U17252 (N_17252,N_14935,N_15698);
xnor U17253 (N_17253,N_14766,N_15449);
and U17254 (N_17254,N_14087,N_14395);
nor U17255 (N_17255,N_15504,N_15659);
nor U17256 (N_17256,N_14593,N_14440);
xor U17257 (N_17257,N_15540,N_15856);
xor U17258 (N_17258,N_15853,N_15123);
and U17259 (N_17259,N_15892,N_14243);
nor U17260 (N_17260,N_15041,N_14110);
nor U17261 (N_17261,N_15483,N_14351);
nor U17262 (N_17262,N_14162,N_14474);
xor U17263 (N_17263,N_15315,N_14832);
and U17264 (N_17264,N_15636,N_15455);
xnor U17265 (N_17265,N_14637,N_15087);
or U17266 (N_17266,N_15344,N_14126);
nor U17267 (N_17267,N_15796,N_14505);
nor U17268 (N_17268,N_14517,N_15921);
nand U17269 (N_17269,N_14768,N_15859);
nor U17270 (N_17270,N_15824,N_15005);
xnor U17271 (N_17271,N_15356,N_14063);
xnor U17272 (N_17272,N_14232,N_14386);
and U17273 (N_17273,N_14983,N_15785);
and U17274 (N_17274,N_15389,N_14253);
and U17275 (N_17275,N_15980,N_15291);
nand U17276 (N_17276,N_15611,N_14220);
nand U17277 (N_17277,N_15907,N_14915);
and U17278 (N_17278,N_14376,N_15332);
nor U17279 (N_17279,N_15619,N_14661);
xor U17280 (N_17280,N_14017,N_15427);
xor U17281 (N_17281,N_14252,N_15351);
or U17282 (N_17282,N_15603,N_15985);
nor U17283 (N_17283,N_15788,N_15456);
and U17284 (N_17284,N_15916,N_14081);
nor U17285 (N_17285,N_15249,N_15192);
xor U17286 (N_17286,N_15496,N_15350);
and U17287 (N_17287,N_15977,N_14222);
nor U17288 (N_17288,N_14520,N_14323);
nor U17289 (N_17289,N_15275,N_14961);
and U17290 (N_17290,N_15889,N_14280);
xnor U17291 (N_17291,N_15637,N_14130);
nor U17292 (N_17292,N_15177,N_14920);
nand U17293 (N_17293,N_15120,N_14193);
xnor U17294 (N_17294,N_14560,N_15956);
nor U17295 (N_17295,N_14113,N_14481);
nor U17296 (N_17296,N_15866,N_15275);
nor U17297 (N_17297,N_15964,N_14058);
nand U17298 (N_17298,N_14630,N_15147);
nand U17299 (N_17299,N_14084,N_14484);
nand U17300 (N_17300,N_15193,N_15369);
nand U17301 (N_17301,N_15455,N_14237);
nand U17302 (N_17302,N_15130,N_15311);
nor U17303 (N_17303,N_15054,N_15228);
nor U17304 (N_17304,N_14182,N_15166);
or U17305 (N_17305,N_14498,N_14334);
nand U17306 (N_17306,N_14672,N_14499);
nor U17307 (N_17307,N_14888,N_15660);
and U17308 (N_17308,N_14197,N_14883);
nand U17309 (N_17309,N_14220,N_14802);
nand U17310 (N_17310,N_14289,N_15541);
nor U17311 (N_17311,N_15759,N_15818);
and U17312 (N_17312,N_15735,N_15190);
xor U17313 (N_17313,N_15362,N_15805);
or U17314 (N_17314,N_14820,N_15192);
and U17315 (N_17315,N_14642,N_15889);
nor U17316 (N_17316,N_15643,N_15317);
nor U17317 (N_17317,N_15413,N_14824);
or U17318 (N_17318,N_14823,N_15430);
or U17319 (N_17319,N_15094,N_15881);
nor U17320 (N_17320,N_14100,N_15284);
or U17321 (N_17321,N_15998,N_14236);
nand U17322 (N_17322,N_14471,N_15844);
xnor U17323 (N_17323,N_15657,N_14203);
xor U17324 (N_17324,N_15534,N_15144);
xor U17325 (N_17325,N_14196,N_14568);
xor U17326 (N_17326,N_15012,N_14740);
or U17327 (N_17327,N_15423,N_14771);
xnor U17328 (N_17328,N_15486,N_14106);
nand U17329 (N_17329,N_14772,N_14778);
or U17330 (N_17330,N_14294,N_14817);
nor U17331 (N_17331,N_14262,N_14121);
or U17332 (N_17332,N_15760,N_15323);
or U17333 (N_17333,N_15111,N_15583);
nand U17334 (N_17334,N_14501,N_14696);
nand U17335 (N_17335,N_14273,N_14279);
or U17336 (N_17336,N_15612,N_14698);
nor U17337 (N_17337,N_14219,N_15161);
xor U17338 (N_17338,N_15476,N_14944);
or U17339 (N_17339,N_14251,N_15019);
xnor U17340 (N_17340,N_14515,N_14381);
and U17341 (N_17341,N_14824,N_14441);
nand U17342 (N_17342,N_14644,N_15116);
nand U17343 (N_17343,N_14803,N_14702);
nand U17344 (N_17344,N_15764,N_15185);
nand U17345 (N_17345,N_14702,N_14386);
nand U17346 (N_17346,N_15790,N_14055);
or U17347 (N_17347,N_14839,N_14576);
and U17348 (N_17348,N_15419,N_14137);
nand U17349 (N_17349,N_15811,N_14687);
xnor U17350 (N_17350,N_14873,N_14108);
xor U17351 (N_17351,N_15321,N_15510);
xnor U17352 (N_17352,N_14130,N_14421);
xor U17353 (N_17353,N_15290,N_14557);
xnor U17354 (N_17354,N_15918,N_14173);
nand U17355 (N_17355,N_15803,N_15107);
nor U17356 (N_17356,N_15158,N_14031);
nand U17357 (N_17357,N_14365,N_14970);
and U17358 (N_17358,N_15104,N_14085);
nand U17359 (N_17359,N_14842,N_14609);
and U17360 (N_17360,N_15785,N_15256);
nor U17361 (N_17361,N_14908,N_15771);
xnor U17362 (N_17362,N_14086,N_15629);
nand U17363 (N_17363,N_15571,N_14502);
xnor U17364 (N_17364,N_14569,N_15485);
and U17365 (N_17365,N_15182,N_14118);
and U17366 (N_17366,N_15622,N_14842);
and U17367 (N_17367,N_14815,N_15107);
nor U17368 (N_17368,N_14553,N_15166);
nor U17369 (N_17369,N_14232,N_14553);
or U17370 (N_17370,N_14170,N_15222);
nand U17371 (N_17371,N_15607,N_14696);
nor U17372 (N_17372,N_15054,N_15886);
nor U17373 (N_17373,N_15654,N_14893);
and U17374 (N_17374,N_15256,N_14712);
nand U17375 (N_17375,N_15666,N_15163);
and U17376 (N_17376,N_14542,N_15916);
xnor U17377 (N_17377,N_14894,N_14061);
or U17378 (N_17378,N_15980,N_14631);
nand U17379 (N_17379,N_15720,N_15429);
or U17380 (N_17380,N_15109,N_15329);
nand U17381 (N_17381,N_14558,N_14200);
nor U17382 (N_17382,N_14464,N_14888);
and U17383 (N_17383,N_14023,N_14211);
nor U17384 (N_17384,N_15139,N_14969);
xnor U17385 (N_17385,N_14926,N_14141);
nor U17386 (N_17386,N_14985,N_14689);
nor U17387 (N_17387,N_15782,N_15572);
nor U17388 (N_17388,N_14176,N_14190);
xor U17389 (N_17389,N_15222,N_14015);
and U17390 (N_17390,N_14016,N_15209);
nand U17391 (N_17391,N_14796,N_14293);
and U17392 (N_17392,N_15126,N_14076);
and U17393 (N_17393,N_15787,N_14462);
nor U17394 (N_17394,N_14456,N_15078);
nor U17395 (N_17395,N_14201,N_15544);
nand U17396 (N_17396,N_14475,N_15462);
and U17397 (N_17397,N_14440,N_15611);
or U17398 (N_17398,N_14884,N_15696);
nor U17399 (N_17399,N_14811,N_14395);
nand U17400 (N_17400,N_15035,N_14054);
or U17401 (N_17401,N_15867,N_14050);
or U17402 (N_17402,N_14714,N_14882);
or U17403 (N_17403,N_15150,N_14212);
xnor U17404 (N_17404,N_14851,N_15997);
or U17405 (N_17405,N_15703,N_14580);
nor U17406 (N_17406,N_15620,N_14491);
nor U17407 (N_17407,N_15228,N_14385);
xor U17408 (N_17408,N_14417,N_15199);
xor U17409 (N_17409,N_14375,N_14315);
and U17410 (N_17410,N_14216,N_15175);
or U17411 (N_17411,N_14584,N_15947);
xnor U17412 (N_17412,N_14114,N_15622);
xor U17413 (N_17413,N_14117,N_15657);
and U17414 (N_17414,N_15623,N_14692);
nand U17415 (N_17415,N_14256,N_14594);
nand U17416 (N_17416,N_15314,N_14367);
nor U17417 (N_17417,N_14765,N_14369);
or U17418 (N_17418,N_15320,N_14194);
nand U17419 (N_17419,N_14256,N_14413);
nor U17420 (N_17420,N_15720,N_15602);
and U17421 (N_17421,N_15454,N_14434);
nand U17422 (N_17422,N_15967,N_15044);
nand U17423 (N_17423,N_14268,N_14057);
nor U17424 (N_17424,N_14700,N_14415);
nand U17425 (N_17425,N_14002,N_14395);
nand U17426 (N_17426,N_14114,N_15080);
nor U17427 (N_17427,N_14433,N_14509);
or U17428 (N_17428,N_14322,N_15990);
nor U17429 (N_17429,N_15677,N_15139);
nor U17430 (N_17430,N_14482,N_15770);
nand U17431 (N_17431,N_14734,N_14834);
xnor U17432 (N_17432,N_15265,N_14028);
and U17433 (N_17433,N_15288,N_15534);
nor U17434 (N_17434,N_14564,N_14081);
or U17435 (N_17435,N_14597,N_15551);
and U17436 (N_17436,N_15123,N_14180);
nor U17437 (N_17437,N_15640,N_15897);
or U17438 (N_17438,N_14389,N_14163);
nor U17439 (N_17439,N_14492,N_14112);
xor U17440 (N_17440,N_15435,N_14588);
nor U17441 (N_17441,N_14931,N_15478);
nand U17442 (N_17442,N_14981,N_15358);
nor U17443 (N_17443,N_14609,N_14321);
xnor U17444 (N_17444,N_14518,N_14588);
or U17445 (N_17445,N_15562,N_14873);
xnor U17446 (N_17446,N_15514,N_14138);
xor U17447 (N_17447,N_15216,N_14180);
or U17448 (N_17448,N_15329,N_15606);
nand U17449 (N_17449,N_14339,N_15376);
nor U17450 (N_17450,N_14381,N_14304);
nand U17451 (N_17451,N_14344,N_14357);
or U17452 (N_17452,N_14237,N_14940);
or U17453 (N_17453,N_15488,N_15710);
nand U17454 (N_17454,N_14061,N_14451);
and U17455 (N_17455,N_15071,N_14218);
or U17456 (N_17456,N_14036,N_15023);
nand U17457 (N_17457,N_15669,N_15191);
or U17458 (N_17458,N_14807,N_14790);
nor U17459 (N_17459,N_14198,N_15740);
and U17460 (N_17460,N_14889,N_14794);
xor U17461 (N_17461,N_15282,N_14746);
nand U17462 (N_17462,N_14122,N_14812);
and U17463 (N_17463,N_15065,N_15234);
nand U17464 (N_17464,N_15420,N_15826);
or U17465 (N_17465,N_14799,N_14199);
or U17466 (N_17466,N_15323,N_15431);
nand U17467 (N_17467,N_15007,N_15112);
xor U17468 (N_17468,N_14938,N_14056);
or U17469 (N_17469,N_15272,N_15104);
nor U17470 (N_17470,N_14775,N_15511);
nor U17471 (N_17471,N_14631,N_14858);
and U17472 (N_17472,N_14787,N_15076);
or U17473 (N_17473,N_14526,N_15465);
and U17474 (N_17474,N_14213,N_14889);
and U17475 (N_17475,N_14770,N_15035);
or U17476 (N_17476,N_15071,N_15753);
xor U17477 (N_17477,N_15478,N_14959);
xnor U17478 (N_17478,N_14631,N_15853);
nor U17479 (N_17479,N_15225,N_14807);
xor U17480 (N_17480,N_14648,N_14494);
and U17481 (N_17481,N_14361,N_14936);
xnor U17482 (N_17482,N_14135,N_15863);
and U17483 (N_17483,N_15052,N_14965);
and U17484 (N_17484,N_15885,N_15480);
nor U17485 (N_17485,N_14705,N_15399);
xnor U17486 (N_17486,N_15057,N_14908);
or U17487 (N_17487,N_14028,N_14645);
nand U17488 (N_17488,N_14839,N_15847);
and U17489 (N_17489,N_15903,N_15231);
and U17490 (N_17490,N_14979,N_15851);
or U17491 (N_17491,N_14210,N_14664);
and U17492 (N_17492,N_15849,N_15918);
nand U17493 (N_17493,N_15501,N_15288);
xor U17494 (N_17494,N_15719,N_14539);
xor U17495 (N_17495,N_15567,N_15174);
nor U17496 (N_17496,N_15007,N_14107);
and U17497 (N_17497,N_14349,N_14035);
or U17498 (N_17498,N_14806,N_15650);
and U17499 (N_17499,N_14201,N_14027);
or U17500 (N_17500,N_15005,N_15070);
nand U17501 (N_17501,N_14037,N_14756);
nor U17502 (N_17502,N_15294,N_15885);
or U17503 (N_17503,N_15203,N_14320);
nor U17504 (N_17504,N_14670,N_14283);
and U17505 (N_17505,N_15823,N_14352);
xnor U17506 (N_17506,N_14263,N_15924);
xor U17507 (N_17507,N_15757,N_14631);
nand U17508 (N_17508,N_15398,N_14706);
or U17509 (N_17509,N_15101,N_15401);
nand U17510 (N_17510,N_15461,N_14866);
or U17511 (N_17511,N_14955,N_14128);
or U17512 (N_17512,N_15201,N_14392);
and U17513 (N_17513,N_15489,N_14526);
xnor U17514 (N_17514,N_15648,N_14655);
nand U17515 (N_17515,N_15863,N_15402);
nand U17516 (N_17516,N_14495,N_14710);
xnor U17517 (N_17517,N_14205,N_15848);
nand U17518 (N_17518,N_15998,N_15335);
xor U17519 (N_17519,N_15122,N_14277);
or U17520 (N_17520,N_15675,N_15091);
and U17521 (N_17521,N_15137,N_14706);
nor U17522 (N_17522,N_15088,N_15025);
nor U17523 (N_17523,N_15580,N_15604);
nor U17524 (N_17524,N_15101,N_15253);
or U17525 (N_17525,N_14335,N_15594);
nand U17526 (N_17526,N_15764,N_15098);
or U17527 (N_17527,N_14958,N_14876);
xnor U17528 (N_17528,N_14517,N_14384);
or U17529 (N_17529,N_14622,N_14162);
nor U17530 (N_17530,N_15381,N_14090);
nor U17531 (N_17531,N_14347,N_15418);
or U17532 (N_17532,N_15793,N_15801);
nand U17533 (N_17533,N_15851,N_14722);
nand U17534 (N_17534,N_15898,N_14898);
and U17535 (N_17535,N_14961,N_15444);
xnor U17536 (N_17536,N_15768,N_14122);
nand U17537 (N_17537,N_14932,N_15823);
or U17538 (N_17538,N_15738,N_14557);
xor U17539 (N_17539,N_14612,N_15978);
nand U17540 (N_17540,N_15246,N_14696);
xnor U17541 (N_17541,N_15938,N_14374);
nand U17542 (N_17542,N_15933,N_15130);
and U17543 (N_17543,N_14635,N_15391);
or U17544 (N_17544,N_14032,N_14044);
and U17545 (N_17545,N_15334,N_14115);
and U17546 (N_17546,N_15712,N_15482);
or U17547 (N_17547,N_15475,N_15982);
xnor U17548 (N_17548,N_15627,N_15951);
nor U17549 (N_17549,N_14263,N_14568);
nand U17550 (N_17550,N_14907,N_14070);
or U17551 (N_17551,N_15619,N_15671);
or U17552 (N_17552,N_15689,N_14955);
nor U17553 (N_17553,N_14114,N_15539);
or U17554 (N_17554,N_15096,N_14571);
nor U17555 (N_17555,N_15928,N_14579);
or U17556 (N_17556,N_15076,N_15901);
xnor U17557 (N_17557,N_14163,N_15912);
and U17558 (N_17558,N_15231,N_15434);
nor U17559 (N_17559,N_14219,N_14064);
nor U17560 (N_17560,N_15831,N_14978);
xor U17561 (N_17561,N_15532,N_14906);
nand U17562 (N_17562,N_15383,N_15547);
or U17563 (N_17563,N_15039,N_14418);
and U17564 (N_17564,N_15476,N_15297);
nor U17565 (N_17565,N_14209,N_15956);
xor U17566 (N_17566,N_15318,N_14731);
or U17567 (N_17567,N_15559,N_15457);
nor U17568 (N_17568,N_15292,N_15638);
or U17569 (N_17569,N_14733,N_14157);
xnor U17570 (N_17570,N_14432,N_15981);
or U17571 (N_17571,N_15110,N_14122);
or U17572 (N_17572,N_15478,N_15133);
nor U17573 (N_17573,N_15459,N_15482);
and U17574 (N_17574,N_14359,N_14092);
or U17575 (N_17575,N_15116,N_15966);
nor U17576 (N_17576,N_14542,N_14360);
or U17577 (N_17577,N_15403,N_14496);
or U17578 (N_17578,N_15328,N_14305);
and U17579 (N_17579,N_15330,N_15320);
nand U17580 (N_17580,N_15004,N_15317);
and U17581 (N_17581,N_14683,N_14474);
or U17582 (N_17582,N_14819,N_15282);
nor U17583 (N_17583,N_14558,N_14559);
and U17584 (N_17584,N_15454,N_14994);
nand U17585 (N_17585,N_15432,N_14296);
nor U17586 (N_17586,N_14330,N_15470);
nand U17587 (N_17587,N_15343,N_14109);
and U17588 (N_17588,N_15281,N_15967);
nor U17589 (N_17589,N_14060,N_15509);
nand U17590 (N_17590,N_15361,N_15336);
nor U17591 (N_17591,N_15055,N_15631);
or U17592 (N_17592,N_15007,N_15818);
nor U17593 (N_17593,N_15413,N_15274);
nor U17594 (N_17594,N_15824,N_14531);
nor U17595 (N_17595,N_15893,N_14907);
or U17596 (N_17596,N_15862,N_15284);
nor U17597 (N_17597,N_15124,N_14526);
and U17598 (N_17598,N_15553,N_15591);
or U17599 (N_17599,N_14638,N_15359);
or U17600 (N_17600,N_14644,N_14156);
nand U17601 (N_17601,N_15348,N_15403);
nor U17602 (N_17602,N_15209,N_15654);
xor U17603 (N_17603,N_14927,N_15688);
nand U17604 (N_17604,N_14109,N_15452);
xnor U17605 (N_17605,N_15273,N_15537);
nand U17606 (N_17606,N_15203,N_14257);
and U17607 (N_17607,N_15770,N_14961);
and U17608 (N_17608,N_15563,N_14434);
and U17609 (N_17609,N_15151,N_14589);
and U17610 (N_17610,N_14346,N_15557);
xnor U17611 (N_17611,N_15624,N_14840);
nor U17612 (N_17612,N_15670,N_15160);
and U17613 (N_17613,N_15305,N_15990);
nand U17614 (N_17614,N_15880,N_14164);
nor U17615 (N_17615,N_15474,N_15084);
xnor U17616 (N_17616,N_15915,N_14335);
or U17617 (N_17617,N_14333,N_14547);
or U17618 (N_17618,N_15051,N_15852);
or U17619 (N_17619,N_15927,N_15595);
nand U17620 (N_17620,N_15639,N_14057);
and U17621 (N_17621,N_15114,N_15603);
nor U17622 (N_17622,N_15697,N_14765);
and U17623 (N_17623,N_14822,N_15318);
or U17624 (N_17624,N_15523,N_15796);
and U17625 (N_17625,N_14305,N_14544);
nand U17626 (N_17626,N_14760,N_15286);
or U17627 (N_17627,N_14277,N_15333);
and U17628 (N_17628,N_15044,N_14798);
nor U17629 (N_17629,N_15981,N_15295);
nand U17630 (N_17630,N_14145,N_15953);
nand U17631 (N_17631,N_15610,N_15966);
or U17632 (N_17632,N_15288,N_15465);
xor U17633 (N_17633,N_14997,N_14882);
nand U17634 (N_17634,N_15496,N_14706);
and U17635 (N_17635,N_14855,N_14482);
nand U17636 (N_17636,N_15281,N_14402);
xor U17637 (N_17637,N_15118,N_14747);
or U17638 (N_17638,N_15844,N_14592);
and U17639 (N_17639,N_14887,N_14596);
nand U17640 (N_17640,N_15300,N_15227);
xnor U17641 (N_17641,N_15447,N_14245);
nand U17642 (N_17642,N_14866,N_14379);
nor U17643 (N_17643,N_15544,N_15620);
nand U17644 (N_17644,N_14053,N_15999);
nor U17645 (N_17645,N_14175,N_15581);
nand U17646 (N_17646,N_15679,N_15258);
or U17647 (N_17647,N_15962,N_14036);
and U17648 (N_17648,N_14689,N_14318);
xnor U17649 (N_17649,N_14899,N_15751);
xor U17650 (N_17650,N_14687,N_14902);
or U17651 (N_17651,N_14826,N_14086);
or U17652 (N_17652,N_15193,N_15168);
nor U17653 (N_17653,N_15373,N_14333);
nand U17654 (N_17654,N_14043,N_15757);
nor U17655 (N_17655,N_15981,N_14160);
xor U17656 (N_17656,N_14649,N_15852);
or U17657 (N_17657,N_15556,N_15801);
and U17658 (N_17658,N_15411,N_14724);
xor U17659 (N_17659,N_14037,N_14593);
nand U17660 (N_17660,N_14673,N_15905);
and U17661 (N_17661,N_14318,N_14119);
nand U17662 (N_17662,N_15429,N_14686);
nand U17663 (N_17663,N_14960,N_14216);
xnor U17664 (N_17664,N_15142,N_14367);
nor U17665 (N_17665,N_14233,N_14867);
nor U17666 (N_17666,N_15390,N_15166);
xor U17667 (N_17667,N_15115,N_14613);
nor U17668 (N_17668,N_14805,N_14765);
and U17669 (N_17669,N_15300,N_14255);
nor U17670 (N_17670,N_14381,N_15488);
or U17671 (N_17671,N_14355,N_14149);
nor U17672 (N_17672,N_14536,N_14596);
xor U17673 (N_17673,N_15961,N_15442);
xor U17674 (N_17674,N_14318,N_15103);
and U17675 (N_17675,N_15537,N_15219);
or U17676 (N_17676,N_14399,N_14360);
and U17677 (N_17677,N_14582,N_15665);
nor U17678 (N_17678,N_14726,N_14987);
xor U17679 (N_17679,N_14202,N_14404);
xor U17680 (N_17680,N_14269,N_14629);
nand U17681 (N_17681,N_15841,N_14041);
and U17682 (N_17682,N_15427,N_15541);
nor U17683 (N_17683,N_15617,N_15218);
nand U17684 (N_17684,N_14435,N_14665);
or U17685 (N_17685,N_15561,N_15419);
xor U17686 (N_17686,N_15634,N_15309);
xnor U17687 (N_17687,N_15890,N_14570);
nor U17688 (N_17688,N_14109,N_15655);
and U17689 (N_17689,N_15037,N_14307);
and U17690 (N_17690,N_14075,N_14893);
nor U17691 (N_17691,N_14748,N_14145);
nand U17692 (N_17692,N_14019,N_14469);
xor U17693 (N_17693,N_14229,N_15639);
or U17694 (N_17694,N_15077,N_14711);
xor U17695 (N_17695,N_15157,N_15411);
nand U17696 (N_17696,N_15060,N_15109);
nor U17697 (N_17697,N_15650,N_15210);
nand U17698 (N_17698,N_15338,N_15051);
and U17699 (N_17699,N_14194,N_15525);
xor U17700 (N_17700,N_14552,N_15165);
or U17701 (N_17701,N_15980,N_14084);
or U17702 (N_17702,N_15683,N_14173);
and U17703 (N_17703,N_14667,N_15233);
xor U17704 (N_17704,N_15736,N_15413);
xor U17705 (N_17705,N_14858,N_15561);
xor U17706 (N_17706,N_14502,N_14984);
and U17707 (N_17707,N_15830,N_14033);
nand U17708 (N_17708,N_14151,N_14843);
nand U17709 (N_17709,N_14992,N_15002);
or U17710 (N_17710,N_14070,N_15363);
nor U17711 (N_17711,N_15467,N_15372);
nand U17712 (N_17712,N_15797,N_14356);
nand U17713 (N_17713,N_15924,N_14259);
nand U17714 (N_17714,N_15608,N_14096);
or U17715 (N_17715,N_14082,N_14044);
nand U17716 (N_17716,N_14178,N_15006);
nand U17717 (N_17717,N_14976,N_15892);
nand U17718 (N_17718,N_15126,N_14641);
nand U17719 (N_17719,N_15576,N_15138);
and U17720 (N_17720,N_15605,N_14145);
and U17721 (N_17721,N_14070,N_15234);
nor U17722 (N_17722,N_14262,N_14120);
nand U17723 (N_17723,N_15429,N_14646);
or U17724 (N_17724,N_14532,N_15917);
and U17725 (N_17725,N_14685,N_15943);
or U17726 (N_17726,N_14593,N_14335);
and U17727 (N_17727,N_15952,N_14601);
xnor U17728 (N_17728,N_14203,N_15816);
and U17729 (N_17729,N_15615,N_15157);
xor U17730 (N_17730,N_15541,N_14996);
nand U17731 (N_17731,N_15605,N_14882);
nand U17732 (N_17732,N_14242,N_15584);
and U17733 (N_17733,N_14201,N_14206);
nor U17734 (N_17734,N_14999,N_14733);
nand U17735 (N_17735,N_14295,N_15630);
and U17736 (N_17736,N_14208,N_15098);
xor U17737 (N_17737,N_15728,N_15882);
nand U17738 (N_17738,N_15273,N_15202);
nor U17739 (N_17739,N_15849,N_14010);
nor U17740 (N_17740,N_14346,N_14942);
nor U17741 (N_17741,N_14341,N_14478);
and U17742 (N_17742,N_15257,N_15510);
xnor U17743 (N_17743,N_15978,N_14132);
nor U17744 (N_17744,N_15284,N_14160);
xnor U17745 (N_17745,N_15182,N_14096);
xor U17746 (N_17746,N_15433,N_15586);
nand U17747 (N_17747,N_15275,N_15597);
or U17748 (N_17748,N_15776,N_14889);
nor U17749 (N_17749,N_15956,N_15428);
xnor U17750 (N_17750,N_14298,N_15424);
nand U17751 (N_17751,N_15816,N_14456);
xor U17752 (N_17752,N_15537,N_14602);
nand U17753 (N_17753,N_15385,N_14888);
nor U17754 (N_17754,N_14621,N_15964);
and U17755 (N_17755,N_15093,N_14514);
or U17756 (N_17756,N_15238,N_15547);
xor U17757 (N_17757,N_14689,N_14740);
or U17758 (N_17758,N_15193,N_14360);
or U17759 (N_17759,N_14145,N_15702);
nor U17760 (N_17760,N_14811,N_14046);
and U17761 (N_17761,N_15403,N_15143);
xor U17762 (N_17762,N_15559,N_14542);
and U17763 (N_17763,N_15715,N_15534);
xnor U17764 (N_17764,N_15567,N_15731);
xnor U17765 (N_17765,N_14925,N_15634);
and U17766 (N_17766,N_15007,N_15809);
nand U17767 (N_17767,N_15183,N_14008);
nor U17768 (N_17768,N_15684,N_15848);
nor U17769 (N_17769,N_15544,N_14838);
xor U17770 (N_17770,N_14218,N_14047);
xor U17771 (N_17771,N_15732,N_14464);
nor U17772 (N_17772,N_14938,N_14791);
and U17773 (N_17773,N_14885,N_15942);
and U17774 (N_17774,N_15363,N_14407);
nand U17775 (N_17775,N_14641,N_15544);
or U17776 (N_17776,N_15402,N_15578);
nor U17777 (N_17777,N_14116,N_15937);
nor U17778 (N_17778,N_15808,N_15169);
nand U17779 (N_17779,N_15491,N_14648);
or U17780 (N_17780,N_15556,N_15665);
nor U17781 (N_17781,N_14382,N_14358);
nand U17782 (N_17782,N_14061,N_14199);
and U17783 (N_17783,N_15413,N_14600);
and U17784 (N_17784,N_14427,N_15223);
nand U17785 (N_17785,N_15676,N_15067);
xor U17786 (N_17786,N_14941,N_14905);
or U17787 (N_17787,N_15806,N_14291);
or U17788 (N_17788,N_15784,N_15593);
xnor U17789 (N_17789,N_15829,N_15313);
nor U17790 (N_17790,N_14700,N_15763);
nand U17791 (N_17791,N_15023,N_15306);
xnor U17792 (N_17792,N_14967,N_15975);
and U17793 (N_17793,N_14900,N_14059);
nor U17794 (N_17794,N_15282,N_14572);
and U17795 (N_17795,N_15448,N_14058);
nand U17796 (N_17796,N_14098,N_15965);
nand U17797 (N_17797,N_15107,N_15180);
xor U17798 (N_17798,N_14052,N_14555);
and U17799 (N_17799,N_15289,N_15833);
and U17800 (N_17800,N_14082,N_15232);
xnor U17801 (N_17801,N_15220,N_14280);
xor U17802 (N_17802,N_14207,N_14206);
and U17803 (N_17803,N_15638,N_14606);
and U17804 (N_17804,N_14923,N_14631);
nor U17805 (N_17805,N_15245,N_14944);
and U17806 (N_17806,N_15778,N_15231);
xnor U17807 (N_17807,N_14338,N_14954);
nand U17808 (N_17808,N_14224,N_14456);
xor U17809 (N_17809,N_15433,N_15395);
xnor U17810 (N_17810,N_15672,N_15321);
nand U17811 (N_17811,N_14885,N_15628);
xnor U17812 (N_17812,N_15126,N_14950);
or U17813 (N_17813,N_14558,N_15614);
nor U17814 (N_17814,N_14909,N_14134);
nand U17815 (N_17815,N_14799,N_15334);
xnor U17816 (N_17816,N_15046,N_15050);
or U17817 (N_17817,N_15290,N_15364);
nor U17818 (N_17818,N_14647,N_14521);
or U17819 (N_17819,N_14648,N_15633);
or U17820 (N_17820,N_15345,N_15817);
nand U17821 (N_17821,N_15927,N_14529);
nor U17822 (N_17822,N_15027,N_14512);
or U17823 (N_17823,N_14070,N_15731);
xor U17824 (N_17824,N_15991,N_15547);
xnor U17825 (N_17825,N_14003,N_15871);
xor U17826 (N_17826,N_14364,N_14229);
and U17827 (N_17827,N_14663,N_14891);
nor U17828 (N_17828,N_15149,N_14238);
and U17829 (N_17829,N_15741,N_15097);
nand U17830 (N_17830,N_14771,N_15553);
nand U17831 (N_17831,N_15660,N_15933);
and U17832 (N_17832,N_14857,N_15238);
nand U17833 (N_17833,N_15626,N_14298);
xnor U17834 (N_17834,N_14115,N_14349);
or U17835 (N_17835,N_15117,N_14508);
and U17836 (N_17836,N_14348,N_15574);
xor U17837 (N_17837,N_15246,N_14724);
xor U17838 (N_17838,N_15254,N_14810);
or U17839 (N_17839,N_15266,N_14638);
nor U17840 (N_17840,N_15991,N_14196);
nor U17841 (N_17841,N_15426,N_15734);
or U17842 (N_17842,N_15569,N_14726);
xor U17843 (N_17843,N_14397,N_14431);
or U17844 (N_17844,N_14066,N_14149);
xnor U17845 (N_17845,N_15809,N_15264);
xor U17846 (N_17846,N_14330,N_14477);
or U17847 (N_17847,N_15429,N_14178);
and U17848 (N_17848,N_14466,N_15692);
nand U17849 (N_17849,N_15731,N_14640);
nor U17850 (N_17850,N_14821,N_15967);
and U17851 (N_17851,N_14254,N_14109);
nand U17852 (N_17852,N_15332,N_15288);
nand U17853 (N_17853,N_14983,N_15738);
nand U17854 (N_17854,N_15790,N_15511);
nor U17855 (N_17855,N_14146,N_15275);
xor U17856 (N_17856,N_14584,N_15199);
and U17857 (N_17857,N_14424,N_15424);
nor U17858 (N_17858,N_15331,N_14196);
nor U17859 (N_17859,N_14539,N_15619);
or U17860 (N_17860,N_14928,N_14908);
nor U17861 (N_17861,N_14254,N_15408);
nand U17862 (N_17862,N_15606,N_15990);
nand U17863 (N_17863,N_15276,N_15391);
xor U17864 (N_17864,N_14956,N_15948);
and U17865 (N_17865,N_15752,N_15822);
and U17866 (N_17866,N_14471,N_15440);
or U17867 (N_17867,N_15598,N_15678);
nand U17868 (N_17868,N_14145,N_15372);
and U17869 (N_17869,N_15720,N_14527);
and U17870 (N_17870,N_15972,N_15602);
nor U17871 (N_17871,N_14947,N_15137);
or U17872 (N_17872,N_15857,N_14527);
and U17873 (N_17873,N_15452,N_14367);
nand U17874 (N_17874,N_14077,N_15011);
nor U17875 (N_17875,N_14770,N_14126);
nor U17876 (N_17876,N_15697,N_15900);
nor U17877 (N_17877,N_15569,N_15006);
or U17878 (N_17878,N_14007,N_14086);
nand U17879 (N_17879,N_14202,N_15534);
and U17880 (N_17880,N_15564,N_15782);
or U17881 (N_17881,N_15998,N_14409);
and U17882 (N_17882,N_14305,N_15218);
nor U17883 (N_17883,N_14435,N_15108);
or U17884 (N_17884,N_15916,N_15879);
nor U17885 (N_17885,N_14226,N_15855);
nand U17886 (N_17886,N_15704,N_14386);
nand U17887 (N_17887,N_14240,N_15896);
nand U17888 (N_17888,N_15149,N_14862);
or U17889 (N_17889,N_14298,N_15676);
and U17890 (N_17890,N_15110,N_14865);
nand U17891 (N_17891,N_15202,N_15089);
xor U17892 (N_17892,N_14431,N_14560);
nor U17893 (N_17893,N_14069,N_14832);
nand U17894 (N_17894,N_15489,N_14256);
or U17895 (N_17895,N_14936,N_14618);
nor U17896 (N_17896,N_15754,N_14356);
and U17897 (N_17897,N_14302,N_15618);
xor U17898 (N_17898,N_15877,N_15583);
and U17899 (N_17899,N_14092,N_14041);
xnor U17900 (N_17900,N_14518,N_15971);
xnor U17901 (N_17901,N_15265,N_14524);
and U17902 (N_17902,N_15220,N_15275);
or U17903 (N_17903,N_14971,N_14329);
nor U17904 (N_17904,N_15156,N_15364);
or U17905 (N_17905,N_15393,N_14334);
and U17906 (N_17906,N_14171,N_14867);
nand U17907 (N_17907,N_14813,N_15794);
or U17908 (N_17908,N_15224,N_15809);
nand U17909 (N_17909,N_15566,N_14444);
xor U17910 (N_17910,N_15623,N_14162);
nor U17911 (N_17911,N_14463,N_15478);
nor U17912 (N_17912,N_15703,N_14275);
xor U17913 (N_17913,N_15384,N_14988);
nor U17914 (N_17914,N_14869,N_15611);
nand U17915 (N_17915,N_15618,N_15307);
nand U17916 (N_17916,N_14397,N_14858);
xnor U17917 (N_17917,N_14496,N_14809);
xor U17918 (N_17918,N_14123,N_14305);
nand U17919 (N_17919,N_15494,N_14556);
or U17920 (N_17920,N_14172,N_15766);
xor U17921 (N_17921,N_15734,N_15363);
xnor U17922 (N_17922,N_14184,N_14056);
or U17923 (N_17923,N_14719,N_15657);
xnor U17924 (N_17924,N_14397,N_14765);
nand U17925 (N_17925,N_14757,N_15546);
xor U17926 (N_17926,N_14009,N_15291);
nand U17927 (N_17927,N_15623,N_15132);
and U17928 (N_17928,N_15614,N_14525);
xor U17929 (N_17929,N_14120,N_14329);
or U17930 (N_17930,N_14008,N_14332);
nor U17931 (N_17931,N_14932,N_14061);
nand U17932 (N_17932,N_15363,N_15823);
nand U17933 (N_17933,N_14477,N_14404);
or U17934 (N_17934,N_14580,N_15082);
xnor U17935 (N_17935,N_15865,N_14762);
and U17936 (N_17936,N_15046,N_14362);
and U17937 (N_17937,N_14459,N_14879);
or U17938 (N_17938,N_14795,N_14746);
nand U17939 (N_17939,N_15229,N_14300);
nand U17940 (N_17940,N_15415,N_14313);
nand U17941 (N_17941,N_15534,N_14376);
or U17942 (N_17942,N_14907,N_15118);
xnor U17943 (N_17943,N_14287,N_15444);
xor U17944 (N_17944,N_14056,N_14205);
and U17945 (N_17945,N_15268,N_14096);
xor U17946 (N_17946,N_15159,N_14677);
nor U17947 (N_17947,N_14524,N_14948);
nor U17948 (N_17948,N_15190,N_14168);
xor U17949 (N_17949,N_14385,N_15908);
nand U17950 (N_17950,N_14292,N_15302);
and U17951 (N_17951,N_14331,N_14936);
nor U17952 (N_17952,N_15585,N_15761);
xnor U17953 (N_17953,N_15759,N_15504);
or U17954 (N_17954,N_14721,N_14998);
and U17955 (N_17955,N_15862,N_15031);
nand U17956 (N_17956,N_14892,N_15208);
nand U17957 (N_17957,N_15263,N_15441);
xor U17958 (N_17958,N_15593,N_15317);
and U17959 (N_17959,N_15825,N_14943);
nor U17960 (N_17960,N_15195,N_14393);
nor U17961 (N_17961,N_15210,N_14969);
nand U17962 (N_17962,N_15338,N_15484);
nor U17963 (N_17963,N_14540,N_15756);
xor U17964 (N_17964,N_14621,N_15370);
nand U17965 (N_17965,N_15482,N_15228);
nand U17966 (N_17966,N_15412,N_14195);
or U17967 (N_17967,N_14914,N_15379);
xnor U17968 (N_17968,N_14014,N_14717);
nand U17969 (N_17969,N_14002,N_15162);
or U17970 (N_17970,N_14547,N_14990);
or U17971 (N_17971,N_14421,N_14004);
xor U17972 (N_17972,N_14994,N_15870);
and U17973 (N_17973,N_14936,N_14268);
and U17974 (N_17974,N_14546,N_14129);
nand U17975 (N_17975,N_15650,N_14493);
nor U17976 (N_17976,N_15641,N_14379);
xor U17977 (N_17977,N_15153,N_15120);
and U17978 (N_17978,N_14701,N_14158);
or U17979 (N_17979,N_14365,N_15180);
nand U17980 (N_17980,N_14842,N_14531);
or U17981 (N_17981,N_15995,N_14386);
xnor U17982 (N_17982,N_14938,N_15241);
nand U17983 (N_17983,N_14193,N_14581);
or U17984 (N_17984,N_15277,N_14822);
or U17985 (N_17985,N_14689,N_15840);
or U17986 (N_17986,N_15863,N_15734);
and U17987 (N_17987,N_15672,N_14712);
xnor U17988 (N_17988,N_15162,N_14793);
and U17989 (N_17989,N_14546,N_14901);
xor U17990 (N_17990,N_14961,N_14861);
and U17991 (N_17991,N_15320,N_15452);
nand U17992 (N_17992,N_14491,N_14421);
xnor U17993 (N_17993,N_14016,N_15896);
nand U17994 (N_17994,N_14012,N_15871);
nor U17995 (N_17995,N_15973,N_15979);
nand U17996 (N_17996,N_15421,N_14165);
or U17997 (N_17997,N_14035,N_14040);
and U17998 (N_17998,N_14687,N_15037);
nand U17999 (N_17999,N_14868,N_15762);
and U18000 (N_18000,N_16106,N_17939);
xnor U18001 (N_18001,N_17140,N_16740);
or U18002 (N_18002,N_17531,N_16987);
and U18003 (N_18003,N_17847,N_17527);
and U18004 (N_18004,N_16452,N_16030);
xnor U18005 (N_18005,N_16277,N_16454);
or U18006 (N_18006,N_16958,N_16310);
nand U18007 (N_18007,N_16423,N_17500);
nand U18008 (N_18008,N_16267,N_16535);
xnor U18009 (N_18009,N_16217,N_17228);
and U18010 (N_18010,N_17843,N_17578);
and U18011 (N_18011,N_17923,N_16603);
nand U18012 (N_18012,N_17605,N_16293);
nor U18013 (N_18013,N_17756,N_17060);
xnor U18014 (N_18014,N_16248,N_17055);
or U18015 (N_18015,N_17774,N_17648);
or U18016 (N_18016,N_16013,N_16774);
and U18017 (N_18017,N_16968,N_17088);
nand U18018 (N_18018,N_16048,N_16595);
and U18019 (N_18019,N_17775,N_16533);
and U18020 (N_18020,N_16464,N_17800);
xnor U18021 (N_18021,N_16931,N_17022);
xnor U18022 (N_18022,N_16653,N_16004);
and U18023 (N_18023,N_16144,N_16373);
or U18024 (N_18024,N_16794,N_16566);
nand U18025 (N_18025,N_17600,N_17083);
and U18026 (N_18026,N_17767,N_17721);
nand U18027 (N_18027,N_16238,N_17810);
xnor U18028 (N_18028,N_16342,N_17434);
nand U18029 (N_18029,N_16359,N_16610);
or U18030 (N_18030,N_17248,N_17682);
and U18031 (N_18031,N_16116,N_16509);
or U18032 (N_18032,N_17076,N_16468);
xor U18033 (N_18033,N_17257,N_16350);
or U18034 (N_18034,N_17120,N_16447);
nand U18035 (N_18035,N_16027,N_16531);
or U18036 (N_18036,N_16403,N_17877);
xnor U18037 (N_18037,N_17370,N_16368);
nor U18038 (N_18038,N_17512,N_16646);
or U18039 (N_18039,N_17040,N_16939);
nand U18040 (N_18040,N_17441,N_16916);
xor U18041 (N_18041,N_17301,N_16021);
and U18042 (N_18042,N_16031,N_17121);
xnor U18043 (N_18043,N_16001,N_17156);
nand U18044 (N_18044,N_16126,N_16710);
nor U18045 (N_18045,N_17525,N_16131);
nand U18046 (N_18046,N_16758,N_16019);
or U18047 (N_18047,N_17149,N_17241);
or U18048 (N_18048,N_17322,N_17957);
or U18049 (N_18049,N_17197,N_16210);
nand U18050 (N_18050,N_16572,N_16601);
nand U18051 (N_18051,N_16881,N_17015);
nand U18052 (N_18052,N_16777,N_16216);
or U18053 (N_18053,N_16457,N_16283);
nand U18054 (N_18054,N_17354,N_16755);
or U18055 (N_18055,N_17179,N_17065);
nand U18056 (N_18056,N_16441,N_17908);
nor U18057 (N_18057,N_17757,N_17989);
or U18058 (N_18058,N_17543,N_16686);
xor U18059 (N_18059,N_17987,N_17107);
or U18060 (N_18060,N_17632,N_17675);
or U18061 (N_18061,N_17590,N_16192);
nand U18062 (N_18062,N_16615,N_16049);
xor U18063 (N_18063,N_17876,N_16833);
xnor U18064 (N_18064,N_17177,N_17153);
or U18065 (N_18065,N_17504,N_16235);
nand U18066 (N_18066,N_17075,N_16651);
xor U18067 (N_18067,N_16800,N_17367);
nand U18068 (N_18068,N_16177,N_17548);
or U18069 (N_18069,N_16308,N_16257);
nor U18070 (N_18070,N_17343,N_16772);
or U18071 (N_18071,N_17452,N_16827);
xor U18072 (N_18072,N_17674,N_16547);
nand U18073 (N_18073,N_16874,N_17984);
nor U18074 (N_18074,N_17857,N_16585);
or U18075 (N_18075,N_17313,N_16171);
and U18076 (N_18076,N_16146,N_16934);
xor U18077 (N_18077,N_16024,N_16255);
nor U18078 (N_18078,N_17701,N_16782);
xor U18079 (N_18079,N_17713,N_17379);
or U18080 (N_18080,N_16434,N_17909);
nand U18081 (N_18081,N_16075,N_17681);
or U18082 (N_18082,N_17113,N_17032);
or U18083 (N_18083,N_17489,N_17583);
or U18084 (N_18084,N_16925,N_16839);
nor U18085 (N_18085,N_17031,N_16504);
and U18086 (N_18086,N_17698,N_17192);
nor U18087 (N_18087,N_17263,N_16776);
xnor U18088 (N_18088,N_17850,N_17401);
xnor U18089 (N_18089,N_16885,N_17963);
xnor U18090 (N_18090,N_17959,N_17488);
nor U18091 (N_18091,N_16406,N_16014);
nand U18092 (N_18092,N_17705,N_16204);
and U18093 (N_18093,N_17330,N_17398);
xor U18094 (N_18094,N_16539,N_16395);
nor U18095 (N_18095,N_16424,N_16775);
xor U18096 (N_18096,N_17968,N_16713);
nand U18097 (N_18097,N_17769,N_16570);
nand U18098 (N_18098,N_16440,N_16889);
nor U18099 (N_18099,N_16750,N_16918);
xor U18100 (N_18100,N_17209,N_17509);
and U18101 (N_18101,N_16157,N_17916);
xnor U18102 (N_18102,N_16955,N_17169);
or U18103 (N_18103,N_17455,N_17123);
nor U18104 (N_18104,N_16702,N_17686);
and U18105 (N_18105,N_17715,N_17386);
nor U18106 (N_18106,N_16599,N_16711);
or U18107 (N_18107,N_16767,N_17943);
or U18108 (N_18108,N_16561,N_16695);
and U18109 (N_18109,N_16278,N_17226);
or U18110 (N_18110,N_17889,N_16730);
and U18111 (N_18111,N_16554,N_17298);
or U18112 (N_18112,N_16642,N_16245);
nor U18113 (N_18113,N_17714,N_16816);
nand U18114 (N_18114,N_16505,N_17315);
xnor U18115 (N_18115,N_16297,N_17607);
nor U18116 (N_18116,N_16324,N_17501);
xnor U18117 (N_18117,N_17419,N_17834);
nor U18118 (N_18118,N_16069,N_16002);
nor U18119 (N_18119,N_16924,N_16160);
nand U18120 (N_18120,N_17790,N_17855);
and U18121 (N_18121,N_16296,N_17360);
xnor U18122 (N_18122,N_17744,N_17299);
or U18123 (N_18123,N_17027,N_17069);
xor U18124 (N_18124,N_16648,N_16259);
nand U18125 (N_18125,N_17998,N_17297);
nor U18126 (N_18126,N_16562,N_16633);
or U18127 (N_18127,N_16053,N_16712);
nand U18128 (N_18128,N_16147,N_17026);
nand U18129 (N_18129,N_16335,N_16158);
and U18130 (N_18130,N_17972,N_16071);
nor U18131 (N_18131,N_16046,N_16594);
nand U18132 (N_18132,N_17663,N_17851);
nand U18133 (N_18133,N_16471,N_17584);
nand U18134 (N_18134,N_16841,N_17796);
and U18135 (N_18135,N_16260,N_17278);
or U18136 (N_18136,N_16607,N_17345);
nor U18137 (N_18137,N_16903,N_16307);
and U18138 (N_18138,N_16745,N_16191);
nor U18139 (N_18139,N_16433,N_17090);
nand U18140 (N_18140,N_17001,N_17637);
nand U18141 (N_18141,N_17634,N_17230);
nor U18142 (N_18142,N_16085,N_17164);
nor U18143 (N_18143,N_16929,N_16732);
or U18144 (N_18144,N_16136,N_17567);
nor U18145 (N_18145,N_16386,N_17802);
xor U18146 (N_18146,N_17539,N_17357);
nor U18147 (N_18147,N_16028,N_17025);
nand U18148 (N_18148,N_17021,N_17665);
or U18149 (N_18149,N_17556,N_17372);
and U18150 (N_18150,N_17063,N_16218);
xnor U18151 (N_18151,N_16460,N_17150);
nand U18152 (N_18152,N_16211,N_16806);
and U18153 (N_18153,N_16543,N_17871);
and U18154 (N_18154,N_17560,N_17669);
nor U18155 (N_18155,N_16417,N_16241);
and U18156 (N_18156,N_17717,N_16804);
or U18157 (N_18157,N_17788,N_17945);
nor U18158 (N_18158,N_17450,N_16232);
nor U18159 (N_18159,N_17430,N_17294);
or U18160 (N_18160,N_16995,N_16792);
nor U18161 (N_18161,N_16606,N_16401);
nand U18162 (N_18162,N_16446,N_16220);
xor U18163 (N_18163,N_17824,N_17552);
or U18164 (N_18164,N_16006,N_16033);
xnor U18165 (N_18165,N_16057,N_17125);
nor U18166 (N_18166,N_17251,N_16382);
nand U18167 (N_18167,N_16381,N_17724);
or U18168 (N_18168,N_16518,N_16735);
nor U18169 (N_18169,N_16344,N_16643);
or U18170 (N_18170,N_17384,N_16432);
or U18171 (N_18171,N_17284,N_17059);
nand U18172 (N_18172,N_16528,N_17199);
or U18173 (N_18173,N_16760,N_17348);
nor U18174 (N_18174,N_16664,N_17247);
and U18175 (N_18175,N_16685,N_16279);
nor U18176 (N_18176,N_16835,N_16892);
xor U18177 (N_18177,N_17352,N_17653);
or U18178 (N_18178,N_17128,N_16943);
or U18179 (N_18179,N_16917,N_16938);
nand U18180 (N_18180,N_17630,N_17776);
and U18181 (N_18181,N_17335,N_17493);
and U18182 (N_18182,N_17369,N_17534);
or U18183 (N_18183,N_16761,N_17244);
or U18184 (N_18184,N_17574,N_16020);
nand U18185 (N_18185,N_16997,N_16857);
or U18186 (N_18186,N_16387,N_17816);
xor U18187 (N_18187,N_16356,N_17720);
or U18188 (N_18188,N_17795,N_16207);
xnor U18189 (N_18189,N_17351,N_16465);
and U18190 (N_18190,N_17437,N_16112);
nor U18191 (N_18191,N_16617,N_17426);
or U18192 (N_18192,N_16203,N_17271);
xnor U18193 (N_18193,N_17180,N_16899);
xor U18194 (N_18194,N_16407,N_16583);
nand U18195 (N_18195,N_17087,N_17115);
and U18196 (N_18196,N_17198,N_17141);
and U18197 (N_18197,N_16631,N_16715);
nor U18198 (N_18198,N_17119,N_16265);
and U18199 (N_18199,N_17011,N_16962);
nand U18200 (N_18200,N_16485,N_17570);
nand U18201 (N_18201,N_17741,N_17323);
nor U18202 (N_18202,N_17456,N_17207);
nand U18203 (N_18203,N_17902,N_16280);
xor U18204 (N_18204,N_17884,N_17887);
nand U18205 (N_18205,N_16023,N_16162);
or U18206 (N_18206,N_16757,N_17392);
nor U18207 (N_18207,N_16953,N_17097);
xnor U18208 (N_18208,N_16196,N_16975);
and U18209 (N_18209,N_16513,N_16863);
nor U18210 (N_18210,N_16669,N_17418);
nor U18211 (N_18211,N_16442,N_16329);
xor U18212 (N_18212,N_17738,N_16638);
or U18213 (N_18213,N_16332,N_16809);
nand U18214 (N_18214,N_17371,N_17174);
nand U18215 (N_18215,N_17173,N_17091);
xor U18216 (N_18216,N_16438,N_16898);
and U18217 (N_18217,N_16920,N_16404);
nand U18218 (N_18218,N_16313,N_16627);
xnor U18219 (N_18219,N_16515,N_17894);
nor U18220 (N_18220,N_17865,N_16506);
nor U18221 (N_18221,N_17696,N_16926);
nor U18222 (N_18222,N_17451,N_16243);
xnor U18223 (N_18223,N_16078,N_16682);
nor U18224 (N_18224,N_17007,N_17996);
and U18225 (N_18225,N_16634,N_16834);
xnor U18226 (N_18226,N_17403,N_16036);
xor U18227 (N_18227,N_16054,N_17259);
xor U18228 (N_18228,N_17457,N_17050);
nor U18229 (N_18229,N_16875,N_16910);
nor U18230 (N_18230,N_17240,N_17792);
and U18231 (N_18231,N_16683,N_17073);
nand U18232 (N_18232,N_16070,N_16083);
xor U18233 (N_18233,N_16848,N_16213);
or U18234 (N_18234,N_16529,N_17654);
xor U18235 (N_18235,N_17528,N_16593);
or U18236 (N_18236,N_17289,N_16587);
xnor U18237 (N_18237,N_17707,N_17368);
xor U18238 (N_18238,N_16166,N_16436);
and U18239 (N_18239,N_16309,N_16428);
nand U18240 (N_18240,N_16357,N_17603);
xor U18241 (N_18241,N_17017,N_17978);
nor U18242 (N_18242,N_16110,N_17464);
nor U18243 (N_18243,N_16497,N_17644);
xnor U18244 (N_18244,N_17684,N_16674);
or U18245 (N_18245,N_16392,N_16303);
xnor U18246 (N_18246,N_17411,N_17553);
or U18247 (N_18247,N_16415,N_16676);
nor U18248 (N_18248,N_17549,N_17380);
and U18249 (N_18249,N_16604,N_17471);
xnor U18250 (N_18250,N_16622,N_17186);
and U18251 (N_18251,N_17160,N_16459);
and U18252 (N_18252,N_17893,N_16410);
xor U18253 (N_18253,N_17424,N_17821);
or U18254 (N_18254,N_16005,N_17797);
xor U18255 (N_18255,N_17687,N_17237);
xnor U18256 (N_18256,N_17109,N_17196);
xnor U18257 (N_18257,N_16467,N_16744);
nor U18258 (N_18258,N_17536,N_16950);
xor U18259 (N_18259,N_16668,N_17317);
nand U18260 (N_18260,N_17854,N_17277);
xor U18261 (N_18261,N_16273,N_17117);
nand U18262 (N_18262,N_16319,N_17641);
or U18263 (N_18263,N_16222,N_17729);
or U18264 (N_18264,N_16107,N_17999);
and U18265 (N_18265,N_16705,N_17049);
or U18266 (N_18266,N_16941,N_16065);
nand U18267 (N_18267,N_17291,N_16519);
nand U18268 (N_18268,N_16501,N_17523);
nor U18269 (N_18269,N_17693,N_17416);
nor U18270 (N_18270,N_16261,N_17642);
or U18271 (N_18271,N_17635,N_17918);
nor U18272 (N_18272,N_16099,N_16655);
and U18273 (N_18273,N_16473,N_17949);
or U18274 (N_18274,N_17895,N_16100);
or U18275 (N_18275,N_16236,N_17718);
and U18276 (N_18276,N_16589,N_16117);
xor U18277 (N_18277,N_17429,N_17146);
nand U18278 (N_18278,N_16673,N_17377);
xnor U18279 (N_18279,N_16427,N_16814);
nand U18280 (N_18280,N_17524,N_16853);
nor U18281 (N_18281,N_17236,N_16972);
nor U18282 (N_18282,N_16625,N_16867);
nand U18283 (N_18283,N_16003,N_17563);
xnor U18284 (N_18284,N_16154,N_16068);
or U18285 (N_18285,N_16345,N_17564);
nor U18286 (N_18286,N_16989,N_16797);
or U18287 (N_18287,N_16872,N_16060);
nand U18288 (N_18288,N_16055,N_17829);
xnor U18289 (N_18289,N_16778,N_16185);
or U18290 (N_18290,N_16688,N_16524);
nor U18291 (N_18291,N_16571,N_16487);
nand U18292 (N_18292,N_16591,N_16649);
nand U18293 (N_18293,N_17839,N_17074);
nor U18294 (N_18294,N_16022,N_17766);
and U18295 (N_18295,N_17596,N_17703);
xnor U18296 (N_18296,N_16798,N_16118);
or U18297 (N_18297,N_17608,N_17482);
nand U18298 (N_18298,N_17734,N_17591);
and U18299 (N_18299,N_16544,N_17387);
nand U18300 (N_18300,N_17579,N_16693);
nand U18301 (N_18301,N_17935,N_16275);
nand U18302 (N_18302,N_16064,N_17214);
xnor U18303 (N_18303,N_16720,N_16435);
nand U18304 (N_18304,N_16380,N_17472);
xnor U18305 (N_18305,N_16129,N_16994);
xnor U18306 (N_18306,N_16374,N_16152);
xnor U18307 (N_18307,N_16510,N_16795);
nand U18308 (N_18308,N_17666,N_17185);
nand U18309 (N_18309,N_17053,N_17882);
nor U18310 (N_18310,N_16957,N_17588);
xor U18311 (N_18311,N_16095,N_16907);
nor U18312 (N_18312,N_16305,N_17872);
and U18313 (N_18313,N_16781,N_17043);
and U18314 (N_18314,N_17448,N_16379);
and U18315 (N_18315,N_17012,N_17431);
xnor U18316 (N_18316,N_17933,N_17182);
xor U18317 (N_18317,N_16932,N_16679);
and U18318 (N_18318,N_17395,N_17530);
xor U18319 (N_18319,N_17941,N_17645);
nand U18320 (N_18320,N_17433,N_17167);
xnor U18321 (N_18321,N_16808,N_17436);
and U18322 (N_18322,N_16176,N_17393);
xnor U18323 (N_18323,N_16251,N_17730);
nand U18324 (N_18324,N_17378,N_17709);
xor U18325 (N_18325,N_16829,N_16791);
nor U18326 (N_18326,N_17355,N_16551);
or U18327 (N_18327,N_16480,N_17274);
xor U18328 (N_18328,N_17736,N_16223);
or U18329 (N_18329,N_16090,N_17511);
or U18330 (N_18330,N_16323,N_16680);
nor U18331 (N_18331,N_16658,N_17799);
and U18332 (N_18332,N_16142,N_16790);
nor U18333 (N_18333,N_17390,N_16897);
nor U18334 (N_18334,N_17764,N_16276);
or U18335 (N_18335,N_17901,N_17415);
nand U18336 (N_18336,N_16936,N_17013);
or U18337 (N_18337,N_17005,N_17926);
nor U18338 (N_18338,N_17833,N_17235);
xor U18339 (N_18339,N_17085,N_16352);
and U18340 (N_18340,N_16405,N_17442);
or U18341 (N_18341,N_17510,N_17805);
or U18342 (N_18342,N_16824,N_16895);
or U18343 (N_18343,N_17474,N_16822);
and U18344 (N_18344,N_16179,N_17231);
or U18345 (N_18345,N_16443,N_16224);
or U18346 (N_18346,N_17618,N_16492);
and U18347 (N_18347,N_17147,N_16662);
or U18348 (N_18348,N_17084,N_17897);
and U18349 (N_18349,N_16219,N_17316);
and U18350 (N_18350,N_17745,N_17782);
and U18351 (N_18351,N_17862,N_17320);
nor U18352 (N_18352,N_16449,N_16988);
nand U18353 (N_18353,N_17565,N_16807);
and U18354 (N_18354,N_17879,N_17661);
and U18355 (N_18355,N_17498,N_17157);
or U18356 (N_18356,N_17194,N_16453);
or U18357 (N_18357,N_17212,N_16109);
or U18358 (N_18358,N_16681,N_17658);
and U18359 (N_18359,N_17657,N_17903);
nor U18360 (N_18360,N_16476,N_16696);
nand U18361 (N_18361,N_17914,N_16855);
xor U18362 (N_18362,N_16038,N_16143);
xnor U18363 (N_18363,N_16714,N_16780);
and U18364 (N_18364,N_17815,N_17947);
or U18365 (N_18365,N_17195,N_17203);
nor U18366 (N_18366,N_16281,N_17144);
and U18367 (N_18367,N_17751,N_16115);
xnor U18368 (N_18368,N_17204,N_17062);
or U18369 (N_18369,N_16522,N_17848);
nor U18370 (N_18370,N_16093,N_16151);
xnor U18371 (N_18371,N_16161,N_16418);
nand U18372 (N_18372,N_17628,N_16470);
or U18373 (N_18373,N_16956,N_16256);
nand U18374 (N_18374,N_17760,N_16128);
xor U18375 (N_18375,N_17508,N_17977);
and U18376 (N_18376,N_17242,N_16164);
and U18377 (N_18377,N_16982,N_17626);
or U18378 (N_18378,N_17421,N_17891);
nand U18379 (N_18379,N_16378,N_17706);
nor U18380 (N_18380,N_17470,N_16555);
or U18381 (N_18381,N_16890,N_16516);
nor U18382 (N_18382,N_17809,N_16706);
nand U18383 (N_18383,N_17610,N_17211);
nand U18384 (N_18384,N_16072,N_17422);
nand U18385 (N_18385,N_17708,N_16495);
nor U18386 (N_18386,N_16302,N_17927);
and U18387 (N_18387,N_17814,N_17328);
nor U18388 (N_18388,N_16900,N_16271);
or U18389 (N_18389,N_17159,N_16489);
or U18390 (N_18390,N_17331,N_17621);
nand U18391 (N_18391,N_17417,N_16201);
or U18392 (N_18392,N_17990,N_17719);
and U18393 (N_18393,N_16704,N_16353);
and U18394 (N_18394,N_17443,N_17787);
nand U18395 (N_18395,N_16840,N_16514);
and U18396 (N_18396,N_16865,N_16145);
and U18397 (N_18397,N_17823,N_17000);
xor U18398 (N_18398,N_17223,N_17342);
and U18399 (N_18399,N_17942,N_17318);
or U18400 (N_18400,N_17333,N_16844);
nor U18401 (N_18401,N_17307,N_16878);
xnor U18402 (N_18402,N_16326,N_16960);
or U18403 (N_18403,N_16709,N_17778);
nand U18404 (N_18404,N_16823,N_17620);
and U18405 (N_18405,N_17832,N_16946);
nand U18406 (N_18406,N_16050,N_17071);
or U18407 (N_18407,N_17576,N_17601);
or U18408 (N_18408,N_16333,N_16475);
and U18409 (N_18409,N_16619,N_16092);
xor U18410 (N_18410,N_16450,N_17910);
or U18411 (N_18411,N_16478,N_17688);
or U18412 (N_18412,N_17282,N_17704);
or U18413 (N_18413,N_16175,N_17365);
and U18414 (N_18414,N_17753,N_16067);
or U18415 (N_18415,N_16289,N_16981);
or U18416 (N_18416,N_17826,N_17092);
and U18417 (N_18417,N_17358,N_16237);
nor U18418 (N_18418,N_16748,N_16999);
nor U18419 (N_18419,N_16877,N_17639);
xor U18420 (N_18420,N_16752,N_16376);
and U18421 (N_18421,N_17986,N_17239);
or U18422 (N_18422,N_16206,N_16933);
nand U18423 (N_18423,N_17602,N_17541);
or U18424 (N_18424,N_16061,N_16422);
xor U18425 (N_18425,N_16399,N_17184);
and U18426 (N_18426,N_17699,N_17461);
and U18427 (N_18427,N_16202,N_17400);
nor U18428 (N_18428,N_16596,N_17300);
nand U18429 (N_18429,N_17373,N_16810);
xnor U18430 (N_18430,N_16976,N_17811);
or U18431 (N_18431,N_17232,N_17103);
nand U18432 (N_18432,N_17649,N_17582);
nor U18433 (N_18433,N_16908,N_16194);
and U18434 (N_18434,N_17420,N_16361);
nand U18435 (N_18435,N_17846,N_17038);
nor U18436 (N_18436,N_17225,N_17030);
nand U18437 (N_18437,N_17870,N_17880);
and U18438 (N_18438,N_16198,N_17612);
nand U18439 (N_18439,N_17445,N_17206);
nor U18440 (N_18440,N_17311,N_17780);
nand U18441 (N_18441,N_16212,N_16155);
or U18442 (N_18442,N_16098,N_16541);
or U18443 (N_18443,N_16564,N_16882);
nand U18444 (N_18444,N_16598,N_17727);
or U18445 (N_18445,N_16388,N_16338);
and U18446 (N_18446,N_17773,N_16985);
nand U18447 (N_18447,N_17516,N_17878);
and U18448 (N_18448,N_17490,N_16360);
nor U18449 (N_18449,N_17408,N_16312);
nand U18450 (N_18450,N_16025,N_17992);
or U18451 (N_18451,N_16645,N_16805);
nor U18452 (N_18452,N_17218,N_17733);
xnor U18453 (N_18453,N_17568,N_17670);
or U18454 (N_18454,N_17034,N_17685);
nor U18455 (N_18455,N_17312,N_17633);
and U18456 (N_18456,N_16456,N_16971);
or U18457 (N_18457,N_17382,N_16614);
nor U18458 (N_18458,N_16304,N_17340);
and U18459 (N_18459,N_16860,N_16836);
nand U18460 (N_18460,N_16852,N_17469);
or U18461 (N_18461,N_16828,N_17279);
xnor U18462 (N_18462,N_17965,N_16314);
or U18463 (N_18463,N_17656,N_16773);
or U18464 (N_18464,N_17946,N_17677);
or U18465 (N_18465,N_16940,N_16722);
or U18466 (N_18466,N_17517,N_16121);
nor U18467 (N_18467,N_16383,N_16719);
nand U18468 (N_18468,N_16862,N_16490);
xnor U18469 (N_18469,N_16153,N_17459);
nor U18470 (N_18470,N_16045,N_17252);
nor U18471 (N_18471,N_16992,N_17138);
or U18472 (N_18472,N_16197,N_16851);
or U18473 (N_18473,N_16097,N_16796);
and U18474 (N_18474,N_17555,N_17671);
nand U18475 (N_18475,N_17822,N_16978);
nand U18476 (N_18476,N_17913,N_16486);
and U18477 (N_18477,N_16831,N_17163);
nand U18478 (N_18478,N_17353,N_17495);
nand U18479 (N_18479,N_17726,N_16463);
nor U18480 (N_18480,N_16915,N_16734);
and U18481 (N_18481,N_17246,N_17858);
nor U18482 (N_18482,N_17404,N_17462);
xnor U18483 (N_18483,N_17364,N_17743);
nand U18484 (N_18484,N_16784,N_17638);
or U18485 (N_18485,N_16292,N_17413);
and U18486 (N_18486,N_16743,N_16868);
nor U18487 (N_18487,N_17327,N_16665);
or U18488 (N_18488,N_16412,N_16644);
or U18489 (N_18489,N_16254,N_16409);
nor U18490 (N_18490,N_16728,N_16843);
or U18491 (N_18491,N_16058,N_17347);
nand U18492 (N_18492,N_16268,N_16859);
and U18493 (N_18493,N_16375,N_17310);
nor U18494 (N_18494,N_17366,N_17072);
nand U18495 (N_18495,N_17931,N_16891);
xor U18496 (N_18496,N_17341,N_16911);
xnor U18497 (N_18497,N_16079,N_17142);
nand U18498 (N_18498,N_17794,N_16525);
xnor U18499 (N_18499,N_17079,N_17285);
or U18500 (N_18500,N_17256,N_17808);
nor U18501 (N_18501,N_16788,N_17170);
nor U18502 (N_18502,N_16991,N_17748);
and U18503 (N_18503,N_17956,N_16499);
nor U18504 (N_18504,N_17334,N_16945);
nand U18505 (N_18505,N_17886,N_16508);
nand U18506 (N_18506,N_16842,N_16282);
xor U18507 (N_18507,N_17047,N_17667);
nand U18508 (N_18508,N_17261,N_17036);
or U18509 (N_18509,N_16484,N_17595);
or U18510 (N_18510,N_17414,N_17208);
nand U18511 (N_18511,N_17009,N_16530);
xnor U18512 (N_18512,N_16007,N_17866);
xnor U18513 (N_18513,N_17785,N_16494);
or U18514 (N_18514,N_16239,N_17890);
nor U18515 (N_18515,N_16586,N_17925);
xnor U18516 (N_18516,N_16137,N_16398);
nand U18517 (N_18517,N_17486,N_16870);
and U18518 (N_18518,N_17754,N_16534);
and U18519 (N_18519,N_17483,N_16108);
xnor U18520 (N_18520,N_17216,N_17924);
xor U18521 (N_18521,N_16521,N_17033);
and U18522 (N_18522,N_16819,N_16922);
xnor U18523 (N_18523,N_17221,N_16258);
nand U18524 (N_18524,N_16986,N_17042);
and U18525 (N_18525,N_16536,N_17061);
and U18526 (N_18526,N_17205,N_16849);
nand U18527 (N_18527,N_16545,N_16414);
xnor U18528 (N_18528,N_17836,N_17728);
and U18529 (N_18529,N_16331,N_16608);
xnor U18530 (N_18530,N_17513,N_16017);
or U18531 (N_18531,N_17599,N_16140);
or U18532 (N_18532,N_16700,N_17112);
nor U18533 (N_18533,N_16552,N_16565);
or U18534 (N_18534,N_16466,N_16228);
and U18535 (N_18535,N_17337,N_16419);
and U18536 (N_18536,N_17227,N_17594);
xnor U18537 (N_18537,N_16845,N_17763);
xor U18538 (N_18538,N_16439,N_17132);
and U18539 (N_18539,N_17625,N_17803);
nand U18540 (N_18540,N_16120,N_17680);
nand U18541 (N_18541,N_17692,N_16689);
and U18542 (N_18542,N_17262,N_17917);
and U18543 (N_18543,N_16672,N_16316);
nor U18544 (N_18544,N_17485,N_17269);
nor U18545 (N_18545,N_16032,N_17970);
xnor U18546 (N_18546,N_16663,N_17145);
and U18547 (N_18547,N_16944,N_17016);
and U18548 (N_18548,N_16431,N_16043);
xnor U18549 (N_18549,N_16884,N_17537);
or U18550 (N_18550,N_16385,N_16880);
or U18551 (N_18551,N_17735,N_16052);
xor U18552 (N_18552,N_16741,N_17394);
and U18553 (N_18553,N_16334,N_16726);
nand U18554 (N_18554,N_16445,N_17078);
nor U18555 (N_18555,N_16474,N_17458);
xnor U18556 (N_18556,N_16190,N_17200);
and U18557 (N_18557,N_17971,N_17233);
or U18558 (N_18558,N_16549,N_16600);
nor U18559 (N_18559,N_17427,N_17492);
and U18560 (N_18560,N_16749,N_16336);
xnor U18561 (N_18561,N_16274,N_16974);
xor U18562 (N_18562,N_16847,N_16138);
nor U18563 (N_18563,N_17077,N_17514);
xor U18564 (N_18564,N_16226,N_17961);
and U18565 (N_18565,N_17875,N_17454);
and U18566 (N_18566,N_16089,N_16139);
nor U18567 (N_18567,N_16009,N_17868);
or U18568 (N_18568,N_17039,N_17818);
or U18569 (N_18569,N_17129,N_17616);
and U18570 (N_18570,N_16272,N_16724);
or U18571 (N_18571,N_17349,N_17953);
or U18572 (N_18572,N_16584,N_16738);
xor U18573 (N_18573,N_16725,N_16803);
nand U18574 (N_18574,N_17296,N_17374);
nand U18575 (N_18575,N_17432,N_16718);
nand U18576 (N_18576,N_17673,N_16527);
nor U18577 (N_18577,N_16400,N_17561);
nand U18578 (N_18578,N_16252,N_17215);
or U18579 (N_18579,N_16812,N_16493);
or U18580 (N_18580,N_16815,N_17702);
or U18581 (N_18581,N_17303,N_16074);
nand U18582 (N_18582,N_16670,N_16250);
or U18583 (N_18583,N_16208,N_16701);
xor U18584 (N_18584,N_17165,N_16921);
nand U18585 (N_18585,N_17716,N_17187);
nand U18586 (N_18586,N_17697,N_16180);
nor U18587 (N_18587,N_17280,N_17873);
xnor U18588 (N_18588,N_16284,N_17849);
and U18589 (N_18589,N_16498,N_16654);
nor U18590 (N_18590,N_16635,N_16393);
and U18591 (N_18591,N_16542,N_17975);
nor U18592 (N_18592,N_17210,N_16130);
nand U18593 (N_18593,N_17869,N_16178);
or U18594 (N_18594,N_17272,N_16966);
or U18595 (N_18595,N_17572,N_17484);
and U18596 (N_18596,N_17711,N_17172);
or U18597 (N_18597,N_17951,N_16125);
nand U18598 (N_18598,N_16488,N_17264);
or U18599 (N_18599,N_17002,N_16675);
and U18600 (N_18600,N_16893,N_17095);
xnor U18601 (N_18601,N_16739,N_16390);
and U18602 (N_18602,N_16998,N_17636);
and U18603 (N_18603,N_17275,N_16963);
nand U18604 (N_18604,N_16246,N_17220);
xor U18605 (N_18605,N_17742,N_17573);
nor U18606 (N_18606,N_17041,N_17253);
nand U18607 (N_18607,N_16482,N_17102);
nor U18608 (N_18608,N_16034,N_16896);
and U18609 (N_18609,N_16193,N_17551);
nand U18610 (N_18610,N_16869,N_16073);
xor U18611 (N_18611,N_16270,N_17406);
nor U18612 (N_18612,N_16954,N_16413);
nand U18613 (N_18613,N_16984,N_16967);
nand U18614 (N_18614,N_16573,N_16801);
xor U18615 (N_18615,N_16914,N_17950);
and U18616 (N_18616,N_17771,N_16371);
xnor U18617 (N_18617,N_17245,N_16913);
xnor U18618 (N_18618,N_17896,N_16850);
nand U18619 (N_18619,N_16677,N_17018);
and U18620 (N_18620,N_16318,N_17783);
xor U18621 (N_18621,N_16567,N_17423);
or U18622 (N_18622,N_16609,N_17948);
or U18623 (N_18623,N_17094,N_16621);
nand U18624 (N_18624,N_17389,N_16866);
nand U18625 (N_18625,N_17503,N_16942);
or U18626 (N_18626,N_16477,N_17559);
and U18627 (N_18627,N_17254,N_17359);
and U18628 (N_18628,N_17306,N_17740);
nand U18629 (N_18629,N_17447,N_17798);
xnor U18630 (N_18630,N_17652,N_16507);
nor U18631 (N_18631,N_17466,N_16538);
nand U18632 (N_18632,N_16753,N_16580);
nand U18633 (N_18633,N_16590,N_16768);
nand U18634 (N_18634,N_16298,N_17646);
and U18635 (N_18635,N_17010,N_16930);
nor U18636 (N_18636,N_16579,N_17224);
or U18637 (N_18637,N_16540,N_17250);
or U18638 (N_18638,N_16195,N_16854);
xor U18639 (N_18639,N_17151,N_17892);
nand U18640 (N_18640,N_17428,N_16346);
nor U18641 (N_18641,N_17494,N_17547);
nand U18642 (N_18642,N_16325,N_16691);
xor U18643 (N_18643,N_17407,N_17614);
xor U18644 (N_18644,N_16086,N_17054);
nand U18645 (N_18645,N_17106,N_16173);
and U18646 (N_18646,N_16105,N_17930);
and U18647 (N_18647,N_16262,N_16666);
or U18648 (N_18648,N_16018,N_17028);
or U18649 (N_18649,N_16209,N_17152);
or U18650 (N_18650,N_16548,N_16559);
xor U18651 (N_18651,N_17856,N_16287);
xor U18652 (N_18652,N_17048,N_16592);
or U18653 (N_18653,N_16721,N_17281);
xnor U18654 (N_18654,N_16091,N_16397);
nor U18655 (N_18655,N_17710,N_16708);
nand U18656 (N_18656,N_17081,N_16200);
xnor U18657 (N_18657,N_16010,N_16081);
xnor U18658 (N_18658,N_17070,N_17995);
and U18659 (N_18659,N_17082,N_17465);
xnor U18660 (N_18660,N_16172,N_16170);
xor U18661 (N_18661,N_17356,N_17940);
or U18662 (N_18662,N_16581,N_17014);
nand U18663 (N_18663,N_16123,N_17938);
xnor U18664 (N_18664,N_17188,N_16657);
and U18665 (N_18665,N_17321,N_16817);
or U18666 (N_18666,N_16483,N_16370);
nand U18667 (N_18667,N_17985,N_17905);
or U18668 (N_18668,N_17679,N_16837);
or U18669 (N_18669,N_17440,N_17519);
and U18670 (N_18670,N_17606,N_16163);
xor U18671 (N_18671,N_17801,N_16337);
nand U18672 (N_18672,N_16408,N_17615);
xnor U18673 (N_18673,N_17746,N_16699);
nor U18674 (N_18674,N_16285,N_16630);
and U18675 (N_18675,N_17093,N_17453);
xnor U18676 (N_18676,N_16421,N_17468);
xor U18677 (N_18677,N_17967,N_16327);
or U18678 (N_18678,N_16716,N_16624);
and U18679 (N_18679,N_16134,N_17051);
nor U18680 (N_18680,N_17304,N_16066);
nor U18681 (N_18681,N_17238,N_16029);
or U18682 (N_18682,N_17964,N_16912);
nand U18683 (N_18683,N_16526,N_16765);
xor U18684 (N_18684,N_17604,N_17329);
and U18685 (N_18685,N_17375,N_17497);
nor U18686 (N_18686,N_17758,N_16919);
nand U18687 (N_18687,N_17131,N_17168);
and U18688 (N_18688,N_17587,N_17089);
nand U18689 (N_18689,N_16039,N_16612);
and U18690 (N_18690,N_16149,N_17130);
nand U18691 (N_18691,N_17538,N_16339);
and U18692 (N_18692,N_16299,N_16838);
and U18693 (N_18693,N_17086,N_17955);
and U18694 (N_18694,N_17361,N_17314);
nand U18695 (N_18695,N_16362,N_17828);
or U18696 (N_18696,N_16723,N_16802);
or U18697 (N_18697,N_16044,N_17883);
or U18698 (N_18698,N_16269,N_16183);
or U18699 (N_18699,N_16242,N_17838);
nand U18700 (N_18700,N_16637,N_16793);
xnor U18701 (N_18701,N_16087,N_17781);
and U18702 (N_18702,N_16826,N_17283);
xnor U18703 (N_18703,N_16341,N_17267);
and U18704 (N_18704,N_16351,N_17617);
xnor U18705 (N_18705,N_16159,N_16035);
and U18706 (N_18706,N_16830,N_16214);
nand U18707 (N_18707,N_16879,N_16873);
nand U18708 (N_18708,N_17155,N_17319);
nand U18709 (N_18709,N_17906,N_16461);
nor U18710 (N_18710,N_16391,N_16229);
xor U18711 (N_18711,N_17888,N_17566);
or U18712 (N_18712,N_16948,N_17597);
nand U18713 (N_18713,N_16629,N_17308);
nor U18714 (N_18714,N_17363,N_17885);
xor U18715 (N_18715,N_16472,N_17881);
nor U18716 (N_18716,N_17479,N_17487);
nor U18717 (N_18717,N_17920,N_17045);
xnor U18718 (N_18718,N_16951,N_17396);
or U18719 (N_18719,N_17859,N_16692);
nand U18720 (N_18720,N_17362,N_16636);
xnor U18721 (N_18721,N_16372,N_16184);
nand U18722 (N_18722,N_16113,N_16959);
nand U18723 (N_18723,N_16626,N_16187);
nor U18724 (N_18724,N_16785,N_17105);
and U18725 (N_18725,N_17700,N_17806);
and U18726 (N_18726,N_17660,N_17505);
xnor U18727 (N_18727,N_16783,N_17664);
nor U18728 (N_18728,N_17183,N_16244);
xnor U18729 (N_18729,N_17982,N_16503);
nand U18730 (N_18730,N_16040,N_16639);
and U18731 (N_18731,N_17438,N_16569);
nor U18732 (N_18732,N_17325,N_16977);
or U18733 (N_18733,N_17629,N_16575);
nand U18734 (N_18734,N_16306,N_17266);
nand U18735 (N_18735,N_16056,N_16563);
xnor U18736 (N_18736,N_17581,N_16354);
or U18737 (N_18737,N_17932,N_17478);
or U18738 (N_18738,N_17983,N_16558);
nand U18739 (N_18739,N_17154,N_16756);
or U18740 (N_18740,N_16221,N_17739);
and U18741 (N_18741,N_16577,N_17518);
nand U18742 (N_18742,N_17911,N_17623);
nor U18743 (N_18743,N_16647,N_16970);
and U18744 (N_18744,N_17598,N_16980);
nand U18745 (N_18745,N_17004,N_17162);
nand U18746 (N_18746,N_17326,N_16632);
xor U18747 (N_18747,N_16887,N_17752);
and U18748 (N_18748,N_16141,N_16253);
nor U18749 (N_18749,N_16167,N_17481);
xnor U18750 (N_18750,N_17339,N_17974);
nor U18751 (N_18751,N_17842,N_17288);
nand U18752 (N_18752,N_17860,N_16500);
nand U18753 (N_18753,N_17820,N_17258);
and U18754 (N_18754,N_16656,N_16684);
or U18755 (N_18755,N_16451,N_17234);
nor U18756 (N_18756,N_17817,N_16717);
xor U18757 (N_18757,N_17841,N_16080);
or U18758 (N_18758,N_16377,N_17668);
and U18759 (N_18759,N_17067,N_17577);
nand U18760 (N_18760,N_16042,N_16122);
xnor U18761 (N_18761,N_16789,N_16553);
or U18762 (N_18762,N_16328,N_17324);
nor U18763 (N_18763,N_16729,N_16935);
or U18764 (N_18764,N_16952,N_17934);
nor U18765 (N_18765,N_16512,N_16928);
and U18766 (N_18766,N_16537,N_17651);
nand U18767 (N_18767,N_17243,N_17019);
nand U18768 (N_18768,N_16340,N_17958);
nor U18769 (N_18769,N_17056,N_16225);
nand U18770 (N_18770,N_16813,N_17295);
nand U18771 (N_18771,N_16008,N_17921);
nor U18772 (N_18772,N_16641,N_16084);
nand U18773 (N_18773,N_17683,N_16077);
or U18774 (N_18774,N_17643,N_16894);
nand U18775 (N_18775,N_17399,N_17813);
or U18776 (N_18776,N_16965,N_17912);
nor U18777 (N_18777,N_17825,N_16883);
nor U18778 (N_18778,N_17265,N_17737);
nand U18779 (N_18779,N_16628,N_17580);
or U18780 (N_18780,N_17557,N_16343);
nand U18781 (N_18781,N_16469,N_16059);
xor U18782 (N_18782,N_17864,N_17023);
nand U18783 (N_18783,N_17997,N_17190);
nor U18784 (N_18784,N_17402,N_17249);
xnor U18785 (N_18785,N_17475,N_16367);
and U18786 (N_18786,N_17108,N_17550);
nor U18787 (N_18787,N_17861,N_16396);
xnor U18788 (N_18788,N_17302,N_17952);
xnor U18789 (N_18789,N_16737,N_17219);
nand U18790 (N_18790,N_16902,N_16355);
and U18791 (N_18791,N_16247,N_17867);
or U18792 (N_18792,N_16611,N_17346);
and U18793 (N_18793,N_17133,N_16240);
nor U18794 (N_18794,N_17672,N_16909);
or U18795 (N_18795,N_17202,N_16697);
or U18796 (N_18796,N_17135,N_17586);
xor U18797 (N_18797,N_17960,N_16746);
or U18798 (N_18798,N_16886,N_16520);
nand U18799 (N_18799,N_16671,N_17383);
xor U18800 (N_18800,N_17928,N_17292);
or U18801 (N_18801,N_17793,N_16311);
and U18802 (N_18802,N_16063,N_16818);
xor U18803 (N_18803,N_17178,N_17546);
or U18804 (N_18804,N_17919,N_16186);
or U18805 (N_18805,N_16416,N_17217);
nor U18806 (N_18806,N_17690,N_17840);
nand U18807 (N_18807,N_16568,N_17558);
nor U18808 (N_18808,N_17830,N_16731);
nor U18809 (N_18809,N_17046,N_17229);
and U18810 (N_18810,N_16047,N_17533);
nor U18811 (N_18811,N_17520,N_16888);
and U18812 (N_18812,N_16188,N_17585);
xnor U18813 (N_18813,N_16000,N_17678);
or U18814 (N_18814,N_16317,N_17732);
and U18815 (N_18815,N_16779,N_16769);
nand U18816 (N_18816,N_17114,N_17755);
xnor U18817 (N_18817,N_16016,N_16444);
xor U18818 (N_18818,N_16365,N_16437);
or U18819 (N_18819,N_17640,N_17148);
and U18820 (N_18820,N_17966,N_17143);
nand U18821 (N_18821,N_16703,N_17554);
nand U18822 (N_18822,N_16295,N_16249);
nand U18823 (N_18823,N_17874,N_16300);
nand U18824 (N_18824,N_17029,N_16263);
or U18825 (N_18825,N_17175,N_16961);
nor U18826 (N_18826,N_17695,N_17405);
or U18827 (N_18827,N_16111,N_16182);
or U18828 (N_18828,N_17589,N_17286);
nand U18829 (N_18829,N_17057,N_17176);
or U18830 (N_18830,N_17691,N_17260);
xor U18831 (N_18831,N_17309,N_17731);
xnor U18832 (N_18832,N_17845,N_16366);
nor U18833 (N_18833,N_16747,N_16904);
xnor U18834 (N_18834,N_16652,N_16876);
xor U18835 (N_18835,N_17622,N_17008);
and U18836 (N_18836,N_17255,N_16759);
and U18837 (N_18837,N_16291,N_16727);
and U18838 (N_18838,N_17480,N_16205);
and U18839 (N_18839,N_16076,N_17064);
nor U18840 (N_18840,N_16811,N_16199);
and U18841 (N_18841,N_17988,N_16481);
and U18842 (N_18842,N_16949,N_17522);
and U18843 (N_18843,N_17499,N_17058);
and U18844 (N_18844,N_16347,N_16861);
xor U18845 (N_18845,N_17305,N_17772);
nor U18846 (N_18846,N_16358,N_17900);
nor U18847 (N_18847,N_17768,N_16426);
nand U18848 (N_18848,N_16234,N_16215);
xor U18849 (N_18849,N_16659,N_17571);
nand U18850 (N_18850,N_17831,N_16787);
nor U18851 (N_18851,N_16290,N_16640);
or U18852 (N_18852,N_17827,N_17098);
nor U18853 (N_18853,N_17136,N_17111);
xnor U18854 (N_18854,N_17689,N_16582);
nand U18855 (N_18855,N_16082,N_16320);
nand U18856 (N_18856,N_16402,N_16101);
nand U18857 (N_18857,N_17898,N_16858);
xnor U18858 (N_18858,N_17922,N_17544);
or U18859 (N_18859,N_17863,N_16011);
and U18860 (N_18860,N_17290,N_17789);
or U18861 (N_18861,N_16479,N_16288);
xor U18862 (N_18862,N_16156,N_16429);
and U18863 (N_18863,N_16937,N_16766);
or U18864 (N_18864,N_17762,N_16771);
or U18865 (N_18865,N_17270,N_17540);
xor U18866 (N_18866,N_16062,N_16462);
xnor U18867 (N_18867,N_17460,N_16694);
nand U18868 (N_18868,N_17562,N_17189);
or U18869 (N_18869,N_16799,N_17024);
nor U18870 (N_18870,N_17171,N_17287);
nor U18871 (N_18871,N_17507,N_17954);
xor U18872 (N_18872,N_16104,N_17344);
or U18873 (N_18873,N_16491,N_16550);
nand U18874 (N_18874,N_17068,N_17201);
xnor U18875 (N_18875,N_17722,N_17213);
nand U18876 (N_18876,N_17962,N_16094);
xor U18877 (N_18877,N_17777,N_16411);
or U18878 (N_18878,N_16993,N_17137);
xor U18879 (N_18879,N_17819,N_16687);
or U18880 (N_18880,N_16321,N_16384);
and U18881 (N_18881,N_17593,N_16041);
or U18882 (N_18882,N_17477,N_16458);
nand U18883 (N_18883,N_17409,N_17980);
xor U18884 (N_18884,N_17609,N_16560);
xnor U18885 (N_18885,N_17293,N_17979);
and U18886 (N_18886,N_16650,N_17969);
nand U18887 (N_18887,N_17655,N_17613);
and U18888 (N_18888,N_17981,N_17545);
and U18889 (N_18889,N_17631,N_16502);
xnor U18890 (N_18890,N_17749,N_16051);
nand U18891 (N_18891,N_17496,N_16661);
nor U18892 (N_18892,N_16096,N_17725);
or U18893 (N_18893,N_16864,N_16168);
nor U18894 (N_18894,N_17592,N_16605);
nand U18895 (N_18895,N_16420,N_16088);
xor U18896 (N_18896,N_16532,N_16294);
nor U18897 (N_18897,N_17439,N_16133);
nand U18898 (N_18898,N_16266,N_17435);
and U18899 (N_18899,N_16588,N_17619);
nor U18900 (N_18900,N_17193,N_16430);
nand U18901 (N_18901,N_17268,N_16227);
and U18902 (N_18902,N_17035,N_16969);
xnor U18903 (N_18903,N_17976,N_17937);
xor U18904 (N_18904,N_16315,N_17388);
xor U18905 (N_18905,N_17532,N_16770);
nand U18906 (N_18906,N_17770,N_16707);
and U18907 (N_18907,N_16369,N_17139);
nor U18908 (N_18908,N_17812,N_16905);
xor U18909 (N_18909,N_17779,N_17676);
nand U18910 (N_18910,N_17336,N_16015);
nand U18911 (N_18911,N_17134,N_17624);
and U18912 (N_18912,N_16996,N_17161);
or U18913 (N_18913,N_16832,N_17381);
xnor U18914 (N_18914,N_17127,N_17929);
nor U18915 (N_18915,N_17191,N_16119);
and U18916 (N_18916,N_16523,N_17222);
xnor U18917 (N_18917,N_16906,N_16602);
or U18918 (N_18918,N_17412,N_17575);
xnor U18919 (N_18919,N_17627,N_17350);
xnor U18920 (N_18920,N_16620,N_17124);
nor U18921 (N_18921,N_16233,N_16165);
xnor U18922 (N_18922,N_16363,N_16455);
or U18923 (N_18923,N_17907,N_17126);
nand U18924 (N_18924,N_16546,N_16181);
xnor U18925 (N_18925,N_17535,N_16148);
and U18926 (N_18926,N_16264,N_16102);
xnor U18927 (N_18927,N_17502,N_17476);
nor U18928 (N_18928,N_17526,N_17747);
or U18929 (N_18929,N_16927,N_17611);
and U18930 (N_18930,N_17273,N_16114);
nand U18931 (N_18931,N_17723,N_17020);
xnor U18932 (N_18932,N_16286,N_17391);
nand U18933 (N_18933,N_16990,N_17449);
nand U18934 (N_18934,N_17765,N_16871);
xor U18935 (N_18935,N_16103,N_16394);
or U18936 (N_18936,N_17397,N_16348);
xnor U18937 (N_18937,N_16448,N_16330);
nor U18938 (N_18938,N_16322,N_16825);
nand U18939 (N_18939,N_17904,N_16425);
xnor U18940 (N_18940,N_17791,N_17521);
xnor U18941 (N_18941,N_17569,N_16762);
and U18942 (N_18942,N_16576,N_16820);
or U18943 (N_18943,N_16135,N_17991);
nor U18944 (N_18944,N_17936,N_17659);
and U18945 (N_18945,N_16736,N_17759);
xor U18946 (N_18946,N_17037,N_17181);
xor U18947 (N_18947,N_16557,N_16132);
and U18948 (N_18948,N_16698,N_17506);
nor U18949 (N_18949,N_17786,N_17467);
nand U18950 (N_18950,N_16597,N_17052);
nor U18951 (N_18951,N_17712,N_16846);
or U18952 (N_18952,N_16496,N_16973);
or U18953 (N_18953,N_16923,N_17542);
nand U18954 (N_18954,N_16301,N_17650);
xnor U18955 (N_18955,N_17444,N_16517);
and U18956 (N_18956,N_16901,N_16983);
or U18957 (N_18957,N_16742,N_17425);
nor U18958 (N_18958,N_17100,N_16667);
nor U18959 (N_18959,N_16124,N_17101);
or U18960 (N_18960,N_16947,N_16012);
xor U18961 (N_18961,N_17852,N_17529);
or U18962 (N_18962,N_16230,N_16964);
nor U18963 (N_18963,N_16231,N_17385);
and U18964 (N_18964,N_16763,N_17853);
nand U18965 (N_18965,N_17761,N_17446);
and U18966 (N_18966,N_17110,N_16616);
nor U18967 (N_18967,N_17844,N_16578);
nand U18968 (N_18968,N_16349,N_17122);
nor U18969 (N_18969,N_17338,N_16733);
or U18970 (N_18970,N_17463,N_16660);
or U18971 (N_18971,N_17006,N_16556);
nand U18972 (N_18972,N_16678,N_17491);
nand U18973 (N_18973,N_16821,N_17835);
and U18974 (N_18974,N_16364,N_17376);
nand U18975 (N_18975,N_17915,N_17003);
or U18976 (N_18976,N_16189,N_16174);
or U18977 (N_18977,N_16690,N_16979);
xnor U18978 (N_18978,N_17804,N_16150);
nand U18979 (N_18979,N_16856,N_17973);
and U18980 (N_18980,N_16613,N_17944);
or U18981 (N_18981,N_17096,N_16169);
xnor U18982 (N_18982,N_17276,N_17166);
or U18983 (N_18983,N_17158,N_17515);
nor U18984 (N_18984,N_17473,N_17116);
or U18985 (N_18985,N_17118,N_16127);
or U18986 (N_18986,N_16511,N_17066);
nor U18987 (N_18987,N_16026,N_17994);
or U18988 (N_18988,N_17647,N_17784);
nand U18989 (N_18989,N_17993,N_17899);
nor U18990 (N_18990,N_17410,N_17807);
or U18991 (N_18991,N_17694,N_16764);
nor U18992 (N_18992,N_17750,N_17837);
xnor U18993 (N_18993,N_16037,N_17044);
nand U18994 (N_18994,N_16751,N_17662);
nor U18995 (N_18995,N_17332,N_16389);
nand U18996 (N_18996,N_16754,N_17099);
or U18997 (N_18997,N_16574,N_16623);
nor U18998 (N_18998,N_17080,N_16618);
xnor U18999 (N_18999,N_17104,N_16786);
and U19000 (N_19000,N_17167,N_16587);
or U19001 (N_19001,N_16308,N_16174);
xnor U19002 (N_19002,N_17777,N_17022);
and U19003 (N_19003,N_16633,N_17718);
and U19004 (N_19004,N_16707,N_16381);
and U19005 (N_19005,N_16449,N_17744);
xor U19006 (N_19006,N_17054,N_16890);
nor U19007 (N_19007,N_16720,N_16770);
and U19008 (N_19008,N_17941,N_17471);
xor U19009 (N_19009,N_17441,N_16764);
xor U19010 (N_19010,N_17545,N_16558);
nand U19011 (N_19011,N_16557,N_17642);
or U19012 (N_19012,N_17864,N_17878);
nand U19013 (N_19013,N_17920,N_16739);
nand U19014 (N_19014,N_16978,N_16355);
and U19015 (N_19015,N_17739,N_17212);
and U19016 (N_19016,N_17125,N_16765);
xor U19017 (N_19017,N_16440,N_17921);
or U19018 (N_19018,N_16622,N_16840);
nor U19019 (N_19019,N_17272,N_16675);
nor U19020 (N_19020,N_17920,N_16204);
nand U19021 (N_19021,N_17039,N_16108);
nand U19022 (N_19022,N_17970,N_16651);
xor U19023 (N_19023,N_16138,N_16144);
xor U19024 (N_19024,N_17112,N_16317);
nand U19025 (N_19025,N_17735,N_16542);
nor U19026 (N_19026,N_16147,N_16539);
or U19027 (N_19027,N_17861,N_16748);
nand U19028 (N_19028,N_16528,N_17100);
or U19029 (N_19029,N_17603,N_17109);
xnor U19030 (N_19030,N_17233,N_17880);
xor U19031 (N_19031,N_16592,N_17832);
or U19032 (N_19032,N_17562,N_16943);
xnor U19033 (N_19033,N_16925,N_16672);
nand U19034 (N_19034,N_17800,N_17449);
nor U19035 (N_19035,N_17576,N_16939);
and U19036 (N_19036,N_16732,N_17817);
xor U19037 (N_19037,N_17070,N_17504);
and U19038 (N_19038,N_17179,N_17857);
nor U19039 (N_19039,N_17118,N_16873);
xnor U19040 (N_19040,N_16238,N_17007);
nor U19041 (N_19041,N_16763,N_16123);
xnor U19042 (N_19042,N_16987,N_16591);
nor U19043 (N_19043,N_17505,N_17435);
nor U19044 (N_19044,N_17258,N_16925);
nand U19045 (N_19045,N_16459,N_17146);
nor U19046 (N_19046,N_16179,N_17609);
and U19047 (N_19047,N_17945,N_17802);
and U19048 (N_19048,N_17562,N_16112);
xor U19049 (N_19049,N_16468,N_17727);
or U19050 (N_19050,N_16237,N_17739);
nor U19051 (N_19051,N_16464,N_17789);
xnor U19052 (N_19052,N_16319,N_17891);
nand U19053 (N_19053,N_16403,N_16597);
nor U19054 (N_19054,N_16790,N_17310);
xor U19055 (N_19055,N_17482,N_16226);
or U19056 (N_19056,N_16528,N_16941);
and U19057 (N_19057,N_16236,N_17384);
and U19058 (N_19058,N_16607,N_16264);
and U19059 (N_19059,N_16337,N_16986);
nor U19060 (N_19060,N_16347,N_16978);
nor U19061 (N_19061,N_17291,N_17504);
and U19062 (N_19062,N_16296,N_17481);
and U19063 (N_19063,N_16037,N_17939);
xor U19064 (N_19064,N_16411,N_16625);
and U19065 (N_19065,N_17991,N_17208);
xor U19066 (N_19066,N_17729,N_16282);
nand U19067 (N_19067,N_17096,N_16485);
or U19068 (N_19068,N_16613,N_17791);
xnor U19069 (N_19069,N_17259,N_17757);
and U19070 (N_19070,N_17536,N_17846);
xnor U19071 (N_19071,N_17591,N_17876);
nor U19072 (N_19072,N_17848,N_17807);
or U19073 (N_19073,N_17647,N_16984);
and U19074 (N_19074,N_16124,N_16897);
or U19075 (N_19075,N_17068,N_17006);
or U19076 (N_19076,N_17810,N_16009);
and U19077 (N_19077,N_16936,N_16310);
xor U19078 (N_19078,N_16602,N_17212);
nand U19079 (N_19079,N_17105,N_16072);
or U19080 (N_19080,N_16804,N_16154);
nor U19081 (N_19081,N_16532,N_17297);
xor U19082 (N_19082,N_16293,N_17984);
and U19083 (N_19083,N_17404,N_17950);
nand U19084 (N_19084,N_16584,N_16090);
nor U19085 (N_19085,N_17871,N_17057);
and U19086 (N_19086,N_16864,N_17332);
or U19087 (N_19087,N_17625,N_17042);
nand U19088 (N_19088,N_16671,N_16704);
xor U19089 (N_19089,N_17046,N_17817);
nor U19090 (N_19090,N_16837,N_17704);
nand U19091 (N_19091,N_16678,N_17679);
or U19092 (N_19092,N_16372,N_16239);
nand U19093 (N_19093,N_17056,N_17124);
nand U19094 (N_19094,N_17198,N_16144);
nand U19095 (N_19095,N_16227,N_17843);
xor U19096 (N_19096,N_16524,N_16599);
nor U19097 (N_19097,N_16115,N_16760);
xnor U19098 (N_19098,N_16346,N_17322);
nand U19099 (N_19099,N_16776,N_16301);
or U19100 (N_19100,N_16809,N_16417);
nor U19101 (N_19101,N_17601,N_17846);
xnor U19102 (N_19102,N_16605,N_17123);
or U19103 (N_19103,N_16501,N_16248);
nand U19104 (N_19104,N_16780,N_17873);
nor U19105 (N_19105,N_17390,N_17388);
xnor U19106 (N_19106,N_17949,N_17335);
xor U19107 (N_19107,N_16594,N_16269);
or U19108 (N_19108,N_17449,N_16682);
or U19109 (N_19109,N_16056,N_16080);
and U19110 (N_19110,N_17093,N_17043);
and U19111 (N_19111,N_17645,N_16936);
and U19112 (N_19112,N_16827,N_16791);
xnor U19113 (N_19113,N_16626,N_17220);
and U19114 (N_19114,N_17690,N_17181);
nand U19115 (N_19115,N_17536,N_17919);
nand U19116 (N_19116,N_16619,N_17010);
or U19117 (N_19117,N_16747,N_16836);
xnor U19118 (N_19118,N_16553,N_17996);
xnor U19119 (N_19119,N_16881,N_16593);
and U19120 (N_19120,N_17769,N_16502);
nand U19121 (N_19121,N_16017,N_16705);
xnor U19122 (N_19122,N_16514,N_17102);
xor U19123 (N_19123,N_17779,N_17796);
nor U19124 (N_19124,N_16780,N_17200);
nand U19125 (N_19125,N_17085,N_16640);
nor U19126 (N_19126,N_16337,N_17896);
and U19127 (N_19127,N_17863,N_17488);
xnor U19128 (N_19128,N_17293,N_16509);
nand U19129 (N_19129,N_17762,N_17654);
and U19130 (N_19130,N_17907,N_16332);
nor U19131 (N_19131,N_17941,N_16940);
nor U19132 (N_19132,N_16216,N_17390);
nor U19133 (N_19133,N_17226,N_16517);
xnor U19134 (N_19134,N_16249,N_17615);
or U19135 (N_19135,N_16682,N_16953);
and U19136 (N_19136,N_17234,N_16651);
nand U19137 (N_19137,N_16636,N_17602);
and U19138 (N_19138,N_17724,N_17406);
nor U19139 (N_19139,N_17081,N_17430);
nand U19140 (N_19140,N_17401,N_17305);
xnor U19141 (N_19141,N_16788,N_16009);
nor U19142 (N_19142,N_16916,N_16001);
nand U19143 (N_19143,N_16947,N_16451);
nor U19144 (N_19144,N_16503,N_17091);
and U19145 (N_19145,N_17742,N_17231);
nor U19146 (N_19146,N_16968,N_16202);
xor U19147 (N_19147,N_16204,N_16427);
nand U19148 (N_19148,N_16526,N_17055);
nor U19149 (N_19149,N_17871,N_16439);
xor U19150 (N_19150,N_17482,N_17615);
and U19151 (N_19151,N_17990,N_16198);
nand U19152 (N_19152,N_16651,N_16091);
nor U19153 (N_19153,N_16824,N_17924);
xnor U19154 (N_19154,N_16701,N_17824);
nand U19155 (N_19155,N_17071,N_17736);
or U19156 (N_19156,N_17889,N_16395);
xnor U19157 (N_19157,N_16119,N_17475);
or U19158 (N_19158,N_17433,N_17980);
nor U19159 (N_19159,N_17068,N_17298);
nor U19160 (N_19160,N_17383,N_17887);
nor U19161 (N_19161,N_17052,N_17981);
and U19162 (N_19162,N_17710,N_16375);
nor U19163 (N_19163,N_16425,N_17686);
and U19164 (N_19164,N_17778,N_16508);
xnor U19165 (N_19165,N_16094,N_16483);
xnor U19166 (N_19166,N_17973,N_17797);
xor U19167 (N_19167,N_17882,N_17020);
xnor U19168 (N_19168,N_16247,N_16799);
and U19169 (N_19169,N_17740,N_17174);
nand U19170 (N_19170,N_17929,N_16861);
nor U19171 (N_19171,N_16706,N_16695);
nand U19172 (N_19172,N_17093,N_17793);
xor U19173 (N_19173,N_16080,N_16546);
and U19174 (N_19174,N_17182,N_17563);
and U19175 (N_19175,N_16065,N_16840);
and U19176 (N_19176,N_17972,N_16615);
nor U19177 (N_19177,N_16523,N_16351);
nand U19178 (N_19178,N_17747,N_16512);
nand U19179 (N_19179,N_16348,N_17452);
and U19180 (N_19180,N_17127,N_17627);
or U19181 (N_19181,N_17494,N_17735);
nand U19182 (N_19182,N_16463,N_17934);
or U19183 (N_19183,N_17371,N_17086);
xor U19184 (N_19184,N_16413,N_17161);
xnor U19185 (N_19185,N_17964,N_17722);
or U19186 (N_19186,N_16272,N_17298);
nor U19187 (N_19187,N_17625,N_17565);
xor U19188 (N_19188,N_17438,N_16853);
or U19189 (N_19189,N_16630,N_17154);
nor U19190 (N_19190,N_17321,N_16132);
nand U19191 (N_19191,N_17063,N_17413);
and U19192 (N_19192,N_16444,N_17906);
or U19193 (N_19193,N_16187,N_17848);
or U19194 (N_19194,N_17827,N_17089);
or U19195 (N_19195,N_16406,N_16313);
and U19196 (N_19196,N_16403,N_17057);
nor U19197 (N_19197,N_17231,N_17884);
xor U19198 (N_19198,N_17882,N_16834);
and U19199 (N_19199,N_16979,N_17273);
nand U19200 (N_19200,N_16675,N_17268);
and U19201 (N_19201,N_16479,N_16255);
or U19202 (N_19202,N_17109,N_16660);
nor U19203 (N_19203,N_16695,N_16423);
or U19204 (N_19204,N_16534,N_17396);
or U19205 (N_19205,N_17833,N_17209);
nor U19206 (N_19206,N_17002,N_17530);
nor U19207 (N_19207,N_16973,N_16759);
nand U19208 (N_19208,N_17045,N_16734);
or U19209 (N_19209,N_17890,N_17195);
nand U19210 (N_19210,N_16744,N_16112);
and U19211 (N_19211,N_17813,N_17608);
nor U19212 (N_19212,N_16825,N_16070);
nor U19213 (N_19213,N_17568,N_16201);
and U19214 (N_19214,N_17269,N_17140);
and U19215 (N_19215,N_17203,N_17290);
nor U19216 (N_19216,N_16062,N_17902);
nand U19217 (N_19217,N_16310,N_17927);
nor U19218 (N_19218,N_17274,N_16122);
xor U19219 (N_19219,N_17903,N_16388);
or U19220 (N_19220,N_17594,N_17146);
nand U19221 (N_19221,N_16122,N_17373);
xnor U19222 (N_19222,N_16334,N_17474);
nand U19223 (N_19223,N_17584,N_17379);
nand U19224 (N_19224,N_16531,N_16826);
nand U19225 (N_19225,N_16143,N_16603);
xor U19226 (N_19226,N_16368,N_16116);
or U19227 (N_19227,N_16867,N_16116);
xor U19228 (N_19228,N_17804,N_16172);
and U19229 (N_19229,N_16884,N_16005);
or U19230 (N_19230,N_17254,N_16654);
and U19231 (N_19231,N_16581,N_17556);
nor U19232 (N_19232,N_17378,N_16649);
nor U19233 (N_19233,N_16221,N_16679);
nor U19234 (N_19234,N_16676,N_16336);
nor U19235 (N_19235,N_17556,N_16643);
or U19236 (N_19236,N_16346,N_16747);
nor U19237 (N_19237,N_16396,N_17161);
or U19238 (N_19238,N_16460,N_16713);
nand U19239 (N_19239,N_17608,N_17126);
nor U19240 (N_19240,N_16050,N_17375);
and U19241 (N_19241,N_17693,N_17940);
and U19242 (N_19242,N_17039,N_16295);
and U19243 (N_19243,N_16210,N_17831);
nand U19244 (N_19244,N_16910,N_16160);
and U19245 (N_19245,N_16440,N_16712);
nor U19246 (N_19246,N_17620,N_17085);
xnor U19247 (N_19247,N_16276,N_17829);
and U19248 (N_19248,N_17914,N_16967);
xnor U19249 (N_19249,N_16889,N_17985);
or U19250 (N_19250,N_17668,N_17532);
nand U19251 (N_19251,N_16249,N_17192);
nand U19252 (N_19252,N_16728,N_17620);
nand U19253 (N_19253,N_16183,N_17356);
and U19254 (N_19254,N_16564,N_17501);
nor U19255 (N_19255,N_17986,N_16442);
nand U19256 (N_19256,N_16649,N_16348);
or U19257 (N_19257,N_17280,N_16918);
or U19258 (N_19258,N_16244,N_17475);
xnor U19259 (N_19259,N_16113,N_17288);
and U19260 (N_19260,N_17982,N_17740);
nor U19261 (N_19261,N_16516,N_17794);
or U19262 (N_19262,N_17501,N_17565);
nor U19263 (N_19263,N_17019,N_17609);
or U19264 (N_19264,N_17062,N_17416);
nand U19265 (N_19265,N_17837,N_16802);
xor U19266 (N_19266,N_16757,N_17092);
and U19267 (N_19267,N_16728,N_16766);
nor U19268 (N_19268,N_17595,N_17109);
nand U19269 (N_19269,N_16436,N_17380);
nand U19270 (N_19270,N_17963,N_17055);
or U19271 (N_19271,N_16179,N_17095);
xor U19272 (N_19272,N_17838,N_17943);
nand U19273 (N_19273,N_16982,N_17943);
and U19274 (N_19274,N_16515,N_17959);
xnor U19275 (N_19275,N_16196,N_16167);
xor U19276 (N_19276,N_16101,N_16965);
xnor U19277 (N_19277,N_17933,N_17085);
nor U19278 (N_19278,N_16983,N_16163);
xnor U19279 (N_19279,N_17222,N_17983);
and U19280 (N_19280,N_17884,N_17284);
xor U19281 (N_19281,N_17741,N_17363);
xnor U19282 (N_19282,N_17041,N_17576);
and U19283 (N_19283,N_17723,N_17195);
and U19284 (N_19284,N_16408,N_17917);
xnor U19285 (N_19285,N_16672,N_16668);
xor U19286 (N_19286,N_16864,N_16942);
or U19287 (N_19287,N_17094,N_17277);
xor U19288 (N_19288,N_16144,N_16608);
nor U19289 (N_19289,N_16883,N_16489);
nor U19290 (N_19290,N_16224,N_17191);
or U19291 (N_19291,N_16675,N_17916);
and U19292 (N_19292,N_16270,N_17934);
nor U19293 (N_19293,N_16443,N_16908);
or U19294 (N_19294,N_17169,N_17552);
nor U19295 (N_19295,N_17394,N_16479);
and U19296 (N_19296,N_17224,N_17992);
and U19297 (N_19297,N_17493,N_16715);
and U19298 (N_19298,N_16922,N_16195);
or U19299 (N_19299,N_17158,N_16128);
or U19300 (N_19300,N_17307,N_16875);
xor U19301 (N_19301,N_16373,N_16526);
nand U19302 (N_19302,N_16017,N_17161);
xor U19303 (N_19303,N_16943,N_16737);
and U19304 (N_19304,N_17858,N_16396);
xnor U19305 (N_19305,N_17968,N_17414);
xnor U19306 (N_19306,N_17869,N_17553);
nor U19307 (N_19307,N_16658,N_16347);
nor U19308 (N_19308,N_16326,N_17892);
xor U19309 (N_19309,N_17942,N_17063);
or U19310 (N_19310,N_16670,N_17068);
nor U19311 (N_19311,N_17424,N_17202);
and U19312 (N_19312,N_16632,N_17189);
nor U19313 (N_19313,N_17379,N_16493);
and U19314 (N_19314,N_16126,N_16031);
xor U19315 (N_19315,N_17193,N_16332);
and U19316 (N_19316,N_16705,N_16015);
nand U19317 (N_19317,N_16093,N_16507);
nand U19318 (N_19318,N_17990,N_17379);
xnor U19319 (N_19319,N_17713,N_16358);
nand U19320 (N_19320,N_17380,N_16416);
xnor U19321 (N_19321,N_16912,N_17307);
xnor U19322 (N_19322,N_16871,N_16801);
nand U19323 (N_19323,N_17807,N_17870);
xnor U19324 (N_19324,N_17583,N_16408);
and U19325 (N_19325,N_16171,N_17223);
or U19326 (N_19326,N_16358,N_17758);
and U19327 (N_19327,N_17530,N_17993);
or U19328 (N_19328,N_17547,N_16397);
nand U19329 (N_19329,N_16367,N_16317);
or U19330 (N_19330,N_16175,N_17958);
nand U19331 (N_19331,N_16169,N_17664);
nor U19332 (N_19332,N_16273,N_17996);
or U19333 (N_19333,N_16151,N_16651);
and U19334 (N_19334,N_17810,N_16164);
nand U19335 (N_19335,N_16552,N_16215);
and U19336 (N_19336,N_16232,N_17313);
or U19337 (N_19337,N_17981,N_16601);
xnor U19338 (N_19338,N_16602,N_17198);
nor U19339 (N_19339,N_17863,N_16333);
xor U19340 (N_19340,N_16520,N_16938);
nand U19341 (N_19341,N_17001,N_16178);
and U19342 (N_19342,N_16573,N_16313);
xor U19343 (N_19343,N_16252,N_16241);
xnor U19344 (N_19344,N_17233,N_16016);
and U19345 (N_19345,N_16183,N_17190);
nor U19346 (N_19346,N_17038,N_16609);
nor U19347 (N_19347,N_17946,N_17374);
xnor U19348 (N_19348,N_17801,N_17991);
and U19349 (N_19349,N_16776,N_16925);
nand U19350 (N_19350,N_17956,N_16486);
or U19351 (N_19351,N_16138,N_17373);
or U19352 (N_19352,N_16365,N_17722);
and U19353 (N_19353,N_16143,N_16540);
or U19354 (N_19354,N_17894,N_16323);
or U19355 (N_19355,N_17117,N_17676);
and U19356 (N_19356,N_17931,N_16769);
and U19357 (N_19357,N_16811,N_17614);
or U19358 (N_19358,N_17489,N_17815);
xor U19359 (N_19359,N_17018,N_16930);
or U19360 (N_19360,N_17070,N_17222);
xor U19361 (N_19361,N_17194,N_17722);
and U19362 (N_19362,N_17275,N_16705);
nor U19363 (N_19363,N_16089,N_16209);
xnor U19364 (N_19364,N_16736,N_16882);
nor U19365 (N_19365,N_17891,N_17449);
nand U19366 (N_19366,N_16591,N_17009);
nand U19367 (N_19367,N_16837,N_16925);
xnor U19368 (N_19368,N_16652,N_16364);
and U19369 (N_19369,N_16718,N_16898);
nand U19370 (N_19370,N_17145,N_16572);
and U19371 (N_19371,N_16349,N_17076);
or U19372 (N_19372,N_16558,N_16554);
or U19373 (N_19373,N_17876,N_17997);
xor U19374 (N_19374,N_16760,N_16465);
nand U19375 (N_19375,N_16957,N_16287);
or U19376 (N_19376,N_17006,N_17103);
xnor U19377 (N_19377,N_16868,N_16555);
xor U19378 (N_19378,N_16493,N_17645);
and U19379 (N_19379,N_17876,N_17211);
or U19380 (N_19380,N_16837,N_16713);
and U19381 (N_19381,N_16575,N_17901);
xnor U19382 (N_19382,N_16716,N_17267);
or U19383 (N_19383,N_17397,N_17669);
or U19384 (N_19384,N_16974,N_17113);
and U19385 (N_19385,N_16523,N_17440);
nand U19386 (N_19386,N_16237,N_16391);
nand U19387 (N_19387,N_17214,N_16551);
xor U19388 (N_19388,N_16255,N_17452);
nand U19389 (N_19389,N_17017,N_17763);
xor U19390 (N_19390,N_17715,N_17764);
nand U19391 (N_19391,N_16935,N_16085);
xnor U19392 (N_19392,N_16073,N_16928);
nand U19393 (N_19393,N_17329,N_17958);
or U19394 (N_19394,N_16561,N_17471);
or U19395 (N_19395,N_17651,N_17384);
and U19396 (N_19396,N_17810,N_17892);
nor U19397 (N_19397,N_16665,N_16139);
xor U19398 (N_19398,N_16623,N_17388);
nor U19399 (N_19399,N_17483,N_16083);
and U19400 (N_19400,N_16519,N_17467);
nor U19401 (N_19401,N_17869,N_16807);
nor U19402 (N_19402,N_16396,N_16769);
nor U19403 (N_19403,N_16373,N_16135);
nand U19404 (N_19404,N_16061,N_16872);
or U19405 (N_19405,N_16127,N_16870);
or U19406 (N_19406,N_17375,N_16264);
or U19407 (N_19407,N_16922,N_17034);
or U19408 (N_19408,N_17745,N_17278);
xor U19409 (N_19409,N_16439,N_16750);
or U19410 (N_19410,N_17712,N_17313);
and U19411 (N_19411,N_17818,N_17539);
and U19412 (N_19412,N_16794,N_16959);
and U19413 (N_19413,N_17110,N_16446);
and U19414 (N_19414,N_17038,N_17789);
or U19415 (N_19415,N_16899,N_16685);
xnor U19416 (N_19416,N_17066,N_17896);
nor U19417 (N_19417,N_17061,N_17343);
nor U19418 (N_19418,N_17083,N_17933);
and U19419 (N_19419,N_17624,N_16143);
xnor U19420 (N_19420,N_17779,N_16433);
nor U19421 (N_19421,N_16345,N_17526);
and U19422 (N_19422,N_17096,N_17848);
xor U19423 (N_19423,N_16264,N_16959);
or U19424 (N_19424,N_16798,N_16869);
or U19425 (N_19425,N_17258,N_16273);
nor U19426 (N_19426,N_16046,N_16948);
or U19427 (N_19427,N_17547,N_17004);
and U19428 (N_19428,N_17235,N_17227);
or U19429 (N_19429,N_17253,N_17463);
or U19430 (N_19430,N_16670,N_17330);
nand U19431 (N_19431,N_17729,N_16257);
nand U19432 (N_19432,N_16162,N_17163);
or U19433 (N_19433,N_16580,N_16552);
or U19434 (N_19434,N_17461,N_17290);
nand U19435 (N_19435,N_16387,N_17841);
nor U19436 (N_19436,N_17473,N_16990);
or U19437 (N_19437,N_16189,N_16269);
or U19438 (N_19438,N_16523,N_17929);
nand U19439 (N_19439,N_16031,N_17981);
and U19440 (N_19440,N_17595,N_16495);
and U19441 (N_19441,N_17593,N_17290);
nand U19442 (N_19442,N_16054,N_17514);
or U19443 (N_19443,N_17475,N_17428);
nand U19444 (N_19444,N_17054,N_16376);
and U19445 (N_19445,N_17925,N_17865);
nor U19446 (N_19446,N_17151,N_17311);
nand U19447 (N_19447,N_16346,N_16884);
and U19448 (N_19448,N_16662,N_16829);
and U19449 (N_19449,N_16570,N_16372);
nor U19450 (N_19450,N_17166,N_17063);
xnor U19451 (N_19451,N_16698,N_17641);
and U19452 (N_19452,N_16213,N_17161);
and U19453 (N_19453,N_16639,N_17259);
xor U19454 (N_19454,N_16119,N_17690);
or U19455 (N_19455,N_16253,N_16437);
nor U19456 (N_19456,N_17112,N_16661);
nor U19457 (N_19457,N_16578,N_16481);
and U19458 (N_19458,N_17810,N_16034);
or U19459 (N_19459,N_16158,N_17445);
or U19460 (N_19460,N_16540,N_17702);
or U19461 (N_19461,N_16108,N_16700);
or U19462 (N_19462,N_16576,N_17321);
nand U19463 (N_19463,N_16238,N_17025);
nand U19464 (N_19464,N_16588,N_16661);
nand U19465 (N_19465,N_16483,N_16824);
or U19466 (N_19466,N_16606,N_17258);
nand U19467 (N_19467,N_17136,N_17741);
or U19468 (N_19468,N_17662,N_16049);
and U19469 (N_19469,N_17713,N_16297);
nand U19470 (N_19470,N_16880,N_16671);
xor U19471 (N_19471,N_17120,N_16395);
or U19472 (N_19472,N_17049,N_17141);
or U19473 (N_19473,N_16040,N_17081);
nor U19474 (N_19474,N_16875,N_16051);
xnor U19475 (N_19475,N_17774,N_16552);
or U19476 (N_19476,N_17252,N_17540);
or U19477 (N_19477,N_17371,N_17472);
nand U19478 (N_19478,N_17471,N_16512);
nand U19479 (N_19479,N_17438,N_17407);
nor U19480 (N_19480,N_17311,N_16815);
xnor U19481 (N_19481,N_17429,N_17507);
xnor U19482 (N_19482,N_17839,N_16782);
and U19483 (N_19483,N_16657,N_17892);
or U19484 (N_19484,N_17417,N_17908);
nand U19485 (N_19485,N_16703,N_16423);
nor U19486 (N_19486,N_17490,N_16709);
or U19487 (N_19487,N_16619,N_16695);
xor U19488 (N_19488,N_17553,N_16536);
nor U19489 (N_19489,N_16556,N_16993);
or U19490 (N_19490,N_16842,N_17681);
and U19491 (N_19491,N_17890,N_16249);
or U19492 (N_19492,N_16517,N_16859);
and U19493 (N_19493,N_16416,N_16618);
nor U19494 (N_19494,N_16523,N_17053);
nand U19495 (N_19495,N_17782,N_16527);
nand U19496 (N_19496,N_16677,N_16611);
xor U19497 (N_19497,N_16742,N_16706);
or U19498 (N_19498,N_16718,N_17809);
nor U19499 (N_19499,N_17798,N_17552);
or U19500 (N_19500,N_16671,N_17101);
nor U19501 (N_19501,N_16542,N_16332);
nand U19502 (N_19502,N_16313,N_16183);
or U19503 (N_19503,N_16762,N_16967);
or U19504 (N_19504,N_17487,N_17851);
xnor U19505 (N_19505,N_16210,N_16033);
nor U19506 (N_19506,N_16480,N_17656);
xnor U19507 (N_19507,N_16744,N_16302);
nor U19508 (N_19508,N_17357,N_17503);
and U19509 (N_19509,N_16576,N_17358);
nand U19510 (N_19510,N_17626,N_17106);
and U19511 (N_19511,N_16865,N_16473);
nand U19512 (N_19512,N_16318,N_17066);
and U19513 (N_19513,N_16720,N_17919);
xor U19514 (N_19514,N_17574,N_17455);
or U19515 (N_19515,N_16537,N_16574);
and U19516 (N_19516,N_17275,N_16427);
and U19517 (N_19517,N_17023,N_17292);
nor U19518 (N_19518,N_17653,N_17198);
xor U19519 (N_19519,N_17558,N_17990);
and U19520 (N_19520,N_16619,N_16114);
or U19521 (N_19521,N_16785,N_16263);
or U19522 (N_19522,N_17766,N_17792);
nand U19523 (N_19523,N_16384,N_16341);
and U19524 (N_19524,N_17175,N_16056);
and U19525 (N_19525,N_17633,N_17551);
nor U19526 (N_19526,N_17814,N_16447);
and U19527 (N_19527,N_17188,N_16268);
nand U19528 (N_19528,N_17545,N_17012);
or U19529 (N_19529,N_16278,N_16229);
nor U19530 (N_19530,N_16181,N_17322);
or U19531 (N_19531,N_17687,N_17070);
xnor U19532 (N_19532,N_16837,N_17008);
nand U19533 (N_19533,N_16833,N_16148);
nor U19534 (N_19534,N_16397,N_16039);
or U19535 (N_19535,N_17752,N_16758);
xor U19536 (N_19536,N_17675,N_17168);
and U19537 (N_19537,N_17607,N_16623);
or U19538 (N_19538,N_17059,N_16628);
xor U19539 (N_19539,N_16456,N_16816);
nand U19540 (N_19540,N_17652,N_17062);
nor U19541 (N_19541,N_17127,N_16248);
nor U19542 (N_19542,N_16655,N_17080);
and U19543 (N_19543,N_17186,N_16285);
nor U19544 (N_19544,N_16793,N_16012);
or U19545 (N_19545,N_16556,N_16332);
and U19546 (N_19546,N_17558,N_16458);
nand U19547 (N_19547,N_17378,N_16690);
nand U19548 (N_19548,N_17305,N_16821);
nor U19549 (N_19549,N_16677,N_16111);
and U19550 (N_19550,N_17230,N_16575);
nand U19551 (N_19551,N_17179,N_17723);
or U19552 (N_19552,N_17868,N_17242);
nand U19553 (N_19553,N_17974,N_17135);
nor U19554 (N_19554,N_17664,N_16674);
xnor U19555 (N_19555,N_17475,N_17946);
and U19556 (N_19556,N_16853,N_16309);
nand U19557 (N_19557,N_17016,N_16992);
nor U19558 (N_19558,N_16696,N_17501);
nand U19559 (N_19559,N_16532,N_16159);
xnor U19560 (N_19560,N_16947,N_16507);
nand U19561 (N_19561,N_16546,N_16444);
and U19562 (N_19562,N_17154,N_16131);
and U19563 (N_19563,N_16583,N_16964);
or U19564 (N_19564,N_17632,N_17496);
or U19565 (N_19565,N_16560,N_17121);
xnor U19566 (N_19566,N_16115,N_17670);
or U19567 (N_19567,N_17610,N_17111);
nor U19568 (N_19568,N_16463,N_17716);
or U19569 (N_19569,N_17652,N_17304);
xor U19570 (N_19570,N_17652,N_17629);
xnor U19571 (N_19571,N_16164,N_17382);
and U19572 (N_19572,N_17002,N_17212);
xor U19573 (N_19573,N_17979,N_17210);
and U19574 (N_19574,N_16282,N_16293);
and U19575 (N_19575,N_17595,N_16346);
xnor U19576 (N_19576,N_16052,N_17724);
xnor U19577 (N_19577,N_16800,N_16364);
nand U19578 (N_19578,N_17972,N_17435);
or U19579 (N_19579,N_17525,N_17262);
xor U19580 (N_19580,N_17642,N_16279);
xnor U19581 (N_19581,N_17697,N_17082);
nor U19582 (N_19582,N_17304,N_16335);
nand U19583 (N_19583,N_17527,N_17839);
nand U19584 (N_19584,N_16920,N_16219);
xnor U19585 (N_19585,N_16471,N_17704);
or U19586 (N_19586,N_16253,N_17631);
nand U19587 (N_19587,N_16710,N_17436);
nor U19588 (N_19588,N_16881,N_17430);
or U19589 (N_19589,N_17908,N_17695);
xor U19590 (N_19590,N_17485,N_16236);
nand U19591 (N_19591,N_17341,N_16079);
xor U19592 (N_19592,N_16905,N_16913);
nor U19593 (N_19593,N_17485,N_16588);
nor U19594 (N_19594,N_17104,N_16205);
and U19595 (N_19595,N_16594,N_17134);
and U19596 (N_19596,N_17392,N_17728);
nand U19597 (N_19597,N_16011,N_16922);
nand U19598 (N_19598,N_16913,N_17040);
nor U19599 (N_19599,N_17293,N_17976);
nor U19600 (N_19600,N_16859,N_16217);
nor U19601 (N_19601,N_17075,N_16795);
or U19602 (N_19602,N_17526,N_17577);
and U19603 (N_19603,N_16647,N_16190);
or U19604 (N_19604,N_17178,N_16373);
nand U19605 (N_19605,N_17128,N_17748);
nor U19606 (N_19606,N_16931,N_17413);
nand U19607 (N_19607,N_16721,N_17430);
xor U19608 (N_19608,N_16484,N_16392);
or U19609 (N_19609,N_17435,N_16861);
or U19610 (N_19610,N_17365,N_16846);
xnor U19611 (N_19611,N_16856,N_16943);
nor U19612 (N_19612,N_16107,N_16444);
nand U19613 (N_19613,N_17069,N_16579);
nor U19614 (N_19614,N_16261,N_16032);
and U19615 (N_19615,N_17620,N_17400);
nor U19616 (N_19616,N_17581,N_16263);
and U19617 (N_19617,N_16755,N_17108);
and U19618 (N_19618,N_17529,N_17651);
nor U19619 (N_19619,N_16203,N_17201);
xnor U19620 (N_19620,N_17471,N_17952);
nand U19621 (N_19621,N_17162,N_16249);
xor U19622 (N_19622,N_17767,N_16130);
nand U19623 (N_19623,N_16076,N_17938);
xnor U19624 (N_19624,N_17874,N_17468);
nand U19625 (N_19625,N_16504,N_17244);
and U19626 (N_19626,N_17596,N_17295);
nand U19627 (N_19627,N_17934,N_16744);
xnor U19628 (N_19628,N_17379,N_16555);
xnor U19629 (N_19629,N_16627,N_16998);
xor U19630 (N_19630,N_17101,N_16865);
xnor U19631 (N_19631,N_16296,N_16672);
and U19632 (N_19632,N_16392,N_16065);
and U19633 (N_19633,N_17537,N_17303);
nor U19634 (N_19634,N_17953,N_17396);
or U19635 (N_19635,N_17127,N_17633);
or U19636 (N_19636,N_16788,N_17325);
nand U19637 (N_19637,N_16216,N_17013);
and U19638 (N_19638,N_17858,N_16359);
nor U19639 (N_19639,N_16053,N_16120);
and U19640 (N_19640,N_16811,N_17977);
xor U19641 (N_19641,N_17840,N_16188);
nand U19642 (N_19642,N_16228,N_16187);
and U19643 (N_19643,N_17316,N_17898);
and U19644 (N_19644,N_16549,N_17736);
nand U19645 (N_19645,N_16979,N_16060);
nor U19646 (N_19646,N_16606,N_17373);
and U19647 (N_19647,N_16094,N_17157);
and U19648 (N_19648,N_16384,N_17637);
and U19649 (N_19649,N_16261,N_16395);
nand U19650 (N_19650,N_16813,N_17591);
xnor U19651 (N_19651,N_17193,N_16679);
or U19652 (N_19652,N_16061,N_17806);
or U19653 (N_19653,N_17801,N_17376);
nand U19654 (N_19654,N_16445,N_16725);
and U19655 (N_19655,N_16171,N_17467);
nand U19656 (N_19656,N_17730,N_16276);
nor U19657 (N_19657,N_16043,N_17498);
or U19658 (N_19658,N_17781,N_17170);
or U19659 (N_19659,N_17368,N_17928);
nor U19660 (N_19660,N_17702,N_17963);
nor U19661 (N_19661,N_17605,N_17874);
xor U19662 (N_19662,N_17157,N_16614);
nor U19663 (N_19663,N_17003,N_17757);
or U19664 (N_19664,N_16015,N_16858);
nand U19665 (N_19665,N_16601,N_17456);
xnor U19666 (N_19666,N_16893,N_16111);
xor U19667 (N_19667,N_16547,N_17994);
xnor U19668 (N_19668,N_16881,N_16769);
and U19669 (N_19669,N_17373,N_17486);
nand U19670 (N_19670,N_17102,N_16810);
or U19671 (N_19671,N_16815,N_16048);
nand U19672 (N_19672,N_16320,N_17245);
and U19673 (N_19673,N_16485,N_16729);
xor U19674 (N_19674,N_16670,N_16984);
or U19675 (N_19675,N_17744,N_17767);
nor U19676 (N_19676,N_17206,N_17513);
xor U19677 (N_19677,N_17602,N_17999);
nor U19678 (N_19678,N_16580,N_16073);
nor U19679 (N_19679,N_16296,N_17751);
or U19680 (N_19680,N_16200,N_16118);
xnor U19681 (N_19681,N_16608,N_16200);
xor U19682 (N_19682,N_17923,N_16528);
and U19683 (N_19683,N_17084,N_17926);
nand U19684 (N_19684,N_16924,N_17921);
nand U19685 (N_19685,N_16613,N_17735);
or U19686 (N_19686,N_16855,N_16899);
and U19687 (N_19687,N_16267,N_17243);
and U19688 (N_19688,N_16124,N_17354);
nor U19689 (N_19689,N_17148,N_17451);
nor U19690 (N_19690,N_16744,N_16437);
and U19691 (N_19691,N_16097,N_16646);
nor U19692 (N_19692,N_16378,N_16368);
nor U19693 (N_19693,N_16796,N_16521);
and U19694 (N_19694,N_17194,N_17480);
xor U19695 (N_19695,N_17014,N_17409);
or U19696 (N_19696,N_17746,N_17581);
or U19697 (N_19697,N_16354,N_17680);
nand U19698 (N_19698,N_17334,N_16476);
and U19699 (N_19699,N_17119,N_16353);
nor U19700 (N_19700,N_17971,N_16005);
or U19701 (N_19701,N_17079,N_17042);
nand U19702 (N_19702,N_16836,N_17772);
nand U19703 (N_19703,N_16020,N_17067);
nand U19704 (N_19704,N_16120,N_17293);
xnor U19705 (N_19705,N_16011,N_17186);
xnor U19706 (N_19706,N_16399,N_16347);
nor U19707 (N_19707,N_16733,N_17917);
and U19708 (N_19708,N_17253,N_16404);
or U19709 (N_19709,N_17905,N_17733);
nor U19710 (N_19710,N_17003,N_17735);
nor U19711 (N_19711,N_16073,N_17328);
nand U19712 (N_19712,N_17883,N_17742);
xnor U19713 (N_19713,N_16273,N_16515);
nand U19714 (N_19714,N_16019,N_17536);
or U19715 (N_19715,N_16126,N_17219);
and U19716 (N_19716,N_16420,N_17112);
nor U19717 (N_19717,N_17744,N_16548);
xor U19718 (N_19718,N_16338,N_17029);
or U19719 (N_19719,N_17223,N_17345);
xnor U19720 (N_19720,N_17894,N_17065);
xnor U19721 (N_19721,N_17666,N_17689);
and U19722 (N_19722,N_16367,N_17677);
or U19723 (N_19723,N_16925,N_16336);
or U19724 (N_19724,N_17910,N_16477);
or U19725 (N_19725,N_16246,N_16685);
xnor U19726 (N_19726,N_17073,N_17121);
and U19727 (N_19727,N_16332,N_16107);
and U19728 (N_19728,N_16348,N_17747);
and U19729 (N_19729,N_16265,N_16361);
and U19730 (N_19730,N_16544,N_16113);
or U19731 (N_19731,N_16351,N_17952);
or U19732 (N_19732,N_16935,N_16757);
and U19733 (N_19733,N_17196,N_16665);
or U19734 (N_19734,N_16094,N_16557);
xor U19735 (N_19735,N_16687,N_16598);
nor U19736 (N_19736,N_17281,N_17394);
xnor U19737 (N_19737,N_17909,N_16322);
or U19738 (N_19738,N_17719,N_16344);
and U19739 (N_19739,N_16959,N_17274);
and U19740 (N_19740,N_17695,N_16116);
nor U19741 (N_19741,N_16609,N_17402);
and U19742 (N_19742,N_16576,N_17965);
and U19743 (N_19743,N_17442,N_16084);
and U19744 (N_19744,N_16628,N_16191);
and U19745 (N_19745,N_17489,N_16812);
xnor U19746 (N_19746,N_17390,N_16641);
xor U19747 (N_19747,N_17167,N_16415);
and U19748 (N_19748,N_17119,N_16266);
xor U19749 (N_19749,N_16514,N_17989);
or U19750 (N_19750,N_16015,N_17996);
and U19751 (N_19751,N_17069,N_17615);
nor U19752 (N_19752,N_16368,N_17010);
or U19753 (N_19753,N_17688,N_16239);
nor U19754 (N_19754,N_16784,N_16266);
nand U19755 (N_19755,N_17334,N_16543);
nand U19756 (N_19756,N_16289,N_17141);
nand U19757 (N_19757,N_17393,N_17109);
nor U19758 (N_19758,N_16423,N_16682);
and U19759 (N_19759,N_16141,N_16713);
nand U19760 (N_19760,N_17217,N_17131);
nand U19761 (N_19761,N_17344,N_17779);
or U19762 (N_19762,N_17446,N_17615);
and U19763 (N_19763,N_16145,N_16963);
xnor U19764 (N_19764,N_17651,N_17933);
xnor U19765 (N_19765,N_16398,N_16899);
or U19766 (N_19766,N_16328,N_17077);
nand U19767 (N_19767,N_17439,N_17563);
nand U19768 (N_19768,N_16966,N_16748);
and U19769 (N_19769,N_17979,N_16413);
nor U19770 (N_19770,N_16031,N_16191);
or U19771 (N_19771,N_17196,N_16295);
nand U19772 (N_19772,N_17384,N_16936);
xor U19773 (N_19773,N_16151,N_16472);
and U19774 (N_19774,N_17275,N_17269);
or U19775 (N_19775,N_17345,N_16027);
nor U19776 (N_19776,N_17098,N_17143);
nand U19777 (N_19777,N_16968,N_17694);
or U19778 (N_19778,N_16701,N_17740);
or U19779 (N_19779,N_17821,N_17453);
xnor U19780 (N_19780,N_16541,N_17654);
or U19781 (N_19781,N_17222,N_16074);
or U19782 (N_19782,N_17043,N_16137);
xor U19783 (N_19783,N_17370,N_17986);
nor U19784 (N_19784,N_16519,N_17514);
xnor U19785 (N_19785,N_16860,N_16065);
nor U19786 (N_19786,N_17467,N_17656);
or U19787 (N_19787,N_17533,N_17603);
and U19788 (N_19788,N_16494,N_16695);
and U19789 (N_19789,N_17146,N_17180);
and U19790 (N_19790,N_17851,N_17928);
and U19791 (N_19791,N_16138,N_16949);
xor U19792 (N_19792,N_17754,N_17215);
or U19793 (N_19793,N_16179,N_16929);
xnor U19794 (N_19794,N_17228,N_17798);
and U19795 (N_19795,N_16948,N_17918);
or U19796 (N_19796,N_17814,N_17100);
and U19797 (N_19797,N_17492,N_16426);
nand U19798 (N_19798,N_17435,N_17589);
and U19799 (N_19799,N_17752,N_17516);
nor U19800 (N_19800,N_16636,N_16504);
xor U19801 (N_19801,N_17849,N_16786);
nand U19802 (N_19802,N_16876,N_16640);
or U19803 (N_19803,N_17310,N_17666);
and U19804 (N_19804,N_16049,N_16425);
nor U19805 (N_19805,N_16776,N_16256);
and U19806 (N_19806,N_17796,N_17072);
and U19807 (N_19807,N_16580,N_17446);
nand U19808 (N_19808,N_17517,N_17739);
and U19809 (N_19809,N_17068,N_17134);
xnor U19810 (N_19810,N_17208,N_17635);
or U19811 (N_19811,N_17605,N_16220);
xor U19812 (N_19812,N_16933,N_17708);
nor U19813 (N_19813,N_16358,N_17802);
or U19814 (N_19814,N_16811,N_17777);
or U19815 (N_19815,N_16891,N_17306);
nor U19816 (N_19816,N_17810,N_16730);
nor U19817 (N_19817,N_16009,N_16343);
or U19818 (N_19818,N_17086,N_16193);
or U19819 (N_19819,N_17753,N_16973);
and U19820 (N_19820,N_17143,N_16637);
nand U19821 (N_19821,N_17733,N_17240);
nand U19822 (N_19822,N_16474,N_17531);
nor U19823 (N_19823,N_17787,N_16372);
nor U19824 (N_19824,N_16738,N_17152);
nand U19825 (N_19825,N_17117,N_17996);
or U19826 (N_19826,N_16447,N_16577);
nor U19827 (N_19827,N_17042,N_16772);
and U19828 (N_19828,N_16736,N_17724);
or U19829 (N_19829,N_16844,N_16955);
nor U19830 (N_19830,N_16604,N_16178);
or U19831 (N_19831,N_16322,N_17493);
or U19832 (N_19832,N_17830,N_17625);
nor U19833 (N_19833,N_17774,N_16600);
or U19834 (N_19834,N_16741,N_16247);
nand U19835 (N_19835,N_17306,N_17747);
nor U19836 (N_19836,N_16021,N_16756);
xnor U19837 (N_19837,N_16587,N_16968);
nor U19838 (N_19838,N_17141,N_17421);
nand U19839 (N_19839,N_17380,N_16139);
nor U19840 (N_19840,N_16269,N_17349);
xor U19841 (N_19841,N_16941,N_17036);
or U19842 (N_19842,N_16491,N_16941);
nor U19843 (N_19843,N_17977,N_17010);
and U19844 (N_19844,N_16317,N_17248);
or U19845 (N_19845,N_17273,N_17356);
nor U19846 (N_19846,N_17192,N_17629);
and U19847 (N_19847,N_17241,N_17053);
and U19848 (N_19848,N_16614,N_17488);
xor U19849 (N_19849,N_16757,N_17389);
and U19850 (N_19850,N_17451,N_16318);
nand U19851 (N_19851,N_16724,N_16741);
and U19852 (N_19852,N_17519,N_16088);
xnor U19853 (N_19853,N_17823,N_17311);
nand U19854 (N_19854,N_17406,N_16517);
nand U19855 (N_19855,N_17749,N_16719);
or U19856 (N_19856,N_16506,N_16082);
xnor U19857 (N_19857,N_17490,N_17955);
nand U19858 (N_19858,N_16909,N_16363);
nand U19859 (N_19859,N_17296,N_16635);
nor U19860 (N_19860,N_17862,N_17846);
and U19861 (N_19861,N_16297,N_17915);
or U19862 (N_19862,N_17510,N_16332);
and U19863 (N_19863,N_17589,N_17651);
and U19864 (N_19864,N_16343,N_16270);
or U19865 (N_19865,N_16644,N_16115);
and U19866 (N_19866,N_16004,N_16024);
xnor U19867 (N_19867,N_17986,N_17792);
xnor U19868 (N_19868,N_16045,N_17327);
or U19869 (N_19869,N_16222,N_17440);
nor U19870 (N_19870,N_16740,N_17411);
nand U19871 (N_19871,N_16918,N_16532);
or U19872 (N_19872,N_17989,N_16303);
nand U19873 (N_19873,N_17227,N_17490);
nor U19874 (N_19874,N_17868,N_16136);
and U19875 (N_19875,N_17016,N_17996);
nand U19876 (N_19876,N_16130,N_16495);
nand U19877 (N_19877,N_16735,N_17745);
nor U19878 (N_19878,N_17593,N_16913);
nand U19879 (N_19879,N_16705,N_16494);
nand U19880 (N_19880,N_17638,N_16005);
or U19881 (N_19881,N_17365,N_16983);
nand U19882 (N_19882,N_16495,N_16489);
nand U19883 (N_19883,N_17605,N_16758);
xnor U19884 (N_19884,N_17336,N_17479);
nand U19885 (N_19885,N_17896,N_16098);
nand U19886 (N_19886,N_17219,N_17397);
xor U19887 (N_19887,N_17546,N_16068);
nor U19888 (N_19888,N_17820,N_17156);
and U19889 (N_19889,N_16281,N_17009);
nor U19890 (N_19890,N_16162,N_16493);
nand U19891 (N_19891,N_16674,N_16363);
or U19892 (N_19892,N_17428,N_17238);
xnor U19893 (N_19893,N_16821,N_16840);
nor U19894 (N_19894,N_16727,N_16643);
xor U19895 (N_19895,N_17780,N_17349);
or U19896 (N_19896,N_16530,N_17625);
and U19897 (N_19897,N_17710,N_16437);
xnor U19898 (N_19898,N_17136,N_17024);
or U19899 (N_19899,N_16434,N_16285);
and U19900 (N_19900,N_17828,N_17098);
nor U19901 (N_19901,N_16795,N_17672);
nor U19902 (N_19902,N_16390,N_16636);
nor U19903 (N_19903,N_17484,N_17547);
nor U19904 (N_19904,N_16167,N_17872);
nand U19905 (N_19905,N_16460,N_16133);
nand U19906 (N_19906,N_16250,N_17695);
xnor U19907 (N_19907,N_16462,N_16935);
nand U19908 (N_19908,N_16343,N_17625);
and U19909 (N_19909,N_17619,N_17215);
nor U19910 (N_19910,N_17469,N_17375);
or U19911 (N_19911,N_16449,N_16050);
nor U19912 (N_19912,N_17681,N_16419);
and U19913 (N_19913,N_17907,N_16072);
and U19914 (N_19914,N_17922,N_17006);
nor U19915 (N_19915,N_16192,N_16463);
nand U19916 (N_19916,N_16509,N_16780);
xnor U19917 (N_19917,N_17421,N_17794);
or U19918 (N_19918,N_17293,N_16935);
and U19919 (N_19919,N_17772,N_17354);
nor U19920 (N_19920,N_17393,N_17218);
or U19921 (N_19921,N_17848,N_17661);
and U19922 (N_19922,N_17780,N_16169);
xor U19923 (N_19923,N_17399,N_16609);
xnor U19924 (N_19924,N_17276,N_17180);
and U19925 (N_19925,N_16218,N_16686);
nand U19926 (N_19926,N_16639,N_16207);
xor U19927 (N_19927,N_17576,N_17366);
and U19928 (N_19928,N_16198,N_17138);
or U19929 (N_19929,N_17101,N_17544);
and U19930 (N_19930,N_17732,N_16999);
nor U19931 (N_19931,N_16959,N_16121);
nor U19932 (N_19932,N_17991,N_16472);
and U19933 (N_19933,N_17857,N_16748);
nor U19934 (N_19934,N_17491,N_16423);
xnor U19935 (N_19935,N_16613,N_16382);
and U19936 (N_19936,N_16434,N_16446);
or U19937 (N_19937,N_17505,N_17820);
nand U19938 (N_19938,N_17564,N_17382);
nor U19939 (N_19939,N_16753,N_16848);
nor U19940 (N_19940,N_16713,N_16421);
xnor U19941 (N_19941,N_16246,N_17686);
and U19942 (N_19942,N_16874,N_16015);
nor U19943 (N_19943,N_17703,N_16125);
nor U19944 (N_19944,N_17735,N_17516);
or U19945 (N_19945,N_17524,N_17671);
and U19946 (N_19946,N_16906,N_17581);
xor U19947 (N_19947,N_16786,N_17198);
xor U19948 (N_19948,N_16308,N_17342);
xnor U19949 (N_19949,N_16870,N_17367);
xnor U19950 (N_19950,N_16567,N_17290);
and U19951 (N_19951,N_16334,N_16057);
and U19952 (N_19952,N_16755,N_16628);
nor U19953 (N_19953,N_17719,N_16446);
and U19954 (N_19954,N_17446,N_16333);
xnor U19955 (N_19955,N_16068,N_16501);
xor U19956 (N_19956,N_17998,N_17719);
nor U19957 (N_19957,N_16546,N_17392);
or U19958 (N_19958,N_16436,N_16760);
nand U19959 (N_19959,N_17890,N_16506);
and U19960 (N_19960,N_17265,N_16157);
nand U19961 (N_19961,N_17175,N_17639);
or U19962 (N_19962,N_17807,N_16798);
xnor U19963 (N_19963,N_16170,N_16197);
or U19964 (N_19964,N_16928,N_17719);
xnor U19965 (N_19965,N_17755,N_17602);
and U19966 (N_19966,N_17475,N_17751);
nor U19967 (N_19967,N_16513,N_17987);
xnor U19968 (N_19968,N_17740,N_16292);
xor U19969 (N_19969,N_17300,N_16297);
nand U19970 (N_19970,N_16568,N_16102);
nand U19971 (N_19971,N_16772,N_16766);
nand U19972 (N_19972,N_16750,N_16148);
and U19973 (N_19973,N_16016,N_17646);
nor U19974 (N_19974,N_17234,N_17264);
nor U19975 (N_19975,N_17206,N_16060);
or U19976 (N_19976,N_17889,N_17320);
nand U19977 (N_19977,N_17519,N_16750);
and U19978 (N_19978,N_16478,N_16605);
or U19979 (N_19979,N_17758,N_16304);
or U19980 (N_19980,N_16337,N_16537);
nor U19981 (N_19981,N_17805,N_17238);
and U19982 (N_19982,N_17997,N_16746);
and U19983 (N_19983,N_17190,N_17943);
or U19984 (N_19984,N_17753,N_17278);
xnor U19985 (N_19985,N_16160,N_16473);
nor U19986 (N_19986,N_17251,N_17453);
and U19987 (N_19987,N_16327,N_17579);
xnor U19988 (N_19988,N_16865,N_17827);
or U19989 (N_19989,N_16913,N_17391);
and U19990 (N_19990,N_17364,N_17549);
or U19991 (N_19991,N_17939,N_16764);
xor U19992 (N_19992,N_17541,N_16673);
xor U19993 (N_19993,N_16983,N_17464);
nor U19994 (N_19994,N_16751,N_17036);
nor U19995 (N_19995,N_16917,N_17678);
and U19996 (N_19996,N_17761,N_16585);
or U19997 (N_19997,N_17195,N_17185);
nor U19998 (N_19998,N_16467,N_17078);
or U19999 (N_19999,N_16462,N_17448);
nor UO_0 (O_0,N_19884,N_19302);
nand UO_1 (O_1,N_18845,N_19938);
or UO_2 (O_2,N_18448,N_18937);
or UO_3 (O_3,N_19596,N_18792);
nor UO_4 (O_4,N_19284,N_19294);
nor UO_5 (O_5,N_19799,N_18411);
nor UO_6 (O_6,N_18446,N_19949);
xor UO_7 (O_7,N_18739,N_18763);
nor UO_8 (O_8,N_19271,N_18035);
nand UO_9 (O_9,N_19202,N_19575);
nor UO_10 (O_10,N_19703,N_18017);
or UO_11 (O_11,N_18588,N_18677);
and UO_12 (O_12,N_18084,N_19570);
or UO_13 (O_13,N_19732,N_18460);
and UO_14 (O_14,N_19822,N_19680);
nand UO_15 (O_15,N_18082,N_19819);
and UO_16 (O_16,N_18001,N_18389);
nand UO_17 (O_17,N_19869,N_18108);
xnor UO_18 (O_18,N_19129,N_19356);
nand UO_19 (O_19,N_19487,N_19228);
or UO_20 (O_20,N_18644,N_18440);
or UO_21 (O_21,N_18343,N_19465);
and UO_22 (O_22,N_18226,N_18847);
nand UO_23 (O_23,N_18419,N_18351);
nand UO_24 (O_24,N_18072,N_18224);
xnor UO_25 (O_25,N_19892,N_18135);
and UO_26 (O_26,N_19577,N_19675);
or UO_27 (O_27,N_18578,N_19134);
nand UO_28 (O_28,N_18742,N_18882);
nand UO_29 (O_29,N_19462,N_18597);
or UO_30 (O_30,N_19082,N_18934);
nor UO_31 (O_31,N_19138,N_18012);
and UO_32 (O_32,N_18288,N_19880);
nor UO_33 (O_33,N_18488,N_19063);
and UO_34 (O_34,N_19497,N_19486);
and UO_35 (O_35,N_18561,N_18788);
and UO_36 (O_36,N_18817,N_18933);
or UO_37 (O_37,N_18799,N_18136);
nand UO_38 (O_38,N_18965,N_19862);
nand UO_39 (O_39,N_19427,N_19917);
or UO_40 (O_40,N_19641,N_18856);
or UO_41 (O_41,N_18380,N_18600);
nand UO_42 (O_42,N_18397,N_19968);
and UO_43 (O_43,N_18852,N_18829);
and UO_44 (O_44,N_19125,N_18137);
xnor UO_45 (O_45,N_19760,N_19094);
or UO_46 (O_46,N_19708,N_19610);
nor UO_47 (O_47,N_18276,N_19064);
xor UO_48 (O_48,N_18443,N_18944);
and UO_49 (O_49,N_19519,N_18245);
nor UO_50 (O_50,N_18275,N_18549);
and UO_51 (O_51,N_19456,N_19752);
nand UO_52 (O_52,N_18257,N_18144);
nand UO_53 (O_53,N_19906,N_19077);
nor UO_54 (O_54,N_19816,N_18004);
nor UO_55 (O_55,N_18326,N_19208);
nand UO_56 (O_56,N_18114,N_18761);
xnor UO_57 (O_57,N_18370,N_19721);
nor UO_58 (O_58,N_19972,N_19056);
or UO_59 (O_59,N_19369,N_18489);
nand UO_60 (O_60,N_19429,N_18943);
or UO_61 (O_61,N_18348,N_19672);
and UO_62 (O_62,N_19850,N_19395);
and UO_63 (O_63,N_18520,N_19109);
nand UO_64 (O_64,N_18731,N_18790);
xnor UO_65 (O_65,N_19644,N_18220);
nand UO_66 (O_66,N_19414,N_18773);
or UO_67 (O_67,N_19691,N_19155);
and UO_68 (O_68,N_18005,N_18759);
and UO_69 (O_69,N_18422,N_19120);
xor UO_70 (O_70,N_18703,N_19187);
nand UO_71 (O_71,N_19670,N_18715);
or UO_72 (O_72,N_19236,N_19810);
and UO_73 (O_73,N_19866,N_18320);
nor UO_74 (O_74,N_18734,N_19081);
nor UO_75 (O_75,N_19458,N_18212);
and UO_76 (O_76,N_19964,N_18795);
nand UO_77 (O_77,N_19553,N_18307);
nor UO_78 (O_78,N_19558,N_18689);
xnor UO_79 (O_79,N_18096,N_18719);
or UO_80 (O_80,N_19279,N_18431);
and UO_81 (O_81,N_18936,N_19740);
or UO_82 (O_82,N_18755,N_18639);
or UO_83 (O_83,N_19895,N_18736);
or UO_84 (O_84,N_19940,N_18093);
or UO_85 (O_85,N_18319,N_19591);
or UO_86 (O_86,N_19009,N_19190);
xor UO_87 (O_87,N_18453,N_18045);
or UO_88 (O_88,N_19368,N_18194);
xor UO_89 (O_89,N_18304,N_18570);
or UO_90 (O_90,N_18798,N_19923);
or UO_91 (O_91,N_18808,N_18617);
nand UO_92 (O_92,N_19903,N_19909);
and UO_93 (O_93,N_19253,N_18985);
xor UO_94 (O_94,N_19100,N_19153);
nand UO_95 (O_95,N_18113,N_18784);
nor UO_96 (O_96,N_18071,N_18328);
nor UO_97 (O_97,N_19685,N_19256);
xnor UO_98 (O_98,N_19426,N_18993);
or UO_99 (O_99,N_19882,N_18608);
nor UO_100 (O_100,N_19742,N_18880);
xnor UO_101 (O_101,N_18503,N_18718);
and UO_102 (O_102,N_18474,N_19332);
and UO_103 (O_103,N_19551,N_19212);
nor UO_104 (O_104,N_18458,N_18381);
nor UO_105 (O_105,N_19635,N_18014);
and UO_106 (O_106,N_19258,N_18191);
and UO_107 (O_107,N_19461,N_18804);
or UO_108 (O_108,N_19029,N_18160);
nand UO_109 (O_109,N_19615,N_18626);
and UO_110 (O_110,N_18374,N_19043);
and UO_111 (O_111,N_18657,N_19702);
nor UO_112 (O_112,N_18636,N_18674);
nand UO_113 (O_113,N_19586,N_19965);
nand UO_114 (O_114,N_19539,N_18055);
nor UO_115 (O_115,N_19375,N_18182);
nor UO_116 (O_116,N_18438,N_19676);
nand UO_117 (O_117,N_18415,N_19144);
or UO_118 (O_118,N_18185,N_19027);
or UO_119 (O_119,N_18686,N_19993);
or UO_120 (O_120,N_18498,N_18913);
nor UO_121 (O_121,N_19677,N_18254);
nand UO_122 (O_122,N_18080,N_18065);
nand UO_123 (O_123,N_19700,N_19441);
or UO_124 (O_124,N_18234,N_19418);
nor UO_125 (O_125,N_19582,N_18542);
xor UO_126 (O_126,N_18083,N_19197);
or UO_127 (O_127,N_18372,N_19560);
and UO_128 (O_128,N_18339,N_19154);
nor UO_129 (O_129,N_19446,N_19374);
or UO_130 (O_130,N_18584,N_19899);
or UO_131 (O_131,N_18537,N_18586);
nand UO_132 (O_132,N_18623,N_19734);
nand UO_133 (O_133,N_18420,N_19293);
xor UO_134 (O_134,N_18454,N_18764);
nor UO_135 (O_135,N_19436,N_18874);
xor UO_136 (O_136,N_19058,N_18078);
xor UO_137 (O_137,N_18541,N_19412);
or UO_138 (O_138,N_18692,N_19124);
xnor UO_139 (O_139,N_19597,N_18827);
nor UO_140 (O_140,N_18655,N_18059);
nor UO_141 (O_141,N_19218,N_19180);
xnor UO_142 (O_142,N_18138,N_18289);
and UO_143 (O_143,N_18077,N_18189);
nand UO_144 (O_144,N_19142,N_19706);
or UO_145 (O_145,N_18910,N_18412);
or UO_146 (O_146,N_18293,N_18949);
xnor UO_147 (O_147,N_19921,N_19074);
nand UO_148 (O_148,N_18352,N_18610);
nor UO_149 (O_149,N_18831,N_18346);
nand UO_150 (O_150,N_18252,N_18063);
nor UO_151 (O_151,N_18101,N_19765);
or UO_152 (O_152,N_19744,N_18920);
or UO_153 (O_153,N_19380,N_18511);
nor UO_154 (O_154,N_19699,N_19737);
nand UO_155 (O_155,N_18268,N_19502);
nor UO_156 (O_156,N_19969,N_18482);
and UO_157 (O_157,N_19847,N_19557);
or UO_158 (O_158,N_19546,N_18721);
and UO_159 (O_159,N_19001,N_18475);
or UO_160 (O_160,N_18039,N_18955);
and UO_161 (O_161,N_19995,N_18513);
or UO_162 (O_162,N_18879,N_19397);
and UO_163 (O_163,N_19612,N_18914);
xnor UO_164 (O_164,N_18036,N_19894);
nor UO_165 (O_165,N_19164,N_19196);
nor UO_166 (O_166,N_19114,N_19472);
xor UO_167 (O_167,N_19123,N_18557);
and UO_168 (O_168,N_19751,N_19337);
or UO_169 (O_169,N_18204,N_19851);
and UO_170 (O_170,N_19014,N_19898);
nand UO_171 (O_171,N_19363,N_18461);
nor UO_172 (O_172,N_18786,N_19747);
nor UO_173 (O_173,N_18368,N_19915);
xor UO_174 (O_174,N_18669,N_19046);
nand UO_175 (O_175,N_19119,N_18400);
or UO_176 (O_176,N_18118,N_18890);
xor UO_177 (O_177,N_19085,N_18291);
and UO_178 (O_178,N_18873,N_18439);
xnor UO_179 (O_179,N_19891,N_19825);
nand UO_180 (O_180,N_18067,N_19592);
nand UO_181 (O_181,N_19645,N_18818);
and UO_182 (O_182,N_18553,N_19836);
nand UO_183 (O_183,N_18158,N_18297);
nor UO_184 (O_184,N_18162,N_19952);
nor UO_185 (O_185,N_19606,N_19494);
xor UO_186 (O_186,N_19070,N_19311);
nor UO_187 (O_187,N_19693,N_19352);
and UO_188 (O_188,N_19372,N_18382);
nand UO_189 (O_189,N_18978,N_19888);
xor UO_190 (O_190,N_19926,N_18208);
nor UO_191 (O_191,N_18909,N_18337);
nor UO_192 (O_192,N_19141,N_19096);
nand UO_193 (O_193,N_18714,N_19299);
xor UO_194 (O_194,N_18848,N_19562);
xnor UO_195 (O_195,N_19957,N_19581);
nor UO_196 (O_196,N_18170,N_19629);
or UO_197 (O_197,N_19479,N_18865);
or UO_198 (O_198,N_19541,N_19460);
and UO_199 (O_199,N_18505,N_18813);
or UO_200 (O_200,N_18637,N_19285);
and UO_201 (O_201,N_18127,N_18793);
and UO_202 (O_202,N_18668,N_18535);
nor UO_203 (O_203,N_19997,N_19942);
or UO_204 (O_204,N_18311,N_18760);
and UO_205 (O_205,N_18534,N_19841);
or UO_206 (O_206,N_18595,N_19314);
and UO_207 (O_207,N_18390,N_18075);
nand UO_208 (O_208,N_19687,N_19291);
nor UO_209 (O_209,N_19470,N_18531);
or UO_210 (O_210,N_18926,N_19049);
and UO_211 (O_211,N_18551,N_18086);
and UO_212 (O_212,N_19767,N_19053);
nor UO_213 (O_213,N_19468,N_19286);
xor UO_214 (O_214,N_19726,N_19445);
or UO_215 (O_215,N_18302,N_18956);
or UO_216 (O_216,N_18952,N_18049);
and UO_217 (O_217,N_19944,N_19137);
xnor UO_218 (O_218,N_19733,N_18215);
or UO_219 (O_219,N_18230,N_19878);
or UO_220 (O_220,N_18277,N_19107);
nand UO_221 (O_221,N_18652,N_18839);
nor UO_222 (O_222,N_19438,N_19994);
or UO_223 (O_223,N_18394,N_19370);
xor UO_224 (O_224,N_19607,N_18476);
or UO_225 (O_225,N_19268,N_18425);
nand UO_226 (O_226,N_19391,N_18164);
nand UO_227 (O_227,N_18213,N_18305);
nand UO_228 (O_228,N_18332,N_18423);
and UO_229 (O_229,N_19229,N_19201);
nand UO_230 (O_230,N_18457,N_18960);
nand UO_231 (O_231,N_19867,N_18698);
xnor UO_232 (O_232,N_18941,N_19413);
or UO_233 (O_233,N_19147,N_18050);
nor UO_234 (O_234,N_18139,N_18508);
and UO_235 (O_235,N_19642,N_18768);
or UO_236 (O_236,N_18079,N_19755);
xnor UO_237 (O_237,N_18727,N_18969);
nand UO_238 (O_238,N_18340,N_18321);
or UO_239 (O_239,N_19222,N_19934);
nand UO_240 (O_240,N_18591,N_18860);
or UO_241 (O_241,N_18497,N_19624);
or UO_242 (O_242,N_18814,N_18911);
or UO_243 (O_243,N_19110,N_19879);
and UO_244 (O_244,N_18056,N_19179);
and UO_245 (O_245,N_19240,N_18717);
or UO_246 (O_246,N_18587,N_19861);
or UO_247 (O_247,N_19140,N_18616);
and UO_248 (O_248,N_19051,N_19312);
and UO_249 (O_249,N_18809,N_18762);
or UO_250 (O_250,N_19274,N_19695);
and UO_251 (O_251,N_18579,N_19627);
nor UO_252 (O_252,N_19566,N_18507);
nand UO_253 (O_253,N_19555,N_18525);
xor UO_254 (O_254,N_18026,N_19349);
and UO_255 (O_255,N_19501,N_19617);
nand UO_256 (O_256,N_18436,N_19233);
and UO_257 (O_257,N_18885,N_18621);
xor UO_258 (O_258,N_19628,N_18115);
or UO_259 (O_259,N_19287,N_18950);
xor UO_260 (O_260,N_18961,N_19908);
or UO_261 (O_261,N_19408,N_19450);
nor UO_262 (O_262,N_19168,N_19219);
or UO_263 (O_263,N_19792,N_19556);
nand UO_264 (O_264,N_18068,N_18401);
nor UO_265 (O_265,N_18463,N_18735);
nor UO_266 (O_266,N_19317,N_18408);
nor UO_267 (O_267,N_19812,N_18317);
xnor UO_268 (O_268,N_19843,N_19184);
nand UO_269 (O_269,N_19636,N_19748);
nor UO_270 (O_270,N_18824,N_18875);
nand UO_271 (O_271,N_18345,N_19975);
and UO_272 (O_272,N_18679,N_18925);
xnor UO_273 (O_273,N_19528,N_18713);
xnor UO_274 (O_274,N_19913,N_19604);
or UO_275 (O_275,N_18939,N_19336);
nor UO_276 (O_276,N_18061,N_18152);
and UO_277 (O_277,N_18833,N_18267);
nand UO_278 (O_278,N_18938,N_19055);
nor UO_279 (O_279,N_18119,N_19045);
and UO_280 (O_280,N_18266,N_18310);
nand UO_281 (O_281,N_18524,N_18362);
and UO_282 (O_282,N_18968,N_18177);
and UO_283 (O_283,N_19378,N_19736);
and UO_284 (O_284,N_18878,N_19933);
or UO_285 (O_285,N_19002,N_19743);
nor UO_286 (O_286,N_18414,N_19531);
nor UO_287 (O_287,N_18855,N_19105);
nand UO_288 (O_288,N_18986,N_19814);
or UO_289 (O_289,N_18556,N_18284);
xor UO_290 (O_290,N_18881,N_18173);
nor UO_291 (O_291,N_19037,N_19951);
nor UO_292 (O_292,N_19663,N_19651);
nor UO_293 (O_293,N_19326,N_19015);
or UO_294 (O_294,N_18494,N_19243);
xnor UO_295 (O_295,N_18815,N_18104);
xor UO_296 (O_296,N_18546,N_19488);
or UO_297 (O_297,N_19999,N_18020);
nand UO_298 (O_298,N_18218,N_18514);
xor UO_299 (O_299,N_18201,N_18782);
nand UO_300 (O_300,N_18239,N_18749);
or UO_301 (O_301,N_19741,N_19455);
nor UO_302 (O_302,N_18812,N_18977);
nand UO_303 (O_303,N_19000,N_19621);
and UO_304 (O_304,N_19571,N_18334);
nor UO_305 (O_305,N_19221,N_19080);
nor UO_306 (O_306,N_18298,N_19602);
xnor UO_307 (O_307,N_18000,N_18583);
or UO_308 (O_308,N_19682,N_19102);
nor UO_309 (O_309,N_19204,N_18603);
xor UO_310 (O_310,N_19381,N_18921);
and UO_311 (O_311,N_18009,N_19247);
nor UO_312 (O_312,N_18540,N_18386);
and UO_313 (O_313,N_18073,N_18918);
nand UO_314 (O_314,N_19669,N_19855);
and UO_315 (O_315,N_18738,N_19276);
nand UO_316 (O_316,N_19265,N_19665);
xnor UO_317 (O_317,N_19170,N_18350);
xnor UO_318 (O_318,N_19595,N_18601);
nor UO_319 (O_319,N_18145,N_19637);
or UO_320 (O_320,N_19333,N_18406);
or UO_321 (O_321,N_19829,N_18013);
nand UO_322 (O_322,N_19377,N_19321);
nand UO_323 (O_323,N_19347,N_18258);
or UO_324 (O_324,N_18744,N_18512);
and UO_325 (O_325,N_18479,N_18046);
and UO_326 (O_326,N_19515,N_19773);
nand UO_327 (O_327,N_18244,N_18629);
nand UO_328 (O_328,N_18342,N_18264);
nand UO_329 (O_329,N_18702,N_18990);
xor UO_330 (O_330,N_19873,N_18450);
xor UO_331 (O_331,N_19630,N_18445);
or UO_332 (O_332,N_18757,N_19513);
xnor UO_333 (O_333,N_19133,N_18923);
or UO_334 (O_334,N_18867,N_19342);
and UO_335 (O_335,N_19146,N_19424);
or UO_336 (O_336,N_19684,N_19567);
nand UO_337 (O_337,N_18746,N_19984);
nor UO_338 (O_338,N_19076,N_18642);
or UO_339 (O_339,N_19805,N_18286);
and UO_340 (O_340,N_19626,N_18772);
and UO_341 (O_341,N_18037,N_19303);
and UO_342 (O_342,N_19970,N_18146);
nor UO_343 (O_343,N_19778,N_19028);
nor UO_344 (O_344,N_18946,N_19503);
xnor UO_345 (O_345,N_19537,N_18199);
xor UO_346 (O_346,N_19690,N_18861);
and UO_347 (O_347,N_18271,N_18912);
xnor UO_348 (O_348,N_19713,N_18331);
or UO_349 (O_349,N_18560,N_19393);
or UO_350 (O_350,N_18700,N_18002);
xnor UO_351 (O_351,N_18504,N_19603);
and UO_352 (O_352,N_19067,N_19280);
xor UO_353 (O_353,N_18997,N_19648);
or UO_354 (O_354,N_18087,N_19833);
xnor UO_355 (O_355,N_18929,N_19200);
nand UO_356 (O_356,N_19191,N_18859);
nand UO_357 (O_357,N_18052,N_19764);
and UO_358 (O_358,N_18519,N_18243);
nor UO_359 (O_359,N_18095,N_19887);
and UO_360 (O_360,N_19667,N_18970);
nor UO_361 (O_361,N_18898,N_19937);
nand UO_362 (O_362,N_18708,N_19121);
nand UO_363 (O_363,N_18336,N_18236);
and UO_364 (O_364,N_19505,N_19674);
and UO_365 (O_365,N_18521,N_19533);
nand UO_366 (O_366,N_18041,N_18850);
and UO_367 (O_367,N_18441,N_18159);
nor UO_368 (O_368,N_19453,N_18424);
and UO_369 (O_369,N_18982,N_18229);
and UO_370 (O_370,N_19139,N_18132);
and UO_371 (O_371,N_19206,N_18030);
xor UO_372 (O_372,N_19784,N_18251);
and UO_373 (O_373,N_18870,N_19485);
nand UO_374 (O_374,N_19012,N_18558);
and UO_375 (O_375,N_18043,N_19731);
nor UO_376 (O_376,N_18681,N_19449);
xor UO_377 (O_377,N_18186,N_18038);
nor UO_378 (O_378,N_18958,N_19839);
xor UO_379 (O_379,N_19774,N_19868);
xor UO_380 (O_380,N_18031,N_19289);
or UO_381 (O_381,N_18754,N_19152);
xor UO_382 (O_382,N_18076,N_19217);
and UO_383 (O_383,N_19955,N_19463);
and UO_384 (O_384,N_18491,N_19283);
nand UO_385 (O_385,N_18712,N_19366);
or UO_386 (O_386,N_18573,N_19019);
or UO_387 (O_387,N_18948,N_18427);
nand UO_388 (O_388,N_18989,N_18435);
or UO_389 (O_389,N_19480,N_18327);
or UO_390 (O_390,N_18680,N_18205);
and UO_391 (O_391,N_19950,N_18315);
xor UO_392 (O_392,N_18274,N_19335);
and UO_393 (O_393,N_18906,N_19145);
or UO_394 (O_394,N_18641,N_19264);
and UO_395 (O_395,N_19116,N_19504);
or UO_396 (O_396,N_18193,N_19569);
and UO_397 (O_397,N_18722,N_19495);
or UO_398 (O_398,N_19203,N_18018);
nand UO_399 (O_399,N_18613,N_19820);
and UO_400 (O_400,N_19579,N_18255);
or UO_401 (O_401,N_18697,N_19404);
nor UO_402 (O_402,N_19182,N_19789);
nor UO_403 (O_403,N_19163,N_19960);
and UO_404 (O_404,N_18140,N_19447);
xor UO_405 (O_405,N_19749,N_18515);
xnor UO_406 (O_406,N_19988,N_19981);
nand UO_407 (O_407,N_19787,N_19547);
nor UO_408 (O_408,N_19300,N_19739);
and UO_409 (O_409,N_18647,N_19392);
nand UO_410 (O_410,N_19098,N_19935);
and UO_411 (O_411,N_19664,N_19719);
nand UO_412 (O_412,N_18092,N_19273);
or UO_413 (O_413,N_18147,N_19160);
or UO_414 (O_414,N_19007,N_19267);
and UO_415 (O_415,N_19410,N_19471);
xor UO_416 (O_416,N_18869,N_18029);
xor UO_417 (O_417,N_18842,N_19167);
or UO_418 (O_418,N_19622,N_19018);
nor UO_419 (O_419,N_18103,N_19351);
or UO_420 (O_420,N_18499,N_18957);
and UO_421 (O_421,N_19928,N_18606);
nand UO_422 (O_422,N_18783,N_18306);
nand UO_423 (O_423,N_19039,N_18375);
nand UO_424 (O_424,N_19662,N_18574);
and UO_425 (O_425,N_18429,N_18330);
nand UO_426 (O_426,N_19788,N_19756);
nor UO_427 (O_427,N_19428,N_18976);
xor UO_428 (O_428,N_18094,N_19069);
nand UO_429 (O_429,N_19339,N_19260);
nand UO_430 (O_430,N_19440,N_18568);
nand UO_431 (O_431,N_19842,N_19172);
and UO_432 (O_432,N_19901,N_18893);
nand UO_433 (O_433,N_19982,N_19681);
xor UO_434 (O_434,N_18467,N_19930);
and UO_435 (O_435,N_19697,N_18575);
and UO_436 (O_436,N_18884,N_18901);
and UO_437 (O_437,N_19493,N_19239);
or UO_438 (O_438,N_18971,N_18111);
nor UO_439 (O_439,N_18577,N_18559);
or UO_440 (O_440,N_18016,N_19771);
nand UO_441 (O_441,N_18858,N_19931);
xor UO_442 (O_442,N_18635,N_19978);
nor UO_443 (O_443,N_18379,N_18235);
xor UO_444 (O_444,N_19897,N_18270);
xnor UO_445 (O_445,N_18572,N_19097);
and UO_446 (O_446,N_18733,N_19729);
or UO_447 (O_447,N_19896,N_19384);
and UO_448 (O_448,N_18344,N_18518);
xnor UO_449 (O_449,N_19156,N_18387);
or UO_450 (O_450,N_19047,N_19980);
nor UO_451 (O_451,N_19815,N_18025);
nand UO_452 (O_452,N_18886,N_18273);
nand UO_453 (O_453,N_19091,N_19623);
or UO_454 (O_454,N_19126,N_18751);
nand UO_455 (O_455,N_18979,N_18769);
xor UO_456 (O_456,N_18384,N_19529);
or UO_457 (O_457,N_18922,N_19824);
or UO_458 (O_458,N_19709,N_19827);
or UO_459 (O_459,N_18154,N_18027);
xor UO_460 (O_460,N_18047,N_18042);
nand UO_461 (O_461,N_19176,N_18149);
or UO_462 (O_462,N_19945,N_18688);
nor UO_463 (O_463,N_19220,N_18807);
or UO_464 (O_464,N_19244,N_18483);
or UO_465 (O_465,N_18192,N_18180);
nor UO_466 (O_466,N_19334,N_18709);
xor UO_467 (O_467,N_19041,N_19157);
nand UO_468 (O_468,N_19956,N_18527);
or UO_469 (O_469,N_18155,N_18896);
or UO_470 (O_470,N_18278,N_19409);
or UO_471 (O_471,N_19315,N_19671);
nor UO_472 (O_472,N_18596,N_19376);
nand UO_473 (O_473,N_18385,N_19532);
xor UO_474 (O_474,N_19946,N_19927);
nor UO_475 (O_475,N_18417,N_19506);
xor UO_476 (O_476,N_18023,N_19213);
nor UO_477 (O_477,N_18260,N_18720);
or UO_478 (O_478,N_19389,N_18355);
xnor UO_479 (O_479,N_19166,N_18353);
nand UO_480 (O_480,N_18219,N_19095);
or UO_481 (O_481,N_19211,N_18991);
or UO_482 (O_482,N_19360,N_19534);
and UO_483 (O_483,N_18231,N_19373);
nor UO_484 (O_484,N_18699,N_18951);
xor UO_485 (O_485,N_18820,N_18428);
nor UO_486 (O_486,N_19990,N_18410);
xor UO_487 (O_487,N_18007,N_18843);
xnor UO_488 (O_488,N_18032,N_19893);
nor UO_489 (O_489,N_19297,N_18631);
nor UO_490 (O_490,N_19275,N_18416);
nand UO_491 (O_491,N_19136,N_18089);
and UO_492 (O_492,N_19728,N_18543);
nand UO_493 (O_493,N_18667,N_18369);
nor UO_494 (O_494,N_18464,N_19912);
or UO_495 (O_495,N_18241,N_18857);
xor UO_496 (O_496,N_19905,N_19073);
nand UO_497 (O_497,N_18455,N_19989);
xnor UO_498 (O_498,N_18724,N_19590);
and UO_499 (O_499,N_18544,N_18102);
or UO_500 (O_500,N_19177,N_19775);
nor UO_501 (O_501,N_18085,N_19158);
and UO_502 (O_502,N_19593,N_19407);
nor UO_503 (O_503,N_19161,N_18183);
xnor UO_504 (O_504,N_19904,N_18396);
nand UO_505 (O_505,N_18547,N_18123);
nor UO_506 (O_506,N_19023,N_19763);
and UO_507 (O_507,N_18341,N_19178);
nand UO_508 (O_508,N_18308,N_18179);
and UO_509 (O_509,N_18725,N_18862);
and UO_510 (O_510,N_19712,N_19338);
or UO_511 (O_511,N_18200,N_19242);
nand UO_512 (O_512,N_19044,N_18645);
xor UO_513 (O_513,N_19288,N_19099);
and UO_514 (O_514,N_19075,N_19341);
nand UO_515 (O_515,N_18116,N_18643);
or UO_516 (O_516,N_18178,N_19481);
and UO_517 (O_517,N_19402,N_18444);
nand UO_518 (O_518,N_19795,N_18282);
nand UO_519 (O_519,N_18054,N_19552);
and UO_520 (O_520,N_18552,N_19886);
and UO_521 (O_521,N_18983,N_18625);
and UO_522 (O_522,N_19406,N_18391);
nand UO_523 (O_523,N_19848,N_18388);
xnor UO_524 (O_524,N_19151,N_19722);
or UO_525 (O_525,N_18548,N_18409);
nand UO_526 (O_526,N_19521,N_19359);
nand UO_527 (O_527,N_18916,N_19425);
xor UO_528 (O_528,N_18377,N_18051);
and UO_529 (O_529,N_19772,N_19601);
xor UO_530 (O_530,N_18675,N_18484);
nand UO_531 (O_531,N_19199,N_18188);
or UO_532 (O_532,N_19710,N_18227);
nor UO_533 (O_533,N_18040,N_18432);
xnor UO_534 (O_534,N_18705,N_18452);
and UO_535 (O_535,N_19522,N_19507);
nand UO_536 (O_536,N_18301,N_18648);
or UO_537 (O_537,N_19840,N_18285);
nor UO_538 (O_538,N_18854,N_19062);
or UO_539 (O_539,N_18981,N_19159);
and UO_540 (O_540,N_19396,N_19962);
xor UO_541 (O_541,N_19459,N_18895);
or UO_542 (O_542,N_19542,N_18840);
nand UO_543 (O_543,N_19066,N_19004);
or UO_544 (O_544,N_18221,N_19250);
and UO_545 (O_545,N_19226,N_18805);
nor UO_546 (O_546,N_18128,N_19800);
and UO_547 (O_547,N_19512,N_19929);
xnor UO_548 (O_548,N_19545,N_19089);
xnor UO_549 (O_549,N_19216,N_18313);
nand UO_550 (O_550,N_18184,N_19059);
and UO_551 (O_551,N_18133,N_19292);
xor UO_552 (O_552,N_18516,N_18758);
xnor UO_553 (O_553,N_19966,N_18582);
and UO_554 (O_554,N_18902,N_18299);
or UO_555 (O_555,N_19423,N_19103);
or UO_556 (O_556,N_19162,N_18994);
xnor UO_557 (O_557,N_19563,N_19809);
or UO_558 (O_558,N_19794,N_18329);
or UO_559 (O_559,N_18710,N_19011);
xnor UO_560 (O_560,N_18671,N_19259);
or UO_561 (O_561,N_18034,N_18202);
nand UO_562 (O_562,N_18003,N_18653);
nor UO_563 (O_563,N_18261,N_18737);
xor UO_564 (O_564,N_18661,N_18048);
and UO_565 (O_565,N_18849,N_18581);
nor UO_566 (O_566,N_18066,N_19768);
nand UO_567 (O_567,N_18743,N_18565);
nand UO_568 (O_568,N_18130,N_18413);
nand UO_569 (O_569,N_19169,N_19065);
nand UO_570 (O_570,N_19245,N_18728);
or UO_571 (O_571,N_19776,N_19050);
nor UO_572 (O_572,N_19186,N_18395);
and UO_573 (O_573,N_19821,N_18917);
nor UO_574 (O_574,N_19826,N_18117);
nor UO_575 (O_575,N_18609,N_19498);
xor UO_576 (O_576,N_18673,N_18373);
nand UO_577 (O_577,N_19738,N_19467);
nand UO_578 (O_578,N_19727,N_18682);
nand UO_579 (O_579,N_18607,N_19278);
xnor UO_580 (O_580,N_18090,N_19261);
and UO_581 (O_581,N_18908,N_19026);
xnor UO_582 (O_582,N_18566,N_19415);
or UO_583 (O_583,N_18888,N_18325);
or UO_584 (O_584,N_19885,N_18676);
nor UO_585 (O_585,N_18774,N_18172);
or UO_586 (O_586,N_18915,N_19362);
nor UO_587 (O_587,N_18614,N_19785);
xnor UO_588 (O_588,N_18502,N_19122);
xnor UO_589 (O_589,N_19345,N_18070);
xnor UO_590 (O_590,N_19967,N_19354);
and UO_591 (O_591,N_18405,N_19036);
or UO_592 (O_592,N_18835,N_19769);
xnor UO_593 (O_593,N_19319,N_19705);
nor UO_594 (O_594,N_19694,N_19650);
nand UO_595 (O_595,N_19022,N_18168);
and UO_596 (O_596,N_19783,N_18562);
nor UO_597 (O_597,N_19195,N_18624);
nand UO_598 (O_598,N_18841,N_19421);
nand UO_599 (O_599,N_18947,N_19620);
xor UO_600 (O_600,N_18864,N_18290);
xnor UO_601 (O_601,N_19818,N_18228);
and UO_602 (O_602,N_19350,N_18354);
nor UO_603 (O_603,N_18576,N_19698);
and UO_604 (O_604,N_18602,N_18265);
nand UO_605 (O_605,N_18752,N_18402);
nand UO_606 (O_606,N_18998,N_18195);
xnor UO_607 (O_607,N_19306,N_19594);
and UO_608 (O_608,N_19974,N_19327);
and UO_609 (O_609,N_19422,N_19524);
nand UO_610 (O_610,N_18501,N_19666);
or UO_611 (O_611,N_18207,N_19500);
nand UO_612 (O_612,N_18333,N_19270);
nand UO_613 (O_613,N_19578,N_18638);
xor UO_614 (O_614,N_19390,N_18684);
nand UO_615 (O_615,N_18124,N_19365);
xor UO_616 (O_616,N_18404,N_19108);
nand UO_617 (O_617,N_19490,N_19536);
and UO_618 (O_618,N_19496,N_19246);
and UO_619 (O_619,N_19943,N_19093);
nor UO_620 (O_620,N_18153,N_19416);
or UO_621 (O_621,N_19430,N_18832);
nand UO_622 (O_622,N_19516,N_19757);
nor UO_623 (O_623,N_18953,N_18361);
nor UO_624 (O_624,N_18690,N_19492);
or UO_625 (O_625,N_19985,N_19499);
and UO_626 (O_626,N_19872,N_19858);
nand UO_627 (O_627,N_19323,N_19013);
and UO_628 (O_628,N_19673,N_18564);
and UO_629 (O_629,N_19084,N_18555);
nand UO_630 (O_630,N_19527,N_19254);
xnor UO_631 (O_631,N_18165,N_19346);
xor UO_632 (O_632,N_19735,N_19780);
or UO_633 (O_633,N_18778,N_18563);
nor UO_634 (O_634,N_18287,N_19754);
nor UO_635 (O_635,N_19474,N_18903);
nand UO_636 (O_636,N_19277,N_18660);
xnor UO_637 (O_637,N_19837,N_19976);
and UO_638 (O_638,N_19305,N_19638);
or UO_639 (O_639,N_18604,N_19544);
nor UO_640 (O_640,N_18796,N_18646);
nor UO_641 (O_641,N_19932,N_19616);
nor UO_642 (O_642,N_18421,N_19394);
or UO_643 (O_643,N_19031,N_19432);
xor UO_644 (O_644,N_18592,N_19106);
nand UO_645 (O_645,N_19585,N_18371);
or UO_646 (O_646,N_19443,N_19979);
xor UO_647 (O_647,N_18176,N_18434);
and UO_648 (O_648,N_19295,N_19707);
or UO_649 (O_649,N_19225,N_18365);
nand UO_650 (O_650,N_19464,N_18612);
and UO_651 (O_651,N_19251,N_18593);
and UO_652 (O_652,N_19540,N_18967);
nand UO_653 (O_653,N_19796,N_18403);
and UO_654 (O_654,N_18246,N_18148);
nand UO_655 (O_655,N_19234,N_19807);
or UO_656 (O_656,N_18279,N_19518);
nor UO_657 (O_657,N_18318,N_19678);
or UO_658 (O_658,N_19649,N_18358);
or UO_659 (O_659,N_18834,N_18569);
or UO_660 (O_660,N_18821,N_19227);
and UO_661 (O_661,N_19865,N_18530);
or UO_662 (O_662,N_18142,N_19398);
or UO_663 (O_663,N_19954,N_18889);
nor UO_664 (O_664,N_19006,N_19241);
and UO_665 (O_665,N_18335,N_18081);
and UO_666 (O_666,N_19790,N_19489);
nand UO_667 (O_667,N_18940,N_19654);
xnor UO_668 (O_668,N_19576,N_18495);
nand UO_669 (O_669,N_19770,N_18984);
nor UO_670 (O_670,N_19853,N_18223);
nand UO_671 (O_671,N_19696,N_18876);
or UO_672 (O_672,N_19589,N_18141);
and UO_673 (O_673,N_18487,N_18987);
or UO_674 (O_674,N_19877,N_19090);
nor UO_675 (O_675,N_18300,N_18785);
or UO_676 (O_676,N_18656,N_19996);
xor UO_677 (O_677,N_19572,N_18791);
nand UO_678 (O_678,N_18797,N_19625);
nor UO_679 (O_679,N_18741,N_19793);
and UO_680 (O_680,N_19282,N_19835);
xor UO_681 (O_681,N_19008,N_19173);
and UO_682 (O_682,N_19875,N_18190);
xnor UO_683 (O_683,N_18263,N_18044);
xor UO_684 (O_684,N_19411,N_18585);
or UO_685 (O_685,N_19307,N_19587);
and UO_686 (O_686,N_19523,N_18174);
xnor UO_687 (O_687,N_18471,N_18605);
xnor UO_688 (O_688,N_18167,N_18678);
and UO_689 (O_689,N_19874,N_19448);
xor UO_690 (O_690,N_19631,N_19520);
nand UO_691 (O_691,N_18486,N_18776);
nand UO_692 (O_692,N_19549,N_18863);
and UO_693 (O_693,N_19003,N_18019);
nor UO_694 (O_694,N_19661,N_19210);
or UO_695 (O_695,N_18459,N_19801);
nor UO_696 (O_696,N_18707,N_19668);
nand UO_697 (O_697,N_18181,N_19902);
xor UO_698 (O_698,N_19309,N_18649);
and UO_699 (O_699,N_18099,N_19911);
nand UO_700 (O_700,N_18312,N_18134);
xnor UO_701 (O_701,N_19613,N_18567);
or UO_702 (O_702,N_18357,N_19652);
nand UO_703 (O_703,N_19061,N_18846);
nand UO_704 (O_704,N_18169,N_18780);
nand UO_705 (O_705,N_19399,N_19188);
or UO_706 (O_706,N_18129,N_18539);
and UO_707 (O_707,N_18622,N_19588);
nand UO_708 (O_708,N_19030,N_19478);
or UO_709 (O_709,N_19653,N_19068);
nor UO_710 (O_710,N_19598,N_19849);
or UO_711 (O_711,N_19194,N_18309);
xnor UO_712 (O_712,N_18650,N_18554);
xnor UO_713 (O_713,N_19491,N_19040);
xnor UO_714 (O_714,N_19079,N_18249);
xnor UO_715 (O_715,N_19343,N_19101);
and UO_716 (O_716,N_19535,N_19659);
xor UO_717 (O_717,N_19117,N_18619);
nand UO_718 (O_718,N_18233,N_18877);
nand UO_719 (O_719,N_18932,N_19806);
and UO_720 (O_720,N_19174,N_19561);
and UO_721 (O_721,N_19883,N_18256);
and UO_722 (O_722,N_18496,N_19786);
nand UO_723 (O_723,N_18838,N_18618);
or UO_724 (O_724,N_19991,N_19331);
xnor UO_725 (O_725,N_19301,N_18992);
nor UO_726 (O_726,N_18693,N_18024);
nor UO_727 (O_727,N_18242,N_19048);
nand UO_728 (O_728,N_19482,N_19526);
xnor UO_729 (O_729,N_19318,N_18701);
or UO_730 (O_730,N_18122,N_18074);
nor UO_731 (O_731,N_19811,N_18166);
nor UO_732 (O_732,N_18069,N_18262);
nor UO_733 (O_733,N_19618,N_18171);
xnor UO_734 (O_734,N_18894,N_18426);
nand UO_735 (O_735,N_19961,N_19088);
nor UO_736 (O_736,N_18010,N_19320);
nand UO_737 (O_737,N_19185,N_19758);
or UO_738 (O_738,N_19823,N_19914);
xor UO_739 (O_739,N_18634,N_19922);
and UO_740 (O_740,N_19025,N_19580);
nor UO_741 (O_741,N_18058,N_19640);
nand UO_742 (O_742,N_18057,N_19881);
nand UO_743 (O_743,N_19033,N_18250);
or UO_744 (O_744,N_19112,N_19475);
nand UO_745 (O_745,N_18580,N_19554);
or UO_746 (O_746,N_19435,N_19688);
and UO_747 (O_747,N_19714,N_19599);
and UO_748 (O_748,N_19401,N_19686);
nor UO_749 (O_749,N_18928,N_19633);
and UO_750 (O_750,N_19224,N_18945);
and UO_751 (O_751,N_18615,N_18935);
nand UO_752 (O_752,N_18109,N_19207);
and UO_753 (O_753,N_18106,N_19175);
nor UO_754 (O_754,N_19798,N_18545);
and UO_755 (O_755,N_19953,N_19511);
or UO_756 (O_756,N_18478,N_19400);
or UO_757 (O_757,N_19564,N_19550);
nor UO_758 (O_758,N_19750,N_18418);
nand UO_759 (O_759,N_18830,N_18359);
or UO_760 (O_760,N_18897,N_19237);
xnor UO_761 (O_761,N_19149,N_18816);
xor UO_762 (O_762,N_19730,N_19042);
nor UO_763 (O_763,N_18775,N_19936);
xnor UO_764 (O_764,N_19992,N_19466);
or UO_765 (O_765,N_19348,N_19998);
or UO_766 (O_766,N_19683,N_18323);
xor UO_767 (O_767,N_18053,N_19803);
nand UO_768 (O_768,N_19609,N_19388);
and UO_769 (O_769,N_18651,N_18696);
and UO_770 (O_770,N_18383,N_18466);
nor UO_771 (O_771,N_19782,N_18338);
and UO_772 (O_772,N_19514,N_18216);
xnor UO_773 (O_773,N_19417,N_18098);
nor UO_774 (O_774,N_19330,N_18811);
nor UO_775 (O_775,N_19052,N_19660);
xor UO_776 (O_776,N_18765,N_18740);
nand UO_777 (O_777,N_18393,N_18974);
and UO_778 (O_778,N_19403,N_19340);
xnor UO_779 (O_779,N_18211,N_18611);
nor UO_780 (O_780,N_19405,N_18015);
nand UO_781 (O_781,N_18972,N_19746);
xnor UO_782 (O_782,N_18028,N_18753);
or UO_783 (O_783,N_18500,N_18248);
and UO_784 (O_784,N_19808,N_19361);
xor UO_785 (O_785,N_19308,N_18995);
nor UO_786 (O_786,N_19433,N_18490);
and UO_787 (O_787,N_18767,N_18105);
and UO_788 (O_788,N_19804,N_19131);
xor UO_789 (O_789,N_19437,N_19759);
xor UO_790 (O_790,N_18206,N_19844);
and UO_791 (O_791,N_18789,N_19647);
or UO_792 (O_792,N_19387,N_19165);
and UO_793 (O_793,N_19761,N_19530);
nand UO_794 (O_794,N_18100,N_19715);
nor UO_795 (O_795,N_19723,N_19367);
or UO_796 (O_796,N_19477,N_19322);
nor UO_797 (O_797,N_18347,N_18151);
and UO_798 (O_798,N_18322,N_18819);
and UO_799 (O_799,N_18529,N_19845);
nand UO_800 (O_800,N_18021,N_19057);
or UO_801 (O_801,N_19543,N_19890);
nor UO_802 (O_802,N_19716,N_19262);
or UO_803 (O_803,N_19344,N_19857);
nor UO_804 (O_804,N_18931,N_19215);
or UO_805 (O_805,N_19452,N_18517);
xnor UO_806 (O_806,N_18451,N_18283);
or UO_807 (O_807,N_19509,N_18794);
or UO_808 (O_808,N_19135,N_19235);
and UO_809 (O_809,N_18481,N_18253);
nor UO_810 (O_810,N_18851,N_18157);
or UO_811 (O_811,N_19745,N_18214);
nand UO_812 (O_812,N_19924,N_18871);
xor UO_813 (O_813,N_19828,N_19918);
nor UO_814 (O_814,N_19171,N_19379);
and UO_815 (O_815,N_19451,N_19484);
nor UO_816 (O_816,N_18670,N_19434);
nand UO_817 (O_817,N_18472,N_19958);
nand UO_818 (O_818,N_18280,N_19634);
and UO_819 (O_819,N_18506,N_19021);
and UO_820 (O_820,N_19864,N_18161);
nor UO_821 (O_821,N_18823,N_19983);
and UO_822 (O_822,N_19024,N_18694);
or UO_823 (O_823,N_18803,N_18533);
nand UO_824 (O_824,N_18662,N_19232);
or UO_825 (O_825,N_19724,N_18887);
nand UO_826 (O_826,N_18022,N_19444);
or UO_827 (O_827,N_18745,N_18672);
nand UO_828 (O_828,N_19209,N_19353);
nand UO_829 (O_829,N_19838,N_19889);
nor UO_830 (O_830,N_18837,N_19941);
nand UO_831 (O_831,N_19476,N_19632);
nand UO_832 (O_832,N_19762,N_18599);
or UO_833 (O_833,N_18966,N_18836);
nor UO_834 (O_834,N_18485,N_18060);
and UO_835 (O_835,N_18756,N_19017);
nand UO_836 (O_836,N_18349,N_19920);
xnor UO_837 (O_837,N_18732,N_18924);
xor UO_838 (O_838,N_19948,N_18522);
xor UO_839 (O_839,N_18532,N_18726);
nor UO_840 (O_840,N_18447,N_19658);
nor UO_841 (O_841,N_18779,N_18008);
and UO_842 (O_842,N_19963,N_18633);
or UO_843 (O_843,N_18598,N_19086);
xor UO_844 (O_844,N_19469,N_18628);
and UO_845 (O_845,N_19214,N_19183);
or UO_846 (O_846,N_19383,N_19854);
or UO_847 (O_847,N_19859,N_18594);
or UO_848 (O_848,N_18919,N_19656);
nand UO_849 (O_849,N_18125,N_19870);
xor UO_850 (O_850,N_19584,N_19223);
and UO_851 (O_851,N_18963,N_19198);
nand UO_852 (O_852,N_19111,N_19517);
nor UO_853 (O_853,N_18126,N_18006);
and UO_854 (O_854,N_19900,N_18225);
xnor UO_855 (O_855,N_19115,N_18107);
nor UO_856 (O_856,N_19358,N_19304);
nor UO_857 (O_857,N_18473,N_18930);
nor UO_858 (O_858,N_19473,N_18210);
and UO_859 (O_859,N_19371,N_18787);
or UO_860 (O_860,N_18468,N_19701);
and UO_861 (O_861,N_18980,N_18844);
nor UO_862 (O_862,N_18240,N_19987);
nor UO_863 (O_863,N_19104,N_18550);
and UO_864 (O_864,N_19856,N_18747);
or UO_865 (O_865,N_18091,N_19689);
or UO_866 (O_866,N_19329,N_18730);
and UO_867 (O_867,N_18891,N_19010);
or UO_868 (O_868,N_18907,N_18143);
and UO_869 (O_869,N_19032,N_18959);
or UO_870 (O_870,N_19619,N_18480);
nor UO_871 (O_871,N_18711,N_18399);
and UO_872 (O_872,N_19830,N_18238);
xnor UO_873 (O_873,N_18538,N_19614);
and UO_874 (O_874,N_18222,N_18659);
or UO_875 (O_875,N_19230,N_18826);
nor UO_876 (O_876,N_18536,N_18766);
and UO_877 (O_877,N_18296,N_19919);
and UO_878 (O_878,N_19608,N_19087);
nand UO_879 (O_879,N_18729,N_18492);
nor UO_880 (O_880,N_18802,N_19797);
xnor UO_881 (O_881,N_19753,N_19583);
xnor UO_882 (O_882,N_19290,N_18691);
nor UO_883 (O_883,N_19357,N_18462);
or UO_884 (O_884,N_19646,N_19657);
nor UO_885 (O_885,N_18198,N_19454);
nand UO_886 (O_886,N_18685,N_18110);
xor UO_887 (O_887,N_18121,N_18996);
nor UO_888 (O_888,N_19193,N_18962);
nand UO_889 (O_889,N_18033,N_18658);
xor UO_890 (O_890,N_18654,N_18237);
and UO_891 (O_891,N_18112,N_19192);
and UO_892 (O_892,N_19385,N_19766);
nor UO_893 (O_893,N_19281,N_19316);
nor UO_894 (O_894,N_18806,N_18825);
xor UO_895 (O_895,N_19777,N_19711);
nand UO_896 (O_896,N_19483,N_19296);
nand UO_897 (O_897,N_19143,N_18272);
or UO_898 (O_898,N_19324,N_18064);
nand UO_899 (O_899,N_18526,N_18872);
or UO_900 (O_900,N_19181,N_18695);
nor UO_901 (O_901,N_18664,N_18150);
nand UO_902 (O_902,N_18866,N_18590);
or UO_903 (O_903,N_18366,N_19255);
and UO_904 (O_904,N_19419,N_18449);
or UO_905 (O_905,N_18750,N_19817);
and UO_906 (O_906,N_18509,N_19971);
nor UO_907 (O_907,N_18209,N_19205);
and UO_908 (O_908,N_18801,N_18456);
xnor UO_909 (O_909,N_18097,N_19118);
nor UO_910 (O_910,N_19813,N_19639);
nor UO_911 (O_911,N_18367,N_19272);
nand UO_912 (O_912,N_19846,N_18493);
or UO_913 (O_913,N_19643,N_19313);
nor UO_914 (O_914,N_19781,N_18822);
or UO_915 (O_915,N_19834,N_18868);
nor UO_916 (O_916,N_19692,N_19364);
nor UO_917 (O_917,N_18316,N_19238);
or UO_918 (O_918,N_18477,N_18294);
nor UO_919 (O_919,N_19718,N_19078);
nor UO_920 (O_920,N_18892,N_19725);
or UO_921 (O_921,N_19189,N_19257);
nor UO_922 (O_922,N_19876,N_18883);
xor UO_923 (O_923,N_19420,N_18398);
and UO_924 (O_924,N_18748,N_18232);
nand UO_925 (O_925,N_18011,N_19720);
and UO_926 (O_926,N_18665,N_18469);
nor UO_927 (O_927,N_19054,N_18900);
and UO_928 (O_928,N_19802,N_19266);
nand UO_929 (O_929,N_19132,N_19269);
xnor UO_930 (O_930,N_19791,N_19573);
and UO_931 (O_931,N_19457,N_19038);
nand UO_932 (O_932,N_18187,N_19128);
and UO_933 (O_933,N_18131,N_19717);
and UO_934 (O_934,N_18853,N_18363);
xor UO_935 (O_935,N_18295,N_19298);
nor UO_936 (O_936,N_18292,N_18975);
xnor UO_937 (O_937,N_19127,N_18465);
nand UO_938 (O_938,N_19574,N_19568);
nor UO_939 (O_939,N_18247,N_19871);
nand UO_940 (O_940,N_18281,N_19907);
and UO_941 (O_941,N_19916,N_19863);
nand UO_942 (O_942,N_18470,N_18666);
and UO_943 (O_943,N_19559,N_18927);
nand UO_944 (O_944,N_18899,N_18706);
xnor UO_945 (O_945,N_18407,N_18781);
xor UO_946 (O_946,N_18392,N_19852);
xnor UO_947 (O_947,N_19034,N_18810);
nor UO_948 (O_948,N_19249,N_19947);
and UO_949 (O_949,N_18800,N_18904);
nor UO_950 (O_950,N_19860,N_19442);
nand UO_951 (O_951,N_19072,N_19959);
xor UO_952 (O_952,N_18259,N_19382);
nand UO_953 (O_953,N_19925,N_18433);
xnor UO_954 (O_954,N_19831,N_18528);
and UO_955 (O_955,N_18777,N_19832);
nor UO_956 (O_956,N_18430,N_18640);
nand UO_957 (O_957,N_19325,N_18683);
and UO_958 (O_958,N_18942,N_19130);
and UO_959 (O_959,N_18663,N_18196);
nor UO_960 (O_960,N_19035,N_18905);
xor UO_961 (O_961,N_19005,N_19704);
nor UO_962 (O_962,N_19605,N_19148);
or UO_963 (O_963,N_18988,N_19083);
and UO_964 (O_964,N_18620,N_19910);
nand UO_965 (O_965,N_19565,N_19386);
xnor UO_966 (O_966,N_18571,N_19510);
nor UO_967 (O_967,N_19310,N_19508);
nor UO_968 (O_968,N_18723,N_19150);
nand UO_969 (O_969,N_18999,N_19231);
or UO_970 (O_970,N_18589,N_18314);
xor UO_971 (O_971,N_19060,N_19600);
nand UO_972 (O_972,N_18828,N_18630);
and UO_973 (O_973,N_18269,N_18163);
and UO_974 (O_974,N_18062,N_19252);
or UO_975 (O_975,N_18364,N_18973);
xor UO_976 (O_976,N_19431,N_19977);
xnor UO_977 (O_977,N_18217,N_18376);
nand UO_978 (O_978,N_19092,N_19973);
xor UO_979 (O_979,N_18770,N_18771);
xnor UO_980 (O_980,N_19525,N_19248);
nand UO_981 (O_981,N_18356,N_19538);
and UO_982 (O_982,N_19113,N_18716);
nand UO_983 (O_983,N_19439,N_19071);
nand UO_984 (O_984,N_19020,N_18360);
or UO_985 (O_985,N_19016,N_18324);
and UO_986 (O_986,N_19779,N_18704);
xor UO_987 (O_987,N_19355,N_19328);
nor UO_988 (O_988,N_18437,N_18954);
nand UO_989 (O_989,N_18964,N_18627);
nor UO_990 (O_990,N_18303,N_19548);
nor UO_991 (O_991,N_19679,N_18523);
xor UO_992 (O_992,N_19611,N_18088);
nand UO_993 (O_993,N_18120,N_18175);
xnor UO_994 (O_994,N_19939,N_19263);
nor UO_995 (O_995,N_18510,N_19986);
and UO_996 (O_996,N_18687,N_18378);
and UO_997 (O_997,N_19655,N_18156);
or UO_998 (O_998,N_18197,N_18442);
nor UO_999 (O_999,N_18632,N_18203);
nand UO_1000 (O_1000,N_18827,N_19527);
nor UO_1001 (O_1001,N_18445,N_19354);
xnor UO_1002 (O_1002,N_19895,N_18551);
xor UO_1003 (O_1003,N_18073,N_19169);
and UO_1004 (O_1004,N_18729,N_19547);
and UO_1005 (O_1005,N_19857,N_18666);
xnor UO_1006 (O_1006,N_18398,N_19861);
xnor UO_1007 (O_1007,N_19532,N_19302);
nand UO_1008 (O_1008,N_19105,N_18350);
nand UO_1009 (O_1009,N_19037,N_19649);
and UO_1010 (O_1010,N_19502,N_19374);
or UO_1011 (O_1011,N_18633,N_18653);
or UO_1012 (O_1012,N_19909,N_18158);
and UO_1013 (O_1013,N_18561,N_19246);
nor UO_1014 (O_1014,N_18763,N_19617);
and UO_1015 (O_1015,N_18697,N_19502);
xnor UO_1016 (O_1016,N_19384,N_19556);
and UO_1017 (O_1017,N_18930,N_19585);
xor UO_1018 (O_1018,N_18139,N_19910);
and UO_1019 (O_1019,N_18410,N_19077);
nand UO_1020 (O_1020,N_19020,N_18061);
nor UO_1021 (O_1021,N_18369,N_18197);
nor UO_1022 (O_1022,N_18319,N_19939);
or UO_1023 (O_1023,N_19723,N_19713);
and UO_1024 (O_1024,N_19754,N_19391);
nor UO_1025 (O_1025,N_19034,N_18241);
nand UO_1026 (O_1026,N_19330,N_18836);
or UO_1027 (O_1027,N_18223,N_18347);
nor UO_1028 (O_1028,N_19578,N_18442);
nand UO_1029 (O_1029,N_18129,N_18501);
nand UO_1030 (O_1030,N_18643,N_19074);
xnor UO_1031 (O_1031,N_19879,N_18955);
or UO_1032 (O_1032,N_18093,N_19340);
nand UO_1033 (O_1033,N_19270,N_19383);
xnor UO_1034 (O_1034,N_19633,N_19909);
xnor UO_1035 (O_1035,N_18336,N_18563);
and UO_1036 (O_1036,N_18266,N_19394);
or UO_1037 (O_1037,N_18362,N_19105);
nor UO_1038 (O_1038,N_19774,N_19652);
nand UO_1039 (O_1039,N_18054,N_18281);
and UO_1040 (O_1040,N_18488,N_18289);
nor UO_1041 (O_1041,N_18956,N_19187);
nor UO_1042 (O_1042,N_18499,N_19513);
or UO_1043 (O_1043,N_19274,N_18128);
or UO_1044 (O_1044,N_19834,N_18822);
or UO_1045 (O_1045,N_19976,N_19009);
or UO_1046 (O_1046,N_19431,N_19947);
and UO_1047 (O_1047,N_18617,N_18933);
nor UO_1048 (O_1048,N_18777,N_19057);
nand UO_1049 (O_1049,N_18196,N_19426);
and UO_1050 (O_1050,N_19323,N_18572);
xnor UO_1051 (O_1051,N_18733,N_18683);
and UO_1052 (O_1052,N_19922,N_18191);
xnor UO_1053 (O_1053,N_18066,N_18646);
nor UO_1054 (O_1054,N_18577,N_19202);
or UO_1055 (O_1055,N_18936,N_19781);
nand UO_1056 (O_1056,N_19315,N_19939);
or UO_1057 (O_1057,N_19554,N_18819);
nand UO_1058 (O_1058,N_18232,N_19231);
and UO_1059 (O_1059,N_18446,N_19279);
nand UO_1060 (O_1060,N_18501,N_19047);
nor UO_1061 (O_1061,N_19450,N_18837);
nand UO_1062 (O_1062,N_18573,N_18288);
or UO_1063 (O_1063,N_19293,N_19567);
nand UO_1064 (O_1064,N_18520,N_18875);
or UO_1065 (O_1065,N_18448,N_19697);
and UO_1066 (O_1066,N_18448,N_18534);
nand UO_1067 (O_1067,N_18350,N_18071);
or UO_1068 (O_1068,N_19040,N_18214);
or UO_1069 (O_1069,N_18477,N_19616);
xnor UO_1070 (O_1070,N_18059,N_18860);
nor UO_1071 (O_1071,N_19439,N_18836);
and UO_1072 (O_1072,N_18550,N_19433);
and UO_1073 (O_1073,N_18325,N_18289);
and UO_1074 (O_1074,N_19444,N_19937);
or UO_1075 (O_1075,N_19772,N_19646);
or UO_1076 (O_1076,N_19334,N_19322);
nand UO_1077 (O_1077,N_18815,N_18607);
nand UO_1078 (O_1078,N_18731,N_19566);
nor UO_1079 (O_1079,N_18057,N_18527);
nand UO_1080 (O_1080,N_18903,N_18332);
or UO_1081 (O_1081,N_19421,N_19801);
nor UO_1082 (O_1082,N_18576,N_18411);
nor UO_1083 (O_1083,N_18719,N_19180);
xnor UO_1084 (O_1084,N_18511,N_19366);
and UO_1085 (O_1085,N_18760,N_19264);
xnor UO_1086 (O_1086,N_19943,N_18009);
xnor UO_1087 (O_1087,N_19766,N_19047);
and UO_1088 (O_1088,N_18022,N_18874);
nor UO_1089 (O_1089,N_18047,N_18976);
nand UO_1090 (O_1090,N_18094,N_18447);
and UO_1091 (O_1091,N_18808,N_18720);
nand UO_1092 (O_1092,N_18360,N_19523);
nor UO_1093 (O_1093,N_18197,N_19009);
and UO_1094 (O_1094,N_18792,N_19924);
or UO_1095 (O_1095,N_18905,N_19800);
or UO_1096 (O_1096,N_18509,N_18523);
nand UO_1097 (O_1097,N_18240,N_18420);
and UO_1098 (O_1098,N_18566,N_19168);
and UO_1099 (O_1099,N_18658,N_18647);
or UO_1100 (O_1100,N_18072,N_19506);
xnor UO_1101 (O_1101,N_18051,N_18875);
xnor UO_1102 (O_1102,N_19214,N_19228);
and UO_1103 (O_1103,N_18232,N_19447);
xor UO_1104 (O_1104,N_18647,N_18858);
nor UO_1105 (O_1105,N_19510,N_19268);
and UO_1106 (O_1106,N_19450,N_19644);
nor UO_1107 (O_1107,N_18231,N_19010);
xor UO_1108 (O_1108,N_18266,N_19225);
and UO_1109 (O_1109,N_19430,N_18193);
or UO_1110 (O_1110,N_19901,N_19538);
xnor UO_1111 (O_1111,N_18609,N_18516);
and UO_1112 (O_1112,N_19008,N_18917);
and UO_1113 (O_1113,N_19745,N_19453);
and UO_1114 (O_1114,N_18923,N_19266);
nand UO_1115 (O_1115,N_19610,N_18867);
and UO_1116 (O_1116,N_19016,N_19727);
and UO_1117 (O_1117,N_19576,N_18606);
and UO_1118 (O_1118,N_19045,N_18057);
xor UO_1119 (O_1119,N_19069,N_19617);
nor UO_1120 (O_1120,N_18919,N_18003);
nor UO_1121 (O_1121,N_19355,N_18233);
or UO_1122 (O_1122,N_19320,N_19031);
xor UO_1123 (O_1123,N_18450,N_19632);
or UO_1124 (O_1124,N_18302,N_19576);
and UO_1125 (O_1125,N_19243,N_19857);
nor UO_1126 (O_1126,N_18965,N_18926);
xnor UO_1127 (O_1127,N_19553,N_18144);
and UO_1128 (O_1128,N_18284,N_19027);
nand UO_1129 (O_1129,N_19648,N_18248);
or UO_1130 (O_1130,N_19611,N_19839);
xnor UO_1131 (O_1131,N_19574,N_19174);
or UO_1132 (O_1132,N_18392,N_19663);
or UO_1133 (O_1133,N_19602,N_18029);
and UO_1134 (O_1134,N_18636,N_19460);
or UO_1135 (O_1135,N_19956,N_19154);
nand UO_1136 (O_1136,N_18757,N_18729);
nor UO_1137 (O_1137,N_19382,N_19248);
xnor UO_1138 (O_1138,N_19425,N_18305);
nand UO_1139 (O_1139,N_19861,N_18782);
nand UO_1140 (O_1140,N_18195,N_19773);
nor UO_1141 (O_1141,N_19842,N_19376);
xnor UO_1142 (O_1142,N_19270,N_19622);
nor UO_1143 (O_1143,N_19520,N_19326);
nand UO_1144 (O_1144,N_19787,N_18778);
xnor UO_1145 (O_1145,N_18013,N_19452);
or UO_1146 (O_1146,N_19462,N_18452);
nor UO_1147 (O_1147,N_19573,N_18308);
xnor UO_1148 (O_1148,N_18670,N_19495);
and UO_1149 (O_1149,N_19186,N_18710);
xor UO_1150 (O_1150,N_18462,N_18517);
nor UO_1151 (O_1151,N_18700,N_19737);
nand UO_1152 (O_1152,N_19711,N_18357);
xor UO_1153 (O_1153,N_19059,N_18420);
and UO_1154 (O_1154,N_18613,N_18086);
nor UO_1155 (O_1155,N_19487,N_18791);
or UO_1156 (O_1156,N_18829,N_18564);
xor UO_1157 (O_1157,N_19371,N_18544);
nand UO_1158 (O_1158,N_18496,N_19925);
nor UO_1159 (O_1159,N_19308,N_19339);
nand UO_1160 (O_1160,N_19187,N_19149);
or UO_1161 (O_1161,N_18941,N_18472);
and UO_1162 (O_1162,N_18353,N_18167);
nand UO_1163 (O_1163,N_19254,N_19100);
and UO_1164 (O_1164,N_18184,N_18984);
nor UO_1165 (O_1165,N_18462,N_18101);
xor UO_1166 (O_1166,N_18126,N_19185);
or UO_1167 (O_1167,N_18548,N_19912);
nor UO_1168 (O_1168,N_18848,N_18651);
and UO_1169 (O_1169,N_18698,N_18995);
xor UO_1170 (O_1170,N_18346,N_18757);
and UO_1171 (O_1171,N_19337,N_19134);
nor UO_1172 (O_1172,N_18085,N_18915);
nand UO_1173 (O_1173,N_19552,N_18677);
or UO_1174 (O_1174,N_18778,N_19594);
nor UO_1175 (O_1175,N_19061,N_19886);
nand UO_1176 (O_1176,N_18567,N_18339);
nand UO_1177 (O_1177,N_19463,N_19576);
nor UO_1178 (O_1178,N_18394,N_19047);
and UO_1179 (O_1179,N_18083,N_19922);
or UO_1180 (O_1180,N_18505,N_18016);
nand UO_1181 (O_1181,N_18888,N_18193);
or UO_1182 (O_1182,N_18259,N_19829);
nor UO_1183 (O_1183,N_18885,N_19242);
nor UO_1184 (O_1184,N_19957,N_19547);
or UO_1185 (O_1185,N_19433,N_19477);
nor UO_1186 (O_1186,N_19145,N_19569);
xor UO_1187 (O_1187,N_18630,N_19905);
xnor UO_1188 (O_1188,N_18837,N_19650);
and UO_1189 (O_1189,N_18570,N_19719);
xnor UO_1190 (O_1190,N_19297,N_18854);
and UO_1191 (O_1191,N_18822,N_18792);
nand UO_1192 (O_1192,N_19648,N_18400);
and UO_1193 (O_1193,N_19398,N_18573);
or UO_1194 (O_1194,N_19382,N_19068);
nor UO_1195 (O_1195,N_19087,N_18458);
and UO_1196 (O_1196,N_18130,N_18022);
and UO_1197 (O_1197,N_19839,N_18136);
nand UO_1198 (O_1198,N_19008,N_18679);
xor UO_1199 (O_1199,N_19817,N_19427);
xor UO_1200 (O_1200,N_18923,N_19822);
xnor UO_1201 (O_1201,N_19228,N_18342);
nand UO_1202 (O_1202,N_18906,N_18078);
or UO_1203 (O_1203,N_19493,N_18098);
or UO_1204 (O_1204,N_18197,N_18861);
nand UO_1205 (O_1205,N_18559,N_18437);
or UO_1206 (O_1206,N_18770,N_19786);
nor UO_1207 (O_1207,N_18011,N_19520);
xor UO_1208 (O_1208,N_18314,N_18891);
nor UO_1209 (O_1209,N_18303,N_19277);
and UO_1210 (O_1210,N_19666,N_18498);
nand UO_1211 (O_1211,N_18174,N_18438);
or UO_1212 (O_1212,N_18155,N_19982);
or UO_1213 (O_1213,N_18620,N_19348);
nand UO_1214 (O_1214,N_18836,N_19224);
xor UO_1215 (O_1215,N_18098,N_19603);
xor UO_1216 (O_1216,N_18606,N_18985);
nand UO_1217 (O_1217,N_19533,N_19157);
nor UO_1218 (O_1218,N_19767,N_18461);
or UO_1219 (O_1219,N_19790,N_19595);
or UO_1220 (O_1220,N_18153,N_19184);
xnor UO_1221 (O_1221,N_19525,N_19004);
xnor UO_1222 (O_1222,N_19424,N_18121);
nor UO_1223 (O_1223,N_18653,N_18802);
xnor UO_1224 (O_1224,N_19200,N_18138);
xnor UO_1225 (O_1225,N_18414,N_18154);
or UO_1226 (O_1226,N_19257,N_18850);
and UO_1227 (O_1227,N_19902,N_19615);
xnor UO_1228 (O_1228,N_18116,N_18182);
nor UO_1229 (O_1229,N_18632,N_18162);
or UO_1230 (O_1230,N_18388,N_19410);
nand UO_1231 (O_1231,N_18434,N_18254);
nor UO_1232 (O_1232,N_19414,N_19250);
nor UO_1233 (O_1233,N_19756,N_18800);
nand UO_1234 (O_1234,N_18646,N_18072);
nand UO_1235 (O_1235,N_18422,N_18781);
and UO_1236 (O_1236,N_19162,N_19327);
nand UO_1237 (O_1237,N_19678,N_18545);
nand UO_1238 (O_1238,N_19302,N_19373);
xnor UO_1239 (O_1239,N_19388,N_18181);
xnor UO_1240 (O_1240,N_19037,N_18401);
and UO_1241 (O_1241,N_18726,N_18319);
or UO_1242 (O_1242,N_18030,N_19394);
and UO_1243 (O_1243,N_18050,N_19138);
nand UO_1244 (O_1244,N_19969,N_19431);
nand UO_1245 (O_1245,N_19662,N_19953);
xor UO_1246 (O_1246,N_18126,N_19869);
nor UO_1247 (O_1247,N_19280,N_19519);
and UO_1248 (O_1248,N_19672,N_19969);
or UO_1249 (O_1249,N_18258,N_19061);
or UO_1250 (O_1250,N_18141,N_19178);
xnor UO_1251 (O_1251,N_18033,N_19375);
nand UO_1252 (O_1252,N_19381,N_19634);
nand UO_1253 (O_1253,N_19126,N_18055);
and UO_1254 (O_1254,N_18884,N_18348);
or UO_1255 (O_1255,N_19862,N_19409);
nand UO_1256 (O_1256,N_19214,N_19368);
xor UO_1257 (O_1257,N_19327,N_19924);
nand UO_1258 (O_1258,N_18412,N_18920);
xor UO_1259 (O_1259,N_19114,N_18543);
nor UO_1260 (O_1260,N_18426,N_18112);
nor UO_1261 (O_1261,N_19451,N_18828);
xor UO_1262 (O_1262,N_19624,N_18058);
and UO_1263 (O_1263,N_19426,N_18547);
xor UO_1264 (O_1264,N_19897,N_18518);
nand UO_1265 (O_1265,N_19446,N_18529);
nor UO_1266 (O_1266,N_19477,N_19367);
nor UO_1267 (O_1267,N_19551,N_19310);
nand UO_1268 (O_1268,N_19361,N_18465);
nor UO_1269 (O_1269,N_19356,N_19744);
or UO_1270 (O_1270,N_18023,N_18019);
or UO_1271 (O_1271,N_19006,N_19272);
nand UO_1272 (O_1272,N_18255,N_19586);
or UO_1273 (O_1273,N_19360,N_18916);
nand UO_1274 (O_1274,N_19855,N_18808);
nand UO_1275 (O_1275,N_18597,N_19201);
and UO_1276 (O_1276,N_19425,N_18688);
or UO_1277 (O_1277,N_18483,N_19115);
nand UO_1278 (O_1278,N_18715,N_18248);
xor UO_1279 (O_1279,N_19221,N_19760);
and UO_1280 (O_1280,N_18516,N_19143);
or UO_1281 (O_1281,N_19687,N_19118);
nand UO_1282 (O_1282,N_19323,N_19862);
nor UO_1283 (O_1283,N_18681,N_18646);
and UO_1284 (O_1284,N_18665,N_19756);
nor UO_1285 (O_1285,N_18001,N_18591);
nand UO_1286 (O_1286,N_19260,N_19473);
nand UO_1287 (O_1287,N_19306,N_19084);
and UO_1288 (O_1288,N_18648,N_19095);
xnor UO_1289 (O_1289,N_19239,N_19552);
nand UO_1290 (O_1290,N_18529,N_19641);
and UO_1291 (O_1291,N_18450,N_18469);
nand UO_1292 (O_1292,N_19666,N_19198);
and UO_1293 (O_1293,N_18633,N_18398);
nor UO_1294 (O_1294,N_19191,N_19122);
or UO_1295 (O_1295,N_19115,N_18818);
xor UO_1296 (O_1296,N_19125,N_19795);
nand UO_1297 (O_1297,N_19734,N_18512);
and UO_1298 (O_1298,N_18957,N_18481);
nand UO_1299 (O_1299,N_18328,N_19938);
xnor UO_1300 (O_1300,N_18813,N_19764);
or UO_1301 (O_1301,N_19948,N_19517);
nor UO_1302 (O_1302,N_19467,N_18100);
nand UO_1303 (O_1303,N_18000,N_18870);
and UO_1304 (O_1304,N_19559,N_18170);
nor UO_1305 (O_1305,N_19598,N_18499);
or UO_1306 (O_1306,N_18560,N_18526);
xor UO_1307 (O_1307,N_18100,N_18672);
or UO_1308 (O_1308,N_19870,N_19938);
nand UO_1309 (O_1309,N_19791,N_18468);
or UO_1310 (O_1310,N_19630,N_18063);
nand UO_1311 (O_1311,N_19670,N_18018);
nand UO_1312 (O_1312,N_19292,N_18553);
xnor UO_1313 (O_1313,N_18394,N_18401);
and UO_1314 (O_1314,N_18856,N_18375);
or UO_1315 (O_1315,N_18560,N_18476);
xnor UO_1316 (O_1316,N_18568,N_18244);
or UO_1317 (O_1317,N_19629,N_18842);
or UO_1318 (O_1318,N_19504,N_18088);
nand UO_1319 (O_1319,N_19390,N_18909);
nand UO_1320 (O_1320,N_18047,N_19929);
xor UO_1321 (O_1321,N_19746,N_19429);
nor UO_1322 (O_1322,N_19895,N_19466);
nand UO_1323 (O_1323,N_19303,N_18088);
nor UO_1324 (O_1324,N_19737,N_19658);
xor UO_1325 (O_1325,N_19525,N_18881);
xor UO_1326 (O_1326,N_19263,N_18775);
nand UO_1327 (O_1327,N_18164,N_19951);
xor UO_1328 (O_1328,N_19942,N_18774);
or UO_1329 (O_1329,N_19657,N_18331);
nor UO_1330 (O_1330,N_18604,N_19540);
nand UO_1331 (O_1331,N_19739,N_18436);
or UO_1332 (O_1332,N_18235,N_19432);
nor UO_1333 (O_1333,N_19076,N_19402);
nand UO_1334 (O_1334,N_19285,N_18597);
nand UO_1335 (O_1335,N_19541,N_18079);
or UO_1336 (O_1336,N_18318,N_18870);
nand UO_1337 (O_1337,N_18377,N_19805);
and UO_1338 (O_1338,N_18354,N_19427);
nor UO_1339 (O_1339,N_18430,N_18765);
nor UO_1340 (O_1340,N_18257,N_19644);
xnor UO_1341 (O_1341,N_18642,N_18449);
and UO_1342 (O_1342,N_19258,N_19900);
nor UO_1343 (O_1343,N_18244,N_18034);
or UO_1344 (O_1344,N_19769,N_18245);
and UO_1345 (O_1345,N_18644,N_18773);
nand UO_1346 (O_1346,N_19185,N_19069);
and UO_1347 (O_1347,N_18199,N_19101);
nor UO_1348 (O_1348,N_18019,N_18609);
and UO_1349 (O_1349,N_19470,N_19612);
nand UO_1350 (O_1350,N_19353,N_18910);
nand UO_1351 (O_1351,N_18729,N_19891);
and UO_1352 (O_1352,N_19395,N_19571);
and UO_1353 (O_1353,N_18786,N_19318);
and UO_1354 (O_1354,N_18880,N_18326);
nand UO_1355 (O_1355,N_18056,N_19395);
or UO_1356 (O_1356,N_19528,N_19979);
nor UO_1357 (O_1357,N_19751,N_19922);
nand UO_1358 (O_1358,N_19610,N_18087);
and UO_1359 (O_1359,N_18109,N_19863);
nor UO_1360 (O_1360,N_18129,N_19812);
nand UO_1361 (O_1361,N_18720,N_18568);
and UO_1362 (O_1362,N_18568,N_19942);
nor UO_1363 (O_1363,N_19320,N_19689);
nor UO_1364 (O_1364,N_19246,N_18018);
and UO_1365 (O_1365,N_19548,N_18690);
and UO_1366 (O_1366,N_19004,N_19827);
nor UO_1367 (O_1367,N_19939,N_19573);
or UO_1368 (O_1368,N_18900,N_19280);
or UO_1369 (O_1369,N_18971,N_19271);
nand UO_1370 (O_1370,N_19385,N_18275);
or UO_1371 (O_1371,N_18220,N_19737);
xnor UO_1372 (O_1372,N_18423,N_18179);
or UO_1373 (O_1373,N_18228,N_19299);
or UO_1374 (O_1374,N_18645,N_19152);
xor UO_1375 (O_1375,N_19014,N_18886);
nand UO_1376 (O_1376,N_19587,N_18294);
and UO_1377 (O_1377,N_19693,N_18465);
nor UO_1378 (O_1378,N_18013,N_18401);
or UO_1379 (O_1379,N_18785,N_18196);
or UO_1380 (O_1380,N_18002,N_19843);
nand UO_1381 (O_1381,N_19285,N_19279);
nand UO_1382 (O_1382,N_18107,N_19155);
or UO_1383 (O_1383,N_19787,N_18059);
nor UO_1384 (O_1384,N_19676,N_19441);
and UO_1385 (O_1385,N_19039,N_18053);
xor UO_1386 (O_1386,N_18333,N_19669);
or UO_1387 (O_1387,N_19266,N_19183);
nor UO_1388 (O_1388,N_19494,N_19416);
nor UO_1389 (O_1389,N_18735,N_18588);
and UO_1390 (O_1390,N_18889,N_19046);
and UO_1391 (O_1391,N_18091,N_18685);
and UO_1392 (O_1392,N_18681,N_18857);
and UO_1393 (O_1393,N_18226,N_19080);
and UO_1394 (O_1394,N_19411,N_18613);
nor UO_1395 (O_1395,N_19654,N_18699);
nor UO_1396 (O_1396,N_19708,N_18347);
xnor UO_1397 (O_1397,N_19274,N_19001);
nand UO_1398 (O_1398,N_19308,N_18605);
and UO_1399 (O_1399,N_19029,N_18506);
and UO_1400 (O_1400,N_19143,N_18897);
nand UO_1401 (O_1401,N_19139,N_18467);
nand UO_1402 (O_1402,N_18676,N_18953);
xor UO_1403 (O_1403,N_18348,N_19170);
nand UO_1404 (O_1404,N_19511,N_19279);
and UO_1405 (O_1405,N_19682,N_18411);
xnor UO_1406 (O_1406,N_18668,N_19410);
xor UO_1407 (O_1407,N_18797,N_19368);
nor UO_1408 (O_1408,N_18928,N_18448);
or UO_1409 (O_1409,N_18791,N_18189);
xor UO_1410 (O_1410,N_18319,N_19138);
xnor UO_1411 (O_1411,N_19734,N_18664);
and UO_1412 (O_1412,N_19739,N_19018);
xnor UO_1413 (O_1413,N_19134,N_18467);
and UO_1414 (O_1414,N_19052,N_19581);
xnor UO_1415 (O_1415,N_18398,N_18199);
xnor UO_1416 (O_1416,N_19274,N_19030);
or UO_1417 (O_1417,N_19822,N_18221);
nor UO_1418 (O_1418,N_18442,N_19186);
xor UO_1419 (O_1419,N_18351,N_18196);
nand UO_1420 (O_1420,N_18744,N_18682);
and UO_1421 (O_1421,N_19364,N_18349);
nor UO_1422 (O_1422,N_19036,N_18338);
nand UO_1423 (O_1423,N_18951,N_19259);
nand UO_1424 (O_1424,N_18285,N_19102);
nor UO_1425 (O_1425,N_19924,N_18999);
or UO_1426 (O_1426,N_18187,N_19113);
and UO_1427 (O_1427,N_18281,N_18564);
nand UO_1428 (O_1428,N_18949,N_18762);
and UO_1429 (O_1429,N_19536,N_19746);
nand UO_1430 (O_1430,N_18532,N_18989);
nor UO_1431 (O_1431,N_18330,N_18622);
nand UO_1432 (O_1432,N_19151,N_18174);
nor UO_1433 (O_1433,N_19475,N_18088);
xor UO_1434 (O_1434,N_18601,N_19990);
or UO_1435 (O_1435,N_19307,N_19923);
or UO_1436 (O_1436,N_19016,N_19416);
nor UO_1437 (O_1437,N_19282,N_18169);
nor UO_1438 (O_1438,N_18319,N_19894);
or UO_1439 (O_1439,N_19722,N_19680);
nand UO_1440 (O_1440,N_18901,N_19022);
or UO_1441 (O_1441,N_18906,N_18294);
or UO_1442 (O_1442,N_18906,N_19315);
and UO_1443 (O_1443,N_18933,N_18443);
xor UO_1444 (O_1444,N_18986,N_18384);
and UO_1445 (O_1445,N_18183,N_19751);
or UO_1446 (O_1446,N_19720,N_19290);
or UO_1447 (O_1447,N_19037,N_18764);
xnor UO_1448 (O_1448,N_18078,N_18981);
nor UO_1449 (O_1449,N_18518,N_19564);
and UO_1450 (O_1450,N_19960,N_19306);
and UO_1451 (O_1451,N_19222,N_18906);
nor UO_1452 (O_1452,N_18215,N_19903);
nand UO_1453 (O_1453,N_18026,N_18384);
nor UO_1454 (O_1454,N_19208,N_18980);
nor UO_1455 (O_1455,N_19000,N_18990);
nor UO_1456 (O_1456,N_18041,N_18840);
nor UO_1457 (O_1457,N_18805,N_19441);
xnor UO_1458 (O_1458,N_19122,N_18141);
or UO_1459 (O_1459,N_18610,N_18281);
xor UO_1460 (O_1460,N_18156,N_18701);
and UO_1461 (O_1461,N_19514,N_19176);
or UO_1462 (O_1462,N_19070,N_19001);
and UO_1463 (O_1463,N_18586,N_19386);
and UO_1464 (O_1464,N_18628,N_19703);
and UO_1465 (O_1465,N_18164,N_19677);
nand UO_1466 (O_1466,N_19847,N_19127);
or UO_1467 (O_1467,N_19106,N_19956);
and UO_1468 (O_1468,N_18958,N_18269);
or UO_1469 (O_1469,N_19303,N_19232);
and UO_1470 (O_1470,N_19243,N_19242);
nor UO_1471 (O_1471,N_18897,N_18344);
xnor UO_1472 (O_1472,N_18206,N_19425);
nor UO_1473 (O_1473,N_19725,N_18866);
nand UO_1474 (O_1474,N_18834,N_19355);
nor UO_1475 (O_1475,N_18716,N_19000);
nand UO_1476 (O_1476,N_18363,N_18116);
xnor UO_1477 (O_1477,N_19804,N_18867);
and UO_1478 (O_1478,N_18228,N_18660);
nand UO_1479 (O_1479,N_19483,N_18525);
nor UO_1480 (O_1480,N_18878,N_18464);
nand UO_1481 (O_1481,N_18979,N_18969);
and UO_1482 (O_1482,N_18926,N_19235);
nand UO_1483 (O_1483,N_18753,N_18810);
nor UO_1484 (O_1484,N_19906,N_18294);
xor UO_1485 (O_1485,N_18720,N_19199);
nor UO_1486 (O_1486,N_19408,N_19535);
or UO_1487 (O_1487,N_19321,N_19464);
xnor UO_1488 (O_1488,N_18599,N_18548);
and UO_1489 (O_1489,N_18434,N_18383);
and UO_1490 (O_1490,N_19285,N_19706);
xnor UO_1491 (O_1491,N_18272,N_19731);
or UO_1492 (O_1492,N_18709,N_19843);
and UO_1493 (O_1493,N_18956,N_18241);
xnor UO_1494 (O_1494,N_19905,N_18787);
and UO_1495 (O_1495,N_19947,N_18946);
nor UO_1496 (O_1496,N_19315,N_18347);
or UO_1497 (O_1497,N_19229,N_19604);
or UO_1498 (O_1498,N_19450,N_19190);
xnor UO_1499 (O_1499,N_18790,N_18402);
and UO_1500 (O_1500,N_18757,N_18746);
nand UO_1501 (O_1501,N_18392,N_18529);
xor UO_1502 (O_1502,N_18042,N_19198);
xnor UO_1503 (O_1503,N_19528,N_18936);
or UO_1504 (O_1504,N_18093,N_19733);
or UO_1505 (O_1505,N_19626,N_18277);
nand UO_1506 (O_1506,N_18614,N_19131);
nor UO_1507 (O_1507,N_19546,N_18876);
or UO_1508 (O_1508,N_19743,N_18772);
nor UO_1509 (O_1509,N_18952,N_18727);
xnor UO_1510 (O_1510,N_18519,N_18689);
nand UO_1511 (O_1511,N_19571,N_19653);
xnor UO_1512 (O_1512,N_19187,N_18918);
xnor UO_1513 (O_1513,N_18674,N_19090);
or UO_1514 (O_1514,N_19246,N_19429);
and UO_1515 (O_1515,N_18443,N_18584);
nor UO_1516 (O_1516,N_18002,N_19723);
xor UO_1517 (O_1517,N_18577,N_18159);
xor UO_1518 (O_1518,N_19312,N_19826);
or UO_1519 (O_1519,N_18383,N_18663);
xor UO_1520 (O_1520,N_19815,N_19465);
nor UO_1521 (O_1521,N_19071,N_18565);
nor UO_1522 (O_1522,N_19330,N_18159);
or UO_1523 (O_1523,N_18839,N_19068);
nand UO_1524 (O_1524,N_19557,N_19207);
xor UO_1525 (O_1525,N_19621,N_18260);
nand UO_1526 (O_1526,N_19714,N_19125);
xor UO_1527 (O_1527,N_19422,N_19683);
or UO_1528 (O_1528,N_18540,N_19373);
xnor UO_1529 (O_1529,N_18891,N_19844);
nand UO_1530 (O_1530,N_18489,N_18497);
or UO_1531 (O_1531,N_19019,N_18366);
or UO_1532 (O_1532,N_19253,N_19429);
and UO_1533 (O_1533,N_18692,N_19520);
nand UO_1534 (O_1534,N_19079,N_18239);
and UO_1535 (O_1535,N_19195,N_19148);
and UO_1536 (O_1536,N_19949,N_19830);
and UO_1537 (O_1537,N_19790,N_18993);
or UO_1538 (O_1538,N_19473,N_19780);
nand UO_1539 (O_1539,N_18186,N_19152);
nand UO_1540 (O_1540,N_18778,N_18176);
xor UO_1541 (O_1541,N_18233,N_18581);
and UO_1542 (O_1542,N_18231,N_19076);
nand UO_1543 (O_1543,N_18496,N_18861);
and UO_1544 (O_1544,N_18304,N_19495);
or UO_1545 (O_1545,N_19266,N_19332);
or UO_1546 (O_1546,N_18752,N_18677);
nand UO_1547 (O_1547,N_18217,N_18189);
or UO_1548 (O_1548,N_19579,N_18849);
nand UO_1549 (O_1549,N_19636,N_18251);
nor UO_1550 (O_1550,N_19576,N_19543);
xor UO_1551 (O_1551,N_19365,N_19003);
xor UO_1552 (O_1552,N_18082,N_18716);
nor UO_1553 (O_1553,N_19199,N_18833);
nand UO_1554 (O_1554,N_18139,N_19979);
and UO_1555 (O_1555,N_19019,N_19883);
and UO_1556 (O_1556,N_18819,N_19973);
xnor UO_1557 (O_1557,N_19988,N_19240);
or UO_1558 (O_1558,N_18939,N_19191);
nand UO_1559 (O_1559,N_18722,N_19843);
xnor UO_1560 (O_1560,N_19726,N_18658);
nor UO_1561 (O_1561,N_19989,N_19786);
nor UO_1562 (O_1562,N_19064,N_19182);
or UO_1563 (O_1563,N_19706,N_19057);
or UO_1564 (O_1564,N_18883,N_19976);
nor UO_1565 (O_1565,N_19621,N_18292);
nand UO_1566 (O_1566,N_18057,N_18485);
and UO_1567 (O_1567,N_19374,N_18704);
nor UO_1568 (O_1568,N_18555,N_18988);
nand UO_1569 (O_1569,N_19357,N_19263);
nand UO_1570 (O_1570,N_18393,N_18858);
nand UO_1571 (O_1571,N_19396,N_19224);
and UO_1572 (O_1572,N_18353,N_18186);
and UO_1573 (O_1573,N_18095,N_19967);
nor UO_1574 (O_1574,N_19608,N_18976);
nor UO_1575 (O_1575,N_19403,N_19433);
xor UO_1576 (O_1576,N_18674,N_18522);
xor UO_1577 (O_1577,N_19093,N_19640);
and UO_1578 (O_1578,N_19178,N_18982);
xnor UO_1579 (O_1579,N_19833,N_18873);
xor UO_1580 (O_1580,N_19033,N_18648);
and UO_1581 (O_1581,N_19805,N_18925);
nor UO_1582 (O_1582,N_18151,N_18830);
or UO_1583 (O_1583,N_19667,N_19628);
or UO_1584 (O_1584,N_18594,N_18363);
and UO_1585 (O_1585,N_18550,N_18025);
nand UO_1586 (O_1586,N_18611,N_18077);
nand UO_1587 (O_1587,N_18869,N_19044);
nor UO_1588 (O_1588,N_19000,N_18761);
nand UO_1589 (O_1589,N_19624,N_19577);
xnor UO_1590 (O_1590,N_18039,N_19662);
nor UO_1591 (O_1591,N_18564,N_18210);
and UO_1592 (O_1592,N_18294,N_18502);
or UO_1593 (O_1593,N_18907,N_19588);
nand UO_1594 (O_1594,N_19778,N_19958);
nor UO_1595 (O_1595,N_18680,N_18863);
nor UO_1596 (O_1596,N_18974,N_18137);
nor UO_1597 (O_1597,N_18322,N_18207);
nand UO_1598 (O_1598,N_19618,N_18756);
xor UO_1599 (O_1599,N_19000,N_18911);
nand UO_1600 (O_1600,N_18704,N_19754);
nor UO_1601 (O_1601,N_18852,N_19007);
or UO_1602 (O_1602,N_18534,N_18445);
and UO_1603 (O_1603,N_18452,N_18371);
and UO_1604 (O_1604,N_18429,N_18506);
or UO_1605 (O_1605,N_19958,N_18622);
and UO_1606 (O_1606,N_18476,N_19185);
nand UO_1607 (O_1607,N_18099,N_19135);
nor UO_1608 (O_1608,N_18243,N_19391);
or UO_1609 (O_1609,N_18749,N_18566);
xnor UO_1610 (O_1610,N_18340,N_19128);
or UO_1611 (O_1611,N_19705,N_18585);
and UO_1612 (O_1612,N_18298,N_18964);
and UO_1613 (O_1613,N_19630,N_19403);
or UO_1614 (O_1614,N_19741,N_19714);
and UO_1615 (O_1615,N_18951,N_19085);
nor UO_1616 (O_1616,N_19340,N_18205);
or UO_1617 (O_1617,N_19040,N_18362);
xnor UO_1618 (O_1618,N_19812,N_18830);
and UO_1619 (O_1619,N_18881,N_19803);
nor UO_1620 (O_1620,N_18094,N_19770);
nand UO_1621 (O_1621,N_19964,N_19090);
xor UO_1622 (O_1622,N_18156,N_18890);
nor UO_1623 (O_1623,N_19454,N_18613);
nand UO_1624 (O_1624,N_18675,N_19593);
nand UO_1625 (O_1625,N_19864,N_19752);
or UO_1626 (O_1626,N_18451,N_19343);
nor UO_1627 (O_1627,N_19856,N_18800);
nand UO_1628 (O_1628,N_18758,N_19050);
or UO_1629 (O_1629,N_18346,N_19870);
and UO_1630 (O_1630,N_18894,N_19182);
or UO_1631 (O_1631,N_19109,N_19347);
and UO_1632 (O_1632,N_19883,N_19055);
and UO_1633 (O_1633,N_19801,N_19721);
xnor UO_1634 (O_1634,N_18762,N_19313);
nor UO_1635 (O_1635,N_19331,N_18525);
and UO_1636 (O_1636,N_19205,N_18655);
or UO_1637 (O_1637,N_18304,N_18254);
nor UO_1638 (O_1638,N_18802,N_19506);
nor UO_1639 (O_1639,N_19635,N_19643);
or UO_1640 (O_1640,N_18612,N_18434);
nor UO_1641 (O_1641,N_18213,N_18974);
and UO_1642 (O_1642,N_19463,N_18917);
or UO_1643 (O_1643,N_18884,N_18595);
and UO_1644 (O_1644,N_18735,N_19174);
xor UO_1645 (O_1645,N_18641,N_19528);
and UO_1646 (O_1646,N_19487,N_18592);
nor UO_1647 (O_1647,N_18069,N_18502);
nor UO_1648 (O_1648,N_18998,N_19234);
or UO_1649 (O_1649,N_18179,N_18519);
nor UO_1650 (O_1650,N_19544,N_19122);
and UO_1651 (O_1651,N_18935,N_18619);
xnor UO_1652 (O_1652,N_19209,N_19625);
or UO_1653 (O_1653,N_18044,N_18321);
and UO_1654 (O_1654,N_18624,N_18979);
xnor UO_1655 (O_1655,N_19233,N_19654);
and UO_1656 (O_1656,N_18140,N_18717);
or UO_1657 (O_1657,N_19349,N_18759);
xnor UO_1658 (O_1658,N_18270,N_18938);
nand UO_1659 (O_1659,N_18186,N_18022);
or UO_1660 (O_1660,N_19419,N_19415);
nor UO_1661 (O_1661,N_18390,N_19178);
or UO_1662 (O_1662,N_18769,N_19566);
and UO_1663 (O_1663,N_18688,N_19334);
nand UO_1664 (O_1664,N_18334,N_19677);
xnor UO_1665 (O_1665,N_19018,N_18211);
and UO_1666 (O_1666,N_19909,N_18552);
or UO_1667 (O_1667,N_19915,N_19789);
nand UO_1668 (O_1668,N_18114,N_18892);
nand UO_1669 (O_1669,N_19503,N_18587);
nor UO_1670 (O_1670,N_18794,N_19022);
or UO_1671 (O_1671,N_18345,N_19637);
or UO_1672 (O_1672,N_18793,N_19213);
xor UO_1673 (O_1673,N_19056,N_19286);
or UO_1674 (O_1674,N_19003,N_19251);
nand UO_1675 (O_1675,N_19392,N_19082);
and UO_1676 (O_1676,N_19152,N_18595);
xor UO_1677 (O_1677,N_18455,N_18512);
xnor UO_1678 (O_1678,N_18997,N_18897);
xor UO_1679 (O_1679,N_18650,N_19787);
xnor UO_1680 (O_1680,N_18024,N_19524);
xnor UO_1681 (O_1681,N_19869,N_19822);
and UO_1682 (O_1682,N_18865,N_18647);
nand UO_1683 (O_1683,N_18165,N_18150);
xnor UO_1684 (O_1684,N_19663,N_18946);
xor UO_1685 (O_1685,N_19661,N_19250);
and UO_1686 (O_1686,N_18978,N_18138);
nand UO_1687 (O_1687,N_19002,N_18304);
xnor UO_1688 (O_1688,N_18129,N_18100);
or UO_1689 (O_1689,N_18020,N_19737);
nor UO_1690 (O_1690,N_18640,N_19118);
nor UO_1691 (O_1691,N_18680,N_18996);
or UO_1692 (O_1692,N_18918,N_18259);
and UO_1693 (O_1693,N_18099,N_19211);
nor UO_1694 (O_1694,N_19064,N_18882);
nand UO_1695 (O_1695,N_19906,N_18084);
nor UO_1696 (O_1696,N_18191,N_19588);
and UO_1697 (O_1697,N_19732,N_19734);
or UO_1698 (O_1698,N_18404,N_19541);
nor UO_1699 (O_1699,N_18636,N_18067);
nand UO_1700 (O_1700,N_19273,N_18207);
and UO_1701 (O_1701,N_19139,N_19839);
nor UO_1702 (O_1702,N_18907,N_19830);
nor UO_1703 (O_1703,N_19124,N_18123);
nand UO_1704 (O_1704,N_18549,N_18415);
nand UO_1705 (O_1705,N_19531,N_19617);
and UO_1706 (O_1706,N_19729,N_18655);
xor UO_1707 (O_1707,N_18655,N_18384);
nand UO_1708 (O_1708,N_19987,N_18416);
xor UO_1709 (O_1709,N_18820,N_19158);
xor UO_1710 (O_1710,N_19631,N_19183);
nor UO_1711 (O_1711,N_18590,N_19298);
or UO_1712 (O_1712,N_19019,N_18955);
or UO_1713 (O_1713,N_19897,N_18638);
and UO_1714 (O_1714,N_19751,N_19841);
xor UO_1715 (O_1715,N_19111,N_18707);
or UO_1716 (O_1716,N_19582,N_18435);
xor UO_1717 (O_1717,N_18050,N_18785);
or UO_1718 (O_1718,N_19813,N_19742);
nand UO_1719 (O_1719,N_19912,N_18863);
nand UO_1720 (O_1720,N_18192,N_18104);
and UO_1721 (O_1721,N_18141,N_18679);
nor UO_1722 (O_1722,N_19919,N_18903);
nor UO_1723 (O_1723,N_19384,N_18421);
and UO_1724 (O_1724,N_18763,N_18644);
nand UO_1725 (O_1725,N_19226,N_18550);
xnor UO_1726 (O_1726,N_18596,N_18797);
nor UO_1727 (O_1727,N_18712,N_19908);
nand UO_1728 (O_1728,N_18258,N_18695);
nor UO_1729 (O_1729,N_18977,N_18432);
nand UO_1730 (O_1730,N_18775,N_18505);
or UO_1731 (O_1731,N_19373,N_18658);
xnor UO_1732 (O_1732,N_18841,N_18692);
xnor UO_1733 (O_1733,N_18291,N_18551);
xnor UO_1734 (O_1734,N_18803,N_18722);
nor UO_1735 (O_1735,N_18299,N_19322);
or UO_1736 (O_1736,N_18156,N_18292);
and UO_1737 (O_1737,N_19250,N_19275);
xnor UO_1738 (O_1738,N_18103,N_18108);
or UO_1739 (O_1739,N_18654,N_19514);
nand UO_1740 (O_1740,N_19950,N_18224);
or UO_1741 (O_1741,N_19874,N_19780);
xnor UO_1742 (O_1742,N_18433,N_19799);
nand UO_1743 (O_1743,N_19746,N_19322);
and UO_1744 (O_1744,N_19545,N_18819);
nor UO_1745 (O_1745,N_19276,N_18756);
xnor UO_1746 (O_1746,N_18937,N_19078);
xor UO_1747 (O_1747,N_18581,N_18609);
or UO_1748 (O_1748,N_18815,N_18049);
nand UO_1749 (O_1749,N_19449,N_19697);
xor UO_1750 (O_1750,N_19626,N_19147);
nand UO_1751 (O_1751,N_18311,N_18557);
or UO_1752 (O_1752,N_19708,N_18528);
xnor UO_1753 (O_1753,N_19582,N_19667);
xnor UO_1754 (O_1754,N_19214,N_19443);
xor UO_1755 (O_1755,N_18502,N_18147);
and UO_1756 (O_1756,N_19241,N_19091);
xnor UO_1757 (O_1757,N_18398,N_18555);
nor UO_1758 (O_1758,N_18129,N_18127);
or UO_1759 (O_1759,N_19686,N_19788);
and UO_1760 (O_1760,N_19778,N_18743);
nor UO_1761 (O_1761,N_18466,N_19351);
xnor UO_1762 (O_1762,N_18545,N_19082);
nor UO_1763 (O_1763,N_18646,N_18979);
nor UO_1764 (O_1764,N_19932,N_19105);
or UO_1765 (O_1765,N_19171,N_19239);
and UO_1766 (O_1766,N_19516,N_18923);
and UO_1767 (O_1767,N_18192,N_18027);
nand UO_1768 (O_1768,N_18683,N_18190);
nand UO_1769 (O_1769,N_18383,N_18547);
nor UO_1770 (O_1770,N_19886,N_19252);
nand UO_1771 (O_1771,N_18158,N_19142);
xor UO_1772 (O_1772,N_19529,N_19331);
nand UO_1773 (O_1773,N_19019,N_19232);
nand UO_1774 (O_1774,N_18299,N_19769);
xor UO_1775 (O_1775,N_19082,N_19458);
nor UO_1776 (O_1776,N_18128,N_19607);
nor UO_1777 (O_1777,N_18120,N_18689);
and UO_1778 (O_1778,N_19417,N_18115);
xor UO_1779 (O_1779,N_18667,N_18775);
nor UO_1780 (O_1780,N_19434,N_18585);
xnor UO_1781 (O_1781,N_19390,N_18028);
and UO_1782 (O_1782,N_19192,N_19904);
or UO_1783 (O_1783,N_19244,N_19076);
nor UO_1784 (O_1784,N_18397,N_18768);
nand UO_1785 (O_1785,N_18511,N_18972);
and UO_1786 (O_1786,N_19286,N_18159);
xnor UO_1787 (O_1787,N_18357,N_19428);
nand UO_1788 (O_1788,N_18929,N_19984);
and UO_1789 (O_1789,N_18382,N_19517);
nor UO_1790 (O_1790,N_18560,N_18042);
nor UO_1791 (O_1791,N_19268,N_19247);
xor UO_1792 (O_1792,N_19053,N_19043);
nor UO_1793 (O_1793,N_18879,N_19860);
nor UO_1794 (O_1794,N_18079,N_19123);
nand UO_1795 (O_1795,N_19165,N_18311);
nor UO_1796 (O_1796,N_18740,N_19047);
xnor UO_1797 (O_1797,N_18816,N_18969);
nor UO_1798 (O_1798,N_18862,N_19177);
and UO_1799 (O_1799,N_19513,N_18173);
nand UO_1800 (O_1800,N_19395,N_19832);
and UO_1801 (O_1801,N_18463,N_19667);
nand UO_1802 (O_1802,N_19754,N_19592);
xnor UO_1803 (O_1803,N_18009,N_19348);
and UO_1804 (O_1804,N_18824,N_19937);
or UO_1805 (O_1805,N_18807,N_19521);
nor UO_1806 (O_1806,N_19059,N_19637);
xor UO_1807 (O_1807,N_19766,N_19156);
and UO_1808 (O_1808,N_18732,N_19435);
or UO_1809 (O_1809,N_19423,N_18995);
or UO_1810 (O_1810,N_19086,N_19182);
xor UO_1811 (O_1811,N_18337,N_18531);
or UO_1812 (O_1812,N_19896,N_18867);
and UO_1813 (O_1813,N_19339,N_19133);
or UO_1814 (O_1814,N_19717,N_19372);
nor UO_1815 (O_1815,N_18067,N_18120);
xnor UO_1816 (O_1816,N_18030,N_19687);
or UO_1817 (O_1817,N_19393,N_18750);
nand UO_1818 (O_1818,N_19476,N_19091);
xor UO_1819 (O_1819,N_18097,N_18877);
and UO_1820 (O_1820,N_18086,N_19278);
or UO_1821 (O_1821,N_18971,N_18381);
xor UO_1822 (O_1822,N_18471,N_18969);
nand UO_1823 (O_1823,N_18933,N_18326);
nor UO_1824 (O_1824,N_18581,N_19688);
and UO_1825 (O_1825,N_19798,N_18833);
xnor UO_1826 (O_1826,N_18237,N_19336);
or UO_1827 (O_1827,N_18869,N_19098);
nand UO_1828 (O_1828,N_19453,N_19886);
and UO_1829 (O_1829,N_19142,N_18314);
or UO_1830 (O_1830,N_19020,N_18691);
or UO_1831 (O_1831,N_18311,N_19034);
nor UO_1832 (O_1832,N_19216,N_18818);
nand UO_1833 (O_1833,N_18573,N_18545);
or UO_1834 (O_1834,N_18955,N_19490);
and UO_1835 (O_1835,N_18837,N_19764);
or UO_1836 (O_1836,N_19131,N_18159);
nand UO_1837 (O_1837,N_19325,N_18669);
xor UO_1838 (O_1838,N_18923,N_18296);
nand UO_1839 (O_1839,N_18551,N_18941);
and UO_1840 (O_1840,N_19420,N_18131);
nand UO_1841 (O_1841,N_18413,N_18282);
and UO_1842 (O_1842,N_18044,N_18744);
nor UO_1843 (O_1843,N_19573,N_18688);
nor UO_1844 (O_1844,N_19202,N_19941);
xnor UO_1845 (O_1845,N_19341,N_19704);
and UO_1846 (O_1846,N_18635,N_19746);
or UO_1847 (O_1847,N_18140,N_18247);
and UO_1848 (O_1848,N_18516,N_19188);
and UO_1849 (O_1849,N_18659,N_19487);
xnor UO_1850 (O_1850,N_19076,N_18665);
xor UO_1851 (O_1851,N_19456,N_18425);
or UO_1852 (O_1852,N_18692,N_18206);
nand UO_1853 (O_1853,N_18760,N_19032);
or UO_1854 (O_1854,N_18850,N_19863);
nor UO_1855 (O_1855,N_19497,N_19913);
nor UO_1856 (O_1856,N_19911,N_18834);
or UO_1857 (O_1857,N_19107,N_18944);
nor UO_1858 (O_1858,N_19326,N_18484);
nand UO_1859 (O_1859,N_18777,N_18744);
xor UO_1860 (O_1860,N_18238,N_19792);
and UO_1861 (O_1861,N_18219,N_18032);
xor UO_1862 (O_1862,N_18853,N_18931);
or UO_1863 (O_1863,N_18719,N_19336);
or UO_1864 (O_1864,N_19069,N_19034);
nand UO_1865 (O_1865,N_19971,N_18754);
nand UO_1866 (O_1866,N_19877,N_18555);
or UO_1867 (O_1867,N_18361,N_19076);
or UO_1868 (O_1868,N_19755,N_19370);
nor UO_1869 (O_1869,N_19660,N_18524);
or UO_1870 (O_1870,N_18725,N_19579);
xor UO_1871 (O_1871,N_18590,N_18760);
nor UO_1872 (O_1872,N_18850,N_19392);
nor UO_1873 (O_1873,N_18116,N_18544);
nand UO_1874 (O_1874,N_18802,N_18183);
nor UO_1875 (O_1875,N_18638,N_18950);
or UO_1876 (O_1876,N_19187,N_18000);
or UO_1877 (O_1877,N_18941,N_18262);
or UO_1878 (O_1878,N_19592,N_19574);
nor UO_1879 (O_1879,N_18401,N_18428);
xnor UO_1880 (O_1880,N_18414,N_19770);
nand UO_1881 (O_1881,N_19633,N_19500);
nand UO_1882 (O_1882,N_19810,N_18466);
or UO_1883 (O_1883,N_19205,N_18734);
or UO_1884 (O_1884,N_18107,N_18984);
nand UO_1885 (O_1885,N_19692,N_18640);
and UO_1886 (O_1886,N_19707,N_19244);
xor UO_1887 (O_1887,N_19123,N_19624);
nand UO_1888 (O_1888,N_18870,N_18729);
or UO_1889 (O_1889,N_19763,N_18132);
xor UO_1890 (O_1890,N_18869,N_18914);
xor UO_1891 (O_1891,N_18303,N_18008);
nand UO_1892 (O_1892,N_18779,N_18510);
or UO_1893 (O_1893,N_18981,N_19730);
or UO_1894 (O_1894,N_18661,N_19152);
nand UO_1895 (O_1895,N_19993,N_18963);
nor UO_1896 (O_1896,N_19262,N_19259);
or UO_1897 (O_1897,N_19287,N_18919);
xor UO_1898 (O_1898,N_19378,N_18951);
and UO_1899 (O_1899,N_19297,N_19661);
xor UO_1900 (O_1900,N_18595,N_19490);
and UO_1901 (O_1901,N_18556,N_19320);
nand UO_1902 (O_1902,N_19933,N_18233);
nor UO_1903 (O_1903,N_19655,N_18780);
and UO_1904 (O_1904,N_19283,N_18803);
nand UO_1905 (O_1905,N_18352,N_18229);
xor UO_1906 (O_1906,N_19252,N_18258);
and UO_1907 (O_1907,N_19999,N_18428);
nand UO_1908 (O_1908,N_18649,N_18906);
xnor UO_1909 (O_1909,N_18604,N_18595);
xor UO_1910 (O_1910,N_18805,N_19216);
xor UO_1911 (O_1911,N_19442,N_18315);
or UO_1912 (O_1912,N_19029,N_18716);
nand UO_1913 (O_1913,N_19341,N_18270);
xnor UO_1914 (O_1914,N_18325,N_19591);
nor UO_1915 (O_1915,N_18216,N_18736);
or UO_1916 (O_1916,N_19566,N_19726);
or UO_1917 (O_1917,N_19845,N_19516);
and UO_1918 (O_1918,N_18724,N_18569);
xnor UO_1919 (O_1919,N_18408,N_19307);
nor UO_1920 (O_1920,N_19791,N_18393);
and UO_1921 (O_1921,N_19668,N_19339);
and UO_1922 (O_1922,N_19594,N_18426);
and UO_1923 (O_1923,N_19375,N_19413);
nand UO_1924 (O_1924,N_19606,N_18413);
and UO_1925 (O_1925,N_19191,N_18097);
nor UO_1926 (O_1926,N_19010,N_18148);
and UO_1927 (O_1927,N_19708,N_19746);
and UO_1928 (O_1928,N_19867,N_18565);
nor UO_1929 (O_1929,N_18912,N_18188);
or UO_1930 (O_1930,N_19554,N_19769);
xnor UO_1931 (O_1931,N_19345,N_18478);
and UO_1932 (O_1932,N_19622,N_18258);
nand UO_1933 (O_1933,N_18491,N_18891);
or UO_1934 (O_1934,N_18196,N_19382);
nor UO_1935 (O_1935,N_18844,N_19004);
or UO_1936 (O_1936,N_18088,N_18245);
nand UO_1937 (O_1937,N_18276,N_18137);
and UO_1938 (O_1938,N_19231,N_18992);
nor UO_1939 (O_1939,N_19522,N_18890);
nand UO_1940 (O_1940,N_18317,N_19690);
or UO_1941 (O_1941,N_18297,N_18416);
xor UO_1942 (O_1942,N_19867,N_19047);
xor UO_1943 (O_1943,N_19292,N_18488);
nor UO_1944 (O_1944,N_18904,N_19639);
nand UO_1945 (O_1945,N_18021,N_19358);
xor UO_1946 (O_1946,N_19934,N_18372);
nor UO_1947 (O_1947,N_19230,N_19227);
and UO_1948 (O_1948,N_18069,N_18361);
xor UO_1949 (O_1949,N_18470,N_19748);
and UO_1950 (O_1950,N_19944,N_18963);
or UO_1951 (O_1951,N_19642,N_18152);
or UO_1952 (O_1952,N_18514,N_19011);
nand UO_1953 (O_1953,N_19408,N_19155);
xnor UO_1954 (O_1954,N_18661,N_19931);
xnor UO_1955 (O_1955,N_18907,N_18132);
nand UO_1956 (O_1956,N_19959,N_18426);
xor UO_1957 (O_1957,N_18360,N_18970);
nand UO_1958 (O_1958,N_19700,N_19367);
and UO_1959 (O_1959,N_18726,N_19431);
nand UO_1960 (O_1960,N_19405,N_18095);
and UO_1961 (O_1961,N_19054,N_18579);
nand UO_1962 (O_1962,N_19980,N_19324);
and UO_1963 (O_1963,N_19701,N_19607);
xnor UO_1964 (O_1964,N_18940,N_18734);
nand UO_1965 (O_1965,N_18122,N_19463);
and UO_1966 (O_1966,N_18806,N_19700);
nor UO_1967 (O_1967,N_18368,N_19306);
nand UO_1968 (O_1968,N_18781,N_19958);
xor UO_1969 (O_1969,N_19072,N_19567);
xor UO_1970 (O_1970,N_18904,N_19905);
and UO_1971 (O_1971,N_18100,N_18298);
and UO_1972 (O_1972,N_18984,N_19994);
xor UO_1973 (O_1973,N_19012,N_18591);
nor UO_1974 (O_1974,N_18069,N_19762);
nand UO_1975 (O_1975,N_19802,N_19004);
and UO_1976 (O_1976,N_19887,N_19577);
or UO_1977 (O_1977,N_19322,N_18515);
and UO_1978 (O_1978,N_19804,N_18309);
or UO_1979 (O_1979,N_19169,N_18252);
and UO_1980 (O_1980,N_18674,N_19672);
nor UO_1981 (O_1981,N_18934,N_18406);
or UO_1982 (O_1982,N_18082,N_19334);
xor UO_1983 (O_1983,N_19542,N_18307);
nor UO_1984 (O_1984,N_18715,N_18933);
nor UO_1985 (O_1985,N_18433,N_19793);
or UO_1986 (O_1986,N_18700,N_19452);
xnor UO_1987 (O_1987,N_18194,N_19224);
nor UO_1988 (O_1988,N_19870,N_18045);
nand UO_1989 (O_1989,N_19660,N_19028);
nor UO_1990 (O_1990,N_19936,N_19198);
xnor UO_1991 (O_1991,N_19223,N_18304);
or UO_1992 (O_1992,N_18393,N_18873);
xnor UO_1993 (O_1993,N_19639,N_18763);
nor UO_1994 (O_1994,N_19979,N_19292);
xnor UO_1995 (O_1995,N_19442,N_18762);
and UO_1996 (O_1996,N_19981,N_19798);
and UO_1997 (O_1997,N_19888,N_19913);
nor UO_1998 (O_1998,N_19413,N_19806);
or UO_1999 (O_1999,N_18627,N_19066);
nand UO_2000 (O_2000,N_18176,N_19182);
nor UO_2001 (O_2001,N_19379,N_19907);
xnor UO_2002 (O_2002,N_19104,N_19362);
nand UO_2003 (O_2003,N_18034,N_19975);
xor UO_2004 (O_2004,N_19417,N_19536);
and UO_2005 (O_2005,N_18080,N_19277);
xor UO_2006 (O_2006,N_19129,N_18115);
nand UO_2007 (O_2007,N_19263,N_18160);
and UO_2008 (O_2008,N_19444,N_18556);
xor UO_2009 (O_2009,N_18487,N_18131);
nand UO_2010 (O_2010,N_18960,N_19275);
nand UO_2011 (O_2011,N_19848,N_19219);
nor UO_2012 (O_2012,N_18485,N_18273);
xnor UO_2013 (O_2013,N_19192,N_19996);
nand UO_2014 (O_2014,N_18181,N_19897);
nand UO_2015 (O_2015,N_18954,N_19507);
nand UO_2016 (O_2016,N_19853,N_18572);
nor UO_2017 (O_2017,N_19669,N_18360);
xor UO_2018 (O_2018,N_19403,N_19907);
nor UO_2019 (O_2019,N_19750,N_18148);
nand UO_2020 (O_2020,N_19747,N_18606);
nand UO_2021 (O_2021,N_18981,N_19668);
nand UO_2022 (O_2022,N_18610,N_18249);
xnor UO_2023 (O_2023,N_18075,N_19466);
xor UO_2024 (O_2024,N_19195,N_18424);
and UO_2025 (O_2025,N_18113,N_18675);
xor UO_2026 (O_2026,N_19320,N_19050);
and UO_2027 (O_2027,N_19157,N_19489);
or UO_2028 (O_2028,N_19526,N_18917);
xor UO_2029 (O_2029,N_18694,N_19254);
nand UO_2030 (O_2030,N_19517,N_19797);
xnor UO_2031 (O_2031,N_19516,N_19452);
or UO_2032 (O_2032,N_18916,N_19977);
xor UO_2033 (O_2033,N_19307,N_18787);
xnor UO_2034 (O_2034,N_19165,N_19294);
or UO_2035 (O_2035,N_19163,N_19793);
and UO_2036 (O_2036,N_18799,N_19058);
or UO_2037 (O_2037,N_19148,N_18087);
or UO_2038 (O_2038,N_19904,N_19457);
xor UO_2039 (O_2039,N_19787,N_18060);
nor UO_2040 (O_2040,N_19640,N_18148);
and UO_2041 (O_2041,N_19993,N_18669);
nor UO_2042 (O_2042,N_18908,N_19069);
and UO_2043 (O_2043,N_19214,N_18831);
and UO_2044 (O_2044,N_19322,N_19752);
nand UO_2045 (O_2045,N_19552,N_18435);
or UO_2046 (O_2046,N_18377,N_19595);
nand UO_2047 (O_2047,N_18112,N_18700);
nand UO_2048 (O_2048,N_19076,N_18120);
or UO_2049 (O_2049,N_19955,N_19991);
or UO_2050 (O_2050,N_19984,N_18869);
xor UO_2051 (O_2051,N_19196,N_19573);
nor UO_2052 (O_2052,N_19395,N_18161);
nand UO_2053 (O_2053,N_18150,N_18292);
and UO_2054 (O_2054,N_18332,N_19939);
or UO_2055 (O_2055,N_19665,N_18901);
nand UO_2056 (O_2056,N_19447,N_19144);
nand UO_2057 (O_2057,N_19032,N_18912);
nand UO_2058 (O_2058,N_19357,N_18292);
or UO_2059 (O_2059,N_19742,N_19475);
xnor UO_2060 (O_2060,N_18286,N_18230);
xnor UO_2061 (O_2061,N_19911,N_18647);
or UO_2062 (O_2062,N_18785,N_19142);
or UO_2063 (O_2063,N_19998,N_18101);
xor UO_2064 (O_2064,N_19645,N_18240);
and UO_2065 (O_2065,N_19700,N_18878);
nor UO_2066 (O_2066,N_18807,N_18100);
nand UO_2067 (O_2067,N_19695,N_19939);
nor UO_2068 (O_2068,N_19274,N_18885);
nand UO_2069 (O_2069,N_19490,N_19603);
nor UO_2070 (O_2070,N_19028,N_19609);
or UO_2071 (O_2071,N_18331,N_19864);
xnor UO_2072 (O_2072,N_18501,N_19012);
or UO_2073 (O_2073,N_18586,N_19622);
or UO_2074 (O_2074,N_18857,N_18566);
nand UO_2075 (O_2075,N_19493,N_19069);
or UO_2076 (O_2076,N_19144,N_18216);
xor UO_2077 (O_2077,N_18505,N_18636);
xor UO_2078 (O_2078,N_19414,N_18713);
nor UO_2079 (O_2079,N_18496,N_18950);
or UO_2080 (O_2080,N_18767,N_18452);
or UO_2081 (O_2081,N_18692,N_19705);
nor UO_2082 (O_2082,N_18433,N_18762);
and UO_2083 (O_2083,N_18972,N_18575);
nor UO_2084 (O_2084,N_19603,N_19664);
and UO_2085 (O_2085,N_19818,N_18315);
xnor UO_2086 (O_2086,N_18485,N_18698);
nor UO_2087 (O_2087,N_19476,N_18448);
and UO_2088 (O_2088,N_19359,N_19560);
xor UO_2089 (O_2089,N_18501,N_18112);
and UO_2090 (O_2090,N_19647,N_18078);
nand UO_2091 (O_2091,N_19501,N_19603);
nor UO_2092 (O_2092,N_18936,N_18704);
xor UO_2093 (O_2093,N_18715,N_19980);
nand UO_2094 (O_2094,N_19011,N_18808);
or UO_2095 (O_2095,N_18799,N_19702);
nand UO_2096 (O_2096,N_18914,N_19180);
nor UO_2097 (O_2097,N_19685,N_19542);
or UO_2098 (O_2098,N_18050,N_18391);
nor UO_2099 (O_2099,N_18996,N_19956);
nor UO_2100 (O_2100,N_19163,N_19671);
and UO_2101 (O_2101,N_18281,N_18306);
nor UO_2102 (O_2102,N_18770,N_18265);
xor UO_2103 (O_2103,N_19768,N_19879);
or UO_2104 (O_2104,N_18445,N_19863);
nor UO_2105 (O_2105,N_18056,N_19277);
xor UO_2106 (O_2106,N_19037,N_19170);
nor UO_2107 (O_2107,N_19429,N_19009);
and UO_2108 (O_2108,N_19718,N_18280);
nor UO_2109 (O_2109,N_19825,N_18617);
and UO_2110 (O_2110,N_19503,N_18655);
nor UO_2111 (O_2111,N_19013,N_18789);
nand UO_2112 (O_2112,N_19361,N_18020);
xnor UO_2113 (O_2113,N_18492,N_18883);
nand UO_2114 (O_2114,N_19946,N_19536);
nor UO_2115 (O_2115,N_19419,N_19251);
xor UO_2116 (O_2116,N_19421,N_19365);
or UO_2117 (O_2117,N_19571,N_19420);
or UO_2118 (O_2118,N_18908,N_19431);
and UO_2119 (O_2119,N_19783,N_18792);
nand UO_2120 (O_2120,N_18574,N_18862);
nor UO_2121 (O_2121,N_18619,N_19267);
and UO_2122 (O_2122,N_19969,N_18971);
and UO_2123 (O_2123,N_19513,N_19870);
or UO_2124 (O_2124,N_19934,N_18724);
or UO_2125 (O_2125,N_19665,N_18482);
or UO_2126 (O_2126,N_19787,N_19183);
xnor UO_2127 (O_2127,N_18304,N_19342);
or UO_2128 (O_2128,N_18577,N_19656);
xnor UO_2129 (O_2129,N_19020,N_19812);
and UO_2130 (O_2130,N_18393,N_18635);
xnor UO_2131 (O_2131,N_18647,N_18923);
and UO_2132 (O_2132,N_19197,N_19100);
and UO_2133 (O_2133,N_19480,N_18379);
nor UO_2134 (O_2134,N_18486,N_18679);
xnor UO_2135 (O_2135,N_18846,N_19499);
nor UO_2136 (O_2136,N_18351,N_18418);
xnor UO_2137 (O_2137,N_18299,N_19588);
xnor UO_2138 (O_2138,N_18244,N_18186);
or UO_2139 (O_2139,N_19108,N_19475);
nand UO_2140 (O_2140,N_18667,N_18056);
or UO_2141 (O_2141,N_18880,N_18662);
and UO_2142 (O_2142,N_19124,N_19557);
or UO_2143 (O_2143,N_19787,N_19132);
xor UO_2144 (O_2144,N_18907,N_19364);
and UO_2145 (O_2145,N_18678,N_18546);
xnor UO_2146 (O_2146,N_18239,N_19591);
or UO_2147 (O_2147,N_18515,N_18725);
xnor UO_2148 (O_2148,N_19726,N_18097);
or UO_2149 (O_2149,N_18811,N_18426);
nand UO_2150 (O_2150,N_18646,N_19045);
nor UO_2151 (O_2151,N_19925,N_19844);
xnor UO_2152 (O_2152,N_19511,N_18080);
nor UO_2153 (O_2153,N_18076,N_18578);
or UO_2154 (O_2154,N_19228,N_19250);
or UO_2155 (O_2155,N_18893,N_18596);
nand UO_2156 (O_2156,N_19429,N_19235);
xor UO_2157 (O_2157,N_19070,N_18472);
nor UO_2158 (O_2158,N_18387,N_19906);
xnor UO_2159 (O_2159,N_18633,N_19264);
nand UO_2160 (O_2160,N_18406,N_18624);
xor UO_2161 (O_2161,N_19993,N_19056);
nand UO_2162 (O_2162,N_18518,N_18010);
or UO_2163 (O_2163,N_19613,N_19062);
xnor UO_2164 (O_2164,N_19703,N_18782);
or UO_2165 (O_2165,N_18254,N_19005);
and UO_2166 (O_2166,N_18533,N_19122);
or UO_2167 (O_2167,N_18503,N_18867);
nand UO_2168 (O_2168,N_18333,N_19111);
nor UO_2169 (O_2169,N_19629,N_18385);
nand UO_2170 (O_2170,N_18223,N_19535);
xor UO_2171 (O_2171,N_19536,N_19124);
xor UO_2172 (O_2172,N_19400,N_18788);
and UO_2173 (O_2173,N_18101,N_19433);
and UO_2174 (O_2174,N_18193,N_18083);
or UO_2175 (O_2175,N_19050,N_18913);
nor UO_2176 (O_2176,N_19941,N_18851);
nand UO_2177 (O_2177,N_19184,N_19177);
nand UO_2178 (O_2178,N_18667,N_18305);
and UO_2179 (O_2179,N_18625,N_18975);
nor UO_2180 (O_2180,N_19206,N_19284);
xnor UO_2181 (O_2181,N_18838,N_19786);
nand UO_2182 (O_2182,N_18291,N_18220);
or UO_2183 (O_2183,N_19850,N_19817);
or UO_2184 (O_2184,N_18458,N_18748);
nand UO_2185 (O_2185,N_19483,N_19482);
nor UO_2186 (O_2186,N_19058,N_19388);
and UO_2187 (O_2187,N_19042,N_18176);
and UO_2188 (O_2188,N_19959,N_18775);
or UO_2189 (O_2189,N_19306,N_18391);
nor UO_2190 (O_2190,N_19837,N_19866);
nand UO_2191 (O_2191,N_18365,N_19943);
nand UO_2192 (O_2192,N_18362,N_19929);
xnor UO_2193 (O_2193,N_18000,N_18406);
and UO_2194 (O_2194,N_18801,N_18594);
or UO_2195 (O_2195,N_18514,N_18200);
nand UO_2196 (O_2196,N_19064,N_19087);
nor UO_2197 (O_2197,N_19589,N_19976);
or UO_2198 (O_2198,N_18258,N_18039);
xnor UO_2199 (O_2199,N_19227,N_18767);
or UO_2200 (O_2200,N_19333,N_19643);
and UO_2201 (O_2201,N_18476,N_18488);
or UO_2202 (O_2202,N_18570,N_18675);
and UO_2203 (O_2203,N_19988,N_19874);
nor UO_2204 (O_2204,N_18287,N_19058);
nand UO_2205 (O_2205,N_18048,N_18333);
and UO_2206 (O_2206,N_19571,N_19073);
nand UO_2207 (O_2207,N_19228,N_19866);
xnor UO_2208 (O_2208,N_19753,N_18664);
nand UO_2209 (O_2209,N_18499,N_18417);
nor UO_2210 (O_2210,N_19857,N_18754);
nor UO_2211 (O_2211,N_19564,N_19541);
xnor UO_2212 (O_2212,N_18208,N_19562);
nor UO_2213 (O_2213,N_18086,N_18242);
and UO_2214 (O_2214,N_18522,N_19813);
nand UO_2215 (O_2215,N_19024,N_19665);
nor UO_2216 (O_2216,N_18204,N_19498);
or UO_2217 (O_2217,N_19712,N_18760);
and UO_2218 (O_2218,N_18929,N_18007);
or UO_2219 (O_2219,N_19233,N_18878);
nor UO_2220 (O_2220,N_19806,N_18004);
or UO_2221 (O_2221,N_18008,N_19381);
nand UO_2222 (O_2222,N_19151,N_18503);
nand UO_2223 (O_2223,N_19314,N_18821);
and UO_2224 (O_2224,N_18232,N_19296);
xnor UO_2225 (O_2225,N_19050,N_19422);
or UO_2226 (O_2226,N_19907,N_19716);
nand UO_2227 (O_2227,N_18403,N_19386);
or UO_2228 (O_2228,N_18882,N_18904);
xnor UO_2229 (O_2229,N_18953,N_19405);
nand UO_2230 (O_2230,N_19200,N_18279);
nor UO_2231 (O_2231,N_19752,N_18706);
nor UO_2232 (O_2232,N_18993,N_18887);
nor UO_2233 (O_2233,N_18365,N_19143);
xor UO_2234 (O_2234,N_18974,N_18049);
xor UO_2235 (O_2235,N_19930,N_19249);
and UO_2236 (O_2236,N_18203,N_19376);
nand UO_2237 (O_2237,N_19851,N_18601);
xor UO_2238 (O_2238,N_18911,N_19008);
nor UO_2239 (O_2239,N_18272,N_19939);
xnor UO_2240 (O_2240,N_19970,N_18743);
nand UO_2241 (O_2241,N_19846,N_18998);
and UO_2242 (O_2242,N_19099,N_18916);
nand UO_2243 (O_2243,N_18712,N_19033);
and UO_2244 (O_2244,N_19180,N_18174);
nor UO_2245 (O_2245,N_19772,N_19357);
and UO_2246 (O_2246,N_18686,N_18161);
and UO_2247 (O_2247,N_19225,N_19354);
xor UO_2248 (O_2248,N_18380,N_19765);
nor UO_2249 (O_2249,N_18864,N_19618);
or UO_2250 (O_2250,N_18197,N_18489);
and UO_2251 (O_2251,N_18975,N_19599);
nand UO_2252 (O_2252,N_19569,N_19272);
or UO_2253 (O_2253,N_18400,N_18308);
nand UO_2254 (O_2254,N_19347,N_18219);
or UO_2255 (O_2255,N_19657,N_18269);
xor UO_2256 (O_2256,N_19292,N_19904);
and UO_2257 (O_2257,N_19402,N_19168);
xnor UO_2258 (O_2258,N_18318,N_18312);
and UO_2259 (O_2259,N_18898,N_18682);
xnor UO_2260 (O_2260,N_18956,N_18444);
xnor UO_2261 (O_2261,N_19679,N_19672);
or UO_2262 (O_2262,N_19882,N_19018);
xnor UO_2263 (O_2263,N_18771,N_19793);
nor UO_2264 (O_2264,N_19972,N_19950);
xor UO_2265 (O_2265,N_18776,N_18566);
or UO_2266 (O_2266,N_18848,N_19628);
and UO_2267 (O_2267,N_19706,N_18273);
xor UO_2268 (O_2268,N_19258,N_19563);
and UO_2269 (O_2269,N_18054,N_19649);
xnor UO_2270 (O_2270,N_18296,N_18693);
xor UO_2271 (O_2271,N_18028,N_18483);
and UO_2272 (O_2272,N_18263,N_19916);
nand UO_2273 (O_2273,N_18630,N_18011);
and UO_2274 (O_2274,N_19927,N_18061);
nor UO_2275 (O_2275,N_19649,N_18972);
nand UO_2276 (O_2276,N_18092,N_19492);
nor UO_2277 (O_2277,N_18911,N_19170);
or UO_2278 (O_2278,N_18728,N_18777);
xor UO_2279 (O_2279,N_18138,N_19718);
nand UO_2280 (O_2280,N_18701,N_19269);
xor UO_2281 (O_2281,N_19949,N_18153);
nor UO_2282 (O_2282,N_18906,N_18890);
nor UO_2283 (O_2283,N_18987,N_18383);
or UO_2284 (O_2284,N_19893,N_18347);
or UO_2285 (O_2285,N_19742,N_18733);
nor UO_2286 (O_2286,N_18047,N_18543);
nand UO_2287 (O_2287,N_18818,N_19120);
xnor UO_2288 (O_2288,N_19270,N_18932);
or UO_2289 (O_2289,N_19555,N_18189);
nand UO_2290 (O_2290,N_19494,N_18861);
xnor UO_2291 (O_2291,N_19364,N_19565);
nor UO_2292 (O_2292,N_19458,N_18034);
xor UO_2293 (O_2293,N_18210,N_18403);
or UO_2294 (O_2294,N_19041,N_18896);
or UO_2295 (O_2295,N_18395,N_19074);
and UO_2296 (O_2296,N_19564,N_18670);
nand UO_2297 (O_2297,N_19924,N_18870);
nor UO_2298 (O_2298,N_19330,N_19658);
nor UO_2299 (O_2299,N_18551,N_18533);
xor UO_2300 (O_2300,N_18817,N_18898);
xnor UO_2301 (O_2301,N_19856,N_19297);
nand UO_2302 (O_2302,N_18876,N_19525);
xor UO_2303 (O_2303,N_18563,N_18499);
nor UO_2304 (O_2304,N_19411,N_18662);
xor UO_2305 (O_2305,N_19900,N_18450);
nand UO_2306 (O_2306,N_19452,N_18876);
nand UO_2307 (O_2307,N_19819,N_19180);
nor UO_2308 (O_2308,N_18382,N_18202);
xnor UO_2309 (O_2309,N_19826,N_19810);
xor UO_2310 (O_2310,N_18581,N_19100);
nand UO_2311 (O_2311,N_19288,N_18962);
nor UO_2312 (O_2312,N_18301,N_19976);
or UO_2313 (O_2313,N_19590,N_18233);
or UO_2314 (O_2314,N_18127,N_19999);
nand UO_2315 (O_2315,N_18178,N_18151);
xor UO_2316 (O_2316,N_19544,N_18877);
xor UO_2317 (O_2317,N_18494,N_18392);
or UO_2318 (O_2318,N_19089,N_18419);
nor UO_2319 (O_2319,N_19047,N_19818);
nor UO_2320 (O_2320,N_18810,N_19452);
nand UO_2321 (O_2321,N_18381,N_19034);
or UO_2322 (O_2322,N_18285,N_18048);
nand UO_2323 (O_2323,N_18587,N_19152);
xnor UO_2324 (O_2324,N_19132,N_18490);
nand UO_2325 (O_2325,N_19326,N_19301);
or UO_2326 (O_2326,N_19175,N_18994);
nor UO_2327 (O_2327,N_18165,N_19855);
nor UO_2328 (O_2328,N_19428,N_18805);
nand UO_2329 (O_2329,N_18625,N_19157);
nand UO_2330 (O_2330,N_18325,N_19386);
and UO_2331 (O_2331,N_18831,N_19295);
or UO_2332 (O_2332,N_18066,N_19948);
xnor UO_2333 (O_2333,N_19875,N_19105);
nand UO_2334 (O_2334,N_18305,N_19940);
or UO_2335 (O_2335,N_19488,N_19572);
or UO_2336 (O_2336,N_18151,N_19375);
and UO_2337 (O_2337,N_19302,N_18663);
and UO_2338 (O_2338,N_18766,N_18938);
nor UO_2339 (O_2339,N_18789,N_18113);
nor UO_2340 (O_2340,N_19803,N_19413);
or UO_2341 (O_2341,N_18095,N_18525);
nor UO_2342 (O_2342,N_18652,N_19531);
and UO_2343 (O_2343,N_18899,N_19604);
and UO_2344 (O_2344,N_18011,N_19056);
xnor UO_2345 (O_2345,N_19602,N_19973);
nor UO_2346 (O_2346,N_18591,N_18612);
and UO_2347 (O_2347,N_18167,N_18032);
nand UO_2348 (O_2348,N_19996,N_19998);
xor UO_2349 (O_2349,N_18152,N_19663);
xnor UO_2350 (O_2350,N_19097,N_19343);
nor UO_2351 (O_2351,N_18290,N_19008);
and UO_2352 (O_2352,N_18714,N_19102);
and UO_2353 (O_2353,N_19524,N_19905);
or UO_2354 (O_2354,N_18532,N_18968);
xor UO_2355 (O_2355,N_18312,N_18996);
nor UO_2356 (O_2356,N_18041,N_19026);
nand UO_2357 (O_2357,N_19337,N_18387);
and UO_2358 (O_2358,N_19224,N_18089);
or UO_2359 (O_2359,N_18963,N_19709);
and UO_2360 (O_2360,N_19389,N_18646);
nand UO_2361 (O_2361,N_19962,N_18621);
or UO_2362 (O_2362,N_18324,N_19388);
and UO_2363 (O_2363,N_19608,N_19744);
or UO_2364 (O_2364,N_19638,N_18796);
and UO_2365 (O_2365,N_18757,N_19234);
and UO_2366 (O_2366,N_18567,N_18893);
xor UO_2367 (O_2367,N_18619,N_19811);
nor UO_2368 (O_2368,N_19840,N_18800);
xnor UO_2369 (O_2369,N_18593,N_18544);
xnor UO_2370 (O_2370,N_18223,N_19527);
nor UO_2371 (O_2371,N_19047,N_18224);
xnor UO_2372 (O_2372,N_18957,N_18719);
or UO_2373 (O_2373,N_19422,N_18923);
and UO_2374 (O_2374,N_19843,N_19765);
or UO_2375 (O_2375,N_19076,N_19844);
and UO_2376 (O_2376,N_19293,N_19162);
nor UO_2377 (O_2377,N_18466,N_19905);
and UO_2378 (O_2378,N_18991,N_19935);
or UO_2379 (O_2379,N_18429,N_19268);
and UO_2380 (O_2380,N_19359,N_19748);
or UO_2381 (O_2381,N_18002,N_19426);
and UO_2382 (O_2382,N_18152,N_18470);
xor UO_2383 (O_2383,N_19871,N_19563);
or UO_2384 (O_2384,N_19314,N_18195);
or UO_2385 (O_2385,N_19240,N_18939);
and UO_2386 (O_2386,N_18562,N_19940);
nor UO_2387 (O_2387,N_18666,N_19075);
nor UO_2388 (O_2388,N_18383,N_18346);
xor UO_2389 (O_2389,N_18015,N_18803);
and UO_2390 (O_2390,N_18482,N_18760);
and UO_2391 (O_2391,N_18759,N_18530);
xor UO_2392 (O_2392,N_19226,N_18008);
nor UO_2393 (O_2393,N_19474,N_19092);
or UO_2394 (O_2394,N_18161,N_18070);
nor UO_2395 (O_2395,N_18286,N_19715);
nand UO_2396 (O_2396,N_18534,N_19743);
and UO_2397 (O_2397,N_19149,N_19427);
xor UO_2398 (O_2398,N_19172,N_19305);
nor UO_2399 (O_2399,N_18954,N_19370);
nor UO_2400 (O_2400,N_19227,N_19399);
xnor UO_2401 (O_2401,N_18813,N_18173);
nand UO_2402 (O_2402,N_18618,N_19103);
nand UO_2403 (O_2403,N_18369,N_19766);
and UO_2404 (O_2404,N_18547,N_19166);
and UO_2405 (O_2405,N_18476,N_19197);
nor UO_2406 (O_2406,N_19059,N_19990);
and UO_2407 (O_2407,N_18281,N_19231);
xnor UO_2408 (O_2408,N_19629,N_18145);
nand UO_2409 (O_2409,N_19848,N_19658);
or UO_2410 (O_2410,N_19233,N_18056);
xnor UO_2411 (O_2411,N_18090,N_19659);
and UO_2412 (O_2412,N_18795,N_19441);
and UO_2413 (O_2413,N_18600,N_18386);
xnor UO_2414 (O_2414,N_18082,N_18334);
or UO_2415 (O_2415,N_18477,N_18507);
nor UO_2416 (O_2416,N_18911,N_19719);
and UO_2417 (O_2417,N_19250,N_19480);
or UO_2418 (O_2418,N_19375,N_19262);
xor UO_2419 (O_2419,N_18025,N_18792);
xor UO_2420 (O_2420,N_19109,N_19302);
xor UO_2421 (O_2421,N_19749,N_18034);
or UO_2422 (O_2422,N_19719,N_19466);
nor UO_2423 (O_2423,N_19867,N_19121);
nand UO_2424 (O_2424,N_18359,N_19036);
nor UO_2425 (O_2425,N_19228,N_18084);
or UO_2426 (O_2426,N_18664,N_18313);
or UO_2427 (O_2427,N_18435,N_18655);
or UO_2428 (O_2428,N_18328,N_18598);
or UO_2429 (O_2429,N_19182,N_18253);
xor UO_2430 (O_2430,N_19029,N_18456);
or UO_2431 (O_2431,N_18745,N_19697);
and UO_2432 (O_2432,N_19000,N_19564);
xnor UO_2433 (O_2433,N_19724,N_18442);
xor UO_2434 (O_2434,N_19462,N_18703);
and UO_2435 (O_2435,N_18121,N_19176);
and UO_2436 (O_2436,N_18649,N_18658);
nor UO_2437 (O_2437,N_19677,N_19122);
nand UO_2438 (O_2438,N_18162,N_18607);
and UO_2439 (O_2439,N_19516,N_19386);
or UO_2440 (O_2440,N_19908,N_18590);
xnor UO_2441 (O_2441,N_18008,N_18734);
xnor UO_2442 (O_2442,N_19420,N_18235);
and UO_2443 (O_2443,N_18750,N_18059);
and UO_2444 (O_2444,N_18774,N_19307);
and UO_2445 (O_2445,N_19028,N_19505);
or UO_2446 (O_2446,N_19095,N_19969);
nand UO_2447 (O_2447,N_19097,N_19749);
nand UO_2448 (O_2448,N_18824,N_18518);
or UO_2449 (O_2449,N_18988,N_19836);
and UO_2450 (O_2450,N_19065,N_19010);
nor UO_2451 (O_2451,N_19850,N_18916);
nand UO_2452 (O_2452,N_18777,N_18013);
and UO_2453 (O_2453,N_18486,N_18556);
xor UO_2454 (O_2454,N_18200,N_19576);
nand UO_2455 (O_2455,N_19213,N_18383);
xnor UO_2456 (O_2456,N_19165,N_18593);
nor UO_2457 (O_2457,N_19627,N_19574);
or UO_2458 (O_2458,N_18935,N_18873);
or UO_2459 (O_2459,N_19481,N_18343);
xnor UO_2460 (O_2460,N_19423,N_18472);
and UO_2461 (O_2461,N_18180,N_19089);
or UO_2462 (O_2462,N_19791,N_18950);
or UO_2463 (O_2463,N_18679,N_19920);
and UO_2464 (O_2464,N_18038,N_18628);
or UO_2465 (O_2465,N_18844,N_18565);
and UO_2466 (O_2466,N_19732,N_18088);
or UO_2467 (O_2467,N_18941,N_19357);
and UO_2468 (O_2468,N_19526,N_19890);
xor UO_2469 (O_2469,N_18889,N_19606);
nor UO_2470 (O_2470,N_18873,N_18201);
and UO_2471 (O_2471,N_18240,N_18050);
and UO_2472 (O_2472,N_19906,N_19051);
and UO_2473 (O_2473,N_18016,N_19916);
nor UO_2474 (O_2474,N_18968,N_18951);
nand UO_2475 (O_2475,N_18257,N_18974);
nand UO_2476 (O_2476,N_18223,N_19900);
and UO_2477 (O_2477,N_19457,N_19935);
or UO_2478 (O_2478,N_18648,N_18633);
xnor UO_2479 (O_2479,N_18352,N_19878);
nand UO_2480 (O_2480,N_18149,N_19914);
nor UO_2481 (O_2481,N_19354,N_18760);
xnor UO_2482 (O_2482,N_18014,N_18421);
xor UO_2483 (O_2483,N_19814,N_19640);
nand UO_2484 (O_2484,N_18663,N_19502);
or UO_2485 (O_2485,N_18707,N_19021);
nor UO_2486 (O_2486,N_18741,N_18057);
nand UO_2487 (O_2487,N_18035,N_19979);
nand UO_2488 (O_2488,N_19689,N_19268);
or UO_2489 (O_2489,N_18199,N_18314);
or UO_2490 (O_2490,N_18262,N_19808);
xnor UO_2491 (O_2491,N_19383,N_18059);
xnor UO_2492 (O_2492,N_19917,N_19707);
or UO_2493 (O_2493,N_18923,N_18165);
nor UO_2494 (O_2494,N_19947,N_19224);
and UO_2495 (O_2495,N_19190,N_18022);
xnor UO_2496 (O_2496,N_18498,N_19457);
or UO_2497 (O_2497,N_19850,N_18543);
or UO_2498 (O_2498,N_19121,N_18534);
and UO_2499 (O_2499,N_19825,N_18863);
endmodule