module basic_500_3000_500_50_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_253,In_7);
or U1 (N_1,In_469,In_490);
and U2 (N_2,In_224,In_42);
and U3 (N_3,In_291,In_105);
nand U4 (N_4,In_242,In_416);
and U5 (N_5,In_395,In_399);
and U6 (N_6,In_166,In_362);
and U7 (N_7,In_431,In_27);
and U8 (N_8,In_10,In_491);
or U9 (N_9,In_227,In_121);
and U10 (N_10,In_355,In_363);
or U11 (N_11,In_436,In_71);
or U12 (N_12,In_422,In_251);
and U13 (N_13,In_204,In_111);
or U14 (N_14,In_454,In_290);
or U15 (N_15,In_228,In_384);
nor U16 (N_16,In_274,In_2);
nand U17 (N_17,In_225,In_243);
and U18 (N_18,In_137,In_221);
nand U19 (N_19,In_34,In_223);
xnor U20 (N_20,In_423,In_350);
and U21 (N_21,In_18,In_282);
xnor U22 (N_22,In_284,In_323);
and U23 (N_23,In_39,In_267);
or U24 (N_24,In_307,In_13);
and U25 (N_25,In_463,In_161);
or U26 (N_26,In_180,In_73);
and U27 (N_27,In_75,In_257);
xor U28 (N_28,In_96,In_170);
and U29 (N_29,In_114,In_345);
nor U30 (N_30,In_460,In_88);
or U31 (N_31,In_182,In_474);
and U32 (N_32,In_276,In_342);
nor U33 (N_33,In_373,In_210);
nor U34 (N_34,In_91,In_132);
nor U35 (N_35,In_53,In_92);
or U36 (N_36,In_277,In_354);
nand U37 (N_37,In_478,In_25);
nand U38 (N_38,In_179,In_472);
nor U39 (N_39,In_237,In_32);
nand U40 (N_40,In_101,In_29);
and U41 (N_41,In_112,In_434);
nor U42 (N_42,In_409,In_181);
and U43 (N_43,In_299,In_167);
nand U44 (N_44,In_270,In_459);
or U45 (N_45,In_364,In_231);
nand U46 (N_46,In_293,In_370);
nor U47 (N_47,In_216,In_497);
nor U48 (N_48,In_302,In_286);
or U49 (N_49,In_489,In_326);
nand U50 (N_50,In_184,In_470);
or U51 (N_51,In_341,In_99);
nand U52 (N_52,In_209,In_448);
and U53 (N_53,In_402,In_318);
nor U54 (N_54,In_58,In_427);
nand U55 (N_55,In_68,In_174);
nand U56 (N_56,In_313,In_393);
nor U57 (N_57,In_254,In_70);
nand U58 (N_58,In_109,In_337);
nand U59 (N_59,In_213,In_201);
nor U60 (N_60,In_211,In_455);
nor U61 (N_61,In_76,In_433);
or U62 (N_62,In_205,In_406);
nor U63 (N_63,In_330,In_273);
nor U64 (N_64,In_141,In_259);
nor U65 (N_65,In_100,In_155);
nor U66 (N_66,N_39,In_171);
nand U67 (N_67,In_61,In_429);
nand U68 (N_68,In_21,In_298);
nor U69 (N_69,In_308,In_106);
xor U70 (N_70,N_9,In_415);
or U71 (N_71,In_206,In_312);
or U72 (N_72,In_360,In_336);
nand U73 (N_73,In_5,In_359);
and U74 (N_74,In_219,In_482);
and U75 (N_75,In_378,In_374);
and U76 (N_76,In_28,N_34);
or U77 (N_77,In_388,N_31);
or U78 (N_78,In_410,In_98);
or U79 (N_79,In_240,N_42);
and U80 (N_80,In_80,In_120);
and U81 (N_81,In_315,In_306);
nor U82 (N_82,In_339,In_102);
nor U83 (N_83,In_380,In_115);
and U84 (N_84,In_493,In_450);
or U85 (N_85,In_22,In_208);
or U86 (N_86,In_165,In_218);
and U87 (N_87,In_122,N_49);
nor U88 (N_88,In_54,In_325);
xor U89 (N_89,In_371,In_358);
and U90 (N_90,In_94,In_62);
or U91 (N_91,N_58,In_3);
or U92 (N_92,N_18,N_4);
nand U93 (N_93,In_351,In_334);
and U94 (N_94,N_33,In_63);
or U95 (N_95,In_485,In_379);
nor U96 (N_96,In_258,In_239);
or U97 (N_97,In_142,In_456);
nor U98 (N_98,In_348,In_66);
and U99 (N_99,In_191,In_278);
or U100 (N_100,In_249,In_139);
and U101 (N_101,In_81,In_496);
or U102 (N_102,N_44,In_300);
nand U103 (N_103,In_499,In_382);
nor U104 (N_104,In_473,In_294);
nor U105 (N_105,In_133,In_391);
nand U106 (N_106,N_27,In_344);
or U107 (N_107,In_156,In_432);
or U108 (N_108,In_397,In_245);
and U109 (N_109,N_14,In_262);
xor U110 (N_110,In_435,In_30);
and U111 (N_111,In_26,In_11);
and U112 (N_112,In_495,In_305);
or U113 (N_113,In_420,In_458);
or U114 (N_114,In_494,In_439);
and U115 (N_115,N_56,In_60);
nand U116 (N_116,In_38,In_126);
nor U117 (N_117,N_3,In_387);
and U118 (N_118,N_7,In_236);
and U119 (N_119,In_215,In_84);
or U120 (N_120,In_235,In_361);
or U121 (N_121,In_16,In_83);
nor U122 (N_122,In_197,In_449);
and U123 (N_123,N_50,In_214);
nor U124 (N_124,In_9,In_193);
or U125 (N_125,In_173,In_346);
and U126 (N_126,In_95,In_479);
nor U127 (N_127,In_189,N_46);
and U128 (N_128,In_125,In_385);
nand U129 (N_129,N_91,In_220);
nor U130 (N_130,In_368,N_55);
and U131 (N_131,In_404,In_104);
or U132 (N_132,N_53,In_401);
nor U133 (N_133,In_176,In_281);
nor U134 (N_134,In_481,In_78);
nand U135 (N_135,N_70,In_64);
and U136 (N_136,N_117,In_110);
nor U137 (N_137,In_244,In_107);
nand U138 (N_138,In_357,In_116);
or U139 (N_139,In_241,N_108);
or U140 (N_140,In_56,In_8);
nand U141 (N_141,In_272,N_116);
nor U142 (N_142,N_37,In_314);
nor U143 (N_143,In_202,In_430);
nand U144 (N_144,In_1,N_96);
nand U145 (N_145,In_252,N_2);
or U146 (N_146,N_61,In_295);
nor U147 (N_147,In_266,In_175);
nor U148 (N_148,In_353,In_400);
and U149 (N_149,N_15,In_288);
or U150 (N_150,In_263,In_292);
nand U151 (N_151,In_418,In_349);
nor U152 (N_152,In_203,In_199);
nand U153 (N_153,In_198,N_79);
nor U154 (N_154,In_50,In_413);
or U155 (N_155,In_261,In_452);
and U156 (N_156,In_367,N_65);
nand U157 (N_157,N_102,In_123);
or U158 (N_158,In_335,N_5);
nor U159 (N_159,N_118,N_20);
or U160 (N_160,N_23,In_289);
or U161 (N_161,N_104,In_285);
nand U162 (N_162,N_115,N_41);
nand U163 (N_163,In_152,In_117);
and U164 (N_164,In_322,In_394);
nand U165 (N_165,In_327,In_160);
nor U166 (N_166,In_466,In_19);
and U167 (N_167,In_147,N_67);
nand U168 (N_168,In_408,In_383);
and U169 (N_169,In_301,N_95);
nor U170 (N_170,N_51,In_453);
nor U171 (N_171,In_398,In_333);
or U172 (N_172,In_407,In_366);
nand U173 (N_173,In_6,In_85);
and U174 (N_174,In_12,In_309);
nor U175 (N_175,In_138,N_63);
nor U176 (N_176,In_169,In_149);
nand U177 (N_177,In_69,In_287);
nor U178 (N_178,N_75,In_465);
and U179 (N_179,In_477,In_36);
and U180 (N_180,In_119,In_74);
or U181 (N_181,In_185,In_338);
or U182 (N_182,In_157,In_372);
nor U183 (N_183,N_82,N_8);
nand U184 (N_184,N_12,In_48);
or U185 (N_185,In_194,In_47);
and U186 (N_186,In_24,N_13);
nand U187 (N_187,In_77,In_303);
nand U188 (N_188,In_212,N_103);
and U189 (N_189,N_73,N_134);
nor U190 (N_190,N_119,In_178);
or U191 (N_191,In_238,In_381);
nand U192 (N_192,In_424,In_15);
and U193 (N_193,N_101,N_35);
and U194 (N_194,In_234,In_438);
xnor U195 (N_195,N_133,N_124);
and U196 (N_196,In_49,N_94);
nand U197 (N_197,N_161,In_46);
nand U198 (N_198,N_16,N_145);
nor U199 (N_199,N_57,N_110);
nand U200 (N_200,N_76,In_352);
and U201 (N_201,N_156,In_467);
or U202 (N_202,In_396,In_414);
and U203 (N_203,In_283,In_340);
or U204 (N_204,In_154,In_0);
nor U205 (N_205,N_36,In_124);
nand U206 (N_206,N_25,In_67);
nor U207 (N_207,In_37,N_81);
and U208 (N_208,In_457,N_141);
and U209 (N_209,In_190,N_17);
nor U210 (N_210,In_444,In_331);
nor U211 (N_211,N_85,In_72);
and U212 (N_212,In_20,In_128);
nand U213 (N_213,N_136,In_475);
and U214 (N_214,In_51,In_43);
nor U215 (N_215,N_90,In_375);
and U216 (N_216,In_144,In_377);
nand U217 (N_217,In_140,In_230);
nand U218 (N_218,N_172,In_89);
and U219 (N_219,In_172,In_412);
nand U220 (N_220,N_99,N_129);
and U221 (N_221,N_84,In_311);
nand U222 (N_222,N_120,In_268);
or U223 (N_223,N_174,In_164);
or U224 (N_224,In_476,N_64);
or U225 (N_225,N_143,N_140);
xor U226 (N_226,In_498,N_128);
or U227 (N_227,N_123,N_159);
or U228 (N_228,In_127,In_87);
nor U229 (N_229,In_163,In_40);
nor U230 (N_230,In_369,N_0);
and U231 (N_231,N_69,N_158);
and U232 (N_232,In_279,N_97);
and U233 (N_233,In_343,In_296);
nand U234 (N_234,N_77,N_131);
nor U235 (N_235,In_134,In_462);
and U236 (N_236,N_157,In_419);
and U237 (N_237,N_6,N_176);
nand U238 (N_238,In_447,N_113);
or U239 (N_239,N_164,In_14);
xor U240 (N_240,N_130,In_390);
nand U241 (N_241,N_199,N_86);
nor U242 (N_242,In_44,N_144);
or U243 (N_243,N_151,In_192);
and U244 (N_244,In_17,In_442);
nand U245 (N_245,N_29,In_250);
or U246 (N_246,N_216,N_59);
or U247 (N_247,N_232,In_59);
nand U248 (N_248,In_183,In_484);
or U249 (N_249,In_275,In_403);
or U250 (N_250,N_109,N_155);
nand U251 (N_251,N_32,In_389);
or U252 (N_252,In_97,N_218);
nor U253 (N_253,N_211,In_188);
nand U254 (N_254,N_221,N_47);
nor U255 (N_255,N_88,N_173);
and U256 (N_256,In_153,In_145);
and U257 (N_257,In_222,In_23);
nand U258 (N_258,N_80,N_206);
nor U259 (N_259,In_280,In_269);
nand U260 (N_260,N_40,N_193);
nor U261 (N_261,N_45,N_114);
and U262 (N_262,In_65,N_19);
nand U263 (N_263,In_332,In_437);
nand U264 (N_264,In_411,In_187);
nor U265 (N_265,N_87,N_62);
or U266 (N_266,In_159,N_239);
and U267 (N_267,In_451,N_201);
nor U268 (N_268,N_78,N_89);
and U269 (N_269,N_183,N_150);
nand U270 (N_270,N_160,N_204);
and U271 (N_271,N_222,N_83);
nand U272 (N_272,N_233,In_196);
and U273 (N_273,N_213,N_190);
nor U274 (N_274,N_163,N_30);
nor U275 (N_275,In_445,N_138);
nor U276 (N_276,N_217,N_209);
nand U277 (N_277,In_31,N_228);
nand U278 (N_278,N_142,N_238);
nand U279 (N_279,In_405,In_229);
nor U280 (N_280,In_417,In_264);
nor U281 (N_281,N_184,N_167);
and U282 (N_282,In_90,In_151);
nand U283 (N_283,In_392,In_135);
and U284 (N_284,N_181,N_179);
or U285 (N_285,N_169,In_324);
nand U286 (N_286,N_139,In_186);
or U287 (N_287,In_486,In_246);
or U288 (N_288,N_212,In_55);
nand U289 (N_289,N_71,In_82);
nor U290 (N_290,In_440,N_214);
nand U291 (N_291,N_147,N_122);
nand U292 (N_292,N_178,N_191);
and U293 (N_293,N_162,N_166);
or U294 (N_294,In_260,N_66);
nor U295 (N_295,N_175,In_41);
nand U296 (N_296,N_48,N_135);
nor U297 (N_297,In_162,In_265);
nor U298 (N_298,N_126,In_57);
or U299 (N_299,In_195,In_441);
nand U300 (N_300,N_168,N_52);
or U301 (N_301,N_262,N_298);
nor U302 (N_302,N_286,N_272);
nand U303 (N_303,N_182,N_220);
and U304 (N_304,N_273,In_130);
nor U305 (N_305,N_250,N_254);
or U306 (N_306,In_468,N_282);
nand U307 (N_307,In_207,N_259);
and U308 (N_308,N_92,N_68);
and U309 (N_309,N_149,N_121);
nor U310 (N_310,N_264,N_185);
and U311 (N_311,N_188,N_279);
and U312 (N_312,In_428,N_281);
xnor U313 (N_313,N_285,In_426);
nand U314 (N_314,N_287,N_292);
xor U315 (N_315,In_446,N_219);
or U316 (N_316,In_487,N_268);
nand U317 (N_317,N_43,In_113);
and U318 (N_318,N_277,N_11);
and U319 (N_319,N_255,N_112);
nor U320 (N_320,N_165,In_316);
nand U321 (N_321,N_171,In_271);
nor U322 (N_322,N_106,In_319);
and U323 (N_323,N_54,In_129);
nand U324 (N_324,In_226,N_297);
nand U325 (N_325,N_275,N_291);
nor U326 (N_326,N_207,N_241);
nor U327 (N_327,N_98,N_240);
nor U328 (N_328,N_295,N_153);
nor U329 (N_329,N_263,N_229);
xnor U330 (N_330,N_274,N_284);
and U331 (N_331,In_480,N_290);
xnor U332 (N_332,In_200,N_215);
nor U333 (N_333,N_245,N_177);
and U334 (N_334,N_107,N_247);
nand U335 (N_335,In_256,In_425);
nor U336 (N_336,N_195,N_252);
and U337 (N_337,N_28,In_304);
nand U338 (N_338,In_386,In_421);
nor U339 (N_339,In_317,In_33);
and U340 (N_340,In_365,N_186);
nand U341 (N_341,In_328,N_137);
or U342 (N_342,N_289,N_203);
nand U343 (N_343,N_296,N_170);
xnor U344 (N_344,In_45,N_251);
nor U345 (N_345,N_271,N_223);
nand U346 (N_346,In_232,N_100);
or U347 (N_347,In_233,N_198);
or U348 (N_348,In_131,In_168);
xnor U349 (N_349,N_243,N_246);
nand U350 (N_350,In_158,In_488);
nand U351 (N_351,N_24,N_154);
and U352 (N_352,N_132,N_205);
or U353 (N_353,In_86,In_320);
nand U354 (N_354,N_127,In_356);
nor U355 (N_355,N_74,In_255);
and U356 (N_356,N_265,In_247);
nor U357 (N_357,N_261,N_280);
nand U358 (N_358,In_35,N_236);
and U359 (N_359,N_200,N_225);
or U360 (N_360,N_329,In_148);
nor U361 (N_361,N_315,N_231);
or U362 (N_362,In_143,N_301);
nand U363 (N_363,N_316,In_177);
nand U364 (N_364,N_302,N_111);
or U365 (N_365,In_310,In_79);
nor U366 (N_366,N_260,N_343);
and U367 (N_367,N_189,N_346);
and U368 (N_368,N_347,N_253);
or U369 (N_369,N_334,N_359);
or U370 (N_370,N_326,N_354);
and U371 (N_371,N_21,N_257);
nand U372 (N_372,In_464,In_329);
and U373 (N_373,N_72,In_217);
nand U374 (N_374,N_105,N_93);
nor U375 (N_375,In_347,In_248);
or U376 (N_376,N_336,N_305);
and U377 (N_377,N_269,N_356);
nand U378 (N_378,N_26,N_202);
nor U379 (N_379,N_303,N_349);
or U380 (N_380,N_249,In_150);
nand U381 (N_381,N_267,N_266);
and U382 (N_382,N_306,N_60);
nand U383 (N_383,N_320,N_324);
nand U384 (N_384,In_93,N_283);
and U385 (N_385,In_321,N_317);
and U386 (N_386,N_148,N_300);
or U387 (N_387,N_332,N_196);
nand U388 (N_388,N_180,In_103);
nand U389 (N_389,N_333,N_321);
and U390 (N_390,N_22,N_288);
nand U391 (N_391,N_234,In_376);
nand U392 (N_392,N_327,In_108);
and U393 (N_393,N_348,N_325);
nand U394 (N_394,In_146,N_210);
nor U395 (N_395,N_350,N_337);
or U396 (N_396,In_136,N_248);
and U397 (N_397,N_319,N_278);
and U398 (N_398,In_461,In_52);
and U399 (N_399,N_353,In_297);
and U400 (N_400,N_197,N_1);
or U401 (N_401,N_323,N_351);
and U402 (N_402,N_358,In_118);
nand U403 (N_403,N_187,N_293);
nand U404 (N_404,N_313,N_10);
and U405 (N_405,N_330,N_322);
and U406 (N_406,In_4,N_308);
nor U407 (N_407,In_492,In_471);
nor U408 (N_408,N_256,N_357);
and U409 (N_409,N_152,N_331);
or U410 (N_410,N_340,N_258);
and U411 (N_411,N_270,N_224);
nand U412 (N_412,N_125,N_299);
nand U413 (N_413,N_318,N_338);
nand U414 (N_414,N_146,N_355);
or U415 (N_415,N_235,N_328);
nor U416 (N_416,N_311,N_192);
nor U417 (N_417,N_309,N_208);
or U418 (N_418,N_242,N_244);
or U419 (N_419,N_230,N_276);
nand U420 (N_420,In_483,N_383);
and U421 (N_421,N_361,N_400);
or U422 (N_422,N_371,N_404);
nand U423 (N_423,N_352,N_341);
or U424 (N_424,N_389,N_385);
xnor U425 (N_425,N_307,N_374);
nor U426 (N_426,N_344,N_393);
nand U427 (N_427,N_413,N_418);
and U428 (N_428,N_412,N_360);
or U429 (N_429,N_339,N_401);
xor U430 (N_430,N_226,N_386);
nand U431 (N_431,N_391,N_382);
nor U432 (N_432,N_407,N_342);
nor U433 (N_433,N_376,N_417);
and U434 (N_434,N_414,N_384);
nand U435 (N_435,N_409,N_304);
or U436 (N_436,N_310,N_408);
nor U437 (N_437,N_373,N_377);
and U438 (N_438,N_365,N_411);
or U439 (N_439,N_345,N_399);
nor U440 (N_440,N_394,N_392);
or U441 (N_441,N_415,N_406);
and U442 (N_442,N_388,N_370);
and U443 (N_443,N_405,N_314);
nand U444 (N_444,N_368,N_403);
and U445 (N_445,N_419,N_397);
nand U446 (N_446,N_367,N_380);
nand U447 (N_447,N_395,N_194);
nor U448 (N_448,N_366,N_396);
nor U449 (N_449,N_379,In_443);
or U450 (N_450,N_378,N_38);
nand U451 (N_451,N_416,N_387);
and U452 (N_452,N_335,N_312);
or U453 (N_453,N_369,N_398);
nand U454 (N_454,N_381,N_363);
and U455 (N_455,N_402,N_364);
nand U456 (N_456,N_375,N_237);
or U457 (N_457,N_410,N_362);
or U458 (N_458,N_294,N_372);
nor U459 (N_459,N_390,N_227);
or U460 (N_460,N_369,N_415);
nand U461 (N_461,N_335,N_407);
nor U462 (N_462,N_366,N_360);
nor U463 (N_463,N_399,N_382);
and U464 (N_464,N_342,N_375);
and U465 (N_465,N_419,N_312);
or U466 (N_466,N_415,N_395);
nor U467 (N_467,N_386,N_381);
nor U468 (N_468,N_415,N_345);
or U469 (N_469,N_373,N_362);
nor U470 (N_470,N_394,N_345);
nor U471 (N_471,N_388,N_367);
and U472 (N_472,N_400,N_399);
or U473 (N_473,N_418,N_397);
and U474 (N_474,N_388,N_392);
nand U475 (N_475,N_416,N_392);
and U476 (N_476,N_412,N_376);
or U477 (N_477,N_365,N_294);
and U478 (N_478,N_360,N_194);
nor U479 (N_479,N_418,N_341);
nand U480 (N_480,N_459,N_421);
nor U481 (N_481,N_475,N_429);
nand U482 (N_482,N_445,N_449);
xor U483 (N_483,N_430,N_472);
nand U484 (N_484,N_440,N_447);
xor U485 (N_485,N_423,N_434);
nor U486 (N_486,N_425,N_476);
nor U487 (N_487,N_426,N_456);
and U488 (N_488,N_441,N_436);
nor U489 (N_489,N_461,N_442);
and U490 (N_490,N_428,N_448);
or U491 (N_491,N_432,N_455);
and U492 (N_492,N_463,N_451);
and U493 (N_493,N_435,N_439);
or U494 (N_494,N_479,N_444);
nor U495 (N_495,N_446,N_465);
nand U496 (N_496,N_470,N_452);
or U497 (N_497,N_471,N_468);
nor U498 (N_498,N_457,N_466);
and U499 (N_499,N_453,N_454);
and U500 (N_500,N_477,N_424);
and U501 (N_501,N_431,N_443);
and U502 (N_502,N_422,N_450);
or U503 (N_503,N_460,N_420);
and U504 (N_504,N_467,N_438);
nand U505 (N_505,N_474,N_464);
or U506 (N_506,N_437,N_458);
or U507 (N_507,N_473,N_427);
nor U508 (N_508,N_433,N_469);
or U509 (N_509,N_462,N_478);
and U510 (N_510,N_463,N_456);
or U511 (N_511,N_465,N_471);
nor U512 (N_512,N_433,N_451);
nor U513 (N_513,N_447,N_476);
and U514 (N_514,N_451,N_450);
or U515 (N_515,N_473,N_432);
nand U516 (N_516,N_429,N_450);
and U517 (N_517,N_427,N_425);
nor U518 (N_518,N_463,N_460);
and U519 (N_519,N_422,N_443);
and U520 (N_520,N_476,N_424);
and U521 (N_521,N_452,N_464);
and U522 (N_522,N_427,N_465);
xor U523 (N_523,N_474,N_440);
and U524 (N_524,N_426,N_469);
or U525 (N_525,N_470,N_463);
nor U526 (N_526,N_458,N_455);
and U527 (N_527,N_450,N_444);
or U528 (N_528,N_476,N_450);
nor U529 (N_529,N_425,N_445);
and U530 (N_530,N_475,N_427);
or U531 (N_531,N_463,N_447);
or U532 (N_532,N_475,N_462);
or U533 (N_533,N_454,N_422);
xor U534 (N_534,N_445,N_428);
or U535 (N_535,N_442,N_428);
nand U536 (N_536,N_451,N_421);
and U537 (N_537,N_460,N_425);
or U538 (N_538,N_454,N_433);
or U539 (N_539,N_445,N_436);
or U540 (N_540,N_538,N_517);
and U541 (N_541,N_484,N_481);
nand U542 (N_542,N_513,N_499);
or U543 (N_543,N_515,N_532);
xor U544 (N_544,N_535,N_500);
or U545 (N_545,N_492,N_523);
nor U546 (N_546,N_536,N_527);
or U547 (N_547,N_534,N_539);
and U548 (N_548,N_487,N_531);
and U549 (N_549,N_502,N_503);
nor U550 (N_550,N_508,N_489);
nor U551 (N_551,N_516,N_529);
and U552 (N_552,N_530,N_488);
and U553 (N_553,N_483,N_480);
nand U554 (N_554,N_522,N_506);
or U555 (N_555,N_509,N_505);
nor U556 (N_556,N_486,N_491);
and U557 (N_557,N_514,N_521);
nor U558 (N_558,N_510,N_525);
nor U559 (N_559,N_518,N_512);
or U560 (N_560,N_498,N_485);
and U561 (N_561,N_526,N_524);
or U562 (N_562,N_507,N_511);
nor U563 (N_563,N_520,N_497);
nor U564 (N_564,N_504,N_528);
and U565 (N_565,N_519,N_482);
or U566 (N_566,N_496,N_501);
nor U567 (N_567,N_493,N_494);
or U568 (N_568,N_537,N_490);
or U569 (N_569,N_533,N_495);
nor U570 (N_570,N_504,N_533);
and U571 (N_571,N_482,N_524);
nor U572 (N_572,N_492,N_499);
and U573 (N_573,N_486,N_493);
and U574 (N_574,N_480,N_538);
nor U575 (N_575,N_498,N_488);
nand U576 (N_576,N_515,N_485);
nand U577 (N_577,N_481,N_507);
or U578 (N_578,N_487,N_480);
nand U579 (N_579,N_536,N_493);
nor U580 (N_580,N_504,N_521);
nand U581 (N_581,N_486,N_531);
nand U582 (N_582,N_480,N_510);
nor U583 (N_583,N_523,N_518);
or U584 (N_584,N_533,N_515);
nand U585 (N_585,N_532,N_500);
xor U586 (N_586,N_535,N_491);
and U587 (N_587,N_538,N_495);
nor U588 (N_588,N_523,N_525);
xnor U589 (N_589,N_495,N_517);
nand U590 (N_590,N_500,N_533);
and U591 (N_591,N_515,N_495);
nand U592 (N_592,N_500,N_526);
or U593 (N_593,N_507,N_502);
and U594 (N_594,N_526,N_520);
nor U595 (N_595,N_499,N_493);
or U596 (N_596,N_527,N_493);
nand U597 (N_597,N_530,N_531);
or U598 (N_598,N_525,N_517);
nand U599 (N_599,N_509,N_506);
or U600 (N_600,N_562,N_546);
nand U601 (N_601,N_570,N_545);
or U602 (N_602,N_598,N_555);
nor U603 (N_603,N_599,N_594);
and U604 (N_604,N_577,N_588);
nand U605 (N_605,N_568,N_557);
nand U606 (N_606,N_586,N_561);
and U607 (N_607,N_548,N_558);
nor U608 (N_608,N_596,N_551);
nor U609 (N_609,N_597,N_550);
nand U610 (N_610,N_556,N_559);
nand U611 (N_611,N_541,N_563);
nor U612 (N_612,N_585,N_576);
or U613 (N_613,N_573,N_595);
and U614 (N_614,N_552,N_567);
and U615 (N_615,N_542,N_543);
nand U616 (N_616,N_554,N_590);
and U617 (N_617,N_565,N_582);
and U618 (N_618,N_540,N_560);
xnor U619 (N_619,N_547,N_583);
nor U620 (N_620,N_572,N_587);
and U621 (N_621,N_566,N_544);
and U622 (N_622,N_569,N_578);
nand U623 (N_623,N_592,N_593);
nand U624 (N_624,N_584,N_564);
xor U625 (N_625,N_575,N_580);
or U626 (N_626,N_581,N_589);
nor U627 (N_627,N_549,N_579);
and U628 (N_628,N_591,N_574);
or U629 (N_629,N_553,N_571);
nor U630 (N_630,N_567,N_574);
nand U631 (N_631,N_564,N_542);
nor U632 (N_632,N_577,N_592);
nor U633 (N_633,N_573,N_581);
and U634 (N_634,N_551,N_582);
or U635 (N_635,N_551,N_549);
and U636 (N_636,N_588,N_550);
and U637 (N_637,N_593,N_598);
nor U638 (N_638,N_568,N_553);
or U639 (N_639,N_540,N_595);
and U640 (N_640,N_555,N_543);
nor U641 (N_641,N_585,N_599);
nor U642 (N_642,N_583,N_540);
and U643 (N_643,N_549,N_568);
nor U644 (N_644,N_593,N_574);
nand U645 (N_645,N_566,N_583);
nor U646 (N_646,N_587,N_571);
and U647 (N_647,N_587,N_597);
nand U648 (N_648,N_559,N_551);
xor U649 (N_649,N_554,N_598);
or U650 (N_650,N_558,N_540);
nand U651 (N_651,N_584,N_599);
or U652 (N_652,N_577,N_549);
nor U653 (N_653,N_590,N_595);
nor U654 (N_654,N_550,N_586);
or U655 (N_655,N_584,N_553);
xor U656 (N_656,N_573,N_557);
nand U657 (N_657,N_551,N_547);
nand U658 (N_658,N_591,N_569);
or U659 (N_659,N_596,N_557);
or U660 (N_660,N_645,N_632);
nand U661 (N_661,N_629,N_639);
or U662 (N_662,N_649,N_659);
and U663 (N_663,N_643,N_623);
and U664 (N_664,N_630,N_653);
and U665 (N_665,N_641,N_658);
nand U666 (N_666,N_611,N_614);
or U667 (N_667,N_635,N_652);
and U668 (N_668,N_655,N_620);
or U669 (N_669,N_610,N_650);
nand U670 (N_670,N_637,N_624);
nand U671 (N_671,N_612,N_644);
or U672 (N_672,N_616,N_626);
nand U673 (N_673,N_651,N_647);
nor U674 (N_674,N_622,N_646);
nand U675 (N_675,N_615,N_654);
nor U676 (N_676,N_642,N_607);
or U677 (N_677,N_638,N_621);
and U678 (N_678,N_605,N_640);
and U679 (N_679,N_602,N_603);
and U680 (N_680,N_600,N_601);
and U681 (N_681,N_606,N_634);
nor U682 (N_682,N_656,N_618);
or U683 (N_683,N_604,N_628);
or U684 (N_684,N_609,N_627);
nand U685 (N_685,N_633,N_648);
or U686 (N_686,N_625,N_613);
or U687 (N_687,N_608,N_636);
nand U688 (N_688,N_657,N_617);
or U689 (N_689,N_631,N_619);
and U690 (N_690,N_636,N_639);
nand U691 (N_691,N_606,N_616);
nor U692 (N_692,N_628,N_641);
nor U693 (N_693,N_635,N_634);
and U694 (N_694,N_624,N_628);
nor U695 (N_695,N_648,N_629);
or U696 (N_696,N_608,N_602);
nand U697 (N_697,N_640,N_601);
or U698 (N_698,N_642,N_658);
nand U699 (N_699,N_641,N_618);
or U700 (N_700,N_641,N_647);
or U701 (N_701,N_642,N_619);
and U702 (N_702,N_645,N_627);
nand U703 (N_703,N_628,N_607);
nor U704 (N_704,N_646,N_610);
and U705 (N_705,N_656,N_600);
and U706 (N_706,N_602,N_632);
nand U707 (N_707,N_615,N_646);
or U708 (N_708,N_618,N_619);
or U709 (N_709,N_628,N_610);
nand U710 (N_710,N_607,N_639);
nor U711 (N_711,N_617,N_658);
or U712 (N_712,N_621,N_606);
nor U713 (N_713,N_618,N_640);
nand U714 (N_714,N_606,N_633);
and U715 (N_715,N_605,N_607);
nor U716 (N_716,N_608,N_657);
or U717 (N_717,N_616,N_623);
nor U718 (N_718,N_620,N_634);
or U719 (N_719,N_646,N_626);
nand U720 (N_720,N_694,N_687);
nand U721 (N_721,N_691,N_705);
nor U722 (N_722,N_675,N_670);
or U723 (N_723,N_692,N_676);
nor U724 (N_724,N_707,N_700);
nand U725 (N_725,N_703,N_671);
nor U726 (N_726,N_663,N_662);
or U727 (N_727,N_689,N_688);
or U728 (N_728,N_690,N_717);
xnor U729 (N_729,N_677,N_699);
or U730 (N_730,N_710,N_665);
nand U731 (N_731,N_660,N_706);
and U732 (N_732,N_704,N_719);
and U733 (N_733,N_709,N_715);
or U734 (N_734,N_674,N_693);
nor U735 (N_735,N_695,N_683);
nor U736 (N_736,N_667,N_685);
nand U737 (N_737,N_711,N_714);
or U738 (N_738,N_681,N_672);
nor U739 (N_739,N_686,N_678);
xnor U740 (N_740,N_716,N_679);
and U741 (N_741,N_702,N_680);
and U742 (N_742,N_661,N_713);
nand U743 (N_743,N_697,N_664);
nand U744 (N_744,N_708,N_696);
nand U745 (N_745,N_666,N_684);
nor U746 (N_746,N_698,N_701);
or U747 (N_747,N_669,N_668);
and U748 (N_748,N_712,N_673);
nand U749 (N_749,N_718,N_682);
xnor U750 (N_750,N_702,N_699);
or U751 (N_751,N_674,N_687);
nand U752 (N_752,N_719,N_692);
and U753 (N_753,N_717,N_661);
or U754 (N_754,N_664,N_702);
nand U755 (N_755,N_716,N_707);
and U756 (N_756,N_678,N_696);
nor U757 (N_757,N_696,N_709);
nand U758 (N_758,N_716,N_697);
nand U759 (N_759,N_713,N_719);
or U760 (N_760,N_700,N_666);
nor U761 (N_761,N_707,N_706);
nor U762 (N_762,N_685,N_677);
nor U763 (N_763,N_694,N_664);
nor U764 (N_764,N_707,N_674);
and U765 (N_765,N_715,N_687);
and U766 (N_766,N_690,N_667);
nor U767 (N_767,N_673,N_668);
and U768 (N_768,N_679,N_667);
or U769 (N_769,N_698,N_682);
xor U770 (N_770,N_702,N_670);
nor U771 (N_771,N_661,N_672);
nor U772 (N_772,N_700,N_668);
nor U773 (N_773,N_693,N_695);
nand U774 (N_774,N_684,N_677);
nand U775 (N_775,N_711,N_683);
xnor U776 (N_776,N_685,N_717);
nand U777 (N_777,N_672,N_671);
or U778 (N_778,N_714,N_718);
and U779 (N_779,N_664,N_687);
nand U780 (N_780,N_722,N_772);
or U781 (N_781,N_733,N_751);
nor U782 (N_782,N_746,N_773);
nor U783 (N_783,N_726,N_743);
and U784 (N_784,N_754,N_775);
nor U785 (N_785,N_724,N_757);
nand U786 (N_786,N_756,N_738);
and U787 (N_787,N_759,N_727);
nor U788 (N_788,N_763,N_778);
nand U789 (N_789,N_758,N_760);
nand U790 (N_790,N_777,N_734);
nor U791 (N_791,N_741,N_765);
and U792 (N_792,N_767,N_770);
nand U793 (N_793,N_766,N_761);
nor U794 (N_794,N_748,N_725);
nand U795 (N_795,N_768,N_747);
nor U796 (N_796,N_771,N_735);
nand U797 (N_797,N_728,N_721);
nor U798 (N_798,N_769,N_753);
nor U799 (N_799,N_774,N_745);
nand U800 (N_800,N_737,N_752);
nand U801 (N_801,N_776,N_729);
and U802 (N_802,N_720,N_764);
or U803 (N_803,N_755,N_744);
and U804 (N_804,N_736,N_731);
nor U805 (N_805,N_732,N_742);
or U806 (N_806,N_750,N_749);
nand U807 (N_807,N_739,N_723);
nand U808 (N_808,N_730,N_762);
or U809 (N_809,N_779,N_740);
nand U810 (N_810,N_724,N_771);
or U811 (N_811,N_728,N_776);
xor U812 (N_812,N_743,N_763);
nor U813 (N_813,N_726,N_770);
and U814 (N_814,N_730,N_726);
or U815 (N_815,N_756,N_779);
or U816 (N_816,N_762,N_723);
nand U817 (N_817,N_761,N_736);
nor U818 (N_818,N_772,N_770);
nor U819 (N_819,N_745,N_746);
nor U820 (N_820,N_721,N_762);
nand U821 (N_821,N_744,N_726);
nor U822 (N_822,N_765,N_729);
and U823 (N_823,N_772,N_731);
or U824 (N_824,N_735,N_736);
and U825 (N_825,N_764,N_775);
or U826 (N_826,N_732,N_722);
or U827 (N_827,N_730,N_725);
nor U828 (N_828,N_779,N_722);
nor U829 (N_829,N_777,N_753);
nor U830 (N_830,N_761,N_752);
or U831 (N_831,N_741,N_758);
and U832 (N_832,N_761,N_760);
and U833 (N_833,N_751,N_767);
nor U834 (N_834,N_736,N_741);
and U835 (N_835,N_777,N_771);
and U836 (N_836,N_722,N_756);
nor U837 (N_837,N_729,N_773);
nor U838 (N_838,N_762,N_769);
or U839 (N_839,N_779,N_727);
xor U840 (N_840,N_839,N_797);
xnor U841 (N_841,N_837,N_803);
nor U842 (N_842,N_782,N_786);
and U843 (N_843,N_823,N_807);
or U844 (N_844,N_793,N_806);
and U845 (N_845,N_802,N_812);
and U846 (N_846,N_791,N_792);
nor U847 (N_847,N_789,N_781);
nor U848 (N_848,N_796,N_799);
nor U849 (N_849,N_787,N_831);
nor U850 (N_850,N_809,N_800);
xnor U851 (N_851,N_832,N_813);
and U852 (N_852,N_827,N_785);
nand U853 (N_853,N_830,N_833);
nand U854 (N_854,N_816,N_795);
nor U855 (N_855,N_822,N_801);
and U856 (N_856,N_819,N_814);
nand U857 (N_857,N_815,N_838);
and U858 (N_858,N_828,N_824);
or U859 (N_859,N_825,N_834);
nand U860 (N_860,N_804,N_817);
and U861 (N_861,N_836,N_798);
nor U862 (N_862,N_820,N_783);
or U863 (N_863,N_810,N_818);
nand U864 (N_864,N_808,N_826);
and U865 (N_865,N_780,N_794);
nand U866 (N_866,N_821,N_829);
nor U867 (N_867,N_811,N_788);
and U868 (N_868,N_790,N_835);
nand U869 (N_869,N_784,N_805);
or U870 (N_870,N_809,N_785);
or U871 (N_871,N_829,N_824);
nand U872 (N_872,N_802,N_821);
nor U873 (N_873,N_820,N_804);
nor U874 (N_874,N_794,N_802);
or U875 (N_875,N_838,N_832);
nor U876 (N_876,N_826,N_806);
nor U877 (N_877,N_822,N_799);
or U878 (N_878,N_814,N_787);
nand U879 (N_879,N_824,N_833);
nor U880 (N_880,N_838,N_795);
or U881 (N_881,N_835,N_811);
nor U882 (N_882,N_788,N_803);
nand U883 (N_883,N_786,N_826);
and U884 (N_884,N_813,N_805);
nand U885 (N_885,N_791,N_828);
and U886 (N_886,N_805,N_786);
and U887 (N_887,N_801,N_813);
or U888 (N_888,N_792,N_806);
nor U889 (N_889,N_780,N_812);
nor U890 (N_890,N_816,N_794);
or U891 (N_891,N_781,N_782);
nor U892 (N_892,N_814,N_826);
nand U893 (N_893,N_829,N_813);
nand U894 (N_894,N_786,N_781);
nand U895 (N_895,N_786,N_811);
nor U896 (N_896,N_810,N_837);
nand U897 (N_897,N_834,N_827);
nand U898 (N_898,N_828,N_832);
xnor U899 (N_899,N_826,N_782);
and U900 (N_900,N_879,N_863);
or U901 (N_901,N_877,N_840);
nor U902 (N_902,N_896,N_853);
or U903 (N_903,N_844,N_852);
or U904 (N_904,N_846,N_842);
and U905 (N_905,N_870,N_892);
nand U906 (N_906,N_878,N_889);
or U907 (N_907,N_859,N_843);
and U908 (N_908,N_880,N_874);
nand U909 (N_909,N_895,N_887);
or U910 (N_910,N_862,N_890);
nand U911 (N_911,N_869,N_849);
nand U912 (N_912,N_858,N_851);
and U913 (N_913,N_871,N_876);
nand U914 (N_914,N_847,N_884);
nor U915 (N_915,N_891,N_854);
and U916 (N_916,N_881,N_897);
or U917 (N_917,N_872,N_865);
nor U918 (N_918,N_885,N_886);
nand U919 (N_919,N_894,N_845);
nor U920 (N_920,N_860,N_898);
and U921 (N_921,N_861,N_899);
and U922 (N_922,N_841,N_850);
or U923 (N_923,N_855,N_888);
and U924 (N_924,N_868,N_848);
nor U925 (N_925,N_866,N_883);
and U926 (N_926,N_864,N_857);
nand U927 (N_927,N_856,N_873);
and U928 (N_928,N_882,N_875);
or U929 (N_929,N_893,N_867);
nand U930 (N_930,N_869,N_863);
and U931 (N_931,N_851,N_856);
and U932 (N_932,N_874,N_856);
nand U933 (N_933,N_887,N_871);
and U934 (N_934,N_848,N_889);
nor U935 (N_935,N_897,N_857);
and U936 (N_936,N_876,N_884);
and U937 (N_937,N_877,N_857);
nand U938 (N_938,N_841,N_865);
or U939 (N_939,N_851,N_874);
nor U940 (N_940,N_872,N_851);
nand U941 (N_941,N_896,N_844);
nor U942 (N_942,N_887,N_881);
or U943 (N_943,N_871,N_892);
nand U944 (N_944,N_840,N_868);
nand U945 (N_945,N_875,N_887);
nor U946 (N_946,N_870,N_856);
and U947 (N_947,N_866,N_875);
and U948 (N_948,N_895,N_890);
nor U949 (N_949,N_849,N_863);
nor U950 (N_950,N_881,N_885);
nor U951 (N_951,N_845,N_890);
nor U952 (N_952,N_858,N_862);
and U953 (N_953,N_890,N_876);
nor U954 (N_954,N_887,N_858);
or U955 (N_955,N_863,N_861);
and U956 (N_956,N_873,N_850);
nor U957 (N_957,N_844,N_867);
and U958 (N_958,N_882,N_843);
or U959 (N_959,N_854,N_870);
nand U960 (N_960,N_900,N_934);
nand U961 (N_961,N_912,N_906);
or U962 (N_962,N_949,N_908);
or U963 (N_963,N_946,N_956);
and U964 (N_964,N_951,N_914);
or U965 (N_965,N_920,N_936);
nor U966 (N_966,N_941,N_939);
nor U967 (N_967,N_937,N_957);
or U968 (N_968,N_919,N_953);
nand U969 (N_969,N_929,N_942);
nand U970 (N_970,N_940,N_950);
or U971 (N_971,N_911,N_927);
or U972 (N_972,N_917,N_947);
nand U973 (N_973,N_907,N_915);
nand U974 (N_974,N_925,N_916);
nand U975 (N_975,N_935,N_933);
nor U976 (N_976,N_938,N_943);
and U977 (N_977,N_902,N_905);
or U978 (N_978,N_903,N_954);
and U979 (N_979,N_922,N_928);
nor U980 (N_980,N_924,N_958);
or U981 (N_981,N_948,N_904);
nand U982 (N_982,N_921,N_931);
nand U983 (N_983,N_923,N_909);
and U984 (N_984,N_913,N_910);
or U985 (N_985,N_955,N_945);
nor U986 (N_986,N_926,N_959);
nand U987 (N_987,N_930,N_944);
and U988 (N_988,N_952,N_932);
or U989 (N_989,N_901,N_918);
nor U990 (N_990,N_941,N_919);
nand U991 (N_991,N_933,N_941);
nor U992 (N_992,N_916,N_946);
and U993 (N_993,N_940,N_955);
nand U994 (N_994,N_931,N_915);
and U995 (N_995,N_906,N_957);
nor U996 (N_996,N_957,N_901);
nor U997 (N_997,N_910,N_934);
or U998 (N_998,N_934,N_919);
or U999 (N_999,N_903,N_919);
or U1000 (N_1000,N_929,N_947);
nor U1001 (N_1001,N_957,N_947);
or U1002 (N_1002,N_958,N_937);
or U1003 (N_1003,N_931,N_923);
and U1004 (N_1004,N_944,N_941);
or U1005 (N_1005,N_939,N_936);
nand U1006 (N_1006,N_907,N_946);
nand U1007 (N_1007,N_910,N_908);
and U1008 (N_1008,N_905,N_929);
nor U1009 (N_1009,N_915,N_910);
or U1010 (N_1010,N_931,N_926);
nand U1011 (N_1011,N_952,N_950);
or U1012 (N_1012,N_926,N_932);
nor U1013 (N_1013,N_920,N_956);
nand U1014 (N_1014,N_903,N_907);
nand U1015 (N_1015,N_949,N_917);
nand U1016 (N_1016,N_936,N_906);
or U1017 (N_1017,N_906,N_945);
nor U1018 (N_1018,N_921,N_946);
nand U1019 (N_1019,N_918,N_930);
nor U1020 (N_1020,N_985,N_1018);
nand U1021 (N_1021,N_980,N_978);
and U1022 (N_1022,N_992,N_964);
and U1023 (N_1023,N_1005,N_1002);
nor U1024 (N_1024,N_997,N_1003);
xor U1025 (N_1025,N_962,N_984);
or U1026 (N_1026,N_1016,N_988);
or U1027 (N_1027,N_968,N_1014);
nand U1028 (N_1028,N_983,N_999);
and U1029 (N_1029,N_972,N_979);
xnor U1030 (N_1030,N_975,N_1000);
nand U1031 (N_1031,N_987,N_974);
or U1032 (N_1032,N_1019,N_1007);
xor U1033 (N_1033,N_982,N_976);
nor U1034 (N_1034,N_996,N_995);
nor U1035 (N_1035,N_986,N_981);
or U1036 (N_1036,N_990,N_960);
nand U1037 (N_1037,N_969,N_977);
nor U1038 (N_1038,N_1012,N_1009);
or U1039 (N_1039,N_1001,N_965);
or U1040 (N_1040,N_1017,N_1015);
or U1041 (N_1041,N_971,N_1004);
nor U1042 (N_1042,N_991,N_967);
and U1043 (N_1043,N_1011,N_966);
or U1044 (N_1044,N_993,N_1013);
nand U1045 (N_1045,N_970,N_998);
or U1046 (N_1046,N_1006,N_961);
nand U1047 (N_1047,N_1008,N_989);
and U1048 (N_1048,N_963,N_994);
and U1049 (N_1049,N_973,N_1010);
nor U1050 (N_1050,N_972,N_967);
or U1051 (N_1051,N_983,N_976);
nand U1052 (N_1052,N_978,N_965);
nand U1053 (N_1053,N_967,N_997);
or U1054 (N_1054,N_1014,N_963);
and U1055 (N_1055,N_971,N_1012);
and U1056 (N_1056,N_1005,N_1018);
nand U1057 (N_1057,N_1016,N_963);
or U1058 (N_1058,N_1012,N_991);
nand U1059 (N_1059,N_1005,N_993);
nor U1060 (N_1060,N_975,N_965);
nor U1061 (N_1061,N_1007,N_997);
or U1062 (N_1062,N_982,N_992);
and U1063 (N_1063,N_1007,N_985);
or U1064 (N_1064,N_998,N_1012);
nand U1065 (N_1065,N_970,N_972);
nand U1066 (N_1066,N_995,N_968);
and U1067 (N_1067,N_981,N_973);
and U1068 (N_1068,N_1010,N_1002);
or U1069 (N_1069,N_1012,N_1014);
nand U1070 (N_1070,N_978,N_1013);
nand U1071 (N_1071,N_1006,N_977);
or U1072 (N_1072,N_1016,N_997);
and U1073 (N_1073,N_976,N_974);
nor U1074 (N_1074,N_1001,N_984);
nand U1075 (N_1075,N_964,N_967);
xnor U1076 (N_1076,N_992,N_1001);
nor U1077 (N_1077,N_1000,N_995);
nand U1078 (N_1078,N_967,N_966);
nor U1079 (N_1079,N_1005,N_1013);
nor U1080 (N_1080,N_1054,N_1062);
and U1081 (N_1081,N_1047,N_1027);
and U1082 (N_1082,N_1032,N_1071);
nand U1083 (N_1083,N_1045,N_1041);
and U1084 (N_1084,N_1053,N_1070);
nor U1085 (N_1085,N_1042,N_1046);
or U1086 (N_1086,N_1060,N_1037);
nor U1087 (N_1087,N_1051,N_1056);
nor U1088 (N_1088,N_1079,N_1058);
or U1089 (N_1089,N_1030,N_1055);
nand U1090 (N_1090,N_1065,N_1044);
nor U1091 (N_1091,N_1064,N_1021);
xnor U1092 (N_1092,N_1052,N_1076);
nor U1093 (N_1093,N_1033,N_1039);
nand U1094 (N_1094,N_1073,N_1077);
nand U1095 (N_1095,N_1049,N_1059);
and U1096 (N_1096,N_1067,N_1040);
or U1097 (N_1097,N_1028,N_1038);
and U1098 (N_1098,N_1069,N_1043);
or U1099 (N_1099,N_1057,N_1029);
nand U1100 (N_1100,N_1034,N_1036);
nand U1101 (N_1101,N_1068,N_1072);
nand U1102 (N_1102,N_1061,N_1031);
and U1103 (N_1103,N_1048,N_1023);
nor U1104 (N_1104,N_1026,N_1075);
nand U1105 (N_1105,N_1066,N_1078);
and U1106 (N_1106,N_1050,N_1074);
nor U1107 (N_1107,N_1063,N_1035);
nor U1108 (N_1108,N_1025,N_1020);
or U1109 (N_1109,N_1024,N_1022);
or U1110 (N_1110,N_1038,N_1061);
and U1111 (N_1111,N_1044,N_1046);
nor U1112 (N_1112,N_1061,N_1055);
and U1113 (N_1113,N_1027,N_1078);
nand U1114 (N_1114,N_1077,N_1046);
nand U1115 (N_1115,N_1048,N_1053);
nand U1116 (N_1116,N_1031,N_1034);
or U1117 (N_1117,N_1056,N_1048);
nor U1118 (N_1118,N_1066,N_1073);
nor U1119 (N_1119,N_1024,N_1062);
or U1120 (N_1120,N_1025,N_1059);
nand U1121 (N_1121,N_1063,N_1073);
nor U1122 (N_1122,N_1031,N_1044);
or U1123 (N_1123,N_1067,N_1030);
nor U1124 (N_1124,N_1022,N_1026);
and U1125 (N_1125,N_1042,N_1039);
nand U1126 (N_1126,N_1022,N_1040);
and U1127 (N_1127,N_1063,N_1061);
and U1128 (N_1128,N_1056,N_1020);
and U1129 (N_1129,N_1038,N_1078);
or U1130 (N_1130,N_1078,N_1065);
and U1131 (N_1131,N_1067,N_1023);
nor U1132 (N_1132,N_1063,N_1054);
nand U1133 (N_1133,N_1035,N_1046);
and U1134 (N_1134,N_1063,N_1048);
and U1135 (N_1135,N_1046,N_1073);
or U1136 (N_1136,N_1046,N_1020);
nor U1137 (N_1137,N_1067,N_1052);
nand U1138 (N_1138,N_1031,N_1048);
and U1139 (N_1139,N_1074,N_1055);
nand U1140 (N_1140,N_1101,N_1112);
and U1141 (N_1141,N_1105,N_1116);
nand U1142 (N_1142,N_1108,N_1134);
or U1143 (N_1143,N_1110,N_1137);
and U1144 (N_1144,N_1089,N_1125);
xnor U1145 (N_1145,N_1139,N_1133);
nand U1146 (N_1146,N_1081,N_1097);
or U1147 (N_1147,N_1102,N_1121);
nor U1148 (N_1148,N_1138,N_1080);
nor U1149 (N_1149,N_1100,N_1087);
and U1150 (N_1150,N_1088,N_1083);
or U1151 (N_1151,N_1092,N_1130);
nand U1152 (N_1152,N_1094,N_1095);
and U1153 (N_1153,N_1104,N_1086);
nor U1154 (N_1154,N_1096,N_1126);
nor U1155 (N_1155,N_1132,N_1113);
nand U1156 (N_1156,N_1118,N_1091);
or U1157 (N_1157,N_1128,N_1090);
or U1158 (N_1158,N_1119,N_1124);
or U1159 (N_1159,N_1123,N_1114);
nor U1160 (N_1160,N_1103,N_1115);
nand U1161 (N_1161,N_1085,N_1127);
and U1162 (N_1162,N_1120,N_1099);
or U1163 (N_1163,N_1109,N_1136);
or U1164 (N_1164,N_1098,N_1082);
xnor U1165 (N_1165,N_1129,N_1107);
nor U1166 (N_1166,N_1106,N_1111);
and U1167 (N_1167,N_1135,N_1084);
nor U1168 (N_1168,N_1117,N_1122);
and U1169 (N_1169,N_1131,N_1093);
nor U1170 (N_1170,N_1117,N_1098);
nand U1171 (N_1171,N_1102,N_1111);
nor U1172 (N_1172,N_1107,N_1122);
and U1173 (N_1173,N_1090,N_1088);
nand U1174 (N_1174,N_1096,N_1105);
and U1175 (N_1175,N_1119,N_1105);
nor U1176 (N_1176,N_1117,N_1091);
and U1177 (N_1177,N_1081,N_1091);
or U1178 (N_1178,N_1081,N_1139);
nor U1179 (N_1179,N_1090,N_1121);
nand U1180 (N_1180,N_1098,N_1122);
nor U1181 (N_1181,N_1111,N_1104);
nand U1182 (N_1182,N_1133,N_1116);
and U1183 (N_1183,N_1129,N_1121);
nand U1184 (N_1184,N_1124,N_1086);
nand U1185 (N_1185,N_1136,N_1094);
nor U1186 (N_1186,N_1083,N_1123);
nand U1187 (N_1187,N_1102,N_1123);
nand U1188 (N_1188,N_1134,N_1128);
and U1189 (N_1189,N_1085,N_1105);
or U1190 (N_1190,N_1109,N_1132);
or U1191 (N_1191,N_1135,N_1115);
nor U1192 (N_1192,N_1098,N_1083);
and U1193 (N_1193,N_1130,N_1105);
nor U1194 (N_1194,N_1098,N_1106);
nand U1195 (N_1195,N_1115,N_1134);
or U1196 (N_1196,N_1098,N_1114);
nor U1197 (N_1197,N_1085,N_1134);
or U1198 (N_1198,N_1083,N_1139);
nand U1199 (N_1199,N_1086,N_1105);
or U1200 (N_1200,N_1199,N_1182);
nand U1201 (N_1201,N_1171,N_1178);
nand U1202 (N_1202,N_1168,N_1189);
nand U1203 (N_1203,N_1164,N_1157);
nand U1204 (N_1204,N_1154,N_1158);
nand U1205 (N_1205,N_1167,N_1192);
nand U1206 (N_1206,N_1147,N_1191);
nand U1207 (N_1207,N_1196,N_1141);
nor U1208 (N_1208,N_1180,N_1179);
and U1209 (N_1209,N_1152,N_1159);
nor U1210 (N_1210,N_1184,N_1181);
or U1211 (N_1211,N_1197,N_1150);
nand U1212 (N_1212,N_1169,N_1142);
or U1213 (N_1213,N_1153,N_1175);
and U1214 (N_1214,N_1170,N_1151);
nand U1215 (N_1215,N_1155,N_1174);
and U1216 (N_1216,N_1148,N_1186);
nor U1217 (N_1217,N_1160,N_1156);
nand U1218 (N_1218,N_1188,N_1177);
nand U1219 (N_1219,N_1166,N_1140);
nand U1220 (N_1220,N_1149,N_1146);
nor U1221 (N_1221,N_1172,N_1195);
xnor U1222 (N_1222,N_1161,N_1187);
nor U1223 (N_1223,N_1162,N_1176);
or U1224 (N_1224,N_1145,N_1173);
xor U1225 (N_1225,N_1183,N_1194);
nand U1226 (N_1226,N_1165,N_1163);
or U1227 (N_1227,N_1193,N_1190);
xnor U1228 (N_1228,N_1143,N_1144);
or U1229 (N_1229,N_1198,N_1185);
nand U1230 (N_1230,N_1165,N_1190);
or U1231 (N_1231,N_1181,N_1176);
nor U1232 (N_1232,N_1191,N_1184);
nor U1233 (N_1233,N_1190,N_1194);
nand U1234 (N_1234,N_1150,N_1189);
or U1235 (N_1235,N_1149,N_1186);
nor U1236 (N_1236,N_1186,N_1155);
nand U1237 (N_1237,N_1155,N_1187);
nand U1238 (N_1238,N_1149,N_1167);
nand U1239 (N_1239,N_1182,N_1179);
and U1240 (N_1240,N_1160,N_1185);
and U1241 (N_1241,N_1148,N_1193);
or U1242 (N_1242,N_1180,N_1140);
or U1243 (N_1243,N_1172,N_1156);
nand U1244 (N_1244,N_1183,N_1162);
or U1245 (N_1245,N_1180,N_1152);
and U1246 (N_1246,N_1164,N_1151);
nor U1247 (N_1247,N_1177,N_1186);
and U1248 (N_1248,N_1154,N_1179);
and U1249 (N_1249,N_1160,N_1179);
and U1250 (N_1250,N_1195,N_1160);
nand U1251 (N_1251,N_1163,N_1149);
and U1252 (N_1252,N_1172,N_1189);
nor U1253 (N_1253,N_1154,N_1143);
nor U1254 (N_1254,N_1179,N_1143);
and U1255 (N_1255,N_1165,N_1182);
and U1256 (N_1256,N_1158,N_1196);
and U1257 (N_1257,N_1148,N_1171);
nand U1258 (N_1258,N_1156,N_1142);
or U1259 (N_1259,N_1179,N_1147);
nand U1260 (N_1260,N_1256,N_1220);
and U1261 (N_1261,N_1252,N_1254);
nand U1262 (N_1262,N_1222,N_1249);
and U1263 (N_1263,N_1217,N_1242);
or U1264 (N_1264,N_1251,N_1235);
and U1265 (N_1265,N_1224,N_1246);
and U1266 (N_1266,N_1223,N_1215);
and U1267 (N_1267,N_1237,N_1211);
and U1268 (N_1268,N_1230,N_1212);
or U1269 (N_1269,N_1258,N_1241);
or U1270 (N_1270,N_1203,N_1213);
nand U1271 (N_1271,N_1208,N_1236);
nand U1272 (N_1272,N_1201,N_1234);
nor U1273 (N_1273,N_1233,N_1225);
or U1274 (N_1274,N_1219,N_1243);
or U1275 (N_1275,N_1240,N_1207);
and U1276 (N_1276,N_1221,N_1204);
nand U1277 (N_1277,N_1239,N_1244);
nand U1278 (N_1278,N_1206,N_1210);
nor U1279 (N_1279,N_1255,N_1248);
and U1280 (N_1280,N_1209,N_1231);
and U1281 (N_1281,N_1202,N_1228);
nor U1282 (N_1282,N_1218,N_1205);
nand U1283 (N_1283,N_1229,N_1253);
nand U1284 (N_1284,N_1245,N_1216);
nand U1285 (N_1285,N_1257,N_1250);
and U1286 (N_1286,N_1238,N_1214);
or U1287 (N_1287,N_1259,N_1227);
or U1288 (N_1288,N_1232,N_1247);
nor U1289 (N_1289,N_1226,N_1200);
or U1290 (N_1290,N_1231,N_1259);
nand U1291 (N_1291,N_1217,N_1251);
and U1292 (N_1292,N_1252,N_1221);
nand U1293 (N_1293,N_1203,N_1216);
nand U1294 (N_1294,N_1216,N_1258);
nor U1295 (N_1295,N_1237,N_1238);
nor U1296 (N_1296,N_1230,N_1225);
nand U1297 (N_1297,N_1257,N_1214);
or U1298 (N_1298,N_1238,N_1203);
and U1299 (N_1299,N_1259,N_1229);
and U1300 (N_1300,N_1207,N_1220);
nand U1301 (N_1301,N_1249,N_1217);
nor U1302 (N_1302,N_1228,N_1230);
and U1303 (N_1303,N_1200,N_1229);
xor U1304 (N_1304,N_1215,N_1210);
nand U1305 (N_1305,N_1221,N_1215);
xor U1306 (N_1306,N_1241,N_1236);
nand U1307 (N_1307,N_1257,N_1236);
or U1308 (N_1308,N_1234,N_1213);
nand U1309 (N_1309,N_1211,N_1228);
nand U1310 (N_1310,N_1214,N_1253);
nand U1311 (N_1311,N_1243,N_1221);
nor U1312 (N_1312,N_1218,N_1248);
nor U1313 (N_1313,N_1256,N_1229);
nor U1314 (N_1314,N_1234,N_1224);
nor U1315 (N_1315,N_1259,N_1233);
or U1316 (N_1316,N_1252,N_1205);
and U1317 (N_1317,N_1237,N_1207);
or U1318 (N_1318,N_1220,N_1241);
and U1319 (N_1319,N_1204,N_1249);
nor U1320 (N_1320,N_1269,N_1302);
and U1321 (N_1321,N_1291,N_1285);
nand U1322 (N_1322,N_1309,N_1298);
and U1323 (N_1323,N_1292,N_1293);
nor U1324 (N_1324,N_1281,N_1290);
nor U1325 (N_1325,N_1300,N_1314);
and U1326 (N_1326,N_1267,N_1299);
and U1327 (N_1327,N_1264,N_1270);
nor U1328 (N_1328,N_1276,N_1271);
nand U1329 (N_1329,N_1310,N_1260);
and U1330 (N_1330,N_1295,N_1273);
or U1331 (N_1331,N_1275,N_1318);
or U1332 (N_1332,N_1315,N_1301);
or U1333 (N_1333,N_1265,N_1274);
nand U1334 (N_1334,N_1303,N_1283);
and U1335 (N_1335,N_1278,N_1294);
and U1336 (N_1336,N_1263,N_1305);
or U1337 (N_1337,N_1289,N_1287);
nor U1338 (N_1338,N_1286,N_1266);
or U1339 (N_1339,N_1280,N_1262);
or U1340 (N_1340,N_1317,N_1272);
and U1341 (N_1341,N_1311,N_1279);
and U1342 (N_1342,N_1304,N_1288);
nand U1343 (N_1343,N_1306,N_1282);
nand U1344 (N_1344,N_1277,N_1284);
nor U1345 (N_1345,N_1319,N_1261);
or U1346 (N_1346,N_1316,N_1307);
nor U1347 (N_1347,N_1313,N_1268);
nor U1348 (N_1348,N_1308,N_1312);
nand U1349 (N_1349,N_1297,N_1296);
and U1350 (N_1350,N_1311,N_1262);
nor U1351 (N_1351,N_1263,N_1302);
and U1352 (N_1352,N_1305,N_1271);
nand U1353 (N_1353,N_1271,N_1273);
or U1354 (N_1354,N_1295,N_1308);
nor U1355 (N_1355,N_1313,N_1314);
nor U1356 (N_1356,N_1305,N_1296);
nor U1357 (N_1357,N_1291,N_1269);
nand U1358 (N_1358,N_1294,N_1279);
nand U1359 (N_1359,N_1319,N_1291);
and U1360 (N_1360,N_1277,N_1261);
nand U1361 (N_1361,N_1296,N_1282);
nor U1362 (N_1362,N_1299,N_1318);
and U1363 (N_1363,N_1260,N_1271);
nor U1364 (N_1364,N_1293,N_1308);
or U1365 (N_1365,N_1309,N_1283);
or U1366 (N_1366,N_1281,N_1288);
and U1367 (N_1367,N_1302,N_1292);
or U1368 (N_1368,N_1275,N_1298);
and U1369 (N_1369,N_1286,N_1296);
or U1370 (N_1370,N_1260,N_1279);
nand U1371 (N_1371,N_1295,N_1312);
and U1372 (N_1372,N_1317,N_1290);
or U1373 (N_1373,N_1261,N_1286);
or U1374 (N_1374,N_1280,N_1298);
and U1375 (N_1375,N_1279,N_1284);
or U1376 (N_1376,N_1317,N_1274);
nor U1377 (N_1377,N_1279,N_1288);
and U1378 (N_1378,N_1310,N_1317);
or U1379 (N_1379,N_1274,N_1302);
nor U1380 (N_1380,N_1358,N_1336);
nor U1381 (N_1381,N_1372,N_1350);
and U1382 (N_1382,N_1327,N_1338);
nand U1383 (N_1383,N_1339,N_1321);
and U1384 (N_1384,N_1366,N_1377);
nor U1385 (N_1385,N_1328,N_1357);
nand U1386 (N_1386,N_1378,N_1342);
and U1387 (N_1387,N_1326,N_1363);
nand U1388 (N_1388,N_1364,N_1330);
or U1389 (N_1389,N_1352,N_1351);
nor U1390 (N_1390,N_1376,N_1322);
and U1391 (N_1391,N_1343,N_1331);
and U1392 (N_1392,N_1346,N_1365);
nand U1393 (N_1393,N_1345,N_1347);
nor U1394 (N_1394,N_1349,N_1341);
or U1395 (N_1395,N_1375,N_1340);
or U1396 (N_1396,N_1369,N_1334);
or U1397 (N_1397,N_1329,N_1325);
nand U1398 (N_1398,N_1362,N_1359);
and U1399 (N_1399,N_1354,N_1335);
nor U1400 (N_1400,N_1379,N_1323);
nand U1401 (N_1401,N_1324,N_1367);
xnor U1402 (N_1402,N_1361,N_1337);
or U1403 (N_1403,N_1344,N_1333);
nor U1404 (N_1404,N_1356,N_1355);
nand U1405 (N_1405,N_1320,N_1332);
and U1406 (N_1406,N_1371,N_1368);
and U1407 (N_1407,N_1374,N_1360);
and U1408 (N_1408,N_1353,N_1348);
nor U1409 (N_1409,N_1370,N_1373);
nand U1410 (N_1410,N_1356,N_1358);
and U1411 (N_1411,N_1364,N_1336);
nand U1412 (N_1412,N_1377,N_1368);
nand U1413 (N_1413,N_1354,N_1358);
nor U1414 (N_1414,N_1356,N_1345);
nor U1415 (N_1415,N_1365,N_1359);
or U1416 (N_1416,N_1372,N_1351);
nand U1417 (N_1417,N_1327,N_1356);
and U1418 (N_1418,N_1364,N_1361);
or U1419 (N_1419,N_1369,N_1333);
and U1420 (N_1420,N_1369,N_1371);
nand U1421 (N_1421,N_1359,N_1350);
or U1422 (N_1422,N_1357,N_1340);
nand U1423 (N_1423,N_1369,N_1329);
nand U1424 (N_1424,N_1339,N_1332);
and U1425 (N_1425,N_1344,N_1334);
nand U1426 (N_1426,N_1347,N_1367);
and U1427 (N_1427,N_1323,N_1359);
nor U1428 (N_1428,N_1367,N_1374);
and U1429 (N_1429,N_1337,N_1360);
nor U1430 (N_1430,N_1353,N_1328);
or U1431 (N_1431,N_1339,N_1335);
nor U1432 (N_1432,N_1375,N_1332);
nor U1433 (N_1433,N_1336,N_1368);
nand U1434 (N_1434,N_1374,N_1364);
nand U1435 (N_1435,N_1368,N_1326);
or U1436 (N_1436,N_1368,N_1334);
xnor U1437 (N_1437,N_1375,N_1372);
and U1438 (N_1438,N_1331,N_1368);
nand U1439 (N_1439,N_1346,N_1350);
and U1440 (N_1440,N_1417,N_1415);
nor U1441 (N_1441,N_1381,N_1398);
nand U1442 (N_1442,N_1401,N_1418);
or U1443 (N_1443,N_1426,N_1403);
nor U1444 (N_1444,N_1413,N_1431);
and U1445 (N_1445,N_1438,N_1400);
and U1446 (N_1446,N_1407,N_1425);
nand U1447 (N_1447,N_1394,N_1423);
nor U1448 (N_1448,N_1422,N_1390);
nand U1449 (N_1449,N_1385,N_1416);
nand U1450 (N_1450,N_1414,N_1396);
nand U1451 (N_1451,N_1383,N_1430);
nor U1452 (N_1452,N_1391,N_1437);
or U1453 (N_1453,N_1380,N_1412);
and U1454 (N_1454,N_1402,N_1427);
nand U1455 (N_1455,N_1393,N_1405);
or U1456 (N_1456,N_1388,N_1395);
nor U1457 (N_1457,N_1421,N_1424);
xnor U1458 (N_1458,N_1410,N_1432);
and U1459 (N_1459,N_1389,N_1406);
or U1460 (N_1460,N_1436,N_1408);
nor U1461 (N_1461,N_1428,N_1409);
or U1462 (N_1462,N_1420,N_1434);
and U1463 (N_1463,N_1439,N_1411);
and U1464 (N_1464,N_1386,N_1387);
and U1465 (N_1465,N_1435,N_1404);
nor U1466 (N_1466,N_1399,N_1429);
and U1467 (N_1467,N_1419,N_1384);
nand U1468 (N_1468,N_1397,N_1392);
or U1469 (N_1469,N_1382,N_1433);
or U1470 (N_1470,N_1412,N_1430);
and U1471 (N_1471,N_1412,N_1388);
nand U1472 (N_1472,N_1420,N_1415);
and U1473 (N_1473,N_1427,N_1390);
and U1474 (N_1474,N_1407,N_1386);
nand U1475 (N_1475,N_1408,N_1420);
or U1476 (N_1476,N_1416,N_1390);
and U1477 (N_1477,N_1430,N_1397);
nand U1478 (N_1478,N_1409,N_1437);
or U1479 (N_1479,N_1409,N_1413);
nand U1480 (N_1480,N_1426,N_1414);
or U1481 (N_1481,N_1395,N_1434);
or U1482 (N_1482,N_1400,N_1411);
nor U1483 (N_1483,N_1438,N_1415);
or U1484 (N_1484,N_1414,N_1415);
nor U1485 (N_1485,N_1438,N_1412);
nor U1486 (N_1486,N_1419,N_1394);
and U1487 (N_1487,N_1393,N_1385);
xnor U1488 (N_1488,N_1394,N_1386);
nand U1489 (N_1489,N_1399,N_1411);
or U1490 (N_1490,N_1430,N_1389);
or U1491 (N_1491,N_1428,N_1382);
nor U1492 (N_1492,N_1402,N_1394);
nand U1493 (N_1493,N_1415,N_1429);
and U1494 (N_1494,N_1410,N_1414);
nand U1495 (N_1495,N_1399,N_1439);
nor U1496 (N_1496,N_1422,N_1393);
nor U1497 (N_1497,N_1432,N_1402);
and U1498 (N_1498,N_1431,N_1388);
and U1499 (N_1499,N_1407,N_1390);
and U1500 (N_1500,N_1490,N_1452);
or U1501 (N_1501,N_1483,N_1468);
nor U1502 (N_1502,N_1477,N_1446);
or U1503 (N_1503,N_1471,N_1481);
nor U1504 (N_1504,N_1461,N_1475);
nor U1505 (N_1505,N_1476,N_1453);
nor U1506 (N_1506,N_1469,N_1458);
nand U1507 (N_1507,N_1442,N_1450);
and U1508 (N_1508,N_1467,N_1495);
nor U1509 (N_1509,N_1457,N_1440);
nand U1510 (N_1510,N_1464,N_1482);
nor U1511 (N_1511,N_1478,N_1445);
nor U1512 (N_1512,N_1448,N_1463);
and U1513 (N_1513,N_1447,N_1472);
nand U1514 (N_1514,N_1462,N_1474);
and U1515 (N_1515,N_1498,N_1441);
nor U1516 (N_1516,N_1499,N_1496);
nand U1517 (N_1517,N_1454,N_1493);
and U1518 (N_1518,N_1480,N_1459);
and U1519 (N_1519,N_1456,N_1479);
nor U1520 (N_1520,N_1486,N_1492);
nand U1521 (N_1521,N_1444,N_1488);
and U1522 (N_1522,N_1460,N_1485);
and U1523 (N_1523,N_1473,N_1449);
nand U1524 (N_1524,N_1455,N_1487);
nor U1525 (N_1525,N_1470,N_1494);
nor U1526 (N_1526,N_1443,N_1491);
nor U1527 (N_1527,N_1497,N_1451);
and U1528 (N_1528,N_1466,N_1484);
nand U1529 (N_1529,N_1489,N_1465);
xnor U1530 (N_1530,N_1473,N_1499);
and U1531 (N_1531,N_1474,N_1471);
and U1532 (N_1532,N_1452,N_1458);
and U1533 (N_1533,N_1448,N_1475);
and U1534 (N_1534,N_1470,N_1446);
or U1535 (N_1535,N_1455,N_1486);
nor U1536 (N_1536,N_1458,N_1467);
nor U1537 (N_1537,N_1473,N_1463);
or U1538 (N_1538,N_1467,N_1449);
or U1539 (N_1539,N_1492,N_1470);
and U1540 (N_1540,N_1456,N_1468);
nor U1541 (N_1541,N_1483,N_1469);
nand U1542 (N_1542,N_1459,N_1483);
or U1543 (N_1543,N_1496,N_1487);
nand U1544 (N_1544,N_1451,N_1447);
and U1545 (N_1545,N_1457,N_1464);
or U1546 (N_1546,N_1465,N_1453);
nand U1547 (N_1547,N_1441,N_1496);
nor U1548 (N_1548,N_1466,N_1446);
and U1549 (N_1549,N_1460,N_1495);
nor U1550 (N_1550,N_1467,N_1498);
nor U1551 (N_1551,N_1476,N_1460);
nand U1552 (N_1552,N_1492,N_1459);
and U1553 (N_1553,N_1442,N_1468);
nor U1554 (N_1554,N_1474,N_1475);
or U1555 (N_1555,N_1496,N_1452);
xnor U1556 (N_1556,N_1486,N_1499);
nand U1557 (N_1557,N_1449,N_1495);
or U1558 (N_1558,N_1468,N_1453);
nor U1559 (N_1559,N_1447,N_1440);
nor U1560 (N_1560,N_1529,N_1508);
and U1561 (N_1561,N_1518,N_1549);
nor U1562 (N_1562,N_1557,N_1525);
xor U1563 (N_1563,N_1539,N_1548);
nand U1564 (N_1564,N_1538,N_1542);
or U1565 (N_1565,N_1507,N_1500);
or U1566 (N_1566,N_1510,N_1553);
and U1567 (N_1567,N_1530,N_1514);
nand U1568 (N_1568,N_1502,N_1535);
xnor U1569 (N_1569,N_1552,N_1536);
nand U1570 (N_1570,N_1540,N_1545);
nand U1571 (N_1571,N_1520,N_1551);
nand U1572 (N_1572,N_1547,N_1555);
nand U1573 (N_1573,N_1503,N_1519);
nand U1574 (N_1574,N_1527,N_1558);
nor U1575 (N_1575,N_1528,N_1521);
and U1576 (N_1576,N_1506,N_1516);
nor U1577 (N_1577,N_1541,N_1559);
and U1578 (N_1578,N_1534,N_1544);
nand U1579 (N_1579,N_1509,N_1537);
nor U1580 (N_1580,N_1515,N_1501);
and U1581 (N_1581,N_1556,N_1504);
and U1582 (N_1582,N_1517,N_1533);
nand U1583 (N_1583,N_1546,N_1543);
or U1584 (N_1584,N_1513,N_1554);
nor U1585 (N_1585,N_1505,N_1526);
nor U1586 (N_1586,N_1511,N_1512);
and U1587 (N_1587,N_1523,N_1531);
nor U1588 (N_1588,N_1524,N_1522);
nor U1589 (N_1589,N_1550,N_1532);
nand U1590 (N_1590,N_1514,N_1520);
xor U1591 (N_1591,N_1541,N_1507);
or U1592 (N_1592,N_1528,N_1543);
nor U1593 (N_1593,N_1552,N_1500);
nand U1594 (N_1594,N_1528,N_1519);
and U1595 (N_1595,N_1544,N_1553);
nor U1596 (N_1596,N_1558,N_1529);
or U1597 (N_1597,N_1540,N_1550);
nand U1598 (N_1598,N_1540,N_1552);
and U1599 (N_1599,N_1540,N_1531);
and U1600 (N_1600,N_1522,N_1559);
or U1601 (N_1601,N_1527,N_1506);
nor U1602 (N_1602,N_1531,N_1519);
or U1603 (N_1603,N_1529,N_1537);
and U1604 (N_1604,N_1537,N_1528);
or U1605 (N_1605,N_1525,N_1556);
nor U1606 (N_1606,N_1543,N_1554);
nor U1607 (N_1607,N_1536,N_1540);
or U1608 (N_1608,N_1555,N_1554);
or U1609 (N_1609,N_1514,N_1528);
nor U1610 (N_1610,N_1537,N_1550);
nor U1611 (N_1611,N_1514,N_1549);
nor U1612 (N_1612,N_1505,N_1530);
or U1613 (N_1613,N_1546,N_1557);
nor U1614 (N_1614,N_1514,N_1505);
nor U1615 (N_1615,N_1538,N_1524);
nor U1616 (N_1616,N_1512,N_1555);
and U1617 (N_1617,N_1539,N_1557);
nand U1618 (N_1618,N_1509,N_1552);
and U1619 (N_1619,N_1515,N_1549);
or U1620 (N_1620,N_1577,N_1562);
xnor U1621 (N_1621,N_1593,N_1600);
and U1622 (N_1622,N_1566,N_1586);
and U1623 (N_1623,N_1585,N_1597);
or U1624 (N_1624,N_1564,N_1565);
and U1625 (N_1625,N_1584,N_1598);
or U1626 (N_1626,N_1568,N_1614);
nand U1627 (N_1627,N_1604,N_1610);
nor U1628 (N_1628,N_1607,N_1574);
or U1629 (N_1629,N_1560,N_1587);
xor U1630 (N_1630,N_1606,N_1609);
and U1631 (N_1631,N_1580,N_1592);
and U1632 (N_1632,N_1575,N_1567);
or U1633 (N_1633,N_1578,N_1608);
or U1634 (N_1634,N_1591,N_1589);
and U1635 (N_1635,N_1582,N_1576);
or U1636 (N_1636,N_1596,N_1617);
and U1637 (N_1637,N_1601,N_1603);
and U1638 (N_1638,N_1581,N_1602);
nor U1639 (N_1639,N_1605,N_1613);
nor U1640 (N_1640,N_1571,N_1573);
nor U1641 (N_1641,N_1594,N_1569);
nor U1642 (N_1642,N_1618,N_1579);
nand U1643 (N_1643,N_1595,N_1588);
nor U1644 (N_1644,N_1616,N_1611);
nor U1645 (N_1645,N_1619,N_1570);
nor U1646 (N_1646,N_1563,N_1583);
nand U1647 (N_1647,N_1572,N_1615);
nor U1648 (N_1648,N_1561,N_1590);
nor U1649 (N_1649,N_1599,N_1612);
nor U1650 (N_1650,N_1609,N_1605);
nor U1651 (N_1651,N_1593,N_1611);
or U1652 (N_1652,N_1589,N_1614);
and U1653 (N_1653,N_1562,N_1611);
nand U1654 (N_1654,N_1586,N_1585);
and U1655 (N_1655,N_1585,N_1601);
nand U1656 (N_1656,N_1598,N_1605);
nor U1657 (N_1657,N_1593,N_1564);
nor U1658 (N_1658,N_1590,N_1607);
nand U1659 (N_1659,N_1609,N_1560);
nor U1660 (N_1660,N_1607,N_1581);
nand U1661 (N_1661,N_1576,N_1613);
nand U1662 (N_1662,N_1586,N_1561);
or U1663 (N_1663,N_1576,N_1610);
and U1664 (N_1664,N_1581,N_1605);
or U1665 (N_1665,N_1587,N_1581);
or U1666 (N_1666,N_1566,N_1611);
nor U1667 (N_1667,N_1598,N_1575);
or U1668 (N_1668,N_1589,N_1618);
nand U1669 (N_1669,N_1601,N_1578);
or U1670 (N_1670,N_1581,N_1597);
nor U1671 (N_1671,N_1603,N_1605);
or U1672 (N_1672,N_1602,N_1599);
and U1673 (N_1673,N_1579,N_1600);
nor U1674 (N_1674,N_1602,N_1605);
nor U1675 (N_1675,N_1585,N_1573);
and U1676 (N_1676,N_1604,N_1573);
and U1677 (N_1677,N_1567,N_1583);
nor U1678 (N_1678,N_1582,N_1607);
and U1679 (N_1679,N_1566,N_1565);
nor U1680 (N_1680,N_1670,N_1673);
and U1681 (N_1681,N_1635,N_1642);
nand U1682 (N_1682,N_1621,N_1643);
or U1683 (N_1683,N_1623,N_1657);
nor U1684 (N_1684,N_1662,N_1676);
nor U1685 (N_1685,N_1656,N_1627);
nor U1686 (N_1686,N_1653,N_1649);
nor U1687 (N_1687,N_1675,N_1658);
nor U1688 (N_1688,N_1644,N_1634);
or U1689 (N_1689,N_1629,N_1672);
nor U1690 (N_1690,N_1678,N_1630);
nor U1691 (N_1691,N_1622,N_1628);
or U1692 (N_1692,N_1659,N_1645);
nand U1693 (N_1693,N_1661,N_1625);
and U1694 (N_1694,N_1654,N_1647);
nand U1695 (N_1695,N_1636,N_1640);
and U1696 (N_1696,N_1665,N_1638);
nand U1697 (N_1697,N_1639,N_1674);
nor U1698 (N_1698,N_1669,N_1668);
and U1699 (N_1699,N_1648,N_1637);
xnor U1700 (N_1700,N_1631,N_1671);
nor U1701 (N_1701,N_1641,N_1651);
or U1702 (N_1702,N_1655,N_1620);
or U1703 (N_1703,N_1667,N_1677);
nand U1704 (N_1704,N_1652,N_1633);
nand U1705 (N_1705,N_1650,N_1666);
and U1706 (N_1706,N_1679,N_1646);
nand U1707 (N_1707,N_1660,N_1632);
nand U1708 (N_1708,N_1664,N_1626);
nor U1709 (N_1709,N_1663,N_1624);
or U1710 (N_1710,N_1674,N_1635);
nand U1711 (N_1711,N_1634,N_1667);
nor U1712 (N_1712,N_1623,N_1639);
and U1713 (N_1713,N_1634,N_1674);
nand U1714 (N_1714,N_1655,N_1629);
nor U1715 (N_1715,N_1662,N_1650);
and U1716 (N_1716,N_1651,N_1668);
or U1717 (N_1717,N_1653,N_1628);
and U1718 (N_1718,N_1638,N_1631);
nand U1719 (N_1719,N_1643,N_1665);
nand U1720 (N_1720,N_1626,N_1667);
nor U1721 (N_1721,N_1654,N_1675);
nand U1722 (N_1722,N_1669,N_1654);
nand U1723 (N_1723,N_1676,N_1629);
nand U1724 (N_1724,N_1670,N_1677);
nor U1725 (N_1725,N_1637,N_1664);
nor U1726 (N_1726,N_1661,N_1660);
or U1727 (N_1727,N_1667,N_1673);
nand U1728 (N_1728,N_1649,N_1679);
and U1729 (N_1729,N_1654,N_1640);
nor U1730 (N_1730,N_1630,N_1664);
nand U1731 (N_1731,N_1630,N_1625);
and U1732 (N_1732,N_1639,N_1657);
and U1733 (N_1733,N_1654,N_1671);
nor U1734 (N_1734,N_1667,N_1669);
nor U1735 (N_1735,N_1658,N_1669);
or U1736 (N_1736,N_1674,N_1660);
nor U1737 (N_1737,N_1644,N_1668);
nand U1738 (N_1738,N_1664,N_1675);
or U1739 (N_1739,N_1621,N_1624);
or U1740 (N_1740,N_1696,N_1685);
nand U1741 (N_1741,N_1686,N_1734);
and U1742 (N_1742,N_1681,N_1680);
and U1743 (N_1743,N_1739,N_1701);
nor U1744 (N_1744,N_1692,N_1738);
or U1745 (N_1745,N_1724,N_1730);
nor U1746 (N_1746,N_1712,N_1693);
or U1747 (N_1747,N_1699,N_1711);
xnor U1748 (N_1748,N_1715,N_1736);
nor U1749 (N_1749,N_1705,N_1684);
xor U1750 (N_1750,N_1718,N_1716);
or U1751 (N_1751,N_1700,N_1710);
and U1752 (N_1752,N_1726,N_1731);
and U1753 (N_1753,N_1735,N_1720);
nor U1754 (N_1754,N_1707,N_1683);
and U1755 (N_1755,N_1698,N_1703);
or U1756 (N_1756,N_1725,N_1708);
nand U1757 (N_1757,N_1723,N_1706);
or U1758 (N_1758,N_1721,N_1737);
and U1759 (N_1759,N_1728,N_1722);
nand U1760 (N_1760,N_1694,N_1727);
and U1761 (N_1761,N_1695,N_1709);
and U1762 (N_1762,N_1713,N_1688);
and U1763 (N_1763,N_1682,N_1704);
nor U1764 (N_1764,N_1689,N_1719);
nor U1765 (N_1765,N_1687,N_1690);
nor U1766 (N_1766,N_1729,N_1717);
nand U1767 (N_1767,N_1732,N_1702);
and U1768 (N_1768,N_1691,N_1714);
nand U1769 (N_1769,N_1697,N_1733);
and U1770 (N_1770,N_1710,N_1739);
nand U1771 (N_1771,N_1686,N_1715);
nand U1772 (N_1772,N_1729,N_1698);
or U1773 (N_1773,N_1711,N_1726);
nor U1774 (N_1774,N_1720,N_1721);
and U1775 (N_1775,N_1730,N_1689);
nor U1776 (N_1776,N_1704,N_1734);
nand U1777 (N_1777,N_1720,N_1705);
and U1778 (N_1778,N_1735,N_1716);
nor U1779 (N_1779,N_1708,N_1699);
or U1780 (N_1780,N_1702,N_1680);
nor U1781 (N_1781,N_1703,N_1697);
or U1782 (N_1782,N_1680,N_1698);
nand U1783 (N_1783,N_1707,N_1739);
nor U1784 (N_1784,N_1687,N_1698);
nand U1785 (N_1785,N_1705,N_1716);
nor U1786 (N_1786,N_1705,N_1693);
or U1787 (N_1787,N_1705,N_1721);
or U1788 (N_1788,N_1730,N_1702);
xor U1789 (N_1789,N_1706,N_1717);
and U1790 (N_1790,N_1689,N_1733);
nand U1791 (N_1791,N_1703,N_1708);
nor U1792 (N_1792,N_1711,N_1694);
or U1793 (N_1793,N_1720,N_1683);
or U1794 (N_1794,N_1701,N_1728);
nand U1795 (N_1795,N_1712,N_1728);
nand U1796 (N_1796,N_1681,N_1728);
and U1797 (N_1797,N_1703,N_1712);
nand U1798 (N_1798,N_1717,N_1712);
and U1799 (N_1799,N_1724,N_1711);
or U1800 (N_1800,N_1794,N_1761);
nor U1801 (N_1801,N_1747,N_1742);
or U1802 (N_1802,N_1785,N_1795);
nor U1803 (N_1803,N_1753,N_1789);
or U1804 (N_1804,N_1788,N_1783);
and U1805 (N_1805,N_1786,N_1745);
nor U1806 (N_1806,N_1782,N_1767);
nor U1807 (N_1807,N_1778,N_1757);
or U1808 (N_1808,N_1780,N_1762);
nor U1809 (N_1809,N_1743,N_1769);
nor U1810 (N_1810,N_1760,N_1772);
nand U1811 (N_1811,N_1775,N_1758);
or U1812 (N_1812,N_1746,N_1744);
or U1813 (N_1813,N_1799,N_1787);
or U1814 (N_1814,N_1749,N_1764);
nand U1815 (N_1815,N_1740,N_1748);
nand U1816 (N_1816,N_1779,N_1751);
nand U1817 (N_1817,N_1752,N_1797);
or U1818 (N_1818,N_1770,N_1756);
or U1819 (N_1819,N_1773,N_1765);
nand U1820 (N_1820,N_1784,N_1759);
nand U1821 (N_1821,N_1754,N_1750);
and U1822 (N_1822,N_1771,N_1741);
nand U1823 (N_1823,N_1774,N_1792);
nand U1824 (N_1824,N_1781,N_1791);
nand U1825 (N_1825,N_1796,N_1766);
or U1826 (N_1826,N_1790,N_1776);
nand U1827 (N_1827,N_1793,N_1763);
nor U1828 (N_1828,N_1768,N_1755);
nand U1829 (N_1829,N_1798,N_1777);
nand U1830 (N_1830,N_1775,N_1762);
and U1831 (N_1831,N_1771,N_1791);
nor U1832 (N_1832,N_1740,N_1799);
and U1833 (N_1833,N_1784,N_1775);
nor U1834 (N_1834,N_1794,N_1786);
or U1835 (N_1835,N_1740,N_1798);
and U1836 (N_1836,N_1795,N_1757);
nand U1837 (N_1837,N_1765,N_1745);
nor U1838 (N_1838,N_1794,N_1789);
nor U1839 (N_1839,N_1771,N_1748);
and U1840 (N_1840,N_1766,N_1789);
or U1841 (N_1841,N_1749,N_1784);
and U1842 (N_1842,N_1778,N_1742);
and U1843 (N_1843,N_1757,N_1753);
nor U1844 (N_1844,N_1766,N_1788);
and U1845 (N_1845,N_1741,N_1788);
and U1846 (N_1846,N_1780,N_1767);
nor U1847 (N_1847,N_1769,N_1768);
nand U1848 (N_1848,N_1785,N_1776);
nor U1849 (N_1849,N_1776,N_1742);
nor U1850 (N_1850,N_1766,N_1748);
nand U1851 (N_1851,N_1791,N_1798);
and U1852 (N_1852,N_1756,N_1740);
and U1853 (N_1853,N_1760,N_1779);
and U1854 (N_1854,N_1780,N_1799);
nand U1855 (N_1855,N_1792,N_1797);
nor U1856 (N_1856,N_1765,N_1761);
or U1857 (N_1857,N_1773,N_1748);
or U1858 (N_1858,N_1796,N_1795);
nor U1859 (N_1859,N_1770,N_1798);
or U1860 (N_1860,N_1841,N_1839);
or U1861 (N_1861,N_1858,N_1853);
or U1862 (N_1862,N_1859,N_1817);
nand U1863 (N_1863,N_1813,N_1849);
nor U1864 (N_1864,N_1847,N_1821);
and U1865 (N_1865,N_1838,N_1844);
or U1866 (N_1866,N_1830,N_1814);
nor U1867 (N_1867,N_1843,N_1842);
nor U1868 (N_1868,N_1845,N_1804);
nand U1869 (N_1869,N_1827,N_1831);
nand U1870 (N_1870,N_1802,N_1837);
xor U1871 (N_1871,N_1832,N_1856);
and U1872 (N_1872,N_1820,N_1810);
xnor U1873 (N_1873,N_1852,N_1850);
nor U1874 (N_1874,N_1840,N_1836);
nand U1875 (N_1875,N_1829,N_1809);
nor U1876 (N_1876,N_1819,N_1855);
nor U1877 (N_1877,N_1833,N_1801);
and U1878 (N_1878,N_1826,N_1806);
nor U1879 (N_1879,N_1825,N_1851);
nor U1880 (N_1880,N_1812,N_1846);
nor U1881 (N_1881,N_1823,N_1828);
or U1882 (N_1882,N_1803,N_1835);
nor U1883 (N_1883,N_1808,N_1848);
nand U1884 (N_1884,N_1857,N_1816);
or U1885 (N_1885,N_1807,N_1854);
and U1886 (N_1886,N_1824,N_1822);
and U1887 (N_1887,N_1818,N_1805);
or U1888 (N_1888,N_1815,N_1811);
or U1889 (N_1889,N_1800,N_1834);
nand U1890 (N_1890,N_1837,N_1815);
or U1891 (N_1891,N_1812,N_1841);
and U1892 (N_1892,N_1836,N_1807);
xnor U1893 (N_1893,N_1828,N_1806);
or U1894 (N_1894,N_1817,N_1812);
nor U1895 (N_1895,N_1820,N_1856);
or U1896 (N_1896,N_1816,N_1829);
nor U1897 (N_1897,N_1803,N_1850);
nand U1898 (N_1898,N_1852,N_1859);
nand U1899 (N_1899,N_1839,N_1842);
nor U1900 (N_1900,N_1835,N_1844);
nor U1901 (N_1901,N_1831,N_1851);
and U1902 (N_1902,N_1803,N_1820);
or U1903 (N_1903,N_1819,N_1806);
nor U1904 (N_1904,N_1848,N_1842);
and U1905 (N_1905,N_1827,N_1806);
or U1906 (N_1906,N_1835,N_1818);
nor U1907 (N_1907,N_1807,N_1847);
nor U1908 (N_1908,N_1812,N_1851);
nand U1909 (N_1909,N_1834,N_1848);
nand U1910 (N_1910,N_1831,N_1850);
nand U1911 (N_1911,N_1818,N_1827);
nor U1912 (N_1912,N_1814,N_1820);
and U1913 (N_1913,N_1823,N_1814);
nor U1914 (N_1914,N_1857,N_1800);
nand U1915 (N_1915,N_1848,N_1855);
nor U1916 (N_1916,N_1848,N_1815);
and U1917 (N_1917,N_1827,N_1811);
nand U1918 (N_1918,N_1842,N_1859);
nor U1919 (N_1919,N_1823,N_1809);
or U1920 (N_1920,N_1862,N_1861);
or U1921 (N_1921,N_1897,N_1905);
nand U1922 (N_1922,N_1884,N_1874);
and U1923 (N_1923,N_1889,N_1871);
nand U1924 (N_1924,N_1877,N_1864);
nand U1925 (N_1925,N_1895,N_1865);
nor U1926 (N_1926,N_1869,N_1885);
nand U1927 (N_1927,N_1913,N_1898);
nor U1928 (N_1928,N_1919,N_1917);
nand U1929 (N_1929,N_1879,N_1914);
or U1930 (N_1930,N_1915,N_1866);
nor U1931 (N_1931,N_1873,N_1909);
or U1932 (N_1932,N_1880,N_1860);
nand U1933 (N_1933,N_1907,N_1902);
nand U1934 (N_1934,N_1908,N_1867);
and U1935 (N_1935,N_1901,N_1887);
and U1936 (N_1936,N_1875,N_1886);
nor U1937 (N_1937,N_1863,N_1896);
or U1938 (N_1938,N_1868,N_1872);
and U1939 (N_1939,N_1882,N_1888);
nor U1940 (N_1940,N_1899,N_1894);
or U1941 (N_1941,N_1878,N_1916);
nor U1942 (N_1942,N_1890,N_1892);
nand U1943 (N_1943,N_1876,N_1893);
and U1944 (N_1944,N_1900,N_1918);
nand U1945 (N_1945,N_1903,N_1870);
nor U1946 (N_1946,N_1906,N_1904);
and U1947 (N_1947,N_1911,N_1883);
or U1948 (N_1948,N_1910,N_1881);
nor U1949 (N_1949,N_1912,N_1891);
and U1950 (N_1950,N_1917,N_1914);
or U1951 (N_1951,N_1890,N_1914);
nand U1952 (N_1952,N_1906,N_1895);
nor U1953 (N_1953,N_1860,N_1900);
or U1954 (N_1954,N_1892,N_1901);
nor U1955 (N_1955,N_1867,N_1898);
nor U1956 (N_1956,N_1897,N_1864);
nor U1957 (N_1957,N_1864,N_1865);
nor U1958 (N_1958,N_1882,N_1867);
and U1959 (N_1959,N_1892,N_1860);
nand U1960 (N_1960,N_1896,N_1878);
nand U1961 (N_1961,N_1885,N_1862);
nand U1962 (N_1962,N_1905,N_1914);
nor U1963 (N_1963,N_1881,N_1905);
xnor U1964 (N_1964,N_1871,N_1873);
or U1965 (N_1965,N_1891,N_1918);
and U1966 (N_1966,N_1887,N_1875);
nand U1967 (N_1967,N_1877,N_1870);
nor U1968 (N_1968,N_1919,N_1883);
nand U1969 (N_1969,N_1886,N_1908);
and U1970 (N_1970,N_1896,N_1897);
nor U1971 (N_1971,N_1897,N_1918);
nand U1972 (N_1972,N_1915,N_1907);
nor U1973 (N_1973,N_1860,N_1865);
nor U1974 (N_1974,N_1918,N_1908);
nand U1975 (N_1975,N_1902,N_1889);
nand U1976 (N_1976,N_1902,N_1891);
nand U1977 (N_1977,N_1897,N_1915);
or U1978 (N_1978,N_1875,N_1866);
nand U1979 (N_1979,N_1876,N_1895);
nand U1980 (N_1980,N_1965,N_1967);
and U1981 (N_1981,N_1949,N_1974);
or U1982 (N_1982,N_1963,N_1926);
and U1983 (N_1983,N_1935,N_1947);
nor U1984 (N_1984,N_1978,N_1933);
and U1985 (N_1985,N_1951,N_1964);
nor U1986 (N_1986,N_1971,N_1943);
nor U1987 (N_1987,N_1958,N_1946);
or U1988 (N_1988,N_1975,N_1938);
and U1989 (N_1989,N_1970,N_1928);
nand U1990 (N_1990,N_1957,N_1948);
or U1991 (N_1991,N_1972,N_1931);
xnor U1992 (N_1992,N_1959,N_1930);
nand U1993 (N_1993,N_1962,N_1945);
nor U1994 (N_1994,N_1927,N_1953);
and U1995 (N_1995,N_1923,N_1954);
nand U1996 (N_1996,N_1929,N_1921);
or U1997 (N_1997,N_1976,N_1924);
and U1998 (N_1998,N_1955,N_1956);
or U1999 (N_1999,N_1973,N_1937);
or U2000 (N_2000,N_1969,N_1950);
or U2001 (N_2001,N_1936,N_1942);
nand U2002 (N_2002,N_1932,N_1944);
nor U2003 (N_2003,N_1939,N_1920);
or U2004 (N_2004,N_1922,N_1966);
nand U2005 (N_2005,N_1934,N_1952);
and U2006 (N_2006,N_1925,N_1977);
and U2007 (N_2007,N_1960,N_1941);
nor U2008 (N_2008,N_1979,N_1940);
and U2009 (N_2009,N_1968,N_1961);
or U2010 (N_2010,N_1978,N_1956);
nand U2011 (N_2011,N_1942,N_1974);
nor U2012 (N_2012,N_1947,N_1954);
and U2013 (N_2013,N_1955,N_1960);
or U2014 (N_2014,N_1922,N_1974);
or U2015 (N_2015,N_1924,N_1972);
and U2016 (N_2016,N_1921,N_1963);
or U2017 (N_2017,N_1977,N_1923);
nor U2018 (N_2018,N_1970,N_1923);
or U2019 (N_2019,N_1939,N_1935);
xnor U2020 (N_2020,N_1931,N_1965);
nand U2021 (N_2021,N_1971,N_1950);
or U2022 (N_2022,N_1952,N_1945);
nor U2023 (N_2023,N_1933,N_1927);
and U2024 (N_2024,N_1967,N_1971);
nor U2025 (N_2025,N_1955,N_1923);
nor U2026 (N_2026,N_1928,N_1947);
and U2027 (N_2027,N_1956,N_1964);
and U2028 (N_2028,N_1947,N_1962);
or U2029 (N_2029,N_1944,N_1948);
or U2030 (N_2030,N_1929,N_1963);
nor U2031 (N_2031,N_1936,N_1952);
nand U2032 (N_2032,N_1934,N_1936);
and U2033 (N_2033,N_1935,N_1925);
nand U2034 (N_2034,N_1949,N_1935);
and U2035 (N_2035,N_1921,N_1932);
nand U2036 (N_2036,N_1966,N_1978);
nor U2037 (N_2037,N_1951,N_1952);
nand U2038 (N_2038,N_1932,N_1970);
or U2039 (N_2039,N_1978,N_1972);
and U2040 (N_2040,N_1992,N_2000);
nand U2041 (N_2041,N_2037,N_1980);
nor U2042 (N_2042,N_2016,N_2026);
or U2043 (N_2043,N_1995,N_1991);
nand U2044 (N_2044,N_2015,N_2020);
nand U2045 (N_2045,N_2024,N_2019);
and U2046 (N_2046,N_2014,N_2012);
nor U2047 (N_2047,N_1988,N_2033);
nor U2048 (N_2048,N_2010,N_1981);
xnor U2049 (N_2049,N_2017,N_2013);
or U2050 (N_2050,N_1984,N_2008);
nand U2051 (N_2051,N_1990,N_2038);
and U2052 (N_2052,N_2005,N_2006);
and U2053 (N_2053,N_2021,N_2039);
nor U2054 (N_2054,N_2035,N_1999);
and U2055 (N_2055,N_1993,N_2029);
and U2056 (N_2056,N_2023,N_1983);
or U2057 (N_2057,N_2009,N_2027);
and U2058 (N_2058,N_1994,N_1986);
nor U2059 (N_2059,N_1998,N_2031);
nand U2060 (N_2060,N_2034,N_2007);
and U2061 (N_2061,N_2025,N_2011);
and U2062 (N_2062,N_2018,N_2001);
nor U2063 (N_2063,N_2028,N_1982);
nand U2064 (N_2064,N_2003,N_1989);
nand U2065 (N_2065,N_2022,N_2004);
or U2066 (N_2066,N_1997,N_2032);
nor U2067 (N_2067,N_2036,N_1987);
and U2068 (N_2068,N_1985,N_2002);
and U2069 (N_2069,N_1996,N_2030);
and U2070 (N_2070,N_2032,N_1999);
nand U2071 (N_2071,N_2007,N_2024);
nand U2072 (N_2072,N_1987,N_2039);
nand U2073 (N_2073,N_2017,N_1984);
and U2074 (N_2074,N_2025,N_2039);
nand U2075 (N_2075,N_2033,N_2005);
and U2076 (N_2076,N_2018,N_2003);
nor U2077 (N_2077,N_2014,N_2005);
nor U2078 (N_2078,N_2021,N_2025);
nor U2079 (N_2079,N_2027,N_2024);
or U2080 (N_2080,N_2006,N_2030);
and U2081 (N_2081,N_1998,N_2002);
and U2082 (N_2082,N_2037,N_1986);
nand U2083 (N_2083,N_1981,N_1991);
nor U2084 (N_2084,N_2032,N_1984);
and U2085 (N_2085,N_2019,N_2016);
nand U2086 (N_2086,N_1980,N_2034);
nand U2087 (N_2087,N_2026,N_2019);
and U2088 (N_2088,N_1986,N_2034);
and U2089 (N_2089,N_2036,N_1984);
nand U2090 (N_2090,N_2003,N_1993);
nand U2091 (N_2091,N_2028,N_2022);
nand U2092 (N_2092,N_1993,N_2027);
nor U2093 (N_2093,N_2030,N_2014);
or U2094 (N_2094,N_2015,N_2030);
and U2095 (N_2095,N_1995,N_1994);
nand U2096 (N_2096,N_2020,N_1985);
and U2097 (N_2097,N_2024,N_2002);
nor U2098 (N_2098,N_2017,N_1995);
nor U2099 (N_2099,N_2007,N_1995);
or U2100 (N_2100,N_2091,N_2070);
or U2101 (N_2101,N_2065,N_2087);
xnor U2102 (N_2102,N_2088,N_2071);
or U2103 (N_2103,N_2099,N_2050);
nor U2104 (N_2104,N_2054,N_2081);
nor U2105 (N_2105,N_2043,N_2083);
or U2106 (N_2106,N_2045,N_2041);
nand U2107 (N_2107,N_2058,N_2095);
or U2108 (N_2108,N_2049,N_2079);
nor U2109 (N_2109,N_2063,N_2076);
and U2110 (N_2110,N_2072,N_2046);
and U2111 (N_2111,N_2060,N_2064);
nor U2112 (N_2112,N_2084,N_2082);
xnor U2113 (N_2113,N_2086,N_2097);
nand U2114 (N_2114,N_2048,N_2074);
or U2115 (N_2115,N_2059,N_2055);
or U2116 (N_2116,N_2062,N_2042);
nand U2117 (N_2117,N_2094,N_2096);
and U2118 (N_2118,N_2075,N_2080);
and U2119 (N_2119,N_2090,N_2061);
nand U2120 (N_2120,N_2040,N_2053);
nor U2121 (N_2121,N_2077,N_2078);
or U2122 (N_2122,N_2057,N_2089);
and U2123 (N_2123,N_2056,N_2092);
and U2124 (N_2124,N_2051,N_2093);
nand U2125 (N_2125,N_2052,N_2044);
nor U2126 (N_2126,N_2047,N_2067);
or U2127 (N_2127,N_2069,N_2066);
nor U2128 (N_2128,N_2098,N_2085);
nor U2129 (N_2129,N_2073,N_2068);
or U2130 (N_2130,N_2077,N_2063);
xnor U2131 (N_2131,N_2068,N_2066);
or U2132 (N_2132,N_2074,N_2097);
nor U2133 (N_2133,N_2040,N_2050);
nand U2134 (N_2134,N_2071,N_2090);
or U2135 (N_2135,N_2062,N_2057);
nor U2136 (N_2136,N_2042,N_2065);
or U2137 (N_2137,N_2080,N_2054);
nand U2138 (N_2138,N_2080,N_2071);
and U2139 (N_2139,N_2094,N_2041);
nand U2140 (N_2140,N_2080,N_2099);
and U2141 (N_2141,N_2082,N_2068);
or U2142 (N_2142,N_2061,N_2049);
and U2143 (N_2143,N_2073,N_2078);
and U2144 (N_2144,N_2063,N_2060);
nand U2145 (N_2145,N_2063,N_2043);
nor U2146 (N_2146,N_2086,N_2099);
nand U2147 (N_2147,N_2062,N_2074);
nand U2148 (N_2148,N_2084,N_2085);
or U2149 (N_2149,N_2064,N_2077);
or U2150 (N_2150,N_2049,N_2042);
nor U2151 (N_2151,N_2066,N_2097);
or U2152 (N_2152,N_2057,N_2070);
and U2153 (N_2153,N_2046,N_2073);
or U2154 (N_2154,N_2080,N_2061);
nand U2155 (N_2155,N_2091,N_2057);
and U2156 (N_2156,N_2072,N_2090);
or U2157 (N_2157,N_2085,N_2045);
or U2158 (N_2158,N_2040,N_2051);
and U2159 (N_2159,N_2080,N_2097);
xor U2160 (N_2160,N_2151,N_2142);
nand U2161 (N_2161,N_2128,N_2141);
or U2162 (N_2162,N_2123,N_2137);
nand U2163 (N_2163,N_2153,N_2158);
nand U2164 (N_2164,N_2126,N_2109);
xnor U2165 (N_2165,N_2134,N_2101);
and U2166 (N_2166,N_2148,N_2102);
nor U2167 (N_2167,N_2150,N_2127);
and U2168 (N_2168,N_2136,N_2125);
and U2169 (N_2169,N_2135,N_2145);
nand U2170 (N_2170,N_2157,N_2122);
nand U2171 (N_2171,N_2114,N_2138);
or U2172 (N_2172,N_2118,N_2113);
and U2173 (N_2173,N_2146,N_2143);
and U2174 (N_2174,N_2149,N_2154);
xor U2175 (N_2175,N_2108,N_2103);
and U2176 (N_2176,N_2156,N_2132);
nand U2177 (N_2177,N_2147,N_2111);
and U2178 (N_2178,N_2129,N_2119);
and U2179 (N_2179,N_2121,N_2112);
xor U2180 (N_2180,N_2100,N_2115);
nand U2181 (N_2181,N_2133,N_2130);
nand U2182 (N_2182,N_2105,N_2131);
or U2183 (N_2183,N_2124,N_2144);
or U2184 (N_2184,N_2152,N_2159);
nor U2185 (N_2185,N_2107,N_2117);
nor U2186 (N_2186,N_2140,N_2106);
and U2187 (N_2187,N_2120,N_2139);
nor U2188 (N_2188,N_2104,N_2155);
and U2189 (N_2189,N_2110,N_2116);
and U2190 (N_2190,N_2138,N_2111);
or U2191 (N_2191,N_2159,N_2156);
nor U2192 (N_2192,N_2123,N_2103);
xnor U2193 (N_2193,N_2142,N_2145);
nand U2194 (N_2194,N_2151,N_2125);
nor U2195 (N_2195,N_2118,N_2107);
or U2196 (N_2196,N_2115,N_2148);
or U2197 (N_2197,N_2102,N_2114);
and U2198 (N_2198,N_2129,N_2134);
and U2199 (N_2199,N_2121,N_2143);
or U2200 (N_2200,N_2124,N_2141);
xnor U2201 (N_2201,N_2108,N_2154);
or U2202 (N_2202,N_2113,N_2117);
xnor U2203 (N_2203,N_2122,N_2132);
nor U2204 (N_2204,N_2101,N_2118);
and U2205 (N_2205,N_2137,N_2101);
nor U2206 (N_2206,N_2109,N_2150);
nand U2207 (N_2207,N_2119,N_2133);
and U2208 (N_2208,N_2127,N_2133);
nand U2209 (N_2209,N_2111,N_2136);
nand U2210 (N_2210,N_2117,N_2105);
or U2211 (N_2211,N_2146,N_2141);
or U2212 (N_2212,N_2113,N_2124);
or U2213 (N_2213,N_2148,N_2151);
nor U2214 (N_2214,N_2101,N_2130);
and U2215 (N_2215,N_2101,N_2140);
nand U2216 (N_2216,N_2127,N_2111);
nor U2217 (N_2217,N_2105,N_2158);
nor U2218 (N_2218,N_2138,N_2113);
nand U2219 (N_2219,N_2106,N_2128);
nor U2220 (N_2220,N_2218,N_2197);
and U2221 (N_2221,N_2192,N_2186);
or U2222 (N_2222,N_2176,N_2168);
nor U2223 (N_2223,N_2215,N_2195);
and U2224 (N_2224,N_2178,N_2219);
or U2225 (N_2225,N_2211,N_2165);
or U2226 (N_2226,N_2191,N_2189);
or U2227 (N_2227,N_2177,N_2194);
or U2228 (N_2228,N_2183,N_2203);
nand U2229 (N_2229,N_2198,N_2217);
and U2230 (N_2230,N_2209,N_2206);
and U2231 (N_2231,N_2210,N_2166);
nor U2232 (N_2232,N_2208,N_2167);
or U2233 (N_2233,N_2164,N_2202);
xor U2234 (N_2234,N_2170,N_2205);
nand U2235 (N_2235,N_2172,N_2182);
and U2236 (N_2236,N_2171,N_2162);
nand U2237 (N_2237,N_2161,N_2173);
and U2238 (N_2238,N_2212,N_2184);
or U2239 (N_2239,N_2188,N_2193);
and U2240 (N_2240,N_2180,N_2196);
and U2241 (N_2241,N_2179,N_2216);
nor U2242 (N_2242,N_2204,N_2163);
nand U2243 (N_2243,N_2207,N_2199);
nor U2244 (N_2244,N_2214,N_2213);
or U2245 (N_2245,N_2181,N_2201);
nand U2246 (N_2246,N_2185,N_2174);
xnor U2247 (N_2247,N_2187,N_2160);
nor U2248 (N_2248,N_2175,N_2169);
nor U2249 (N_2249,N_2200,N_2190);
or U2250 (N_2250,N_2170,N_2160);
and U2251 (N_2251,N_2176,N_2204);
and U2252 (N_2252,N_2203,N_2162);
or U2253 (N_2253,N_2215,N_2217);
nand U2254 (N_2254,N_2191,N_2218);
nor U2255 (N_2255,N_2173,N_2218);
nand U2256 (N_2256,N_2168,N_2191);
and U2257 (N_2257,N_2186,N_2199);
and U2258 (N_2258,N_2207,N_2170);
nand U2259 (N_2259,N_2190,N_2193);
nand U2260 (N_2260,N_2172,N_2183);
nor U2261 (N_2261,N_2192,N_2183);
nand U2262 (N_2262,N_2215,N_2160);
nor U2263 (N_2263,N_2190,N_2173);
nand U2264 (N_2264,N_2193,N_2167);
nor U2265 (N_2265,N_2186,N_2178);
nand U2266 (N_2266,N_2216,N_2173);
or U2267 (N_2267,N_2202,N_2183);
nor U2268 (N_2268,N_2169,N_2213);
nand U2269 (N_2269,N_2197,N_2177);
and U2270 (N_2270,N_2213,N_2171);
nand U2271 (N_2271,N_2169,N_2189);
or U2272 (N_2272,N_2178,N_2163);
and U2273 (N_2273,N_2175,N_2160);
and U2274 (N_2274,N_2204,N_2191);
or U2275 (N_2275,N_2193,N_2179);
nand U2276 (N_2276,N_2181,N_2217);
or U2277 (N_2277,N_2186,N_2176);
nor U2278 (N_2278,N_2214,N_2203);
nand U2279 (N_2279,N_2209,N_2203);
and U2280 (N_2280,N_2223,N_2258);
nor U2281 (N_2281,N_2273,N_2267);
and U2282 (N_2282,N_2276,N_2277);
xor U2283 (N_2283,N_2227,N_2261);
or U2284 (N_2284,N_2249,N_2259);
or U2285 (N_2285,N_2270,N_2236);
or U2286 (N_2286,N_2274,N_2248);
nand U2287 (N_2287,N_2246,N_2265);
or U2288 (N_2288,N_2224,N_2257);
nand U2289 (N_2289,N_2244,N_2275);
nor U2290 (N_2290,N_2243,N_2263);
nand U2291 (N_2291,N_2269,N_2262);
nor U2292 (N_2292,N_2255,N_2245);
nor U2293 (N_2293,N_2252,N_2251);
nor U2294 (N_2294,N_2222,N_2266);
or U2295 (N_2295,N_2225,N_2226);
and U2296 (N_2296,N_2279,N_2231);
and U2297 (N_2297,N_2271,N_2247);
nor U2298 (N_2298,N_2230,N_2229);
or U2299 (N_2299,N_2253,N_2233);
nor U2300 (N_2300,N_2228,N_2278);
nor U2301 (N_2301,N_2268,N_2272);
or U2302 (N_2302,N_2235,N_2250);
or U2303 (N_2303,N_2260,N_2237);
and U2304 (N_2304,N_2256,N_2220);
nor U2305 (N_2305,N_2241,N_2221);
and U2306 (N_2306,N_2239,N_2234);
nor U2307 (N_2307,N_2242,N_2238);
nand U2308 (N_2308,N_2240,N_2264);
nor U2309 (N_2309,N_2254,N_2232);
and U2310 (N_2310,N_2264,N_2248);
nor U2311 (N_2311,N_2236,N_2258);
nor U2312 (N_2312,N_2233,N_2274);
and U2313 (N_2313,N_2264,N_2266);
nand U2314 (N_2314,N_2268,N_2229);
and U2315 (N_2315,N_2267,N_2265);
nor U2316 (N_2316,N_2273,N_2256);
or U2317 (N_2317,N_2262,N_2243);
nand U2318 (N_2318,N_2243,N_2249);
and U2319 (N_2319,N_2236,N_2249);
nor U2320 (N_2320,N_2229,N_2275);
nand U2321 (N_2321,N_2226,N_2252);
and U2322 (N_2322,N_2277,N_2236);
nor U2323 (N_2323,N_2236,N_2265);
nand U2324 (N_2324,N_2260,N_2279);
and U2325 (N_2325,N_2236,N_2228);
nand U2326 (N_2326,N_2266,N_2256);
nand U2327 (N_2327,N_2229,N_2227);
and U2328 (N_2328,N_2257,N_2274);
nor U2329 (N_2329,N_2273,N_2236);
nor U2330 (N_2330,N_2256,N_2225);
or U2331 (N_2331,N_2227,N_2277);
nand U2332 (N_2332,N_2230,N_2221);
nor U2333 (N_2333,N_2230,N_2279);
nand U2334 (N_2334,N_2243,N_2274);
nand U2335 (N_2335,N_2226,N_2266);
and U2336 (N_2336,N_2257,N_2266);
and U2337 (N_2337,N_2268,N_2264);
nand U2338 (N_2338,N_2245,N_2226);
and U2339 (N_2339,N_2273,N_2259);
nand U2340 (N_2340,N_2288,N_2286);
nor U2341 (N_2341,N_2325,N_2301);
or U2342 (N_2342,N_2309,N_2339);
nor U2343 (N_2343,N_2338,N_2317);
or U2344 (N_2344,N_2330,N_2332);
or U2345 (N_2345,N_2335,N_2289);
nand U2346 (N_2346,N_2304,N_2302);
and U2347 (N_2347,N_2298,N_2280);
and U2348 (N_2348,N_2326,N_2336);
xor U2349 (N_2349,N_2331,N_2337);
or U2350 (N_2350,N_2316,N_2311);
nand U2351 (N_2351,N_2283,N_2292);
nor U2352 (N_2352,N_2333,N_2306);
or U2353 (N_2353,N_2297,N_2305);
and U2354 (N_2354,N_2321,N_2285);
or U2355 (N_2355,N_2320,N_2287);
and U2356 (N_2356,N_2314,N_2323);
or U2357 (N_2357,N_2307,N_2290);
and U2358 (N_2358,N_2294,N_2281);
xor U2359 (N_2359,N_2329,N_2322);
and U2360 (N_2360,N_2295,N_2313);
nand U2361 (N_2361,N_2328,N_2303);
nor U2362 (N_2362,N_2315,N_2291);
or U2363 (N_2363,N_2324,N_2293);
nand U2364 (N_2364,N_2296,N_2318);
nor U2365 (N_2365,N_2284,N_2312);
nor U2366 (N_2366,N_2282,N_2308);
or U2367 (N_2367,N_2319,N_2334);
nor U2368 (N_2368,N_2327,N_2310);
and U2369 (N_2369,N_2299,N_2300);
and U2370 (N_2370,N_2339,N_2287);
or U2371 (N_2371,N_2322,N_2291);
nand U2372 (N_2372,N_2288,N_2306);
nor U2373 (N_2373,N_2297,N_2301);
or U2374 (N_2374,N_2327,N_2286);
nor U2375 (N_2375,N_2338,N_2334);
nor U2376 (N_2376,N_2314,N_2313);
and U2377 (N_2377,N_2305,N_2339);
nand U2378 (N_2378,N_2289,N_2290);
nor U2379 (N_2379,N_2318,N_2339);
or U2380 (N_2380,N_2281,N_2337);
nand U2381 (N_2381,N_2315,N_2280);
nor U2382 (N_2382,N_2328,N_2316);
or U2383 (N_2383,N_2323,N_2318);
or U2384 (N_2384,N_2331,N_2289);
xor U2385 (N_2385,N_2301,N_2324);
nor U2386 (N_2386,N_2296,N_2289);
nor U2387 (N_2387,N_2290,N_2300);
and U2388 (N_2388,N_2312,N_2291);
nand U2389 (N_2389,N_2301,N_2290);
nor U2390 (N_2390,N_2282,N_2336);
or U2391 (N_2391,N_2303,N_2304);
nand U2392 (N_2392,N_2338,N_2320);
or U2393 (N_2393,N_2324,N_2320);
nor U2394 (N_2394,N_2325,N_2306);
or U2395 (N_2395,N_2314,N_2334);
nand U2396 (N_2396,N_2313,N_2305);
nand U2397 (N_2397,N_2335,N_2288);
or U2398 (N_2398,N_2330,N_2303);
nand U2399 (N_2399,N_2301,N_2310);
nand U2400 (N_2400,N_2398,N_2391);
nor U2401 (N_2401,N_2373,N_2384);
nor U2402 (N_2402,N_2377,N_2366);
and U2403 (N_2403,N_2362,N_2363);
xor U2404 (N_2404,N_2370,N_2346);
and U2405 (N_2405,N_2395,N_2347);
or U2406 (N_2406,N_2396,N_2358);
nand U2407 (N_2407,N_2368,N_2367);
nand U2408 (N_2408,N_2399,N_2382);
and U2409 (N_2409,N_2387,N_2350);
nand U2410 (N_2410,N_2374,N_2351);
nand U2411 (N_2411,N_2383,N_2380);
or U2412 (N_2412,N_2371,N_2356);
nor U2413 (N_2413,N_2361,N_2360);
xor U2414 (N_2414,N_2340,N_2390);
nand U2415 (N_2415,N_2365,N_2389);
nor U2416 (N_2416,N_2386,N_2369);
or U2417 (N_2417,N_2375,N_2354);
and U2418 (N_2418,N_2343,N_2379);
xnor U2419 (N_2419,N_2353,N_2345);
nor U2420 (N_2420,N_2372,N_2348);
or U2421 (N_2421,N_2394,N_2359);
nand U2422 (N_2422,N_2393,N_2364);
nand U2423 (N_2423,N_2392,N_2378);
or U2424 (N_2424,N_2352,N_2342);
nor U2425 (N_2425,N_2341,N_2397);
nor U2426 (N_2426,N_2355,N_2349);
or U2427 (N_2427,N_2381,N_2344);
nor U2428 (N_2428,N_2388,N_2376);
and U2429 (N_2429,N_2385,N_2357);
nor U2430 (N_2430,N_2358,N_2341);
and U2431 (N_2431,N_2382,N_2358);
and U2432 (N_2432,N_2393,N_2365);
nor U2433 (N_2433,N_2397,N_2346);
and U2434 (N_2434,N_2385,N_2362);
and U2435 (N_2435,N_2397,N_2387);
or U2436 (N_2436,N_2364,N_2353);
or U2437 (N_2437,N_2347,N_2357);
nand U2438 (N_2438,N_2380,N_2381);
nand U2439 (N_2439,N_2389,N_2395);
and U2440 (N_2440,N_2383,N_2363);
nand U2441 (N_2441,N_2358,N_2340);
and U2442 (N_2442,N_2354,N_2344);
nand U2443 (N_2443,N_2349,N_2391);
nor U2444 (N_2444,N_2343,N_2355);
nor U2445 (N_2445,N_2393,N_2380);
nand U2446 (N_2446,N_2394,N_2355);
nand U2447 (N_2447,N_2340,N_2373);
nor U2448 (N_2448,N_2382,N_2376);
nor U2449 (N_2449,N_2395,N_2388);
and U2450 (N_2450,N_2373,N_2390);
or U2451 (N_2451,N_2341,N_2344);
nor U2452 (N_2452,N_2397,N_2377);
or U2453 (N_2453,N_2352,N_2371);
nand U2454 (N_2454,N_2387,N_2344);
and U2455 (N_2455,N_2378,N_2362);
and U2456 (N_2456,N_2358,N_2399);
nor U2457 (N_2457,N_2382,N_2364);
nand U2458 (N_2458,N_2399,N_2375);
nor U2459 (N_2459,N_2387,N_2343);
or U2460 (N_2460,N_2418,N_2408);
and U2461 (N_2461,N_2452,N_2413);
and U2462 (N_2462,N_2431,N_2441);
and U2463 (N_2463,N_2459,N_2407);
nor U2464 (N_2464,N_2430,N_2426);
or U2465 (N_2465,N_2410,N_2438);
or U2466 (N_2466,N_2414,N_2437);
nand U2467 (N_2467,N_2435,N_2428);
nor U2468 (N_2468,N_2444,N_2447);
nand U2469 (N_2469,N_2457,N_2450);
nor U2470 (N_2470,N_2419,N_2446);
or U2471 (N_2471,N_2432,N_2443);
or U2472 (N_2472,N_2400,N_2412);
nor U2473 (N_2473,N_2453,N_2458);
and U2474 (N_2474,N_2405,N_2422);
nand U2475 (N_2475,N_2449,N_2406);
nor U2476 (N_2476,N_2424,N_2436);
nor U2477 (N_2477,N_2403,N_2425);
and U2478 (N_2478,N_2439,N_2429);
and U2479 (N_2479,N_2451,N_2433);
and U2480 (N_2480,N_2416,N_2415);
nand U2481 (N_2481,N_2445,N_2434);
and U2482 (N_2482,N_2454,N_2417);
or U2483 (N_2483,N_2401,N_2442);
nand U2484 (N_2484,N_2402,N_2448);
and U2485 (N_2485,N_2455,N_2456);
and U2486 (N_2486,N_2427,N_2411);
or U2487 (N_2487,N_2404,N_2440);
and U2488 (N_2488,N_2409,N_2423);
nor U2489 (N_2489,N_2420,N_2421);
or U2490 (N_2490,N_2422,N_2428);
or U2491 (N_2491,N_2427,N_2452);
nand U2492 (N_2492,N_2420,N_2440);
nand U2493 (N_2493,N_2417,N_2435);
nor U2494 (N_2494,N_2409,N_2415);
or U2495 (N_2495,N_2457,N_2422);
and U2496 (N_2496,N_2425,N_2412);
nor U2497 (N_2497,N_2457,N_2410);
or U2498 (N_2498,N_2405,N_2444);
xnor U2499 (N_2499,N_2406,N_2409);
nor U2500 (N_2500,N_2412,N_2402);
and U2501 (N_2501,N_2406,N_2430);
nor U2502 (N_2502,N_2405,N_2407);
nand U2503 (N_2503,N_2417,N_2447);
and U2504 (N_2504,N_2400,N_2441);
and U2505 (N_2505,N_2423,N_2433);
nor U2506 (N_2506,N_2426,N_2459);
and U2507 (N_2507,N_2405,N_2453);
nand U2508 (N_2508,N_2443,N_2444);
nand U2509 (N_2509,N_2430,N_2417);
and U2510 (N_2510,N_2443,N_2436);
or U2511 (N_2511,N_2426,N_2423);
and U2512 (N_2512,N_2408,N_2419);
and U2513 (N_2513,N_2457,N_2403);
nand U2514 (N_2514,N_2432,N_2411);
or U2515 (N_2515,N_2417,N_2429);
and U2516 (N_2516,N_2410,N_2446);
nor U2517 (N_2517,N_2416,N_2449);
nand U2518 (N_2518,N_2403,N_2419);
nand U2519 (N_2519,N_2438,N_2420);
nor U2520 (N_2520,N_2489,N_2509);
and U2521 (N_2521,N_2484,N_2470);
nand U2522 (N_2522,N_2500,N_2467);
nand U2523 (N_2523,N_2517,N_2497);
nor U2524 (N_2524,N_2487,N_2519);
nand U2525 (N_2525,N_2512,N_2478);
and U2526 (N_2526,N_2515,N_2506);
or U2527 (N_2527,N_2511,N_2460);
and U2528 (N_2528,N_2462,N_2516);
and U2529 (N_2529,N_2491,N_2471);
and U2530 (N_2530,N_2501,N_2488);
nand U2531 (N_2531,N_2496,N_2464);
nand U2532 (N_2532,N_2499,N_2510);
and U2533 (N_2533,N_2508,N_2474);
nor U2534 (N_2534,N_2472,N_2503);
nor U2535 (N_2535,N_2514,N_2493);
nand U2536 (N_2536,N_2498,N_2492);
and U2537 (N_2537,N_2473,N_2494);
or U2538 (N_2538,N_2518,N_2466);
and U2539 (N_2539,N_2486,N_2469);
or U2540 (N_2540,N_2463,N_2465);
nand U2541 (N_2541,N_2495,N_2479);
and U2542 (N_2542,N_2505,N_2502);
nor U2543 (N_2543,N_2461,N_2504);
nand U2544 (N_2544,N_2490,N_2468);
or U2545 (N_2545,N_2507,N_2513);
nand U2546 (N_2546,N_2482,N_2485);
nor U2547 (N_2547,N_2476,N_2481);
nor U2548 (N_2548,N_2480,N_2477);
nand U2549 (N_2549,N_2483,N_2475);
nand U2550 (N_2550,N_2462,N_2495);
nand U2551 (N_2551,N_2504,N_2515);
or U2552 (N_2552,N_2494,N_2517);
xor U2553 (N_2553,N_2475,N_2479);
and U2554 (N_2554,N_2460,N_2461);
and U2555 (N_2555,N_2493,N_2503);
nand U2556 (N_2556,N_2478,N_2491);
or U2557 (N_2557,N_2467,N_2493);
nor U2558 (N_2558,N_2519,N_2490);
and U2559 (N_2559,N_2489,N_2494);
or U2560 (N_2560,N_2470,N_2471);
nor U2561 (N_2561,N_2513,N_2476);
and U2562 (N_2562,N_2494,N_2475);
nor U2563 (N_2563,N_2512,N_2488);
or U2564 (N_2564,N_2487,N_2460);
nor U2565 (N_2565,N_2511,N_2476);
nor U2566 (N_2566,N_2478,N_2516);
nand U2567 (N_2567,N_2472,N_2479);
nor U2568 (N_2568,N_2518,N_2514);
nand U2569 (N_2569,N_2500,N_2462);
nor U2570 (N_2570,N_2505,N_2471);
or U2571 (N_2571,N_2466,N_2484);
or U2572 (N_2572,N_2487,N_2483);
or U2573 (N_2573,N_2487,N_2500);
and U2574 (N_2574,N_2467,N_2519);
nor U2575 (N_2575,N_2492,N_2511);
nor U2576 (N_2576,N_2460,N_2472);
nand U2577 (N_2577,N_2480,N_2519);
nand U2578 (N_2578,N_2499,N_2498);
nor U2579 (N_2579,N_2493,N_2504);
nor U2580 (N_2580,N_2537,N_2568);
nor U2581 (N_2581,N_2565,N_2564);
and U2582 (N_2582,N_2530,N_2557);
nand U2583 (N_2583,N_2524,N_2521);
and U2584 (N_2584,N_2563,N_2548);
or U2585 (N_2585,N_2578,N_2570);
and U2586 (N_2586,N_2544,N_2571);
nor U2587 (N_2587,N_2527,N_2573);
or U2588 (N_2588,N_2555,N_2535);
nand U2589 (N_2589,N_2534,N_2556);
xnor U2590 (N_2590,N_2558,N_2561);
or U2591 (N_2591,N_2545,N_2550);
or U2592 (N_2592,N_2538,N_2575);
nand U2593 (N_2593,N_2525,N_2522);
or U2594 (N_2594,N_2569,N_2540);
or U2595 (N_2595,N_2546,N_2523);
and U2596 (N_2596,N_2539,N_2528);
nand U2597 (N_2597,N_2552,N_2566);
nand U2598 (N_2598,N_2559,N_2531);
or U2599 (N_2599,N_2562,N_2560);
and U2600 (N_2600,N_2572,N_2520);
nor U2601 (N_2601,N_2551,N_2579);
nand U2602 (N_2602,N_2532,N_2526);
nor U2603 (N_2603,N_2542,N_2536);
xnor U2604 (N_2604,N_2554,N_2543);
nand U2605 (N_2605,N_2576,N_2529);
and U2606 (N_2606,N_2567,N_2549);
or U2607 (N_2607,N_2533,N_2553);
nor U2608 (N_2608,N_2541,N_2577);
or U2609 (N_2609,N_2574,N_2547);
nand U2610 (N_2610,N_2565,N_2575);
nand U2611 (N_2611,N_2576,N_2546);
nor U2612 (N_2612,N_2535,N_2540);
or U2613 (N_2613,N_2529,N_2553);
and U2614 (N_2614,N_2538,N_2522);
nand U2615 (N_2615,N_2571,N_2554);
nand U2616 (N_2616,N_2547,N_2536);
nor U2617 (N_2617,N_2549,N_2535);
nand U2618 (N_2618,N_2548,N_2579);
and U2619 (N_2619,N_2557,N_2533);
nor U2620 (N_2620,N_2566,N_2558);
xor U2621 (N_2621,N_2573,N_2547);
nor U2622 (N_2622,N_2527,N_2550);
or U2623 (N_2623,N_2545,N_2577);
nand U2624 (N_2624,N_2529,N_2544);
and U2625 (N_2625,N_2541,N_2547);
nor U2626 (N_2626,N_2579,N_2535);
and U2627 (N_2627,N_2571,N_2528);
nand U2628 (N_2628,N_2575,N_2551);
nand U2629 (N_2629,N_2551,N_2560);
nand U2630 (N_2630,N_2556,N_2527);
or U2631 (N_2631,N_2576,N_2568);
and U2632 (N_2632,N_2530,N_2577);
nand U2633 (N_2633,N_2521,N_2522);
and U2634 (N_2634,N_2566,N_2573);
and U2635 (N_2635,N_2566,N_2553);
or U2636 (N_2636,N_2578,N_2546);
nor U2637 (N_2637,N_2524,N_2558);
or U2638 (N_2638,N_2547,N_2523);
nor U2639 (N_2639,N_2574,N_2531);
nand U2640 (N_2640,N_2605,N_2603);
nor U2641 (N_2641,N_2638,N_2610);
nand U2642 (N_2642,N_2593,N_2587);
or U2643 (N_2643,N_2596,N_2584);
nand U2644 (N_2644,N_2619,N_2598);
nand U2645 (N_2645,N_2630,N_2583);
and U2646 (N_2646,N_2607,N_2623);
nand U2647 (N_2647,N_2606,N_2621);
and U2648 (N_2648,N_2594,N_2586);
and U2649 (N_2649,N_2613,N_2588);
xor U2650 (N_2650,N_2626,N_2614);
nand U2651 (N_2651,N_2634,N_2612);
and U2652 (N_2652,N_2618,N_2635);
or U2653 (N_2653,N_2595,N_2633);
and U2654 (N_2654,N_2625,N_2636);
and U2655 (N_2655,N_2589,N_2604);
nand U2656 (N_2656,N_2608,N_2609);
nand U2657 (N_2657,N_2600,N_2632);
nand U2658 (N_2658,N_2631,N_2611);
nor U2659 (N_2659,N_2615,N_2616);
nor U2660 (N_2660,N_2590,N_2602);
nand U2661 (N_2661,N_2592,N_2585);
nand U2662 (N_2662,N_2617,N_2624);
or U2663 (N_2663,N_2627,N_2582);
and U2664 (N_2664,N_2597,N_2580);
or U2665 (N_2665,N_2581,N_2637);
and U2666 (N_2666,N_2639,N_2628);
or U2667 (N_2667,N_2591,N_2599);
nor U2668 (N_2668,N_2629,N_2622);
and U2669 (N_2669,N_2620,N_2601);
or U2670 (N_2670,N_2611,N_2587);
nand U2671 (N_2671,N_2584,N_2580);
or U2672 (N_2672,N_2609,N_2591);
and U2673 (N_2673,N_2612,N_2623);
nor U2674 (N_2674,N_2629,N_2583);
or U2675 (N_2675,N_2616,N_2603);
nand U2676 (N_2676,N_2605,N_2586);
nand U2677 (N_2677,N_2581,N_2629);
or U2678 (N_2678,N_2637,N_2621);
nor U2679 (N_2679,N_2587,N_2580);
nor U2680 (N_2680,N_2582,N_2632);
and U2681 (N_2681,N_2615,N_2637);
nor U2682 (N_2682,N_2617,N_2595);
and U2683 (N_2683,N_2618,N_2617);
and U2684 (N_2684,N_2623,N_2630);
nand U2685 (N_2685,N_2600,N_2617);
nand U2686 (N_2686,N_2613,N_2602);
or U2687 (N_2687,N_2616,N_2635);
and U2688 (N_2688,N_2580,N_2628);
and U2689 (N_2689,N_2595,N_2601);
or U2690 (N_2690,N_2628,N_2595);
or U2691 (N_2691,N_2587,N_2583);
or U2692 (N_2692,N_2620,N_2618);
nor U2693 (N_2693,N_2602,N_2580);
and U2694 (N_2694,N_2626,N_2619);
and U2695 (N_2695,N_2600,N_2606);
nand U2696 (N_2696,N_2582,N_2585);
nand U2697 (N_2697,N_2623,N_2589);
and U2698 (N_2698,N_2627,N_2626);
and U2699 (N_2699,N_2615,N_2601);
and U2700 (N_2700,N_2668,N_2666);
or U2701 (N_2701,N_2694,N_2654);
and U2702 (N_2702,N_2656,N_2676);
nand U2703 (N_2703,N_2646,N_2660);
or U2704 (N_2704,N_2661,N_2653);
nor U2705 (N_2705,N_2674,N_2672);
nand U2706 (N_2706,N_2669,N_2687);
and U2707 (N_2707,N_2698,N_2695);
or U2708 (N_2708,N_2682,N_2640);
nor U2709 (N_2709,N_2658,N_2697);
nor U2710 (N_2710,N_2696,N_2648);
nand U2711 (N_2711,N_2689,N_2699);
and U2712 (N_2712,N_2684,N_2691);
nor U2713 (N_2713,N_2652,N_2663);
and U2714 (N_2714,N_2657,N_2651);
nand U2715 (N_2715,N_2680,N_2673);
nand U2716 (N_2716,N_2692,N_2679);
and U2717 (N_2717,N_2665,N_2675);
nor U2718 (N_2718,N_2664,N_2683);
or U2719 (N_2719,N_2681,N_2650);
xor U2720 (N_2720,N_2686,N_2647);
or U2721 (N_2721,N_2671,N_2655);
nand U2722 (N_2722,N_2662,N_2677);
nor U2723 (N_2723,N_2641,N_2645);
or U2724 (N_2724,N_2678,N_2688);
nand U2725 (N_2725,N_2670,N_2693);
nand U2726 (N_2726,N_2649,N_2643);
or U2727 (N_2727,N_2685,N_2659);
or U2728 (N_2728,N_2690,N_2667);
or U2729 (N_2729,N_2644,N_2642);
nand U2730 (N_2730,N_2690,N_2661);
nor U2731 (N_2731,N_2690,N_2650);
or U2732 (N_2732,N_2644,N_2676);
xor U2733 (N_2733,N_2689,N_2661);
or U2734 (N_2734,N_2687,N_2655);
xor U2735 (N_2735,N_2683,N_2665);
nand U2736 (N_2736,N_2665,N_2693);
or U2737 (N_2737,N_2679,N_2652);
nand U2738 (N_2738,N_2690,N_2654);
or U2739 (N_2739,N_2680,N_2684);
or U2740 (N_2740,N_2671,N_2642);
nand U2741 (N_2741,N_2641,N_2669);
or U2742 (N_2742,N_2648,N_2651);
nor U2743 (N_2743,N_2696,N_2665);
nand U2744 (N_2744,N_2675,N_2640);
nand U2745 (N_2745,N_2663,N_2651);
nor U2746 (N_2746,N_2691,N_2697);
and U2747 (N_2747,N_2677,N_2654);
nor U2748 (N_2748,N_2657,N_2664);
or U2749 (N_2749,N_2676,N_2669);
and U2750 (N_2750,N_2667,N_2650);
nand U2751 (N_2751,N_2654,N_2693);
nand U2752 (N_2752,N_2641,N_2685);
and U2753 (N_2753,N_2689,N_2664);
nor U2754 (N_2754,N_2668,N_2684);
and U2755 (N_2755,N_2651,N_2649);
or U2756 (N_2756,N_2694,N_2650);
nand U2757 (N_2757,N_2696,N_2698);
and U2758 (N_2758,N_2672,N_2693);
nor U2759 (N_2759,N_2659,N_2697);
nor U2760 (N_2760,N_2756,N_2755);
nor U2761 (N_2761,N_2724,N_2717);
or U2762 (N_2762,N_2752,N_2703);
and U2763 (N_2763,N_2749,N_2741);
nand U2764 (N_2764,N_2757,N_2747);
and U2765 (N_2765,N_2715,N_2745);
nor U2766 (N_2766,N_2750,N_2729);
and U2767 (N_2767,N_2744,N_2710);
nor U2768 (N_2768,N_2738,N_2707);
and U2769 (N_2769,N_2702,N_2725);
nand U2770 (N_2770,N_2728,N_2742);
nor U2771 (N_2771,N_2705,N_2706);
or U2772 (N_2772,N_2721,N_2740);
nor U2773 (N_2773,N_2758,N_2746);
and U2774 (N_2774,N_2712,N_2700);
and U2775 (N_2775,N_2734,N_2730);
nor U2776 (N_2776,N_2714,N_2720);
xor U2777 (N_2777,N_2722,N_2704);
nand U2778 (N_2778,N_2713,N_2733);
nor U2779 (N_2779,N_2735,N_2726);
nor U2780 (N_2780,N_2711,N_2737);
and U2781 (N_2781,N_2719,N_2723);
nor U2782 (N_2782,N_2716,N_2718);
nor U2783 (N_2783,N_2759,N_2701);
nor U2784 (N_2784,N_2748,N_2751);
or U2785 (N_2785,N_2736,N_2731);
nor U2786 (N_2786,N_2709,N_2727);
xnor U2787 (N_2787,N_2753,N_2739);
nor U2788 (N_2788,N_2708,N_2754);
xor U2789 (N_2789,N_2732,N_2743);
nand U2790 (N_2790,N_2726,N_2723);
nor U2791 (N_2791,N_2703,N_2704);
and U2792 (N_2792,N_2710,N_2709);
xnor U2793 (N_2793,N_2747,N_2730);
and U2794 (N_2794,N_2718,N_2703);
or U2795 (N_2795,N_2714,N_2732);
and U2796 (N_2796,N_2706,N_2717);
and U2797 (N_2797,N_2718,N_2722);
or U2798 (N_2798,N_2710,N_2747);
or U2799 (N_2799,N_2751,N_2755);
nor U2800 (N_2800,N_2756,N_2748);
nor U2801 (N_2801,N_2705,N_2715);
or U2802 (N_2802,N_2727,N_2734);
nand U2803 (N_2803,N_2756,N_2734);
nor U2804 (N_2804,N_2722,N_2701);
nor U2805 (N_2805,N_2751,N_2720);
and U2806 (N_2806,N_2739,N_2758);
nand U2807 (N_2807,N_2758,N_2716);
nor U2808 (N_2808,N_2752,N_2712);
nand U2809 (N_2809,N_2709,N_2717);
nand U2810 (N_2810,N_2719,N_2717);
nand U2811 (N_2811,N_2744,N_2757);
nor U2812 (N_2812,N_2707,N_2758);
or U2813 (N_2813,N_2752,N_2704);
nor U2814 (N_2814,N_2735,N_2751);
xor U2815 (N_2815,N_2737,N_2746);
and U2816 (N_2816,N_2721,N_2730);
or U2817 (N_2817,N_2701,N_2735);
nand U2818 (N_2818,N_2737,N_2732);
nand U2819 (N_2819,N_2735,N_2740);
nand U2820 (N_2820,N_2804,N_2817);
and U2821 (N_2821,N_2818,N_2794);
or U2822 (N_2822,N_2775,N_2776);
nand U2823 (N_2823,N_2796,N_2810);
or U2824 (N_2824,N_2764,N_2819);
and U2825 (N_2825,N_2799,N_2781);
and U2826 (N_2826,N_2768,N_2790);
nor U2827 (N_2827,N_2770,N_2761);
nand U2828 (N_2828,N_2783,N_2809);
nand U2829 (N_2829,N_2782,N_2798);
and U2830 (N_2830,N_2784,N_2773);
or U2831 (N_2831,N_2786,N_2785);
nor U2832 (N_2832,N_2779,N_2772);
nor U2833 (N_2833,N_2812,N_2793);
and U2834 (N_2834,N_2771,N_2797);
nand U2835 (N_2835,N_2800,N_2760);
or U2836 (N_2836,N_2791,N_2805);
xnor U2837 (N_2837,N_2765,N_2763);
nand U2838 (N_2838,N_2816,N_2807);
or U2839 (N_2839,N_2789,N_2778);
and U2840 (N_2840,N_2780,N_2815);
xnor U2841 (N_2841,N_2811,N_2801);
and U2842 (N_2842,N_2766,N_2767);
and U2843 (N_2843,N_2795,N_2806);
or U2844 (N_2844,N_2803,N_2774);
and U2845 (N_2845,N_2777,N_2808);
xnor U2846 (N_2846,N_2813,N_2802);
or U2847 (N_2847,N_2769,N_2787);
and U2848 (N_2848,N_2814,N_2762);
nor U2849 (N_2849,N_2792,N_2788);
nand U2850 (N_2850,N_2794,N_2762);
nor U2851 (N_2851,N_2789,N_2793);
nor U2852 (N_2852,N_2781,N_2766);
or U2853 (N_2853,N_2810,N_2814);
nand U2854 (N_2854,N_2806,N_2788);
and U2855 (N_2855,N_2762,N_2813);
and U2856 (N_2856,N_2809,N_2779);
nand U2857 (N_2857,N_2763,N_2807);
and U2858 (N_2858,N_2776,N_2766);
nand U2859 (N_2859,N_2803,N_2762);
and U2860 (N_2860,N_2810,N_2764);
or U2861 (N_2861,N_2803,N_2777);
or U2862 (N_2862,N_2783,N_2796);
nand U2863 (N_2863,N_2764,N_2775);
nand U2864 (N_2864,N_2761,N_2790);
or U2865 (N_2865,N_2772,N_2769);
nor U2866 (N_2866,N_2813,N_2788);
nand U2867 (N_2867,N_2771,N_2791);
nand U2868 (N_2868,N_2819,N_2791);
nand U2869 (N_2869,N_2771,N_2768);
or U2870 (N_2870,N_2798,N_2816);
nand U2871 (N_2871,N_2777,N_2763);
and U2872 (N_2872,N_2805,N_2766);
or U2873 (N_2873,N_2765,N_2798);
or U2874 (N_2874,N_2807,N_2784);
or U2875 (N_2875,N_2795,N_2774);
nor U2876 (N_2876,N_2802,N_2792);
nand U2877 (N_2877,N_2779,N_2767);
or U2878 (N_2878,N_2762,N_2810);
or U2879 (N_2879,N_2801,N_2768);
nor U2880 (N_2880,N_2866,N_2851);
nand U2881 (N_2881,N_2841,N_2860);
nor U2882 (N_2882,N_2856,N_2847);
nor U2883 (N_2883,N_2850,N_2821);
nor U2884 (N_2884,N_2824,N_2835);
or U2885 (N_2885,N_2868,N_2855);
or U2886 (N_2886,N_2874,N_2837);
nand U2887 (N_2887,N_2834,N_2867);
and U2888 (N_2888,N_2873,N_2829);
or U2889 (N_2889,N_2823,N_2869);
or U2890 (N_2890,N_2848,N_2859);
and U2891 (N_2891,N_2875,N_2822);
or U2892 (N_2892,N_2836,N_2830);
nand U2893 (N_2893,N_2877,N_2854);
and U2894 (N_2894,N_2828,N_2827);
or U2895 (N_2895,N_2870,N_2826);
and U2896 (N_2896,N_2864,N_2820);
nor U2897 (N_2897,N_2853,N_2840);
or U2898 (N_2898,N_2876,N_2831);
and U2899 (N_2899,N_2865,N_2852);
nand U2900 (N_2900,N_2871,N_2842);
and U2901 (N_2901,N_2838,N_2849);
and U2902 (N_2902,N_2839,N_2872);
or U2903 (N_2903,N_2832,N_2843);
and U2904 (N_2904,N_2857,N_2845);
or U2905 (N_2905,N_2833,N_2862);
nand U2906 (N_2906,N_2878,N_2846);
or U2907 (N_2907,N_2861,N_2879);
nand U2908 (N_2908,N_2825,N_2844);
nor U2909 (N_2909,N_2858,N_2863);
nand U2910 (N_2910,N_2868,N_2858);
or U2911 (N_2911,N_2876,N_2874);
or U2912 (N_2912,N_2820,N_2821);
or U2913 (N_2913,N_2858,N_2836);
xnor U2914 (N_2914,N_2865,N_2866);
nor U2915 (N_2915,N_2861,N_2855);
nor U2916 (N_2916,N_2843,N_2857);
nand U2917 (N_2917,N_2848,N_2831);
nand U2918 (N_2918,N_2840,N_2830);
or U2919 (N_2919,N_2869,N_2848);
nand U2920 (N_2920,N_2867,N_2846);
nor U2921 (N_2921,N_2869,N_2856);
or U2922 (N_2922,N_2879,N_2847);
nor U2923 (N_2923,N_2836,N_2853);
nor U2924 (N_2924,N_2832,N_2834);
or U2925 (N_2925,N_2861,N_2853);
nand U2926 (N_2926,N_2867,N_2850);
or U2927 (N_2927,N_2851,N_2848);
and U2928 (N_2928,N_2863,N_2840);
or U2929 (N_2929,N_2828,N_2821);
nand U2930 (N_2930,N_2829,N_2831);
nand U2931 (N_2931,N_2866,N_2834);
and U2932 (N_2932,N_2823,N_2862);
nand U2933 (N_2933,N_2839,N_2823);
or U2934 (N_2934,N_2862,N_2855);
and U2935 (N_2935,N_2853,N_2868);
or U2936 (N_2936,N_2855,N_2846);
nand U2937 (N_2937,N_2842,N_2821);
nand U2938 (N_2938,N_2840,N_2824);
and U2939 (N_2939,N_2877,N_2863);
or U2940 (N_2940,N_2926,N_2920);
nor U2941 (N_2941,N_2909,N_2897);
or U2942 (N_2942,N_2913,N_2902);
and U2943 (N_2943,N_2923,N_2890);
nand U2944 (N_2944,N_2894,N_2887);
nor U2945 (N_2945,N_2892,N_2921);
and U2946 (N_2946,N_2881,N_2932);
or U2947 (N_2947,N_2937,N_2912);
or U2948 (N_2948,N_2899,N_2882);
or U2949 (N_2949,N_2934,N_2901);
nand U2950 (N_2950,N_2930,N_2918);
nor U2951 (N_2951,N_2910,N_2922);
or U2952 (N_2952,N_2907,N_2935);
nor U2953 (N_2953,N_2886,N_2900);
nor U2954 (N_2954,N_2919,N_2938);
and U2955 (N_2955,N_2925,N_2895);
and U2956 (N_2956,N_2884,N_2927);
nand U2957 (N_2957,N_2905,N_2914);
nand U2958 (N_2958,N_2916,N_2893);
and U2959 (N_2959,N_2936,N_2889);
nand U2960 (N_2960,N_2898,N_2880);
nand U2961 (N_2961,N_2931,N_2928);
nand U2962 (N_2962,N_2906,N_2915);
nor U2963 (N_2963,N_2929,N_2904);
and U2964 (N_2964,N_2888,N_2939);
nor U2965 (N_2965,N_2883,N_2891);
nand U2966 (N_2966,N_2911,N_2933);
or U2967 (N_2967,N_2885,N_2903);
and U2968 (N_2968,N_2896,N_2917);
and U2969 (N_2969,N_2924,N_2908);
nand U2970 (N_2970,N_2935,N_2916);
nand U2971 (N_2971,N_2897,N_2917);
nor U2972 (N_2972,N_2939,N_2902);
or U2973 (N_2973,N_2918,N_2905);
and U2974 (N_2974,N_2939,N_2935);
or U2975 (N_2975,N_2896,N_2912);
and U2976 (N_2976,N_2890,N_2932);
nor U2977 (N_2977,N_2925,N_2894);
or U2978 (N_2978,N_2911,N_2885);
and U2979 (N_2979,N_2907,N_2897);
nor U2980 (N_2980,N_2902,N_2938);
nor U2981 (N_2981,N_2914,N_2927);
and U2982 (N_2982,N_2916,N_2930);
or U2983 (N_2983,N_2918,N_2892);
nand U2984 (N_2984,N_2902,N_2894);
and U2985 (N_2985,N_2887,N_2890);
nand U2986 (N_2986,N_2917,N_2889);
nor U2987 (N_2987,N_2902,N_2921);
nor U2988 (N_2988,N_2909,N_2882);
and U2989 (N_2989,N_2915,N_2913);
nor U2990 (N_2990,N_2926,N_2888);
and U2991 (N_2991,N_2893,N_2918);
nand U2992 (N_2992,N_2935,N_2936);
and U2993 (N_2993,N_2898,N_2924);
nand U2994 (N_2994,N_2910,N_2917);
nand U2995 (N_2995,N_2926,N_2934);
or U2996 (N_2996,N_2886,N_2927);
xor U2997 (N_2997,N_2899,N_2897);
nand U2998 (N_2998,N_2901,N_2895);
or U2999 (N_2999,N_2893,N_2931);
nor UO_0 (O_0,N_2976,N_2975);
and UO_1 (O_1,N_2974,N_2988);
or UO_2 (O_2,N_2968,N_2959);
nor UO_3 (O_3,N_2950,N_2999);
nand UO_4 (O_4,N_2971,N_2982);
or UO_5 (O_5,N_2996,N_2964);
and UO_6 (O_6,N_2993,N_2987);
nor UO_7 (O_7,N_2990,N_2981);
and UO_8 (O_8,N_2957,N_2953);
and UO_9 (O_9,N_2942,N_2958);
nor UO_10 (O_10,N_2970,N_2969);
nand UO_11 (O_11,N_2956,N_2949);
nor UO_12 (O_12,N_2946,N_2985);
and UO_13 (O_13,N_2992,N_2947);
and UO_14 (O_14,N_2997,N_2995);
or UO_15 (O_15,N_2944,N_2967);
nor UO_16 (O_16,N_2998,N_2940);
nor UO_17 (O_17,N_2943,N_2960);
nor UO_18 (O_18,N_2965,N_2952);
xor UO_19 (O_19,N_2973,N_2979);
nor UO_20 (O_20,N_2991,N_2972);
nand UO_21 (O_21,N_2955,N_2989);
nor UO_22 (O_22,N_2951,N_2961);
nand UO_23 (O_23,N_2966,N_2978);
xnor UO_24 (O_24,N_2948,N_2954);
nor UO_25 (O_25,N_2963,N_2994);
or UO_26 (O_26,N_2984,N_2941);
and UO_27 (O_27,N_2962,N_2983);
nand UO_28 (O_28,N_2945,N_2986);
nor UO_29 (O_29,N_2977,N_2980);
nor UO_30 (O_30,N_2949,N_2978);
nand UO_31 (O_31,N_2974,N_2986);
nand UO_32 (O_32,N_2980,N_2974);
and UO_33 (O_33,N_2941,N_2978);
xnor UO_34 (O_34,N_2984,N_2947);
or UO_35 (O_35,N_2950,N_2965);
nor UO_36 (O_36,N_2984,N_2976);
or UO_37 (O_37,N_2985,N_2995);
nor UO_38 (O_38,N_2981,N_2995);
or UO_39 (O_39,N_2947,N_2967);
and UO_40 (O_40,N_2968,N_2961);
and UO_41 (O_41,N_2946,N_2997);
and UO_42 (O_42,N_2978,N_2943);
and UO_43 (O_43,N_2998,N_2992);
and UO_44 (O_44,N_2983,N_2946);
and UO_45 (O_45,N_2955,N_2963);
or UO_46 (O_46,N_2984,N_2944);
nor UO_47 (O_47,N_2943,N_2950);
nor UO_48 (O_48,N_2959,N_2955);
xor UO_49 (O_49,N_2945,N_2952);
and UO_50 (O_50,N_2970,N_2946);
or UO_51 (O_51,N_2951,N_2965);
and UO_52 (O_52,N_2978,N_2971);
or UO_53 (O_53,N_2962,N_2991);
or UO_54 (O_54,N_2985,N_2958);
nor UO_55 (O_55,N_2997,N_2949);
nand UO_56 (O_56,N_2993,N_2957);
or UO_57 (O_57,N_2960,N_2982);
nor UO_58 (O_58,N_2998,N_2951);
and UO_59 (O_59,N_2997,N_2975);
nor UO_60 (O_60,N_2940,N_2988);
nand UO_61 (O_61,N_2973,N_2948);
and UO_62 (O_62,N_2990,N_2984);
nor UO_63 (O_63,N_2943,N_2966);
xor UO_64 (O_64,N_2951,N_2945);
and UO_65 (O_65,N_2962,N_2955);
xor UO_66 (O_66,N_2962,N_2984);
or UO_67 (O_67,N_2947,N_2953);
or UO_68 (O_68,N_2962,N_2946);
or UO_69 (O_69,N_2948,N_2974);
and UO_70 (O_70,N_2991,N_2955);
nand UO_71 (O_71,N_2947,N_2949);
nand UO_72 (O_72,N_2980,N_2946);
or UO_73 (O_73,N_2983,N_2942);
or UO_74 (O_74,N_2999,N_2952);
nor UO_75 (O_75,N_2955,N_2974);
nand UO_76 (O_76,N_2962,N_2952);
nand UO_77 (O_77,N_2991,N_2971);
nand UO_78 (O_78,N_2968,N_2942);
and UO_79 (O_79,N_2971,N_2985);
and UO_80 (O_80,N_2966,N_2991);
and UO_81 (O_81,N_2974,N_2997);
or UO_82 (O_82,N_2975,N_2971);
nor UO_83 (O_83,N_2967,N_2998);
or UO_84 (O_84,N_2989,N_2997);
nand UO_85 (O_85,N_2980,N_2992);
nor UO_86 (O_86,N_2995,N_2979);
or UO_87 (O_87,N_2997,N_2981);
and UO_88 (O_88,N_2989,N_2966);
and UO_89 (O_89,N_2968,N_2997);
nor UO_90 (O_90,N_2964,N_2989);
nand UO_91 (O_91,N_2964,N_2979);
and UO_92 (O_92,N_2997,N_2993);
or UO_93 (O_93,N_2950,N_2973);
nor UO_94 (O_94,N_2992,N_2994);
nand UO_95 (O_95,N_2974,N_2976);
nand UO_96 (O_96,N_2994,N_2976);
or UO_97 (O_97,N_2990,N_2991);
or UO_98 (O_98,N_2965,N_2999);
or UO_99 (O_99,N_2949,N_2941);
or UO_100 (O_100,N_2974,N_2973);
and UO_101 (O_101,N_2966,N_2979);
nand UO_102 (O_102,N_2949,N_2946);
nor UO_103 (O_103,N_2959,N_2997);
and UO_104 (O_104,N_2964,N_2956);
xor UO_105 (O_105,N_2968,N_2955);
and UO_106 (O_106,N_2970,N_2981);
or UO_107 (O_107,N_2997,N_2952);
nand UO_108 (O_108,N_2948,N_2989);
nand UO_109 (O_109,N_2954,N_2996);
or UO_110 (O_110,N_2992,N_2976);
nand UO_111 (O_111,N_2976,N_2965);
or UO_112 (O_112,N_2963,N_2993);
and UO_113 (O_113,N_2946,N_2950);
or UO_114 (O_114,N_2963,N_2965);
nor UO_115 (O_115,N_2959,N_2953);
nand UO_116 (O_116,N_2976,N_2986);
nand UO_117 (O_117,N_2992,N_2952);
or UO_118 (O_118,N_2984,N_2999);
nor UO_119 (O_119,N_2975,N_2992);
and UO_120 (O_120,N_2944,N_2945);
nand UO_121 (O_121,N_2979,N_2976);
or UO_122 (O_122,N_2971,N_2987);
nand UO_123 (O_123,N_2964,N_2992);
nor UO_124 (O_124,N_2981,N_2956);
or UO_125 (O_125,N_2983,N_2958);
nor UO_126 (O_126,N_2942,N_2982);
and UO_127 (O_127,N_2980,N_2993);
or UO_128 (O_128,N_2968,N_2994);
and UO_129 (O_129,N_2986,N_2965);
and UO_130 (O_130,N_2944,N_2947);
nand UO_131 (O_131,N_2976,N_2949);
nand UO_132 (O_132,N_2995,N_2959);
nand UO_133 (O_133,N_2954,N_2994);
or UO_134 (O_134,N_2973,N_2981);
nand UO_135 (O_135,N_2977,N_2986);
and UO_136 (O_136,N_2979,N_2959);
nand UO_137 (O_137,N_2948,N_2942);
nor UO_138 (O_138,N_2955,N_2941);
and UO_139 (O_139,N_2989,N_2973);
nor UO_140 (O_140,N_2972,N_2994);
nor UO_141 (O_141,N_2984,N_2961);
or UO_142 (O_142,N_2963,N_2940);
xnor UO_143 (O_143,N_2953,N_2944);
nand UO_144 (O_144,N_2948,N_2975);
nand UO_145 (O_145,N_2953,N_2955);
or UO_146 (O_146,N_2984,N_2992);
or UO_147 (O_147,N_2955,N_2999);
or UO_148 (O_148,N_2954,N_2945);
and UO_149 (O_149,N_2985,N_2961);
and UO_150 (O_150,N_2950,N_2961);
nor UO_151 (O_151,N_2969,N_2992);
nor UO_152 (O_152,N_2983,N_2978);
or UO_153 (O_153,N_2961,N_2986);
nor UO_154 (O_154,N_2943,N_2996);
nor UO_155 (O_155,N_2979,N_2965);
nand UO_156 (O_156,N_2963,N_2981);
or UO_157 (O_157,N_2948,N_2977);
nor UO_158 (O_158,N_2941,N_2982);
nor UO_159 (O_159,N_2954,N_2999);
or UO_160 (O_160,N_2982,N_2946);
nor UO_161 (O_161,N_2994,N_2964);
nand UO_162 (O_162,N_2940,N_2990);
nand UO_163 (O_163,N_2953,N_2951);
and UO_164 (O_164,N_2968,N_2979);
and UO_165 (O_165,N_2999,N_2957);
xnor UO_166 (O_166,N_2983,N_2971);
nor UO_167 (O_167,N_2999,N_2945);
nor UO_168 (O_168,N_2976,N_2960);
or UO_169 (O_169,N_2967,N_2976);
and UO_170 (O_170,N_2951,N_2949);
and UO_171 (O_171,N_2945,N_2953);
xnor UO_172 (O_172,N_2993,N_2966);
or UO_173 (O_173,N_2960,N_2954);
xor UO_174 (O_174,N_2953,N_2940);
or UO_175 (O_175,N_2942,N_2969);
nor UO_176 (O_176,N_2965,N_2954);
or UO_177 (O_177,N_2949,N_2975);
and UO_178 (O_178,N_2961,N_2998);
or UO_179 (O_179,N_2944,N_2983);
and UO_180 (O_180,N_2960,N_2956);
nand UO_181 (O_181,N_2980,N_2958);
nand UO_182 (O_182,N_2940,N_2976);
or UO_183 (O_183,N_2984,N_2949);
or UO_184 (O_184,N_2945,N_2997);
or UO_185 (O_185,N_2982,N_2945);
or UO_186 (O_186,N_2993,N_2971);
nand UO_187 (O_187,N_2962,N_2992);
or UO_188 (O_188,N_2973,N_2958);
and UO_189 (O_189,N_2996,N_2945);
or UO_190 (O_190,N_2967,N_2994);
nand UO_191 (O_191,N_2957,N_2989);
nand UO_192 (O_192,N_2989,N_2976);
or UO_193 (O_193,N_2994,N_2952);
or UO_194 (O_194,N_2984,N_2973);
nand UO_195 (O_195,N_2956,N_2948);
and UO_196 (O_196,N_2961,N_2949);
nor UO_197 (O_197,N_2941,N_2968);
nand UO_198 (O_198,N_2951,N_2982);
and UO_199 (O_199,N_2947,N_2990);
nand UO_200 (O_200,N_2982,N_2965);
nand UO_201 (O_201,N_2951,N_2962);
or UO_202 (O_202,N_2968,N_2953);
nand UO_203 (O_203,N_2994,N_2986);
and UO_204 (O_204,N_2941,N_2999);
nor UO_205 (O_205,N_2990,N_2961);
or UO_206 (O_206,N_2995,N_2966);
xnor UO_207 (O_207,N_2981,N_2986);
and UO_208 (O_208,N_2971,N_2941);
nor UO_209 (O_209,N_2987,N_2961);
nand UO_210 (O_210,N_2996,N_2950);
and UO_211 (O_211,N_2977,N_2987);
and UO_212 (O_212,N_2974,N_2971);
and UO_213 (O_213,N_2998,N_2995);
and UO_214 (O_214,N_2997,N_2971);
or UO_215 (O_215,N_2960,N_2968);
or UO_216 (O_216,N_2951,N_2996);
nand UO_217 (O_217,N_2997,N_2958);
or UO_218 (O_218,N_2964,N_2945);
nand UO_219 (O_219,N_2995,N_2984);
and UO_220 (O_220,N_2996,N_2957);
nor UO_221 (O_221,N_2946,N_2955);
nor UO_222 (O_222,N_2988,N_2960);
or UO_223 (O_223,N_2958,N_2955);
or UO_224 (O_224,N_2973,N_2951);
nand UO_225 (O_225,N_2978,N_2953);
or UO_226 (O_226,N_2996,N_2992);
or UO_227 (O_227,N_2997,N_2953);
and UO_228 (O_228,N_2987,N_2946);
or UO_229 (O_229,N_2956,N_2975);
or UO_230 (O_230,N_2948,N_2957);
and UO_231 (O_231,N_2953,N_2973);
and UO_232 (O_232,N_2969,N_2974);
nand UO_233 (O_233,N_2987,N_2968);
and UO_234 (O_234,N_2997,N_2942);
or UO_235 (O_235,N_2972,N_2946);
or UO_236 (O_236,N_2958,N_2987);
nor UO_237 (O_237,N_2975,N_2957);
nand UO_238 (O_238,N_2979,N_2963);
or UO_239 (O_239,N_2941,N_2964);
nor UO_240 (O_240,N_2983,N_2965);
or UO_241 (O_241,N_2990,N_2986);
nand UO_242 (O_242,N_2959,N_2957);
nor UO_243 (O_243,N_2950,N_2959);
nand UO_244 (O_244,N_2947,N_2956);
or UO_245 (O_245,N_2948,N_2971);
or UO_246 (O_246,N_2953,N_2948);
nand UO_247 (O_247,N_2957,N_2940);
nand UO_248 (O_248,N_2976,N_2973);
nor UO_249 (O_249,N_2976,N_2997);
nor UO_250 (O_250,N_2965,N_2941);
or UO_251 (O_251,N_2945,N_2991);
nor UO_252 (O_252,N_2947,N_2982);
xor UO_253 (O_253,N_2956,N_2944);
nand UO_254 (O_254,N_2992,N_2960);
or UO_255 (O_255,N_2948,N_2946);
and UO_256 (O_256,N_2985,N_2984);
nand UO_257 (O_257,N_2990,N_2941);
nor UO_258 (O_258,N_2962,N_2969);
or UO_259 (O_259,N_2963,N_2960);
or UO_260 (O_260,N_2975,N_2950);
and UO_261 (O_261,N_2984,N_2963);
nor UO_262 (O_262,N_2986,N_2946);
nor UO_263 (O_263,N_2961,N_2975);
or UO_264 (O_264,N_2943,N_2959);
nor UO_265 (O_265,N_2957,N_2965);
or UO_266 (O_266,N_2999,N_2972);
nand UO_267 (O_267,N_2988,N_2971);
nand UO_268 (O_268,N_2977,N_2994);
nor UO_269 (O_269,N_2991,N_2952);
nor UO_270 (O_270,N_2988,N_2946);
nor UO_271 (O_271,N_2951,N_2967);
nor UO_272 (O_272,N_2999,N_2958);
and UO_273 (O_273,N_2991,N_2947);
and UO_274 (O_274,N_2947,N_2973);
nor UO_275 (O_275,N_2951,N_2970);
and UO_276 (O_276,N_2947,N_2972);
and UO_277 (O_277,N_2970,N_2948);
nand UO_278 (O_278,N_2965,N_2970);
and UO_279 (O_279,N_2957,N_2964);
and UO_280 (O_280,N_2981,N_2958);
nand UO_281 (O_281,N_2960,N_2941);
and UO_282 (O_282,N_2956,N_2995);
nand UO_283 (O_283,N_2980,N_2988);
or UO_284 (O_284,N_2992,N_2968);
and UO_285 (O_285,N_2984,N_2980);
nor UO_286 (O_286,N_2997,N_2992);
nand UO_287 (O_287,N_2944,N_2942);
or UO_288 (O_288,N_2991,N_2998);
and UO_289 (O_289,N_2946,N_2959);
and UO_290 (O_290,N_2967,N_2983);
xor UO_291 (O_291,N_2999,N_2992);
or UO_292 (O_292,N_2966,N_2997);
and UO_293 (O_293,N_2948,N_2941);
and UO_294 (O_294,N_2968,N_2980);
nor UO_295 (O_295,N_2965,N_2964);
or UO_296 (O_296,N_2997,N_2969);
and UO_297 (O_297,N_2997,N_2986);
or UO_298 (O_298,N_2957,N_2945);
or UO_299 (O_299,N_2954,N_2980);
or UO_300 (O_300,N_2972,N_2973);
nand UO_301 (O_301,N_2957,N_2991);
nor UO_302 (O_302,N_2944,N_2991);
and UO_303 (O_303,N_2960,N_2990);
nor UO_304 (O_304,N_2962,N_2945);
or UO_305 (O_305,N_2958,N_2965);
xor UO_306 (O_306,N_2946,N_2963);
nor UO_307 (O_307,N_2955,N_2985);
or UO_308 (O_308,N_2979,N_2940);
and UO_309 (O_309,N_2957,N_2988);
nand UO_310 (O_310,N_2967,N_2984);
or UO_311 (O_311,N_2964,N_2952);
and UO_312 (O_312,N_2986,N_2959);
and UO_313 (O_313,N_2972,N_2988);
and UO_314 (O_314,N_2940,N_2967);
and UO_315 (O_315,N_2960,N_2991);
and UO_316 (O_316,N_2940,N_2955);
nand UO_317 (O_317,N_2949,N_2970);
nor UO_318 (O_318,N_2943,N_2994);
and UO_319 (O_319,N_2952,N_2958);
xor UO_320 (O_320,N_2956,N_2945);
nor UO_321 (O_321,N_2941,N_2981);
and UO_322 (O_322,N_2971,N_2968);
or UO_323 (O_323,N_2971,N_2950);
nand UO_324 (O_324,N_2940,N_2980);
nand UO_325 (O_325,N_2994,N_2941);
nor UO_326 (O_326,N_2947,N_2993);
nand UO_327 (O_327,N_2984,N_2953);
or UO_328 (O_328,N_2979,N_2996);
nor UO_329 (O_329,N_2969,N_2973);
or UO_330 (O_330,N_2949,N_2986);
nor UO_331 (O_331,N_2999,N_2949);
or UO_332 (O_332,N_2941,N_2987);
nor UO_333 (O_333,N_2985,N_2954);
or UO_334 (O_334,N_2969,N_2945);
xor UO_335 (O_335,N_2972,N_2985);
or UO_336 (O_336,N_2992,N_2971);
and UO_337 (O_337,N_2967,N_2954);
and UO_338 (O_338,N_2996,N_2969);
nand UO_339 (O_339,N_2979,N_2952);
and UO_340 (O_340,N_2992,N_2954);
or UO_341 (O_341,N_2987,N_2956);
nor UO_342 (O_342,N_2994,N_2957);
and UO_343 (O_343,N_2951,N_2950);
and UO_344 (O_344,N_2973,N_2999);
nand UO_345 (O_345,N_2977,N_2976);
nor UO_346 (O_346,N_2968,N_2970);
nand UO_347 (O_347,N_2975,N_2955);
nand UO_348 (O_348,N_2985,N_2996);
and UO_349 (O_349,N_2950,N_2958);
nor UO_350 (O_350,N_2973,N_2993);
or UO_351 (O_351,N_2944,N_2971);
nand UO_352 (O_352,N_2945,N_2987);
and UO_353 (O_353,N_2951,N_2943);
nand UO_354 (O_354,N_2943,N_2971);
and UO_355 (O_355,N_2962,N_2998);
or UO_356 (O_356,N_2976,N_2991);
xnor UO_357 (O_357,N_2989,N_2991);
nor UO_358 (O_358,N_2976,N_2983);
nor UO_359 (O_359,N_2957,N_2966);
nand UO_360 (O_360,N_2943,N_2998);
nor UO_361 (O_361,N_2974,N_2946);
nor UO_362 (O_362,N_2975,N_2940);
xor UO_363 (O_363,N_2964,N_2988);
nand UO_364 (O_364,N_2961,N_2995);
and UO_365 (O_365,N_2991,N_2958);
nand UO_366 (O_366,N_2994,N_2948);
or UO_367 (O_367,N_2954,N_2941);
nor UO_368 (O_368,N_2942,N_2980);
and UO_369 (O_369,N_2946,N_2992);
nand UO_370 (O_370,N_2974,N_2999);
or UO_371 (O_371,N_2989,N_2943);
xnor UO_372 (O_372,N_2985,N_2952);
or UO_373 (O_373,N_2972,N_2965);
nor UO_374 (O_374,N_2975,N_2965);
nor UO_375 (O_375,N_2948,N_2945);
or UO_376 (O_376,N_2964,N_2961);
or UO_377 (O_377,N_2962,N_2978);
nand UO_378 (O_378,N_2964,N_2940);
or UO_379 (O_379,N_2942,N_2967);
and UO_380 (O_380,N_2952,N_2963);
nand UO_381 (O_381,N_2960,N_2984);
and UO_382 (O_382,N_2982,N_2987);
nor UO_383 (O_383,N_2988,N_2992);
and UO_384 (O_384,N_2994,N_2959);
and UO_385 (O_385,N_2944,N_2996);
nor UO_386 (O_386,N_2988,N_2958);
or UO_387 (O_387,N_2961,N_2970);
and UO_388 (O_388,N_2961,N_2988);
nand UO_389 (O_389,N_2958,N_2945);
or UO_390 (O_390,N_2995,N_2973);
and UO_391 (O_391,N_2941,N_2992);
and UO_392 (O_392,N_2988,N_2967);
or UO_393 (O_393,N_2968,N_2950);
and UO_394 (O_394,N_2979,N_2992);
or UO_395 (O_395,N_2940,N_2989);
nor UO_396 (O_396,N_2974,N_2996);
xor UO_397 (O_397,N_2962,N_2965);
nor UO_398 (O_398,N_2992,N_2943);
nor UO_399 (O_399,N_2987,N_2951);
nand UO_400 (O_400,N_2966,N_2948);
or UO_401 (O_401,N_2963,N_2982);
or UO_402 (O_402,N_2958,N_2984);
nand UO_403 (O_403,N_2993,N_2944);
or UO_404 (O_404,N_2993,N_2967);
and UO_405 (O_405,N_2944,N_2969);
nor UO_406 (O_406,N_2957,N_2973);
nand UO_407 (O_407,N_2996,N_2970);
and UO_408 (O_408,N_2977,N_2968);
nand UO_409 (O_409,N_2960,N_2997);
or UO_410 (O_410,N_2985,N_2947);
or UO_411 (O_411,N_2961,N_2969);
xor UO_412 (O_412,N_2943,N_2977);
nand UO_413 (O_413,N_2959,N_2940);
or UO_414 (O_414,N_2985,N_2941);
nand UO_415 (O_415,N_2988,N_2954);
nand UO_416 (O_416,N_2943,N_2995);
or UO_417 (O_417,N_2960,N_2993);
nor UO_418 (O_418,N_2998,N_2993);
xor UO_419 (O_419,N_2966,N_2952);
and UO_420 (O_420,N_2947,N_2978);
nand UO_421 (O_421,N_2968,N_2943);
nor UO_422 (O_422,N_2951,N_2954);
nand UO_423 (O_423,N_2949,N_2965);
xor UO_424 (O_424,N_2961,N_2955);
and UO_425 (O_425,N_2991,N_2987);
nand UO_426 (O_426,N_2969,N_2966);
nand UO_427 (O_427,N_2979,N_2978);
nor UO_428 (O_428,N_2944,N_2999);
and UO_429 (O_429,N_2957,N_2983);
nand UO_430 (O_430,N_2992,N_2953);
nand UO_431 (O_431,N_2945,N_2976);
and UO_432 (O_432,N_2946,N_2977);
nor UO_433 (O_433,N_2958,N_2947);
nand UO_434 (O_434,N_2975,N_2960);
and UO_435 (O_435,N_2960,N_2961);
and UO_436 (O_436,N_2953,N_2969);
nor UO_437 (O_437,N_2982,N_2958);
nand UO_438 (O_438,N_2943,N_2957);
or UO_439 (O_439,N_2956,N_2959);
and UO_440 (O_440,N_2950,N_2948);
or UO_441 (O_441,N_2945,N_2943);
xnor UO_442 (O_442,N_2984,N_2974);
and UO_443 (O_443,N_2989,N_2996);
and UO_444 (O_444,N_2957,N_2942);
and UO_445 (O_445,N_2985,N_2977);
or UO_446 (O_446,N_2999,N_2997);
nor UO_447 (O_447,N_2985,N_2960);
and UO_448 (O_448,N_2950,N_2990);
or UO_449 (O_449,N_2970,N_2977);
nand UO_450 (O_450,N_2993,N_2999);
and UO_451 (O_451,N_2999,N_2969);
or UO_452 (O_452,N_2978,N_2987);
nand UO_453 (O_453,N_2977,N_2941);
or UO_454 (O_454,N_2979,N_2985);
and UO_455 (O_455,N_2973,N_2977);
nand UO_456 (O_456,N_2990,N_2993);
and UO_457 (O_457,N_2989,N_2993);
nand UO_458 (O_458,N_2944,N_2981);
or UO_459 (O_459,N_2961,N_2994);
and UO_460 (O_460,N_2953,N_2989);
and UO_461 (O_461,N_2974,N_2949);
and UO_462 (O_462,N_2953,N_2982);
and UO_463 (O_463,N_2999,N_2987);
or UO_464 (O_464,N_2959,N_2944);
and UO_465 (O_465,N_2974,N_2982);
or UO_466 (O_466,N_2980,N_2943);
nor UO_467 (O_467,N_2987,N_2983);
nor UO_468 (O_468,N_2977,N_2963);
nand UO_469 (O_469,N_2955,N_2981);
nand UO_470 (O_470,N_2942,N_2975);
xnor UO_471 (O_471,N_2978,N_2975);
or UO_472 (O_472,N_2944,N_2955);
and UO_473 (O_473,N_2945,N_2993);
or UO_474 (O_474,N_2979,N_2967);
nand UO_475 (O_475,N_2989,N_2945);
and UO_476 (O_476,N_2996,N_2976);
nand UO_477 (O_477,N_2974,N_2944);
nor UO_478 (O_478,N_2985,N_2980);
and UO_479 (O_479,N_2997,N_2998);
and UO_480 (O_480,N_2984,N_2987);
and UO_481 (O_481,N_2945,N_2985);
and UO_482 (O_482,N_2970,N_2947);
or UO_483 (O_483,N_2959,N_2991);
and UO_484 (O_484,N_2955,N_2942);
or UO_485 (O_485,N_2986,N_2995);
and UO_486 (O_486,N_2972,N_2983);
and UO_487 (O_487,N_2941,N_2975);
and UO_488 (O_488,N_2998,N_2941);
or UO_489 (O_489,N_2973,N_2956);
and UO_490 (O_490,N_2980,N_2999);
nor UO_491 (O_491,N_2953,N_2990);
nor UO_492 (O_492,N_2961,N_2947);
nor UO_493 (O_493,N_2946,N_2952);
nand UO_494 (O_494,N_2975,N_2962);
and UO_495 (O_495,N_2994,N_2974);
nor UO_496 (O_496,N_2986,N_2963);
nand UO_497 (O_497,N_2942,N_2965);
and UO_498 (O_498,N_2986,N_2998);
nor UO_499 (O_499,N_2986,N_2985);
endmodule